module basic_5000_50000_5000_25_levels_10xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999,N_30000,N_30001,N_30002,N_30003,N_30004,N_30005,N_30006,N_30007,N_30008,N_30009,N_30010,N_30011,N_30012,N_30013,N_30014,N_30015,N_30016,N_30017,N_30018,N_30019,N_30020,N_30021,N_30022,N_30023,N_30024,N_30025,N_30026,N_30027,N_30028,N_30029,N_30030,N_30031,N_30032,N_30033,N_30034,N_30035,N_30036,N_30037,N_30038,N_30039,N_30040,N_30041,N_30042,N_30043,N_30044,N_30045,N_30046,N_30047,N_30048,N_30049,N_30050,N_30051,N_30052,N_30053,N_30054,N_30055,N_30056,N_30057,N_30058,N_30059,N_30060,N_30061,N_30062,N_30063,N_30064,N_30065,N_30066,N_30067,N_30068,N_30069,N_30070,N_30071,N_30072,N_30073,N_30074,N_30075,N_30076,N_30077,N_30078,N_30079,N_30080,N_30081,N_30082,N_30083,N_30084,N_30085,N_30086,N_30087,N_30088,N_30089,N_30090,N_30091,N_30092,N_30093,N_30094,N_30095,N_30096,N_30097,N_30098,N_30099,N_30100,N_30101,N_30102,N_30103,N_30104,N_30105,N_30106,N_30107,N_30108,N_30109,N_30110,N_30111,N_30112,N_30113,N_30114,N_30115,N_30116,N_30117,N_30118,N_30119,N_30120,N_30121,N_30122,N_30123,N_30124,N_30125,N_30126,N_30127,N_30128,N_30129,N_30130,N_30131,N_30132,N_30133,N_30134,N_30135,N_30136,N_30137,N_30138,N_30139,N_30140,N_30141,N_30142,N_30143,N_30144,N_30145,N_30146,N_30147,N_30148,N_30149,N_30150,N_30151,N_30152,N_30153,N_30154,N_30155,N_30156,N_30157,N_30158,N_30159,N_30160,N_30161,N_30162,N_30163,N_30164,N_30165,N_30166,N_30167,N_30168,N_30169,N_30170,N_30171,N_30172,N_30173,N_30174,N_30175,N_30176,N_30177,N_30178,N_30179,N_30180,N_30181,N_30182,N_30183,N_30184,N_30185,N_30186,N_30187,N_30188,N_30189,N_30190,N_30191,N_30192,N_30193,N_30194,N_30195,N_30196,N_30197,N_30198,N_30199,N_30200,N_30201,N_30202,N_30203,N_30204,N_30205,N_30206,N_30207,N_30208,N_30209,N_30210,N_30211,N_30212,N_30213,N_30214,N_30215,N_30216,N_30217,N_30218,N_30219,N_30220,N_30221,N_30222,N_30223,N_30224,N_30225,N_30226,N_30227,N_30228,N_30229,N_30230,N_30231,N_30232,N_30233,N_30234,N_30235,N_30236,N_30237,N_30238,N_30239,N_30240,N_30241,N_30242,N_30243,N_30244,N_30245,N_30246,N_30247,N_30248,N_30249,N_30250,N_30251,N_30252,N_30253,N_30254,N_30255,N_30256,N_30257,N_30258,N_30259,N_30260,N_30261,N_30262,N_30263,N_30264,N_30265,N_30266,N_30267,N_30268,N_30269,N_30270,N_30271,N_30272,N_30273,N_30274,N_30275,N_30276,N_30277,N_30278,N_30279,N_30280,N_30281,N_30282,N_30283,N_30284,N_30285,N_30286,N_30287,N_30288,N_30289,N_30290,N_30291,N_30292,N_30293,N_30294,N_30295,N_30296,N_30297,N_30298,N_30299,N_30300,N_30301,N_30302,N_30303,N_30304,N_30305,N_30306,N_30307,N_30308,N_30309,N_30310,N_30311,N_30312,N_30313,N_30314,N_30315,N_30316,N_30317,N_30318,N_30319,N_30320,N_30321,N_30322,N_30323,N_30324,N_30325,N_30326,N_30327,N_30328,N_30329,N_30330,N_30331,N_30332,N_30333,N_30334,N_30335,N_30336,N_30337,N_30338,N_30339,N_30340,N_30341,N_30342,N_30343,N_30344,N_30345,N_30346,N_30347,N_30348,N_30349,N_30350,N_30351,N_30352,N_30353,N_30354,N_30355,N_30356,N_30357,N_30358,N_30359,N_30360,N_30361,N_30362,N_30363,N_30364,N_30365,N_30366,N_30367,N_30368,N_30369,N_30370,N_30371,N_30372,N_30373,N_30374,N_30375,N_30376,N_30377,N_30378,N_30379,N_30380,N_30381,N_30382,N_30383,N_30384,N_30385,N_30386,N_30387,N_30388,N_30389,N_30390,N_30391,N_30392,N_30393,N_30394,N_30395,N_30396,N_30397,N_30398,N_30399,N_30400,N_30401,N_30402,N_30403,N_30404,N_30405,N_30406,N_30407,N_30408,N_30409,N_30410,N_30411,N_30412,N_30413,N_30414,N_30415,N_30416,N_30417,N_30418,N_30419,N_30420,N_30421,N_30422,N_30423,N_30424,N_30425,N_30426,N_30427,N_30428,N_30429,N_30430,N_30431,N_30432,N_30433,N_30434,N_30435,N_30436,N_30437,N_30438,N_30439,N_30440,N_30441,N_30442,N_30443,N_30444,N_30445,N_30446,N_30447,N_30448,N_30449,N_30450,N_30451,N_30452,N_30453,N_30454,N_30455,N_30456,N_30457,N_30458,N_30459,N_30460,N_30461,N_30462,N_30463,N_30464,N_30465,N_30466,N_30467,N_30468,N_30469,N_30470,N_30471,N_30472,N_30473,N_30474,N_30475,N_30476,N_30477,N_30478,N_30479,N_30480,N_30481,N_30482,N_30483,N_30484,N_30485,N_30486,N_30487,N_30488,N_30489,N_30490,N_30491,N_30492,N_30493,N_30494,N_30495,N_30496,N_30497,N_30498,N_30499,N_30500,N_30501,N_30502,N_30503,N_30504,N_30505,N_30506,N_30507,N_30508,N_30509,N_30510,N_30511,N_30512,N_30513,N_30514,N_30515,N_30516,N_30517,N_30518,N_30519,N_30520,N_30521,N_30522,N_30523,N_30524,N_30525,N_30526,N_30527,N_30528,N_30529,N_30530,N_30531,N_30532,N_30533,N_30534,N_30535,N_30536,N_30537,N_30538,N_30539,N_30540,N_30541,N_30542,N_30543,N_30544,N_30545,N_30546,N_30547,N_30548,N_30549,N_30550,N_30551,N_30552,N_30553,N_30554,N_30555,N_30556,N_30557,N_30558,N_30559,N_30560,N_30561,N_30562,N_30563,N_30564,N_30565,N_30566,N_30567,N_30568,N_30569,N_30570,N_30571,N_30572,N_30573,N_30574,N_30575,N_30576,N_30577,N_30578,N_30579,N_30580,N_30581,N_30582,N_30583,N_30584,N_30585,N_30586,N_30587,N_30588,N_30589,N_30590,N_30591,N_30592,N_30593,N_30594,N_30595,N_30596,N_30597,N_30598,N_30599,N_30600,N_30601,N_30602,N_30603,N_30604,N_30605,N_30606,N_30607,N_30608,N_30609,N_30610,N_30611,N_30612,N_30613,N_30614,N_30615,N_30616,N_30617,N_30618,N_30619,N_30620,N_30621,N_30622,N_30623,N_30624,N_30625,N_30626,N_30627,N_30628,N_30629,N_30630,N_30631,N_30632,N_30633,N_30634,N_30635,N_30636,N_30637,N_30638,N_30639,N_30640,N_30641,N_30642,N_30643,N_30644,N_30645,N_30646,N_30647,N_30648,N_30649,N_30650,N_30651,N_30652,N_30653,N_30654,N_30655,N_30656,N_30657,N_30658,N_30659,N_30660,N_30661,N_30662,N_30663,N_30664,N_30665,N_30666,N_30667,N_30668,N_30669,N_30670,N_30671,N_30672,N_30673,N_30674,N_30675,N_30676,N_30677,N_30678,N_30679,N_30680,N_30681,N_30682,N_30683,N_30684,N_30685,N_30686,N_30687,N_30688,N_30689,N_30690,N_30691,N_30692,N_30693,N_30694,N_30695,N_30696,N_30697,N_30698,N_30699,N_30700,N_30701,N_30702,N_30703,N_30704,N_30705,N_30706,N_30707,N_30708,N_30709,N_30710,N_30711,N_30712,N_30713,N_30714,N_30715,N_30716,N_30717,N_30718,N_30719,N_30720,N_30721,N_30722,N_30723,N_30724,N_30725,N_30726,N_30727,N_30728,N_30729,N_30730,N_30731,N_30732,N_30733,N_30734,N_30735,N_30736,N_30737,N_30738,N_30739,N_30740,N_30741,N_30742,N_30743,N_30744,N_30745,N_30746,N_30747,N_30748,N_30749,N_30750,N_30751,N_30752,N_30753,N_30754,N_30755,N_30756,N_30757,N_30758,N_30759,N_30760,N_30761,N_30762,N_30763,N_30764,N_30765,N_30766,N_30767,N_30768,N_30769,N_30770,N_30771,N_30772,N_30773,N_30774,N_30775,N_30776,N_30777,N_30778,N_30779,N_30780,N_30781,N_30782,N_30783,N_30784,N_30785,N_30786,N_30787,N_30788,N_30789,N_30790,N_30791,N_30792,N_30793,N_30794,N_30795,N_30796,N_30797,N_30798,N_30799,N_30800,N_30801,N_30802,N_30803,N_30804,N_30805,N_30806,N_30807,N_30808,N_30809,N_30810,N_30811,N_30812,N_30813,N_30814,N_30815,N_30816,N_30817,N_30818,N_30819,N_30820,N_30821,N_30822,N_30823,N_30824,N_30825,N_30826,N_30827,N_30828,N_30829,N_30830,N_30831,N_30832,N_30833,N_30834,N_30835,N_30836,N_30837,N_30838,N_30839,N_30840,N_30841,N_30842,N_30843,N_30844,N_30845,N_30846,N_30847,N_30848,N_30849,N_30850,N_30851,N_30852,N_30853,N_30854,N_30855,N_30856,N_30857,N_30858,N_30859,N_30860,N_30861,N_30862,N_30863,N_30864,N_30865,N_30866,N_30867,N_30868,N_30869,N_30870,N_30871,N_30872,N_30873,N_30874,N_30875,N_30876,N_30877,N_30878,N_30879,N_30880,N_30881,N_30882,N_30883,N_30884,N_30885,N_30886,N_30887,N_30888,N_30889,N_30890,N_30891,N_30892,N_30893,N_30894,N_30895,N_30896,N_30897,N_30898,N_30899,N_30900,N_30901,N_30902,N_30903,N_30904,N_30905,N_30906,N_30907,N_30908,N_30909,N_30910,N_30911,N_30912,N_30913,N_30914,N_30915,N_30916,N_30917,N_30918,N_30919,N_30920,N_30921,N_30922,N_30923,N_30924,N_30925,N_30926,N_30927,N_30928,N_30929,N_30930,N_30931,N_30932,N_30933,N_30934,N_30935,N_30936,N_30937,N_30938,N_30939,N_30940,N_30941,N_30942,N_30943,N_30944,N_30945,N_30946,N_30947,N_30948,N_30949,N_30950,N_30951,N_30952,N_30953,N_30954,N_30955,N_30956,N_30957,N_30958,N_30959,N_30960,N_30961,N_30962,N_30963,N_30964,N_30965,N_30966,N_30967,N_30968,N_30969,N_30970,N_30971,N_30972,N_30973,N_30974,N_30975,N_30976,N_30977,N_30978,N_30979,N_30980,N_30981,N_30982,N_30983,N_30984,N_30985,N_30986,N_30987,N_30988,N_30989,N_30990,N_30991,N_30992,N_30993,N_30994,N_30995,N_30996,N_30997,N_30998,N_30999,N_31000,N_31001,N_31002,N_31003,N_31004,N_31005,N_31006,N_31007,N_31008,N_31009,N_31010,N_31011,N_31012,N_31013,N_31014,N_31015,N_31016,N_31017,N_31018,N_31019,N_31020,N_31021,N_31022,N_31023,N_31024,N_31025,N_31026,N_31027,N_31028,N_31029,N_31030,N_31031,N_31032,N_31033,N_31034,N_31035,N_31036,N_31037,N_31038,N_31039,N_31040,N_31041,N_31042,N_31043,N_31044,N_31045,N_31046,N_31047,N_31048,N_31049,N_31050,N_31051,N_31052,N_31053,N_31054,N_31055,N_31056,N_31057,N_31058,N_31059,N_31060,N_31061,N_31062,N_31063,N_31064,N_31065,N_31066,N_31067,N_31068,N_31069,N_31070,N_31071,N_31072,N_31073,N_31074,N_31075,N_31076,N_31077,N_31078,N_31079,N_31080,N_31081,N_31082,N_31083,N_31084,N_31085,N_31086,N_31087,N_31088,N_31089,N_31090,N_31091,N_31092,N_31093,N_31094,N_31095,N_31096,N_31097,N_31098,N_31099,N_31100,N_31101,N_31102,N_31103,N_31104,N_31105,N_31106,N_31107,N_31108,N_31109,N_31110,N_31111,N_31112,N_31113,N_31114,N_31115,N_31116,N_31117,N_31118,N_31119,N_31120,N_31121,N_31122,N_31123,N_31124,N_31125,N_31126,N_31127,N_31128,N_31129,N_31130,N_31131,N_31132,N_31133,N_31134,N_31135,N_31136,N_31137,N_31138,N_31139,N_31140,N_31141,N_31142,N_31143,N_31144,N_31145,N_31146,N_31147,N_31148,N_31149,N_31150,N_31151,N_31152,N_31153,N_31154,N_31155,N_31156,N_31157,N_31158,N_31159,N_31160,N_31161,N_31162,N_31163,N_31164,N_31165,N_31166,N_31167,N_31168,N_31169,N_31170,N_31171,N_31172,N_31173,N_31174,N_31175,N_31176,N_31177,N_31178,N_31179,N_31180,N_31181,N_31182,N_31183,N_31184,N_31185,N_31186,N_31187,N_31188,N_31189,N_31190,N_31191,N_31192,N_31193,N_31194,N_31195,N_31196,N_31197,N_31198,N_31199,N_31200,N_31201,N_31202,N_31203,N_31204,N_31205,N_31206,N_31207,N_31208,N_31209,N_31210,N_31211,N_31212,N_31213,N_31214,N_31215,N_31216,N_31217,N_31218,N_31219,N_31220,N_31221,N_31222,N_31223,N_31224,N_31225,N_31226,N_31227,N_31228,N_31229,N_31230,N_31231,N_31232,N_31233,N_31234,N_31235,N_31236,N_31237,N_31238,N_31239,N_31240,N_31241,N_31242,N_31243,N_31244,N_31245,N_31246,N_31247,N_31248,N_31249,N_31250,N_31251,N_31252,N_31253,N_31254,N_31255,N_31256,N_31257,N_31258,N_31259,N_31260,N_31261,N_31262,N_31263,N_31264,N_31265,N_31266,N_31267,N_31268,N_31269,N_31270,N_31271,N_31272,N_31273,N_31274,N_31275,N_31276,N_31277,N_31278,N_31279,N_31280,N_31281,N_31282,N_31283,N_31284,N_31285,N_31286,N_31287,N_31288,N_31289,N_31290,N_31291,N_31292,N_31293,N_31294,N_31295,N_31296,N_31297,N_31298,N_31299,N_31300,N_31301,N_31302,N_31303,N_31304,N_31305,N_31306,N_31307,N_31308,N_31309,N_31310,N_31311,N_31312,N_31313,N_31314,N_31315,N_31316,N_31317,N_31318,N_31319,N_31320,N_31321,N_31322,N_31323,N_31324,N_31325,N_31326,N_31327,N_31328,N_31329,N_31330,N_31331,N_31332,N_31333,N_31334,N_31335,N_31336,N_31337,N_31338,N_31339,N_31340,N_31341,N_31342,N_31343,N_31344,N_31345,N_31346,N_31347,N_31348,N_31349,N_31350,N_31351,N_31352,N_31353,N_31354,N_31355,N_31356,N_31357,N_31358,N_31359,N_31360,N_31361,N_31362,N_31363,N_31364,N_31365,N_31366,N_31367,N_31368,N_31369,N_31370,N_31371,N_31372,N_31373,N_31374,N_31375,N_31376,N_31377,N_31378,N_31379,N_31380,N_31381,N_31382,N_31383,N_31384,N_31385,N_31386,N_31387,N_31388,N_31389,N_31390,N_31391,N_31392,N_31393,N_31394,N_31395,N_31396,N_31397,N_31398,N_31399,N_31400,N_31401,N_31402,N_31403,N_31404,N_31405,N_31406,N_31407,N_31408,N_31409,N_31410,N_31411,N_31412,N_31413,N_31414,N_31415,N_31416,N_31417,N_31418,N_31419,N_31420,N_31421,N_31422,N_31423,N_31424,N_31425,N_31426,N_31427,N_31428,N_31429,N_31430,N_31431,N_31432,N_31433,N_31434,N_31435,N_31436,N_31437,N_31438,N_31439,N_31440,N_31441,N_31442,N_31443,N_31444,N_31445,N_31446,N_31447,N_31448,N_31449,N_31450,N_31451,N_31452,N_31453,N_31454,N_31455,N_31456,N_31457,N_31458,N_31459,N_31460,N_31461,N_31462,N_31463,N_31464,N_31465,N_31466,N_31467,N_31468,N_31469,N_31470,N_31471,N_31472,N_31473,N_31474,N_31475,N_31476,N_31477,N_31478,N_31479,N_31480,N_31481,N_31482,N_31483,N_31484,N_31485,N_31486,N_31487,N_31488,N_31489,N_31490,N_31491,N_31492,N_31493,N_31494,N_31495,N_31496,N_31497,N_31498,N_31499,N_31500,N_31501,N_31502,N_31503,N_31504,N_31505,N_31506,N_31507,N_31508,N_31509,N_31510,N_31511,N_31512,N_31513,N_31514,N_31515,N_31516,N_31517,N_31518,N_31519,N_31520,N_31521,N_31522,N_31523,N_31524,N_31525,N_31526,N_31527,N_31528,N_31529,N_31530,N_31531,N_31532,N_31533,N_31534,N_31535,N_31536,N_31537,N_31538,N_31539,N_31540,N_31541,N_31542,N_31543,N_31544,N_31545,N_31546,N_31547,N_31548,N_31549,N_31550,N_31551,N_31552,N_31553,N_31554,N_31555,N_31556,N_31557,N_31558,N_31559,N_31560,N_31561,N_31562,N_31563,N_31564,N_31565,N_31566,N_31567,N_31568,N_31569,N_31570,N_31571,N_31572,N_31573,N_31574,N_31575,N_31576,N_31577,N_31578,N_31579,N_31580,N_31581,N_31582,N_31583,N_31584,N_31585,N_31586,N_31587,N_31588,N_31589,N_31590,N_31591,N_31592,N_31593,N_31594,N_31595,N_31596,N_31597,N_31598,N_31599,N_31600,N_31601,N_31602,N_31603,N_31604,N_31605,N_31606,N_31607,N_31608,N_31609,N_31610,N_31611,N_31612,N_31613,N_31614,N_31615,N_31616,N_31617,N_31618,N_31619,N_31620,N_31621,N_31622,N_31623,N_31624,N_31625,N_31626,N_31627,N_31628,N_31629,N_31630,N_31631,N_31632,N_31633,N_31634,N_31635,N_31636,N_31637,N_31638,N_31639,N_31640,N_31641,N_31642,N_31643,N_31644,N_31645,N_31646,N_31647,N_31648,N_31649,N_31650,N_31651,N_31652,N_31653,N_31654,N_31655,N_31656,N_31657,N_31658,N_31659,N_31660,N_31661,N_31662,N_31663,N_31664,N_31665,N_31666,N_31667,N_31668,N_31669,N_31670,N_31671,N_31672,N_31673,N_31674,N_31675,N_31676,N_31677,N_31678,N_31679,N_31680,N_31681,N_31682,N_31683,N_31684,N_31685,N_31686,N_31687,N_31688,N_31689,N_31690,N_31691,N_31692,N_31693,N_31694,N_31695,N_31696,N_31697,N_31698,N_31699,N_31700,N_31701,N_31702,N_31703,N_31704,N_31705,N_31706,N_31707,N_31708,N_31709,N_31710,N_31711,N_31712,N_31713,N_31714,N_31715,N_31716,N_31717,N_31718,N_31719,N_31720,N_31721,N_31722,N_31723,N_31724,N_31725,N_31726,N_31727,N_31728,N_31729,N_31730,N_31731,N_31732,N_31733,N_31734,N_31735,N_31736,N_31737,N_31738,N_31739,N_31740,N_31741,N_31742,N_31743,N_31744,N_31745,N_31746,N_31747,N_31748,N_31749,N_31750,N_31751,N_31752,N_31753,N_31754,N_31755,N_31756,N_31757,N_31758,N_31759,N_31760,N_31761,N_31762,N_31763,N_31764,N_31765,N_31766,N_31767,N_31768,N_31769,N_31770,N_31771,N_31772,N_31773,N_31774,N_31775,N_31776,N_31777,N_31778,N_31779,N_31780,N_31781,N_31782,N_31783,N_31784,N_31785,N_31786,N_31787,N_31788,N_31789,N_31790,N_31791,N_31792,N_31793,N_31794,N_31795,N_31796,N_31797,N_31798,N_31799,N_31800,N_31801,N_31802,N_31803,N_31804,N_31805,N_31806,N_31807,N_31808,N_31809,N_31810,N_31811,N_31812,N_31813,N_31814,N_31815,N_31816,N_31817,N_31818,N_31819,N_31820,N_31821,N_31822,N_31823,N_31824,N_31825,N_31826,N_31827,N_31828,N_31829,N_31830,N_31831,N_31832,N_31833,N_31834,N_31835,N_31836,N_31837,N_31838,N_31839,N_31840,N_31841,N_31842,N_31843,N_31844,N_31845,N_31846,N_31847,N_31848,N_31849,N_31850,N_31851,N_31852,N_31853,N_31854,N_31855,N_31856,N_31857,N_31858,N_31859,N_31860,N_31861,N_31862,N_31863,N_31864,N_31865,N_31866,N_31867,N_31868,N_31869,N_31870,N_31871,N_31872,N_31873,N_31874,N_31875,N_31876,N_31877,N_31878,N_31879,N_31880,N_31881,N_31882,N_31883,N_31884,N_31885,N_31886,N_31887,N_31888,N_31889,N_31890,N_31891,N_31892,N_31893,N_31894,N_31895,N_31896,N_31897,N_31898,N_31899,N_31900,N_31901,N_31902,N_31903,N_31904,N_31905,N_31906,N_31907,N_31908,N_31909,N_31910,N_31911,N_31912,N_31913,N_31914,N_31915,N_31916,N_31917,N_31918,N_31919,N_31920,N_31921,N_31922,N_31923,N_31924,N_31925,N_31926,N_31927,N_31928,N_31929,N_31930,N_31931,N_31932,N_31933,N_31934,N_31935,N_31936,N_31937,N_31938,N_31939,N_31940,N_31941,N_31942,N_31943,N_31944,N_31945,N_31946,N_31947,N_31948,N_31949,N_31950,N_31951,N_31952,N_31953,N_31954,N_31955,N_31956,N_31957,N_31958,N_31959,N_31960,N_31961,N_31962,N_31963,N_31964,N_31965,N_31966,N_31967,N_31968,N_31969,N_31970,N_31971,N_31972,N_31973,N_31974,N_31975,N_31976,N_31977,N_31978,N_31979,N_31980,N_31981,N_31982,N_31983,N_31984,N_31985,N_31986,N_31987,N_31988,N_31989,N_31990,N_31991,N_31992,N_31993,N_31994,N_31995,N_31996,N_31997,N_31998,N_31999,N_32000,N_32001,N_32002,N_32003,N_32004,N_32005,N_32006,N_32007,N_32008,N_32009,N_32010,N_32011,N_32012,N_32013,N_32014,N_32015,N_32016,N_32017,N_32018,N_32019,N_32020,N_32021,N_32022,N_32023,N_32024,N_32025,N_32026,N_32027,N_32028,N_32029,N_32030,N_32031,N_32032,N_32033,N_32034,N_32035,N_32036,N_32037,N_32038,N_32039,N_32040,N_32041,N_32042,N_32043,N_32044,N_32045,N_32046,N_32047,N_32048,N_32049,N_32050,N_32051,N_32052,N_32053,N_32054,N_32055,N_32056,N_32057,N_32058,N_32059,N_32060,N_32061,N_32062,N_32063,N_32064,N_32065,N_32066,N_32067,N_32068,N_32069,N_32070,N_32071,N_32072,N_32073,N_32074,N_32075,N_32076,N_32077,N_32078,N_32079,N_32080,N_32081,N_32082,N_32083,N_32084,N_32085,N_32086,N_32087,N_32088,N_32089,N_32090,N_32091,N_32092,N_32093,N_32094,N_32095,N_32096,N_32097,N_32098,N_32099,N_32100,N_32101,N_32102,N_32103,N_32104,N_32105,N_32106,N_32107,N_32108,N_32109,N_32110,N_32111,N_32112,N_32113,N_32114,N_32115,N_32116,N_32117,N_32118,N_32119,N_32120,N_32121,N_32122,N_32123,N_32124,N_32125,N_32126,N_32127,N_32128,N_32129,N_32130,N_32131,N_32132,N_32133,N_32134,N_32135,N_32136,N_32137,N_32138,N_32139,N_32140,N_32141,N_32142,N_32143,N_32144,N_32145,N_32146,N_32147,N_32148,N_32149,N_32150,N_32151,N_32152,N_32153,N_32154,N_32155,N_32156,N_32157,N_32158,N_32159,N_32160,N_32161,N_32162,N_32163,N_32164,N_32165,N_32166,N_32167,N_32168,N_32169,N_32170,N_32171,N_32172,N_32173,N_32174,N_32175,N_32176,N_32177,N_32178,N_32179,N_32180,N_32181,N_32182,N_32183,N_32184,N_32185,N_32186,N_32187,N_32188,N_32189,N_32190,N_32191,N_32192,N_32193,N_32194,N_32195,N_32196,N_32197,N_32198,N_32199,N_32200,N_32201,N_32202,N_32203,N_32204,N_32205,N_32206,N_32207,N_32208,N_32209,N_32210,N_32211,N_32212,N_32213,N_32214,N_32215,N_32216,N_32217,N_32218,N_32219,N_32220,N_32221,N_32222,N_32223,N_32224,N_32225,N_32226,N_32227,N_32228,N_32229,N_32230,N_32231,N_32232,N_32233,N_32234,N_32235,N_32236,N_32237,N_32238,N_32239,N_32240,N_32241,N_32242,N_32243,N_32244,N_32245,N_32246,N_32247,N_32248,N_32249,N_32250,N_32251,N_32252,N_32253,N_32254,N_32255,N_32256,N_32257,N_32258,N_32259,N_32260,N_32261,N_32262,N_32263,N_32264,N_32265,N_32266,N_32267,N_32268,N_32269,N_32270,N_32271,N_32272,N_32273,N_32274,N_32275,N_32276,N_32277,N_32278,N_32279,N_32280,N_32281,N_32282,N_32283,N_32284,N_32285,N_32286,N_32287,N_32288,N_32289,N_32290,N_32291,N_32292,N_32293,N_32294,N_32295,N_32296,N_32297,N_32298,N_32299,N_32300,N_32301,N_32302,N_32303,N_32304,N_32305,N_32306,N_32307,N_32308,N_32309,N_32310,N_32311,N_32312,N_32313,N_32314,N_32315,N_32316,N_32317,N_32318,N_32319,N_32320,N_32321,N_32322,N_32323,N_32324,N_32325,N_32326,N_32327,N_32328,N_32329,N_32330,N_32331,N_32332,N_32333,N_32334,N_32335,N_32336,N_32337,N_32338,N_32339,N_32340,N_32341,N_32342,N_32343,N_32344,N_32345,N_32346,N_32347,N_32348,N_32349,N_32350,N_32351,N_32352,N_32353,N_32354,N_32355,N_32356,N_32357,N_32358,N_32359,N_32360,N_32361,N_32362,N_32363,N_32364,N_32365,N_32366,N_32367,N_32368,N_32369,N_32370,N_32371,N_32372,N_32373,N_32374,N_32375,N_32376,N_32377,N_32378,N_32379,N_32380,N_32381,N_32382,N_32383,N_32384,N_32385,N_32386,N_32387,N_32388,N_32389,N_32390,N_32391,N_32392,N_32393,N_32394,N_32395,N_32396,N_32397,N_32398,N_32399,N_32400,N_32401,N_32402,N_32403,N_32404,N_32405,N_32406,N_32407,N_32408,N_32409,N_32410,N_32411,N_32412,N_32413,N_32414,N_32415,N_32416,N_32417,N_32418,N_32419,N_32420,N_32421,N_32422,N_32423,N_32424,N_32425,N_32426,N_32427,N_32428,N_32429,N_32430,N_32431,N_32432,N_32433,N_32434,N_32435,N_32436,N_32437,N_32438,N_32439,N_32440,N_32441,N_32442,N_32443,N_32444,N_32445,N_32446,N_32447,N_32448,N_32449,N_32450,N_32451,N_32452,N_32453,N_32454,N_32455,N_32456,N_32457,N_32458,N_32459,N_32460,N_32461,N_32462,N_32463,N_32464,N_32465,N_32466,N_32467,N_32468,N_32469,N_32470,N_32471,N_32472,N_32473,N_32474,N_32475,N_32476,N_32477,N_32478,N_32479,N_32480,N_32481,N_32482,N_32483,N_32484,N_32485,N_32486,N_32487,N_32488,N_32489,N_32490,N_32491,N_32492,N_32493,N_32494,N_32495,N_32496,N_32497,N_32498,N_32499,N_32500,N_32501,N_32502,N_32503,N_32504,N_32505,N_32506,N_32507,N_32508,N_32509,N_32510,N_32511,N_32512,N_32513,N_32514,N_32515,N_32516,N_32517,N_32518,N_32519,N_32520,N_32521,N_32522,N_32523,N_32524,N_32525,N_32526,N_32527,N_32528,N_32529,N_32530,N_32531,N_32532,N_32533,N_32534,N_32535,N_32536,N_32537,N_32538,N_32539,N_32540,N_32541,N_32542,N_32543,N_32544,N_32545,N_32546,N_32547,N_32548,N_32549,N_32550,N_32551,N_32552,N_32553,N_32554,N_32555,N_32556,N_32557,N_32558,N_32559,N_32560,N_32561,N_32562,N_32563,N_32564,N_32565,N_32566,N_32567,N_32568,N_32569,N_32570,N_32571,N_32572,N_32573,N_32574,N_32575,N_32576,N_32577,N_32578,N_32579,N_32580,N_32581,N_32582,N_32583,N_32584,N_32585,N_32586,N_32587,N_32588,N_32589,N_32590,N_32591,N_32592,N_32593,N_32594,N_32595,N_32596,N_32597,N_32598,N_32599,N_32600,N_32601,N_32602,N_32603,N_32604,N_32605,N_32606,N_32607,N_32608,N_32609,N_32610,N_32611,N_32612,N_32613,N_32614,N_32615,N_32616,N_32617,N_32618,N_32619,N_32620,N_32621,N_32622,N_32623,N_32624,N_32625,N_32626,N_32627,N_32628,N_32629,N_32630,N_32631,N_32632,N_32633,N_32634,N_32635,N_32636,N_32637,N_32638,N_32639,N_32640,N_32641,N_32642,N_32643,N_32644,N_32645,N_32646,N_32647,N_32648,N_32649,N_32650,N_32651,N_32652,N_32653,N_32654,N_32655,N_32656,N_32657,N_32658,N_32659,N_32660,N_32661,N_32662,N_32663,N_32664,N_32665,N_32666,N_32667,N_32668,N_32669,N_32670,N_32671,N_32672,N_32673,N_32674,N_32675,N_32676,N_32677,N_32678,N_32679,N_32680,N_32681,N_32682,N_32683,N_32684,N_32685,N_32686,N_32687,N_32688,N_32689,N_32690,N_32691,N_32692,N_32693,N_32694,N_32695,N_32696,N_32697,N_32698,N_32699,N_32700,N_32701,N_32702,N_32703,N_32704,N_32705,N_32706,N_32707,N_32708,N_32709,N_32710,N_32711,N_32712,N_32713,N_32714,N_32715,N_32716,N_32717,N_32718,N_32719,N_32720,N_32721,N_32722,N_32723,N_32724,N_32725,N_32726,N_32727,N_32728,N_32729,N_32730,N_32731,N_32732,N_32733,N_32734,N_32735,N_32736,N_32737,N_32738,N_32739,N_32740,N_32741,N_32742,N_32743,N_32744,N_32745,N_32746,N_32747,N_32748,N_32749,N_32750,N_32751,N_32752,N_32753,N_32754,N_32755,N_32756,N_32757,N_32758,N_32759,N_32760,N_32761,N_32762,N_32763,N_32764,N_32765,N_32766,N_32767,N_32768,N_32769,N_32770,N_32771,N_32772,N_32773,N_32774,N_32775,N_32776,N_32777,N_32778,N_32779,N_32780,N_32781,N_32782,N_32783,N_32784,N_32785,N_32786,N_32787,N_32788,N_32789,N_32790,N_32791,N_32792,N_32793,N_32794,N_32795,N_32796,N_32797,N_32798,N_32799,N_32800,N_32801,N_32802,N_32803,N_32804,N_32805,N_32806,N_32807,N_32808,N_32809,N_32810,N_32811,N_32812,N_32813,N_32814,N_32815,N_32816,N_32817,N_32818,N_32819,N_32820,N_32821,N_32822,N_32823,N_32824,N_32825,N_32826,N_32827,N_32828,N_32829,N_32830,N_32831,N_32832,N_32833,N_32834,N_32835,N_32836,N_32837,N_32838,N_32839,N_32840,N_32841,N_32842,N_32843,N_32844,N_32845,N_32846,N_32847,N_32848,N_32849,N_32850,N_32851,N_32852,N_32853,N_32854,N_32855,N_32856,N_32857,N_32858,N_32859,N_32860,N_32861,N_32862,N_32863,N_32864,N_32865,N_32866,N_32867,N_32868,N_32869,N_32870,N_32871,N_32872,N_32873,N_32874,N_32875,N_32876,N_32877,N_32878,N_32879,N_32880,N_32881,N_32882,N_32883,N_32884,N_32885,N_32886,N_32887,N_32888,N_32889,N_32890,N_32891,N_32892,N_32893,N_32894,N_32895,N_32896,N_32897,N_32898,N_32899,N_32900,N_32901,N_32902,N_32903,N_32904,N_32905,N_32906,N_32907,N_32908,N_32909,N_32910,N_32911,N_32912,N_32913,N_32914,N_32915,N_32916,N_32917,N_32918,N_32919,N_32920,N_32921,N_32922,N_32923,N_32924,N_32925,N_32926,N_32927,N_32928,N_32929,N_32930,N_32931,N_32932,N_32933,N_32934,N_32935,N_32936,N_32937,N_32938,N_32939,N_32940,N_32941,N_32942,N_32943,N_32944,N_32945,N_32946,N_32947,N_32948,N_32949,N_32950,N_32951,N_32952,N_32953,N_32954,N_32955,N_32956,N_32957,N_32958,N_32959,N_32960,N_32961,N_32962,N_32963,N_32964,N_32965,N_32966,N_32967,N_32968,N_32969,N_32970,N_32971,N_32972,N_32973,N_32974,N_32975,N_32976,N_32977,N_32978,N_32979,N_32980,N_32981,N_32982,N_32983,N_32984,N_32985,N_32986,N_32987,N_32988,N_32989,N_32990,N_32991,N_32992,N_32993,N_32994,N_32995,N_32996,N_32997,N_32998,N_32999,N_33000,N_33001,N_33002,N_33003,N_33004,N_33005,N_33006,N_33007,N_33008,N_33009,N_33010,N_33011,N_33012,N_33013,N_33014,N_33015,N_33016,N_33017,N_33018,N_33019,N_33020,N_33021,N_33022,N_33023,N_33024,N_33025,N_33026,N_33027,N_33028,N_33029,N_33030,N_33031,N_33032,N_33033,N_33034,N_33035,N_33036,N_33037,N_33038,N_33039,N_33040,N_33041,N_33042,N_33043,N_33044,N_33045,N_33046,N_33047,N_33048,N_33049,N_33050,N_33051,N_33052,N_33053,N_33054,N_33055,N_33056,N_33057,N_33058,N_33059,N_33060,N_33061,N_33062,N_33063,N_33064,N_33065,N_33066,N_33067,N_33068,N_33069,N_33070,N_33071,N_33072,N_33073,N_33074,N_33075,N_33076,N_33077,N_33078,N_33079,N_33080,N_33081,N_33082,N_33083,N_33084,N_33085,N_33086,N_33087,N_33088,N_33089,N_33090,N_33091,N_33092,N_33093,N_33094,N_33095,N_33096,N_33097,N_33098,N_33099,N_33100,N_33101,N_33102,N_33103,N_33104,N_33105,N_33106,N_33107,N_33108,N_33109,N_33110,N_33111,N_33112,N_33113,N_33114,N_33115,N_33116,N_33117,N_33118,N_33119,N_33120,N_33121,N_33122,N_33123,N_33124,N_33125,N_33126,N_33127,N_33128,N_33129,N_33130,N_33131,N_33132,N_33133,N_33134,N_33135,N_33136,N_33137,N_33138,N_33139,N_33140,N_33141,N_33142,N_33143,N_33144,N_33145,N_33146,N_33147,N_33148,N_33149,N_33150,N_33151,N_33152,N_33153,N_33154,N_33155,N_33156,N_33157,N_33158,N_33159,N_33160,N_33161,N_33162,N_33163,N_33164,N_33165,N_33166,N_33167,N_33168,N_33169,N_33170,N_33171,N_33172,N_33173,N_33174,N_33175,N_33176,N_33177,N_33178,N_33179,N_33180,N_33181,N_33182,N_33183,N_33184,N_33185,N_33186,N_33187,N_33188,N_33189,N_33190,N_33191,N_33192,N_33193,N_33194,N_33195,N_33196,N_33197,N_33198,N_33199,N_33200,N_33201,N_33202,N_33203,N_33204,N_33205,N_33206,N_33207,N_33208,N_33209,N_33210,N_33211,N_33212,N_33213,N_33214,N_33215,N_33216,N_33217,N_33218,N_33219,N_33220,N_33221,N_33222,N_33223,N_33224,N_33225,N_33226,N_33227,N_33228,N_33229,N_33230,N_33231,N_33232,N_33233,N_33234,N_33235,N_33236,N_33237,N_33238,N_33239,N_33240,N_33241,N_33242,N_33243,N_33244,N_33245,N_33246,N_33247,N_33248,N_33249,N_33250,N_33251,N_33252,N_33253,N_33254,N_33255,N_33256,N_33257,N_33258,N_33259,N_33260,N_33261,N_33262,N_33263,N_33264,N_33265,N_33266,N_33267,N_33268,N_33269,N_33270,N_33271,N_33272,N_33273,N_33274,N_33275,N_33276,N_33277,N_33278,N_33279,N_33280,N_33281,N_33282,N_33283,N_33284,N_33285,N_33286,N_33287,N_33288,N_33289,N_33290,N_33291,N_33292,N_33293,N_33294,N_33295,N_33296,N_33297,N_33298,N_33299,N_33300,N_33301,N_33302,N_33303,N_33304,N_33305,N_33306,N_33307,N_33308,N_33309,N_33310,N_33311,N_33312,N_33313,N_33314,N_33315,N_33316,N_33317,N_33318,N_33319,N_33320,N_33321,N_33322,N_33323,N_33324,N_33325,N_33326,N_33327,N_33328,N_33329,N_33330,N_33331,N_33332,N_33333,N_33334,N_33335,N_33336,N_33337,N_33338,N_33339,N_33340,N_33341,N_33342,N_33343,N_33344,N_33345,N_33346,N_33347,N_33348,N_33349,N_33350,N_33351,N_33352,N_33353,N_33354,N_33355,N_33356,N_33357,N_33358,N_33359,N_33360,N_33361,N_33362,N_33363,N_33364,N_33365,N_33366,N_33367,N_33368,N_33369,N_33370,N_33371,N_33372,N_33373,N_33374,N_33375,N_33376,N_33377,N_33378,N_33379,N_33380,N_33381,N_33382,N_33383,N_33384,N_33385,N_33386,N_33387,N_33388,N_33389,N_33390,N_33391,N_33392,N_33393,N_33394,N_33395,N_33396,N_33397,N_33398,N_33399,N_33400,N_33401,N_33402,N_33403,N_33404,N_33405,N_33406,N_33407,N_33408,N_33409,N_33410,N_33411,N_33412,N_33413,N_33414,N_33415,N_33416,N_33417,N_33418,N_33419,N_33420,N_33421,N_33422,N_33423,N_33424,N_33425,N_33426,N_33427,N_33428,N_33429,N_33430,N_33431,N_33432,N_33433,N_33434,N_33435,N_33436,N_33437,N_33438,N_33439,N_33440,N_33441,N_33442,N_33443,N_33444,N_33445,N_33446,N_33447,N_33448,N_33449,N_33450,N_33451,N_33452,N_33453,N_33454,N_33455,N_33456,N_33457,N_33458,N_33459,N_33460,N_33461,N_33462,N_33463,N_33464,N_33465,N_33466,N_33467,N_33468,N_33469,N_33470,N_33471,N_33472,N_33473,N_33474,N_33475,N_33476,N_33477,N_33478,N_33479,N_33480,N_33481,N_33482,N_33483,N_33484,N_33485,N_33486,N_33487,N_33488,N_33489,N_33490,N_33491,N_33492,N_33493,N_33494,N_33495,N_33496,N_33497,N_33498,N_33499,N_33500,N_33501,N_33502,N_33503,N_33504,N_33505,N_33506,N_33507,N_33508,N_33509,N_33510,N_33511,N_33512,N_33513,N_33514,N_33515,N_33516,N_33517,N_33518,N_33519,N_33520,N_33521,N_33522,N_33523,N_33524,N_33525,N_33526,N_33527,N_33528,N_33529,N_33530,N_33531,N_33532,N_33533,N_33534,N_33535,N_33536,N_33537,N_33538,N_33539,N_33540,N_33541,N_33542,N_33543,N_33544,N_33545,N_33546,N_33547,N_33548,N_33549,N_33550,N_33551,N_33552,N_33553,N_33554,N_33555,N_33556,N_33557,N_33558,N_33559,N_33560,N_33561,N_33562,N_33563,N_33564,N_33565,N_33566,N_33567,N_33568,N_33569,N_33570,N_33571,N_33572,N_33573,N_33574,N_33575,N_33576,N_33577,N_33578,N_33579,N_33580,N_33581,N_33582,N_33583,N_33584,N_33585,N_33586,N_33587,N_33588,N_33589,N_33590,N_33591,N_33592,N_33593,N_33594,N_33595,N_33596,N_33597,N_33598,N_33599,N_33600,N_33601,N_33602,N_33603,N_33604,N_33605,N_33606,N_33607,N_33608,N_33609,N_33610,N_33611,N_33612,N_33613,N_33614,N_33615,N_33616,N_33617,N_33618,N_33619,N_33620,N_33621,N_33622,N_33623,N_33624,N_33625,N_33626,N_33627,N_33628,N_33629,N_33630,N_33631,N_33632,N_33633,N_33634,N_33635,N_33636,N_33637,N_33638,N_33639,N_33640,N_33641,N_33642,N_33643,N_33644,N_33645,N_33646,N_33647,N_33648,N_33649,N_33650,N_33651,N_33652,N_33653,N_33654,N_33655,N_33656,N_33657,N_33658,N_33659,N_33660,N_33661,N_33662,N_33663,N_33664,N_33665,N_33666,N_33667,N_33668,N_33669,N_33670,N_33671,N_33672,N_33673,N_33674,N_33675,N_33676,N_33677,N_33678,N_33679,N_33680,N_33681,N_33682,N_33683,N_33684,N_33685,N_33686,N_33687,N_33688,N_33689,N_33690,N_33691,N_33692,N_33693,N_33694,N_33695,N_33696,N_33697,N_33698,N_33699,N_33700,N_33701,N_33702,N_33703,N_33704,N_33705,N_33706,N_33707,N_33708,N_33709,N_33710,N_33711,N_33712,N_33713,N_33714,N_33715,N_33716,N_33717,N_33718,N_33719,N_33720,N_33721,N_33722,N_33723,N_33724,N_33725,N_33726,N_33727,N_33728,N_33729,N_33730,N_33731,N_33732,N_33733,N_33734,N_33735,N_33736,N_33737,N_33738,N_33739,N_33740,N_33741,N_33742,N_33743,N_33744,N_33745,N_33746,N_33747,N_33748,N_33749,N_33750,N_33751,N_33752,N_33753,N_33754,N_33755,N_33756,N_33757,N_33758,N_33759,N_33760,N_33761,N_33762,N_33763,N_33764,N_33765,N_33766,N_33767,N_33768,N_33769,N_33770,N_33771,N_33772,N_33773,N_33774,N_33775,N_33776,N_33777,N_33778,N_33779,N_33780,N_33781,N_33782,N_33783,N_33784,N_33785,N_33786,N_33787,N_33788,N_33789,N_33790,N_33791,N_33792,N_33793,N_33794,N_33795,N_33796,N_33797,N_33798,N_33799,N_33800,N_33801,N_33802,N_33803,N_33804,N_33805,N_33806,N_33807,N_33808,N_33809,N_33810,N_33811,N_33812,N_33813,N_33814,N_33815,N_33816,N_33817,N_33818,N_33819,N_33820,N_33821,N_33822,N_33823,N_33824,N_33825,N_33826,N_33827,N_33828,N_33829,N_33830,N_33831,N_33832,N_33833,N_33834,N_33835,N_33836,N_33837,N_33838,N_33839,N_33840,N_33841,N_33842,N_33843,N_33844,N_33845,N_33846,N_33847,N_33848,N_33849,N_33850,N_33851,N_33852,N_33853,N_33854,N_33855,N_33856,N_33857,N_33858,N_33859,N_33860,N_33861,N_33862,N_33863,N_33864,N_33865,N_33866,N_33867,N_33868,N_33869,N_33870,N_33871,N_33872,N_33873,N_33874,N_33875,N_33876,N_33877,N_33878,N_33879,N_33880,N_33881,N_33882,N_33883,N_33884,N_33885,N_33886,N_33887,N_33888,N_33889,N_33890,N_33891,N_33892,N_33893,N_33894,N_33895,N_33896,N_33897,N_33898,N_33899,N_33900,N_33901,N_33902,N_33903,N_33904,N_33905,N_33906,N_33907,N_33908,N_33909,N_33910,N_33911,N_33912,N_33913,N_33914,N_33915,N_33916,N_33917,N_33918,N_33919,N_33920,N_33921,N_33922,N_33923,N_33924,N_33925,N_33926,N_33927,N_33928,N_33929,N_33930,N_33931,N_33932,N_33933,N_33934,N_33935,N_33936,N_33937,N_33938,N_33939,N_33940,N_33941,N_33942,N_33943,N_33944,N_33945,N_33946,N_33947,N_33948,N_33949,N_33950,N_33951,N_33952,N_33953,N_33954,N_33955,N_33956,N_33957,N_33958,N_33959,N_33960,N_33961,N_33962,N_33963,N_33964,N_33965,N_33966,N_33967,N_33968,N_33969,N_33970,N_33971,N_33972,N_33973,N_33974,N_33975,N_33976,N_33977,N_33978,N_33979,N_33980,N_33981,N_33982,N_33983,N_33984,N_33985,N_33986,N_33987,N_33988,N_33989,N_33990,N_33991,N_33992,N_33993,N_33994,N_33995,N_33996,N_33997,N_33998,N_33999,N_34000,N_34001,N_34002,N_34003,N_34004,N_34005,N_34006,N_34007,N_34008,N_34009,N_34010,N_34011,N_34012,N_34013,N_34014,N_34015,N_34016,N_34017,N_34018,N_34019,N_34020,N_34021,N_34022,N_34023,N_34024,N_34025,N_34026,N_34027,N_34028,N_34029,N_34030,N_34031,N_34032,N_34033,N_34034,N_34035,N_34036,N_34037,N_34038,N_34039,N_34040,N_34041,N_34042,N_34043,N_34044,N_34045,N_34046,N_34047,N_34048,N_34049,N_34050,N_34051,N_34052,N_34053,N_34054,N_34055,N_34056,N_34057,N_34058,N_34059,N_34060,N_34061,N_34062,N_34063,N_34064,N_34065,N_34066,N_34067,N_34068,N_34069,N_34070,N_34071,N_34072,N_34073,N_34074,N_34075,N_34076,N_34077,N_34078,N_34079,N_34080,N_34081,N_34082,N_34083,N_34084,N_34085,N_34086,N_34087,N_34088,N_34089,N_34090,N_34091,N_34092,N_34093,N_34094,N_34095,N_34096,N_34097,N_34098,N_34099,N_34100,N_34101,N_34102,N_34103,N_34104,N_34105,N_34106,N_34107,N_34108,N_34109,N_34110,N_34111,N_34112,N_34113,N_34114,N_34115,N_34116,N_34117,N_34118,N_34119,N_34120,N_34121,N_34122,N_34123,N_34124,N_34125,N_34126,N_34127,N_34128,N_34129,N_34130,N_34131,N_34132,N_34133,N_34134,N_34135,N_34136,N_34137,N_34138,N_34139,N_34140,N_34141,N_34142,N_34143,N_34144,N_34145,N_34146,N_34147,N_34148,N_34149,N_34150,N_34151,N_34152,N_34153,N_34154,N_34155,N_34156,N_34157,N_34158,N_34159,N_34160,N_34161,N_34162,N_34163,N_34164,N_34165,N_34166,N_34167,N_34168,N_34169,N_34170,N_34171,N_34172,N_34173,N_34174,N_34175,N_34176,N_34177,N_34178,N_34179,N_34180,N_34181,N_34182,N_34183,N_34184,N_34185,N_34186,N_34187,N_34188,N_34189,N_34190,N_34191,N_34192,N_34193,N_34194,N_34195,N_34196,N_34197,N_34198,N_34199,N_34200,N_34201,N_34202,N_34203,N_34204,N_34205,N_34206,N_34207,N_34208,N_34209,N_34210,N_34211,N_34212,N_34213,N_34214,N_34215,N_34216,N_34217,N_34218,N_34219,N_34220,N_34221,N_34222,N_34223,N_34224,N_34225,N_34226,N_34227,N_34228,N_34229,N_34230,N_34231,N_34232,N_34233,N_34234,N_34235,N_34236,N_34237,N_34238,N_34239,N_34240,N_34241,N_34242,N_34243,N_34244,N_34245,N_34246,N_34247,N_34248,N_34249,N_34250,N_34251,N_34252,N_34253,N_34254,N_34255,N_34256,N_34257,N_34258,N_34259,N_34260,N_34261,N_34262,N_34263,N_34264,N_34265,N_34266,N_34267,N_34268,N_34269,N_34270,N_34271,N_34272,N_34273,N_34274,N_34275,N_34276,N_34277,N_34278,N_34279,N_34280,N_34281,N_34282,N_34283,N_34284,N_34285,N_34286,N_34287,N_34288,N_34289,N_34290,N_34291,N_34292,N_34293,N_34294,N_34295,N_34296,N_34297,N_34298,N_34299,N_34300,N_34301,N_34302,N_34303,N_34304,N_34305,N_34306,N_34307,N_34308,N_34309,N_34310,N_34311,N_34312,N_34313,N_34314,N_34315,N_34316,N_34317,N_34318,N_34319,N_34320,N_34321,N_34322,N_34323,N_34324,N_34325,N_34326,N_34327,N_34328,N_34329,N_34330,N_34331,N_34332,N_34333,N_34334,N_34335,N_34336,N_34337,N_34338,N_34339,N_34340,N_34341,N_34342,N_34343,N_34344,N_34345,N_34346,N_34347,N_34348,N_34349,N_34350,N_34351,N_34352,N_34353,N_34354,N_34355,N_34356,N_34357,N_34358,N_34359,N_34360,N_34361,N_34362,N_34363,N_34364,N_34365,N_34366,N_34367,N_34368,N_34369,N_34370,N_34371,N_34372,N_34373,N_34374,N_34375,N_34376,N_34377,N_34378,N_34379,N_34380,N_34381,N_34382,N_34383,N_34384,N_34385,N_34386,N_34387,N_34388,N_34389,N_34390,N_34391,N_34392,N_34393,N_34394,N_34395,N_34396,N_34397,N_34398,N_34399,N_34400,N_34401,N_34402,N_34403,N_34404,N_34405,N_34406,N_34407,N_34408,N_34409,N_34410,N_34411,N_34412,N_34413,N_34414,N_34415,N_34416,N_34417,N_34418,N_34419,N_34420,N_34421,N_34422,N_34423,N_34424,N_34425,N_34426,N_34427,N_34428,N_34429,N_34430,N_34431,N_34432,N_34433,N_34434,N_34435,N_34436,N_34437,N_34438,N_34439,N_34440,N_34441,N_34442,N_34443,N_34444,N_34445,N_34446,N_34447,N_34448,N_34449,N_34450,N_34451,N_34452,N_34453,N_34454,N_34455,N_34456,N_34457,N_34458,N_34459,N_34460,N_34461,N_34462,N_34463,N_34464,N_34465,N_34466,N_34467,N_34468,N_34469,N_34470,N_34471,N_34472,N_34473,N_34474,N_34475,N_34476,N_34477,N_34478,N_34479,N_34480,N_34481,N_34482,N_34483,N_34484,N_34485,N_34486,N_34487,N_34488,N_34489,N_34490,N_34491,N_34492,N_34493,N_34494,N_34495,N_34496,N_34497,N_34498,N_34499,N_34500,N_34501,N_34502,N_34503,N_34504,N_34505,N_34506,N_34507,N_34508,N_34509,N_34510,N_34511,N_34512,N_34513,N_34514,N_34515,N_34516,N_34517,N_34518,N_34519,N_34520,N_34521,N_34522,N_34523,N_34524,N_34525,N_34526,N_34527,N_34528,N_34529,N_34530,N_34531,N_34532,N_34533,N_34534,N_34535,N_34536,N_34537,N_34538,N_34539,N_34540,N_34541,N_34542,N_34543,N_34544,N_34545,N_34546,N_34547,N_34548,N_34549,N_34550,N_34551,N_34552,N_34553,N_34554,N_34555,N_34556,N_34557,N_34558,N_34559,N_34560,N_34561,N_34562,N_34563,N_34564,N_34565,N_34566,N_34567,N_34568,N_34569,N_34570,N_34571,N_34572,N_34573,N_34574,N_34575,N_34576,N_34577,N_34578,N_34579,N_34580,N_34581,N_34582,N_34583,N_34584,N_34585,N_34586,N_34587,N_34588,N_34589,N_34590,N_34591,N_34592,N_34593,N_34594,N_34595,N_34596,N_34597,N_34598,N_34599,N_34600,N_34601,N_34602,N_34603,N_34604,N_34605,N_34606,N_34607,N_34608,N_34609,N_34610,N_34611,N_34612,N_34613,N_34614,N_34615,N_34616,N_34617,N_34618,N_34619,N_34620,N_34621,N_34622,N_34623,N_34624,N_34625,N_34626,N_34627,N_34628,N_34629,N_34630,N_34631,N_34632,N_34633,N_34634,N_34635,N_34636,N_34637,N_34638,N_34639,N_34640,N_34641,N_34642,N_34643,N_34644,N_34645,N_34646,N_34647,N_34648,N_34649,N_34650,N_34651,N_34652,N_34653,N_34654,N_34655,N_34656,N_34657,N_34658,N_34659,N_34660,N_34661,N_34662,N_34663,N_34664,N_34665,N_34666,N_34667,N_34668,N_34669,N_34670,N_34671,N_34672,N_34673,N_34674,N_34675,N_34676,N_34677,N_34678,N_34679,N_34680,N_34681,N_34682,N_34683,N_34684,N_34685,N_34686,N_34687,N_34688,N_34689,N_34690,N_34691,N_34692,N_34693,N_34694,N_34695,N_34696,N_34697,N_34698,N_34699,N_34700,N_34701,N_34702,N_34703,N_34704,N_34705,N_34706,N_34707,N_34708,N_34709,N_34710,N_34711,N_34712,N_34713,N_34714,N_34715,N_34716,N_34717,N_34718,N_34719,N_34720,N_34721,N_34722,N_34723,N_34724,N_34725,N_34726,N_34727,N_34728,N_34729,N_34730,N_34731,N_34732,N_34733,N_34734,N_34735,N_34736,N_34737,N_34738,N_34739,N_34740,N_34741,N_34742,N_34743,N_34744,N_34745,N_34746,N_34747,N_34748,N_34749,N_34750,N_34751,N_34752,N_34753,N_34754,N_34755,N_34756,N_34757,N_34758,N_34759,N_34760,N_34761,N_34762,N_34763,N_34764,N_34765,N_34766,N_34767,N_34768,N_34769,N_34770,N_34771,N_34772,N_34773,N_34774,N_34775,N_34776,N_34777,N_34778,N_34779,N_34780,N_34781,N_34782,N_34783,N_34784,N_34785,N_34786,N_34787,N_34788,N_34789,N_34790,N_34791,N_34792,N_34793,N_34794,N_34795,N_34796,N_34797,N_34798,N_34799,N_34800,N_34801,N_34802,N_34803,N_34804,N_34805,N_34806,N_34807,N_34808,N_34809,N_34810,N_34811,N_34812,N_34813,N_34814,N_34815,N_34816,N_34817,N_34818,N_34819,N_34820,N_34821,N_34822,N_34823,N_34824,N_34825,N_34826,N_34827,N_34828,N_34829,N_34830,N_34831,N_34832,N_34833,N_34834,N_34835,N_34836,N_34837,N_34838,N_34839,N_34840,N_34841,N_34842,N_34843,N_34844,N_34845,N_34846,N_34847,N_34848,N_34849,N_34850,N_34851,N_34852,N_34853,N_34854,N_34855,N_34856,N_34857,N_34858,N_34859,N_34860,N_34861,N_34862,N_34863,N_34864,N_34865,N_34866,N_34867,N_34868,N_34869,N_34870,N_34871,N_34872,N_34873,N_34874,N_34875,N_34876,N_34877,N_34878,N_34879,N_34880,N_34881,N_34882,N_34883,N_34884,N_34885,N_34886,N_34887,N_34888,N_34889,N_34890,N_34891,N_34892,N_34893,N_34894,N_34895,N_34896,N_34897,N_34898,N_34899,N_34900,N_34901,N_34902,N_34903,N_34904,N_34905,N_34906,N_34907,N_34908,N_34909,N_34910,N_34911,N_34912,N_34913,N_34914,N_34915,N_34916,N_34917,N_34918,N_34919,N_34920,N_34921,N_34922,N_34923,N_34924,N_34925,N_34926,N_34927,N_34928,N_34929,N_34930,N_34931,N_34932,N_34933,N_34934,N_34935,N_34936,N_34937,N_34938,N_34939,N_34940,N_34941,N_34942,N_34943,N_34944,N_34945,N_34946,N_34947,N_34948,N_34949,N_34950,N_34951,N_34952,N_34953,N_34954,N_34955,N_34956,N_34957,N_34958,N_34959,N_34960,N_34961,N_34962,N_34963,N_34964,N_34965,N_34966,N_34967,N_34968,N_34969,N_34970,N_34971,N_34972,N_34973,N_34974,N_34975,N_34976,N_34977,N_34978,N_34979,N_34980,N_34981,N_34982,N_34983,N_34984,N_34985,N_34986,N_34987,N_34988,N_34989,N_34990,N_34991,N_34992,N_34993,N_34994,N_34995,N_34996,N_34997,N_34998,N_34999,N_35000,N_35001,N_35002,N_35003,N_35004,N_35005,N_35006,N_35007,N_35008,N_35009,N_35010,N_35011,N_35012,N_35013,N_35014,N_35015,N_35016,N_35017,N_35018,N_35019,N_35020,N_35021,N_35022,N_35023,N_35024,N_35025,N_35026,N_35027,N_35028,N_35029,N_35030,N_35031,N_35032,N_35033,N_35034,N_35035,N_35036,N_35037,N_35038,N_35039,N_35040,N_35041,N_35042,N_35043,N_35044,N_35045,N_35046,N_35047,N_35048,N_35049,N_35050,N_35051,N_35052,N_35053,N_35054,N_35055,N_35056,N_35057,N_35058,N_35059,N_35060,N_35061,N_35062,N_35063,N_35064,N_35065,N_35066,N_35067,N_35068,N_35069,N_35070,N_35071,N_35072,N_35073,N_35074,N_35075,N_35076,N_35077,N_35078,N_35079,N_35080,N_35081,N_35082,N_35083,N_35084,N_35085,N_35086,N_35087,N_35088,N_35089,N_35090,N_35091,N_35092,N_35093,N_35094,N_35095,N_35096,N_35097,N_35098,N_35099,N_35100,N_35101,N_35102,N_35103,N_35104,N_35105,N_35106,N_35107,N_35108,N_35109,N_35110,N_35111,N_35112,N_35113,N_35114,N_35115,N_35116,N_35117,N_35118,N_35119,N_35120,N_35121,N_35122,N_35123,N_35124,N_35125,N_35126,N_35127,N_35128,N_35129,N_35130,N_35131,N_35132,N_35133,N_35134,N_35135,N_35136,N_35137,N_35138,N_35139,N_35140,N_35141,N_35142,N_35143,N_35144,N_35145,N_35146,N_35147,N_35148,N_35149,N_35150,N_35151,N_35152,N_35153,N_35154,N_35155,N_35156,N_35157,N_35158,N_35159,N_35160,N_35161,N_35162,N_35163,N_35164,N_35165,N_35166,N_35167,N_35168,N_35169,N_35170,N_35171,N_35172,N_35173,N_35174,N_35175,N_35176,N_35177,N_35178,N_35179,N_35180,N_35181,N_35182,N_35183,N_35184,N_35185,N_35186,N_35187,N_35188,N_35189,N_35190,N_35191,N_35192,N_35193,N_35194,N_35195,N_35196,N_35197,N_35198,N_35199,N_35200,N_35201,N_35202,N_35203,N_35204,N_35205,N_35206,N_35207,N_35208,N_35209,N_35210,N_35211,N_35212,N_35213,N_35214,N_35215,N_35216,N_35217,N_35218,N_35219,N_35220,N_35221,N_35222,N_35223,N_35224,N_35225,N_35226,N_35227,N_35228,N_35229,N_35230,N_35231,N_35232,N_35233,N_35234,N_35235,N_35236,N_35237,N_35238,N_35239,N_35240,N_35241,N_35242,N_35243,N_35244,N_35245,N_35246,N_35247,N_35248,N_35249,N_35250,N_35251,N_35252,N_35253,N_35254,N_35255,N_35256,N_35257,N_35258,N_35259,N_35260,N_35261,N_35262,N_35263,N_35264,N_35265,N_35266,N_35267,N_35268,N_35269,N_35270,N_35271,N_35272,N_35273,N_35274,N_35275,N_35276,N_35277,N_35278,N_35279,N_35280,N_35281,N_35282,N_35283,N_35284,N_35285,N_35286,N_35287,N_35288,N_35289,N_35290,N_35291,N_35292,N_35293,N_35294,N_35295,N_35296,N_35297,N_35298,N_35299,N_35300,N_35301,N_35302,N_35303,N_35304,N_35305,N_35306,N_35307,N_35308,N_35309,N_35310,N_35311,N_35312,N_35313,N_35314,N_35315,N_35316,N_35317,N_35318,N_35319,N_35320,N_35321,N_35322,N_35323,N_35324,N_35325,N_35326,N_35327,N_35328,N_35329,N_35330,N_35331,N_35332,N_35333,N_35334,N_35335,N_35336,N_35337,N_35338,N_35339,N_35340,N_35341,N_35342,N_35343,N_35344,N_35345,N_35346,N_35347,N_35348,N_35349,N_35350,N_35351,N_35352,N_35353,N_35354,N_35355,N_35356,N_35357,N_35358,N_35359,N_35360,N_35361,N_35362,N_35363,N_35364,N_35365,N_35366,N_35367,N_35368,N_35369,N_35370,N_35371,N_35372,N_35373,N_35374,N_35375,N_35376,N_35377,N_35378,N_35379,N_35380,N_35381,N_35382,N_35383,N_35384,N_35385,N_35386,N_35387,N_35388,N_35389,N_35390,N_35391,N_35392,N_35393,N_35394,N_35395,N_35396,N_35397,N_35398,N_35399,N_35400,N_35401,N_35402,N_35403,N_35404,N_35405,N_35406,N_35407,N_35408,N_35409,N_35410,N_35411,N_35412,N_35413,N_35414,N_35415,N_35416,N_35417,N_35418,N_35419,N_35420,N_35421,N_35422,N_35423,N_35424,N_35425,N_35426,N_35427,N_35428,N_35429,N_35430,N_35431,N_35432,N_35433,N_35434,N_35435,N_35436,N_35437,N_35438,N_35439,N_35440,N_35441,N_35442,N_35443,N_35444,N_35445,N_35446,N_35447,N_35448,N_35449,N_35450,N_35451,N_35452,N_35453,N_35454,N_35455,N_35456,N_35457,N_35458,N_35459,N_35460,N_35461,N_35462,N_35463,N_35464,N_35465,N_35466,N_35467,N_35468,N_35469,N_35470,N_35471,N_35472,N_35473,N_35474,N_35475,N_35476,N_35477,N_35478,N_35479,N_35480,N_35481,N_35482,N_35483,N_35484,N_35485,N_35486,N_35487,N_35488,N_35489,N_35490,N_35491,N_35492,N_35493,N_35494,N_35495,N_35496,N_35497,N_35498,N_35499,N_35500,N_35501,N_35502,N_35503,N_35504,N_35505,N_35506,N_35507,N_35508,N_35509,N_35510,N_35511,N_35512,N_35513,N_35514,N_35515,N_35516,N_35517,N_35518,N_35519,N_35520,N_35521,N_35522,N_35523,N_35524,N_35525,N_35526,N_35527,N_35528,N_35529,N_35530,N_35531,N_35532,N_35533,N_35534,N_35535,N_35536,N_35537,N_35538,N_35539,N_35540,N_35541,N_35542,N_35543,N_35544,N_35545,N_35546,N_35547,N_35548,N_35549,N_35550,N_35551,N_35552,N_35553,N_35554,N_35555,N_35556,N_35557,N_35558,N_35559,N_35560,N_35561,N_35562,N_35563,N_35564,N_35565,N_35566,N_35567,N_35568,N_35569,N_35570,N_35571,N_35572,N_35573,N_35574,N_35575,N_35576,N_35577,N_35578,N_35579,N_35580,N_35581,N_35582,N_35583,N_35584,N_35585,N_35586,N_35587,N_35588,N_35589,N_35590,N_35591,N_35592,N_35593,N_35594,N_35595,N_35596,N_35597,N_35598,N_35599,N_35600,N_35601,N_35602,N_35603,N_35604,N_35605,N_35606,N_35607,N_35608,N_35609,N_35610,N_35611,N_35612,N_35613,N_35614,N_35615,N_35616,N_35617,N_35618,N_35619,N_35620,N_35621,N_35622,N_35623,N_35624,N_35625,N_35626,N_35627,N_35628,N_35629,N_35630,N_35631,N_35632,N_35633,N_35634,N_35635,N_35636,N_35637,N_35638,N_35639,N_35640,N_35641,N_35642,N_35643,N_35644,N_35645,N_35646,N_35647,N_35648,N_35649,N_35650,N_35651,N_35652,N_35653,N_35654,N_35655,N_35656,N_35657,N_35658,N_35659,N_35660,N_35661,N_35662,N_35663,N_35664,N_35665,N_35666,N_35667,N_35668,N_35669,N_35670,N_35671,N_35672,N_35673,N_35674,N_35675,N_35676,N_35677,N_35678,N_35679,N_35680,N_35681,N_35682,N_35683,N_35684,N_35685,N_35686,N_35687,N_35688,N_35689,N_35690,N_35691,N_35692,N_35693,N_35694,N_35695,N_35696,N_35697,N_35698,N_35699,N_35700,N_35701,N_35702,N_35703,N_35704,N_35705,N_35706,N_35707,N_35708,N_35709,N_35710,N_35711,N_35712,N_35713,N_35714,N_35715,N_35716,N_35717,N_35718,N_35719,N_35720,N_35721,N_35722,N_35723,N_35724,N_35725,N_35726,N_35727,N_35728,N_35729,N_35730,N_35731,N_35732,N_35733,N_35734,N_35735,N_35736,N_35737,N_35738,N_35739,N_35740,N_35741,N_35742,N_35743,N_35744,N_35745,N_35746,N_35747,N_35748,N_35749,N_35750,N_35751,N_35752,N_35753,N_35754,N_35755,N_35756,N_35757,N_35758,N_35759,N_35760,N_35761,N_35762,N_35763,N_35764,N_35765,N_35766,N_35767,N_35768,N_35769,N_35770,N_35771,N_35772,N_35773,N_35774,N_35775,N_35776,N_35777,N_35778,N_35779,N_35780,N_35781,N_35782,N_35783,N_35784,N_35785,N_35786,N_35787,N_35788,N_35789,N_35790,N_35791,N_35792,N_35793,N_35794,N_35795,N_35796,N_35797,N_35798,N_35799,N_35800,N_35801,N_35802,N_35803,N_35804,N_35805,N_35806,N_35807,N_35808,N_35809,N_35810,N_35811,N_35812,N_35813,N_35814,N_35815,N_35816,N_35817,N_35818,N_35819,N_35820,N_35821,N_35822,N_35823,N_35824,N_35825,N_35826,N_35827,N_35828,N_35829,N_35830,N_35831,N_35832,N_35833,N_35834,N_35835,N_35836,N_35837,N_35838,N_35839,N_35840,N_35841,N_35842,N_35843,N_35844,N_35845,N_35846,N_35847,N_35848,N_35849,N_35850,N_35851,N_35852,N_35853,N_35854,N_35855,N_35856,N_35857,N_35858,N_35859,N_35860,N_35861,N_35862,N_35863,N_35864,N_35865,N_35866,N_35867,N_35868,N_35869,N_35870,N_35871,N_35872,N_35873,N_35874,N_35875,N_35876,N_35877,N_35878,N_35879,N_35880,N_35881,N_35882,N_35883,N_35884,N_35885,N_35886,N_35887,N_35888,N_35889,N_35890,N_35891,N_35892,N_35893,N_35894,N_35895,N_35896,N_35897,N_35898,N_35899,N_35900,N_35901,N_35902,N_35903,N_35904,N_35905,N_35906,N_35907,N_35908,N_35909,N_35910,N_35911,N_35912,N_35913,N_35914,N_35915,N_35916,N_35917,N_35918,N_35919,N_35920,N_35921,N_35922,N_35923,N_35924,N_35925,N_35926,N_35927,N_35928,N_35929,N_35930,N_35931,N_35932,N_35933,N_35934,N_35935,N_35936,N_35937,N_35938,N_35939,N_35940,N_35941,N_35942,N_35943,N_35944,N_35945,N_35946,N_35947,N_35948,N_35949,N_35950,N_35951,N_35952,N_35953,N_35954,N_35955,N_35956,N_35957,N_35958,N_35959,N_35960,N_35961,N_35962,N_35963,N_35964,N_35965,N_35966,N_35967,N_35968,N_35969,N_35970,N_35971,N_35972,N_35973,N_35974,N_35975,N_35976,N_35977,N_35978,N_35979,N_35980,N_35981,N_35982,N_35983,N_35984,N_35985,N_35986,N_35987,N_35988,N_35989,N_35990,N_35991,N_35992,N_35993,N_35994,N_35995,N_35996,N_35997,N_35998,N_35999,N_36000,N_36001,N_36002,N_36003,N_36004,N_36005,N_36006,N_36007,N_36008,N_36009,N_36010,N_36011,N_36012,N_36013,N_36014,N_36015,N_36016,N_36017,N_36018,N_36019,N_36020,N_36021,N_36022,N_36023,N_36024,N_36025,N_36026,N_36027,N_36028,N_36029,N_36030,N_36031,N_36032,N_36033,N_36034,N_36035,N_36036,N_36037,N_36038,N_36039,N_36040,N_36041,N_36042,N_36043,N_36044,N_36045,N_36046,N_36047,N_36048,N_36049,N_36050,N_36051,N_36052,N_36053,N_36054,N_36055,N_36056,N_36057,N_36058,N_36059,N_36060,N_36061,N_36062,N_36063,N_36064,N_36065,N_36066,N_36067,N_36068,N_36069,N_36070,N_36071,N_36072,N_36073,N_36074,N_36075,N_36076,N_36077,N_36078,N_36079,N_36080,N_36081,N_36082,N_36083,N_36084,N_36085,N_36086,N_36087,N_36088,N_36089,N_36090,N_36091,N_36092,N_36093,N_36094,N_36095,N_36096,N_36097,N_36098,N_36099,N_36100,N_36101,N_36102,N_36103,N_36104,N_36105,N_36106,N_36107,N_36108,N_36109,N_36110,N_36111,N_36112,N_36113,N_36114,N_36115,N_36116,N_36117,N_36118,N_36119,N_36120,N_36121,N_36122,N_36123,N_36124,N_36125,N_36126,N_36127,N_36128,N_36129,N_36130,N_36131,N_36132,N_36133,N_36134,N_36135,N_36136,N_36137,N_36138,N_36139,N_36140,N_36141,N_36142,N_36143,N_36144,N_36145,N_36146,N_36147,N_36148,N_36149,N_36150,N_36151,N_36152,N_36153,N_36154,N_36155,N_36156,N_36157,N_36158,N_36159,N_36160,N_36161,N_36162,N_36163,N_36164,N_36165,N_36166,N_36167,N_36168,N_36169,N_36170,N_36171,N_36172,N_36173,N_36174,N_36175,N_36176,N_36177,N_36178,N_36179,N_36180,N_36181,N_36182,N_36183,N_36184,N_36185,N_36186,N_36187,N_36188,N_36189,N_36190,N_36191,N_36192,N_36193,N_36194,N_36195,N_36196,N_36197,N_36198,N_36199,N_36200,N_36201,N_36202,N_36203,N_36204,N_36205,N_36206,N_36207,N_36208,N_36209,N_36210,N_36211,N_36212,N_36213,N_36214,N_36215,N_36216,N_36217,N_36218,N_36219,N_36220,N_36221,N_36222,N_36223,N_36224,N_36225,N_36226,N_36227,N_36228,N_36229,N_36230,N_36231,N_36232,N_36233,N_36234,N_36235,N_36236,N_36237,N_36238,N_36239,N_36240,N_36241,N_36242,N_36243,N_36244,N_36245,N_36246,N_36247,N_36248,N_36249,N_36250,N_36251,N_36252,N_36253,N_36254,N_36255,N_36256,N_36257,N_36258,N_36259,N_36260,N_36261,N_36262,N_36263,N_36264,N_36265,N_36266,N_36267,N_36268,N_36269,N_36270,N_36271,N_36272,N_36273,N_36274,N_36275,N_36276,N_36277,N_36278,N_36279,N_36280,N_36281,N_36282,N_36283,N_36284,N_36285,N_36286,N_36287,N_36288,N_36289,N_36290,N_36291,N_36292,N_36293,N_36294,N_36295,N_36296,N_36297,N_36298,N_36299,N_36300,N_36301,N_36302,N_36303,N_36304,N_36305,N_36306,N_36307,N_36308,N_36309,N_36310,N_36311,N_36312,N_36313,N_36314,N_36315,N_36316,N_36317,N_36318,N_36319,N_36320,N_36321,N_36322,N_36323,N_36324,N_36325,N_36326,N_36327,N_36328,N_36329,N_36330,N_36331,N_36332,N_36333,N_36334,N_36335,N_36336,N_36337,N_36338,N_36339,N_36340,N_36341,N_36342,N_36343,N_36344,N_36345,N_36346,N_36347,N_36348,N_36349,N_36350,N_36351,N_36352,N_36353,N_36354,N_36355,N_36356,N_36357,N_36358,N_36359,N_36360,N_36361,N_36362,N_36363,N_36364,N_36365,N_36366,N_36367,N_36368,N_36369,N_36370,N_36371,N_36372,N_36373,N_36374,N_36375,N_36376,N_36377,N_36378,N_36379,N_36380,N_36381,N_36382,N_36383,N_36384,N_36385,N_36386,N_36387,N_36388,N_36389,N_36390,N_36391,N_36392,N_36393,N_36394,N_36395,N_36396,N_36397,N_36398,N_36399,N_36400,N_36401,N_36402,N_36403,N_36404,N_36405,N_36406,N_36407,N_36408,N_36409,N_36410,N_36411,N_36412,N_36413,N_36414,N_36415,N_36416,N_36417,N_36418,N_36419,N_36420,N_36421,N_36422,N_36423,N_36424,N_36425,N_36426,N_36427,N_36428,N_36429,N_36430,N_36431,N_36432,N_36433,N_36434,N_36435,N_36436,N_36437,N_36438,N_36439,N_36440,N_36441,N_36442,N_36443,N_36444,N_36445,N_36446,N_36447,N_36448,N_36449,N_36450,N_36451,N_36452,N_36453,N_36454,N_36455,N_36456,N_36457,N_36458,N_36459,N_36460,N_36461,N_36462,N_36463,N_36464,N_36465,N_36466,N_36467,N_36468,N_36469,N_36470,N_36471,N_36472,N_36473,N_36474,N_36475,N_36476,N_36477,N_36478,N_36479,N_36480,N_36481,N_36482,N_36483,N_36484,N_36485,N_36486,N_36487,N_36488,N_36489,N_36490,N_36491,N_36492,N_36493,N_36494,N_36495,N_36496,N_36497,N_36498,N_36499,N_36500,N_36501,N_36502,N_36503,N_36504,N_36505,N_36506,N_36507,N_36508,N_36509,N_36510,N_36511,N_36512,N_36513,N_36514,N_36515,N_36516,N_36517,N_36518,N_36519,N_36520,N_36521,N_36522,N_36523,N_36524,N_36525,N_36526,N_36527,N_36528,N_36529,N_36530,N_36531,N_36532,N_36533,N_36534,N_36535,N_36536,N_36537,N_36538,N_36539,N_36540,N_36541,N_36542,N_36543,N_36544,N_36545,N_36546,N_36547,N_36548,N_36549,N_36550,N_36551,N_36552,N_36553,N_36554,N_36555,N_36556,N_36557,N_36558,N_36559,N_36560,N_36561,N_36562,N_36563,N_36564,N_36565,N_36566,N_36567,N_36568,N_36569,N_36570,N_36571,N_36572,N_36573,N_36574,N_36575,N_36576,N_36577,N_36578,N_36579,N_36580,N_36581,N_36582,N_36583,N_36584,N_36585,N_36586,N_36587,N_36588,N_36589,N_36590,N_36591,N_36592,N_36593,N_36594,N_36595,N_36596,N_36597,N_36598,N_36599,N_36600,N_36601,N_36602,N_36603,N_36604,N_36605,N_36606,N_36607,N_36608,N_36609,N_36610,N_36611,N_36612,N_36613,N_36614,N_36615,N_36616,N_36617,N_36618,N_36619,N_36620,N_36621,N_36622,N_36623,N_36624,N_36625,N_36626,N_36627,N_36628,N_36629,N_36630,N_36631,N_36632,N_36633,N_36634,N_36635,N_36636,N_36637,N_36638,N_36639,N_36640,N_36641,N_36642,N_36643,N_36644,N_36645,N_36646,N_36647,N_36648,N_36649,N_36650,N_36651,N_36652,N_36653,N_36654,N_36655,N_36656,N_36657,N_36658,N_36659,N_36660,N_36661,N_36662,N_36663,N_36664,N_36665,N_36666,N_36667,N_36668,N_36669,N_36670,N_36671,N_36672,N_36673,N_36674,N_36675,N_36676,N_36677,N_36678,N_36679,N_36680,N_36681,N_36682,N_36683,N_36684,N_36685,N_36686,N_36687,N_36688,N_36689,N_36690,N_36691,N_36692,N_36693,N_36694,N_36695,N_36696,N_36697,N_36698,N_36699,N_36700,N_36701,N_36702,N_36703,N_36704,N_36705,N_36706,N_36707,N_36708,N_36709,N_36710,N_36711,N_36712,N_36713,N_36714,N_36715,N_36716,N_36717,N_36718,N_36719,N_36720,N_36721,N_36722,N_36723,N_36724,N_36725,N_36726,N_36727,N_36728,N_36729,N_36730,N_36731,N_36732,N_36733,N_36734,N_36735,N_36736,N_36737,N_36738,N_36739,N_36740,N_36741,N_36742,N_36743,N_36744,N_36745,N_36746,N_36747,N_36748,N_36749,N_36750,N_36751,N_36752,N_36753,N_36754,N_36755,N_36756,N_36757,N_36758,N_36759,N_36760,N_36761,N_36762,N_36763,N_36764,N_36765,N_36766,N_36767,N_36768,N_36769,N_36770,N_36771,N_36772,N_36773,N_36774,N_36775,N_36776,N_36777,N_36778,N_36779,N_36780,N_36781,N_36782,N_36783,N_36784,N_36785,N_36786,N_36787,N_36788,N_36789,N_36790,N_36791,N_36792,N_36793,N_36794,N_36795,N_36796,N_36797,N_36798,N_36799,N_36800,N_36801,N_36802,N_36803,N_36804,N_36805,N_36806,N_36807,N_36808,N_36809,N_36810,N_36811,N_36812,N_36813,N_36814,N_36815,N_36816,N_36817,N_36818,N_36819,N_36820,N_36821,N_36822,N_36823,N_36824,N_36825,N_36826,N_36827,N_36828,N_36829,N_36830,N_36831,N_36832,N_36833,N_36834,N_36835,N_36836,N_36837,N_36838,N_36839,N_36840,N_36841,N_36842,N_36843,N_36844,N_36845,N_36846,N_36847,N_36848,N_36849,N_36850,N_36851,N_36852,N_36853,N_36854,N_36855,N_36856,N_36857,N_36858,N_36859,N_36860,N_36861,N_36862,N_36863,N_36864,N_36865,N_36866,N_36867,N_36868,N_36869,N_36870,N_36871,N_36872,N_36873,N_36874,N_36875,N_36876,N_36877,N_36878,N_36879,N_36880,N_36881,N_36882,N_36883,N_36884,N_36885,N_36886,N_36887,N_36888,N_36889,N_36890,N_36891,N_36892,N_36893,N_36894,N_36895,N_36896,N_36897,N_36898,N_36899,N_36900,N_36901,N_36902,N_36903,N_36904,N_36905,N_36906,N_36907,N_36908,N_36909,N_36910,N_36911,N_36912,N_36913,N_36914,N_36915,N_36916,N_36917,N_36918,N_36919,N_36920,N_36921,N_36922,N_36923,N_36924,N_36925,N_36926,N_36927,N_36928,N_36929,N_36930,N_36931,N_36932,N_36933,N_36934,N_36935,N_36936,N_36937,N_36938,N_36939,N_36940,N_36941,N_36942,N_36943,N_36944,N_36945,N_36946,N_36947,N_36948,N_36949,N_36950,N_36951,N_36952,N_36953,N_36954,N_36955,N_36956,N_36957,N_36958,N_36959,N_36960,N_36961,N_36962,N_36963,N_36964,N_36965,N_36966,N_36967,N_36968,N_36969,N_36970,N_36971,N_36972,N_36973,N_36974,N_36975,N_36976,N_36977,N_36978,N_36979,N_36980,N_36981,N_36982,N_36983,N_36984,N_36985,N_36986,N_36987,N_36988,N_36989,N_36990,N_36991,N_36992,N_36993,N_36994,N_36995,N_36996,N_36997,N_36998,N_36999,N_37000,N_37001,N_37002,N_37003,N_37004,N_37005,N_37006,N_37007,N_37008,N_37009,N_37010,N_37011,N_37012,N_37013,N_37014,N_37015,N_37016,N_37017,N_37018,N_37019,N_37020,N_37021,N_37022,N_37023,N_37024,N_37025,N_37026,N_37027,N_37028,N_37029,N_37030,N_37031,N_37032,N_37033,N_37034,N_37035,N_37036,N_37037,N_37038,N_37039,N_37040,N_37041,N_37042,N_37043,N_37044,N_37045,N_37046,N_37047,N_37048,N_37049,N_37050,N_37051,N_37052,N_37053,N_37054,N_37055,N_37056,N_37057,N_37058,N_37059,N_37060,N_37061,N_37062,N_37063,N_37064,N_37065,N_37066,N_37067,N_37068,N_37069,N_37070,N_37071,N_37072,N_37073,N_37074,N_37075,N_37076,N_37077,N_37078,N_37079,N_37080,N_37081,N_37082,N_37083,N_37084,N_37085,N_37086,N_37087,N_37088,N_37089,N_37090,N_37091,N_37092,N_37093,N_37094,N_37095,N_37096,N_37097,N_37098,N_37099,N_37100,N_37101,N_37102,N_37103,N_37104,N_37105,N_37106,N_37107,N_37108,N_37109,N_37110,N_37111,N_37112,N_37113,N_37114,N_37115,N_37116,N_37117,N_37118,N_37119,N_37120,N_37121,N_37122,N_37123,N_37124,N_37125,N_37126,N_37127,N_37128,N_37129,N_37130,N_37131,N_37132,N_37133,N_37134,N_37135,N_37136,N_37137,N_37138,N_37139,N_37140,N_37141,N_37142,N_37143,N_37144,N_37145,N_37146,N_37147,N_37148,N_37149,N_37150,N_37151,N_37152,N_37153,N_37154,N_37155,N_37156,N_37157,N_37158,N_37159,N_37160,N_37161,N_37162,N_37163,N_37164,N_37165,N_37166,N_37167,N_37168,N_37169,N_37170,N_37171,N_37172,N_37173,N_37174,N_37175,N_37176,N_37177,N_37178,N_37179,N_37180,N_37181,N_37182,N_37183,N_37184,N_37185,N_37186,N_37187,N_37188,N_37189,N_37190,N_37191,N_37192,N_37193,N_37194,N_37195,N_37196,N_37197,N_37198,N_37199,N_37200,N_37201,N_37202,N_37203,N_37204,N_37205,N_37206,N_37207,N_37208,N_37209,N_37210,N_37211,N_37212,N_37213,N_37214,N_37215,N_37216,N_37217,N_37218,N_37219,N_37220,N_37221,N_37222,N_37223,N_37224,N_37225,N_37226,N_37227,N_37228,N_37229,N_37230,N_37231,N_37232,N_37233,N_37234,N_37235,N_37236,N_37237,N_37238,N_37239,N_37240,N_37241,N_37242,N_37243,N_37244,N_37245,N_37246,N_37247,N_37248,N_37249,N_37250,N_37251,N_37252,N_37253,N_37254,N_37255,N_37256,N_37257,N_37258,N_37259,N_37260,N_37261,N_37262,N_37263,N_37264,N_37265,N_37266,N_37267,N_37268,N_37269,N_37270,N_37271,N_37272,N_37273,N_37274,N_37275,N_37276,N_37277,N_37278,N_37279,N_37280,N_37281,N_37282,N_37283,N_37284,N_37285,N_37286,N_37287,N_37288,N_37289,N_37290,N_37291,N_37292,N_37293,N_37294,N_37295,N_37296,N_37297,N_37298,N_37299,N_37300,N_37301,N_37302,N_37303,N_37304,N_37305,N_37306,N_37307,N_37308,N_37309,N_37310,N_37311,N_37312,N_37313,N_37314,N_37315,N_37316,N_37317,N_37318,N_37319,N_37320,N_37321,N_37322,N_37323,N_37324,N_37325,N_37326,N_37327,N_37328,N_37329,N_37330,N_37331,N_37332,N_37333,N_37334,N_37335,N_37336,N_37337,N_37338,N_37339,N_37340,N_37341,N_37342,N_37343,N_37344,N_37345,N_37346,N_37347,N_37348,N_37349,N_37350,N_37351,N_37352,N_37353,N_37354,N_37355,N_37356,N_37357,N_37358,N_37359,N_37360,N_37361,N_37362,N_37363,N_37364,N_37365,N_37366,N_37367,N_37368,N_37369,N_37370,N_37371,N_37372,N_37373,N_37374,N_37375,N_37376,N_37377,N_37378,N_37379,N_37380,N_37381,N_37382,N_37383,N_37384,N_37385,N_37386,N_37387,N_37388,N_37389,N_37390,N_37391,N_37392,N_37393,N_37394,N_37395,N_37396,N_37397,N_37398,N_37399,N_37400,N_37401,N_37402,N_37403,N_37404,N_37405,N_37406,N_37407,N_37408,N_37409,N_37410,N_37411,N_37412,N_37413,N_37414,N_37415,N_37416,N_37417,N_37418,N_37419,N_37420,N_37421,N_37422,N_37423,N_37424,N_37425,N_37426,N_37427,N_37428,N_37429,N_37430,N_37431,N_37432,N_37433,N_37434,N_37435,N_37436,N_37437,N_37438,N_37439,N_37440,N_37441,N_37442,N_37443,N_37444,N_37445,N_37446,N_37447,N_37448,N_37449,N_37450,N_37451,N_37452,N_37453,N_37454,N_37455,N_37456,N_37457,N_37458,N_37459,N_37460,N_37461,N_37462,N_37463,N_37464,N_37465,N_37466,N_37467,N_37468,N_37469,N_37470,N_37471,N_37472,N_37473,N_37474,N_37475,N_37476,N_37477,N_37478,N_37479,N_37480,N_37481,N_37482,N_37483,N_37484,N_37485,N_37486,N_37487,N_37488,N_37489,N_37490,N_37491,N_37492,N_37493,N_37494,N_37495,N_37496,N_37497,N_37498,N_37499,N_37500,N_37501,N_37502,N_37503,N_37504,N_37505,N_37506,N_37507,N_37508,N_37509,N_37510,N_37511,N_37512,N_37513,N_37514,N_37515,N_37516,N_37517,N_37518,N_37519,N_37520,N_37521,N_37522,N_37523,N_37524,N_37525,N_37526,N_37527,N_37528,N_37529,N_37530,N_37531,N_37532,N_37533,N_37534,N_37535,N_37536,N_37537,N_37538,N_37539,N_37540,N_37541,N_37542,N_37543,N_37544,N_37545,N_37546,N_37547,N_37548,N_37549,N_37550,N_37551,N_37552,N_37553,N_37554,N_37555,N_37556,N_37557,N_37558,N_37559,N_37560,N_37561,N_37562,N_37563,N_37564,N_37565,N_37566,N_37567,N_37568,N_37569,N_37570,N_37571,N_37572,N_37573,N_37574,N_37575,N_37576,N_37577,N_37578,N_37579,N_37580,N_37581,N_37582,N_37583,N_37584,N_37585,N_37586,N_37587,N_37588,N_37589,N_37590,N_37591,N_37592,N_37593,N_37594,N_37595,N_37596,N_37597,N_37598,N_37599,N_37600,N_37601,N_37602,N_37603,N_37604,N_37605,N_37606,N_37607,N_37608,N_37609,N_37610,N_37611,N_37612,N_37613,N_37614,N_37615,N_37616,N_37617,N_37618,N_37619,N_37620,N_37621,N_37622,N_37623,N_37624,N_37625,N_37626,N_37627,N_37628,N_37629,N_37630,N_37631,N_37632,N_37633,N_37634,N_37635,N_37636,N_37637,N_37638,N_37639,N_37640,N_37641,N_37642,N_37643,N_37644,N_37645,N_37646,N_37647,N_37648,N_37649,N_37650,N_37651,N_37652,N_37653,N_37654,N_37655,N_37656,N_37657,N_37658,N_37659,N_37660,N_37661,N_37662,N_37663,N_37664,N_37665,N_37666,N_37667,N_37668,N_37669,N_37670,N_37671,N_37672,N_37673,N_37674,N_37675,N_37676,N_37677,N_37678,N_37679,N_37680,N_37681,N_37682,N_37683,N_37684,N_37685,N_37686,N_37687,N_37688,N_37689,N_37690,N_37691,N_37692,N_37693,N_37694,N_37695,N_37696,N_37697,N_37698,N_37699,N_37700,N_37701,N_37702,N_37703,N_37704,N_37705,N_37706,N_37707,N_37708,N_37709,N_37710,N_37711,N_37712,N_37713,N_37714,N_37715,N_37716,N_37717,N_37718,N_37719,N_37720,N_37721,N_37722,N_37723,N_37724,N_37725,N_37726,N_37727,N_37728,N_37729,N_37730,N_37731,N_37732,N_37733,N_37734,N_37735,N_37736,N_37737,N_37738,N_37739,N_37740,N_37741,N_37742,N_37743,N_37744,N_37745,N_37746,N_37747,N_37748,N_37749,N_37750,N_37751,N_37752,N_37753,N_37754,N_37755,N_37756,N_37757,N_37758,N_37759,N_37760,N_37761,N_37762,N_37763,N_37764,N_37765,N_37766,N_37767,N_37768,N_37769,N_37770,N_37771,N_37772,N_37773,N_37774,N_37775,N_37776,N_37777,N_37778,N_37779,N_37780,N_37781,N_37782,N_37783,N_37784,N_37785,N_37786,N_37787,N_37788,N_37789,N_37790,N_37791,N_37792,N_37793,N_37794,N_37795,N_37796,N_37797,N_37798,N_37799,N_37800,N_37801,N_37802,N_37803,N_37804,N_37805,N_37806,N_37807,N_37808,N_37809,N_37810,N_37811,N_37812,N_37813,N_37814,N_37815,N_37816,N_37817,N_37818,N_37819,N_37820,N_37821,N_37822,N_37823,N_37824,N_37825,N_37826,N_37827,N_37828,N_37829,N_37830,N_37831,N_37832,N_37833,N_37834,N_37835,N_37836,N_37837,N_37838,N_37839,N_37840,N_37841,N_37842,N_37843,N_37844,N_37845,N_37846,N_37847,N_37848,N_37849,N_37850,N_37851,N_37852,N_37853,N_37854,N_37855,N_37856,N_37857,N_37858,N_37859,N_37860,N_37861,N_37862,N_37863,N_37864,N_37865,N_37866,N_37867,N_37868,N_37869,N_37870,N_37871,N_37872,N_37873,N_37874,N_37875,N_37876,N_37877,N_37878,N_37879,N_37880,N_37881,N_37882,N_37883,N_37884,N_37885,N_37886,N_37887,N_37888,N_37889,N_37890,N_37891,N_37892,N_37893,N_37894,N_37895,N_37896,N_37897,N_37898,N_37899,N_37900,N_37901,N_37902,N_37903,N_37904,N_37905,N_37906,N_37907,N_37908,N_37909,N_37910,N_37911,N_37912,N_37913,N_37914,N_37915,N_37916,N_37917,N_37918,N_37919,N_37920,N_37921,N_37922,N_37923,N_37924,N_37925,N_37926,N_37927,N_37928,N_37929,N_37930,N_37931,N_37932,N_37933,N_37934,N_37935,N_37936,N_37937,N_37938,N_37939,N_37940,N_37941,N_37942,N_37943,N_37944,N_37945,N_37946,N_37947,N_37948,N_37949,N_37950,N_37951,N_37952,N_37953,N_37954,N_37955,N_37956,N_37957,N_37958,N_37959,N_37960,N_37961,N_37962,N_37963,N_37964,N_37965,N_37966,N_37967,N_37968,N_37969,N_37970,N_37971,N_37972,N_37973,N_37974,N_37975,N_37976,N_37977,N_37978,N_37979,N_37980,N_37981,N_37982,N_37983,N_37984,N_37985,N_37986,N_37987,N_37988,N_37989,N_37990,N_37991,N_37992,N_37993,N_37994,N_37995,N_37996,N_37997,N_37998,N_37999,N_38000,N_38001,N_38002,N_38003,N_38004,N_38005,N_38006,N_38007,N_38008,N_38009,N_38010,N_38011,N_38012,N_38013,N_38014,N_38015,N_38016,N_38017,N_38018,N_38019,N_38020,N_38021,N_38022,N_38023,N_38024,N_38025,N_38026,N_38027,N_38028,N_38029,N_38030,N_38031,N_38032,N_38033,N_38034,N_38035,N_38036,N_38037,N_38038,N_38039,N_38040,N_38041,N_38042,N_38043,N_38044,N_38045,N_38046,N_38047,N_38048,N_38049,N_38050,N_38051,N_38052,N_38053,N_38054,N_38055,N_38056,N_38057,N_38058,N_38059,N_38060,N_38061,N_38062,N_38063,N_38064,N_38065,N_38066,N_38067,N_38068,N_38069,N_38070,N_38071,N_38072,N_38073,N_38074,N_38075,N_38076,N_38077,N_38078,N_38079,N_38080,N_38081,N_38082,N_38083,N_38084,N_38085,N_38086,N_38087,N_38088,N_38089,N_38090,N_38091,N_38092,N_38093,N_38094,N_38095,N_38096,N_38097,N_38098,N_38099,N_38100,N_38101,N_38102,N_38103,N_38104,N_38105,N_38106,N_38107,N_38108,N_38109,N_38110,N_38111,N_38112,N_38113,N_38114,N_38115,N_38116,N_38117,N_38118,N_38119,N_38120,N_38121,N_38122,N_38123,N_38124,N_38125,N_38126,N_38127,N_38128,N_38129,N_38130,N_38131,N_38132,N_38133,N_38134,N_38135,N_38136,N_38137,N_38138,N_38139,N_38140,N_38141,N_38142,N_38143,N_38144,N_38145,N_38146,N_38147,N_38148,N_38149,N_38150,N_38151,N_38152,N_38153,N_38154,N_38155,N_38156,N_38157,N_38158,N_38159,N_38160,N_38161,N_38162,N_38163,N_38164,N_38165,N_38166,N_38167,N_38168,N_38169,N_38170,N_38171,N_38172,N_38173,N_38174,N_38175,N_38176,N_38177,N_38178,N_38179,N_38180,N_38181,N_38182,N_38183,N_38184,N_38185,N_38186,N_38187,N_38188,N_38189,N_38190,N_38191,N_38192,N_38193,N_38194,N_38195,N_38196,N_38197,N_38198,N_38199,N_38200,N_38201,N_38202,N_38203,N_38204,N_38205,N_38206,N_38207,N_38208,N_38209,N_38210,N_38211,N_38212,N_38213,N_38214,N_38215,N_38216,N_38217,N_38218,N_38219,N_38220,N_38221,N_38222,N_38223,N_38224,N_38225,N_38226,N_38227,N_38228,N_38229,N_38230,N_38231,N_38232,N_38233,N_38234,N_38235,N_38236,N_38237,N_38238,N_38239,N_38240,N_38241,N_38242,N_38243,N_38244,N_38245,N_38246,N_38247,N_38248,N_38249,N_38250,N_38251,N_38252,N_38253,N_38254,N_38255,N_38256,N_38257,N_38258,N_38259,N_38260,N_38261,N_38262,N_38263,N_38264,N_38265,N_38266,N_38267,N_38268,N_38269,N_38270,N_38271,N_38272,N_38273,N_38274,N_38275,N_38276,N_38277,N_38278,N_38279,N_38280,N_38281,N_38282,N_38283,N_38284,N_38285,N_38286,N_38287,N_38288,N_38289,N_38290,N_38291,N_38292,N_38293,N_38294,N_38295,N_38296,N_38297,N_38298,N_38299,N_38300,N_38301,N_38302,N_38303,N_38304,N_38305,N_38306,N_38307,N_38308,N_38309,N_38310,N_38311,N_38312,N_38313,N_38314,N_38315,N_38316,N_38317,N_38318,N_38319,N_38320,N_38321,N_38322,N_38323,N_38324,N_38325,N_38326,N_38327,N_38328,N_38329,N_38330,N_38331,N_38332,N_38333,N_38334,N_38335,N_38336,N_38337,N_38338,N_38339,N_38340,N_38341,N_38342,N_38343,N_38344,N_38345,N_38346,N_38347,N_38348,N_38349,N_38350,N_38351,N_38352,N_38353,N_38354,N_38355,N_38356,N_38357,N_38358,N_38359,N_38360,N_38361,N_38362,N_38363,N_38364,N_38365,N_38366,N_38367,N_38368,N_38369,N_38370,N_38371,N_38372,N_38373,N_38374,N_38375,N_38376,N_38377,N_38378,N_38379,N_38380,N_38381,N_38382,N_38383,N_38384,N_38385,N_38386,N_38387,N_38388,N_38389,N_38390,N_38391,N_38392,N_38393,N_38394,N_38395,N_38396,N_38397,N_38398,N_38399,N_38400,N_38401,N_38402,N_38403,N_38404,N_38405,N_38406,N_38407,N_38408,N_38409,N_38410,N_38411,N_38412,N_38413,N_38414,N_38415,N_38416,N_38417,N_38418,N_38419,N_38420,N_38421,N_38422,N_38423,N_38424,N_38425,N_38426,N_38427,N_38428,N_38429,N_38430,N_38431,N_38432,N_38433,N_38434,N_38435,N_38436,N_38437,N_38438,N_38439,N_38440,N_38441,N_38442,N_38443,N_38444,N_38445,N_38446,N_38447,N_38448,N_38449,N_38450,N_38451,N_38452,N_38453,N_38454,N_38455,N_38456,N_38457,N_38458,N_38459,N_38460,N_38461,N_38462,N_38463,N_38464,N_38465,N_38466,N_38467,N_38468,N_38469,N_38470,N_38471,N_38472,N_38473,N_38474,N_38475,N_38476,N_38477,N_38478,N_38479,N_38480,N_38481,N_38482,N_38483,N_38484,N_38485,N_38486,N_38487,N_38488,N_38489,N_38490,N_38491,N_38492,N_38493,N_38494,N_38495,N_38496,N_38497,N_38498,N_38499,N_38500,N_38501,N_38502,N_38503,N_38504,N_38505,N_38506,N_38507,N_38508,N_38509,N_38510,N_38511,N_38512,N_38513,N_38514,N_38515,N_38516,N_38517,N_38518,N_38519,N_38520,N_38521,N_38522,N_38523,N_38524,N_38525,N_38526,N_38527,N_38528,N_38529,N_38530,N_38531,N_38532,N_38533,N_38534,N_38535,N_38536,N_38537,N_38538,N_38539,N_38540,N_38541,N_38542,N_38543,N_38544,N_38545,N_38546,N_38547,N_38548,N_38549,N_38550,N_38551,N_38552,N_38553,N_38554,N_38555,N_38556,N_38557,N_38558,N_38559,N_38560,N_38561,N_38562,N_38563,N_38564,N_38565,N_38566,N_38567,N_38568,N_38569,N_38570,N_38571,N_38572,N_38573,N_38574,N_38575,N_38576,N_38577,N_38578,N_38579,N_38580,N_38581,N_38582,N_38583,N_38584,N_38585,N_38586,N_38587,N_38588,N_38589,N_38590,N_38591,N_38592,N_38593,N_38594,N_38595,N_38596,N_38597,N_38598,N_38599,N_38600,N_38601,N_38602,N_38603,N_38604,N_38605,N_38606,N_38607,N_38608,N_38609,N_38610,N_38611,N_38612,N_38613,N_38614,N_38615,N_38616,N_38617,N_38618,N_38619,N_38620,N_38621,N_38622,N_38623,N_38624,N_38625,N_38626,N_38627,N_38628,N_38629,N_38630,N_38631,N_38632,N_38633,N_38634,N_38635,N_38636,N_38637,N_38638,N_38639,N_38640,N_38641,N_38642,N_38643,N_38644,N_38645,N_38646,N_38647,N_38648,N_38649,N_38650,N_38651,N_38652,N_38653,N_38654,N_38655,N_38656,N_38657,N_38658,N_38659,N_38660,N_38661,N_38662,N_38663,N_38664,N_38665,N_38666,N_38667,N_38668,N_38669,N_38670,N_38671,N_38672,N_38673,N_38674,N_38675,N_38676,N_38677,N_38678,N_38679,N_38680,N_38681,N_38682,N_38683,N_38684,N_38685,N_38686,N_38687,N_38688,N_38689,N_38690,N_38691,N_38692,N_38693,N_38694,N_38695,N_38696,N_38697,N_38698,N_38699,N_38700,N_38701,N_38702,N_38703,N_38704,N_38705,N_38706,N_38707,N_38708,N_38709,N_38710,N_38711,N_38712,N_38713,N_38714,N_38715,N_38716,N_38717,N_38718,N_38719,N_38720,N_38721,N_38722,N_38723,N_38724,N_38725,N_38726,N_38727,N_38728,N_38729,N_38730,N_38731,N_38732,N_38733,N_38734,N_38735,N_38736,N_38737,N_38738,N_38739,N_38740,N_38741,N_38742,N_38743,N_38744,N_38745,N_38746,N_38747,N_38748,N_38749,N_38750,N_38751,N_38752,N_38753,N_38754,N_38755,N_38756,N_38757,N_38758,N_38759,N_38760,N_38761,N_38762,N_38763,N_38764,N_38765,N_38766,N_38767,N_38768,N_38769,N_38770,N_38771,N_38772,N_38773,N_38774,N_38775,N_38776,N_38777,N_38778,N_38779,N_38780,N_38781,N_38782,N_38783,N_38784,N_38785,N_38786,N_38787,N_38788,N_38789,N_38790,N_38791,N_38792,N_38793,N_38794,N_38795,N_38796,N_38797,N_38798,N_38799,N_38800,N_38801,N_38802,N_38803,N_38804,N_38805,N_38806,N_38807,N_38808,N_38809,N_38810,N_38811,N_38812,N_38813,N_38814,N_38815,N_38816,N_38817,N_38818,N_38819,N_38820,N_38821,N_38822,N_38823,N_38824,N_38825,N_38826,N_38827,N_38828,N_38829,N_38830,N_38831,N_38832,N_38833,N_38834,N_38835,N_38836,N_38837,N_38838,N_38839,N_38840,N_38841,N_38842,N_38843,N_38844,N_38845,N_38846,N_38847,N_38848,N_38849,N_38850,N_38851,N_38852,N_38853,N_38854,N_38855,N_38856,N_38857,N_38858,N_38859,N_38860,N_38861,N_38862,N_38863,N_38864,N_38865,N_38866,N_38867,N_38868,N_38869,N_38870,N_38871,N_38872,N_38873,N_38874,N_38875,N_38876,N_38877,N_38878,N_38879,N_38880,N_38881,N_38882,N_38883,N_38884,N_38885,N_38886,N_38887,N_38888,N_38889,N_38890,N_38891,N_38892,N_38893,N_38894,N_38895,N_38896,N_38897,N_38898,N_38899,N_38900,N_38901,N_38902,N_38903,N_38904,N_38905,N_38906,N_38907,N_38908,N_38909,N_38910,N_38911,N_38912,N_38913,N_38914,N_38915,N_38916,N_38917,N_38918,N_38919,N_38920,N_38921,N_38922,N_38923,N_38924,N_38925,N_38926,N_38927,N_38928,N_38929,N_38930,N_38931,N_38932,N_38933,N_38934,N_38935,N_38936,N_38937,N_38938,N_38939,N_38940,N_38941,N_38942,N_38943,N_38944,N_38945,N_38946,N_38947,N_38948,N_38949,N_38950,N_38951,N_38952,N_38953,N_38954,N_38955,N_38956,N_38957,N_38958,N_38959,N_38960,N_38961,N_38962,N_38963,N_38964,N_38965,N_38966,N_38967,N_38968,N_38969,N_38970,N_38971,N_38972,N_38973,N_38974,N_38975,N_38976,N_38977,N_38978,N_38979,N_38980,N_38981,N_38982,N_38983,N_38984,N_38985,N_38986,N_38987,N_38988,N_38989,N_38990,N_38991,N_38992,N_38993,N_38994,N_38995,N_38996,N_38997,N_38998,N_38999,N_39000,N_39001,N_39002,N_39003,N_39004,N_39005,N_39006,N_39007,N_39008,N_39009,N_39010,N_39011,N_39012,N_39013,N_39014,N_39015,N_39016,N_39017,N_39018,N_39019,N_39020,N_39021,N_39022,N_39023,N_39024,N_39025,N_39026,N_39027,N_39028,N_39029,N_39030,N_39031,N_39032,N_39033,N_39034,N_39035,N_39036,N_39037,N_39038,N_39039,N_39040,N_39041,N_39042,N_39043,N_39044,N_39045,N_39046,N_39047,N_39048,N_39049,N_39050,N_39051,N_39052,N_39053,N_39054,N_39055,N_39056,N_39057,N_39058,N_39059,N_39060,N_39061,N_39062,N_39063,N_39064,N_39065,N_39066,N_39067,N_39068,N_39069,N_39070,N_39071,N_39072,N_39073,N_39074,N_39075,N_39076,N_39077,N_39078,N_39079,N_39080,N_39081,N_39082,N_39083,N_39084,N_39085,N_39086,N_39087,N_39088,N_39089,N_39090,N_39091,N_39092,N_39093,N_39094,N_39095,N_39096,N_39097,N_39098,N_39099,N_39100,N_39101,N_39102,N_39103,N_39104,N_39105,N_39106,N_39107,N_39108,N_39109,N_39110,N_39111,N_39112,N_39113,N_39114,N_39115,N_39116,N_39117,N_39118,N_39119,N_39120,N_39121,N_39122,N_39123,N_39124,N_39125,N_39126,N_39127,N_39128,N_39129,N_39130,N_39131,N_39132,N_39133,N_39134,N_39135,N_39136,N_39137,N_39138,N_39139,N_39140,N_39141,N_39142,N_39143,N_39144,N_39145,N_39146,N_39147,N_39148,N_39149,N_39150,N_39151,N_39152,N_39153,N_39154,N_39155,N_39156,N_39157,N_39158,N_39159,N_39160,N_39161,N_39162,N_39163,N_39164,N_39165,N_39166,N_39167,N_39168,N_39169,N_39170,N_39171,N_39172,N_39173,N_39174,N_39175,N_39176,N_39177,N_39178,N_39179,N_39180,N_39181,N_39182,N_39183,N_39184,N_39185,N_39186,N_39187,N_39188,N_39189,N_39190,N_39191,N_39192,N_39193,N_39194,N_39195,N_39196,N_39197,N_39198,N_39199,N_39200,N_39201,N_39202,N_39203,N_39204,N_39205,N_39206,N_39207,N_39208,N_39209,N_39210,N_39211,N_39212,N_39213,N_39214,N_39215,N_39216,N_39217,N_39218,N_39219,N_39220,N_39221,N_39222,N_39223,N_39224,N_39225,N_39226,N_39227,N_39228,N_39229,N_39230,N_39231,N_39232,N_39233,N_39234,N_39235,N_39236,N_39237,N_39238,N_39239,N_39240,N_39241,N_39242,N_39243,N_39244,N_39245,N_39246,N_39247,N_39248,N_39249,N_39250,N_39251,N_39252,N_39253,N_39254,N_39255,N_39256,N_39257,N_39258,N_39259,N_39260,N_39261,N_39262,N_39263,N_39264,N_39265,N_39266,N_39267,N_39268,N_39269,N_39270,N_39271,N_39272,N_39273,N_39274,N_39275,N_39276,N_39277,N_39278,N_39279,N_39280,N_39281,N_39282,N_39283,N_39284,N_39285,N_39286,N_39287,N_39288,N_39289,N_39290,N_39291,N_39292,N_39293,N_39294,N_39295,N_39296,N_39297,N_39298,N_39299,N_39300,N_39301,N_39302,N_39303,N_39304,N_39305,N_39306,N_39307,N_39308,N_39309,N_39310,N_39311,N_39312,N_39313,N_39314,N_39315,N_39316,N_39317,N_39318,N_39319,N_39320,N_39321,N_39322,N_39323,N_39324,N_39325,N_39326,N_39327,N_39328,N_39329,N_39330,N_39331,N_39332,N_39333,N_39334,N_39335,N_39336,N_39337,N_39338,N_39339,N_39340,N_39341,N_39342,N_39343,N_39344,N_39345,N_39346,N_39347,N_39348,N_39349,N_39350,N_39351,N_39352,N_39353,N_39354,N_39355,N_39356,N_39357,N_39358,N_39359,N_39360,N_39361,N_39362,N_39363,N_39364,N_39365,N_39366,N_39367,N_39368,N_39369,N_39370,N_39371,N_39372,N_39373,N_39374,N_39375,N_39376,N_39377,N_39378,N_39379,N_39380,N_39381,N_39382,N_39383,N_39384,N_39385,N_39386,N_39387,N_39388,N_39389,N_39390,N_39391,N_39392,N_39393,N_39394,N_39395,N_39396,N_39397,N_39398,N_39399,N_39400,N_39401,N_39402,N_39403,N_39404,N_39405,N_39406,N_39407,N_39408,N_39409,N_39410,N_39411,N_39412,N_39413,N_39414,N_39415,N_39416,N_39417,N_39418,N_39419,N_39420,N_39421,N_39422,N_39423,N_39424,N_39425,N_39426,N_39427,N_39428,N_39429,N_39430,N_39431,N_39432,N_39433,N_39434,N_39435,N_39436,N_39437,N_39438,N_39439,N_39440,N_39441,N_39442,N_39443,N_39444,N_39445,N_39446,N_39447,N_39448,N_39449,N_39450,N_39451,N_39452,N_39453,N_39454,N_39455,N_39456,N_39457,N_39458,N_39459,N_39460,N_39461,N_39462,N_39463,N_39464,N_39465,N_39466,N_39467,N_39468,N_39469,N_39470,N_39471,N_39472,N_39473,N_39474,N_39475,N_39476,N_39477,N_39478,N_39479,N_39480,N_39481,N_39482,N_39483,N_39484,N_39485,N_39486,N_39487,N_39488,N_39489,N_39490,N_39491,N_39492,N_39493,N_39494,N_39495,N_39496,N_39497,N_39498,N_39499,N_39500,N_39501,N_39502,N_39503,N_39504,N_39505,N_39506,N_39507,N_39508,N_39509,N_39510,N_39511,N_39512,N_39513,N_39514,N_39515,N_39516,N_39517,N_39518,N_39519,N_39520,N_39521,N_39522,N_39523,N_39524,N_39525,N_39526,N_39527,N_39528,N_39529,N_39530,N_39531,N_39532,N_39533,N_39534,N_39535,N_39536,N_39537,N_39538,N_39539,N_39540,N_39541,N_39542,N_39543,N_39544,N_39545,N_39546,N_39547,N_39548,N_39549,N_39550,N_39551,N_39552,N_39553,N_39554,N_39555,N_39556,N_39557,N_39558,N_39559,N_39560,N_39561,N_39562,N_39563,N_39564,N_39565,N_39566,N_39567,N_39568,N_39569,N_39570,N_39571,N_39572,N_39573,N_39574,N_39575,N_39576,N_39577,N_39578,N_39579,N_39580,N_39581,N_39582,N_39583,N_39584,N_39585,N_39586,N_39587,N_39588,N_39589,N_39590,N_39591,N_39592,N_39593,N_39594,N_39595,N_39596,N_39597,N_39598,N_39599,N_39600,N_39601,N_39602,N_39603,N_39604,N_39605,N_39606,N_39607,N_39608,N_39609,N_39610,N_39611,N_39612,N_39613,N_39614,N_39615,N_39616,N_39617,N_39618,N_39619,N_39620,N_39621,N_39622,N_39623,N_39624,N_39625,N_39626,N_39627,N_39628,N_39629,N_39630,N_39631,N_39632,N_39633,N_39634,N_39635,N_39636,N_39637,N_39638,N_39639,N_39640,N_39641,N_39642,N_39643,N_39644,N_39645,N_39646,N_39647,N_39648,N_39649,N_39650,N_39651,N_39652,N_39653,N_39654,N_39655,N_39656,N_39657,N_39658,N_39659,N_39660,N_39661,N_39662,N_39663,N_39664,N_39665,N_39666,N_39667,N_39668,N_39669,N_39670,N_39671,N_39672,N_39673,N_39674,N_39675,N_39676,N_39677,N_39678,N_39679,N_39680,N_39681,N_39682,N_39683,N_39684,N_39685,N_39686,N_39687,N_39688,N_39689,N_39690,N_39691,N_39692,N_39693,N_39694,N_39695,N_39696,N_39697,N_39698,N_39699,N_39700,N_39701,N_39702,N_39703,N_39704,N_39705,N_39706,N_39707,N_39708,N_39709,N_39710,N_39711,N_39712,N_39713,N_39714,N_39715,N_39716,N_39717,N_39718,N_39719,N_39720,N_39721,N_39722,N_39723,N_39724,N_39725,N_39726,N_39727,N_39728,N_39729,N_39730,N_39731,N_39732,N_39733,N_39734,N_39735,N_39736,N_39737,N_39738,N_39739,N_39740,N_39741,N_39742,N_39743,N_39744,N_39745,N_39746,N_39747,N_39748,N_39749,N_39750,N_39751,N_39752,N_39753,N_39754,N_39755,N_39756,N_39757,N_39758,N_39759,N_39760,N_39761,N_39762,N_39763,N_39764,N_39765,N_39766,N_39767,N_39768,N_39769,N_39770,N_39771,N_39772,N_39773,N_39774,N_39775,N_39776,N_39777,N_39778,N_39779,N_39780,N_39781,N_39782,N_39783,N_39784,N_39785,N_39786,N_39787,N_39788,N_39789,N_39790,N_39791,N_39792,N_39793,N_39794,N_39795,N_39796,N_39797,N_39798,N_39799,N_39800,N_39801,N_39802,N_39803,N_39804,N_39805,N_39806,N_39807,N_39808,N_39809,N_39810,N_39811,N_39812,N_39813,N_39814,N_39815,N_39816,N_39817,N_39818,N_39819,N_39820,N_39821,N_39822,N_39823,N_39824,N_39825,N_39826,N_39827,N_39828,N_39829,N_39830,N_39831,N_39832,N_39833,N_39834,N_39835,N_39836,N_39837,N_39838,N_39839,N_39840,N_39841,N_39842,N_39843,N_39844,N_39845,N_39846,N_39847,N_39848,N_39849,N_39850,N_39851,N_39852,N_39853,N_39854,N_39855,N_39856,N_39857,N_39858,N_39859,N_39860,N_39861,N_39862,N_39863,N_39864,N_39865,N_39866,N_39867,N_39868,N_39869,N_39870,N_39871,N_39872,N_39873,N_39874,N_39875,N_39876,N_39877,N_39878,N_39879,N_39880,N_39881,N_39882,N_39883,N_39884,N_39885,N_39886,N_39887,N_39888,N_39889,N_39890,N_39891,N_39892,N_39893,N_39894,N_39895,N_39896,N_39897,N_39898,N_39899,N_39900,N_39901,N_39902,N_39903,N_39904,N_39905,N_39906,N_39907,N_39908,N_39909,N_39910,N_39911,N_39912,N_39913,N_39914,N_39915,N_39916,N_39917,N_39918,N_39919,N_39920,N_39921,N_39922,N_39923,N_39924,N_39925,N_39926,N_39927,N_39928,N_39929,N_39930,N_39931,N_39932,N_39933,N_39934,N_39935,N_39936,N_39937,N_39938,N_39939,N_39940,N_39941,N_39942,N_39943,N_39944,N_39945,N_39946,N_39947,N_39948,N_39949,N_39950,N_39951,N_39952,N_39953,N_39954,N_39955,N_39956,N_39957,N_39958,N_39959,N_39960,N_39961,N_39962,N_39963,N_39964,N_39965,N_39966,N_39967,N_39968,N_39969,N_39970,N_39971,N_39972,N_39973,N_39974,N_39975,N_39976,N_39977,N_39978,N_39979,N_39980,N_39981,N_39982,N_39983,N_39984,N_39985,N_39986,N_39987,N_39988,N_39989,N_39990,N_39991,N_39992,N_39993,N_39994,N_39995,N_39996,N_39997,N_39998,N_39999,N_40000,N_40001,N_40002,N_40003,N_40004,N_40005,N_40006,N_40007,N_40008,N_40009,N_40010,N_40011,N_40012,N_40013,N_40014,N_40015,N_40016,N_40017,N_40018,N_40019,N_40020,N_40021,N_40022,N_40023,N_40024,N_40025,N_40026,N_40027,N_40028,N_40029,N_40030,N_40031,N_40032,N_40033,N_40034,N_40035,N_40036,N_40037,N_40038,N_40039,N_40040,N_40041,N_40042,N_40043,N_40044,N_40045,N_40046,N_40047,N_40048,N_40049,N_40050,N_40051,N_40052,N_40053,N_40054,N_40055,N_40056,N_40057,N_40058,N_40059,N_40060,N_40061,N_40062,N_40063,N_40064,N_40065,N_40066,N_40067,N_40068,N_40069,N_40070,N_40071,N_40072,N_40073,N_40074,N_40075,N_40076,N_40077,N_40078,N_40079,N_40080,N_40081,N_40082,N_40083,N_40084,N_40085,N_40086,N_40087,N_40088,N_40089,N_40090,N_40091,N_40092,N_40093,N_40094,N_40095,N_40096,N_40097,N_40098,N_40099,N_40100,N_40101,N_40102,N_40103,N_40104,N_40105,N_40106,N_40107,N_40108,N_40109,N_40110,N_40111,N_40112,N_40113,N_40114,N_40115,N_40116,N_40117,N_40118,N_40119,N_40120,N_40121,N_40122,N_40123,N_40124,N_40125,N_40126,N_40127,N_40128,N_40129,N_40130,N_40131,N_40132,N_40133,N_40134,N_40135,N_40136,N_40137,N_40138,N_40139,N_40140,N_40141,N_40142,N_40143,N_40144,N_40145,N_40146,N_40147,N_40148,N_40149,N_40150,N_40151,N_40152,N_40153,N_40154,N_40155,N_40156,N_40157,N_40158,N_40159,N_40160,N_40161,N_40162,N_40163,N_40164,N_40165,N_40166,N_40167,N_40168,N_40169,N_40170,N_40171,N_40172,N_40173,N_40174,N_40175,N_40176,N_40177,N_40178,N_40179,N_40180,N_40181,N_40182,N_40183,N_40184,N_40185,N_40186,N_40187,N_40188,N_40189,N_40190,N_40191,N_40192,N_40193,N_40194,N_40195,N_40196,N_40197,N_40198,N_40199,N_40200,N_40201,N_40202,N_40203,N_40204,N_40205,N_40206,N_40207,N_40208,N_40209,N_40210,N_40211,N_40212,N_40213,N_40214,N_40215,N_40216,N_40217,N_40218,N_40219,N_40220,N_40221,N_40222,N_40223,N_40224,N_40225,N_40226,N_40227,N_40228,N_40229,N_40230,N_40231,N_40232,N_40233,N_40234,N_40235,N_40236,N_40237,N_40238,N_40239,N_40240,N_40241,N_40242,N_40243,N_40244,N_40245,N_40246,N_40247,N_40248,N_40249,N_40250,N_40251,N_40252,N_40253,N_40254,N_40255,N_40256,N_40257,N_40258,N_40259,N_40260,N_40261,N_40262,N_40263,N_40264,N_40265,N_40266,N_40267,N_40268,N_40269,N_40270,N_40271,N_40272,N_40273,N_40274,N_40275,N_40276,N_40277,N_40278,N_40279,N_40280,N_40281,N_40282,N_40283,N_40284,N_40285,N_40286,N_40287,N_40288,N_40289,N_40290,N_40291,N_40292,N_40293,N_40294,N_40295,N_40296,N_40297,N_40298,N_40299,N_40300,N_40301,N_40302,N_40303,N_40304,N_40305,N_40306,N_40307,N_40308,N_40309,N_40310,N_40311,N_40312,N_40313,N_40314,N_40315,N_40316,N_40317,N_40318,N_40319,N_40320,N_40321,N_40322,N_40323,N_40324,N_40325,N_40326,N_40327,N_40328,N_40329,N_40330,N_40331,N_40332,N_40333,N_40334,N_40335,N_40336,N_40337,N_40338,N_40339,N_40340,N_40341,N_40342,N_40343,N_40344,N_40345,N_40346,N_40347,N_40348,N_40349,N_40350,N_40351,N_40352,N_40353,N_40354,N_40355,N_40356,N_40357,N_40358,N_40359,N_40360,N_40361,N_40362,N_40363,N_40364,N_40365,N_40366,N_40367,N_40368,N_40369,N_40370,N_40371,N_40372,N_40373,N_40374,N_40375,N_40376,N_40377,N_40378,N_40379,N_40380,N_40381,N_40382,N_40383,N_40384,N_40385,N_40386,N_40387,N_40388,N_40389,N_40390,N_40391,N_40392,N_40393,N_40394,N_40395,N_40396,N_40397,N_40398,N_40399,N_40400,N_40401,N_40402,N_40403,N_40404,N_40405,N_40406,N_40407,N_40408,N_40409,N_40410,N_40411,N_40412,N_40413,N_40414,N_40415,N_40416,N_40417,N_40418,N_40419,N_40420,N_40421,N_40422,N_40423,N_40424,N_40425,N_40426,N_40427,N_40428,N_40429,N_40430,N_40431,N_40432,N_40433,N_40434,N_40435,N_40436,N_40437,N_40438,N_40439,N_40440,N_40441,N_40442,N_40443,N_40444,N_40445,N_40446,N_40447,N_40448,N_40449,N_40450,N_40451,N_40452,N_40453,N_40454,N_40455,N_40456,N_40457,N_40458,N_40459,N_40460,N_40461,N_40462,N_40463,N_40464,N_40465,N_40466,N_40467,N_40468,N_40469,N_40470,N_40471,N_40472,N_40473,N_40474,N_40475,N_40476,N_40477,N_40478,N_40479,N_40480,N_40481,N_40482,N_40483,N_40484,N_40485,N_40486,N_40487,N_40488,N_40489,N_40490,N_40491,N_40492,N_40493,N_40494,N_40495,N_40496,N_40497,N_40498,N_40499,N_40500,N_40501,N_40502,N_40503,N_40504,N_40505,N_40506,N_40507,N_40508,N_40509,N_40510,N_40511,N_40512,N_40513,N_40514,N_40515,N_40516,N_40517,N_40518,N_40519,N_40520,N_40521,N_40522,N_40523,N_40524,N_40525,N_40526,N_40527,N_40528,N_40529,N_40530,N_40531,N_40532,N_40533,N_40534,N_40535,N_40536,N_40537,N_40538,N_40539,N_40540,N_40541,N_40542,N_40543,N_40544,N_40545,N_40546,N_40547,N_40548,N_40549,N_40550,N_40551,N_40552,N_40553,N_40554,N_40555,N_40556,N_40557,N_40558,N_40559,N_40560,N_40561,N_40562,N_40563,N_40564,N_40565,N_40566,N_40567,N_40568,N_40569,N_40570,N_40571,N_40572,N_40573,N_40574,N_40575,N_40576,N_40577,N_40578,N_40579,N_40580,N_40581,N_40582,N_40583,N_40584,N_40585,N_40586,N_40587,N_40588,N_40589,N_40590,N_40591,N_40592,N_40593,N_40594,N_40595,N_40596,N_40597,N_40598,N_40599,N_40600,N_40601,N_40602,N_40603,N_40604,N_40605,N_40606,N_40607,N_40608,N_40609,N_40610,N_40611,N_40612,N_40613,N_40614,N_40615,N_40616,N_40617,N_40618,N_40619,N_40620,N_40621,N_40622,N_40623,N_40624,N_40625,N_40626,N_40627,N_40628,N_40629,N_40630,N_40631,N_40632,N_40633,N_40634,N_40635,N_40636,N_40637,N_40638,N_40639,N_40640,N_40641,N_40642,N_40643,N_40644,N_40645,N_40646,N_40647,N_40648,N_40649,N_40650,N_40651,N_40652,N_40653,N_40654,N_40655,N_40656,N_40657,N_40658,N_40659,N_40660,N_40661,N_40662,N_40663,N_40664,N_40665,N_40666,N_40667,N_40668,N_40669,N_40670,N_40671,N_40672,N_40673,N_40674,N_40675,N_40676,N_40677,N_40678,N_40679,N_40680,N_40681,N_40682,N_40683,N_40684,N_40685,N_40686,N_40687,N_40688,N_40689,N_40690,N_40691,N_40692,N_40693,N_40694,N_40695,N_40696,N_40697,N_40698,N_40699,N_40700,N_40701,N_40702,N_40703,N_40704,N_40705,N_40706,N_40707,N_40708,N_40709,N_40710,N_40711,N_40712,N_40713,N_40714,N_40715,N_40716,N_40717,N_40718,N_40719,N_40720,N_40721,N_40722,N_40723,N_40724,N_40725,N_40726,N_40727,N_40728,N_40729,N_40730,N_40731,N_40732,N_40733,N_40734,N_40735,N_40736,N_40737,N_40738,N_40739,N_40740,N_40741,N_40742,N_40743,N_40744,N_40745,N_40746,N_40747,N_40748,N_40749,N_40750,N_40751,N_40752,N_40753,N_40754,N_40755,N_40756,N_40757,N_40758,N_40759,N_40760,N_40761,N_40762,N_40763,N_40764,N_40765,N_40766,N_40767,N_40768,N_40769,N_40770,N_40771,N_40772,N_40773,N_40774,N_40775,N_40776,N_40777,N_40778,N_40779,N_40780,N_40781,N_40782,N_40783,N_40784,N_40785,N_40786,N_40787,N_40788,N_40789,N_40790,N_40791,N_40792,N_40793,N_40794,N_40795,N_40796,N_40797,N_40798,N_40799,N_40800,N_40801,N_40802,N_40803,N_40804,N_40805,N_40806,N_40807,N_40808,N_40809,N_40810,N_40811,N_40812,N_40813,N_40814,N_40815,N_40816,N_40817,N_40818,N_40819,N_40820,N_40821,N_40822,N_40823,N_40824,N_40825,N_40826,N_40827,N_40828,N_40829,N_40830,N_40831,N_40832,N_40833,N_40834,N_40835,N_40836,N_40837,N_40838,N_40839,N_40840,N_40841,N_40842,N_40843,N_40844,N_40845,N_40846,N_40847,N_40848,N_40849,N_40850,N_40851,N_40852,N_40853,N_40854,N_40855,N_40856,N_40857,N_40858,N_40859,N_40860,N_40861,N_40862,N_40863,N_40864,N_40865,N_40866,N_40867,N_40868,N_40869,N_40870,N_40871,N_40872,N_40873,N_40874,N_40875,N_40876,N_40877,N_40878,N_40879,N_40880,N_40881,N_40882,N_40883,N_40884,N_40885,N_40886,N_40887,N_40888,N_40889,N_40890,N_40891,N_40892,N_40893,N_40894,N_40895,N_40896,N_40897,N_40898,N_40899,N_40900,N_40901,N_40902,N_40903,N_40904,N_40905,N_40906,N_40907,N_40908,N_40909,N_40910,N_40911,N_40912,N_40913,N_40914,N_40915,N_40916,N_40917,N_40918,N_40919,N_40920,N_40921,N_40922,N_40923,N_40924,N_40925,N_40926,N_40927,N_40928,N_40929,N_40930,N_40931,N_40932,N_40933,N_40934,N_40935,N_40936,N_40937,N_40938,N_40939,N_40940,N_40941,N_40942,N_40943,N_40944,N_40945,N_40946,N_40947,N_40948,N_40949,N_40950,N_40951,N_40952,N_40953,N_40954,N_40955,N_40956,N_40957,N_40958,N_40959,N_40960,N_40961,N_40962,N_40963,N_40964,N_40965,N_40966,N_40967,N_40968,N_40969,N_40970,N_40971,N_40972,N_40973,N_40974,N_40975,N_40976,N_40977,N_40978,N_40979,N_40980,N_40981,N_40982,N_40983,N_40984,N_40985,N_40986,N_40987,N_40988,N_40989,N_40990,N_40991,N_40992,N_40993,N_40994,N_40995,N_40996,N_40997,N_40998,N_40999,N_41000,N_41001,N_41002,N_41003,N_41004,N_41005,N_41006,N_41007,N_41008,N_41009,N_41010,N_41011,N_41012,N_41013,N_41014,N_41015,N_41016,N_41017,N_41018,N_41019,N_41020,N_41021,N_41022,N_41023,N_41024,N_41025,N_41026,N_41027,N_41028,N_41029,N_41030,N_41031,N_41032,N_41033,N_41034,N_41035,N_41036,N_41037,N_41038,N_41039,N_41040,N_41041,N_41042,N_41043,N_41044,N_41045,N_41046,N_41047,N_41048,N_41049,N_41050,N_41051,N_41052,N_41053,N_41054,N_41055,N_41056,N_41057,N_41058,N_41059,N_41060,N_41061,N_41062,N_41063,N_41064,N_41065,N_41066,N_41067,N_41068,N_41069,N_41070,N_41071,N_41072,N_41073,N_41074,N_41075,N_41076,N_41077,N_41078,N_41079,N_41080,N_41081,N_41082,N_41083,N_41084,N_41085,N_41086,N_41087,N_41088,N_41089,N_41090,N_41091,N_41092,N_41093,N_41094,N_41095,N_41096,N_41097,N_41098,N_41099,N_41100,N_41101,N_41102,N_41103,N_41104,N_41105,N_41106,N_41107,N_41108,N_41109,N_41110,N_41111,N_41112,N_41113,N_41114,N_41115,N_41116,N_41117,N_41118,N_41119,N_41120,N_41121,N_41122,N_41123,N_41124,N_41125,N_41126,N_41127,N_41128,N_41129,N_41130,N_41131,N_41132,N_41133,N_41134,N_41135,N_41136,N_41137,N_41138,N_41139,N_41140,N_41141,N_41142,N_41143,N_41144,N_41145,N_41146,N_41147,N_41148,N_41149,N_41150,N_41151,N_41152,N_41153,N_41154,N_41155,N_41156,N_41157,N_41158,N_41159,N_41160,N_41161,N_41162,N_41163,N_41164,N_41165,N_41166,N_41167,N_41168,N_41169,N_41170,N_41171,N_41172,N_41173,N_41174,N_41175,N_41176,N_41177,N_41178,N_41179,N_41180,N_41181,N_41182,N_41183,N_41184,N_41185,N_41186,N_41187,N_41188,N_41189,N_41190,N_41191,N_41192,N_41193,N_41194,N_41195,N_41196,N_41197,N_41198,N_41199,N_41200,N_41201,N_41202,N_41203,N_41204,N_41205,N_41206,N_41207,N_41208,N_41209,N_41210,N_41211,N_41212,N_41213,N_41214,N_41215,N_41216,N_41217,N_41218,N_41219,N_41220,N_41221,N_41222,N_41223,N_41224,N_41225,N_41226,N_41227,N_41228,N_41229,N_41230,N_41231,N_41232,N_41233,N_41234,N_41235,N_41236,N_41237,N_41238,N_41239,N_41240,N_41241,N_41242,N_41243,N_41244,N_41245,N_41246,N_41247,N_41248,N_41249,N_41250,N_41251,N_41252,N_41253,N_41254,N_41255,N_41256,N_41257,N_41258,N_41259,N_41260,N_41261,N_41262,N_41263,N_41264,N_41265,N_41266,N_41267,N_41268,N_41269,N_41270,N_41271,N_41272,N_41273,N_41274,N_41275,N_41276,N_41277,N_41278,N_41279,N_41280,N_41281,N_41282,N_41283,N_41284,N_41285,N_41286,N_41287,N_41288,N_41289,N_41290,N_41291,N_41292,N_41293,N_41294,N_41295,N_41296,N_41297,N_41298,N_41299,N_41300,N_41301,N_41302,N_41303,N_41304,N_41305,N_41306,N_41307,N_41308,N_41309,N_41310,N_41311,N_41312,N_41313,N_41314,N_41315,N_41316,N_41317,N_41318,N_41319,N_41320,N_41321,N_41322,N_41323,N_41324,N_41325,N_41326,N_41327,N_41328,N_41329,N_41330,N_41331,N_41332,N_41333,N_41334,N_41335,N_41336,N_41337,N_41338,N_41339,N_41340,N_41341,N_41342,N_41343,N_41344,N_41345,N_41346,N_41347,N_41348,N_41349,N_41350,N_41351,N_41352,N_41353,N_41354,N_41355,N_41356,N_41357,N_41358,N_41359,N_41360,N_41361,N_41362,N_41363,N_41364,N_41365,N_41366,N_41367,N_41368,N_41369,N_41370,N_41371,N_41372,N_41373,N_41374,N_41375,N_41376,N_41377,N_41378,N_41379,N_41380,N_41381,N_41382,N_41383,N_41384,N_41385,N_41386,N_41387,N_41388,N_41389,N_41390,N_41391,N_41392,N_41393,N_41394,N_41395,N_41396,N_41397,N_41398,N_41399,N_41400,N_41401,N_41402,N_41403,N_41404,N_41405,N_41406,N_41407,N_41408,N_41409,N_41410,N_41411,N_41412,N_41413,N_41414,N_41415,N_41416,N_41417,N_41418,N_41419,N_41420,N_41421,N_41422,N_41423,N_41424,N_41425,N_41426,N_41427,N_41428,N_41429,N_41430,N_41431,N_41432,N_41433,N_41434,N_41435,N_41436,N_41437,N_41438,N_41439,N_41440,N_41441,N_41442,N_41443,N_41444,N_41445,N_41446,N_41447,N_41448,N_41449,N_41450,N_41451,N_41452,N_41453,N_41454,N_41455,N_41456,N_41457,N_41458,N_41459,N_41460,N_41461,N_41462,N_41463,N_41464,N_41465,N_41466,N_41467,N_41468,N_41469,N_41470,N_41471,N_41472,N_41473,N_41474,N_41475,N_41476,N_41477,N_41478,N_41479,N_41480,N_41481,N_41482,N_41483,N_41484,N_41485,N_41486,N_41487,N_41488,N_41489,N_41490,N_41491,N_41492,N_41493,N_41494,N_41495,N_41496,N_41497,N_41498,N_41499,N_41500,N_41501,N_41502,N_41503,N_41504,N_41505,N_41506,N_41507,N_41508,N_41509,N_41510,N_41511,N_41512,N_41513,N_41514,N_41515,N_41516,N_41517,N_41518,N_41519,N_41520,N_41521,N_41522,N_41523,N_41524,N_41525,N_41526,N_41527,N_41528,N_41529,N_41530,N_41531,N_41532,N_41533,N_41534,N_41535,N_41536,N_41537,N_41538,N_41539,N_41540,N_41541,N_41542,N_41543,N_41544,N_41545,N_41546,N_41547,N_41548,N_41549,N_41550,N_41551,N_41552,N_41553,N_41554,N_41555,N_41556,N_41557,N_41558,N_41559,N_41560,N_41561,N_41562,N_41563,N_41564,N_41565,N_41566,N_41567,N_41568,N_41569,N_41570,N_41571,N_41572,N_41573,N_41574,N_41575,N_41576,N_41577,N_41578,N_41579,N_41580,N_41581,N_41582,N_41583,N_41584,N_41585,N_41586,N_41587,N_41588,N_41589,N_41590,N_41591,N_41592,N_41593,N_41594,N_41595,N_41596,N_41597,N_41598,N_41599,N_41600,N_41601,N_41602,N_41603,N_41604,N_41605,N_41606,N_41607,N_41608,N_41609,N_41610,N_41611,N_41612,N_41613,N_41614,N_41615,N_41616,N_41617,N_41618,N_41619,N_41620,N_41621,N_41622,N_41623,N_41624,N_41625,N_41626,N_41627,N_41628,N_41629,N_41630,N_41631,N_41632,N_41633,N_41634,N_41635,N_41636,N_41637,N_41638,N_41639,N_41640,N_41641,N_41642,N_41643,N_41644,N_41645,N_41646,N_41647,N_41648,N_41649,N_41650,N_41651,N_41652,N_41653,N_41654,N_41655,N_41656,N_41657,N_41658,N_41659,N_41660,N_41661,N_41662,N_41663,N_41664,N_41665,N_41666,N_41667,N_41668,N_41669,N_41670,N_41671,N_41672,N_41673,N_41674,N_41675,N_41676,N_41677,N_41678,N_41679,N_41680,N_41681,N_41682,N_41683,N_41684,N_41685,N_41686,N_41687,N_41688,N_41689,N_41690,N_41691,N_41692,N_41693,N_41694,N_41695,N_41696,N_41697,N_41698,N_41699,N_41700,N_41701,N_41702,N_41703,N_41704,N_41705,N_41706,N_41707,N_41708,N_41709,N_41710,N_41711,N_41712,N_41713,N_41714,N_41715,N_41716,N_41717,N_41718,N_41719,N_41720,N_41721,N_41722,N_41723,N_41724,N_41725,N_41726,N_41727,N_41728,N_41729,N_41730,N_41731,N_41732,N_41733,N_41734,N_41735,N_41736,N_41737,N_41738,N_41739,N_41740,N_41741,N_41742,N_41743,N_41744,N_41745,N_41746,N_41747,N_41748,N_41749,N_41750,N_41751,N_41752,N_41753,N_41754,N_41755,N_41756,N_41757,N_41758,N_41759,N_41760,N_41761,N_41762,N_41763,N_41764,N_41765,N_41766,N_41767,N_41768,N_41769,N_41770,N_41771,N_41772,N_41773,N_41774,N_41775,N_41776,N_41777,N_41778,N_41779,N_41780,N_41781,N_41782,N_41783,N_41784,N_41785,N_41786,N_41787,N_41788,N_41789,N_41790,N_41791,N_41792,N_41793,N_41794,N_41795,N_41796,N_41797,N_41798,N_41799,N_41800,N_41801,N_41802,N_41803,N_41804,N_41805,N_41806,N_41807,N_41808,N_41809,N_41810,N_41811,N_41812,N_41813,N_41814,N_41815,N_41816,N_41817,N_41818,N_41819,N_41820,N_41821,N_41822,N_41823,N_41824,N_41825,N_41826,N_41827,N_41828,N_41829,N_41830,N_41831,N_41832,N_41833,N_41834,N_41835,N_41836,N_41837,N_41838,N_41839,N_41840,N_41841,N_41842,N_41843,N_41844,N_41845,N_41846,N_41847,N_41848,N_41849,N_41850,N_41851,N_41852,N_41853,N_41854,N_41855,N_41856,N_41857,N_41858,N_41859,N_41860,N_41861,N_41862,N_41863,N_41864,N_41865,N_41866,N_41867,N_41868,N_41869,N_41870,N_41871,N_41872,N_41873,N_41874,N_41875,N_41876,N_41877,N_41878,N_41879,N_41880,N_41881,N_41882,N_41883,N_41884,N_41885,N_41886,N_41887,N_41888,N_41889,N_41890,N_41891,N_41892,N_41893,N_41894,N_41895,N_41896,N_41897,N_41898,N_41899,N_41900,N_41901,N_41902,N_41903,N_41904,N_41905,N_41906,N_41907,N_41908,N_41909,N_41910,N_41911,N_41912,N_41913,N_41914,N_41915,N_41916,N_41917,N_41918,N_41919,N_41920,N_41921,N_41922,N_41923,N_41924,N_41925,N_41926,N_41927,N_41928,N_41929,N_41930,N_41931,N_41932,N_41933,N_41934,N_41935,N_41936,N_41937,N_41938,N_41939,N_41940,N_41941,N_41942,N_41943,N_41944,N_41945,N_41946,N_41947,N_41948,N_41949,N_41950,N_41951,N_41952,N_41953,N_41954,N_41955,N_41956,N_41957,N_41958,N_41959,N_41960,N_41961,N_41962,N_41963,N_41964,N_41965,N_41966,N_41967,N_41968,N_41969,N_41970,N_41971,N_41972,N_41973,N_41974,N_41975,N_41976,N_41977,N_41978,N_41979,N_41980,N_41981,N_41982,N_41983,N_41984,N_41985,N_41986,N_41987,N_41988,N_41989,N_41990,N_41991,N_41992,N_41993,N_41994,N_41995,N_41996,N_41997,N_41998,N_41999,N_42000,N_42001,N_42002,N_42003,N_42004,N_42005,N_42006,N_42007,N_42008,N_42009,N_42010,N_42011,N_42012,N_42013,N_42014,N_42015,N_42016,N_42017,N_42018,N_42019,N_42020,N_42021,N_42022,N_42023,N_42024,N_42025,N_42026,N_42027,N_42028,N_42029,N_42030,N_42031,N_42032,N_42033,N_42034,N_42035,N_42036,N_42037,N_42038,N_42039,N_42040,N_42041,N_42042,N_42043,N_42044,N_42045,N_42046,N_42047,N_42048,N_42049,N_42050,N_42051,N_42052,N_42053,N_42054,N_42055,N_42056,N_42057,N_42058,N_42059,N_42060,N_42061,N_42062,N_42063,N_42064,N_42065,N_42066,N_42067,N_42068,N_42069,N_42070,N_42071,N_42072,N_42073,N_42074,N_42075,N_42076,N_42077,N_42078,N_42079,N_42080,N_42081,N_42082,N_42083,N_42084,N_42085,N_42086,N_42087,N_42088,N_42089,N_42090,N_42091,N_42092,N_42093,N_42094,N_42095,N_42096,N_42097,N_42098,N_42099,N_42100,N_42101,N_42102,N_42103,N_42104,N_42105,N_42106,N_42107,N_42108,N_42109,N_42110,N_42111,N_42112,N_42113,N_42114,N_42115,N_42116,N_42117,N_42118,N_42119,N_42120,N_42121,N_42122,N_42123,N_42124,N_42125,N_42126,N_42127,N_42128,N_42129,N_42130,N_42131,N_42132,N_42133,N_42134,N_42135,N_42136,N_42137,N_42138,N_42139,N_42140,N_42141,N_42142,N_42143,N_42144,N_42145,N_42146,N_42147,N_42148,N_42149,N_42150,N_42151,N_42152,N_42153,N_42154,N_42155,N_42156,N_42157,N_42158,N_42159,N_42160,N_42161,N_42162,N_42163,N_42164,N_42165,N_42166,N_42167,N_42168,N_42169,N_42170,N_42171,N_42172,N_42173,N_42174,N_42175,N_42176,N_42177,N_42178,N_42179,N_42180,N_42181,N_42182,N_42183,N_42184,N_42185,N_42186,N_42187,N_42188,N_42189,N_42190,N_42191,N_42192,N_42193,N_42194,N_42195,N_42196,N_42197,N_42198,N_42199,N_42200,N_42201,N_42202,N_42203,N_42204,N_42205,N_42206,N_42207,N_42208,N_42209,N_42210,N_42211,N_42212,N_42213,N_42214,N_42215,N_42216,N_42217,N_42218,N_42219,N_42220,N_42221,N_42222,N_42223,N_42224,N_42225,N_42226,N_42227,N_42228,N_42229,N_42230,N_42231,N_42232,N_42233,N_42234,N_42235,N_42236,N_42237,N_42238,N_42239,N_42240,N_42241,N_42242,N_42243,N_42244,N_42245,N_42246,N_42247,N_42248,N_42249,N_42250,N_42251,N_42252,N_42253,N_42254,N_42255,N_42256,N_42257,N_42258,N_42259,N_42260,N_42261,N_42262,N_42263,N_42264,N_42265,N_42266,N_42267,N_42268,N_42269,N_42270,N_42271,N_42272,N_42273,N_42274,N_42275,N_42276,N_42277,N_42278,N_42279,N_42280,N_42281,N_42282,N_42283,N_42284,N_42285,N_42286,N_42287,N_42288,N_42289,N_42290,N_42291,N_42292,N_42293,N_42294,N_42295,N_42296,N_42297,N_42298,N_42299,N_42300,N_42301,N_42302,N_42303,N_42304,N_42305,N_42306,N_42307,N_42308,N_42309,N_42310,N_42311,N_42312,N_42313,N_42314,N_42315,N_42316,N_42317,N_42318,N_42319,N_42320,N_42321,N_42322,N_42323,N_42324,N_42325,N_42326,N_42327,N_42328,N_42329,N_42330,N_42331,N_42332,N_42333,N_42334,N_42335,N_42336,N_42337,N_42338,N_42339,N_42340,N_42341,N_42342,N_42343,N_42344,N_42345,N_42346,N_42347,N_42348,N_42349,N_42350,N_42351,N_42352,N_42353,N_42354,N_42355,N_42356,N_42357,N_42358,N_42359,N_42360,N_42361,N_42362,N_42363,N_42364,N_42365,N_42366,N_42367,N_42368,N_42369,N_42370,N_42371,N_42372,N_42373,N_42374,N_42375,N_42376,N_42377,N_42378,N_42379,N_42380,N_42381,N_42382,N_42383,N_42384,N_42385,N_42386,N_42387,N_42388,N_42389,N_42390,N_42391,N_42392,N_42393,N_42394,N_42395,N_42396,N_42397,N_42398,N_42399,N_42400,N_42401,N_42402,N_42403,N_42404,N_42405,N_42406,N_42407,N_42408,N_42409,N_42410,N_42411,N_42412,N_42413,N_42414,N_42415,N_42416,N_42417,N_42418,N_42419,N_42420,N_42421,N_42422,N_42423,N_42424,N_42425,N_42426,N_42427,N_42428,N_42429,N_42430,N_42431,N_42432,N_42433,N_42434,N_42435,N_42436,N_42437,N_42438,N_42439,N_42440,N_42441,N_42442,N_42443,N_42444,N_42445,N_42446,N_42447,N_42448,N_42449,N_42450,N_42451,N_42452,N_42453,N_42454,N_42455,N_42456,N_42457,N_42458,N_42459,N_42460,N_42461,N_42462,N_42463,N_42464,N_42465,N_42466,N_42467,N_42468,N_42469,N_42470,N_42471,N_42472,N_42473,N_42474,N_42475,N_42476,N_42477,N_42478,N_42479,N_42480,N_42481,N_42482,N_42483,N_42484,N_42485,N_42486,N_42487,N_42488,N_42489,N_42490,N_42491,N_42492,N_42493,N_42494,N_42495,N_42496,N_42497,N_42498,N_42499,N_42500,N_42501,N_42502,N_42503,N_42504,N_42505,N_42506,N_42507,N_42508,N_42509,N_42510,N_42511,N_42512,N_42513,N_42514,N_42515,N_42516,N_42517,N_42518,N_42519,N_42520,N_42521,N_42522,N_42523,N_42524,N_42525,N_42526,N_42527,N_42528,N_42529,N_42530,N_42531,N_42532,N_42533,N_42534,N_42535,N_42536,N_42537,N_42538,N_42539,N_42540,N_42541,N_42542,N_42543,N_42544,N_42545,N_42546,N_42547,N_42548,N_42549,N_42550,N_42551,N_42552,N_42553,N_42554,N_42555,N_42556,N_42557,N_42558,N_42559,N_42560,N_42561,N_42562,N_42563,N_42564,N_42565,N_42566,N_42567,N_42568,N_42569,N_42570,N_42571,N_42572,N_42573,N_42574,N_42575,N_42576,N_42577,N_42578,N_42579,N_42580,N_42581,N_42582,N_42583,N_42584,N_42585,N_42586,N_42587,N_42588,N_42589,N_42590,N_42591,N_42592,N_42593,N_42594,N_42595,N_42596,N_42597,N_42598,N_42599,N_42600,N_42601,N_42602,N_42603,N_42604,N_42605,N_42606,N_42607,N_42608,N_42609,N_42610,N_42611,N_42612,N_42613,N_42614,N_42615,N_42616,N_42617,N_42618,N_42619,N_42620,N_42621,N_42622,N_42623,N_42624,N_42625,N_42626,N_42627,N_42628,N_42629,N_42630,N_42631,N_42632,N_42633,N_42634,N_42635,N_42636,N_42637,N_42638,N_42639,N_42640,N_42641,N_42642,N_42643,N_42644,N_42645,N_42646,N_42647,N_42648,N_42649,N_42650,N_42651,N_42652,N_42653,N_42654,N_42655,N_42656,N_42657,N_42658,N_42659,N_42660,N_42661,N_42662,N_42663,N_42664,N_42665,N_42666,N_42667,N_42668,N_42669,N_42670,N_42671,N_42672,N_42673,N_42674,N_42675,N_42676,N_42677,N_42678,N_42679,N_42680,N_42681,N_42682,N_42683,N_42684,N_42685,N_42686,N_42687,N_42688,N_42689,N_42690,N_42691,N_42692,N_42693,N_42694,N_42695,N_42696,N_42697,N_42698,N_42699,N_42700,N_42701,N_42702,N_42703,N_42704,N_42705,N_42706,N_42707,N_42708,N_42709,N_42710,N_42711,N_42712,N_42713,N_42714,N_42715,N_42716,N_42717,N_42718,N_42719,N_42720,N_42721,N_42722,N_42723,N_42724,N_42725,N_42726,N_42727,N_42728,N_42729,N_42730,N_42731,N_42732,N_42733,N_42734,N_42735,N_42736,N_42737,N_42738,N_42739,N_42740,N_42741,N_42742,N_42743,N_42744,N_42745,N_42746,N_42747,N_42748,N_42749,N_42750,N_42751,N_42752,N_42753,N_42754,N_42755,N_42756,N_42757,N_42758,N_42759,N_42760,N_42761,N_42762,N_42763,N_42764,N_42765,N_42766,N_42767,N_42768,N_42769,N_42770,N_42771,N_42772,N_42773,N_42774,N_42775,N_42776,N_42777,N_42778,N_42779,N_42780,N_42781,N_42782,N_42783,N_42784,N_42785,N_42786,N_42787,N_42788,N_42789,N_42790,N_42791,N_42792,N_42793,N_42794,N_42795,N_42796,N_42797,N_42798,N_42799,N_42800,N_42801,N_42802,N_42803,N_42804,N_42805,N_42806,N_42807,N_42808,N_42809,N_42810,N_42811,N_42812,N_42813,N_42814,N_42815,N_42816,N_42817,N_42818,N_42819,N_42820,N_42821,N_42822,N_42823,N_42824,N_42825,N_42826,N_42827,N_42828,N_42829,N_42830,N_42831,N_42832,N_42833,N_42834,N_42835,N_42836,N_42837,N_42838,N_42839,N_42840,N_42841,N_42842,N_42843,N_42844,N_42845,N_42846,N_42847,N_42848,N_42849,N_42850,N_42851,N_42852,N_42853,N_42854,N_42855,N_42856,N_42857,N_42858,N_42859,N_42860,N_42861,N_42862,N_42863,N_42864,N_42865,N_42866,N_42867,N_42868,N_42869,N_42870,N_42871,N_42872,N_42873,N_42874,N_42875,N_42876,N_42877,N_42878,N_42879,N_42880,N_42881,N_42882,N_42883,N_42884,N_42885,N_42886,N_42887,N_42888,N_42889,N_42890,N_42891,N_42892,N_42893,N_42894,N_42895,N_42896,N_42897,N_42898,N_42899,N_42900,N_42901,N_42902,N_42903,N_42904,N_42905,N_42906,N_42907,N_42908,N_42909,N_42910,N_42911,N_42912,N_42913,N_42914,N_42915,N_42916,N_42917,N_42918,N_42919,N_42920,N_42921,N_42922,N_42923,N_42924,N_42925,N_42926,N_42927,N_42928,N_42929,N_42930,N_42931,N_42932,N_42933,N_42934,N_42935,N_42936,N_42937,N_42938,N_42939,N_42940,N_42941,N_42942,N_42943,N_42944,N_42945,N_42946,N_42947,N_42948,N_42949,N_42950,N_42951,N_42952,N_42953,N_42954,N_42955,N_42956,N_42957,N_42958,N_42959,N_42960,N_42961,N_42962,N_42963,N_42964,N_42965,N_42966,N_42967,N_42968,N_42969,N_42970,N_42971,N_42972,N_42973,N_42974,N_42975,N_42976,N_42977,N_42978,N_42979,N_42980,N_42981,N_42982,N_42983,N_42984,N_42985,N_42986,N_42987,N_42988,N_42989,N_42990,N_42991,N_42992,N_42993,N_42994,N_42995,N_42996,N_42997,N_42998,N_42999,N_43000,N_43001,N_43002,N_43003,N_43004,N_43005,N_43006,N_43007,N_43008,N_43009,N_43010,N_43011,N_43012,N_43013,N_43014,N_43015,N_43016,N_43017,N_43018,N_43019,N_43020,N_43021,N_43022,N_43023,N_43024,N_43025,N_43026,N_43027,N_43028,N_43029,N_43030,N_43031,N_43032,N_43033,N_43034,N_43035,N_43036,N_43037,N_43038,N_43039,N_43040,N_43041,N_43042,N_43043,N_43044,N_43045,N_43046,N_43047,N_43048,N_43049,N_43050,N_43051,N_43052,N_43053,N_43054,N_43055,N_43056,N_43057,N_43058,N_43059,N_43060,N_43061,N_43062,N_43063,N_43064,N_43065,N_43066,N_43067,N_43068,N_43069,N_43070,N_43071,N_43072,N_43073,N_43074,N_43075,N_43076,N_43077,N_43078,N_43079,N_43080,N_43081,N_43082,N_43083,N_43084,N_43085,N_43086,N_43087,N_43088,N_43089,N_43090,N_43091,N_43092,N_43093,N_43094,N_43095,N_43096,N_43097,N_43098,N_43099,N_43100,N_43101,N_43102,N_43103,N_43104,N_43105,N_43106,N_43107,N_43108,N_43109,N_43110,N_43111,N_43112,N_43113,N_43114,N_43115,N_43116,N_43117,N_43118,N_43119,N_43120,N_43121,N_43122,N_43123,N_43124,N_43125,N_43126,N_43127,N_43128,N_43129,N_43130,N_43131,N_43132,N_43133,N_43134,N_43135,N_43136,N_43137,N_43138,N_43139,N_43140,N_43141,N_43142,N_43143,N_43144,N_43145,N_43146,N_43147,N_43148,N_43149,N_43150,N_43151,N_43152,N_43153,N_43154,N_43155,N_43156,N_43157,N_43158,N_43159,N_43160,N_43161,N_43162,N_43163,N_43164,N_43165,N_43166,N_43167,N_43168,N_43169,N_43170,N_43171,N_43172,N_43173,N_43174,N_43175,N_43176,N_43177,N_43178,N_43179,N_43180,N_43181,N_43182,N_43183,N_43184,N_43185,N_43186,N_43187,N_43188,N_43189,N_43190,N_43191,N_43192,N_43193,N_43194,N_43195,N_43196,N_43197,N_43198,N_43199,N_43200,N_43201,N_43202,N_43203,N_43204,N_43205,N_43206,N_43207,N_43208,N_43209,N_43210,N_43211,N_43212,N_43213,N_43214,N_43215,N_43216,N_43217,N_43218,N_43219,N_43220,N_43221,N_43222,N_43223,N_43224,N_43225,N_43226,N_43227,N_43228,N_43229,N_43230,N_43231,N_43232,N_43233,N_43234,N_43235,N_43236,N_43237,N_43238,N_43239,N_43240,N_43241,N_43242,N_43243,N_43244,N_43245,N_43246,N_43247,N_43248,N_43249,N_43250,N_43251,N_43252,N_43253,N_43254,N_43255,N_43256,N_43257,N_43258,N_43259,N_43260,N_43261,N_43262,N_43263,N_43264,N_43265,N_43266,N_43267,N_43268,N_43269,N_43270,N_43271,N_43272,N_43273,N_43274,N_43275,N_43276,N_43277,N_43278,N_43279,N_43280,N_43281,N_43282,N_43283,N_43284,N_43285,N_43286,N_43287,N_43288,N_43289,N_43290,N_43291,N_43292,N_43293,N_43294,N_43295,N_43296,N_43297,N_43298,N_43299,N_43300,N_43301,N_43302,N_43303,N_43304,N_43305,N_43306,N_43307,N_43308,N_43309,N_43310,N_43311,N_43312,N_43313,N_43314,N_43315,N_43316,N_43317,N_43318,N_43319,N_43320,N_43321,N_43322,N_43323,N_43324,N_43325,N_43326,N_43327,N_43328,N_43329,N_43330,N_43331,N_43332,N_43333,N_43334,N_43335,N_43336,N_43337,N_43338,N_43339,N_43340,N_43341,N_43342,N_43343,N_43344,N_43345,N_43346,N_43347,N_43348,N_43349,N_43350,N_43351,N_43352,N_43353,N_43354,N_43355,N_43356,N_43357,N_43358,N_43359,N_43360,N_43361,N_43362,N_43363,N_43364,N_43365,N_43366,N_43367,N_43368,N_43369,N_43370,N_43371,N_43372,N_43373,N_43374,N_43375,N_43376,N_43377,N_43378,N_43379,N_43380,N_43381,N_43382,N_43383,N_43384,N_43385,N_43386,N_43387,N_43388,N_43389,N_43390,N_43391,N_43392,N_43393,N_43394,N_43395,N_43396,N_43397,N_43398,N_43399,N_43400,N_43401,N_43402,N_43403,N_43404,N_43405,N_43406,N_43407,N_43408,N_43409,N_43410,N_43411,N_43412,N_43413,N_43414,N_43415,N_43416,N_43417,N_43418,N_43419,N_43420,N_43421,N_43422,N_43423,N_43424,N_43425,N_43426,N_43427,N_43428,N_43429,N_43430,N_43431,N_43432,N_43433,N_43434,N_43435,N_43436,N_43437,N_43438,N_43439,N_43440,N_43441,N_43442,N_43443,N_43444,N_43445,N_43446,N_43447,N_43448,N_43449,N_43450,N_43451,N_43452,N_43453,N_43454,N_43455,N_43456,N_43457,N_43458,N_43459,N_43460,N_43461,N_43462,N_43463,N_43464,N_43465,N_43466,N_43467,N_43468,N_43469,N_43470,N_43471,N_43472,N_43473,N_43474,N_43475,N_43476,N_43477,N_43478,N_43479,N_43480,N_43481,N_43482,N_43483,N_43484,N_43485,N_43486,N_43487,N_43488,N_43489,N_43490,N_43491,N_43492,N_43493,N_43494,N_43495,N_43496,N_43497,N_43498,N_43499,N_43500,N_43501,N_43502,N_43503,N_43504,N_43505,N_43506,N_43507,N_43508,N_43509,N_43510,N_43511,N_43512,N_43513,N_43514,N_43515,N_43516,N_43517,N_43518,N_43519,N_43520,N_43521,N_43522,N_43523,N_43524,N_43525,N_43526,N_43527,N_43528,N_43529,N_43530,N_43531,N_43532,N_43533,N_43534,N_43535,N_43536,N_43537,N_43538,N_43539,N_43540,N_43541,N_43542,N_43543,N_43544,N_43545,N_43546,N_43547,N_43548,N_43549,N_43550,N_43551,N_43552,N_43553,N_43554,N_43555,N_43556,N_43557,N_43558,N_43559,N_43560,N_43561,N_43562,N_43563,N_43564,N_43565,N_43566,N_43567,N_43568,N_43569,N_43570,N_43571,N_43572,N_43573,N_43574,N_43575,N_43576,N_43577,N_43578,N_43579,N_43580,N_43581,N_43582,N_43583,N_43584,N_43585,N_43586,N_43587,N_43588,N_43589,N_43590,N_43591,N_43592,N_43593,N_43594,N_43595,N_43596,N_43597,N_43598,N_43599,N_43600,N_43601,N_43602,N_43603,N_43604,N_43605,N_43606,N_43607,N_43608,N_43609,N_43610,N_43611,N_43612,N_43613,N_43614,N_43615,N_43616,N_43617,N_43618,N_43619,N_43620,N_43621,N_43622,N_43623,N_43624,N_43625,N_43626,N_43627,N_43628,N_43629,N_43630,N_43631,N_43632,N_43633,N_43634,N_43635,N_43636,N_43637,N_43638,N_43639,N_43640,N_43641,N_43642,N_43643,N_43644,N_43645,N_43646,N_43647,N_43648,N_43649,N_43650,N_43651,N_43652,N_43653,N_43654,N_43655,N_43656,N_43657,N_43658,N_43659,N_43660,N_43661,N_43662,N_43663,N_43664,N_43665,N_43666,N_43667,N_43668,N_43669,N_43670,N_43671,N_43672,N_43673,N_43674,N_43675,N_43676,N_43677,N_43678,N_43679,N_43680,N_43681,N_43682,N_43683,N_43684,N_43685,N_43686,N_43687,N_43688,N_43689,N_43690,N_43691,N_43692,N_43693,N_43694,N_43695,N_43696,N_43697,N_43698,N_43699,N_43700,N_43701,N_43702,N_43703,N_43704,N_43705,N_43706,N_43707,N_43708,N_43709,N_43710,N_43711,N_43712,N_43713,N_43714,N_43715,N_43716,N_43717,N_43718,N_43719,N_43720,N_43721,N_43722,N_43723,N_43724,N_43725,N_43726,N_43727,N_43728,N_43729,N_43730,N_43731,N_43732,N_43733,N_43734,N_43735,N_43736,N_43737,N_43738,N_43739,N_43740,N_43741,N_43742,N_43743,N_43744,N_43745,N_43746,N_43747,N_43748,N_43749,N_43750,N_43751,N_43752,N_43753,N_43754,N_43755,N_43756,N_43757,N_43758,N_43759,N_43760,N_43761,N_43762,N_43763,N_43764,N_43765,N_43766,N_43767,N_43768,N_43769,N_43770,N_43771,N_43772,N_43773,N_43774,N_43775,N_43776,N_43777,N_43778,N_43779,N_43780,N_43781,N_43782,N_43783,N_43784,N_43785,N_43786,N_43787,N_43788,N_43789,N_43790,N_43791,N_43792,N_43793,N_43794,N_43795,N_43796,N_43797,N_43798,N_43799,N_43800,N_43801,N_43802,N_43803,N_43804,N_43805,N_43806,N_43807,N_43808,N_43809,N_43810,N_43811,N_43812,N_43813,N_43814,N_43815,N_43816,N_43817,N_43818,N_43819,N_43820,N_43821,N_43822,N_43823,N_43824,N_43825,N_43826,N_43827,N_43828,N_43829,N_43830,N_43831,N_43832,N_43833,N_43834,N_43835,N_43836,N_43837,N_43838,N_43839,N_43840,N_43841,N_43842,N_43843,N_43844,N_43845,N_43846,N_43847,N_43848,N_43849,N_43850,N_43851,N_43852,N_43853,N_43854,N_43855,N_43856,N_43857,N_43858,N_43859,N_43860,N_43861,N_43862,N_43863,N_43864,N_43865,N_43866,N_43867,N_43868,N_43869,N_43870,N_43871,N_43872,N_43873,N_43874,N_43875,N_43876,N_43877,N_43878,N_43879,N_43880,N_43881,N_43882,N_43883,N_43884,N_43885,N_43886,N_43887,N_43888,N_43889,N_43890,N_43891,N_43892,N_43893,N_43894,N_43895,N_43896,N_43897,N_43898,N_43899,N_43900,N_43901,N_43902,N_43903,N_43904,N_43905,N_43906,N_43907,N_43908,N_43909,N_43910,N_43911,N_43912,N_43913,N_43914,N_43915,N_43916,N_43917,N_43918,N_43919,N_43920,N_43921,N_43922,N_43923,N_43924,N_43925,N_43926,N_43927,N_43928,N_43929,N_43930,N_43931,N_43932,N_43933,N_43934,N_43935,N_43936,N_43937,N_43938,N_43939,N_43940,N_43941,N_43942,N_43943,N_43944,N_43945,N_43946,N_43947,N_43948,N_43949,N_43950,N_43951,N_43952,N_43953,N_43954,N_43955,N_43956,N_43957,N_43958,N_43959,N_43960,N_43961,N_43962,N_43963,N_43964,N_43965,N_43966,N_43967,N_43968,N_43969,N_43970,N_43971,N_43972,N_43973,N_43974,N_43975,N_43976,N_43977,N_43978,N_43979,N_43980,N_43981,N_43982,N_43983,N_43984,N_43985,N_43986,N_43987,N_43988,N_43989,N_43990,N_43991,N_43992,N_43993,N_43994,N_43995,N_43996,N_43997,N_43998,N_43999,N_44000,N_44001,N_44002,N_44003,N_44004,N_44005,N_44006,N_44007,N_44008,N_44009,N_44010,N_44011,N_44012,N_44013,N_44014,N_44015,N_44016,N_44017,N_44018,N_44019,N_44020,N_44021,N_44022,N_44023,N_44024,N_44025,N_44026,N_44027,N_44028,N_44029,N_44030,N_44031,N_44032,N_44033,N_44034,N_44035,N_44036,N_44037,N_44038,N_44039,N_44040,N_44041,N_44042,N_44043,N_44044,N_44045,N_44046,N_44047,N_44048,N_44049,N_44050,N_44051,N_44052,N_44053,N_44054,N_44055,N_44056,N_44057,N_44058,N_44059,N_44060,N_44061,N_44062,N_44063,N_44064,N_44065,N_44066,N_44067,N_44068,N_44069,N_44070,N_44071,N_44072,N_44073,N_44074,N_44075,N_44076,N_44077,N_44078,N_44079,N_44080,N_44081,N_44082,N_44083,N_44084,N_44085,N_44086,N_44087,N_44088,N_44089,N_44090,N_44091,N_44092,N_44093,N_44094,N_44095,N_44096,N_44097,N_44098,N_44099,N_44100,N_44101,N_44102,N_44103,N_44104,N_44105,N_44106,N_44107,N_44108,N_44109,N_44110,N_44111,N_44112,N_44113,N_44114,N_44115,N_44116,N_44117,N_44118,N_44119,N_44120,N_44121,N_44122,N_44123,N_44124,N_44125,N_44126,N_44127,N_44128,N_44129,N_44130,N_44131,N_44132,N_44133,N_44134,N_44135,N_44136,N_44137,N_44138,N_44139,N_44140,N_44141,N_44142,N_44143,N_44144,N_44145,N_44146,N_44147,N_44148,N_44149,N_44150,N_44151,N_44152,N_44153,N_44154,N_44155,N_44156,N_44157,N_44158,N_44159,N_44160,N_44161,N_44162,N_44163,N_44164,N_44165,N_44166,N_44167,N_44168,N_44169,N_44170,N_44171,N_44172,N_44173,N_44174,N_44175,N_44176,N_44177,N_44178,N_44179,N_44180,N_44181,N_44182,N_44183,N_44184,N_44185,N_44186,N_44187,N_44188,N_44189,N_44190,N_44191,N_44192,N_44193,N_44194,N_44195,N_44196,N_44197,N_44198,N_44199,N_44200,N_44201,N_44202,N_44203,N_44204,N_44205,N_44206,N_44207,N_44208,N_44209,N_44210,N_44211,N_44212,N_44213,N_44214,N_44215,N_44216,N_44217,N_44218,N_44219,N_44220,N_44221,N_44222,N_44223,N_44224,N_44225,N_44226,N_44227,N_44228,N_44229,N_44230,N_44231,N_44232,N_44233,N_44234,N_44235,N_44236,N_44237,N_44238,N_44239,N_44240,N_44241,N_44242,N_44243,N_44244,N_44245,N_44246,N_44247,N_44248,N_44249,N_44250,N_44251,N_44252,N_44253,N_44254,N_44255,N_44256,N_44257,N_44258,N_44259,N_44260,N_44261,N_44262,N_44263,N_44264,N_44265,N_44266,N_44267,N_44268,N_44269,N_44270,N_44271,N_44272,N_44273,N_44274,N_44275,N_44276,N_44277,N_44278,N_44279,N_44280,N_44281,N_44282,N_44283,N_44284,N_44285,N_44286,N_44287,N_44288,N_44289,N_44290,N_44291,N_44292,N_44293,N_44294,N_44295,N_44296,N_44297,N_44298,N_44299,N_44300,N_44301,N_44302,N_44303,N_44304,N_44305,N_44306,N_44307,N_44308,N_44309,N_44310,N_44311,N_44312,N_44313,N_44314,N_44315,N_44316,N_44317,N_44318,N_44319,N_44320,N_44321,N_44322,N_44323,N_44324,N_44325,N_44326,N_44327,N_44328,N_44329,N_44330,N_44331,N_44332,N_44333,N_44334,N_44335,N_44336,N_44337,N_44338,N_44339,N_44340,N_44341,N_44342,N_44343,N_44344,N_44345,N_44346,N_44347,N_44348,N_44349,N_44350,N_44351,N_44352,N_44353,N_44354,N_44355,N_44356,N_44357,N_44358,N_44359,N_44360,N_44361,N_44362,N_44363,N_44364,N_44365,N_44366,N_44367,N_44368,N_44369,N_44370,N_44371,N_44372,N_44373,N_44374,N_44375,N_44376,N_44377,N_44378,N_44379,N_44380,N_44381,N_44382,N_44383,N_44384,N_44385,N_44386,N_44387,N_44388,N_44389,N_44390,N_44391,N_44392,N_44393,N_44394,N_44395,N_44396,N_44397,N_44398,N_44399,N_44400,N_44401,N_44402,N_44403,N_44404,N_44405,N_44406,N_44407,N_44408,N_44409,N_44410,N_44411,N_44412,N_44413,N_44414,N_44415,N_44416,N_44417,N_44418,N_44419,N_44420,N_44421,N_44422,N_44423,N_44424,N_44425,N_44426,N_44427,N_44428,N_44429,N_44430,N_44431,N_44432,N_44433,N_44434,N_44435,N_44436,N_44437,N_44438,N_44439,N_44440,N_44441,N_44442,N_44443,N_44444,N_44445,N_44446,N_44447,N_44448,N_44449,N_44450,N_44451,N_44452,N_44453,N_44454,N_44455,N_44456,N_44457,N_44458,N_44459,N_44460,N_44461,N_44462,N_44463,N_44464,N_44465,N_44466,N_44467,N_44468,N_44469,N_44470,N_44471,N_44472,N_44473,N_44474,N_44475,N_44476,N_44477,N_44478,N_44479,N_44480,N_44481,N_44482,N_44483,N_44484,N_44485,N_44486,N_44487,N_44488,N_44489,N_44490,N_44491,N_44492,N_44493,N_44494,N_44495,N_44496,N_44497,N_44498,N_44499,N_44500,N_44501,N_44502,N_44503,N_44504,N_44505,N_44506,N_44507,N_44508,N_44509,N_44510,N_44511,N_44512,N_44513,N_44514,N_44515,N_44516,N_44517,N_44518,N_44519,N_44520,N_44521,N_44522,N_44523,N_44524,N_44525,N_44526,N_44527,N_44528,N_44529,N_44530,N_44531,N_44532,N_44533,N_44534,N_44535,N_44536,N_44537,N_44538,N_44539,N_44540,N_44541,N_44542,N_44543,N_44544,N_44545,N_44546,N_44547,N_44548,N_44549,N_44550,N_44551,N_44552,N_44553,N_44554,N_44555,N_44556,N_44557,N_44558,N_44559,N_44560,N_44561,N_44562,N_44563,N_44564,N_44565,N_44566,N_44567,N_44568,N_44569,N_44570,N_44571,N_44572,N_44573,N_44574,N_44575,N_44576,N_44577,N_44578,N_44579,N_44580,N_44581,N_44582,N_44583,N_44584,N_44585,N_44586,N_44587,N_44588,N_44589,N_44590,N_44591,N_44592,N_44593,N_44594,N_44595,N_44596,N_44597,N_44598,N_44599,N_44600,N_44601,N_44602,N_44603,N_44604,N_44605,N_44606,N_44607,N_44608,N_44609,N_44610,N_44611,N_44612,N_44613,N_44614,N_44615,N_44616,N_44617,N_44618,N_44619,N_44620,N_44621,N_44622,N_44623,N_44624,N_44625,N_44626,N_44627,N_44628,N_44629,N_44630,N_44631,N_44632,N_44633,N_44634,N_44635,N_44636,N_44637,N_44638,N_44639,N_44640,N_44641,N_44642,N_44643,N_44644,N_44645,N_44646,N_44647,N_44648,N_44649,N_44650,N_44651,N_44652,N_44653,N_44654,N_44655,N_44656,N_44657,N_44658,N_44659,N_44660,N_44661,N_44662,N_44663,N_44664,N_44665,N_44666,N_44667,N_44668,N_44669,N_44670,N_44671,N_44672,N_44673,N_44674,N_44675,N_44676,N_44677,N_44678,N_44679,N_44680,N_44681,N_44682,N_44683,N_44684,N_44685,N_44686,N_44687,N_44688,N_44689,N_44690,N_44691,N_44692,N_44693,N_44694,N_44695,N_44696,N_44697,N_44698,N_44699,N_44700,N_44701,N_44702,N_44703,N_44704,N_44705,N_44706,N_44707,N_44708,N_44709,N_44710,N_44711,N_44712,N_44713,N_44714,N_44715,N_44716,N_44717,N_44718,N_44719,N_44720,N_44721,N_44722,N_44723,N_44724,N_44725,N_44726,N_44727,N_44728,N_44729,N_44730,N_44731,N_44732,N_44733,N_44734,N_44735,N_44736,N_44737,N_44738,N_44739,N_44740,N_44741,N_44742,N_44743,N_44744,N_44745,N_44746,N_44747,N_44748,N_44749,N_44750,N_44751,N_44752,N_44753,N_44754,N_44755,N_44756,N_44757,N_44758,N_44759,N_44760,N_44761,N_44762,N_44763,N_44764,N_44765,N_44766,N_44767,N_44768,N_44769,N_44770,N_44771,N_44772,N_44773,N_44774,N_44775,N_44776,N_44777,N_44778,N_44779,N_44780,N_44781,N_44782,N_44783,N_44784,N_44785,N_44786,N_44787,N_44788,N_44789,N_44790,N_44791,N_44792,N_44793,N_44794,N_44795,N_44796,N_44797,N_44798,N_44799,N_44800,N_44801,N_44802,N_44803,N_44804,N_44805,N_44806,N_44807,N_44808,N_44809,N_44810,N_44811,N_44812,N_44813,N_44814,N_44815,N_44816,N_44817,N_44818,N_44819,N_44820,N_44821,N_44822,N_44823,N_44824,N_44825,N_44826,N_44827,N_44828,N_44829,N_44830,N_44831,N_44832,N_44833,N_44834,N_44835,N_44836,N_44837,N_44838,N_44839,N_44840,N_44841,N_44842,N_44843,N_44844,N_44845,N_44846,N_44847,N_44848,N_44849,N_44850,N_44851,N_44852,N_44853,N_44854,N_44855,N_44856,N_44857,N_44858,N_44859,N_44860,N_44861,N_44862,N_44863,N_44864,N_44865,N_44866,N_44867,N_44868,N_44869,N_44870,N_44871,N_44872,N_44873,N_44874,N_44875,N_44876,N_44877,N_44878,N_44879,N_44880,N_44881,N_44882,N_44883,N_44884,N_44885,N_44886,N_44887,N_44888,N_44889,N_44890,N_44891,N_44892,N_44893,N_44894,N_44895,N_44896,N_44897,N_44898,N_44899,N_44900,N_44901,N_44902,N_44903,N_44904,N_44905,N_44906,N_44907,N_44908,N_44909,N_44910,N_44911,N_44912,N_44913,N_44914,N_44915,N_44916,N_44917,N_44918,N_44919,N_44920,N_44921,N_44922,N_44923,N_44924,N_44925,N_44926,N_44927,N_44928,N_44929,N_44930,N_44931,N_44932,N_44933,N_44934,N_44935,N_44936,N_44937,N_44938,N_44939,N_44940,N_44941,N_44942,N_44943,N_44944,N_44945,N_44946,N_44947,N_44948,N_44949,N_44950,N_44951,N_44952,N_44953,N_44954,N_44955,N_44956,N_44957,N_44958,N_44959,N_44960,N_44961,N_44962,N_44963,N_44964,N_44965,N_44966,N_44967,N_44968,N_44969,N_44970,N_44971,N_44972,N_44973,N_44974,N_44975,N_44976,N_44977,N_44978,N_44979,N_44980,N_44981,N_44982,N_44983,N_44984,N_44985,N_44986,N_44987,N_44988,N_44989,N_44990,N_44991,N_44992,N_44993,N_44994,N_44995,N_44996,N_44997,N_44998,N_44999,N_45000,N_45001,N_45002,N_45003,N_45004,N_45005,N_45006,N_45007,N_45008,N_45009,N_45010,N_45011,N_45012,N_45013,N_45014,N_45015,N_45016,N_45017,N_45018,N_45019,N_45020,N_45021,N_45022,N_45023,N_45024,N_45025,N_45026,N_45027,N_45028,N_45029,N_45030,N_45031,N_45032,N_45033,N_45034,N_45035,N_45036,N_45037,N_45038,N_45039,N_45040,N_45041,N_45042,N_45043,N_45044,N_45045,N_45046,N_45047,N_45048,N_45049,N_45050,N_45051,N_45052,N_45053,N_45054,N_45055,N_45056,N_45057,N_45058,N_45059,N_45060,N_45061,N_45062,N_45063,N_45064,N_45065,N_45066,N_45067,N_45068,N_45069,N_45070,N_45071,N_45072,N_45073,N_45074,N_45075,N_45076,N_45077,N_45078,N_45079,N_45080,N_45081,N_45082,N_45083,N_45084,N_45085,N_45086,N_45087,N_45088,N_45089,N_45090,N_45091,N_45092,N_45093,N_45094,N_45095,N_45096,N_45097,N_45098,N_45099,N_45100,N_45101,N_45102,N_45103,N_45104,N_45105,N_45106,N_45107,N_45108,N_45109,N_45110,N_45111,N_45112,N_45113,N_45114,N_45115,N_45116,N_45117,N_45118,N_45119,N_45120,N_45121,N_45122,N_45123,N_45124,N_45125,N_45126,N_45127,N_45128,N_45129,N_45130,N_45131,N_45132,N_45133,N_45134,N_45135,N_45136,N_45137,N_45138,N_45139,N_45140,N_45141,N_45142,N_45143,N_45144,N_45145,N_45146,N_45147,N_45148,N_45149,N_45150,N_45151,N_45152,N_45153,N_45154,N_45155,N_45156,N_45157,N_45158,N_45159,N_45160,N_45161,N_45162,N_45163,N_45164,N_45165,N_45166,N_45167,N_45168,N_45169,N_45170,N_45171,N_45172,N_45173,N_45174,N_45175,N_45176,N_45177,N_45178,N_45179,N_45180,N_45181,N_45182,N_45183,N_45184,N_45185,N_45186,N_45187,N_45188,N_45189,N_45190,N_45191,N_45192,N_45193,N_45194,N_45195,N_45196,N_45197,N_45198,N_45199,N_45200,N_45201,N_45202,N_45203,N_45204,N_45205,N_45206,N_45207,N_45208,N_45209,N_45210,N_45211,N_45212,N_45213,N_45214,N_45215,N_45216,N_45217,N_45218,N_45219,N_45220,N_45221,N_45222,N_45223,N_45224,N_45225,N_45226,N_45227,N_45228,N_45229,N_45230,N_45231,N_45232,N_45233,N_45234,N_45235,N_45236,N_45237,N_45238,N_45239,N_45240,N_45241,N_45242,N_45243,N_45244,N_45245,N_45246,N_45247,N_45248,N_45249,N_45250,N_45251,N_45252,N_45253,N_45254,N_45255,N_45256,N_45257,N_45258,N_45259,N_45260,N_45261,N_45262,N_45263,N_45264,N_45265,N_45266,N_45267,N_45268,N_45269,N_45270,N_45271,N_45272,N_45273,N_45274,N_45275,N_45276,N_45277,N_45278,N_45279,N_45280,N_45281,N_45282,N_45283,N_45284,N_45285,N_45286,N_45287,N_45288,N_45289,N_45290,N_45291,N_45292,N_45293,N_45294,N_45295,N_45296,N_45297,N_45298,N_45299,N_45300,N_45301,N_45302,N_45303,N_45304,N_45305,N_45306,N_45307,N_45308,N_45309,N_45310,N_45311,N_45312,N_45313,N_45314,N_45315,N_45316,N_45317,N_45318,N_45319,N_45320,N_45321,N_45322,N_45323,N_45324,N_45325,N_45326,N_45327,N_45328,N_45329,N_45330,N_45331,N_45332,N_45333,N_45334,N_45335,N_45336,N_45337,N_45338,N_45339,N_45340,N_45341,N_45342,N_45343,N_45344,N_45345,N_45346,N_45347,N_45348,N_45349,N_45350,N_45351,N_45352,N_45353,N_45354,N_45355,N_45356,N_45357,N_45358,N_45359,N_45360,N_45361,N_45362,N_45363,N_45364,N_45365,N_45366,N_45367,N_45368,N_45369,N_45370,N_45371,N_45372,N_45373,N_45374,N_45375,N_45376,N_45377,N_45378,N_45379,N_45380,N_45381,N_45382,N_45383,N_45384,N_45385,N_45386,N_45387,N_45388,N_45389,N_45390,N_45391,N_45392,N_45393,N_45394,N_45395,N_45396,N_45397,N_45398,N_45399,N_45400,N_45401,N_45402,N_45403,N_45404,N_45405,N_45406,N_45407,N_45408,N_45409,N_45410,N_45411,N_45412,N_45413,N_45414,N_45415,N_45416,N_45417,N_45418,N_45419,N_45420,N_45421,N_45422,N_45423,N_45424,N_45425,N_45426,N_45427,N_45428,N_45429,N_45430,N_45431,N_45432,N_45433,N_45434,N_45435,N_45436,N_45437,N_45438,N_45439,N_45440,N_45441,N_45442,N_45443,N_45444,N_45445,N_45446,N_45447,N_45448,N_45449,N_45450,N_45451,N_45452,N_45453,N_45454,N_45455,N_45456,N_45457,N_45458,N_45459,N_45460,N_45461,N_45462,N_45463,N_45464,N_45465,N_45466,N_45467,N_45468,N_45469,N_45470,N_45471,N_45472,N_45473,N_45474,N_45475,N_45476,N_45477,N_45478,N_45479,N_45480,N_45481,N_45482,N_45483,N_45484,N_45485,N_45486,N_45487,N_45488,N_45489,N_45490,N_45491,N_45492,N_45493,N_45494,N_45495,N_45496,N_45497,N_45498,N_45499,N_45500,N_45501,N_45502,N_45503,N_45504,N_45505,N_45506,N_45507,N_45508,N_45509,N_45510,N_45511,N_45512,N_45513,N_45514,N_45515,N_45516,N_45517,N_45518,N_45519,N_45520,N_45521,N_45522,N_45523,N_45524,N_45525,N_45526,N_45527,N_45528,N_45529,N_45530,N_45531,N_45532,N_45533,N_45534,N_45535,N_45536,N_45537,N_45538,N_45539,N_45540,N_45541,N_45542,N_45543,N_45544,N_45545,N_45546,N_45547,N_45548,N_45549,N_45550,N_45551,N_45552,N_45553,N_45554,N_45555,N_45556,N_45557,N_45558,N_45559,N_45560,N_45561,N_45562,N_45563,N_45564,N_45565,N_45566,N_45567,N_45568,N_45569,N_45570,N_45571,N_45572,N_45573,N_45574,N_45575,N_45576,N_45577,N_45578,N_45579,N_45580,N_45581,N_45582,N_45583,N_45584,N_45585,N_45586,N_45587,N_45588,N_45589,N_45590,N_45591,N_45592,N_45593,N_45594,N_45595,N_45596,N_45597,N_45598,N_45599,N_45600,N_45601,N_45602,N_45603,N_45604,N_45605,N_45606,N_45607,N_45608,N_45609,N_45610,N_45611,N_45612,N_45613,N_45614,N_45615,N_45616,N_45617,N_45618,N_45619,N_45620,N_45621,N_45622,N_45623,N_45624,N_45625,N_45626,N_45627,N_45628,N_45629,N_45630,N_45631,N_45632,N_45633,N_45634,N_45635,N_45636,N_45637,N_45638,N_45639,N_45640,N_45641,N_45642,N_45643,N_45644,N_45645,N_45646,N_45647,N_45648,N_45649,N_45650,N_45651,N_45652,N_45653,N_45654,N_45655,N_45656,N_45657,N_45658,N_45659,N_45660,N_45661,N_45662,N_45663,N_45664,N_45665,N_45666,N_45667,N_45668,N_45669,N_45670,N_45671,N_45672,N_45673,N_45674,N_45675,N_45676,N_45677,N_45678,N_45679,N_45680,N_45681,N_45682,N_45683,N_45684,N_45685,N_45686,N_45687,N_45688,N_45689,N_45690,N_45691,N_45692,N_45693,N_45694,N_45695,N_45696,N_45697,N_45698,N_45699,N_45700,N_45701,N_45702,N_45703,N_45704,N_45705,N_45706,N_45707,N_45708,N_45709,N_45710,N_45711,N_45712,N_45713,N_45714,N_45715,N_45716,N_45717,N_45718,N_45719,N_45720,N_45721,N_45722,N_45723,N_45724,N_45725,N_45726,N_45727,N_45728,N_45729,N_45730,N_45731,N_45732,N_45733,N_45734,N_45735,N_45736,N_45737,N_45738,N_45739,N_45740,N_45741,N_45742,N_45743,N_45744,N_45745,N_45746,N_45747,N_45748,N_45749,N_45750,N_45751,N_45752,N_45753,N_45754,N_45755,N_45756,N_45757,N_45758,N_45759,N_45760,N_45761,N_45762,N_45763,N_45764,N_45765,N_45766,N_45767,N_45768,N_45769,N_45770,N_45771,N_45772,N_45773,N_45774,N_45775,N_45776,N_45777,N_45778,N_45779,N_45780,N_45781,N_45782,N_45783,N_45784,N_45785,N_45786,N_45787,N_45788,N_45789,N_45790,N_45791,N_45792,N_45793,N_45794,N_45795,N_45796,N_45797,N_45798,N_45799,N_45800,N_45801,N_45802,N_45803,N_45804,N_45805,N_45806,N_45807,N_45808,N_45809,N_45810,N_45811,N_45812,N_45813,N_45814,N_45815,N_45816,N_45817,N_45818,N_45819,N_45820,N_45821,N_45822,N_45823,N_45824,N_45825,N_45826,N_45827,N_45828,N_45829,N_45830,N_45831,N_45832,N_45833,N_45834,N_45835,N_45836,N_45837,N_45838,N_45839,N_45840,N_45841,N_45842,N_45843,N_45844,N_45845,N_45846,N_45847,N_45848,N_45849,N_45850,N_45851,N_45852,N_45853,N_45854,N_45855,N_45856,N_45857,N_45858,N_45859,N_45860,N_45861,N_45862,N_45863,N_45864,N_45865,N_45866,N_45867,N_45868,N_45869,N_45870,N_45871,N_45872,N_45873,N_45874,N_45875,N_45876,N_45877,N_45878,N_45879,N_45880,N_45881,N_45882,N_45883,N_45884,N_45885,N_45886,N_45887,N_45888,N_45889,N_45890,N_45891,N_45892,N_45893,N_45894,N_45895,N_45896,N_45897,N_45898,N_45899,N_45900,N_45901,N_45902,N_45903,N_45904,N_45905,N_45906,N_45907,N_45908,N_45909,N_45910,N_45911,N_45912,N_45913,N_45914,N_45915,N_45916,N_45917,N_45918,N_45919,N_45920,N_45921,N_45922,N_45923,N_45924,N_45925,N_45926,N_45927,N_45928,N_45929,N_45930,N_45931,N_45932,N_45933,N_45934,N_45935,N_45936,N_45937,N_45938,N_45939,N_45940,N_45941,N_45942,N_45943,N_45944,N_45945,N_45946,N_45947,N_45948,N_45949,N_45950,N_45951,N_45952,N_45953,N_45954,N_45955,N_45956,N_45957,N_45958,N_45959,N_45960,N_45961,N_45962,N_45963,N_45964,N_45965,N_45966,N_45967,N_45968,N_45969,N_45970,N_45971,N_45972,N_45973,N_45974,N_45975,N_45976,N_45977,N_45978,N_45979,N_45980,N_45981,N_45982,N_45983,N_45984,N_45985,N_45986,N_45987,N_45988,N_45989,N_45990,N_45991,N_45992,N_45993,N_45994,N_45995,N_45996,N_45997,N_45998,N_45999,N_46000,N_46001,N_46002,N_46003,N_46004,N_46005,N_46006,N_46007,N_46008,N_46009,N_46010,N_46011,N_46012,N_46013,N_46014,N_46015,N_46016,N_46017,N_46018,N_46019,N_46020,N_46021,N_46022,N_46023,N_46024,N_46025,N_46026,N_46027,N_46028,N_46029,N_46030,N_46031,N_46032,N_46033,N_46034,N_46035,N_46036,N_46037,N_46038,N_46039,N_46040,N_46041,N_46042,N_46043,N_46044,N_46045,N_46046,N_46047,N_46048,N_46049,N_46050,N_46051,N_46052,N_46053,N_46054,N_46055,N_46056,N_46057,N_46058,N_46059,N_46060,N_46061,N_46062,N_46063,N_46064,N_46065,N_46066,N_46067,N_46068,N_46069,N_46070,N_46071,N_46072,N_46073,N_46074,N_46075,N_46076,N_46077,N_46078,N_46079,N_46080,N_46081,N_46082,N_46083,N_46084,N_46085,N_46086,N_46087,N_46088,N_46089,N_46090,N_46091,N_46092,N_46093,N_46094,N_46095,N_46096,N_46097,N_46098,N_46099,N_46100,N_46101,N_46102,N_46103,N_46104,N_46105,N_46106,N_46107,N_46108,N_46109,N_46110,N_46111,N_46112,N_46113,N_46114,N_46115,N_46116,N_46117,N_46118,N_46119,N_46120,N_46121,N_46122,N_46123,N_46124,N_46125,N_46126,N_46127,N_46128,N_46129,N_46130,N_46131,N_46132,N_46133,N_46134,N_46135,N_46136,N_46137,N_46138,N_46139,N_46140,N_46141,N_46142,N_46143,N_46144,N_46145,N_46146,N_46147,N_46148,N_46149,N_46150,N_46151,N_46152,N_46153,N_46154,N_46155,N_46156,N_46157,N_46158,N_46159,N_46160,N_46161,N_46162,N_46163,N_46164,N_46165,N_46166,N_46167,N_46168,N_46169,N_46170,N_46171,N_46172,N_46173,N_46174,N_46175,N_46176,N_46177,N_46178,N_46179,N_46180,N_46181,N_46182,N_46183,N_46184,N_46185,N_46186,N_46187,N_46188,N_46189,N_46190,N_46191,N_46192,N_46193,N_46194,N_46195,N_46196,N_46197,N_46198,N_46199,N_46200,N_46201,N_46202,N_46203,N_46204,N_46205,N_46206,N_46207,N_46208,N_46209,N_46210,N_46211,N_46212,N_46213,N_46214,N_46215,N_46216,N_46217,N_46218,N_46219,N_46220,N_46221,N_46222,N_46223,N_46224,N_46225,N_46226,N_46227,N_46228,N_46229,N_46230,N_46231,N_46232,N_46233,N_46234,N_46235,N_46236,N_46237,N_46238,N_46239,N_46240,N_46241,N_46242,N_46243,N_46244,N_46245,N_46246,N_46247,N_46248,N_46249,N_46250,N_46251,N_46252,N_46253,N_46254,N_46255,N_46256,N_46257,N_46258,N_46259,N_46260,N_46261,N_46262,N_46263,N_46264,N_46265,N_46266,N_46267,N_46268,N_46269,N_46270,N_46271,N_46272,N_46273,N_46274,N_46275,N_46276,N_46277,N_46278,N_46279,N_46280,N_46281,N_46282,N_46283,N_46284,N_46285,N_46286,N_46287,N_46288,N_46289,N_46290,N_46291,N_46292,N_46293,N_46294,N_46295,N_46296,N_46297,N_46298,N_46299,N_46300,N_46301,N_46302,N_46303,N_46304,N_46305,N_46306,N_46307,N_46308,N_46309,N_46310,N_46311,N_46312,N_46313,N_46314,N_46315,N_46316,N_46317,N_46318,N_46319,N_46320,N_46321,N_46322,N_46323,N_46324,N_46325,N_46326,N_46327,N_46328,N_46329,N_46330,N_46331,N_46332,N_46333,N_46334,N_46335,N_46336,N_46337,N_46338,N_46339,N_46340,N_46341,N_46342,N_46343,N_46344,N_46345,N_46346,N_46347,N_46348,N_46349,N_46350,N_46351,N_46352,N_46353,N_46354,N_46355,N_46356,N_46357,N_46358,N_46359,N_46360,N_46361,N_46362,N_46363,N_46364,N_46365,N_46366,N_46367,N_46368,N_46369,N_46370,N_46371,N_46372,N_46373,N_46374,N_46375,N_46376,N_46377,N_46378,N_46379,N_46380,N_46381,N_46382,N_46383,N_46384,N_46385,N_46386,N_46387,N_46388,N_46389,N_46390,N_46391,N_46392,N_46393,N_46394,N_46395,N_46396,N_46397,N_46398,N_46399,N_46400,N_46401,N_46402,N_46403,N_46404,N_46405,N_46406,N_46407,N_46408,N_46409,N_46410,N_46411,N_46412,N_46413,N_46414,N_46415,N_46416,N_46417,N_46418,N_46419,N_46420,N_46421,N_46422,N_46423,N_46424,N_46425,N_46426,N_46427,N_46428,N_46429,N_46430,N_46431,N_46432,N_46433,N_46434,N_46435,N_46436,N_46437,N_46438,N_46439,N_46440,N_46441,N_46442,N_46443,N_46444,N_46445,N_46446,N_46447,N_46448,N_46449,N_46450,N_46451,N_46452,N_46453,N_46454,N_46455,N_46456,N_46457,N_46458,N_46459,N_46460,N_46461,N_46462,N_46463,N_46464,N_46465,N_46466,N_46467,N_46468,N_46469,N_46470,N_46471,N_46472,N_46473,N_46474,N_46475,N_46476,N_46477,N_46478,N_46479,N_46480,N_46481,N_46482,N_46483,N_46484,N_46485,N_46486,N_46487,N_46488,N_46489,N_46490,N_46491,N_46492,N_46493,N_46494,N_46495,N_46496,N_46497,N_46498,N_46499,N_46500,N_46501,N_46502,N_46503,N_46504,N_46505,N_46506,N_46507,N_46508,N_46509,N_46510,N_46511,N_46512,N_46513,N_46514,N_46515,N_46516,N_46517,N_46518,N_46519,N_46520,N_46521,N_46522,N_46523,N_46524,N_46525,N_46526,N_46527,N_46528,N_46529,N_46530,N_46531,N_46532,N_46533,N_46534,N_46535,N_46536,N_46537,N_46538,N_46539,N_46540,N_46541,N_46542,N_46543,N_46544,N_46545,N_46546,N_46547,N_46548,N_46549,N_46550,N_46551,N_46552,N_46553,N_46554,N_46555,N_46556,N_46557,N_46558,N_46559,N_46560,N_46561,N_46562,N_46563,N_46564,N_46565,N_46566,N_46567,N_46568,N_46569,N_46570,N_46571,N_46572,N_46573,N_46574,N_46575,N_46576,N_46577,N_46578,N_46579,N_46580,N_46581,N_46582,N_46583,N_46584,N_46585,N_46586,N_46587,N_46588,N_46589,N_46590,N_46591,N_46592,N_46593,N_46594,N_46595,N_46596,N_46597,N_46598,N_46599,N_46600,N_46601,N_46602,N_46603,N_46604,N_46605,N_46606,N_46607,N_46608,N_46609,N_46610,N_46611,N_46612,N_46613,N_46614,N_46615,N_46616,N_46617,N_46618,N_46619,N_46620,N_46621,N_46622,N_46623,N_46624,N_46625,N_46626,N_46627,N_46628,N_46629,N_46630,N_46631,N_46632,N_46633,N_46634,N_46635,N_46636,N_46637,N_46638,N_46639,N_46640,N_46641,N_46642,N_46643,N_46644,N_46645,N_46646,N_46647,N_46648,N_46649,N_46650,N_46651,N_46652,N_46653,N_46654,N_46655,N_46656,N_46657,N_46658,N_46659,N_46660,N_46661,N_46662,N_46663,N_46664,N_46665,N_46666,N_46667,N_46668,N_46669,N_46670,N_46671,N_46672,N_46673,N_46674,N_46675,N_46676,N_46677,N_46678,N_46679,N_46680,N_46681,N_46682,N_46683,N_46684,N_46685,N_46686,N_46687,N_46688,N_46689,N_46690,N_46691,N_46692,N_46693,N_46694,N_46695,N_46696,N_46697,N_46698,N_46699,N_46700,N_46701,N_46702,N_46703,N_46704,N_46705,N_46706,N_46707,N_46708,N_46709,N_46710,N_46711,N_46712,N_46713,N_46714,N_46715,N_46716,N_46717,N_46718,N_46719,N_46720,N_46721,N_46722,N_46723,N_46724,N_46725,N_46726,N_46727,N_46728,N_46729,N_46730,N_46731,N_46732,N_46733,N_46734,N_46735,N_46736,N_46737,N_46738,N_46739,N_46740,N_46741,N_46742,N_46743,N_46744,N_46745,N_46746,N_46747,N_46748,N_46749,N_46750,N_46751,N_46752,N_46753,N_46754,N_46755,N_46756,N_46757,N_46758,N_46759,N_46760,N_46761,N_46762,N_46763,N_46764,N_46765,N_46766,N_46767,N_46768,N_46769,N_46770,N_46771,N_46772,N_46773,N_46774,N_46775,N_46776,N_46777,N_46778,N_46779,N_46780,N_46781,N_46782,N_46783,N_46784,N_46785,N_46786,N_46787,N_46788,N_46789,N_46790,N_46791,N_46792,N_46793,N_46794,N_46795,N_46796,N_46797,N_46798,N_46799,N_46800,N_46801,N_46802,N_46803,N_46804,N_46805,N_46806,N_46807,N_46808,N_46809,N_46810,N_46811,N_46812,N_46813,N_46814,N_46815,N_46816,N_46817,N_46818,N_46819,N_46820,N_46821,N_46822,N_46823,N_46824,N_46825,N_46826,N_46827,N_46828,N_46829,N_46830,N_46831,N_46832,N_46833,N_46834,N_46835,N_46836,N_46837,N_46838,N_46839,N_46840,N_46841,N_46842,N_46843,N_46844,N_46845,N_46846,N_46847,N_46848,N_46849,N_46850,N_46851,N_46852,N_46853,N_46854,N_46855,N_46856,N_46857,N_46858,N_46859,N_46860,N_46861,N_46862,N_46863,N_46864,N_46865,N_46866,N_46867,N_46868,N_46869,N_46870,N_46871,N_46872,N_46873,N_46874,N_46875,N_46876,N_46877,N_46878,N_46879,N_46880,N_46881,N_46882,N_46883,N_46884,N_46885,N_46886,N_46887,N_46888,N_46889,N_46890,N_46891,N_46892,N_46893,N_46894,N_46895,N_46896,N_46897,N_46898,N_46899,N_46900,N_46901,N_46902,N_46903,N_46904,N_46905,N_46906,N_46907,N_46908,N_46909,N_46910,N_46911,N_46912,N_46913,N_46914,N_46915,N_46916,N_46917,N_46918,N_46919,N_46920,N_46921,N_46922,N_46923,N_46924,N_46925,N_46926,N_46927,N_46928,N_46929,N_46930,N_46931,N_46932,N_46933,N_46934,N_46935,N_46936,N_46937,N_46938,N_46939,N_46940,N_46941,N_46942,N_46943,N_46944,N_46945,N_46946,N_46947,N_46948,N_46949,N_46950,N_46951,N_46952,N_46953,N_46954,N_46955,N_46956,N_46957,N_46958,N_46959,N_46960,N_46961,N_46962,N_46963,N_46964,N_46965,N_46966,N_46967,N_46968,N_46969,N_46970,N_46971,N_46972,N_46973,N_46974,N_46975,N_46976,N_46977,N_46978,N_46979,N_46980,N_46981,N_46982,N_46983,N_46984,N_46985,N_46986,N_46987,N_46988,N_46989,N_46990,N_46991,N_46992,N_46993,N_46994,N_46995,N_46996,N_46997,N_46998,N_46999,N_47000,N_47001,N_47002,N_47003,N_47004,N_47005,N_47006,N_47007,N_47008,N_47009,N_47010,N_47011,N_47012,N_47013,N_47014,N_47015,N_47016,N_47017,N_47018,N_47019,N_47020,N_47021,N_47022,N_47023,N_47024,N_47025,N_47026,N_47027,N_47028,N_47029,N_47030,N_47031,N_47032,N_47033,N_47034,N_47035,N_47036,N_47037,N_47038,N_47039,N_47040,N_47041,N_47042,N_47043,N_47044,N_47045,N_47046,N_47047,N_47048,N_47049,N_47050,N_47051,N_47052,N_47053,N_47054,N_47055,N_47056,N_47057,N_47058,N_47059,N_47060,N_47061,N_47062,N_47063,N_47064,N_47065,N_47066,N_47067,N_47068,N_47069,N_47070,N_47071,N_47072,N_47073,N_47074,N_47075,N_47076,N_47077,N_47078,N_47079,N_47080,N_47081,N_47082,N_47083,N_47084,N_47085,N_47086,N_47087,N_47088,N_47089,N_47090,N_47091,N_47092,N_47093,N_47094,N_47095,N_47096,N_47097,N_47098,N_47099,N_47100,N_47101,N_47102,N_47103,N_47104,N_47105,N_47106,N_47107,N_47108,N_47109,N_47110,N_47111,N_47112,N_47113,N_47114,N_47115,N_47116,N_47117,N_47118,N_47119,N_47120,N_47121,N_47122,N_47123,N_47124,N_47125,N_47126,N_47127,N_47128,N_47129,N_47130,N_47131,N_47132,N_47133,N_47134,N_47135,N_47136,N_47137,N_47138,N_47139,N_47140,N_47141,N_47142,N_47143,N_47144,N_47145,N_47146,N_47147,N_47148,N_47149,N_47150,N_47151,N_47152,N_47153,N_47154,N_47155,N_47156,N_47157,N_47158,N_47159,N_47160,N_47161,N_47162,N_47163,N_47164,N_47165,N_47166,N_47167,N_47168,N_47169,N_47170,N_47171,N_47172,N_47173,N_47174,N_47175,N_47176,N_47177,N_47178,N_47179,N_47180,N_47181,N_47182,N_47183,N_47184,N_47185,N_47186,N_47187,N_47188,N_47189,N_47190,N_47191,N_47192,N_47193,N_47194,N_47195,N_47196,N_47197,N_47198,N_47199,N_47200,N_47201,N_47202,N_47203,N_47204,N_47205,N_47206,N_47207,N_47208,N_47209,N_47210,N_47211,N_47212,N_47213,N_47214,N_47215,N_47216,N_47217,N_47218,N_47219,N_47220,N_47221,N_47222,N_47223,N_47224,N_47225,N_47226,N_47227,N_47228,N_47229,N_47230,N_47231,N_47232,N_47233,N_47234,N_47235,N_47236,N_47237,N_47238,N_47239,N_47240,N_47241,N_47242,N_47243,N_47244,N_47245,N_47246,N_47247,N_47248,N_47249,N_47250,N_47251,N_47252,N_47253,N_47254,N_47255,N_47256,N_47257,N_47258,N_47259,N_47260,N_47261,N_47262,N_47263,N_47264,N_47265,N_47266,N_47267,N_47268,N_47269,N_47270,N_47271,N_47272,N_47273,N_47274,N_47275,N_47276,N_47277,N_47278,N_47279,N_47280,N_47281,N_47282,N_47283,N_47284,N_47285,N_47286,N_47287,N_47288,N_47289,N_47290,N_47291,N_47292,N_47293,N_47294,N_47295,N_47296,N_47297,N_47298,N_47299,N_47300,N_47301,N_47302,N_47303,N_47304,N_47305,N_47306,N_47307,N_47308,N_47309,N_47310,N_47311,N_47312,N_47313,N_47314,N_47315,N_47316,N_47317,N_47318,N_47319,N_47320,N_47321,N_47322,N_47323,N_47324,N_47325,N_47326,N_47327,N_47328,N_47329,N_47330,N_47331,N_47332,N_47333,N_47334,N_47335,N_47336,N_47337,N_47338,N_47339,N_47340,N_47341,N_47342,N_47343,N_47344,N_47345,N_47346,N_47347,N_47348,N_47349,N_47350,N_47351,N_47352,N_47353,N_47354,N_47355,N_47356,N_47357,N_47358,N_47359,N_47360,N_47361,N_47362,N_47363,N_47364,N_47365,N_47366,N_47367,N_47368,N_47369,N_47370,N_47371,N_47372,N_47373,N_47374,N_47375,N_47376,N_47377,N_47378,N_47379,N_47380,N_47381,N_47382,N_47383,N_47384,N_47385,N_47386,N_47387,N_47388,N_47389,N_47390,N_47391,N_47392,N_47393,N_47394,N_47395,N_47396,N_47397,N_47398,N_47399,N_47400,N_47401,N_47402,N_47403,N_47404,N_47405,N_47406,N_47407,N_47408,N_47409,N_47410,N_47411,N_47412,N_47413,N_47414,N_47415,N_47416,N_47417,N_47418,N_47419,N_47420,N_47421,N_47422,N_47423,N_47424,N_47425,N_47426,N_47427,N_47428,N_47429,N_47430,N_47431,N_47432,N_47433,N_47434,N_47435,N_47436,N_47437,N_47438,N_47439,N_47440,N_47441,N_47442,N_47443,N_47444,N_47445,N_47446,N_47447,N_47448,N_47449,N_47450,N_47451,N_47452,N_47453,N_47454,N_47455,N_47456,N_47457,N_47458,N_47459,N_47460,N_47461,N_47462,N_47463,N_47464,N_47465,N_47466,N_47467,N_47468,N_47469,N_47470,N_47471,N_47472,N_47473,N_47474,N_47475,N_47476,N_47477,N_47478,N_47479,N_47480,N_47481,N_47482,N_47483,N_47484,N_47485,N_47486,N_47487,N_47488,N_47489,N_47490,N_47491,N_47492,N_47493,N_47494,N_47495,N_47496,N_47497,N_47498,N_47499,N_47500,N_47501,N_47502,N_47503,N_47504,N_47505,N_47506,N_47507,N_47508,N_47509,N_47510,N_47511,N_47512,N_47513,N_47514,N_47515,N_47516,N_47517,N_47518,N_47519,N_47520,N_47521,N_47522,N_47523,N_47524,N_47525,N_47526,N_47527,N_47528,N_47529,N_47530,N_47531,N_47532,N_47533,N_47534,N_47535,N_47536,N_47537,N_47538,N_47539,N_47540,N_47541,N_47542,N_47543,N_47544,N_47545,N_47546,N_47547,N_47548,N_47549,N_47550,N_47551,N_47552,N_47553,N_47554,N_47555,N_47556,N_47557,N_47558,N_47559,N_47560,N_47561,N_47562,N_47563,N_47564,N_47565,N_47566,N_47567,N_47568,N_47569,N_47570,N_47571,N_47572,N_47573,N_47574,N_47575,N_47576,N_47577,N_47578,N_47579,N_47580,N_47581,N_47582,N_47583,N_47584,N_47585,N_47586,N_47587,N_47588,N_47589,N_47590,N_47591,N_47592,N_47593,N_47594,N_47595,N_47596,N_47597,N_47598,N_47599,N_47600,N_47601,N_47602,N_47603,N_47604,N_47605,N_47606,N_47607,N_47608,N_47609,N_47610,N_47611,N_47612,N_47613,N_47614,N_47615,N_47616,N_47617,N_47618,N_47619,N_47620,N_47621,N_47622,N_47623,N_47624,N_47625,N_47626,N_47627,N_47628,N_47629,N_47630,N_47631,N_47632,N_47633,N_47634,N_47635,N_47636,N_47637,N_47638,N_47639,N_47640,N_47641,N_47642,N_47643,N_47644,N_47645,N_47646,N_47647,N_47648,N_47649,N_47650,N_47651,N_47652,N_47653,N_47654,N_47655,N_47656,N_47657,N_47658,N_47659,N_47660,N_47661,N_47662,N_47663,N_47664,N_47665,N_47666,N_47667,N_47668,N_47669,N_47670,N_47671,N_47672,N_47673,N_47674,N_47675,N_47676,N_47677,N_47678,N_47679,N_47680,N_47681,N_47682,N_47683,N_47684,N_47685,N_47686,N_47687,N_47688,N_47689,N_47690,N_47691,N_47692,N_47693,N_47694,N_47695,N_47696,N_47697,N_47698,N_47699,N_47700,N_47701,N_47702,N_47703,N_47704,N_47705,N_47706,N_47707,N_47708,N_47709,N_47710,N_47711,N_47712,N_47713,N_47714,N_47715,N_47716,N_47717,N_47718,N_47719,N_47720,N_47721,N_47722,N_47723,N_47724,N_47725,N_47726,N_47727,N_47728,N_47729,N_47730,N_47731,N_47732,N_47733,N_47734,N_47735,N_47736,N_47737,N_47738,N_47739,N_47740,N_47741,N_47742,N_47743,N_47744,N_47745,N_47746,N_47747,N_47748,N_47749,N_47750,N_47751,N_47752,N_47753,N_47754,N_47755,N_47756,N_47757,N_47758,N_47759,N_47760,N_47761,N_47762,N_47763,N_47764,N_47765,N_47766,N_47767,N_47768,N_47769,N_47770,N_47771,N_47772,N_47773,N_47774,N_47775,N_47776,N_47777,N_47778,N_47779,N_47780,N_47781,N_47782,N_47783,N_47784,N_47785,N_47786,N_47787,N_47788,N_47789,N_47790,N_47791,N_47792,N_47793,N_47794,N_47795,N_47796,N_47797,N_47798,N_47799,N_47800,N_47801,N_47802,N_47803,N_47804,N_47805,N_47806,N_47807,N_47808,N_47809,N_47810,N_47811,N_47812,N_47813,N_47814,N_47815,N_47816,N_47817,N_47818,N_47819,N_47820,N_47821,N_47822,N_47823,N_47824,N_47825,N_47826,N_47827,N_47828,N_47829,N_47830,N_47831,N_47832,N_47833,N_47834,N_47835,N_47836,N_47837,N_47838,N_47839,N_47840,N_47841,N_47842,N_47843,N_47844,N_47845,N_47846,N_47847,N_47848,N_47849,N_47850,N_47851,N_47852,N_47853,N_47854,N_47855,N_47856,N_47857,N_47858,N_47859,N_47860,N_47861,N_47862,N_47863,N_47864,N_47865,N_47866,N_47867,N_47868,N_47869,N_47870,N_47871,N_47872,N_47873,N_47874,N_47875,N_47876,N_47877,N_47878,N_47879,N_47880,N_47881,N_47882,N_47883,N_47884,N_47885,N_47886,N_47887,N_47888,N_47889,N_47890,N_47891,N_47892,N_47893,N_47894,N_47895,N_47896,N_47897,N_47898,N_47899,N_47900,N_47901,N_47902,N_47903,N_47904,N_47905,N_47906,N_47907,N_47908,N_47909,N_47910,N_47911,N_47912,N_47913,N_47914,N_47915,N_47916,N_47917,N_47918,N_47919,N_47920,N_47921,N_47922,N_47923,N_47924,N_47925,N_47926,N_47927,N_47928,N_47929,N_47930,N_47931,N_47932,N_47933,N_47934,N_47935,N_47936,N_47937,N_47938,N_47939,N_47940,N_47941,N_47942,N_47943,N_47944,N_47945,N_47946,N_47947,N_47948,N_47949,N_47950,N_47951,N_47952,N_47953,N_47954,N_47955,N_47956,N_47957,N_47958,N_47959,N_47960,N_47961,N_47962,N_47963,N_47964,N_47965,N_47966,N_47967,N_47968,N_47969,N_47970,N_47971,N_47972,N_47973,N_47974,N_47975,N_47976,N_47977,N_47978,N_47979,N_47980,N_47981,N_47982,N_47983,N_47984,N_47985,N_47986,N_47987,N_47988,N_47989,N_47990,N_47991,N_47992,N_47993,N_47994,N_47995,N_47996,N_47997,N_47998,N_47999,N_48000,N_48001,N_48002,N_48003,N_48004,N_48005,N_48006,N_48007,N_48008,N_48009,N_48010,N_48011,N_48012,N_48013,N_48014,N_48015,N_48016,N_48017,N_48018,N_48019,N_48020,N_48021,N_48022,N_48023,N_48024,N_48025,N_48026,N_48027,N_48028,N_48029,N_48030,N_48031,N_48032,N_48033,N_48034,N_48035,N_48036,N_48037,N_48038,N_48039,N_48040,N_48041,N_48042,N_48043,N_48044,N_48045,N_48046,N_48047,N_48048,N_48049,N_48050,N_48051,N_48052,N_48053,N_48054,N_48055,N_48056,N_48057,N_48058,N_48059,N_48060,N_48061,N_48062,N_48063,N_48064,N_48065,N_48066,N_48067,N_48068,N_48069,N_48070,N_48071,N_48072,N_48073,N_48074,N_48075,N_48076,N_48077,N_48078,N_48079,N_48080,N_48081,N_48082,N_48083,N_48084,N_48085,N_48086,N_48087,N_48088,N_48089,N_48090,N_48091,N_48092,N_48093,N_48094,N_48095,N_48096,N_48097,N_48098,N_48099,N_48100,N_48101,N_48102,N_48103,N_48104,N_48105,N_48106,N_48107,N_48108,N_48109,N_48110,N_48111,N_48112,N_48113,N_48114,N_48115,N_48116,N_48117,N_48118,N_48119,N_48120,N_48121,N_48122,N_48123,N_48124,N_48125,N_48126,N_48127,N_48128,N_48129,N_48130,N_48131,N_48132,N_48133,N_48134,N_48135,N_48136,N_48137,N_48138,N_48139,N_48140,N_48141,N_48142,N_48143,N_48144,N_48145,N_48146,N_48147,N_48148,N_48149,N_48150,N_48151,N_48152,N_48153,N_48154,N_48155,N_48156,N_48157,N_48158,N_48159,N_48160,N_48161,N_48162,N_48163,N_48164,N_48165,N_48166,N_48167,N_48168,N_48169,N_48170,N_48171,N_48172,N_48173,N_48174,N_48175,N_48176,N_48177,N_48178,N_48179,N_48180,N_48181,N_48182,N_48183,N_48184,N_48185,N_48186,N_48187,N_48188,N_48189,N_48190,N_48191,N_48192,N_48193,N_48194,N_48195,N_48196,N_48197,N_48198,N_48199,N_48200,N_48201,N_48202,N_48203,N_48204,N_48205,N_48206,N_48207,N_48208,N_48209,N_48210,N_48211,N_48212,N_48213,N_48214,N_48215,N_48216,N_48217,N_48218,N_48219,N_48220,N_48221,N_48222,N_48223,N_48224,N_48225,N_48226,N_48227,N_48228,N_48229,N_48230,N_48231,N_48232,N_48233,N_48234,N_48235,N_48236,N_48237,N_48238,N_48239,N_48240,N_48241,N_48242,N_48243,N_48244,N_48245,N_48246,N_48247,N_48248,N_48249,N_48250,N_48251,N_48252,N_48253,N_48254,N_48255,N_48256,N_48257,N_48258,N_48259,N_48260,N_48261,N_48262,N_48263,N_48264,N_48265,N_48266,N_48267,N_48268,N_48269,N_48270,N_48271,N_48272,N_48273,N_48274,N_48275,N_48276,N_48277,N_48278,N_48279,N_48280,N_48281,N_48282,N_48283,N_48284,N_48285,N_48286,N_48287,N_48288,N_48289,N_48290,N_48291,N_48292,N_48293,N_48294,N_48295,N_48296,N_48297,N_48298,N_48299,N_48300,N_48301,N_48302,N_48303,N_48304,N_48305,N_48306,N_48307,N_48308,N_48309,N_48310,N_48311,N_48312,N_48313,N_48314,N_48315,N_48316,N_48317,N_48318,N_48319,N_48320,N_48321,N_48322,N_48323,N_48324,N_48325,N_48326,N_48327,N_48328,N_48329,N_48330,N_48331,N_48332,N_48333,N_48334,N_48335,N_48336,N_48337,N_48338,N_48339,N_48340,N_48341,N_48342,N_48343,N_48344,N_48345,N_48346,N_48347,N_48348,N_48349,N_48350,N_48351,N_48352,N_48353,N_48354,N_48355,N_48356,N_48357,N_48358,N_48359,N_48360,N_48361,N_48362,N_48363,N_48364,N_48365,N_48366,N_48367,N_48368,N_48369,N_48370,N_48371,N_48372,N_48373,N_48374,N_48375,N_48376,N_48377,N_48378,N_48379,N_48380,N_48381,N_48382,N_48383,N_48384,N_48385,N_48386,N_48387,N_48388,N_48389,N_48390,N_48391,N_48392,N_48393,N_48394,N_48395,N_48396,N_48397,N_48398,N_48399,N_48400,N_48401,N_48402,N_48403,N_48404,N_48405,N_48406,N_48407,N_48408,N_48409,N_48410,N_48411,N_48412,N_48413,N_48414,N_48415,N_48416,N_48417,N_48418,N_48419,N_48420,N_48421,N_48422,N_48423,N_48424,N_48425,N_48426,N_48427,N_48428,N_48429,N_48430,N_48431,N_48432,N_48433,N_48434,N_48435,N_48436,N_48437,N_48438,N_48439,N_48440,N_48441,N_48442,N_48443,N_48444,N_48445,N_48446,N_48447,N_48448,N_48449,N_48450,N_48451,N_48452,N_48453,N_48454,N_48455,N_48456,N_48457,N_48458,N_48459,N_48460,N_48461,N_48462,N_48463,N_48464,N_48465,N_48466,N_48467,N_48468,N_48469,N_48470,N_48471,N_48472,N_48473,N_48474,N_48475,N_48476,N_48477,N_48478,N_48479,N_48480,N_48481,N_48482,N_48483,N_48484,N_48485,N_48486,N_48487,N_48488,N_48489,N_48490,N_48491,N_48492,N_48493,N_48494,N_48495,N_48496,N_48497,N_48498,N_48499,N_48500,N_48501,N_48502,N_48503,N_48504,N_48505,N_48506,N_48507,N_48508,N_48509,N_48510,N_48511,N_48512,N_48513,N_48514,N_48515,N_48516,N_48517,N_48518,N_48519,N_48520,N_48521,N_48522,N_48523,N_48524,N_48525,N_48526,N_48527,N_48528,N_48529,N_48530,N_48531,N_48532,N_48533,N_48534,N_48535,N_48536,N_48537,N_48538,N_48539,N_48540,N_48541,N_48542,N_48543,N_48544,N_48545,N_48546,N_48547,N_48548,N_48549,N_48550,N_48551,N_48552,N_48553,N_48554,N_48555,N_48556,N_48557,N_48558,N_48559,N_48560,N_48561,N_48562,N_48563,N_48564,N_48565,N_48566,N_48567,N_48568,N_48569,N_48570,N_48571,N_48572,N_48573,N_48574,N_48575,N_48576,N_48577,N_48578,N_48579,N_48580,N_48581,N_48582,N_48583,N_48584,N_48585,N_48586,N_48587,N_48588,N_48589,N_48590,N_48591,N_48592,N_48593,N_48594,N_48595,N_48596,N_48597,N_48598,N_48599,N_48600,N_48601,N_48602,N_48603,N_48604,N_48605,N_48606,N_48607,N_48608,N_48609,N_48610,N_48611,N_48612,N_48613,N_48614,N_48615,N_48616,N_48617,N_48618,N_48619,N_48620,N_48621,N_48622,N_48623,N_48624,N_48625,N_48626,N_48627,N_48628,N_48629,N_48630,N_48631,N_48632,N_48633,N_48634,N_48635,N_48636,N_48637,N_48638,N_48639,N_48640,N_48641,N_48642,N_48643,N_48644,N_48645,N_48646,N_48647,N_48648,N_48649,N_48650,N_48651,N_48652,N_48653,N_48654,N_48655,N_48656,N_48657,N_48658,N_48659,N_48660,N_48661,N_48662,N_48663,N_48664,N_48665,N_48666,N_48667,N_48668,N_48669,N_48670,N_48671,N_48672,N_48673,N_48674,N_48675,N_48676,N_48677,N_48678,N_48679,N_48680,N_48681,N_48682,N_48683,N_48684,N_48685,N_48686,N_48687,N_48688,N_48689,N_48690,N_48691,N_48692,N_48693,N_48694,N_48695,N_48696,N_48697,N_48698,N_48699,N_48700,N_48701,N_48702,N_48703,N_48704,N_48705,N_48706,N_48707,N_48708,N_48709,N_48710,N_48711,N_48712,N_48713,N_48714,N_48715,N_48716,N_48717,N_48718,N_48719,N_48720,N_48721,N_48722,N_48723,N_48724,N_48725,N_48726,N_48727,N_48728,N_48729,N_48730,N_48731,N_48732,N_48733,N_48734,N_48735,N_48736,N_48737,N_48738,N_48739,N_48740,N_48741,N_48742,N_48743,N_48744,N_48745,N_48746,N_48747,N_48748,N_48749,N_48750,N_48751,N_48752,N_48753,N_48754,N_48755,N_48756,N_48757,N_48758,N_48759,N_48760,N_48761,N_48762,N_48763,N_48764,N_48765,N_48766,N_48767,N_48768,N_48769,N_48770,N_48771,N_48772,N_48773,N_48774,N_48775,N_48776,N_48777,N_48778,N_48779,N_48780,N_48781,N_48782,N_48783,N_48784,N_48785,N_48786,N_48787,N_48788,N_48789,N_48790,N_48791,N_48792,N_48793,N_48794,N_48795,N_48796,N_48797,N_48798,N_48799,N_48800,N_48801,N_48802,N_48803,N_48804,N_48805,N_48806,N_48807,N_48808,N_48809,N_48810,N_48811,N_48812,N_48813,N_48814,N_48815,N_48816,N_48817,N_48818,N_48819,N_48820,N_48821,N_48822,N_48823,N_48824,N_48825,N_48826,N_48827,N_48828,N_48829,N_48830,N_48831,N_48832,N_48833,N_48834,N_48835,N_48836,N_48837,N_48838,N_48839,N_48840,N_48841,N_48842,N_48843,N_48844,N_48845,N_48846,N_48847,N_48848,N_48849,N_48850,N_48851,N_48852,N_48853,N_48854,N_48855,N_48856,N_48857,N_48858,N_48859,N_48860,N_48861,N_48862,N_48863,N_48864,N_48865,N_48866,N_48867,N_48868,N_48869,N_48870,N_48871,N_48872,N_48873,N_48874,N_48875,N_48876,N_48877,N_48878,N_48879,N_48880,N_48881,N_48882,N_48883,N_48884,N_48885,N_48886,N_48887,N_48888,N_48889,N_48890,N_48891,N_48892,N_48893,N_48894,N_48895,N_48896,N_48897,N_48898,N_48899,N_48900,N_48901,N_48902,N_48903,N_48904,N_48905,N_48906,N_48907,N_48908,N_48909,N_48910,N_48911,N_48912,N_48913,N_48914,N_48915,N_48916,N_48917,N_48918,N_48919,N_48920,N_48921,N_48922,N_48923,N_48924,N_48925,N_48926,N_48927,N_48928,N_48929,N_48930,N_48931,N_48932,N_48933,N_48934,N_48935,N_48936,N_48937,N_48938,N_48939,N_48940,N_48941,N_48942,N_48943,N_48944,N_48945,N_48946,N_48947,N_48948,N_48949,N_48950,N_48951,N_48952,N_48953,N_48954,N_48955,N_48956,N_48957,N_48958,N_48959,N_48960,N_48961,N_48962,N_48963,N_48964,N_48965,N_48966,N_48967,N_48968,N_48969,N_48970,N_48971,N_48972,N_48973,N_48974,N_48975,N_48976,N_48977,N_48978,N_48979,N_48980,N_48981,N_48982,N_48983,N_48984,N_48985,N_48986,N_48987,N_48988,N_48989,N_48990,N_48991,N_48992,N_48993,N_48994,N_48995,N_48996,N_48997,N_48998,N_48999,N_49000,N_49001,N_49002,N_49003,N_49004,N_49005,N_49006,N_49007,N_49008,N_49009,N_49010,N_49011,N_49012,N_49013,N_49014,N_49015,N_49016,N_49017,N_49018,N_49019,N_49020,N_49021,N_49022,N_49023,N_49024,N_49025,N_49026,N_49027,N_49028,N_49029,N_49030,N_49031,N_49032,N_49033,N_49034,N_49035,N_49036,N_49037,N_49038,N_49039,N_49040,N_49041,N_49042,N_49043,N_49044,N_49045,N_49046,N_49047,N_49048,N_49049,N_49050,N_49051,N_49052,N_49053,N_49054,N_49055,N_49056,N_49057,N_49058,N_49059,N_49060,N_49061,N_49062,N_49063,N_49064,N_49065,N_49066,N_49067,N_49068,N_49069,N_49070,N_49071,N_49072,N_49073,N_49074,N_49075,N_49076,N_49077,N_49078,N_49079,N_49080,N_49081,N_49082,N_49083,N_49084,N_49085,N_49086,N_49087,N_49088,N_49089,N_49090,N_49091,N_49092,N_49093,N_49094,N_49095,N_49096,N_49097,N_49098,N_49099,N_49100,N_49101,N_49102,N_49103,N_49104,N_49105,N_49106,N_49107,N_49108,N_49109,N_49110,N_49111,N_49112,N_49113,N_49114,N_49115,N_49116,N_49117,N_49118,N_49119,N_49120,N_49121,N_49122,N_49123,N_49124,N_49125,N_49126,N_49127,N_49128,N_49129,N_49130,N_49131,N_49132,N_49133,N_49134,N_49135,N_49136,N_49137,N_49138,N_49139,N_49140,N_49141,N_49142,N_49143,N_49144,N_49145,N_49146,N_49147,N_49148,N_49149,N_49150,N_49151,N_49152,N_49153,N_49154,N_49155,N_49156,N_49157,N_49158,N_49159,N_49160,N_49161,N_49162,N_49163,N_49164,N_49165,N_49166,N_49167,N_49168,N_49169,N_49170,N_49171,N_49172,N_49173,N_49174,N_49175,N_49176,N_49177,N_49178,N_49179,N_49180,N_49181,N_49182,N_49183,N_49184,N_49185,N_49186,N_49187,N_49188,N_49189,N_49190,N_49191,N_49192,N_49193,N_49194,N_49195,N_49196,N_49197,N_49198,N_49199,N_49200,N_49201,N_49202,N_49203,N_49204,N_49205,N_49206,N_49207,N_49208,N_49209,N_49210,N_49211,N_49212,N_49213,N_49214,N_49215,N_49216,N_49217,N_49218,N_49219,N_49220,N_49221,N_49222,N_49223,N_49224,N_49225,N_49226,N_49227,N_49228,N_49229,N_49230,N_49231,N_49232,N_49233,N_49234,N_49235,N_49236,N_49237,N_49238,N_49239,N_49240,N_49241,N_49242,N_49243,N_49244,N_49245,N_49246,N_49247,N_49248,N_49249,N_49250,N_49251,N_49252,N_49253,N_49254,N_49255,N_49256,N_49257,N_49258,N_49259,N_49260,N_49261,N_49262,N_49263,N_49264,N_49265,N_49266,N_49267,N_49268,N_49269,N_49270,N_49271,N_49272,N_49273,N_49274,N_49275,N_49276,N_49277,N_49278,N_49279,N_49280,N_49281,N_49282,N_49283,N_49284,N_49285,N_49286,N_49287,N_49288,N_49289,N_49290,N_49291,N_49292,N_49293,N_49294,N_49295,N_49296,N_49297,N_49298,N_49299,N_49300,N_49301,N_49302,N_49303,N_49304,N_49305,N_49306,N_49307,N_49308,N_49309,N_49310,N_49311,N_49312,N_49313,N_49314,N_49315,N_49316,N_49317,N_49318,N_49319,N_49320,N_49321,N_49322,N_49323,N_49324,N_49325,N_49326,N_49327,N_49328,N_49329,N_49330,N_49331,N_49332,N_49333,N_49334,N_49335,N_49336,N_49337,N_49338,N_49339,N_49340,N_49341,N_49342,N_49343,N_49344,N_49345,N_49346,N_49347,N_49348,N_49349,N_49350,N_49351,N_49352,N_49353,N_49354,N_49355,N_49356,N_49357,N_49358,N_49359,N_49360,N_49361,N_49362,N_49363,N_49364,N_49365,N_49366,N_49367,N_49368,N_49369,N_49370,N_49371,N_49372,N_49373,N_49374,N_49375,N_49376,N_49377,N_49378,N_49379,N_49380,N_49381,N_49382,N_49383,N_49384,N_49385,N_49386,N_49387,N_49388,N_49389,N_49390,N_49391,N_49392,N_49393,N_49394,N_49395,N_49396,N_49397,N_49398,N_49399,N_49400,N_49401,N_49402,N_49403,N_49404,N_49405,N_49406,N_49407,N_49408,N_49409,N_49410,N_49411,N_49412,N_49413,N_49414,N_49415,N_49416,N_49417,N_49418,N_49419,N_49420,N_49421,N_49422,N_49423,N_49424,N_49425,N_49426,N_49427,N_49428,N_49429,N_49430,N_49431,N_49432,N_49433,N_49434,N_49435,N_49436,N_49437,N_49438,N_49439,N_49440,N_49441,N_49442,N_49443,N_49444,N_49445,N_49446,N_49447,N_49448,N_49449,N_49450,N_49451,N_49452,N_49453,N_49454,N_49455,N_49456,N_49457,N_49458,N_49459,N_49460,N_49461,N_49462,N_49463,N_49464,N_49465,N_49466,N_49467,N_49468,N_49469,N_49470,N_49471,N_49472,N_49473,N_49474,N_49475,N_49476,N_49477,N_49478,N_49479,N_49480,N_49481,N_49482,N_49483,N_49484,N_49485,N_49486,N_49487,N_49488,N_49489,N_49490,N_49491,N_49492,N_49493,N_49494,N_49495,N_49496,N_49497,N_49498,N_49499,N_49500,N_49501,N_49502,N_49503,N_49504,N_49505,N_49506,N_49507,N_49508,N_49509,N_49510,N_49511,N_49512,N_49513,N_49514,N_49515,N_49516,N_49517,N_49518,N_49519,N_49520,N_49521,N_49522,N_49523,N_49524,N_49525,N_49526,N_49527,N_49528,N_49529,N_49530,N_49531,N_49532,N_49533,N_49534,N_49535,N_49536,N_49537,N_49538,N_49539,N_49540,N_49541,N_49542,N_49543,N_49544,N_49545,N_49546,N_49547,N_49548,N_49549,N_49550,N_49551,N_49552,N_49553,N_49554,N_49555,N_49556,N_49557,N_49558,N_49559,N_49560,N_49561,N_49562,N_49563,N_49564,N_49565,N_49566,N_49567,N_49568,N_49569,N_49570,N_49571,N_49572,N_49573,N_49574,N_49575,N_49576,N_49577,N_49578,N_49579,N_49580,N_49581,N_49582,N_49583,N_49584,N_49585,N_49586,N_49587,N_49588,N_49589,N_49590,N_49591,N_49592,N_49593,N_49594,N_49595,N_49596,N_49597,N_49598,N_49599,N_49600,N_49601,N_49602,N_49603,N_49604,N_49605,N_49606,N_49607,N_49608,N_49609,N_49610,N_49611,N_49612,N_49613,N_49614,N_49615,N_49616,N_49617,N_49618,N_49619,N_49620,N_49621,N_49622,N_49623,N_49624,N_49625,N_49626,N_49627,N_49628,N_49629,N_49630,N_49631,N_49632,N_49633,N_49634,N_49635,N_49636,N_49637,N_49638,N_49639,N_49640,N_49641,N_49642,N_49643,N_49644,N_49645,N_49646,N_49647,N_49648,N_49649,N_49650,N_49651,N_49652,N_49653,N_49654,N_49655,N_49656,N_49657,N_49658,N_49659,N_49660,N_49661,N_49662,N_49663,N_49664,N_49665,N_49666,N_49667,N_49668,N_49669,N_49670,N_49671,N_49672,N_49673,N_49674,N_49675,N_49676,N_49677,N_49678,N_49679,N_49680,N_49681,N_49682,N_49683,N_49684,N_49685,N_49686,N_49687,N_49688,N_49689,N_49690,N_49691,N_49692,N_49693,N_49694,N_49695,N_49696,N_49697,N_49698,N_49699,N_49700,N_49701,N_49702,N_49703,N_49704,N_49705,N_49706,N_49707,N_49708,N_49709,N_49710,N_49711,N_49712,N_49713,N_49714,N_49715,N_49716,N_49717,N_49718,N_49719,N_49720,N_49721,N_49722,N_49723,N_49724,N_49725,N_49726,N_49727,N_49728,N_49729,N_49730,N_49731,N_49732,N_49733,N_49734,N_49735,N_49736,N_49737,N_49738,N_49739,N_49740,N_49741,N_49742,N_49743,N_49744,N_49745,N_49746,N_49747,N_49748,N_49749,N_49750,N_49751,N_49752,N_49753,N_49754,N_49755,N_49756,N_49757,N_49758,N_49759,N_49760,N_49761,N_49762,N_49763,N_49764,N_49765,N_49766,N_49767,N_49768,N_49769,N_49770,N_49771,N_49772,N_49773,N_49774,N_49775,N_49776,N_49777,N_49778,N_49779,N_49780,N_49781,N_49782,N_49783,N_49784,N_49785,N_49786,N_49787,N_49788,N_49789,N_49790,N_49791,N_49792,N_49793,N_49794,N_49795,N_49796,N_49797,N_49798,N_49799,N_49800,N_49801,N_49802,N_49803,N_49804,N_49805,N_49806,N_49807,N_49808,N_49809,N_49810,N_49811,N_49812,N_49813,N_49814,N_49815,N_49816,N_49817,N_49818,N_49819,N_49820,N_49821,N_49822,N_49823,N_49824,N_49825,N_49826,N_49827,N_49828,N_49829,N_49830,N_49831,N_49832,N_49833,N_49834,N_49835,N_49836,N_49837,N_49838,N_49839,N_49840,N_49841,N_49842,N_49843,N_49844,N_49845,N_49846,N_49847,N_49848,N_49849,N_49850,N_49851,N_49852,N_49853,N_49854,N_49855,N_49856,N_49857,N_49858,N_49859,N_49860,N_49861,N_49862,N_49863,N_49864,N_49865,N_49866,N_49867,N_49868,N_49869,N_49870,N_49871,N_49872,N_49873,N_49874,N_49875,N_49876,N_49877,N_49878,N_49879,N_49880,N_49881,N_49882,N_49883,N_49884,N_49885,N_49886,N_49887,N_49888,N_49889,N_49890,N_49891,N_49892,N_49893,N_49894,N_49895,N_49896,N_49897,N_49898,N_49899,N_49900,N_49901,N_49902,N_49903,N_49904,N_49905,N_49906,N_49907,N_49908,N_49909,N_49910,N_49911,N_49912,N_49913,N_49914,N_49915,N_49916,N_49917,N_49918,N_49919,N_49920,N_49921,N_49922,N_49923,N_49924,N_49925,N_49926,N_49927,N_49928,N_49929,N_49930,N_49931,N_49932,N_49933,N_49934,N_49935,N_49936,N_49937,N_49938,N_49939,N_49940,N_49941,N_49942,N_49943,N_49944,N_49945,N_49946,N_49947,N_49948,N_49949,N_49950,N_49951,N_49952,N_49953,N_49954,N_49955,N_49956,N_49957,N_49958,N_49959,N_49960,N_49961,N_49962,N_49963,N_49964,N_49965,N_49966,N_49967,N_49968,N_49969,N_49970,N_49971,N_49972,N_49973,N_49974,N_49975,N_49976,N_49977,N_49978,N_49979,N_49980,N_49981,N_49982,N_49983,N_49984,N_49985,N_49986,N_49987,N_49988,N_49989,N_49990,N_49991,N_49992,N_49993,N_49994,N_49995,N_49996,N_49997,N_49998,N_49999;
nor U0 (N_0,In_4835,In_4236);
and U1 (N_1,In_4,In_3836);
xnor U2 (N_2,In_4673,In_1062);
xnor U3 (N_3,In_1548,In_724);
or U4 (N_4,In_1534,In_1934);
xnor U5 (N_5,In_4275,In_368);
or U6 (N_6,In_4028,In_4553);
and U7 (N_7,In_837,In_3394);
nor U8 (N_8,In_4576,In_4735);
xor U9 (N_9,In_2765,In_476);
or U10 (N_10,In_1948,In_3084);
xnor U11 (N_11,In_258,In_3045);
or U12 (N_12,In_3414,In_452);
nand U13 (N_13,In_1910,In_4093);
or U14 (N_14,In_4448,In_2516);
and U15 (N_15,In_4387,In_2395);
xnor U16 (N_16,In_1086,In_4014);
nor U17 (N_17,In_1848,In_241);
or U18 (N_18,In_2556,In_4377);
xnor U19 (N_19,In_4975,In_60);
xnor U20 (N_20,In_4375,In_1748);
xnor U21 (N_21,In_4096,In_4364);
xnor U22 (N_22,In_2949,In_3993);
or U23 (N_23,In_982,In_612);
xnor U24 (N_24,In_817,In_3453);
and U25 (N_25,In_4786,In_243);
nand U26 (N_26,In_2122,In_1655);
and U27 (N_27,In_4277,In_2164);
or U28 (N_28,In_751,In_1015);
or U29 (N_29,In_25,In_3495);
nand U30 (N_30,In_687,In_4611);
nor U31 (N_31,In_1726,In_1085);
nor U32 (N_32,In_4089,In_2611);
and U33 (N_33,In_2542,In_94);
and U34 (N_34,In_1866,In_3789);
nor U35 (N_35,In_2734,In_2073);
nor U36 (N_36,In_1629,In_2236);
and U37 (N_37,In_4726,In_4680);
and U38 (N_38,In_1800,In_1365);
nor U39 (N_39,In_3118,In_2958);
xor U40 (N_40,In_2002,In_1354);
and U41 (N_41,In_4694,In_2534);
nand U42 (N_42,In_1865,In_522);
xor U43 (N_43,In_1751,In_2440);
and U44 (N_44,In_1216,In_1831);
and U45 (N_45,In_4797,In_4698);
or U46 (N_46,In_1495,In_2400);
nor U47 (N_47,In_3198,In_1307);
nand U48 (N_48,In_1321,In_75);
and U49 (N_49,In_2485,In_4548);
nand U50 (N_50,In_2904,In_119);
or U51 (N_51,In_3123,In_568);
xnor U52 (N_52,In_3380,In_1049);
or U53 (N_53,In_4727,In_4779);
and U54 (N_54,In_2880,In_402);
and U55 (N_55,In_1101,In_1117);
xnor U56 (N_56,In_4101,In_1839);
or U57 (N_57,In_3982,In_3886);
or U58 (N_58,In_4395,In_3905);
xor U59 (N_59,In_1386,In_664);
or U60 (N_60,In_1297,In_1059);
and U61 (N_61,In_2529,In_922);
nor U62 (N_62,In_4469,In_4037);
xor U63 (N_63,In_1561,In_2367);
and U64 (N_64,In_2599,In_1623);
xor U65 (N_65,In_3041,In_3521);
or U66 (N_66,In_4477,In_973);
xor U67 (N_67,In_3857,In_4487);
nand U68 (N_68,In_2205,In_1290);
nor U69 (N_69,In_1731,In_55);
or U70 (N_70,In_2549,In_1652);
and U71 (N_71,In_3861,In_4449);
xor U72 (N_72,In_4517,In_4730);
nor U73 (N_73,In_64,In_2562);
or U74 (N_74,In_1409,In_2499);
nand U75 (N_75,In_2680,In_380);
nor U76 (N_76,In_2279,In_556);
or U77 (N_77,In_252,In_1581);
xnor U78 (N_78,In_4437,In_1378);
nor U79 (N_79,In_2216,In_1334);
xor U80 (N_80,In_533,In_2274);
nor U81 (N_81,In_2442,In_1919);
and U82 (N_82,In_4356,In_3891);
xnor U83 (N_83,In_2342,In_4272);
nand U84 (N_84,In_1638,In_1033);
nand U85 (N_85,In_797,In_1521);
nor U86 (N_86,In_1802,In_3835);
nand U87 (N_87,In_2891,In_4902);
nand U88 (N_88,In_4290,In_1553);
or U89 (N_89,In_3459,In_355);
xor U90 (N_90,In_4015,In_2736);
nand U91 (N_91,In_1864,In_127);
and U92 (N_92,In_4454,In_941);
or U93 (N_93,In_638,In_705);
xor U94 (N_94,In_4087,In_2494);
nand U95 (N_95,In_4905,In_287);
xnor U96 (N_96,In_4910,In_2139);
or U97 (N_97,In_1654,In_1416);
nor U98 (N_98,In_4333,In_2019);
xor U99 (N_99,In_1302,In_877);
nor U100 (N_100,In_1450,In_2441);
and U101 (N_101,In_914,In_2250);
xnor U102 (N_102,In_1459,In_4651);
nand U103 (N_103,In_1110,In_1202);
or U104 (N_104,In_2692,In_4196);
or U105 (N_105,In_501,In_2851);
and U106 (N_106,In_3865,In_459);
and U107 (N_107,In_3725,In_3846);
or U108 (N_108,In_650,In_1901);
and U109 (N_109,In_2328,In_2349);
nand U110 (N_110,In_4816,In_1468);
nor U111 (N_111,In_2835,In_4580);
and U112 (N_112,In_4497,In_4843);
nand U113 (N_113,In_2003,In_1231);
and U114 (N_114,In_330,In_4251);
nand U115 (N_115,In_3574,In_3633);
nor U116 (N_116,In_165,In_3003);
and U117 (N_117,In_1818,In_3183);
nor U118 (N_118,In_4022,In_3837);
xor U119 (N_119,In_2525,In_177);
nand U120 (N_120,In_1769,In_2746);
or U121 (N_121,In_1860,In_2656);
and U122 (N_122,In_1041,In_2900);
nand U123 (N_123,In_4000,In_4465);
or U124 (N_124,In_2951,In_1328);
and U125 (N_125,In_3570,In_3173);
nand U126 (N_126,In_3433,In_1789);
xnor U127 (N_127,In_2100,In_1929);
nand U128 (N_128,In_998,In_630);
nor U129 (N_129,In_611,In_218);
nor U130 (N_130,In_1192,In_1690);
nand U131 (N_131,In_3566,In_4609);
nand U132 (N_132,In_3538,In_1036);
nand U133 (N_133,In_4436,In_4741);
and U134 (N_134,In_111,In_352);
and U135 (N_135,In_178,In_3243);
xor U136 (N_136,In_4083,In_1146);
or U137 (N_137,In_4309,In_2017);
and U138 (N_138,In_3471,In_3941);
or U139 (N_139,In_3502,In_2940);
and U140 (N_140,In_238,In_482);
xor U141 (N_141,In_1657,In_3553);
or U142 (N_142,In_609,In_3297);
nor U143 (N_143,In_4507,In_980);
nor U144 (N_144,In_2316,In_365);
nor U145 (N_145,In_2532,In_1219);
xnor U146 (N_146,In_688,In_583);
xor U147 (N_147,In_1727,In_4388);
nand U148 (N_148,In_2793,In_3673);
and U149 (N_149,In_4008,In_264);
xnor U150 (N_150,In_72,In_4260);
or U151 (N_151,In_1186,In_1026);
and U152 (N_152,In_700,In_1436);
nor U153 (N_153,In_2283,In_2329);
nor U154 (N_154,In_4760,In_2803);
or U155 (N_155,In_1650,In_3540);
xnor U156 (N_156,In_462,In_3143);
nand U157 (N_157,In_2527,In_3631);
xnor U158 (N_158,In_1568,In_3796);
or U159 (N_159,In_3994,In_3577);
xnor U160 (N_160,In_846,In_879);
nand U161 (N_161,In_3293,In_3388);
xnor U162 (N_162,In_2797,In_3013);
nand U163 (N_163,In_1805,In_1244);
or U164 (N_164,In_1614,In_3845);
nor U165 (N_165,In_3944,In_1298);
nor U166 (N_166,In_843,In_4586);
nor U167 (N_167,In_1473,In_2676);
xor U168 (N_168,In_2051,In_1799);
nand U169 (N_169,In_4860,In_1827);
nor U170 (N_170,In_3511,In_406);
xnor U171 (N_171,In_336,In_666);
nand U172 (N_172,In_613,In_607);
nand U173 (N_173,In_2240,In_2927);
xnor U174 (N_174,In_2536,In_4955);
or U175 (N_175,In_4914,In_320);
and U176 (N_176,In_1317,In_1491);
and U177 (N_177,In_4499,In_4850);
nand U178 (N_178,In_433,In_4683);
nand U179 (N_179,In_2507,In_4931);
nand U180 (N_180,In_3456,In_2854);
or U181 (N_181,In_3662,In_1188);
nor U182 (N_182,In_3814,In_4150);
or U183 (N_183,In_2795,In_4259);
or U184 (N_184,In_421,In_3831);
nand U185 (N_185,In_4949,In_3367);
or U186 (N_186,In_1451,In_2173);
or U187 (N_187,In_2526,In_3762);
nand U188 (N_188,In_4307,In_783);
or U189 (N_189,In_2022,In_1607);
and U190 (N_190,In_3099,In_1278);
nor U191 (N_191,In_67,In_1824);
nor U192 (N_192,In_1045,In_4884);
nor U193 (N_193,In_4614,In_3378);
nand U194 (N_194,In_4861,In_793);
nand U195 (N_195,In_261,In_3605);
and U196 (N_196,In_2109,In_624);
nand U197 (N_197,In_3598,In_2588);
or U198 (N_198,In_1636,In_3206);
nor U199 (N_199,In_4264,In_4799);
xor U200 (N_200,In_4879,In_1464);
nor U201 (N_201,In_2917,In_2052);
nor U202 (N_202,In_1631,In_1640);
nor U203 (N_203,In_2212,In_1388);
xnor U204 (N_204,In_557,In_3693);
nor U205 (N_205,In_2114,In_2956);
nor U206 (N_206,In_3343,In_1132);
and U207 (N_207,In_601,In_2254);
or U208 (N_208,In_784,In_172);
or U209 (N_209,In_4643,In_979);
or U210 (N_210,In_734,In_4193);
and U211 (N_211,In_363,In_2089);
nor U212 (N_212,In_310,In_1257);
nor U213 (N_213,In_2024,In_4568);
nor U214 (N_214,In_1155,In_3800);
and U215 (N_215,In_4827,In_847);
nand U216 (N_216,In_4575,In_2626);
or U217 (N_217,In_471,In_3049);
nor U218 (N_218,In_59,In_3204);
xor U219 (N_219,In_4270,In_1465);
xor U220 (N_220,In_3562,In_4175);
xor U221 (N_221,In_4759,In_1516);
nor U222 (N_222,In_1444,In_2975);
nand U223 (N_223,In_1730,In_2308);
nor U224 (N_224,In_3683,In_2571);
nand U225 (N_225,In_547,In_3780);
xor U226 (N_226,In_3520,In_1904);
and U227 (N_227,In_1108,In_2559);
xor U228 (N_228,In_1747,In_4939);
or U229 (N_229,In_2881,In_4572);
nand U230 (N_230,In_4430,In_3549);
nand U231 (N_231,In_2468,In_649);
and U232 (N_232,In_2300,In_3134);
or U233 (N_233,In_3203,In_3954);
xnor U234 (N_234,In_19,In_3628);
nor U235 (N_235,In_46,In_2210);
or U236 (N_236,In_2397,In_4630);
xor U237 (N_237,In_4645,In_256);
xor U238 (N_238,In_248,In_3496);
or U239 (N_239,In_3341,In_3152);
nor U240 (N_240,In_2932,In_2156);
xor U241 (N_241,In_3799,In_210);
or U242 (N_242,In_4899,In_3641);
and U243 (N_243,In_3498,In_962);
xor U244 (N_244,In_440,In_4045);
nand U245 (N_245,In_1279,In_2276);
xor U246 (N_246,In_1137,In_4709);
xnor U247 (N_247,In_564,In_404);
nand U248 (N_248,In_773,In_1977);
nor U249 (N_249,In_3121,In_1738);
nor U250 (N_250,In_4268,In_1874);
xnor U251 (N_251,In_1234,In_254);
or U252 (N_252,In_3389,In_4114);
and U253 (N_253,In_2084,In_1432);
or U254 (N_254,In_3359,In_2477);
xnor U255 (N_255,In_3019,In_4872);
and U256 (N_256,In_324,In_4577);
xnor U257 (N_257,In_3970,In_4353);
xnor U258 (N_258,In_906,In_3869);
nand U259 (N_259,In_1898,In_904);
or U260 (N_260,In_1849,In_4107);
or U261 (N_261,In_3848,In_1793);
nand U262 (N_262,In_3060,In_253);
nor U263 (N_263,In_1499,In_1859);
nand U264 (N_264,In_1744,In_1618);
nor U265 (N_265,In_1458,In_4561);
xnor U266 (N_266,In_3685,In_3113);
nand U267 (N_267,In_3564,In_3786);
and U268 (N_268,In_3427,In_4832);
xnor U269 (N_269,In_2617,In_483);
and U270 (N_270,In_1850,In_2687);
and U271 (N_271,In_4349,In_3002);
nand U272 (N_272,In_10,In_642);
xnor U273 (N_273,In_1713,In_526);
or U274 (N_274,In_4296,In_2422);
xor U275 (N_275,In_480,In_2597);
or U276 (N_276,In_4891,In_4973);
and U277 (N_277,In_4415,In_593);
xnor U278 (N_278,In_2662,In_2393);
nand U279 (N_279,In_1243,In_1689);
xor U280 (N_280,In_4492,In_745);
xnor U281 (N_281,In_4520,In_105);
nor U282 (N_282,In_1983,In_389);
and U283 (N_283,In_4090,In_1455);
or U284 (N_284,In_3038,In_2812);
nor U285 (N_285,In_1175,In_1274);
nand U286 (N_286,In_2818,In_369);
or U287 (N_287,In_1210,In_2739);
and U288 (N_288,In_4941,In_3147);
and U289 (N_289,In_2213,In_303);
or U290 (N_290,In_3475,In_122);
nor U291 (N_291,In_464,In_911);
xnor U292 (N_292,In_893,In_4221);
and U293 (N_293,In_2501,In_2580);
nor U294 (N_294,In_4235,In_623);
and U295 (N_295,In_4053,In_595);
or U296 (N_296,In_1082,In_167);
and U297 (N_297,In_4758,In_1018);
or U298 (N_298,In_1260,In_2869);
nor U299 (N_299,In_545,In_4153);
nand U300 (N_300,In_4341,In_1665);
nor U301 (N_301,In_663,In_3467);
or U302 (N_302,In_1484,In_3301);
nor U303 (N_303,In_4052,In_2633);
or U304 (N_304,In_822,In_1255);
nand U305 (N_305,In_1489,In_1783);
or U306 (N_306,In_3069,In_2321);
xor U307 (N_307,In_3135,In_2941);
or U308 (N_308,In_2874,In_830);
and U309 (N_309,In_1662,In_3751);
nand U310 (N_310,In_2512,In_4171);
xor U311 (N_311,In_3172,In_65);
nand U312 (N_312,In_3852,In_3919);
or U313 (N_313,In_2303,In_2421);
nand U314 (N_314,In_1902,In_1630);
and U315 (N_315,In_983,In_1111);
and U316 (N_316,In_2685,In_3768);
or U317 (N_317,In_3647,In_1542);
xor U318 (N_318,In_658,In_3110);
and U319 (N_319,In_3357,In_196);
and U320 (N_320,In_1953,In_3724);
and U321 (N_321,In_3138,In_4717);
nand U322 (N_322,In_3534,In_2901);
nand U323 (N_323,In_4599,In_4359);
or U324 (N_324,In_2221,In_2876);
nor U325 (N_325,In_1020,In_631);
and U326 (N_326,In_1011,In_1529);
nand U327 (N_327,In_2798,In_2625);
or U328 (N_328,In_1613,In_283);
nor U329 (N_329,In_1501,In_1217);
or U330 (N_330,In_1995,In_230);
or U331 (N_331,In_2804,In_4386);
and U332 (N_332,In_4968,In_3642);
or U333 (N_333,In_3720,In_3913);
nand U334 (N_334,In_1717,In_990);
or U335 (N_335,In_4502,In_4308);
xor U336 (N_336,In_2664,In_3051);
and U337 (N_337,In_891,In_3925);
or U338 (N_338,In_3573,In_3466);
nor U339 (N_339,In_2668,In_2309);
xnor U340 (N_340,In_2132,In_1959);
xnor U341 (N_341,In_2594,In_63);
xor U342 (N_342,In_4862,In_1265);
or U343 (N_343,In_599,In_3080);
nor U344 (N_344,In_1295,In_3743);
and U345 (N_345,In_2053,In_2569);
and U346 (N_346,In_2161,In_213);
or U347 (N_347,In_3961,In_417);
and U348 (N_348,In_401,In_1421);
nor U349 (N_349,In_3807,In_2032);
and U350 (N_350,In_3844,In_1209);
or U351 (N_351,In_2417,In_407);
or U352 (N_352,In_3980,In_900);
or U353 (N_353,In_3165,In_2402);
xnor U354 (N_354,In_1896,In_3094);
xor U355 (N_355,In_1419,In_3684);
and U356 (N_356,In_1152,In_1387);
nand U357 (N_357,In_4523,In_3105);
nand U358 (N_358,In_2377,In_1212);
nand U359 (N_359,In_3130,In_4423);
nand U360 (N_360,In_2973,In_839);
nor U361 (N_361,In_4740,In_4456);
or U362 (N_362,In_1397,In_3352);
xor U363 (N_363,In_4447,In_1541);
xor U364 (N_364,In_2026,In_3753);
nand U365 (N_365,In_1021,In_2688);
nor U366 (N_366,In_4974,In_1304);
nor U367 (N_367,In_4301,In_4432);
xnor U368 (N_368,In_3216,In_4050);
xor U369 (N_369,In_869,In_3981);
nand U370 (N_370,In_1734,In_1720);
xnor U371 (N_371,In_2751,In_4897);
or U372 (N_372,In_1361,In_1935);
nand U373 (N_373,In_4833,In_1475);
nand U374 (N_374,In_4656,In_3958);
xnor U375 (N_375,In_3976,In_3661);
xnor U376 (N_376,In_225,In_3070);
or U377 (N_377,In_1601,In_2163);
nand U378 (N_378,In_946,In_4682);
or U379 (N_379,In_1504,In_798);
and U380 (N_380,In_1068,In_2256);
and U381 (N_381,In_1347,In_2635);
xnor U382 (N_382,In_4230,In_637);
nor U383 (N_383,In_995,In_437);
nor U384 (N_384,In_463,In_1006);
nand U385 (N_385,In_2238,In_3815);
or U386 (N_386,In_3430,In_2614);
nand U387 (N_387,In_168,In_2777);
xor U388 (N_388,In_2370,In_289);
and U389 (N_389,In_4967,In_2394);
and U390 (N_390,In_2604,In_1206);
nor U391 (N_391,In_2754,In_4451);
xor U392 (N_392,In_1031,In_4648);
xnor U393 (N_393,In_342,In_519);
and U394 (N_394,In_3497,In_386);
nand U395 (N_395,In_3748,In_1315);
nand U396 (N_396,In_2353,In_4420);
and U397 (N_397,In_3372,In_1252);
and U398 (N_398,In_3363,In_3505);
and U399 (N_399,In_4882,In_3331);
and U400 (N_400,In_854,In_3667);
nand U401 (N_401,In_2711,In_2574);
or U402 (N_402,In_3851,In_3047);
nor U403 (N_403,In_1215,In_4635);
or U404 (N_404,In_1410,In_2060);
and U405 (N_405,In_1514,In_3530);
nor U406 (N_406,In_3254,In_1166);
and U407 (N_407,In_3756,In_181);
xor U408 (N_408,In_1988,In_4770);
or U409 (N_409,In_4687,In_2607);
nand U410 (N_410,In_3075,In_1233);
or U411 (N_411,In_8,In_373);
nor U412 (N_412,In_1920,In_2272);
or U413 (N_413,In_1582,In_1782);
xnor U414 (N_414,In_4753,In_3499);
nand U415 (N_415,In_1594,In_1398);
and U416 (N_416,In_3847,In_2262);
nand U417 (N_417,In_1362,In_2027);
or U418 (N_418,In_226,In_4393);
nor U419 (N_419,In_2416,In_2769);
nand U420 (N_420,In_2641,In_4329);
or U421 (N_421,In_1998,In_4564);
nor U422 (N_422,In_931,In_222);
and U423 (N_423,In_2552,In_4528);
nor U424 (N_424,In_2045,In_4746);
nor U425 (N_425,In_2282,In_2521);
or U426 (N_426,In_2472,In_3864);
nor U427 (N_427,In_430,In_313);
and U428 (N_428,In_803,In_236);
or U429 (N_429,In_4311,In_4267);
or U430 (N_430,In_2919,In_151);
nand U431 (N_431,In_4453,In_1449);
nor U432 (N_432,In_4594,In_835);
nor U433 (N_433,In_2697,In_2581);
xnor U434 (N_434,In_1722,In_2816);
nor U435 (N_435,In_4152,In_3569);
or U436 (N_436,In_1970,In_275);
nand U437 (N_437,In_4410,In_3151);
xnor U438 (N_438,In_3101,In_1861);
xnor U439 (N_439,In_938,In_3665);
nand U440 (N_440,In_543,In_1885);
nand U441 (N_441,In_1299,In_2177);
nor U442 (N_442,In_422,In_2206);
and U443 (N_443,In_274,In_1550);
or U444 (N_444,In_2101,In_1723);
nor U445 (N_445,In_3531,In_3606);
and U446 (N_446,In_4084,In_617);
and U447 (N_447,In_2194,In_1711);
nand U448 (N_448,In_2341,In_3504);
xnor U449 (N_449,In_3898,In_3649);
nor U450 (N_450,In_3462,In_4186);
and U451 (N_451,In_184,In_2431);
nor U452 (N_452,In_3445,In_2568);
or U453 (N_453,In_3171,In_2129);
nor U454 (N_454,In_1170,In_197);
xor U455 (N_455,In_4757,In_1537);
or U456 (N_456,In_2930,In_1509);
xor U457 (N_457,In_4320,In_738);
nand U458 (N_458,In_3251,In_654);
nand U459 (N_459,In_4701,In_2064);
and U460 (N_460,In_124,In_4640);
and U461 (N_461,In_2371,In_1395);
nor U462 (N_462,In_1172,In_2235);
xnor U463 (N_463,In_4848,In_3654);
or U464 (N_464,In_3938,In_3578);
nor U465 (N_465,In_1570,In_3821);
xnor U466 (N_466,In_1057,In_2879);
xor U467 (N_467,In_36,In_3804);
nand U468 (N_468,In_1051,In_272);
nand U469 (N_469,In_4488,In_360);
xnor U470 (N_470,In_2922,In_3512);
xnor U471 (N_471,In_1169,In_2140);
xnor U472 (N_472,In_2075,In_1060);
xor U473 (N_473,In_3346,In_192);
and U474 (N_474,In_2510,In_4321);
or U475 (N_475,In_2085,In_2498);
nand U476 (N_476,In_903,In_2506);
and U477 (N_477,In_4531,In_2942);
or U478 (N_478,In_1968,In_3207);
and U479 (N_479,In_3387,In_1496);
or U480 (N_480,In_244,In_4143);
and U481 (N_481,In_769,In_145);
nand U482 (N_482,In_4007,In_2373);
xor U483 (N_483,In_2915,In_2304);
or U484 (N_484,In_4178,In_2771);
and U485 (N_485,In_1808,In_1807);
and U486 (N_486,In_4475,In_51);
or U487 (N_487,In_502,In_234);
xor U488 (N_488,In_2106,In_4570);
and U489 (N_489,In_308,In_2558);
xor U490 (N_490,In_214,In_1389);
xnor U491 (N_491,In_4650,In_3421);
nand U492 (N_492,In_864,In_2670);
xnor U493 (N_493,In_1492,In_2091);
nand U494 (N_494,In_4159,In_2450);
and U495 (N_495,In_1912,In_1435);
nand U496 (N_496,In_4039,In_2030);
and U497 (N_497,In_71,In_2155);
nor U498 (N_498,In_3150,In_413);
xor U499 (N_499,In_4422,In_2957);
and U500 (N_500,In_2162,In_87);
or U501 (N_501,In_4722,In_3524);
or U502 (N_502,In_4878,In_600);
nand U503 (N_503,In_4444,In_4498);
xnor U504 (N_504,In_4241,In_2258);
and U505 (N_505,In_4670,In_4092);
xnor U506 (N_506,In_2249,In_756);
xor U507 (N_507,In_2227,In_2492);
or U508 (N_508,In_4486,In_940);
and U509 (N_509,In_559,In_58);
xor U510 (N_510,In_4997,In_2679);
nand U511 (N_511,In_4795,In_575);
or U512 (N_512,In_4985,In_2035);
xor U513 (N_513,In_2288,In_2652);
or U514 (N_514,In_2575,In_3360);
nor U515 (N_515,In_3491,In_393);
nand U516 (N_516,In_43,In_3160);
xnor U517 (N_517,In_1448,In_2307);
and U518 (N_518,In_3650,In_4086);
or U519 (N_519,In_3373,In_2518);
nor U520 (N_520,In_942,In_4242);
or U521 (N_521,In_4592,In_3419);
or U522 (N_522,In_3434,In_1580);
nor U523 (N_523,In_1645,In_808);
and U524 (N_524,In_850,In_4177);
xnor U525 (N_525,In_1044,In_15);
nor U526 (N_526,In_2385,In_4217);
nand U527 (N_527,In_4384,In_3021);
nand U528 (N_528,In_4204,In_3872);
xnor U529 (N_529,In_4831,In_3644);
or U530 (N_530,In_4712,In_3256);
xor U531 (N_531,In_1034,In_810);
nand U532 (N_532,In_974,In_2619);
xnor U533 (N_533,In_2331,In_1074);
nand U534 (N_534,In_3714,In_154);
or U535 (N_535,In_2115,In_1167);
nor U536 (N_536,In_1566,In_3407);
and U537 (N_537,In_3877,In_910);
and U538 (N_538,In_4538,In_4646);
and U539 (N_539,In_2744,In_2128);
xnor U540 (N_540,In_1200,In_766);
xor U541 (N_541,In_4482,In_1527);
xor U542 (N_542,In_520,In_2742);
xnor U543 (N_543,In_113,In_1054);
or U544 (N_544,In_2201,In_1346);
nand U545 (N_545,In_1426,In_3653);
xor U546 (N_546,In_189,In_129);
and U547 (N_547,In_3006,In_2465);
xor U548 (N_548,In_1691,In_3985);
nand U549 (N_549,In_4644,In_1375);
nor U550 (N_550,In_3943,In_4059);
or U551 (N_551,In_3232,In_721);
nor U552 (N_552,In_3237,In_1836);
nand U553 (N_553,In_2346,In_2148);
nand U554 (N_554,In_1164,In_3303);
or U555 (N_555,In_95,In_3563);
and U556 (N_556,In_2996,In_3858);
or U557 (N_557,In_1430,In_2425);
xnor U558 (N_558,In_3946,In_4794);
nor U559 (N_559,In_1014,In_390);
xor U560 (N_560,In_4442,In_2924);
nand U561 (N_561,In_2716,In_3048);
or U562 (N_562,In_4252,In_1797);
xor U563 (N_563,In_4243,In_1149);
nand U564 (N_564,In_1179,In_3518);
or U565 (N_565,In_795,In_2301);
and U566 (N_566,In_3067,In_4881);
xnor U567 (N_567,In_2447,In_4261);
xnor U568 (N_568,In_2124,In_2735);
and U569 (N_569,In_490,In_3826);
or U570 (N_570,In_913,In_4280);
xor U571 (N_571,In_985,In_1900);
or U572 (N_572,In_2523,In_4514);
nor U573 (N_573,In_4291,In_4414);
nor U574 (N_574,In_4334,In_4559);
xor U575 (N_575,In_674,In_2399);
nand U576 (N_576,In_1879,In_626);
and U577 (N_577,In_2583,In_2590);
or U578 (N_578,In_2467,In_1284);
xor U579 (N_579,In_2151,In_3064);
nand U580 (N_580,In_2196,In_4339);
nand U581 (N_581,In_2601,In_4540);
nor U582 (N_582,In_2598,In_3140);
xnor U583 (N_583,In_4549,In_1000);
and U584 (N_584,In_2189,In_1143);
or U585 (N_585,In_4147,In_1724);
nand U586 (N_586,In_3690,In_3175);
xor U587 (N_587,In_1293,In_4588);
nor U588 (N_588,In_2449,In_3537);
or U589 (N_589,In_130,In_1966);
nand U590 (N_590,In_3744,In_1767);
and U591 (N_591,In_44,In_4214);
nor U592 (N_592,In_3432,In_4238);
nor U593 (N_593,In_3109,In_4470);
nor U594 (N_594,In_4773,In_3774);
or U595 (N_595,In_761,In_269);
and U596 (N_596,In_4711,In_3735);
nor U597 (N_597,In_206,In_2411);
xnor U598 (N_598,In_1575,In_3882);
and U599 (N_599,In_2634,In_29);
nor U600 (N_600,In_200,In_1370);
xor U601 (N_601,In_2675,In_706);
nand U602 (N_602,In_4943,In_4710);
nand U603 (N_603,In_3766,In_2119);
and U604 (N_604,In_195,In_529);
and U605 (N_605,In_3991,In_323);
nand U606 (N_606,In_343,In_4637);
and U607 (N_607,In_2678,In_695);
nand U608 (N_608,In_2585,In_1829);
nor U609 (N_609,In_2454,In_2537);
xor U610 (N_610,In_2630,In_957);
nand U611 (N_611,In_2600,In_3881);
nor U612 (N_612,In_659,In_3014);
xnor U613 (N_613,In_579,In_1471);
xnor U614 (N_614,In_4121,In_3458);
and U615 (N_615,In_1335,In_1394);
nor U616 (N_616,In_128,In_1547);
or U617 (N_617,In_295,In_1620);
nand U618 (N_618,In_3745,In_4777);
and U619 (N_619,In_4809,In_3104);
and U620 (N_620,In_1809,In_827);
xor U621 (N_621,In_3945,In_4441);
xnor U622 (N_622,In_2923,In_3694);
nor U623 (N_623,In_3486,In_4621);
nor U624 (N_624,In_3268,In_2497);
and U625 (N_625,In_37,In_1453);
nor U626 (N_626,In_4647,In_629);
xnor U627 (N_627,In_1076,In_3555);
and U628 (N_628,In_585,In_3349);
nand U629 (N_629,In_3634,In_918);
or U630 (N_630,In_3261,In_799);
xor U631 (N_631,In_2759,In_2302);
xnor U632 (N_632,In_3782,In_4960);
nand U633 (N_633,In_657,In_375);
or U634 (N_634,In_2178,In_4871);
xor U635 (N_635,In_2853,In_1753);
and U636 (N_636,In_4825,In_831);
nor U637 (N_637,In_4697,In_1229);
and U638 (N_638,In_4129,In_481);
and U639 (N_639,In_3733,In_584);
nor U640 (N_640,In_1693,In_3613);
or U641 (N_641,In_1437,In_2237);
nand U642 (N_642,In_1123,In_1945);
or U643 (N_643,In_1355,In_2931);
and U644 (N_644,In_2561,In_2884);
or U645 (N_645,In_2348,In_1563);
and U646 (N_646,In_1798,In_1506);
or U647 (N_647,In_3100,In_4027);
xnor U648 (N_648,In_2865,In_1562);
nand U649 (N_649,In_1942,In_3600);
nor U650 (N_650,In_1616,In_2522);
nor U651 (N_651,In_4344,In_894);
nand U652 (N_652,In_828,In_2145);
xor U653 (N_653,In_1083,In_4842);
nand U654 (N_654,In_1889,In_2961);
and U655 (N_655,In_3179,In_66);
xnor U656 (N_656,In_2723,In_1351);
nor U657 (N_657,In_3565,In_4796);
nand U658 (N_658,In_4731,In_2764);
or U659 (N_659,In_3726,In_4811);
or U660 (N_660,In_4091,In_1940);
or U661 (N_661,In_1413,In_4417);
and U662 (N_662,In_2715,In_1221);
xnor U663 (N_663,In_4357,In_4539);
xor U664 (N_664,In_2573,In_746);
and U665 (N_665,In_4789,In_3377);
nor U666 (N_666,In_1736,In_587);
nor U667 (N_667,In_1096,In_1135);
or U668 (N_668,In_4351,In_2482);
and U669 (N_669,In_2118,In_3180);
or U670 (N_670,In_1423,In_1148);
or U671 (N_671,In_3808,In_1578);
xnor U672 (N_672,In_4763,In_2078);
nor U673 (N_673,In_2544,In_2964);
or U674 (N_674,In_1418,In_691);
and U675 (N_675,In_3765,In_3311);
nor U676 (N_676,In_3238,In_2579);
xnor U677 (N_677,In_1637,In_4220);
xnor U678 (N_678,In_1784,In_1978);
nor U679 (N_679,In_2110,In_2832);
xnor U680 (N_680,In_2248,In_3712);
nand U681 (N_681,In_3603,In_2763);
xnor U682 (N_682,In_4612,In_2123);
and U683 (N_683,In_448,In_3214);
or U684 (N_684,In_3035,In_3812);
or U685 (N_685,In_1224,In_1447);
or U686 (N_686,In_432,In_701);
nor U687 (N_687,In_683,In_1721);
xnor U688 (N_688,In_4889,In_221);
nor U689 (N_689,In_439,In_4046);
nor U690 (N_690,In_3556,In_2244);
nor U691 (N_691,In_1883,In_4323);
and U692 (N_692,In_359,In_4608);
xor U693 (N_693,In_778,In_1180);
nand U694 (N_694,In_731,In_1794);
nand U695 (N_695,In_115,In_70);
xor U696 (N_696,In_3689,In_4073);
and U697 (N_697,In_1815,In_220);
nor U698 (N_698,In_3936,In_1554);
nand U699 (N_699,In_32,In_438);
or U700 (N_700,In_1344,In_2786);
nor U701 (N_701,In_3544,In_1084);
and U702 (N_702,In_4255,In_1162);
or U703 (N_703,In_3587,In_4461);
and U704 (N_704,In_4070,In_4666);
or U705 (N_705,In_4057,In_2709);
and U706 (N_706,In_1228,In_591);
nor U707 (N_707,In_709,In_3304);
and U708 (N_708,In_1482,In_2149);
xor U709 (N_709,In_315,In_2047);
nand U710 (N_710,In_1771,In_3408);
nor U711 (N_711,In_1067,In_732);
or U712 (N_712,In_2470,In_376);
xor U713 (N_713,In_3448,In_212);
xor U714 (N_714,In_3154,In_469);
nor U715 (N_715,In_2902,In_454);
and U716 (N_716,In_748,In_4885);
nor U717 (N_717,In_2570,In_3678);
or U718 (N_718,In_3717,In_3999);
xnor U719 (N_719,In_2136,In_2102);
nand U720 (N_720,In_4226,In_3632);
xor U721 (N_721,In_2265,In_4790);
nand U722 (N_722,In_2717,In_17);
xnor U723 (N_723,In_2311,In_4372);
or U724 (N_724,In_1390,In_662);
or U725 (N_725,In_4049,In_468);
xnor U726 (N_726,In_1880,In_3580);
or U727 (N_727,In_3788,In_3630);
xor U728 (N_728,In_4338,In_730);
xnor U729 (N_729,In_286,In_2821);
and U730 (N_730,In_2489,In_4064);
or U731 (N_731,In_1352,In_774);
xor U732 (N_732,In_3476,In_4034);
nand U733 (N_733,In_1190,In_2143);
and U734 (N_734,In_3004,In_4883);
nor U735 (N_735,In_2705,In_1392);
nor U736 (N_736,In_4729,In_2179);
and U737 (N_737,In_3850,In_3220);
nand U738 (N_738,In_2693,In_3056);
xor U739 (N_739,In_3057,In_428);
xor U740 (N_740,In_3942,In_4693);
and U741 (N_741,In_968,In_3126);
nand U742 (N_742,In_4342,In_3939);
nor U743 (N_743,In_377,In_1688);
or U744 (N_744,In_405,In_3166);
xor U745 (N_745,In_1930,In_4810);
xor U746 (N_746,In_1868,In_2603);
or U747 (N_747,In_535,In_2724);
nor U748 (N_748,In_425,In_1682);
and U749 (N_749,In_3257,In_2657);
nor U750 (N_750,In_4996,In_4040);
nor U751 (N_751,In_1144,In_4139);
and U752 (N_752,In_416,In_3025);
xor U753 (N_753,In_3885,In_4187);
nor U754 (N_754,In_326,In_1651);
and U755 (N_755,In_4340,In_2018);
xnor U756 (N_756,In_4890,In_4596);
and U757 (N_757,In_689,In_3889);
nor U758 (N_758,In_4986,In_4819);
and U759 (N_759,In_1735,In_896);
and U760 (N_760,In_3170,In_1647);
or U761 (N_761,In_558,In_3679);
xnor U762 (N_762,In_2937,In_2142);
nor U763 (N_763,In_2990,In_62);
and U764 (N_764,In_4294,In_561);
and U765 (N_765,In_2520,In_1109);
xor U766 (N_766,In_1174,In_4616);
nand U767 (N_767,In_265,In_1916);
nand U768 (N_768,In_1120,In_497);
and U769 (N_769,In_3169,In_97);
nor U770 (N_770,In_3398,In_2352);
nand U771 (N_771,In_4555,In_3440);
nand U772 (N_772,In_2092,In_3589);
xnor U773 (N_773,In_2551,In_3092);
or U774 (N_774,In_2296,In_4380);
nand U775 (N_775,In_1826,In_340);
nand U776 (N_776,In_250,In_565);
xnor U777 (N_777,In_2407,In_1586);
xnor U778 (N_778,In_3132,In_4163);
nor U779 (N_779,In_3975,In_3757);
xnor U780 (N_780,In_3167,In_961);
nand U781 (N_781,In_1584,In_45);
xnor U782 (N_782,In_888,In_3273);
nor U783 (N_783,In_3584,In_2491);
xnor U784 (N_784,In_1705,In_4203);
and U785 (N_785,In_932,In_4081);
and U786 (N_786,In_3288,In_3722);
xor U787 (N_787,In_4946,In_1539);
nand U788 (N_788,In_2883,In_2538);
and U789 (N_789,In_306,In_158);
and U790 (N_790,In_4390,In_1574);
and U791 (N_791,In_106,In_2955);
and U792 (N_792,In_3397,In_4589);
or U793 (N_793,In_1673,In_4133);
xnor U794 (N_794,In_3670,In_4452);
nand U795 (N_795,In_3483,In_1979);
or U796 (N_796,In_1037,In_3455);
nor U797 (N_797,In_4865,In_892);
and U798 (N_798,In_1405,In_3697);
nor U799 (N_799,In_50,In_4745);
xor U800 (N_800,In_4172,In_1127);
nor U801 (N_801,In_2637,In_276);
xor U802 (N_802,In_4613,In_2892);
nand U803 (N_803,In_1565,In_2627);
nor U804 (N_804,In_1207,In_2255);
nor U805 (N_805,In_1081,In_4992);
nand U806 (N_806,In_3155,In_419);
nand U807 (N_807,In_4641,In_4058);
and U808 (N_808,In_2391,In_3318);
nor U809 (N_809,In_1768,In_4667);
or U810 (N_810,In_1258,In_1320);
and U811 (N_811,In_825,In_3874);
nor U812 (N_812,In_1030,In_2040);
xor U813 (N_813,In_4500,In_1947);
or U814 (N_814,In_4804,In_3503);
xor U815 (N_815,In_2935,In_2661);
and U816 (N_816,In_991,In_2197);
or U817 (N_817,In_3390,In_2058);
nand U818 (N_818,In_123,In_2191);
xor U819 (N_819,In_771,In_2010);
nor U820 (N_820,In_765,In_398);
nor U821 (N_821,In_4285,In_887);
or U822 (N_822,In_1262,In_1399);
nand U823 (N_823,In_3,In_872);
nor U824 (N_824,In_1254,In_3674);
and U825 (N_825,In_633,In_4527);
or U826 (N_826,In_2840,In_3820);
nor U827 (N_827,In_1589,In_2609);
xnor U828 (N_828,In_494,In_1967);
or U829 (N_829,In_152,In_92);
xor U830 (N_830,In_2807,In_4684);
or U831 (N_831,In_3963,In_3356);
nand U832 (N_832,In_1598,In_3305);
or U833 (N_833,In_2671,In_4006);
nand U834 (N_834,In_928,In_4298);
and U835 (N_835,In_1749,In_4677);
nand U836 (N_836,In_4003,In_4700);
and U837 (N_837,In_2438,In_201);
xor U838 (N_838,In_101,In_1204);
nor U839 (N_839,In_133,In_2673);
nor U840 (N_840,In_4085,In_1671);
nor U841 (N_841,In_68,In_4579);
and U842 (N_842,In_754,In_1222);
nor U843 (N_843,In_4013,In_4713);
and U844 (N_844,In_53,In_1203);
and U845 (N_845,In_1326,In_2374);
nand U846 (N_846,In_1684,In_4043);
nand U847 (N_847,In_4714,In_4544);
or U848 (N_848,In_1851,In_3809);
or U849 (N_849,In_4971,In_1237);
and U850 (N_850,In_4945,In_965);
nor U851 (N_851,In_4106,In_760);
or U852 (N_852,In_2056,In_592);
nand U853 (N_853,In_1974,In_988);
or U854 (N_854,In_905,In_1938);
nor U855 (N_855,In_73,In_34);
nand U856 (N_856,In_2785,In_857);
and U857 (N_857,In_4915,In_1404);
nand U858 (N_858,In_3107,In_2322);
and U859 (N_859,In_4348,In_4389);
nor U860 (N_860,In_4199,In_3984);
nand U861 (N_861,In_2753,In_3708);
and U862 (N_862,In_3543,In_1070);
or U863 (N_863,In_902,In_298);
and U864 (N_864,In_26,In_4661);
or U865 (N_865,In_3810,In_552);
and U866 (N_866,In_3005,In_4761);
and U867 (N_867,In_4210,In_1716);
xnor U868 (N_868,In_1066,In_229);
nor U869 (N_869,In_4855,In_4715);
nand U870 (N_870,In_1991,In_4625);
xor U871 (N_871,In_3127,In_3468);
xnor U872 (N_872,In_4654,In_3721);
nor U873 (N_873,In_2200,In_1211);
and U874 (N_874,In_1884,In_4148);
nand U875 (N_875,In_4102,In_4183);
or U876 (N_876,In_3230,In_333);
or U877 (N_877,In_137,In_2553);
xor U878 (N_878,In_2423,In_1245);
or U879 (N_879,In_1545,In_3046);
and U880 (N_880,In_2690,In_2667);
nand U881 (N_881,In_544,In_396);
or U882 (N_882,In_4913,In_1596);
nor U883 (N_883,In_54,In_3731);
xor U884 (N_884,In_460,In_3507);
nor U885 (N_885,In_1825,In_4173);
and U886 (N_886,In_4060,In_4462);
and U887 (N_887,In_786,In_1381);
or U888 (N_888,In_3111,In_596);
nand U889 (N_889,In_3489,In_4407);
or U890 (N_890,In_1002,In_2718);
and U891 (N_891,In_2299,In_82);
nand U892 (N_892,In_2211,In_2948);
nor U893 (N_893,In_3802,In_2228);
or U894 (N_894,In_3374,In_1733);
or U895 (N_895,In_2806,In_1551);
nor U896 (N_896,In_3451,In_3250);
xnor U897 (N_897,In_3282,In_672);
xor U898 (N_898,In_1954,In_458);
or U899 (N_899,In_125,In_4869);
nand U900 (N_900,In_3535,In_3755);
or U901 (N_901,In_569,In_3205);
nor U902 (N_902,In_1071,In_3116);
nand U903 (N_903,In_2747,In_3701);
xor U904 (N_904,In_840,In_3443);
xor U905 (N_905,In_3516,In_2207);
xnor U906 (N_906,In_2192,In_4231);
xnor U907 (N_907,In_4299,In_4877);
nor U908 (N_908,In_537,In_2513);
nand U909 (N_909,In_3416,In_3449);
and U910 (N_910,In_4398,In_4021);
xnor U911 (N_911,In_3490,In_4911);
nor U912 (N_912,In_4858,In_2648);
and U913 (N_913,In_3385,In_2672);
nor U914 (N_914,In_4979,In_3907);
nand U915 (N_915,In_1754,In_3671);
nand U916 (N_916,In_3302,In_994);
and U917 (N_917,In_1316,In_1177);
nand U918 (N_918,In_1095,In_532);
and U919 (N_919,In_2219,In_187);
nand U920 (N_920,In_4557,In_199);
xnor U921 (N_921,In_4581,In_1525);
or U922 (N_922,In_327,In_3623);
and U923 (N_923,In_3321,In_4513);
xor U924 (N_924,In_39,In_3062);
xnor U925 (N_925,In_2995,In_1532);
or U926 (N_926,In_959,In_1625);
nor U927 (N_927,In_3369,In_834);
nand U928 (N_928,In_4179,In_3568);
xor U929 (N_929,In_1877,In_1530);
nor U930 (N_930,In_3727,In_4847);
nand U931 (N_931,In_3880,In_1992);
or U932 (N_932,In_4278,In_2455);
and U933 (N_933,In_3262,In_3020);
or U934 (N_934,In_643,In_1440);
or U935 (N_935,In_1745,In_1876);
nor U936 (N_936,In_3995,In_2330);
xnor U937 (N_937,In_3910,In_3236);
or U938 (N_938,In_3229,In_1323);
or U939 (N_939,In_4888,In_2169);
or U940 (N_940,In_1795,In_4781);
and U941 (N_941,In_2981,In_4649);
nor U942 (N_942,In_1053,In_2475);
nand U943 (N_943,In_4747,In_2934);
xnor U944 (N_944,In_1820,In_1844);
or U945 (N_945,In_4483,In_2141);
and U946 (N_946,In_232,In_3415);
xnor U947 (N_947,In_3645,In_2595);
nor U948 (N_948,In_3139,In_2315);
and U949 (N_949,In_2589,In_2669);
nor U950 (N_950,In_3749,In_3191);
xor U951 (N_951,In_3217,In_2896);
xor U952 (N_952,In_3652,In_1380);
xnor U953 (N_953,In_4663,In_2545);
or U954 (N_954,In_950,In_81);
and U955 (N_955,In_142,In_2749);
nor U956 (N_956,In_1025,In_3798);
xnor U957 (N_957,In_1310,In_3921);
nor U958 (N_958,In_1124,In_4304);
nand U959 (N_959,In_1704,In_489);
nor U960 (N_960,In_2025,In_690);
xor U961 (N_961,In_2560,In_2278);
nor U962 (N_962,In_4194,In_4368);
nand U963 (N_963,In_1376,In_371);
and U964 (N_964,In_2287,In_3931);
xor U965 (N_965,In_1439,In_2419);
nand U966 (N_966,In_4273,In_148);
nand U967 (N_967,In_245,In_4036);
xor U968 (N_968,In_4585,In_1976);
or U969 (N_969,In_1515,In_2469);
and U970 (N_970,In_4957,In_4868);
nand U971 (N_971,In_4510,In_1488);
nor U972 (N_972,In_312,In_4736);
nor U973 (N_973,In_3669,In_3300);
nand U974 (N_974,In_3771,In_3319);
and U975 (N_975,In_1357,In_1077);
nor U976 (N_976,In_3940,In_934);
nor U977 (N_977,In_1341,In_249);
and U978 (N_978,In_2639,In_1579);
and U979 (N_979,In_3265,In_4041);
nand U980 (N_980,In_4062,In_4893);
or U981 (N_981,In_2356,In_1664);
and U982 (N_982,In_1564,In_4319);
or U983 (N_983,In_2490,In_1855);
and U984 (N_984,In_499,In_1632);
and U985 (N_985,In_2770,In_1813);
or U986 (N_986,In_61,In_2713);
and U987 (N_987,In_2350,In_2760);
nand U988 (N_988,In_2737,In_1427);
and U989 (N_989,In_4851,In_841);
and U990 (N_990,In_3221,In_865);
nand U991 (N_991,In_614,In_3406);
nor U992 (N_992,In_4489,In_3576);
or U993 (N_993,In_3554,In_3575);
nand U994 (N_994,In_3244,In_2071);
or U995 (N_995,In_1707,In_372);
and U996 (N_996,In_4829,In_4657);
nand U997 (N_997,In_4920,In_2405);
nor U998 (N_998,In_3093,In_4964);
and U999 (N_999,In_2738,In_257);
nand U1000 (N_1000,In_2677,In_2659);
xor U1001 (N_1001,In_3866,In_4257);
nand U1002 (N_1002,In_2007,In_3264);
and U1003 (N_1003,In_4282,In_3839);
xnor U1004 (N_1004,In_3044,In_3868);
nand U1005 (N_1005,In_878,In_972);
xor U1006 (N_1006,In_3522,In_3876);
nand U1007 (N_1007,In_1016,In_3842);
and U1008 (N_1008,In_1642,In_1445);
and U1009 (N_1009,In_3436,In_1615);
nor U1010 (N_1010,In_2345,In_1396);
nor U1011 (N_1011,In_2247,In_4854);
and U1012 (N_1012,In_2241,In_3849);
xor U1013 (N_1013,In_727,In_1588);
nor U1014 (N_1014,In_3635,In_4343);
and U1015 (N_1015,In_4126,In_1743);
nor U1016 (N_1016,In_3494,In_907);
nor U1017 (N_1017,In_2277,In_2230);
nor U1018 (N_1018,In_970,In_1699);
or U1019 (N_1019,In_4189,In_3284);
nor U1020 (N_1020,In_4864,In_38);
nand U1021 (N_1021,In_3235,In_4327);
or U1022 (N_1022,In_2044,In_920);
xor U1023 (N_1023,In_2910,In_3681);
or U1024 (N_1024,In_3953,In_3286);
nand U1025 (N_1025,In_1189,In_1780);
and U1026 (N_1026,In_3480,In_1941);
nand U1027 (N_1027,In_3000,In_2847);
nor U1028 (N_1028,In_3960,In_1055);
nor U1029 (N_1029,In_4485,In_2343);
nor U1030 (N_1030,In_2584,In_138);
nand U1031 (N_1031,In_925,In_2415);
xor U1032 (N_1032,In_2540,In_3883);
xor U1033 (N_1033,In_1533,In_1417);
or U1034 (N_1034,In_4567,In_4426);
nor U1035 (N_1035,In_2001,In_1811);
or U1036 (N_1036,In_2243,In_640);
xnor U1037 (N_1037,In_2293,In_3792);
or U1038 (N_1038,In_636,In_577);
nand U1039 (N_1039,In_652,In_4734);
nor U1040 (N_1040,In_4120,In_668);
nand U1041 (N_1041,In_694,In_3734);
xnor U1042 (N_1042,In_4167,In_3085);
and U1043 (N_1043,In_1814,In_311);
nor U1044 (N_1044,In_2741,In_3601);
or U1045 (N_1045,In_1643,In_2566);
xnor U1046 (N_1046,In_370,In_3382);
nand U1047 (N_1047,In_4875,In_2871);
xor U1048 (N_1048,In_3894,In_40);
nand U1049 (N_1049,In_4306,In_3732);
xnor U1050 (N_1050,In_2029,In_1700);
and U1051 (N_1051,In_3089,In_362);
or U1052 (N_1052,In_2339,In_291);
nand U1053 (N_1053,In_1787,In_3423);
xnor U1054 (N_1054,In_485,In_3627);
and U1055 (N_1055,In_2466,In_3509);
nand U1056 (N_1056,In_4468,In_3365);
xnor U1057 (N_1057,In_4109,In_3296);
nor U1058 (N_1058,In_3951,In_52);
nand U1059 (N_1059,In_1840,In_2624);
nor U1060 (N_1060,In_2722,In_2993);
xor U1061 (N_1061,In_802,In_1706);
nor U1062 (N_1062,In_4728,In_2121);
xor U1063 (N_1063,In_4969,In_1989);
or U1064 (N_1064,In_4841,In_3884);
xnor U1065 (N_1065,In_4530,In_4947);
or U1066 (N_1066,In_1158,In_1519);
xnor U1067 (N_1067,In_509,In_3283);
nor U1068 (N_1068,In_4679,In_477);
xor U1069 (N_1069,In_4922,In_2253);
nand U1070 (N_1070,In_472,In_3193);
nand U1071 (N_1071,In_2808,In_3240);
nand U1072 (N_1072,In_1567,In_1403);
and U1073 (N_1073,In_3911,In_1138);
nand U1074 (N_1074,In_2689,In_3770);
or U1075 (N_1075,In_4970,In_923);
nor U1076 (N_1076,In_3055,In_3822);
or U1077 (N_1077,In_733,In_2555);
xnor U1078 (N_1078,In_3184,In_2587);
and U1079 (N_1079,In_2750,In_1997);
xor U1080 (N_1080,In_507,In_570);
nor U1081 (N_1081,In_2592,In_4593);
nand U1082 (N_1082,In_140,In_4035);
or U1083 (N_1083,In_4801,In_300);
and U1084 (N_1084,In_4830,In_4515);
nor U1085 (N_1085,In_1098,In_2474);
nor U1086 (N_1086,In_1502,In_1980);
nor U1087 (N_1087,In_2062,In_4263);
or U1088 (N_1088,In_671,In_3932);
nand U1089 (N_1089,In_935,In_102);
or U1090 (N_1090,In_2954,In_3558);
xor U1091 (N_1091,In_3873,In_2810);
nand U1092 (N_1092,In_2858,In_1092);
or U1093 (N_1093,In_2873,In_704);
nor U1094 (N_1094,In_741,In_4352);
nor U1095 (N_1095,In_3457,In_1479);
nand U1096 (N_1096,In_2120,In_3492);
and U1097 (N_1097,In_4766,In_2976);
and U1098 (N_1098,In_3223,In_2848);
nor U1099 (N_1099,In_710,In_3008);
or U1100 (N_1100,In_3533,In_4118);
xnor U1101 (N_1101,In_4982,In_279);
nor U1102 (N_1102,In_1079,In_1624);
nor U1103 (N_1103,In_49,In_2602);
nor U1104 (N_1104,In_2259,In_4547);
or U1105 (N_1105,In_3119,In_280);
or U1106 (N_1106,In_2729,In_971);
or U1107 (N_1107,In_204,In_4756);
and U1108 (N_1108,In_4870,In_3548);
nand U1109 (N_1109,In_641,In_4391);
xnor U1110 (N_1110,In_2913,In_3928);
nand U1111 (N_1111,In_4936,In_1182);
or U1112 (N_1112,In_2039,In_1774);
nor U1113 (N_1113,In_2225,In_2969);
xor U1114 (N_1114,In_4791,In_2631);
or U1115 (N_1115,In_2063,In_1946);
or U1116 (N_1116,In_1159,In_1286);
and U1117 (N_1117,In_1558,In_3992);
or U1118 (N_1118,In_4798,In_2435);
xnor U1119 (N_1119,In_3618,In_4211);
xor U1120 (N_1120,In_2028,In_4149);
nor U1121 (N_1121,In_3106,In_1892);
and U1122 (N_1122,In_21,In_239);
nor U1123 (N_1123,In_3675,In_1264);
nand U1124 (N_1124,In_2108,In_1042);
nor U1125 (N_1125,In_3803,In_3895);
and U1126 (N_1126,In_3987,In_1406);
or U1127 (N_1127,In_3625,In_411);
and U1128 (N_1128,In_24,In_193);
nand U1129 (N_1129,In_6,In_4332);
nor U1130 (N_1130,In_4025,In_4620);
nand U1131 (N_1131,In_1373,In_3791);
xor U1132 (N_1132,In_2042,In_1728);
or U1133 (N_1133,In_3927,In_2897);
or U1134 (N_1134,In_109,In_875);
or U1135 (N_1135,In_2857,In_110);
nand U1136 (N_1136,In_3446,In_85);
xnor U1137 (N_1137,In_466,In_2324);
nor U1138 (N_1138,In_3624,In_30);
or U1139 (N_1139,In_1653,In_2776);
or U1140 (N_1140,In_4772,In_3354);
nor U1141 (N_1141,In_4716,In_981);
and U1142 (N_1142,In_3760,In_1485);
or U1143 (N_1143,In_2681,In_2861);
or U1144 (N_1144,In_2514,In_1080);
nand U1145 (N_1145,In_634,In_508);
nor U1146 (N_1146,In_1803,In_3643);
xor U1147 (N_1147,In_530,In_514);
and U1148 (N_1148,In_4328,In_4685);
nor U1149 (N_1149,In_3860,In_91);
nor U1150 (N_1150,In_811,In_1253);
nand U1151 (N_1151,In_1227,In_147);
or U1152 (N_1152,In_2043,In_104);
and U1153 (N_1153,In_622,In_2264);
nand U1154 (N_1154,In_3137,In_3691);
or U1155 (N_1155,In_2172,In_1822);
nand U1156 (N_1156,In_484,In_3696);
or U1157 (N_1157,In_4082,In_2193);
and U1158 (N_1158,In_4094,In_4295);
nor U1159 (N_1159,In_1560,In_680);
and U1160 (N_1160,In_3114,In_3816);
or U1161 (N_1161,In_2814,In_2396);
nand U1162 (N_1162,In_3699,In_921);
xor U1163 (N_1163,In_1401,In_4984);
and U1164 (N_1164,In_2787,In_4458);
nor U1165 (N_1165,In_4495,In_1157);
xnor U1166 (N_1166,In_2208,In_2347);
nand U1167 (N_1167,In_2444,In_1843);
or U1168 (N_1168,In_4509,In_2887);
nor U1169 (N_1169,In_2095,In_4632);
xor U1170 (N_1170,In_1701,In_3306);
nand U1171 (N_1171,In_4607,In_3335);
xnor U1172 (N_1172,In_1369,In_2488);
and U1173 (N_1173,In_4418,In_4005);
and U1174 (N_1174,In_1949,In_1100);
xor U1175 (N_1175,In_1385,In_1981);
nand U1176 (N_1176,In_3097,In_758);
nor U1177 (N_1177,In_3033,In_4154);
xor U1178 (N_1178,In_263,In_742);
nand U1179 (N_1179,In_1923,In_714);
and U1180 (N_1180,In_3470,In_536);
xnor U1181 (N_1181,In_3322,In_4916);
and U1182 (N_1182,In_1680,In_2319);
or U1183 (N_1183,In_302,In_2220);
nor U1184 (N_1184,In_3066,In_1325);
and U1185 (N_1185,In_2888,In_2195);
xnor U1186 (N_1186,In_1005,In_136);
xor U1187 (N_1187,In_3779,In_829);
xnor U1188 (N_1188,In_2950,In_719);
nand U1189 (N_1189,In_28,In_186);
xnor U1190 (N_1190,In_574,In_1330);
nand U1191 (N_1191,In_3108,In_1669);
xnor U1192 (N_1192,In_2090,In_4128);
or U1193 (N_1193,In_1517,In_2628);
and U1194 (N_1194,In_4100,In_4615);
nand U1195 (N_1195,In_3500,In_3201);
xnor U1196 (N_1196,In_806,In_83);
nand U1197 (N_1197,In_1862,In_1823);
and U1198 (N_1198,In_235,In_3010);
xor U1199 (N_1199,In_4642,In_4198);
nor U1200 (N_1200,In_2653,In_2801);
xor U1201 (N_1201,In_4067,In_1612);
or U1202 (N_1202,In_1679,In_898);
or U1203 (N_1203,In_3978,In_814);
nor U1204 (N_1204,In_4130,In_2503);
xor U1205 (N_1205,In_1677,In_1746);
and U1206 (N_1206,In_3053,In_4660);
nand U1207 (N_1207,In_1960,In_1634);
and U1208 (N_1208,In_3610,In_1142);
nor U1209 (N_1209,In_3129,In_2622);
xor U1210 (N_1210,In_444,In_908);
nand U1211 (N_1211,In_1779,In_112);
and U1212 (N_1212,In_1340,In_4662);
xor U1213 (N_1213,In_541,In_2855);
nor U1214 (N_1214,In_134,In_3267);
and U1215 (N_1215,In_2999,In_1617);
nand U1216 (N_1216,In_4427,In_1009);
or U1217 (N_1217,In_4617,In_2800);
xnor U1218 (N_1218,In_4103,In_4634);
and U1219 (N_1219,In_4075,In_2978);
xnor U1220 (N_1220,In_1999,In_722);
xnor U1221 (N_1221,In_1154,In_874);
and U1222 (N_1222,In_18,In_4639);
xor U1223 (N_1223,In_3117,In_2789);
or U1224 (N_1224,In_1223,In_4394);
xnor U1225 (N_1225,In_987,In_954);
or U1226 (N_1226,In_3218,In_538);
and U1227 (N_1227,In_3327,In_4440);
nand U1228 (N_1228,In_2152,In_3189);
nand U1229 (N_1229,In_3178,In_1292);
or U1230 (N_1230,In_2251,In_335);
and U1231 (N_1231,In_2666,In_692);
and U1232 (N_1232,In_4463,In_2130);
nor U1233 (N_1233,In_3146,In_1283);
xnor U1234 (N_1234,In_431,In_1777);
nor U1235 (N_1235,In_1248,In_22);
nand U1236 (N_1236,In_3754,In_4800);
xnor U1237 (N_1237,In_3142,In_2576);
or U1238 (N_1238,In_3337,In_3706);
nand U1239 (N_1239,In_2517,In_826);
nor U1240 (N_1240,In_3029,In_1022);
and U1241 (N_1241,In_1842,In_842);
or U1242 (N_1242,In_2275,In_4886);
nand U1243 (N_1243,In_4834,In_1587);
xor U1244 (N_1244,In_4806,In_4438);
or U1245 (N_1245,In_1318,In_1130);
nor U1246 (N_1246,In_2127,In_789);
xnor U1247 (N_1247,In_866,In_947);
xor U1248 (N_1248,In_3447,In_1911);
or U1249 (N_1249,In_4774,In_3687);
and U1250 (N_1250,In_1819,In_3716);
and U1251 (N_1251,In_4972,In_4933);
nor U1252 (N_1252,In_1277,In_2696);
and U1253 (N_1253,In_3914,In_1905);
xor U1254 (N_1254,In_1963,In_546);
nor U1255 (N_1255,In_3637,In_534);
nand U1256 (N_1256,In_582,In_4490);
nor U1257 (N_1257,In_2921,In_4445);
xnor U1258 (N_1258,In_2031,In_2363);
xor U1259 (N_1259,In_2086,In_1218);
nand U1260 (N_1260,In_301,In_4803);
nor U1261 (N_1261,In_4145,In_712);
and U1262 (N_1262,In_848,In_3959);
and U1263 (N_1263,In_3742,In_2408);
nand U1264 (N_1264,In_2218,In_4156);
or U1265 (N_1265,In_4887,In_4471);
nor U1266 (N_1266,In_4253,In_4582);
nand U1267 (N_1267,In_2184,In_2384);
nor U1268 (N_1268,In_1984,In_3929);
nor U1269 (N_1269,In_47,In_3039);
and U1270 (N_1270,In_1778,In_563);
or U1271 (N_1271,In_3830,In_1870);
and U1272 (N_1272,In_851,In_3604);
nor U1273 (N_1273,In_1213,In_2850);
xnor U1274 (N_1274,In_12,In_3596);
nand U1275 (N_1275,In_90,In_2912);
nand U1276 (N_1276,In_4245,In_1238);
nor U1277 (N_1277,In_1812,In_3651);
nand U1278 (N_1278,In_207,In_2181);
xnor U1279 (N_1279,In_3998,In_2968);
nand U1280 (N_1280,In_3617,In_833);
xor U1281 (N_1281,In_3875,In_1478);
nor U1282 (N_1282,In_2898,In_3312);
nand U1283 (N_1283,In_1555,In_3384);
nand U1284 (N_1284,In_3081,In_4724);
xnor U1285 (N_1285,In_4286,In_505);
xor U1286 (N_1286,In_3752,In_4506);
nand U1287 (N_1287,In_2608,In_2389);
xnor U1288 (N_1288,In_379,In_2686);
nand U1289 (N_1289,In_4206,In_1462);
or U1290 (N_1290,In_3746,In_3040);
nand U1291 (N_1291,In_4601,In_4812);
and U1292 (N_1292,In_4208,In_3529);
and U1293 (N_1293,In_1003,In_616);
and U1294 (N_1294,In_4170,In_4918);
and U1295 (N_1295,In_358,In_284);
nor U1296 (N_1296,In_4460,In_1065);
nor U1297 (N_1297,In_1273,In_4026);
nor U1298 (N_1298,In_1668,In_487);
and U1299 (N_1299,In_4350,In_3059);
xor U1300 (N_1300,In_4079,In_1348);
xor U1301 (N_1301,In_4948,In_4371);
or U1302 (N_1302,In_4820,In_3950);
nor U1303 (N_1303,In_4708,In_2860);
xnor U1304 (N_1304,In_1908,In_2524);
and U1305 (N_1305,In_1052,In_645);
or U1306 (N_1306,In_395,In_4744);
or U1307 (N_1307,In_2925,In_247);
xor U1308 (N_1308,In_4376,In_4030);
xnor U1309 (N_1309,In_986,In_3923);
xor U1310 (N_1310,In_2452,In_511);
xnor U1311 (N_1311,In_3664,In_1314);
and U1312 (N_1312,In_4197,In_1894);
xnor U1313 (N_1313,In_4963,In_2773);
and U1314 (N_1314,In_4536,In_1893);
xnor U1315 (N_1315,In_2067,In_590);
and U1316 (N_1316,In_1331,In_208);
or U1317 (N_1317,In_3478,In_4099);
or U1318 (N_1318,In_2310,In_84);
nand U1319 (N_1319,In_4055,In_3474);
nand U1320 (N_1320,In_2284,In_174);
or U1321 (N_1321,In_639,In_288);
and U1322 (N_1322,In_1017,In_1881);
xnor U1323 (N_1323,In_3247,In_1486);
nand U1324 (N_1324,In_3222,In_3320);
xnor U1325 (N_1325,In_1141,In_4160);
nor U1326 (N_1326,In_3052,In_4216);
or U1327 (N_1327,In_1697,In_4940);
xnor U1328 (N_1328,In_2992,In_3648);
nand U1329 (N_1329,In_3328,In_1958);
nand U1330 (N_1330,In_1294,In_48);
or U1331 (N_1331,In_4912,In_515);
nand U1332 (N_1332,In_277,In_4325);
nor U1333 (N_1333,In_2214,In_4493);
xnor U1334 (N_1334,In_4001,In_3622);
and U1335 (N_1335,In_1790,In_3593);
and U1336 (N_1336,In_4504,In_597);
nor U1337 (N_1337,In_4192,In_451);
nor U1338 (N_1338,In_446,In_2636);
nand U1339 (N_1339,In_2895,In_3636);
and U1340 (N_1340,In_3386,In_2844);
and U1341 (N_1341,In_4023,In_1063);
or U1342 (N_1342,In_2457,In_2591);
or U1343 (N_1343,In_4016,In_2312);
and U1344 (N_1344,In_4903,In_1858);
or U1345 (N_1345,In_496,In_3750);
nand U1346 (N_1346,In_4597,In_2945);
nor U1347 (N_1347,In_191,In_1914);
nand U1348 (N_1348,In_205,In_956);
and U1349 (N_1349,In_493,In_915);
and U1350 (N_1350,In_4069,In_3656);
nor U1351 (N_1351,In_3245,In_2000);
and U1352 (N_1352,In_4950,In_618);
nand U1353 (N_1353,In_1364,In_4989);
nand U1354 (N_1354,In_3718,In_478);
and U1355 (N_1355,In_1336,In_2432);
xor U1356 (N_1356,In_4098,In_2147);
and U1357 (N_1357,In_3211,In_2463);
or U1358 (N_1358,In_1667,In_1535);
xnor U1359 (N_1359,In_2048,In_779);
nand U1360 (N_1360,In_1116,In_2204);
or U1361 (N_1361,In_2546,In_3098);
nor U1362 (N_1362,In_653,In_924);
nand U1363 (N_1363,In_2783,In_1621);
or U1364 (N_1364,In_3011,In_1133);
nor U1365 (N_1365,In_3655,In_3290);
xnor U1366 (N_1366,In_2458,In_246);
or U1367 (N_1367,In_1750,In_4472);
xnor U1368 (N_1368,In_2325,In_2427);
nor U1369 (N_1369,In_409,In_2065);
and U1370 (N_1370,In_3424,In_1239);
nand U1371 (N_1371,In_4077,In_3263);
and U1372 (N_1372,In_1757,In_1856);
and U1373 (N_1373,In_3163,In_2712);
xnor U1374 (N_1374,In_2009,In_1205);
and U1375 (N_1375,In_849,In_3228);
or U1376 (N_1376,In_2418,In_1922);
nand U1377 (N_1377,In_1272,In_467);
nor U1378 (N_1378,In_3208,In_4752);
xnor U1379 (N_1379,In_2126,In_1770);
and U1380 (N_1380,In_750,In_4123);
or U1381 (N_1381,In_1796,In_912);
or U1382 (N_1382,In_1240,In_4503);
nor U1383 (N_1383,In_4409,In_3202);
and U1384 (N_1384,In_2752,In_2768);
and U1385 (N_1385,In_984,In_1863);
and U1386 (N_1386,In_1360,In_2180);
xor U1387 (N_1387,In_1428,In_4604);
xor U1388 (N_1388,In_2326,In_334);
nand U1389 (N_1389,In_4652,In_2623);
and U1390 (N_1390,In_580,In_717);
and U1391 (N_1391,In_116,In_2856);
xnor U1392 (N_1392,In_4904,In_2825);
and U1393 (N_1393,In_2242,In_527);
and U1394 (N_1394,In_4924,In_4266);
and U1395 (N_1395,In_3773,In_4355);
xor U1396 (N_1396,In_2340,In_3469);
xor U1397 (N_1397,In_4450,In_4424);
nor U1398 (N_1398,In_4033,In_4725);
xor U1399 (N_1399,In_1696,In_159);
nor U1400 (N_1400,In_4958,In_1708);
xnor U1401 (N_1401,In_3162,In_1038);
xnor U1402 (N_1402,In_976,In_2104);
xnor U1403 (N_1403,In_328,In_815);
xnor U1404 (N_1404,In_787,In_4565);
or U1405 (N_1405,In_1275,In_4240);
and U1406 (N_1406,In_173,In_2984);
or U1407 (N_1407,In_3867,In_1467);
nor U1408 (N_1408,In_676,In_3785);
xnor U1409 (N_1409,In_455,In_3729);
and U1410 (N_1410,In_1129,In_884);
nand U1411 (N_1411,In_1128,In_4704);
xnor U1412 (N_1412,In_2023,In_3280);
nor U1413 (N_1413,In_3315,In_1755);
or U1414 (N_1414,In_3986,In_3859);
nand U1415 (N_1415,In_767,In_3781);
nand U1416 (N_1416,In_792,In_853);
and U1417 (N_1417,In_4876,In_3168);
nor U1418 (N_1418,In_1106,In_3713);
nand U1419 (N_1419,In_1443,In_33);
nand U1420 (N_1420,In_3903,In_1058);
nand U1421 (N_1421,In_3279,In_804);
xor U1422 (N_1422,In_2226,In_3112);
xor U1423 (N_1423,In_2926,In_3213);
and U1424 (N_1424,In_929,In_307);
and U1425 (N_1425,In_1924,In_410);
or U1426 (N_1426,In_3351,In_4292);
or U1427 (N_1427,In_3893,In_4926);
or U1428 (N_1428,In_388,In_384);
and U1429 (N_1429,In_3824,In_2543);
nand U1430 (N_1430,In_2261,In_3324);
nand U1431 (N_1431,In_739,In_4161);
xor U1432 (N_1432,In_2986,In_2016);
or U1433 (N_1433,In_3829,In_3935);
nand U1434 (N_1434,In_776,In_2333);
nand U1435 (N_1435,In_1024,In_86);
xnor U1436 (N_1436,In_2909,In_3375);
nor U1437 (N_1437,In_2380,In_2229);
or U1438 (N_1438,In_820,In_818);
or U1439 (N_1439,In_1470,In_4554);
nor U1440 (N_1440,In_293,In_4071);
nand U1441 (N_1441,In_4188,In_2269);
or U1442 (N_1442,In_2967,In_1590);
nor U1443 (N_1443,In_2703,In_1288);
and U1444 (N_1444,In_2368,In_1936);
or U1445 (N_1445,In_4134,In_449);
nand U1446 (N_1446,In_441,In_2663);
or U1447 (N_1447,In_890,In_2962);
and U1448 (N_1448,In_2146,In_3646);
xnor U1449 (N_1449,In_400,In_693);
nand U1450 (N_1450,In_4117,In_2412);
xor U1451 (N_1451,In_3186,In_1973);
nand U1452 (N_1452,In_2541,In_2079);
and U1453 (N_1453,In_3579,In_2076);
nor U1454 (N_1454,In_3362,In_3122);
and U1455 (N_1455,In_4951,In_486);
xor U1456 (N_1456,In_1312,In_3396);
and U1457 (N_1457,In_1760,In_632);
and U1458 (N_1458,In_4562,In_2578);
nand U1459 (N_1459,In_4900,In_135);
xnor U1460 (N_1460,In_3342,In_3761);
nand U1461 (N_1461,In_4733,In_41);
xnor U1462 (N_1462,In_4529,In_434);
xor U1463 (N_1463,In_23,In_4782);
or U1464 (N_1464,In_3711,In_1477);
xnor U1465 (N_1465,In_3192,In_266);
nor U1466 (N_1466,In_3325,In_4769);
nor U1467 (N_1467,In_2471,In_2813);
or U1468 (N_1468,In_3666,In_566);
nor U1469 (N_1469,In_3901,In_2809);
nor U1470 (N_1470,In_3068,In_2554);
nor U1471 (N_1471,In_3361,In_3188);
nand U1472 (N_1472,In_1990,In_3444);
nor U1473 (N_1473,In_1408,In_4750);
xnor U1474 (N_1474,In_1644,In_1115);
nand U1475 (N_1475,In_2778,In_753);
nand U1476 (N_1476,In_3429,In_952);
xor U1477 (N_1477,In_1102,In_781);
xnor U1478 (N_1478,In_1569,In_2977);
xor U1479 (N_1479,In_1737,In_1256);
nand U1480 (N_1480,In_1512,In_3676);
and U1481 (N_1481,In_2231,In_1393);
nand U1482 (N_1482,In_2721,In_1384);
xor U1483 (N_1483,In_316,In_4653);
and U1484 (N_1484,In_2144,In_1943);
nor U1485 (N_1485,In_1895,In_2239);
or U1486 (N_1486,In_2480,In_2433);
or U1487 (N_1487,In_3707,In_3260);
xnor U1488 (N_1488,In_2695,In_2390);
xnor U1489 (N_1489,In_4600,In_2382);
nor U1490 (N_1490,In_4239,In_1306);
nand U1491 (N_1491,In_4457,In_2223);
or U1492 (N_1492,In_1841,In_711);
or U1493 (N_1493,In_3550,In_4142);
or U1494 (N_1494,In_139,In_2257);
nor U1495 (N_1495,In_3344,In_881);
or U1496 (N_1496,In_3438,In_3968);
nand U1497 (N_1497,In_4633,In_461);
nand U1498 (N_1498,In_2361,In_1639);
and U1499 (N_1499,In_4400,In_4866);
and U1500 (N_1500,In_223,In_4401);
or U1501 (N_1501,In_2036,In_3581);
nor U1502 (N_1502,In_423,In_408);
xor U1503 (N_1503,In_3078,In_1882);
and U1504 (N_1504,In_2116,In_2327);
and U1505 (N_1505,In_175,In_2182);
nor U1506 (N_1506,In_1764,In_3811);
xor U1507 (N_1507,In_2318,In_3128);
nor U1508 (N_1508,In_3908,In_382);
xor U1509 (N_1509,In_1507,In_4668);
xor U1510 (N_1510,In_1171,In_321);
xor U1511 (N_1511,In_2320,In_3513);
and U1512 (N_1512,In_2388,In_4563);
or U1513 (N_1513,In_2020,In_1531);
or U1514 (N_1514,In_2936,In_1425);
xnor U1515 (N_1515,In_2351,In_2112);
or U1516 (N_1516,In_1853,In_2660);
or U1517 (N_1517,In_4771,In_161);
nor U1518 (N_1518,In_4873,In_268);
or U1519 (N_1519,In_1493,In_2004);
or U1520 (N_1520,In_1628,In_391);
nand U1521 (N_1521,In_3930,In_2271);
xor U1522 (N_1522,In_4692,In_4399);
xor U1523 (N_1523,In_4952,In_4953);
or U1524 (N_1524,In_1422,In_2187);
and U1525 (N_1525,In_4274,In_3015);
nor U1526 (N_1526,In_1327,In_775);
or U1527 (N_1527,In_2837,In_743);
nand U1528 (N_1528,In_3454,In_4335);
and U1529 (N_1529,In_4909,In_3912);
and U1530 (N_1530,In_3012,In_3364);
nand U1531 (N_1531,In_3473,In_3759);
nand U1532 (N_1532,In_3358,In_4754);
nor U1533 (N_1533,In_3590,In_3164);
xnor U1534 (N_1534,In_2886,In_445);
and U1535 (N_1535,In_1975,In_1538);
nor U1536 (N_1536,In_322,In_807);
xnor U1537 (N_1537,In_2166,In_385);
or U1538 (N_1538,In_2069,In_2638);
nor U1539 (N_1539,In_4076,In_4466);
nor U1540 (N_1540,In_4494,In_2822);
and U1541 (N_1541,In_2745,In_2872);
nor U1542 (N_1542,In_2305,In_4431);
or U1543 (N_1543,In_4603,In_1505);
nand U1544 (N_1544,In_2426,In_383);
xor U1545 (N_1545,In_1591,In_3464);
nand U1546 (N_1546,In_1184,In_723);
nor U1547 (N_1547,In_4435,In_1456);
nand U1548 (N_1548,In_3700,In_3827);
or U1549 (N_1549,In_2,In_2700);
and U1550 (N_1550,In_4256,In_1891);
nand U1551 (N_1551,In_4993,In_880);
xnor U1552 (N_1552,In_4610,In_2068);
xnor U1553 (N_1553,In_2386,In_816);
nor U1554 (N_1554,In_2845,In_2217);
nand U1555 (N_1555,In_3611,In_728);
nand U1556 (N_1556,In_4209,In_1356);
nor U1557 (N_1557,In_2621,In_1759);
nor U1558 (N_1558,In_2153,In_4990);
or U1559 (N_1559,In_3983,In_1626);
xor U1560 (N_1560,In_604,In_4248);
nor U1561 (N_1561,In_2908,In_1332);
xnor U1562 (N_1562,In_2082,In_4751);
or U1563 (N_1563,In_4317,In_3528);
and U1564 (N_1564,In_1964,In_1043);
xor U1565 (N_1565,In_1391,In_1027);
and U1566 (N_1566,In_4720,In_3079);
nor U1567 (N_1567,In_4370,In_1909);
or U1568 (N_1568,In_796,In_2364);
or U1569 (N_1569,In_2994,In_1197);
nand U1570 (N_1570,In_4127,In_2866);
nand U1571 (N_1571,In_2473,In_3058);
and U1572 (N_1572,In_118,In_945);
and U1573 (N_1573,In_1663,In_2131);
and U1574 (N_1574,In_4315,In_2788);
and U1575 (N_1575,In_3660,In_644);
nor U1576 (N_1576,In_2487,In_3024);
nand U1577 (N_1577,In_1196,In_2889);
or U1578 (N_1578,In_1156,In_3813);
nand U1579 (N_1579,In_4822,In_917);
or U1580 (N_1580,In_4383,In_3823);
nand U1581 (N_1581,In_2833,In_353);
nor U1582 (N_1582,In_4705,In_1772);
nand U1583 (N_1583,In_3915,In_4363);
or U1584 (N_1584,In_1544,In_1576);
nor U1585 (N_1585,In_4168,In_1454);
nand U1586 (N_1586,In_1281,In_3258);
and U1587 (N_1587,In_3767,In_4784);
or U1588 (N_1588,In_3441,In_1039);
xor U1589 (N_1589,In_4318,In_3567);
nor U1590 (N_1590,In_2959,In_4300);
nor U1591 (N_1591,In_1487,In_1296);
or U1592 (N_1592,In_2914,In_685);
and U1593 (N_1593,In_179,In_1287);
nor U1594 (N_1594,In_2867,In_531);
or U1595 (N_1595,In_4999,In_1319);
nand U1596 (N_1596,In_3967,In_3542);
and U1597 (N_1597,In_1126,In_117);
xnor U1598 (N_1598,In_621,In_3887);
nand U1599 (N_1599,In_772,In_4061);
or U1600 (N_1600,In_603,In_2582);
xnor U1601 (N_1601,In_492,In_4480);
xor U1602 (N_1602,In_567,In_1433);
nor U1603 (N_1603,In_1075,In_1480);
nand U1604 (N_1604,In_3728,In_338);
or U1605 (N_1605,In_4998,In_4631);
xor U1606 (N_1606,In_4191,In_273);
nor U1607 (N_1607,In_2094,In_4590);
or U1608 (N_1608,In_2792,In_4743);
and U1609 (N_1609,In_3856,In_4135);
nor U1610 (N_1610,In_1886,In_3777);
and U1611 (N_1611,In_2864,In_2234);
and U1612 (N_1612,In_164,In_3450);
nor U1613 (N_1613,In_4038,In_3252);
xnor U1614 (N_1614,In_4836,In_4928);
and U1615 (N_1615,In_782,In_4987);
or U1616 (N_1616,In_4808,In_4122);
xor U1617 (N_1617,In_2970,In_4695);
and U1618 (N_1618,In_1434,In_4476);
nor U1619 (N_1619,In_1463,In_231);
and U1620 (N_1620,In_4224,In_4965);
or U1621 (N_1621,In_2398,In_3702);
nor U1622 (N_1622,In_2462,In_259);
nor U1623 (N_1623,In_4988,In_4932);
or U1624 (N_1624,In_1420,In_2033);
nand U1625 (N_1625,In_3916,In_1285);
nand U1626 (N_1626,In_2176,In_426);
xnor U1627 (N_1627,In_176,In_1969);
or U1628 (N_1628,In_3269,In_4313);
nor U1629 (N_1629,In_1168,In_1672);
nor U1630 (N_1630,In_4164,In_2756);
or U1631 (N_1631,In_4287,In_1702);
or U1632 (N_1632,In_4181,In_725);
nand U1633 (N_1633,In_3461,In_4228);
or U1634 (N_1634,In_1235,In_3863);
xnor U1635 (N_1635,In_1324,In_1523);
nor U1636 (N_1636,In_2894,In_788);
xor U1637 (N_1637,In_2707,In_4374);
nor U1638 (N_1638,In_4146,In_4545);
and U1639 (N_1639,In_3418,In_757);
xor U1640 (N_1640,In_1592,In_2899);
nand U1641 (N_1641,In_4112,In_2037);
and U1642 (N_1642,In_3539,In_457);
xnor U1643 (N_1643,In_1852,In_1460);
nand U1644 (N_1644,In_1756,In_1791);
or U1645 (N_1645,In_3153,In_415);
xnor U1646 (N_1646,In_1817,In_3657);
or U1647 (N_1647,In_948,In_1585);
nand U1648 (N_1648,In_4367,In_367);
nand U1649 (N_1649,In_989,In_3599);
xor U1650 (N_1650,In_2295,In_791);
nand U1651 (N_1651,In_3969,In_3838);
or U1652 (N_1652,In_2245,In_4824);
and U1653 (N_1653,In_4907,In_1832);
or U1654 (N_1654,In_2952,In_2314);
nor U1655 (N_1655,In_344,In_3329);
nand U1656 (N_1656,In_1741,In_3027);
xnor U1657 (N_1657,In_4144,In_819);
and U1658 (N_1658,In_4852,In_4944);
and U1659 (N_1659,In_442,In_3747);
xor U1660 (N_1660,In_1469,In_4289);
nor U1661 (N_1661,In_3819,In_763);
xor U1662 (N_1662,In_4622,In_1282);
or U1663 (N_1663,In_4511,In_2757);
nand U1664 (N_1664,In_4218,In_926);
xor U1665 (N_1665,In_2280,In_1801);
nor U1666 (N_1666,In_2658,In_3370);
nand U1667 (N_1667,In_2834,In_80);
or U1668 (N_1668,In_3546,In_1710);
and U1669 (N_1669,In_3366,In_737);
nand U1670 (N_1670,In_4379,In_240);
nor U1671 (N_1671,In_1276,In_2077);
nor U1672 (N_1672,In_3917,In_2409);
xor U1673 (N_1673,In_3439,In_4421);
and U1674 (N_1674,In_2985,In_4223);
or U1675 (N_1675,In_3401,In_3042);
nand U1676 (N_1676,In_1520,In_4748);
nor U1677 (N_1677,In_4840,In_2404);
nor U1678 (N_1678,In_1602,In_4688);
nand U1679 (N_1679,In_1353,In_4524);
nor U1680 (N_1680,In_4732,In_4157);
and U1681 (N_1681,In_1225,In_4406);
nor U1682 (N_1682,In_1028,In_2567);
xor U1683 (N_1683,In_4624,In_3144);
xnor U1684 (N_1684,In_3523,In_1007);
and U1685 (N_1685,In_860,In_4669);
xnor U1686 (N_1686,In_4689,In_2334);
or U1687 (N_1687,In_4002,In_4525);
nor U1688 (N_1688,In_2852,In_3077);
nor U1689 (N_1689,In_2997,In_524);
and U1690 (N_1690,In_4534,In_4416);
and U1691 (N_1691,In_1269,In_3277);
nor U1692 (N_1692,In_1259,In_3591);
xnor U1693 (N_1693,In_4425,In_752);
or U1694 (N_1694,In_3465,In_4303);
or U1695 (N_1695,In_4676,In_3594);
xor U1696 (N_1696,In_3103,In_3572);
xnor U1697 (N_1697,In_951,In_267);
and U1698 (N_1698,In_4723,In_2862);
or U1699 (N_1699,In_2772,In_3769);
nor U1700 (N_1700,In_3620,In_3560);
and U1701 (N_1701,In_2183,In_1761);
xor U1702 (N_1702,In_160,In_1994);
or U1703 (N_1703,In_2748,In_4381);
or U1704 (N_1704,In_3698,In_4074);
or U1705 (N_1705,In_2134,In_4573);
or U1706 (N_1706,In_4550,In_456);
and U1707 (N_1707,In_1605,In_3355);
or U1708 (N_1708,In_3629,In_3902);
or U1709 (N_1709,In_2829,In_260);
nor U1710 (N_1710,In_1835,In_4583);
xor U1711 (N_1711,In_99,In_2998);
and U1712 (N_1712,In_3031,In_845);
nor U1713 (N_1713,In_4776,In_3790);
and U1714 (N_1714,In_399,In_4024);
and U1715 (N_1715,In_966,In_2868);
and U1716 (N_1716,In_702,In_3270);
and U1717 (N_1717,In_861,In_2836);
and U1718 (N_1718,In_100,In_901);
xnor U1719 (N_1719,In_679,In_777);
nor U1720 (N_1720,In_4108,In_3658);
xnor U1721 (N_1721,In_2842,In_290);
nor U1722 (N_1722,In_1681,In_1094);
nor U1723 (N_1723,In_3095,In_4346);
or U1724 (N_1724,In_4322,In_1415);
or U1725 (N_1725,In_1107,In_2290);
nand U1726 (N_1726,In_2802,In_2199);
xnor U1727 (N_1727,In_4742,In_4137);
nand U1728 (N_1728,In_2406,In_1194);
and U1729 (N_1729,In_35,In_4284);
and U1730 (N_1730,In_1526,In_3532);
nor U1731 (N_1731,In_2882,In_1556);
nor U1732 (N_1732,In_2863,In_2478);
or U1733 (N_1733,In_3017,In_2758);
nand U1734 (N_1734,In_4512,In_1230);
xnor U1735 (N_1735,In_856,In_3710);
or U1736 (N_1736,In_2008,In_3239);
nor U1737 (N_1737,In_1333,In_4895);
or U1738 (N_1738,In_2618,In_3695);
nor U1739 (N_1739,In_1993,In_3996);
nor U1740 (N_1740,In_2267,In_1828);
nand U1741 (N_1741,In_930,In_3323);
or U1742 (N_1742,In_3979,In_605);
and U1743 (N_1743,In_4856,In_356);
nand U1744 (N_1744,In_3065,In_999);
or U1745 (N_1745,In_2539,In_1867);
and U1746 (N_1746,In_4250,In_3353);
nand U1747 (N_1747,In_2780,In_4283);
or U1748 (N_1748,In_992,In_2338);
nor U1749 (N_1749,In_3190,In_4032);
nand U1750 (N_1750,In_3299,In_183);
and U1751 (N_1751,In_2938,In_1956);
and U1752 (N_1752,In_27,In_4551);
nor U1753 (N_1753,In_3948,In_4403);
nand U1754 (N_1754,In_963,In_2198);
or U1755 (N_1755,In_1090,In_474);
xnor U1756 (N_1756,In_3974,In_242);
or U1757 (N_1757,In_667,In_3515);
nand U1758 (N_1758,In_3460,In_1752);
and U1759 (N_1759,In_2270,In_4185);
or U1760 (N_1760,In_1183,In_681);
xor U1761 (N_1761,In_3412,In_2819);
or U1762 (N_1762,In_4207,In_2730);
xnor U1763 (N_1763,In_3640,In_606);
nor U1764 (N_1764,In_4606,In_1048);
xnor U1765 (N_1765,In_1573,In_3776);
and U1766 (N_1766,In_1374,In_3962);
nor U1767 (N_1767,In_4703,In_11);
nor U1768 (N_1768,In_2081,In_4764);
and U1769 (N_1769,In_3199,In_150);
nor U1770 (N_1770,In_1358,In_2728);
or U1771 (N_1771,In_4382,In_3032);
nand U1772 (N_1772,In_299,In_2006);
xnor U1773 (N_1773,In_1173,In_2963);
nand U1774 (N_1774,In_1382,In_4464);
nand U1775 (N_1775,In_1683,In_2830);
or U1776 (N_1776,In_2610,In_1056);
and U1777 (N_1777,In_1597,In_3007);
xnor U1778 (N_1778,In_403,In_4981);
xnor U1779 (N_1779,In_4162,In_2691);
and U1780 (N_1780,In_4066,In_3888);
nand U1781 (N_1781,In_4558,In_2460);
xor U1782 (N_1782,In_2096,In_3964);
nand U1783 (N_1783,In_1412,In_2699);
or U1784 (N_1784,In_3120,In_3292);
xnor U1785 (N_1785,In_88,In_4048);
nand U1786 (N_1786,In_378,In_4314);
or U1787 (N_1787,In_1766,In_4184);
nand U1788 (N_1788,In_3255,In_677);
nor U1789 (N_1789,In_3054,In_1559);
xor U1790 (N_1790,In_1599,In_1781);
xnor U1791 (N_1791,In_2383,In_2572);
nand U1792 (N_1792,In_3009,In_114);
or U1793 (N_1793,In_1201,In_2710);
and U1794 (N_1794,In_2215,In_4136);
and U1795 (N_1795,In_1903,In_157);
or U1796 (N_1796,In_2376,In_3797);
or U1797 (N_1797,In_2790,In_4681);
nand U1798 (N_1798,In_868,In_503);
nand U1799 (N_1799,In_1648,In_2706);
nand U1800 (N_1800,In_2980,In_2246);
nand U1801 (N_1801,In_3400,In_2381);
or U1802 (N_1802,In_2392,In_281);
nor U1803 (N_1803,In_4522,In_78);
or U1804 (N_1804,In_1046,In_144);
nand U1805 (N_1805,In_4031,In_4125);
nand U1806 (N_1806,In_2080,In_1339);
nor U1807 (N_1807,In_1270,In_3176);
xnor U1808 (N_1808,In_1424,In_1343);
or U1809 (N_1809,In_2483,In_3586);
or U1810 (N_1810,In_3937,In_3615);
xnor U1811 (N_1811,In_4658,In_153);
xnor U1812 (N_1812,In_4837,In_2167);
and U1813 (N_1813,In_2827,In_909);
xnor U1814 (N_1814,In_2781,In_764);
and U1815 (N_1815,In_1788,In_1089);
and U1816 (N_1816,In_4279,In_1280);
and U1817 (N_1817,In_3805,In_4595);
nor U1818 (N_1818,In_3276,In_3368);
or U1819 (N_1819,In_473,In_1010);
nand U1820 (N_1820,In_3828,In_3145);
or U1821 (N_1821,In_1481,In_1061);
nand U1822 (N_1822,In_262,In_1806);
nor U1823 (N_1823,In_4788,In_4780);
xor U1824 (N_1824,In_997,In_1342);
and U1825 (N_1825,In_4029,In_4785);
or U1826 (N_1826,In_1610,In_1915);
and U1827 (N_1827,In_1872,In_2015);
and U1828 (N_1828,In_2358,In_3947);
or U1829 (N_1829,In_1289,In_1160);
nor U1830 (N_1830,In_3764,In_2698);
nand U1831 (N_1831,In_1429,In_1871);
or U1832 (N_1832,In_331,In_2061);
nand U1833 (N_1833,In_13,In_361);
nand U1834 (N_1834,In_4324,In_4845);
nor U1835 (N_1835,In_697,In_4802);
or U1836 (N_1836,In_3517,In_2445);
xnor U1837 (N_1837,In_188,In_4546);
nand U1838 (N_1838,In_325,In_2791);
or U1839 (N_1839,In_2733,In_4119);
nand U1840 (N_1840,In_2366,In_2831);
and U1841 (N_1841,In_699,In_3016);
nand U1842 (N_1842,In_394,In_1338);
or U1843 (N_1843,In_3161,In_3076);
xor U1844 (N_1844,In_4111,In_4088);
and U1845 (N_1845,In_4867,In_978);
and U1846 (N_1846,In_2233,In_4411);
or U1847 (N_1847,In_4659,In_3422);
or U1848 (N_1848,In_3552,In_1013);
xnor U1849 (N_1849,In_2464,In_1918);
nand U1850 (N_1850,In_3141,In_1441);
and U1851 (N_1851,In_1178,In_450);
xnor U1852 (N_1852,In_1131,In_2701);
nand U1853 (N_1853,In_1543,In_1670);
nand U1854 (N_1854,In_2684,In_1987);
or U1855 (N_1855,In_3086,In_919);
xor U1856 (N_1856,In_3547,In_2260);
nand U1857 (N_1857,In_3704,In_2158);
and U1858 (N_1858,In_3224,In_2323);
nand U1859 (N_1859,In_219,In_2083);
nand U1860 (N_1860,In_4176,In_4229);
xor U1861 (N_1861,In_4619,In_4265);
nor U1862 (N_1862,In_3102,In_1411);
and U1863 (N_1863,In_1181,In_2034);
or U1864 (N_1864,In_1739,In_3338);
nand U1865 (N_1865,In_278,In_3519);
nand U1866 (N_1866,In_2577,In_1600);
nand U1867 (N_1867,In_3023,In_651);
and U1868 (N_1868,In_1198,In_2360);
nand U1869 (N_1869,In_3956,In_3371);
nand U1870 (N_1870,In_2041,In_2511);
nor U1871 (N_1871,In_3871,In_3621);
or U1872 (N_1872,In_665,In_2171);
and U1873 (N_1873,In_2720,In_3037);
nor U1874 (N_1874,In_337,In_1368);
xnor U1875 (N_1875,In_871,In_3022);
nor U1876 (N_1876,In_2504,In_3410);
or U1877 (N_1877,In_4227,In_3607);
xnor U1878 (N_1878,In_3043,In_4994);
nor U1879 (N_1879,In_347,In_4496);
and U1880 (N_1880,In_1367,In_4080);
nor U1881 (N_1881,In_1518,In_3619);
nor U1882 (N_1882,In_3241,In_1371);
nor U1883 (N_1883,In_1899,In_3677);
nand U1884 (N_1884,In_2674,In_162);
nand U1885 (N_1885,In_549,In_4358);
xor U1886 (N_1886,In_4428,In_3348);
nor U1887 (N_1887,In_2646,In_2714);
nand U1888 (N_1888,In_1268,In_2885);
nand U1889 (N_1889,In_4977,In_1557);
nor U1890 (N_1890,In_3703,In_2983);
and U1891 (N_1891,In_498,In_1400);
and U1892 (N_1892,In_1072,In_1510);
nand U1893 (N_1893,In_661,In_1187);
and U1894 (N_1894,In_1073,In_4602);
xnor U1895 (N_1895,In_2890,In_3278);
and U1896 (N_1896,In_3608,In_4212);
nand U1897 (N_1897,In_716,In_2332);
xnor U1898 (N_1898,In_3087,In_1577);
nand U1899 (N_1899,In_1926,In_521);
nor U1900 (N_1900,In_2947,In_2794);
and U1901 (N_1901,In_586,In_3709);
xnor U1902 (N_1902,In_1050,In_4326);
nor U1903 (N_1903,In_1147,In_553);
nand U1904 (N_1904,In_3972,In_707);
or U1905 (N_1905,In_4165,In_2365);
nor U1906 (N_1906,In_2414,In_1193);
xor U1907 (N_1907,In_3899,In_1776);
or U1908 (N_1908,In_1595,In_4526);
nand U1909 (N_1909,In_573,In_16);
and U1910 (N_1910,In_759,In_2105);
or U1911 (N_1911,In_3233,In_4234);
or U1912 (N_1912,In_4691,In_2502);
and U1913 (N_1913,In_1834,In_4961);
nand U1914 (N_1914,In_3028,In_3339);
or U1915 (N_1915,In_2550,In_4533);
and U1916 (N_1916,In_1113,In_2965);
nand U1917 (N_1917,In_1105,In_2190);
and U1918 (N_1918,In_684,In_4116);
nor U1919 (N_1919,In_809,In_4378);
or U1920 (N_1920,In_4638,In_3536);
xnor U1921 (N_1921,In_1035,In_1407);
or U1922 (N_1922,In_1134,In_1611);
nand U1923 (N_1923,In_4584,In_523);
nor U1924 (N_1924,In_1220,In_2682);
xor U1925 (N_1925,In_1513,In_4244);
or U1926 (N_1926,In_3772,In_656);
nand U1927 (N_1927,In_3853,In_4405);
xnor U1928 (N_1928,In_939,In_3730);
nand U1929 (N_1929,In_2159,In_79);
nand U1930 (N_1930,In_121,In_3957);
xor U1931 (N_1931,In_2775,In_1097);
or U1932 (N_1932,In_4896,In_3878);
nand U1933 (N_1933,In_4484,In_3892);
nand U1934 (N_1934,In_4518,In_1698);
nand U1935 (N_1935,In_4249,In_1122);
or U1936 (N_1936,In_4434,In_3787);
nand U1937 (N_1937,In_2943,In_2928);
or U1938 (N_1938,In_2038,In_4158);
nor U1939 (N_1939,In_1029,In_1846);
or U1940 (N_1940,In_2878,In_4678);
xor U1941 (N_1941,In_120,In_3595);
or U1942 (N_1942,In_3783,In_4934);
nor U1943 (N_1943,In_2929,In_838);
and U1944 (N_1944,In_4174,In_495);
nand U1945 (N_1945,In_2344,In_1635);
or U1946 (N_1946,In_3557,In_3485);
and U1947 (N_1947,In_1678,In_516);
nand U1948 (N_1948,In_1136,In_4569);
or U1949 (N_1949,In_314,In_57);
or U1950 (N_1950,In_149,In_3571);
nand U1951 (N_1951,In_4215,In_2070);
or U1952 (N_1952,In_2285,In_3177);
or U1953 (N_1953,In_2021,In_1888);
nand U1954 (N_1954,In_1309,In_3501);
xnor U1955 (N_1955,In_2893,In_2057);
nor U1956 (N_1956,In_3583,In_2838);
nand U1957 (N_1957,In_512,In_3626);
xor U1958 (N_1958,In_4232,In_1961);
and U1959 (N_1959,In_1804,In_146);
or U1960 (N_1960,In_3614,In_1875);
nand U1961 (N_1961,In_4213,In_555);
nand U1962 (N_1962,In_2944,In_1641);
nand U1963 (N_1963,In_224,In_3317);
or U1964 (N_1964,In_4105,In_2586);
nor U1965 (N_1965,In_2375,In_696);
xnor U1966 (N_1966,In_1878,In_3715);
xnor U1967 (N_1967,In_1001,In_3526);
and U1968 (N_1968,In_1552,In_698);
xnor U1969 (N_1969,In_2907,In_4288);
or U1970 (N_1970,In_350,In_2612);
nor U1971 (N_1971,In_1718,In_339);
or U1972 (N_1972,In_4508,In_2903);
nand U1973 (N_1973,In_4205,In_1414);
nor U1974 (N_1974,In_4491,In_2596);
xor U1975 (N_1975,In_1646,In_2424);
or U1976 (N_1976,In_3310,In_2593);
or U1977 (N_1977,In_2565,In_3585);
xor U1978 (N_1978,In_548,In_4783);
xor U1979 (N_1979,In_955,In_2266);
nor U1980 (N_1980,In_227,In_3484);
or U1981 (N_1981,In_4535,In_1032);
nand U1982 (N_1982,In_3561,In_4828);
or U1983 (N_1983,In_1008,In_317);
nand U1984 (N_1984,In_4696,In_4775);
xor U1985 (N_1985,In_713,In_2175);
nand U1986 (N_1986,In_387,In_4591);
nor U1987 (N_1987,In_3918,In_2289);
xnor U1988 (N_1988,In_3246,In_572);
xnor U1989 (N_1989,In_3156,In_4201);
or U1990 (N_1990,In_1350,In_4671);
or U1991 (N_1991,In_3616,In_1176);
and U1992 (N_1992,In_4954,In_1498);
or U1993 (N_1993,In_2413,In_3403);
or U1994 (N_1994,In_1494,In_3026);
nor U1995 (N_1995,In_823,In_3274);
and U1996 (N_1996,In_3083,In_2174);
and U1997 (N_1997,In_2911,In_4020);
nor U1998 (N_1998,In_319,In_4880);
nand U1999 (N_1999,In_5,In_3955);
or U2000 (N_2000,In_3248,N_1096);
or U2001 (N_2001,N_938,In_2046);
xnor U2002 (N_2002,N_84,N_1929);
xor U2003 (N_2003,N_1656,In_4571);
or U2004 (N_2004,N_90,In_936);
xnor U2005 (N_2005,In_2137,N_689);
xor U2006 (N_2006,N_1380,N_889);
or U2007 (N_2007,N_57,In_1524);
nor U2008 (N_2008,In_4605,N_1541);
or U2009 (N_2009,N_1359,In_2298);
and U2010 (N_2010,N_957,In_4404);
nand U2011 (N_2011,N_1699,In_198);
or U2012 (N_2012,N_1808,In_1675);
or U2013 (N_2013,In_4542,N_273);
nor U2014 (N_2014,In_1546,In_4844);
nand U2015 (N_2015,N_62,In_2420);
nand U2016 (N_2016,In_93,N_97);
or U2017 (N_2017,N_641,In_4051);
nor U2018 (N_2018,N_1769,N_21);
and U2019 (N_2019,N_1141,N_1817);
nor U2020 (N_2020,In_74,N_1634);
nor U2021 (N_2021,N_284,In_504);
nand U2022 (N_2022,N_1353,N_1293);
xor U2023 (N_2023,N_506,N_569);
nand U2024 (N_2024,N_580,N_1983);
or U2025 (N_2025,N_1498,N_660);
xnor U2026 (N_2026,N_1221,N_192);
xnor U2027 (N_2027,N_605,In_4354);
and U2028 (N_2028,N_619,N_220);
xnor U2029 (N_2029,In_3817,In_156);
nand U2030 (N_2030,N_1282,In_1695);
and U2031 (N_2031,N_1672,N_1200);
nor U2032 (N_2032,N_1617,In_3965);
and U2033 (N_2033,In_2479,N_1532);
nand U2034 (N_2034,N_1098,N_1473);
and U2035 (N_2035,In_647,N_261);
and U2036 (N_2036,N_807,In_3949);
nor U2037 (N_2037,N_433,N_1788);
nand U2038 (N_2038,In_1153,In_528);
and U2039 (N_2039,N_190,N_82);
and U2040 (N_2040,In_2905,N_1618);
nor U2041 (N_2041,In_4598,N_1103);
or U2042 (N_2042,N_814,N_684);
and U2043 (N_2043,In_1972,In_397);
or U2044 (N_2044,N_1657,In_488);
nand U2045 (N_2045,N_932,N_1217);
or U2046 (N_2046,N_670,N_36);
xnor U2047 (N_2047,N_1492,N_1058);
or U2048 (N_2048,N_118,In_2379);
and U2049 (N_2049,In_2443,N_718);
nand U2050 (N_2050,N_625,N_101);
and U2051 (N_2051,N_268,N_747);
or U2052 (N_2052,In_3350,N_757);
nor U2053 (N_2053,In_3795,N_1873);
and U2054 (N_2054,In_4336,N_1362);
xnor U2055 (N_2055,In_883,N_1501);
xnor U2056 (N_2056,In_4104,N_448);
xnor U2057 (N_2057,In_3266,N_637);
and U2058 (N_2058,N_432,In_366);
nand U2059 (N_2059,N_1726,In_744);
and U2060 (N_2060,In_2649,N_1458);
and U2061 (N_2061,In_2533,In_2509);
and U2062 (N_2062,N_967,N_1561);
or U2063 (N_2063,N_1211,N_324);
or U2064 (N_2064,N_672,N_221);
or U2065 (N_2065,In_3639,N_590);
xnor U2066 (N_2066,N_1953,N_1874);
nand U2067 (N_2067,In_550,N_1327);
or U2068 (N_2068,In_4838,N_917);
and U2069 (N_2069,In_3862,In_2826);
nor U2070 (N_2070,In_1466,N_1937);
xor U2071 (N_2071,N_1637,N_617);
and U2072 (N_2072,In_933,N_1785);
and U2073 (N_2073,N_934,N_279);
and U2074 (N_2074,N_736,In_4362);
and U2075 (N_2075,N_1170,In_3740);
xor U2076 (N_2076,N_11,N_965);
xnor U2077 (N_2077,N_642,N_145);
nor U2078 (N_2078,N_1622,N_1895);
and U2079 (N_2079,N_1643,N_1190);
nand U2080 (N_2080,N_979,In_98);
xor U2081 (N_2081,In_3737,In_354);
nor U2082 (N_2082,N_851,In_4938);
nor U2083 (N_2083,N_1497,N_1166);
nor U2084 (N_2084,N_958,In_4628);
xor U2085 (N_2085,In_4269,N_1333);
and U2086 (N_2086,N_1973,N_1163);
and U2087 (N_2087,In_4699,N_150);
or U2088 (N_2088,N_479,N_1340);
nor U2089 (N_2089,N_528,In_1040);
xnor U2090 (N_2090,N_1328,N_1240);
or U2091 (N_2091,In_4543,In_3920);
and U2092 (N_2092,N_3,In_720);
or U2093 (N_2093,N_45,N_547);
or U2094 (N_2094,In_1208,N_1354);
nand U2095 (N_2095,In_194,N_1352);
xor U2096 (N_2096,N_1412,N_1626);
xor U2097 (N_2097,N_1706,N_147);
and U2098 (N_2098,N_1204,N_995);
nor U2099 (N_2099,N_413,N_1140);
nand U2100 (N_2100,N_1631,In_4991);
and U2101 (N_2101,N_1888,N_367);
nand U2102 (N_2102,In_1913,In_3425);
and U2103 (N_2103,In_1714,N_700);
and U2104 (N_2104,In_1962,In_655);
nor U2105 (N_2105,N_1077,N_1958);
nor U2106 (N_2106,N_1736,N_163);
nor U2107 (N_2107,In_4429,In_1472);
or U2108 (N_2108,In_2354,N_792);
nor U2109 (N_2109,N_1214,N_463);
and U2110 (N_2110,N_1148,N_1243);
or U2111 (N_2111,N_833,N_1165);
or U2112 (N_2112,N_293,N_1324);
nand U2113 (N_2113,In_3841,In_2335);
or U2114 (N_2114,N_909,N_1833);
or U2115 (N_2115,N_225,In_3463);
nand U2116 (N_2116,N_464,N_1158);
or U2117 (N_2117,N_505,In_2849);
xor U2118 (N_2118,N_716,N_709);
nand U2119 (N_2119,N_1915,N_1427);
nor U2120 (N_2120,N_89,N_592);
xnor U2121 (N_2121,N_447,N_238);
nand U2122 (N_2122,N_564,N_1731);
and U2123 (N_2123,In_1112,N_1824);
nand U2124 (N_2124,In_2725,N_96);
or U2125 (N_2125,N_1811,In_126);
and U2126 (N_2126,N_196,N_1091);
or U2127 (N_2127,N_1898,N_1287);
xnor U2128 (N_2128,In_993,N_1691);
nor U2129 (N_2129,N_407,N_406);
and U2130 (N_2130,N_1988,N_52);
nor U2131 (N_2131,N_338,N_1518);
nand U2132 (N_2132,N_30,In_2796);
nor U2133 (N_2133,In_729,N_944);
or U2134 (N_2134,N_332,In_2979);
nand U2135 (N_2135,N_632,N_514);
nor U2136 (N_2136,In_3426,N_711);
xor U2137 (N_2137,N_1981,N_1577);
and U2138 (N_2138,N_1993,In_4768);
or U2139 (N_2139,N_576,N_1239);
and U2140 (N_2140,N_1055,N_1080);
xor U2141 (N_2141,N_589,In_4917);
and U2142 (N_2142,In_3136,In_1821);
nand U2143 (N_2143,N_1564,N_263);
nand U2144 (N_2144,N_1703,N_808);
or U2145 (N_2145,N_782,N_8);
nor U2146 (N_2146,N_1,N_305);
nor U2147 (N_2147,N_497,N_556);
nand U2148 (N_2148,In_4141,N_1540);
or U2149 (N_2149,N_160,N_1635);
and U2150 (N_2150,In_602,In_3200);
or U2151 (N_2151,In_2268,N_1343);
nor U2152 (N_2152,N_827,N_167);
nand U2153 (N_2153,N_1692,In_3437);
nand U2154 (N_2154,In_3680,N_910);
nor U2155 (N_2155,N_1432,N_1060);
nor U2156 (N_2156,In_1571,N_188);
or U2157 (N_2157,In_2505,In_3973);
and U2158 (N_2158,N_651,In_3073);
or U2159 (N_2159,N_1265,N_1076);
nand U2160 (N_2160,N_353,In_2055);
nor U2161 (N_2161,In_1604,N_1863);
xor U2162 (N_2162,N_1490,In_3333);
xor U2163 (N_2163,N_1868,N_1329);
nor U2164 (N_2164,N_1321,N_758);
and U2165 (N_2165,In_31,In_2439);
nor U2166 (N_2166,In_4331,In_3922);
or U2167 (N_2167,N_1303,In_953);
or U2168 (N_2168,N_1700,N_1157);
xnor U2169 (N_2169,In_4927,N_210);
nor U2170 (N_2170,N_1482,N_1586);
xor U2171 (N_2171,In_1151,N_1291);
nand U2172 (N_2172,N_1685,N_1297);
and U2173 (N_2173,N_1790,N_1168);
xor U2174 (N_2174,N_1230,N_1809);
nor U2175 (N_2175,In_4385,N_1687);
nor U2176 (N_2176,N_1510,In_2727);
and U2177 (N_2177,N_1308,In_897);
or U2178 (N_2178,N_1526,N_1879);
xor U2179 (N_2179,In_2766,In_2683);
nor U2180 (N_2180,In_1921,In_2500);
nand U2181 (N_2181,N_743,N_1784);
nor U2182 (N_2182,N_319,N_1882);
and U2183 (N_2183,N_760,In_2168);
and U2184 (N_2184,In_447,In_4587);
and U2185 (N_2185,N_896,In_2372);
xnor U2186 (N_2186,In_2606,In_3088);
xor U2187 (N_2187,N_1733,In_3399);
and U2188 (N_2188,In_2655,N_1536);
nor U2189 (N_2189,N_951,N_1529);
xor U2190 (N_2190,N_355,In_3736);
and U2191 (N_2191,N_132,N_955);
nand U2192 (N_2192,In_3313,N_1111);
or U2193 (N_2193,N_1611,In_542);
or U2194 (N_2194,N_1686,N_1894);
xnor U2195 (N_2195,N_1160,In_678);
nand U2196 (N_2196,N_1917,In_4366);
or U2197 (N_2197,N_390,In_3187);
nand U2198 (N_2198,N_1311,In_3934);
nor U2199 (N_2199,In_4521,In_3289);
or U2200 (N_2200,In_2111,N_1557);
and U2201 (N_2201,N_1903,N_1438);
nor U2202 (N_2202,N_1194,N_471);
nand U2203 (N_2203,N_1825,N_173);
or U2204 (N_2204,N_242,In_1121);
xnor U2205 (N_2205,In_736,In_1246);
and U2206 (N_2206,N_1082,N_175);
xor U2207 (N_2207,In_1118,N_1390);
or U2208 (N_2208,N_712,N_1835);
and U2209 (N_2209,N_358,N_1559);
xnor U2210 (N_2210,In_4702,N_1447);
and U2211 (N_2211,N_812,In_1692);
xor U2212 (N_2212,N_140,N_1048);
nor U2213 (N_2213,In_1603,N_1583);
nand U2214 (N_2214,N_538,In_1687);
xor U2215 (N_2215,N_1219,In_4516);
nor U2216 (N_2216,N_230,N_348);
and U2217 (N_2217,N_285,N_1468);
xnor U2218 (N_2218,N_71,N_1695);
and U2219 (N_2219,N_26,N_943);
xor U2220 (N_2220,N_503,N_1227);
or U2221 (N_2221,N_873,N_732);
nand U2222 (N_2222,N_297,N_231);
and U2223 (N_2223,N_1403,N_1511);
and U2224 (N_2224,In_1271,N_1436);
xnor U2225 (N_2225,N_1312,In_3477);
or U2226 (N_2226,N_1999,In_270);
xnor U2227 (N_2227,N_630,In_2966);
xor U2228 (N_2228,In_4195,N_594);
and U2229 (N_2229,N_1451,N_417);
and U2230 (N_2230,N_863,N_733);
or U2231 (N_2231,N_767,N_1112);
nand U2232 (N_2232,In_2726,N_1252);
nor U2233 (N_2233,N_161,In_1004);
nor U2234 (N_2234,N_1885,N_1576);
xnor U2235 (N_2235,In_1087,In_949);
or U2236 (N_2236,N_989,In_4345);
nand U2237 (N_2237,In_2615,In_3061);
xor U2238 (N_2238,N_616,N_1976);
nor U2239 (N_2239,N_855,N_1355);
xor U2240 (N_2240,N_1425,N_1138);
nand U2241 (N_2241,N_690,In_3582);
xnor U2242 (N_2242,N_746,N_1969);
nand U2243 (N_2243,N_1544,N_1269);
nor U2244 (N_2244,N_1787,N_815);
nand U2245 (N_2245,N_1043,N_115);
or U2246 (N_2246,In_4807,N_601);
or U2247 (N_2247,N_42,In_619);
xor U2248 (N_2248,In_3063,In_4898);
nor U2249 (N_2249,In_1431,N_217);
nand U2250 (N_2250,In_4765,N_973);
and U2251 (N_2251,N_1404,N_112);
and U2252 (N_2252,N_1930,N_1244);
nand U2253 (N_2253,N_829,N_510);
nor U2254 (N_2254,N_1857,In_1305);
nor U2255 (N_2255,N_1923,N_201);
nor U2256 (N_2256,N_624,N_1569);
and U2257 (N_2257,In_3391,In_4180);
nor U2258 (N_2258,N_898,N_702);
or U2259 (N_2259,N_1712,In_3036);
nor U2260 (N_2260,N_1250,N_571);
and U2261 (N_2261,N_978,N_1514);
nor U2262 (N_2262,N_202,N_1487);
and U2263 (N_2263,N_780,N_1539);
nand U2264 (N_2264,N_956,N_55);
xor U2265 (N_2265,In_4097,N_22);
or U2266 (N_2266,N_1073,In_4012);
nor U2267 (N_2267,N_890,N_1850);
nand U2268 (N_2268,N_1360,N_195);
nand U2269 (N_2269,N_1476,N_1842);
nand U2270 (N_2270,In_3990,In_2401);
nor U2271 (N_2271,In_2620,In_703);
xnor U2272 (N_2272,In_1191,N_727);
and U2273 (N_2273,N_1800,N_1040);
and U2274 (N_2274,In_4310,N_125);
nand U2275 (N_2275,N_416,In_1241);
nand U2276 (N_2276,In_2548,In_1661);
xnor U2277 (N_2277,N_1548,N_686);
or U2278 (N_2278,N_1867,In_3393);
or U2279 (N_2279,N_1791,N_1053);
nand U2280 (N_2280,In_4627,In_3442);
nor U2281 (N_2281,N_106,In_3663);
and U2282 (N_2282,In_1890,N_46);
xnor U2283 (N_2283,N_903,N_1897);
nor U2284 (N_2284,N_1987,N_1248);
or U2285 (N_2285,N_609,N_1891);
nand U2286 (N_2286,N_1620,In_2493);
or U2287 (N_2287,N_288,N_257);
nand U2288 (N_2288,In_2535,N_1907);
or U2289 (N_2289,In_2823,N_1862);
and U2290 (N_2290,In_2779,N_1374);
nor U2291 (N_2291,N_919,N_611);
or U2292 (N_2292,N_908,N_1609);
and U2293 (N_2293,In_4305,In_2113);
nor U2294 (N_2294,N_489,N_100);
or U2295 (N_2295,In_1732,N_1963);
xor U2296 (N_2296,In_4623,N_1991);
or U2297 (N_2297,In_620,In_4962);
nor U2298 (N_2298,N_557,In_3739);
and U2299 (N_2299,N_467,In_1511);
and U2300 (N_2300,N_1520,In_3234);
and U2301 (N_2301,N_931,N_334);
or U2302 (N_2302,In_2643,In_1446);
nor U2303 (N_2303,N_937,N_404);
nand U2304 (N_2304,N_181,In_3508);
nand U2305 (N_2305,N_618,In_3854);
or U2306 (N_2306,In_132,N_1056);
nand U2307 (N_2307,N_638,In_4813);
or U2308 (N_2308,In_805,N_1491);
xnor U2309 (N_2309,N_382,N_323);
and U2310 (N_2310,In_3933,N_253);
and U2311 (N_2311,In_1869,In_870);
and U2312 (N_2312,N_1286,In_4131);
or U2313 (N_2313,N_549,N_1783);
xnor U2314 (N_2314,In_3281,N_705);
nand U2315 (N_2315,N_1792,N_1603);
nor U2316 (N_2316,N_1274,N_1276);
nand U2317 (N_2317,N_484,In_1522);
xnor U2318 (N_2318,N_1348,N_843);
xnor U2319 (N_2319,In_479,N_737);
xnor U2320 (N_2320,In_2209,In_1247);
nor U2321 (N_2321,N_1639,In_2359);
nor U2322 (N_2322,In_4675,N_1805);
nand U2323 (N_2323,N_43,N_1162);
xnor U2324 (N_2324,In_4566,In_3924);
or U2325 (N_2325,N_176,In_1161);
xor U2326 (N_2326,In_4408,In_2013);
nor U2327 (N_2327,N_1568,In_418);
or U2328 (N_2328,N_1319,N_1300);
and U2329 (N_2329,N_719,N_1046);
and U2330 (N_2330,N_708,In_4560);
xor U2331 (N_2331,In_518,In_2841);
or U2332 (N_2332,N_486,N_120);
nand U2333 (N_2333,N_487,N_316);
xor U2334 (N_2334,N_1992,N_1024);
nand U2335 (N_2335,In_3195,In_1762);
nand U2336 (N_2336,N_1616,N_491);
or U2337 (N_2337,N_1258,N_1718);
or U2338 (N_2338,In_1837,N_1851);
or U2339 (N_2339,N_1592,In_1658);
or U2340 (N_2340,N_1433,N_87);
and U2341 (N_2341,In_203,In_2059);
nor U2342 (N_2342,In_228,N_1499);
nor U2343 (N_2343,N_357,N_1967);
nand U2344 (N_2344,N_880,N_602);
nor U2345 (N_2345,In_4200,In_4467);
and U2346 (N_2346,N_392,N_1453);
xor U2347 (N_2347,N_1384,N_91);
and U2348 (N_2348,N_354,N_1067);
and U2349 (N_2349,In_3174,N_1015);
nor U2350 (N_2350,N_954,N_440);
nand U2351 (N_2351,In_3148,N_1777);
or U2352 (N_2352,In_3345,In_4815);
or U2353 (N_2353,In_1715,N_1011);
and U2354 (N_2354,In_669,In_1758);
xnor U2355 (N_2355,N_1256,N_1180);
and U2356 (N_2356,N_72,In_4863);
nand U2357 (N_2357,In_1833,N_1020);
nand U2358 (N_2358,In_610,In_1649);
xor U2359 (N_2359,N_1780,N_1560);
xor U2360 (N_2360,N_272,N_1475);
xnor U2361 (N_2361,In_4072,In_1091);
xor U2362 (N_2362,In_708,N_1912);
and U2363 (N_2363,N_545,In_443);
or U2364 (N_2364,N_135,N_466);
and U2365 (N_2365,In_996,In_4818);
and U2366 (N_2366,In_1660,N_488);
nor U2367 (N_2367,In_3479,N_1175);
nand U2368 (N_2368,In_718,N_318);
or U2369 (N_2369,N_465,In_2557);
nor U2370 (N_2370,N_19,N_840);
and U2371 (N_2371,In_4826,In_2906);
or U2372 (N_2372,N_986,In_3482);
or U2373 (N_2373,N_523,N_254);
nor U2374 (N_2374,In_1765,N_645);
or U2375 (N_2375,N_543,N_798);
and U2376 (N_2376,N_159,In_4004);
nor U2377 (N_2377,In_346,N_721);
nor U2378 (N_2378,In_2306,N_1773);
nand U2379 (N_2379,N_1387,In_3551);
nand U2380 (N_2380,In_646,N_1749);
or U2381 (N_2381,N_551,N_838);
and U2382 (N_2382,N_1210,N_769);
or U2383 (N_2383,In_3226,In_4505);
nand U2384 (N_2384,In_1917,N_1573);
nor U2385 (N_2385,N_1670,N_29);
and U2386 (N_2386,N_1209,In_4636);
nand U2387 (N_2387,N_1676,N_1830);
xnor U2388 (N_2388,N_1205,N_1813);
nor U2389 (N_2389,In_576,In_1627);
or U2390 (N_2390,In_1719,N_1893);
and U2391 (N_2391,N_61,N_842);
nor U2392 (N_2392,In_2291,N_475);
nor U2393 (N_2393,N_1357,N_93);
xor U2394 (N_2394,In_589,In_3307);
nor U2395 (N_2395,In_2459,In_1927);
and U2396 (N_2396,N_124,N_977);
nand U2397 (N_2397,N_531,In_166);
nand U2398 (N_2398,In_2811,N_1028);
and U2399 (N_2399,In_3609,In_1019);
or U2400 (N_2400,N_982,N_169);
xnor U2401 (N_2401,N_741,N_1723);
nor U2402 (N_2402,In_4901,N_1904);
xor U2403 (N_2403,N_1174,In_1816);
xor U2404 (N_2404,In_3559,In_180);
xor U2405 (N_2405,N_1607,In_4019);
and U2406 (N_2406,N_1262,In_4823);
and U2407 (N_2407,N_1237,N_1644);
and U2408 (N_2408,N_1445,N_1755);
nand U2409 (N_2409,In_1377,N_1588);
xnor U2410 (N_2410,In_873,In_3294);
nand U2411 (N_2411,N_255,N_1302);
and U2412 (N_2412,In_1971,N_0);
or U2413 (N_2413,N_1330,N_371);
and U2414 (N_2414,N_99,N_246);
nor U2415 (N_2415,N_820,In_832);
nor U2416 (N_2416,N_1574,N_56);
nand U2417 (N_2417,In_237,N_541);
and U2418 (N_2418,N_1843,In_3435);
and U2419 (N_2419,N_1645,N_114);
nor U2420 (N_2420,N_1696,N_1507);
nor U2421 (N_2421,N_110,In_348);
nor U2422 (N_2422,N_994,N_717);
nand U2423 (N_2423,N_60,N_184);
xnor U2424 (N_2424,N_1980,N_706);
nor U2425 (N_2425,N_47,In_2369);
nand U2426 (N_2426,N_380,N_1189);
nand U2427 (N_2427,N_935,In_1729);
or U2428 (N_2428,N_1865,In_2991);
or U2429 (N_2429,N_819,In_770);
nor U2430 (N_2430,N_1750,N_1169);
xnor U2431 (N_2431,In_1,N_1605);
xnor U2432 (N_2432,N_810,N_212);
nand U2433 (N_2433,N_1985,N_336);
nor U2434 (N_2434,In_4762,N_1393);
nor U2435 (N_2435,N_94,In_2508);
xor U2436 (N_2436,N_1296,N_1594);
nand U2437 (N_2437,In_424,In_1023);
nand U2438 (N_2438,N_786,N_350);
nor U2439 (N_2439,N_1065,In_42);
and U2440 (N_2440,N_1567,In_202);
nand U2441 (N_2441,N_874,N_1477);
nor U2442 (N_2442,In_794,In_3409);
or U2443 (N_2443,N_349,N_1461);
nor U2444 (N_2444,In_1676,In_4254);
xnor U2445 (N_2445,N_294,N_1062);
and U2446 (N_2446,N_975,N_1565);
nand U2447 (N_2447,In_588,In_292);
nand U2448 (N_2448,N_1932,In_2232);
nand U2449 (N_2449,N_1836,N_1834);
nand U2450 (N_2450,N_1819,N_1094);
nand U2451 (N_2451,In_1712,N_1766);
nand U2452 (N_2452,In_958,N_968);
or U2453 (N_2453,N_1326,In_608);
xnor U2454 (N_2454,N_731,N_772);
nand U2455 (N_2455,N_241,N_813);
nor U2456 (N_2456,N_25,N_247);
or U2457 (N_2457,In_297,In_4935);
xor U2458 (N_2458,N_1251,N_312);
xor U2459 (N_2459,In_1165,N_1849);
nor U2460 (N_2460,In_3904,N_1129);
nor U2461 (N_2461,N_148,N_1488);
or U2462 (N_2462,N_1041,N_209);
xor U2463 (N_2463,In_357,In_4446);
or U2464 (N_2464,In_0,N_1727);
nand U2465 (N_2465,In_3638,N_1376);
nand U2466 (N_2466,N_197,N_1125);
nor U2467 (N_2467,N_1896,N_600);
and U2468 (N_2468,N_905,In_964);
or U2469 (N_2469,In_3686,N_1797);
xnor U2470 (N_2470,In_4956,In_4618);
and U2471 (N_2471,In_9,N_871);
or U2472 (N_2472,N_1309,N_1628);
or U2473 (N_2473,In_4737,N_1386);
and U2474 (N_2474,N_442,In_103);
xor U2475 (N_2475,In_3096,In_2640);
nor U2476 (N_2476,N_1426,N_612);
nor U2477 (N_2477,In_1452,In_1986);
xnor U2478 (N_2478,In_1742,N_142);
xnor U2479 (N_2479,N_468,N_1954);
or U2480 (N_2480,In_3074,N_191);
nor U2481 (N_2481,In_4132,N_575);
nand U2482 (N_2482,In_2428,N_997);
nand U2483 (N_2483,N_1633,N_710);
nand U2484 (N_2484,N_568,N_724);
or U2485 (N_2485,N_1459,N_1457);
nand U2486 (N_2486,N_374,N_728);
xnor U2487 (N_2487,N_1515,In_1996);
or U2488 (N_2488,In_2799,N_226);
and U2489 (N_2489,N_1619,In_4361);
or U2490 (N_2490,In_3793,In_1125);
and U2491 (N_2491,N_587,In_76);
or U2492 (N_2492,In_332,N_826);
nor U2493 (N_2493,In_341,N_280);
nor U2494 (N_2494,N_751,N_1590);
nand U2495 (N_2495,N_68,N_290);
and U2496 (N_2496,N_13,N_1610);
nand U2497 (N_2497,N_566,In_3510);
and U2498 (N_2498,N_330,N_1113);
or U2499 (N_2499,N_275,N_1655);
nand U2500 (N_2500,N_483,N_834);
nor U2501 (N_2501,N_317,In_1907);
or U2502 (N_2502,N_1092,In_2647);
nor U2503 (N_2503,N_570,N_902);
or U2504 (N_2504,N_781,N_1902);
and U2505 (N_2505,N_411,N_1935);
and U2506 (N_2506,In_4894,In_3926);
or U2507 (N_2507,N_1760,In_2828);
nand U2508 (N_2508,In_2088,In_420);
nor U2509 (N_2509,N_1660,N_607);
nor U2510 (N_2510,In_4738,In_1383);
nand U2511 (N_2511,In_855,N_1310);
xor U2512 (N_2512,N_137,N_949);
or U2513 (N_2513,N_203,N_981);
or U2514 (N_2514,N_343,N_1216);
and U2515 (N_2515,In_2097,N_847);
and U2516 (N_2516,In_2099,In_2605);
xor U2517 (N_2517,N_1916,N_723);
or U2518 (N_2518,N_418,N_274);
nand U2519 (N_2519,N_462,In_3545);
nor U2520 (N_2520,In_1139,In_4767);
nor U2521 (N_2521,N_1254,In_3149);
and U2522 (N_2522,N_436,N_495);
nor U2523 (N_2523,N_1083,N_1680);
and U2524 (N_2524,N_1114,In_800);
nor U2525 (N_2525,In_1786,In_4063);
and U2526 (N_2526,N_33,N_1998);
nand U2527 (N_2527,N_1378,In_4857);
nand U2528 (N_2528,N_1747,N_870);
nand U2529 (N_2529,N_1848,N_1922);
nand U2530 (N_2530,N_1346,N_1956);
xor U2531 (N_2531,In_1549,In_3158);
nand U2532 (N_2532,N_1153,In_2708);
nor U2533 (N_2533,N_77,N_1630);
nor U2534 (N_2534,In_4537,N_1272);
or U2535 (N_2535,N_1005,In_927);
xor U2536 (N_2536,N_897,N_1881);
and U2537 (N_2537,In_56,In_4271);
nand U2538 (N_2538,In_3452,In_562);
xor U2539 (N_2539,N_1636,N_400);
nor U2540 (N_2540,N_1295,N_927);
nor U2541 (N_2541,N_1212,In_2446);
and U2542 (N_2542,N_1624,N_963);
xnor U2543 (N_2543,N_453,N_676);
and U2544 (N_2544,In_4044,In_4655);
nand U2545 (N_2545,N_597,N_517);
xor U2546 (N_2546,In_1725,N_1604);
xnor U2547 (N_2547,N_1734,In_3185);
or U2548 (N_2548,N_1012,In_3527);
or U2549 (N_2549,N_675,N_1921);
or U2550 (N_2550,N_846,N_911);
xor U2551 (N_2551,In_3115,N_1572);
or U2552 (N_2552,In_2222,N_877);
xnor U2553 (N_2553,In_4778,In_1937);
xnor U2554 (N_2554,In_2870,N_1648);
and U2555 (N_2555,N_904,N_1156);
xnor U2556 (N_2556,N_375,N_1006);
and U2557 (N_2557,N_1223,N_888);
or U2558 (N_2558,In_3212,N_797);
xor U2559 (N_2559,In_1928,N_1877);
xnor U2560 (N_2560,N_990,In_4169);
or U2561 (N_2561,N_1467,N_40);
or U2562 (N_2562,N_119,N_1106);
nand U2563 (N_2563,N_1016,N_164);
nor U2564 (N_2564,N_243,N_1802);
or U2565 (N_2565,N_697,N_1763);
or U2566 (N_2566,In_4373,N_803);
nand U2567 (N_2567,N_1408,In_2125);
xor U2568 (N_2568,N_869,In_351);
xor U2569 (N_2569,In_937,In_1854);
or U2570 (N_2570,In_2613,N_1948);
nand U2571 (N_2571,N_868,N_482);
nor U2572 (N_2572,In_1363,N_81);
or U2573 (N_2573,In_885,N_153);
nor U2574 (N_2574,In_4739,N_1410);
or U2575 (N_2575,N_1602,In_785);
or U2576 (N_2576,N_791,In_4413);
nand U2577 (N_2577,N_839,N_883);
xor U2578 (N_2578,N_1739,N_755);
nand U2579 (N_2579,N_170,N_837);
xnor U2580 (N_2580,N_693,In_392);
or U2581 (N_2581,N_1423,N_1456);
nor U2582 (N_2582,In_3413,N_959);
and U2583 (N_2583,N_421,N_567);
or U2584 (N_2584,N_1495,N_157);
or U2585 (N_2585,N_740,In_1931);
nand U2586 (N_2586,N_1117,N_527);
or U2587 (N_2587,In_4219,In_4202);
xnor U2588 (N_2588,N_1665,In_2138);
nand U2589 (N_2589,N_1207,N_1960);
or U2590 (N_2590,N_1151,In_2098);
xnor U2591 (N_2591,N_558,In_345);
nor U2592 (N_2592,N_1840,In_4258);
nor U2593 (N_2593,In_2107,N_1290);
and U2594 (N_2594,N_328,N_1122);
nor U2595 (N_2595,N_1064,In_2188);
or U2596 (N_2596,In_1119,N_1553);
and U2597 (N_2597,N_127,N_1100);
or U2598 (N_2598,In_2877,N_1079);
nor U2599 (N_2599,In_578,N_1263);
nor U2600 (N_2600,N_1441,N_596);
and U2601 (N_2601,N_1280,N_364);
xnor U2602 (N_2602,N_1044,In_2974);
nand U2603 (N_2603,In_2740,In_3758);
or U2604 (N_2604,In_2987,N_1220);
nor U2605 (N_2605,N_1858,In_2160);
or U2606 (N_2606,In_3794,N_1193);
and U2607 (N_2607,N_144,N_1335);
or U2608 (N_2608,N_1728,N_1729);
and U2609 (N_2609,N_1679,N_725);
nand U2610 (N_2610,In_4262,In_3285);
nor U2611 (N_2611,N_237,In_836);
nor U2612 (N_2612,In_285,In_2336);
or U2613 (N_2613,N_1332,N_1974);
or U2614 (N_2614,N_730,N_756);
or U2615 (N_2615,N_872,In_4316);
or U2616 (N_2616,N_333,N_849);
nor U2617 (N_2617,N_1743,N_152);
and U2618 (N_2618,N_1247,N_830);
nand U2619 (N_2619,In_255,N_1615);
nand U2620 (N_2620,N_425,N_1994);
or U2621 (N_2621,N_806,N_598);
nand U2622 (N_2622,N_1045,N_313);
or U2623 (N_2623,N_360,N_1029);
xnor U2624 (N_2624,In_3404,In_1952);
and U2625 (N_2625,N_469,In_1214);
and U2626 (N_2626,In_1608,N_1522);
xor U2627 (N_2627,In_4018,N_884);
or U2628 (N_2628,N_1494,In_4017);
and U2629 (N_2629,N_1480,N_1910);
nor U2630 (N_2630,N_831,N_1856);
nand U2631 (N_2631,In_3843,N_1164);
and U2632 (N_2632,N_283,N_1088);
and U2633 (N_2633,In_3275,In_4853);
xnor U2634 (N_2634,N_525,N_1018);
or U2635 (N_2635,N_752,In_4054);
xnor U2636 (N_2636,N_1778,N_533);
nand U2637 (N_2637,In_3778,In_4578);
nor U2638 (N_2638,In_2875,N_1671);
nand U2639 (N_2639,N_1007,N_1523);
or U2640 (N_2640,N_530,In_1291);
or U2641 (N_2641,In_2782,N_864);
or U2642 (N_2642,In_4365,N_351);
or U2643 (N_2643,In_2988,N_635);
nand U2644 (N_2644,N_1756,N_369);
and U2645 (N_2645,N_856,N_1493);
nor U2646 (N_2646,N_337,N_726);
or U2647 (N_2647,N_79,N_1855);
xor U2648 (N_2648,N_1119,In_3215);
or U2649 (N_2649,In_844,In_3392);
or U2650 (N_2650,N_1183,N_1415);
and U2651 (N_2651,N_6,In_2563);
or U2652 (N_2652,N_554,In_859);
and U2653 (N_2653,N_102,In_2224);
xor U2654 (N_2654,In_899,N_1392);
and U2655 (N_2655,In_2387,N_438);
xnor U2656 (N_2656,N_779,N_687);
or U2657 (N_2657,N_1838,N_398);
or U2658 (N_2658,N_969,N_494);
nor U2659 (N_2659,In_2185,N_1762);
or U2660 (N_2660,N_821,N_1229);
and U2661 (N_2661,In_1785,In_510);
and U2662 (N_2662,In_1709,In_1372);
or U2663 (N_2663,N_988,N_1502);
nand U2664 (N_2664,In_3381,N_1500);
or U2665 (N_2665,N_962,N_1177);
nand U2666 (N_2666,N_1349,N_526);
or U2667 (N_2667,In_1593,N_1546);
and U2668 (N_2668,N_1371,N_1496);
and U2669 (N_2669,N_1798,In_1933);
nor U2670 (N_2670,N_98,N_1847);
and U2671 (N_2671,N_1530,N_901);
or U2672 (N_2672,N_947,In_1236);
xor U2673 (N_2673,N_1931,N_1435);
and U2674 (N_2674,N_1759,In_1150);
or U2675 (N_2675,N_1218,N_674);
nor U2676 (N_2676,N_650,In_3896);
nand U2677 (N_2677,N_881,N_377);
or U2678 (N_2678,In_4312,N_1688);
nor U2679 (N_2679,In_3291,N_1010);
xor U2680 (N_2680,In_2203,N_604);
nand U2681 (N_2681,N_1597,N_136);
xnor U2682 (N_2682,N_1213,N_1192);
xnor U2683 (N_2683,N_562,N_205);
or U2684 (N_2684,In_2616,In_3870);
or U2685 (N_2685,In_3072,N_906);
xnor U2686 (N_2686,N_764,N_891);
nand U2687 (N_2687,N_1023,N_269);
xor U2688 (N_2688,In_4347,N_584);
nand U2689 (N_2689,In_1957,N_331);
xnor U2690 (N_2690,In_3159,N_384);
xnor U2691 (N_2691,N_895,N_1884);
nor U2692 (N_2692,In_209,In_2918);
or U2693 (N_2693,N_1641,N_1261);
xor U2694 (N_2694,N_1398,N_1866);
nor U2695 (N_2695,In_3890,N_1066);
xor U2696 (N_2696,N_1249,N_480);
nor U2697 (N_2697,N_368,In_2461);
nor U2698 (N_2698,N_1761,In_1242);
nor U2699 (N_2699,In_2486,N_445);
or U2700 (N_2700,N_1652,In_4937);
and U2701 (N_2701,In_3402,N_1052);
nor U2702 (N_2702,N_366,N_394);
nand U2703 (N_2703,N_1279,In_2843);
or U2704 (N_2704,N_550,N_422);
or U2705 (N_2705,N_1919,N_1677);
or U2706 (N_2706,N_673,N_402);
xor U2707 (N_2707,N_14,N_1707);
nor U2708 (N_2708,N_410,N_439);
and U2709 (N_2709,N_1132,In_3376);
nor U2710 (N_2710,N_1402,In_2005);
xor U2711 (N_2711,N_1955,N_405);
or U2712 (N_2712,In_233,N_1283);
or U2713 (N_2713,N_1547,In_740);
or U2714 (N_2714,In_1703,N_1545);
or U2715 (N_2715,N_428,N_1464);
xnor U2716 (N_2716,In_414,N_1150);
and U2717 (N_2717,N_1899,N_1126);
nor U2718 (N_2718,N_1109,N_862);
nand U2719 (N_2719,N_713,N_1394);
or U2720 (N_2720,In_4532,N_1019);
xor U2721 (N_2721,N_23,N_1854);
and U2722 (N_2722,N_1370,In_4281);
nand U2723 (N_2723,N_768,In_3131);
and U2724 (N_2724,N_1178,N_1191);
nor U2725 (N_2725,N_1225,N_1938);
nand U2726 (N_2726,N_688,N_1187);
or U2727 (N_2727,N_37,In_282);
nor U2728 (N_2728,N_1719,In_4718);
and U2729 (N_2729,N_683,In_4686);
nor U2730 (N_2730,In_4360,In_525);
nand U2731 (N_2731,In_4707,N_1925);
nand U2732 (N_2732,In_2982,In_726);
nand U2733 (N_2733,In_2820,In_3091);
nor U2734 (N_2734,N_522,N_980);
nor U2735 (N_2735,In_1944,N_714);
nor U2736 (N_2736,N_1416,N_1381);
or U2737 (N_2737,In_2784,N_207);
or U2738 (N_2738,N_1417,N_1134);
nand U2739 (N_2739,In_2012,N_1962);
xnor U2740 (N_2740,In_1694,N_1682);
or U2741 (N_2741,N_1057,N_970);
nor U2742 (N_2742,In_4995,N_1042);
and U2743 (N_2743,N_298,In_1985);
and U2744 (N_2744,N_1270,In_3909);
xor U2745 (N_2745,N_1596,In_975);
or U2746 (N_2746,N_249,In_2484);
xnor U2747 (N_2747,In_670,In_821);
nor U2748 (N_2748,N_1528,N_1732);
nor U2749 (N_2749,In_2564,In_4419);
xor U2750 (N_2750,N_649,N_1669);
nand U2751 (N_2751,N_701,N_704);
or U2752 (N_2752,In_4369,N_1504);
and U2753 (N_2753,N_998,N_1764);
nor U2754 (N_2754,In_2946,N_1782);
and U2755 (N_2755,In_4980,In_3834);
nor U2756 (N_2756,N_399,N_753);
xor U2757 (N_2757,In_1379,In_628);
nor U2758 (N_2758,N_386,In_1078);
and U2759 (N_2759,N_1578,N_250);
nor U2760 (N_2760,N_363,N_1683);
xnor U2761 (N_2761,N_952,N_1068);
nor U2762 (N_2762,N_240,N_1632);
or U2763 (N_2763,N_579,In_3071);
or U2764 (N_2764,In_1461,In_1773);
nor U2765 (N_2765,N_1936,N_1259);
or U2766 (N_2766,In_3314,N_857);
or U2767 (N_2767,N_960,N_1009);
nand U2768 (N_2768,N_1906,N_1751);
xnor U2769 (N_2769,In_2817,N_321);
or U2770 (N_2770,N_1924,N_1549);
nor U2771 (N_2771,N_204,N_409);
and U2772 (N_2772,In_1349,In_2292);
and U2773 (N_2773,In_3775,N_1301);
and U2774 (N_2774,In_3541,In_163);
and U2775 (N_2775,N_451,N_1555);
xnor U2776 (N_2776,In_4541,N_373);
nand U2777 (N_2777,In_876,N_481);
nor U2778 (N_2778,In_4556,In_2072);
nor U2779 (N_2779,N_1563,N_1720);
and U2780 (N_2780,N_206,In_2437);
or U2781 (N_2781,N_73,N_1986);
xnor U2782 (N_2782,N_915,In_2429);
and U2783 (N_2783,N_1338,In_2317);
or U2784 (N_2784,In_3989,N_1123);
and U2785 (N_2785,In_2805,N_1186);
or U2786 (N_2786,In_3428,N_738);
or U2787 (N_2787,N_165,N_520);
xnor U2788 (N_2788,N_745,In_3879);
nor U2789 (N_2789,N_1664,N_1668);
nor U2790 (N_2790,N_28,N_1273);
nor U2791 (N_2791,In_3897,In_2719);
nand U2792 (N_2792,N_474,N_985);
nand U2793 (N_2793,N_1710,N_216);
or U2794 (N_2794,N_1022,N_1241);
xnor U2795 (N_2795,N_984,N_1271);
or U2796 (N_2796,N_1880,N_578);
or U2797 (N_2797,In_1303,N_1101);
and U2798 (N_2798,N_1804,In_2530);
xor U2799 (N_2799,N_1543,In_4721);
nor U2800 (N_2800,N_227,In_1810);
nand U2801 (N_2801,In_1329,In_944);
nor U2802 (N_2802,N_1503,N_59);
or U2803 (N_2803,N_655,N_1462);
and U2804 (N_2804,N_1350,N_304);
nand U2805 (N_2805,N_1025,N_1037);
nor U2806 (N_2806,In_215,N_389);
nor U2807 (N_2807,N_458,N_1584);
nor U2808 (N_2808,N_770,N_301);
or U2809 (N_2809,N_1774,N_1509);
and U2810 (N_2810,In_755,N_1342);
xor U2811 (N_2811,In_1250,N_1951);
xnor U2812 (N_2812,N_1325,In_2011);
and U2813 (N_2813,In_1503,In_349);
xnor U2814 (N_2814,N_867,In_1775);
xnor U2815 (N_2815,In_2694,N_885);
xnor U2816 (N_2816,N_824,N_67);
and U2817 (N_2817,N_643,N_1775);
or U2818 (N_2818,N_1516,In_1300);
xnor U2819 (N_2819,N_822,In_2066);
and U2820 (N_2820,N_1253,N_784);
and U2821 (N_2821,N_1965,N_224);
nand U2822 (N_2822,N_88,N_1551);
and U2823 (N_2823,N_691,N_103);
nand U2824 (N_2824,In_7,N_1344);
nand U2825 (N_2825,N_748,N_622);
and U2826 (N_2826,In_2531,In_916);
xnor U2827 (N_2827,N_1002,N_233);
and U2828 (N_2828,N_599,N_1806);
nand U2829 (N_2829,In_4439,N_80);
nand U2830 (N_2830,N_848,In_3719);
xor U2831 (N_2831,In_3133,N_548);
or U2832 (N_2832,In_294,N_631);
or U2833 (N_2833,In_1313,N_122);
or U2834 (N_2834,N_1745,N_139);
or U2835 (N_2835,N_1054,In_4978);
nor U2836 (N_2836,In_4225,In_3253);
or U2837 (N_2837,In_2774,N_500);
or U2838 (N_2838,N_1049,N_341);
or U2839 (N_2839,N_1582,In_3431);
nand U2840 (N_2840,N_720,In_2281);
nand U2841 (N_2841,N_1185,In_2704);
or U2842 (N_2842,N_1171,N_78);
nand U2843 (N_2843,In_318,N_51);
nand U2844 (N_2844,N_1831,N_1322);
or U2845 (N_2845,N_1081,N_844);
or U2846 (N_2846,N_121,N_759);
xnor U2847 (N_2847,N_754,N_1570);
nor U2848 (N_2848,In_4473,In_2761);
and U2849 (N_2849,N_1278,N_289);
and U2850 (N_2850,N_302,In_3668);
or U2851 (N_2851,N_818,N_1448);
and U2852 (N_2852,In_4930,In_1301);
nand U2853 (N_2853,N_178,In_4459);
xnor U2854 (N_2854,N_669,N_1034);
xor U2855 (N_2855,N_430,N_1869);
xor U2856 (N_2856,N_379,In_217);
xnor U2857 (N_2857,In_4247,N_1027);
xnor U2858 (N_2858,In_735,N_1714);
and U2859 (N_2859,N_75,N_1437);
xor U2860 (N_2860,N_1465,N_1939);
or U2861 (N_2861,N_789,In_4302);
nand U2862 (N_2862,N_1289,N_166);
nor U2863 (N_2863,N_559,In_3840);
nor U2864 (N_2864,N_86,N_185);
or U2865 (N_2865,N_252,In_1345);
and U2866 (N_2866,N_671,N_64);
and U2867 (N_2867,N_1198,In_2971);
and U2868 (N_2868,N_1822,N_1385);
or U2869 (N_2869,N_1133,N_925);
nor U2870 (N_2870,N_667,N_1107);
or U2871 (N_2871,N_452,N_972);
xor U2872 (N_2872,N_200,In_1263);
and U2873 (N_2873,N_1977,In_1887);
nand U2874 (N_2874,N_444,N_665);
and U2875 (N_2875,N_1124,N_1820);
and U2876 (N_2876,N_54,In_2434);
and U2877 (N_2877,In_2528,In_4706);
nand U2878 (N_2878,N_339,N_1909);
and U2879 (N_2879,N_1828,N_663);
nand U2880 (N_2880,N_1413,N_524);
or U2881 (N_2881,N_1365,In_2989);
and U2882 (N_2882,In_686,N_1298);
xor U2883 (N_2883,N_563,N_765);
or U2884 (N_2884,N_653,N_1388);
and U2885 (N_2885,N_17,In_3692);
or U2886 (N_2886,In_3420,N_1285);
and U2887 (N_2887,N_1460,N_1399);
xor U2888 (N_2888,N_606,In_1508);
xor U2889 (N_2889,N_1554,N_1595);
nand U2890 (N_2890,In_1950,N_1681);
xnor U2891 (N_2891,In_1955,N_1105);
nor U2892 (N_2892,N_1358,N_776);
and U2893 (N_2893,N_936,N_1199);
or U2894 (N_2894,N_983,In_4821);
or U2895 (N_2895,In_4574,N_239);
nand U2896 (N_2896,N_1621,In_1925);
or U2897 (N_2897,N_512,N_1318);
nor U2898 (N_2898,N_680,In_4929);
nand U2899 (N_2899,In_4479,N_1288);
or U2900 (N_2900,In_749,N_586);
nand U2901 (N_2901,In_4068,N_1486);
xor U2902 (N_2902,N_1208,In_465);
nor U2903 (N_2903,N_1708,N_585);
nand U2904 (N_2904,In_3030,In_412);
or U2905 (N_2905,N_5,N_879);
and U2906 (N_2906,In_2050,In_1442);
nor U2907 (N_2907,N_1004,N_615);
nor U2908 (N_2908,N_1484,N_208);
and U2909 (N_2909,In_3818,N_460);
and U2910 (N_2910,In_3124,N_493);
nand U2911 (N_2911,N_1966,N_292);
xor U2912 (N_2912,N_1527,N_383);
nor U2913 (N_2913,N_1172,N_189);
or U2914 (N_2914,N_1864,N_1823);
nand U2915 (N_2915,N_1698,N_1746);
xor U2916 (N_2916,In_506,In_969);
and U2917 (N_2917,In_3271,N_149);
and U2918 (N_2918,N_1666,N_508);
nand U2919 (N_2919,N_15,N_499);
nor U2920 (N_2920,N_1120,N_265);
nand U2921 (N_2921,N_694,N_1926);
nand U2922 (N_2922,N_1339,In_1199);
or U2923 (N_2923,N_1647,N_1334);
nand U2924 (N_2924,In_790,In_1932);
xor U2925 (N_2925,In_4552,N_681);
or U2926 (N_2926,N_1136,N_588);
xor U2927 (N_2927,N_1748,N_95);
nand U2928 (N_2928,N_560,N_1890);
or U2929 (N_2929,N_516,In_3210);
and U2930 (N_2930,N_926,N_322);
and U2931 (N_2931,In_3738,N_654);
and U2932 (N_2932,N_1434,In_3906);
nand U2933 (N_2933,N_344,N_509);
and U2934 (N_2934,N_1737,In_3050);
nand U2935 (N_2935,N_1740,N_1614);
xor U2936 (N_2936,N_1971,N_1401);
and U2937 (N_2937,N_928,N_1446);
nor U2938 (N_2938,In_3287,N_823);
nor U2939 (N_2939,N_1829,N_155);
nor U2940 (N_2940,N_1928,N_1257);
or U2941 (N_2941,N_1650,N_1268);
and U2942 (N_2942,N_661,In_4787);
xnor U2943 (N_2943,N_774,N_1860);
or U2944 (N_2944,N_1070,In_2960);
or U2945 (N_2945,In_1359,N_668);
or U2946 (N_2946,N_1421,N_454);
and U2947 (N_2947,N_1796,In_1064);
and U2948 (N_2948,N_1950,In_3334);
nand U2949 (N_2949,In_768,N_1450);
xnor U2950 (N_2950,N_376,In_598);
nor U2951 (N_2951,N_1942,In_2337);
or U2952 (N_2952,In_453,N_1181);
xor U2953 (N_2953,N_1411,In_2074);
or U2954 (N_2954,In_2645,N_734);
nor U2955 (N_2955,N_1933,N_750);
xnor U2956 (N_2956,N_109,In_4455);
and U2957 (N_2957,N_1786,N_498);
or U2958 (N_2958,In_4874,In_4749);
nor U2959 (N_2959,In_374,In_3336);
nand U2960 (N_2960,N_696,N_1121);
nand U2961 (N_2961,N_1275,In_2355);
and U2962 (N_2962,In_4942,In_4396);
nor U2963 (N_2963,N_420,N_1418);
xor U2964 (N_2964,In_427,N_1228);
nor U2965 (N_2965,N_329,N_1173);
xor U2966 (N_2966,In_3225,N_92);
or U2967 (N_2967,N_1032,N_1781);
nor U2968 (N_2968,In_4923,N_259);
xor U2969 (N_2969,N_308,N_940);
or U2970 (N_2970,N_1149,N_1638);
xor U2971 (N_2971,In_1572,N_1110);
nor U2972 (N_2972,In_3514,In_251);
nor U2973 (N_2973,In_4293,N_1513);
nor U2974 (N_2974,N_1255,N_146);
nand U2975 (N_2975,N_1377,In_4665);
or U2976 (N_2976,In_4846,N_850);
nand U2977 (N_2977,N_1242,In_1195);
and U2978 (N_2978,In_3181,N_1598);
xnor U2979 (N_2979,In_4433,N_1003);
or U2980 (N_2980,N_882,N_1084);
and U2981 (N_2981,N_156,In_1965);
nor U2982 (N_2982,N_1131,N_692);
nor U2983 (N_2983,In_3506,N_271);
or U2984 (N_2984,N_1089,N_1292);
xor U2985 (N_2985,N_1405,N_311);
xor U2986 (N_2986,In_960,N_1463);
nand U2987 (N_2987,N_582,N_685);
or U2988 (N_2988,In_3194,N_1870);
and U2989 (N_2989,In_3308,In_1583);
or U2990 (N_2990,N_1072,N_1097);
nor U2991 (N_2991,N_715,N_1407);
and U2992 (N_2992,In_2515,N_133);
and U2993 (N_2993,In_4664,N_766);
xor U2994 (N_2994,N_614,N_1409);
and U2995 (N_2995,N_455,N_540);
or U2996 (N_2996,N_634,In_1047);
xor U2997 (N_2997,In_3659,In_4519);
and U2998 (N_2998,N_1952,N_1768);
or U2999 (N_2999,In_3971,N_194);
nor U3000 (N_3000,In_1500,N_1331);
xnor U3001 (N_3001,N_63,In_3209);
xnor U3002 (N_3002,N_1927,N_1431);
or U3003 (N_3003,N_1587,N_1717);
xnor U3004 (N_3004,In_4839,N_544);
or U3005 (N_3005,N_529,N_805);
xnor U3006 (N_3006,N_1566,N_811);
nand U3007 (N_3007,N_1801,N_1914);
and U3008 (N_3008,In_4478,N_327);
nor U3009 (N_3009,N_76,In_171);
nor U3010 (N_3010,N_396,In_2767);
or U3011 (N_3011,N_1395,N_1832);
nor U3012 (N_3012,In_3672,N_707);
and U3013 (N_3013,N_134,N_1085);
nand U3014 (N_3014,N_1591,N_828);
and U3015 (N_3015,N_1238,N_470);
nor U3016 (N_3016,In_3525,N_1744);
and U3017 (N_3017,N_1711,N_395);
or U3018 (N_3018,N_992,N_539);
or U3019 (N_3019,In_2755,In_3723);
xor U3020 (N_3020,N_1892,N_236);
nor U3021 (N_3021,N_658,N_942);
xor U3022 (N_3022,N_1155,N_666);
xnor U3023 (N_3023,N_1693,In_3966);
or U3024 (N_3024,In_1114,N_281);
nor U3025 (N_3025,In_967,N_858);
xnor U3026 (N_3026,N_1872,N_245);
nor U3027 (N_3027,N_1752,In_3481);
xor U3028 (N_3028,N_183,N_1202);
nor U3029 (N_3029,In_3612,N_1188);
or U3030 (N_3030,N_1316,In_89);
and U3031 (N_3031,N_1320,In_2430);
nor U3032 (N_3032,N_778,N_1512);
xnor U3033 (N_3033,N_1771,N_16);
nor U3034 (N_3034,N_143,In_1674);
and U3035 (N_3035,In_4009,In_4906);
or U3036 (N_3036,N_1466,N_496);
nor U3037 (N_3037,N_388,N_659);
nand U3038 (N_3038,N_214,N_492);
nor U3039 (N_3039,N_320,In_4190);
nor U3040 (N_3040,In_4124,N_427);
nand U3041 (N_3041,N_939,N_999);
and U3042 (N_3042,N_424,In_4330);
or U3043 (N_3043,N_244,N_1001);
nor U3044 (N_3044,N_1795,N_408);
and U3045 (N_3045,N_865,In_4078);
xor U3046 (N_3046,N_546,In_2252);
xor U3047 (N_3047,In_4138,N_1419);
xnor U3048 (N_3048,N_561,N_1702);
and U3049 (N_3049,N_809,N_1147);
xnor U3050 (N_3050,N_1878,N_1741);
or U3051 (N_3051,N_1152,N_446);
nor U3052 (N_3052,N_104,In_1847);
nor U3053 (N_3053,N_1095,N_1581);
nor U3054 (N_3054,N_182,N_1039);
xor U3055 (N_3055,N_1901,N_415);
nor U3056 (N_3056,In_2839,N_372);
nand U3057 (N_3057,N_1366,N_1968);
nand U3058 (N_3058,In_3326,N_744);
or U3059 (N_3059,N_414,N_922);
or U3060 (N_3060,In_4474,N_340);
or U3061 (N_3061,N_1372,N_518);
or U3062 (N_3062,In_2135,N_1875);
or U3063 (N_3063,N_307,N_553);
xor U3064 (N_3064,N_362,N_1613);
and U3065 (N_3065,N_260,N_1179);
nor U3066 (N_3066,N_703,In_4047);
and U3067 (N_3067,N_1182,In_824);
nor U3068 (N_3068,N_423,N_130);
and U3069 (N_3069,N_151,N_277);
xor U3070 (N_3070,In_780,N_1483);
nand U3071 (N_3071,N_223,N_1908);
nor U3072 (N_3072,N_267,N_83);
xnor U3073 (N_3073,In_143,N_1485);
nor U3074 (N_3074,N_1640,N_536);
nand U3075 (N_3075,N_1481,N_138);
nor U3076 (N_3076,In_1838,N_4);
xnor U3077 (N_3077,In_305,In_2154);
nor U3078 (N_3078,N_1224,N_1537);
or U3079 (N_3079,In_886,N_1972);
nand U3080 (N_3080,In_2093,In_1609);
nand U3081 (N_3081,N_610,N_1531);
and U3082 (N_3082,In_2859,In_3977);
and U3083 (N_3083,N_1442,In_1656);
or U3084 (N_3084,N_393,N_991);
nor U3085 (N_3085,In_4095,N_1653);
and U3086 (N_3086,N_974,In_1402);
nand U3087 (N_3087,N_1982,N_70);
and U3088 (N_3088,In_1528,In_1763);
nand U3089 (N_3089,N_1845,N_742);
and U3090 (N_3090,N_627,N_1277);
nor U3091 (N_3091,In_1873,In_2362);
and U3092 (N_3092,N_18,N_1765);
nor U3093 (N_3093,In_436,N_1661);
nor U3094 (N_3094,N_1758,In_182);
or U3095 (N_3095,N_235,In_4629);
and U3096 (N_3096,N_841,N_1231);
and U3097 (N_3097,In_364,N_1116);
nor U3098 (N_3098,N_1142,N_1478);
nor U3099 (N_3099,N_1964,N_886);
and U3100 (N_3100,N_1943,N_381);
nor U3101 (N_3101,In_4814,N_1911);
nand U3102 (N_3102,N_1918,In_3763);
nand U3103 (N_3103,N_1827,N_875);
and U3104 (N_3104,N_804,N_628);
nand U3105 (N_3105,In_2133,N_1444);
and U3106 (N_3106,In_2972,In_675);
xor U3107 (N_3107,In_1659,N_35);
or U3108 (N_3108,In_1897,N_1026);
nand U3109 (N_3109,In_1536,In_4337);
nand U3110 (N_3110,N_378,N_1947);
or U3111 (N_3111,N_1266,N_817);
and U3112 (N_3112,In_3383,N_1841);
xnor U3113 (N_3113,N_581,N_773);
xor U3114 (N_3114,N_1443,N_1730);
nor U3115 (N_3115,N_854,N_613);
nor U3116 (N_3116,In_517,In_4626);
nand U3117 (N_3117,N_1684,In_170);
nor U3118 (N_3118,In_4166,N_1807);
xnor U3119 (N_3119,N_1351,N_835);
xor U3120 (N_3120,N_1600,N_1580);
xor U3121 (N_3121,In_682,N_74);
and U3122 (N_3122,N_762,N_315);
nand U3123 (N_3123,In_155,N_621);
nor U3124 (N_3124,In_4919,N_933);
or U3125 (N_3125,N_1074,In_1337);
or U3126 (N_3126,N_603,In_4966);
nor U3127 (N_3127,N_1534,N_1853);
and U3128 (N_3128,In_1232,In_2049);
nor U3129 (N_3129,N_644,N_1674);
xor U3130 (N_3130,In_615,N_131);
xnor U3131 (N_3131,N_832,N_472);
nor U3132 (N_3132,N_930,N_1716);
nor U3133 (N_3133,N_441,In_4412);
or U3134 (N_3134,In_1666,N_1837);
nor U3135 (N_3135,N_1538,N_636);
or U3136 (N_3136,In_2496,N_1770);
nand U3137 (N_3137,N_1146,In_4155);
nand U3138 (N_3138,N_1654,N_1305);
or U3139 (N_3139,N_918,N_1920);
nor U3140 (N_3140,N_1099,In_271);
xor U3141 (N_3141,N_1709,In_747);
nand U3142 (N_3142,N_1889,N_211);
xnor U3143 (N_3143,N_1642,N_652);
nand U3144 (N_3144,N_306,In_2920);
xnor U3145 (N_3145,N_1550,N_1589);
xor U3146 (N_3146,N_1913,N_1341);
or U3147 (N_3147,N_678,In_1267);
nand U3148 (N_3148,N_456,In_3379);
xor U3149 (N_3149,In_2313,N_39);
nor U3150 (N_3150,N_1821,N_1722);
nand U3151 (N_3151,In_2453,N_174);
xnor U3152 (N_3152,In_1249,In_4237);
nand U3153 (N_3153,In_1088,N_7);
xor U3154 (N_3154,N_1997,N_1814);
and U3155 (N_3155,N_457,N_361);
xor U3156 (N_3156,N_787,N_1941);
nor U3157 (N_3157,N_1368,In_1185);
nor U3158 (N_3158,N_385,N_1347);
nand U3159 (N_3159,In_3487,N_1000);
or U3160 (N_3160,N_1701,N_278);
and U3161 (N_3161,In_943,In_4817);
xnor U3162 (N_3162,N_555,In_4110);
and U3163 (N_3163,N_198,N_993);
xor U3164 (N_3164,N_335,N_515);
or U3165 (N_3165,N_1161,N_1361);
or U3166 (N_3166,In_108,In_4010);
nor U3167 (N_3167,In_4892,N_186);
or U3168 (N_3168,N_1115,N_887);
and U3169 (N_3169,In_513,N_111);
xor U3170 (N_3170,In_1226,N_1260);
xor U3171 (N_3171,N_1697,N_866);
nand U3172 (N_3172,N_1127,N_359);
nor U3173 (N_3173,N_542,In_4402);
nand U3174 (N_3174,N_1662,N_1724);
nand U3175 (N_3175,N_623,In_131);
nor U3176 (N_3176,N_1014,N_1246);
nand U3177 (N_3177,In_858,In_3784);
or U3178 (N_3178,In_1474,N_1705);
and U3179 (N_3179,N_53,N_1232);
xnor U3180 (N_3180,In_2403,In_4921);
and U3181 (N_3181,N_802,N_162);
or U3182 (N_3182,In_1490,In_3125);
nand U3183 (N_3183,N_920,In_1140);
and U3184 (N_3184,N_1905,N_1128);
and U3185 (N_3185,In_4397,In_1145);
nand U3186 (N_3186,N_300,N_1506);
xnor U3187 (N_3187,N_1222,N_941);
and U3188 (N_3188,N_450,In_4805);
nand U3189 (N_3189,N_129,In_3997);
or U3190 (N_3190,N_971,N_85);
nor U3191 (N_3191,In_1939,In_4481);
nor U3192 (N_3192,In_2933,N_215);
or U3193 (N_3193,N_921,N_519);
xor U3194 (N_3194,N_860,N_356);
nand U3195 (N_3195,N_775,N_511);
or U3196 (N_3196,In_4276,N_1008);
and U3197 (N_3197,In_2665,In_1982);
nand U3198 (N_3198,N_1979,N_1069);
or U3199 (N_3199,N_303,N_1533);
or U3200 (N_3200,In_3018,In_1308);
xnor U3201 (N_3201,N_532,In_304);
nor U3202 (N_3202,In_69,N_1036);
nand U3203 (N_3203,In_3034,In_190);
nand U3204 (N_3204,N_1455,N_729);
nor U3205 (N_3205,N_179,N_656);
nor U3206 (N_3206,N_1201,N_1663);
nor U3207 (N_3207,In_3833,In_4233);
xnor U3208 (N_3208,N_801,In_1251);
nor U3209 (N_3209,N_1078,N_1989);
and U3210 (N_3210,N_1233,In_3588);
or U3211 (N_3211,N_1779,In_296);
nand U3212 (N_3212,N_325,In_895);
or U3213 (N_3213,N_1449,N_1646);
xor U3214 (N_3214,N_1754,N_1108);
nand U3215 (N_3215,N_1396,N_1772);
nand U3216 (N_3216,In_1366,N_478);
xnor U3217 (N_3217,N_105,In_1483);
and U3218 (N_3218,N_1826,N_1757);
and U3219 (N_3219,N_1063,N_825);
xor U3220 (N_3220,N_1946,In_3825);
nand U3221 (N_3221,N_342,In_2378);
xnor U3222 (N_3222,N_1579,N_1013);
or U3223 (N_3223,N_504,N_391);
or U3224 (N_3224,N_1606,In_500);
xnor U3225 (N_3225,In_435,In_2297);
nand U3226 (N_3226,In_4859,N_1031);
xnor U3227 (N_3227,N_108,In_169);
xnor U3228 (N_3228,In_3259,N_1562);
nand U3229 (N_3229,In_852,N_1859);
xor U3230 (N_3230,N_1317,N_107);
xnor U3231 (N_3231,In_813,N_1304);
nor U3232 (N_3232,In_673,In_4056);
xnor U3233 (N_3233,N_987,N_1489);
or U3234 (N_3234,N_1970,N_1975);
or U3235 (N_3235,N_1336,In_3832);
nor U3236 (N_3236,N_1742,In_1633);
nor U3237 (N_3237,N_964,N_1886);
nor U3238 (N_3238,In_1093,N_295);
nor U3239 (N_3239,N_1887,N_449);
and U3240 (N_3240,N_1794,In_1012);
nor U3241 (N_3241,N_853,N_573);
nand U3242 (N_3242,N_647,In_2263);
or U3243 (N_3243,In_4849,N_1816);
and U3244 (N_3244,In_3227,N_913);
and U3245 (N_3245,N_270,In_3411);
nand U3246 (N_3246,N_193,N_593);
and U3247 (N_3247,N_296,In_2654);
and U3248 (N_3248,N_419,In_3298);
xnor U3249 (N_3249,N_1861,In_1163);
and U3250 (N_3250,In_2731,N_256);
and U3251 (N_3251,N_1871,N_309);
or U3252 (N_3252,N_1704,In_889);
nor U3253 (N_3253,In_3082,N_1075);
or U3254 (N_3254,N_1900,N_9);
nor U3255 (N_3255,N_900,In_4011);
nor U3256 (N_3256,N_948,N_501);
nor U3257 (N_3257,N_799,In_3952);
nor U3258 (N_3258,N_58,In_801);
and U3259 (N_3259,N_777,N_1102);
nand U3260 (N_3260,N_852,N_914);
nand U3261 (N_3261,N_1104,N_1400);
nor U3262 (N_3262,N_1508,N_443);
nand U3263 (N_3263,In_2743,N_199);
or U3264 (N_3264,N_507,In_309);
nor U3265 (N_3265,N_1145,N_572);
or U3266 (N_3266,In_1906,In_3682);
or U3267 (N_3267,In_4674,In_2495);
nand U3268 (N_3268,In_3602,N_141);
and U3269 (N_3269,In_1261,N_1789);
nor U3270 (N_3270,In_2953,N_739);
nor U3271 (N_3271,N_50,In_4042);
or U3272 (N_3272,N_24,In_3688);
nor U3273 (N_3273,N_513,N_352);
or U3274 (N_3274,In_3249,N_476);
and U3275 (N_3275,In_1069,N_1995);
or U3276 (N_3276,N_1406,In_1830);
xnor U3277 (N_3277,In_4672,In_1322);
and U3278 (N_3278,N_1940,In_4113);
and U3279 (N_3279,N_1071,N_1118);
nor U3280 (N_3280,N_177,N_1245);
or U3281 (N_3281,N_1474,N_213);
or U3282 (N_3282,N_1154,N_1812);
nor U3283 (N_3283,In_627,N_945);
xor U3284 (N_3284,N_403,N_793);
xor U3285 (N_3285,N_640,In_635);
nand U3286 (N_3286,N_894,N_1996);
xnor U3287 (N_3287,In_2117,N_783);
nand U3288 (N_3288,In_2702,N_310);
nor U3289 (N_3289,In_3332,In_429);
or U3290 (N_3290,N_698,N_722);
or U3291 (N_3291,N_1093,N_48);
nand U3292 (N_3292,In_4115,N_1519);
and U3293 (N_3293,N_1420,N_679);
nor U3294 (N_3294,In_3347,N_1195);
or U3295 (N_3295,N_1264,In_1857);
nand U3296 (N_3296,N_234,In_3493);
nor U3297 (N_3297,In_4690,N_1571);
or U3298 (N_3298,N_629,N_219);
nand U3299 (N_3299,N_893,N_1345);
xor U3300 (N_3300,N_1389,In_381);
or U3301 (N_3301,N_1307,N_1226);
and U3302 (N_3302,N_1629,N_1130);
xor U3303 (N_3303,N_929,N_1236);
and U3304 (N_3304,In_2165,N_434);
xor U3305 (N_3305,N_1439,N_1337);
nand U3306 (N_3306,N_1846,N_1299);
xnor U3307 (N_3307,N_950,In_2054);
nor U3308 (N_3308,N_1961,N_521);
nor U3309 (N_3309,In_2629,In_4793);
nand U3310 (N_3310,N_878,N_1428);
nor U3311 (N_3311,N_128,In_4719);
and U3312 (N_3312,N_923,N_996);
and U3313 (N_3313,N_431,N_1363);
or U3314 (N_3314,N_1524,N_1035);
or U3315 (N_3315,N_347,N_1690);
xor U3316 (N_3316,In_2157,N_1944);
and U3317 (N_3317,N_795,N_1429);
nand U3318 (N_3318,In_2632,N_1284);
and U3319 (N_3319,N_1612,In_4976);
or U3320 (N_3320,N_1452,N_1803);
nand U3321 (N_3321,N_626,N_1294);
nor U3322 (N_3322,N_1738,N_1852);
and U3323 (N_3323,In_540,N_907);
nand U3324 (N_3324,In_2273,In_3197);
nand U3325 (N_3325,In_648,N_154);
nand U3326 (N_3326,N_1086,In_3090);
and U3327 (N_3327,N_699,N_1367);
nor U3328 (N_3328,In_3219,N_401);
nand U3329 (N_3329,In_3741,N_1649);
or U3330 (N_3330,N_1379,In_2202);
nand U3331 (N_3331,N_1713,N_232);
nand U3332 (N_3332,N_761,N_1315);
or U3333 (N_3333,N_1017,In_3231);
nand U3334 (N_3334,In_4908,N_1422);
nand U3335 (N_3335,N_800,N_1051);
and U3336 (N_3336,N_1542,N_1675);
nor U3337 (N_3337,N_1556,N_535);
nor U3338 (N_3338,In_3855,N_1196);
xnor U3339 (N_3339,N_899,In_594);
or U3340 (N_3340,N_287,In_4246);
nor U3341 (N_3341,N_477,N_1945);
or U3342 (N_3342,N_1558,N_1469);
nor U3343 (N_3343,N_1470,N_286);
and U3344 (N_3344,N_490,In_2448);
nor U3345 (N_3345,In_977,N_1776);
and U3346 (N_3346,N_1552,In_1540);
and U3347 (N_3347,N_38,N_49);
nor U3348 (N_3348,N_1949,In_1266);
and U3349 (N_3349,N_1599,N_861);
and U3350 (N_3350,In_3157,N_591);
xor U3351 (N_3351,N_1689,In_1606);
and U3352 (N_3352,N_1167,In_141);
and U3353 (N_3353,N_1521,N_1144);
or U3354 (N_3354,In_660,In_625);
xor U3355 (N_3355,In_2650,N_264);
xnor U3356 (N_3356,N_1373,N_1137);
or U3357 (N_3357,In_1104,N_1535);
and U3358 (N_3358,N_796,N_387);
and U3359 (N_3359,In_554,N_1658);
and U3360 (N_3360,In_3196,N_314);
and U3361 (N_3361,N_1267,In_107);
xnor U3362 (N_3362,N_749,In_2547);
xnor U3363 (N_3363,In_2815,In_3295);
xnor U3364 (N_3364,In_1619,In_4983);
nand U3365 (N_3365,N_1678,N_41);
or U3366 (N_3366,In_2651,N_845);
nand U3367 (N_3367,In_96,N_10);
and U3368 (N_3368,N_365,In_715);
or U3369 (N_3369,In_3801,N_34);
nand U3370 (N_3370,N_646,N_27);
xnor U3371 (N_3371,N_565,In_1740);
nor U3372 (N_3372,N_1505,In_862);
nand U3373 (N_3373,N_1735,N_1050);
or U3374 (N_3374,N_1839,N_1876);
nand U3375 (N_3375,N_1844,In_551);
and U3376 (N_3376,In_3988,In_3316);
or U3377 (N_3377,N_1391,N_1959);
nand U3378 (N_3378,In_4297,In_2939);
and U3379 (N_3379,N_126,N_1694);
xnor U3380 (N_3380,N_2,N_534);
xor U3381 (N_3381,N_1159,N_912);
or U3382 (N_3382,N_291,N_412);
nand U3383 (N_3383,In_571,In_4443);
nor U3384 (N_3384,In_216,N_1030);
nor U3385 (N_3385,In_4925,N_608);
nand U3386 (N_3386,N_370,N_66);
nor U3387 (N_3387,N_117,In_560);
and U3388 (N_3388,N_735,In_2286);
xnor U3389 (N_3389,N_172,N_836);
or U3390 (N_3390,In_4755,N_1627);
xor U3391 (N_3391,N_639,N_574);
and U3392 (N_3392,N_187,In_3592);
and U3393 (N_3393,N_262,In_2451);
xnor U3394 (N_3394,N_1715,N_473);
xnor U3395 (N_3395,N_1414,In_2436);
and U3396 (N_3396,N_69,N_123);
nand U3397 (N_3397,N_1575,N_1033);
or U3398 (N_3398,N_946,N_657);
or U3399 (N_3399,N_876,N_577);
nor U3400 (N_3400,N_168,In_812);
xor U3401 (N_3401,N_345,N_158);
and U3402 (N_3402,N_1047,N_552);
xnor U3403 (N_3403,N_1059,N_437);
or U3404 (N_3404,N_1725,In_581);
xnor U3405 (N_3405,N_816,In_2846);
or U3406 (N_3406,N_1356,N_1883);
and U3407 (N_3407,N_299,N_924);
or U3408 (N_3408,N_461,N_282);
or U3409 (N_3409,In_77,In_2824);
or U3410 (N_3410,In_1311,In_1951);
nor U3411 (N_3411,N_20,N_116);
nor U3412 (N_3412,N_695,N_1135);
and U3413 (N_3413,N_1313,N_218);
or U3414 (N_3414,N_1306,N_1323);
and U3415 (N_3415,N_326,N_1667);
and U3416 (N_3416,In_4501,N_1479);
nor U3417 (N_3417,In_20,N_1721);
or U3418 (N_3418,In_491,In_1099);
and U3419 (N_3419,In_882,N_1206);
nand U3420 (N_3420,N_1234,N_1184);
nand U3421 (N_3421,N_633,N_1369);
or U3422 (N_3422,N_1375,In_2186);
nand U3423 (N_3423,N_682,N_763);
nand U3424 (N_3424,N_31,N_1383);
nand U3425 (N_3425,N_1651,N_1021);
xnor U3426 (N_3426,N_1623,N_664);
and U3427 (N_3427,N_429,N_537);
and U3428 (N_3428,N_953,N_1454);
and U3429 (N_3429,In_3182,In_2519);
or U3430 (N_3430,N_1673,In_1792);
xor U3431 (N_3431,N_1978,N_171);
or U3432 (N_3432,N_1934,In_2150);
xor U3433 (N_3433,N_1281,In_1497);
xnor U3434 (N_3434,N_1215,N_916);
or U3435 (N_3435,N_961,N_648);
nand U3436 (N_3436,In_3705,N_459);
or U3437 (N_3437,N_1990,N_1139);
xnor U3438 (N_3438,N_228,N_1197);
xor U3439 (N_3439,N_276,N_113);
and U3440 (N_3440,N_180,In_2481);
nand U3441 (N_3441,N_1235,N_1625);
nor U3442 (N_3442,N_1659,N_620);
xor U3443 (N_3443,In_1685,N_397);
or U3444 (N_3444,N_1793,N_1472);
nor U3445 (N_3445,N_966,N_1601);
nor U3446 (N_3446,N_788,N_1799);
nand U3447 (N_3447,N_1430,N_1593);
nor U3448 (N_3448,N_790,In_2170);
or U3449 (N_3449,In_3900,N_1810);
nor U3450 (N_3450,N_771,In_2644);
xnor U3451 (N_3451,N_485,N_248);
xor U3452 (N_3452,N_583,N_1517);
and U3453 (N_3453,N_502,N_892);
nand U3454 (N_3454,N_1176,N_1753);
or U3455 (N_3455,In_4182,In_2916);
xnor U3456 (N_3456,In_1457,In_3309);
and U3457 (N_3457,In_185,N_859);
and U3458 (N_3458,In_2357,N_1525);
and U3459 (N_3459,In_867,In_4151);
or U3460 (N_3460,In_475,N_1957);
nor U3461 (N_3461,In_1438,In_4065);
nor U3462 (N_3462,N_1087,N_222);
xnor U3463 (N_3463,N_677,In_3330);
nand U3464 (N_3464,N_785,N_794);
nand U3465 (N_3465,N_1397,N_1815);
xnor U3466 (N_3466,N_229,In_3472);
nand U3467 (N_3467,In_1686,In_2476);
or U3468 (N_3468,N_1364,In_1845);
nand U3469 (N_3469,N_266,In_3417);
nor U3470 (N_3470,N_44,In_1476);
or U3471 (N_3471,N_1767,N_1471);
nor U3472 (N_3472,N_1440,In_3242);
nor U3473 (N_3473,In_3001,In_4959);
or U3474 (N_3474,N_1585,In_2732);
or U3475 (N_3475,In_3806,N_1818);
nor U3476 (N_3476,In_4792,In_3340);
or U3477 (N_3477,N_1314,In_3405);
nor U3478 (N_3478,In_3272,N_65);
nand U3479 (N_3479,N_1090,In_4140);
or U3480 (N_3480,N_1203,In_2103);
nand U3481 (N_3481,N_258,In_14);
nand U3482 (N_3482,In_2456,N_595);
nor U3483 (N_3483,N_435,N_1061);
nor U3484 (N_3484,N_426,N_1143);
nand U3485 (N_3485,N_12,N_32);
nor U3486 (N_3486,In_4392,In_1622);
nand U3487 (N_3487,In_2294,In_4222);
or U3488 (N_3488,In_2642,In_863);
and U3489 (N_3489,In_2762,In_762);
xnor U3490 (N_3490,N_1382,In_470);
nand U3491 (N_3491,In_329,In_3597);
xnor U3492 (N_3492,In_2014,In_211);
nor U3493 (N_3493,N_1424,In_539);
xnor U3494 (N_3494,In_2087,N_1984);
or U3495 (N_3495,N_1038,N_1608);
xnor U3496 (N_3496,N_251,N_346);
xnor U3497 (N_3497,In_2410,In_3395);
nor U3498 (N_3498,In_1103,N_976);
or U3499 (N_3499,N_662,In_3488);
or U3500 (N_3500,N_1579,In_2654);
and U3501 (N_3501,N_787,N_1471);
nand U3502 (N_3502,N_374,N_275);
and U3503 (N_3503,N_1447,In_251);
xnor U3504 (N_3504,In_4271,N_1336);
nand U3505 (N_3505,N_176,In_3187);
or U3506 (N_3506,N_1787,N_1300);
or U3507 (N_3507,In_4598,N_1283);
and U3508 (N_3508,N_1897,In_1687);
xor U3509 (N_3509,N_1555,N_1459);
xor U3510 (N_3510,N_1077,N_688);
xor U3511 (N_3511,N_1109,N_816);
nand U3512 (N_3512,In_351,N_845);
or U3513 (N_3513,N_1132,N_1544);
xnor U3514 (N_3514,N_870,N_1296);
or U3515 (N_3515,N_645,N_335);
xnor U3516 (N_3516,In_1775,N_1114);
nand U3517 (N_3517,N_449,N_1397);
xnor U3518 (N_3518,N_132,N_585);
or U3519 (N_3519,N_1569,N_1599);
xor U3520 (N_3520,In_768,In_3124);
nand U3521 (N_3521,N_1405,In_855);
and U3522 (N_3522,N_1186,N_1553);
and U3523 (N_3523,In_3091,N_257);
xor U3524 (N_3524,N_118,In_2535);
and U3525 (N_3525,N_158,N_862);
nor U3526 (N_3526,N_716,In_3840);
nand U3527 (N_3527,N_1045,N_1856);
nor U3528 (N_3528,N_847,N_1131);
nand U3529 (N_3529,N_1616,N_1945);
or U3530 (N_3530,N_1383,In_42);
or U3531 (N_3531,In_4095,In_669);
or U3532 (N_3532,N_1628,In_2732);
nor U3533 (N_3533,N_1320,N_662);
or U3534 (N_3534,N_1069,N_1699);
or U3535 (N_3535,N_614,N_269);
and U3536 (N_3536,In_4598,In_3209);
and U3537 (N_3537,N_942,N_1030);
nor U3538 (N_3538,In_3036,N_1427);
nand U3539 (N_3539,In_1250,In_4010);
nand U3540 (N_3540,N_839,N_1592);
or U3541 (N_3541,In_2313,N_845);
nand U3542 (N_3542,N_881,N_1599);
nor U3543 (N_3543,N_1917,In_2632);
or U3544 (N_3544,N_367,N_1589);
xnor U3545 (N_3545,In_3197,In_98);
nand U3546 (N_3546,N_80,In_1540);
nand U3547 (N_3547,In_3639,In_3435);
or U3548 (N_3548,N_226,N_803);
xnor U3549 (N_3549,In_169,N_152);
xor U3550 (N_3550,N_641,In_3174);
nand U3551 (N_3551,In_4481,In_3212);
and U3552 (N_3552,In_1112,In_3399);
or U3553 (N_3553,N_1705,In_3904);
nor U3554 (N_3554,N_1181,N_649);
or U3555 (N_3555,N_779,N_1057);
xor U3556 (N_3556,N_471,N_1459);
or U3557 (N_3557,In_418,N_172);
xnor U3558 (N_3558,N_478,In_3551);
nor U3559 (N_3559,In_2613,In_1659);
xnor U3560 (N_3560,In_3347,N_782);
xnor U3561 (N_3561,N_820,In_4095);
and U3562 (N_3562,In_3395,N_42);
nand U3563 (N_3563,N_1644,In_805);
or U3564 (N_3564,N_1438,In_2533);
or U3565 (N_3565,N_1850,N_1493);
and U3566 (N_3566,N_592,N_1092);
nor U3567 (N_3567,N_1567,N_472);
xor U3568 (N_3568,In_209,In_4560);
and U3569 (N_3569,In_2533,In_4018);
or U3570 (N_3570,N_1493,N_1016);
nand U3571 (N_3571,N_871,N_1461);
or U3572 (N_3572,N_659,In_2291);
xor U3573 (N_3573,N_1355,In_1490);
nor U3574 (N_3574,In_345,N_1554);
and U3575 (N_3575,N_387,N_1465);
and U3576 (N_3576,N_345,In_1763);
xor U3577 (N_3577,N_880,N_256);
nand U3578 (N_3578,In_282,In_1522);
or U3579 (N_3579,N_772,In_3340);
xnor U3580 (N_3580,N_1906,N_260);
nor U3581 (N_3581,In_132,In_4397);
nor U3582 (N_3582,N_1443,N_443);
or U3583 (N_3583,In_4898,N_1146);
and U3584 (N_3584,N_1088,N_483);
nand U3585 (N_3585,N_953,In_4047);
xor U3586 (N_3586,In_3758,N_1893);
nor U3587 (N_3587,In_1933,N_1554);
nor U3588 (N_3588,N_699,In_517);
nand U3589 (N_3589,In_863,N_1581);
and U3590 (N_3590,In_3157,N_885);
and U3591 (N_3591,N_210,In_1383);
xor U3592 (N_3592,N_1921,In_4849);
and U3593 (N_3593,In_4690,N_708);
or U3594 (N_3594,In_2820,N_1422);
or U3595 (N_3595,In_96,In_2615);
or U3596 (N_3596,In_2755,In_4366);
and U3597 (N_3597,N_1659,In_1830);
xor U3598 (N_3598,In_4151,N_712);
xnor U3599 (N_3599,N_1167,N_1315);
nand U3600 (N_3600,In_3253,In_2982);
nor U3601 (N_3601,N_1477,N_108);
nand U3602 (N_3602,N_1408,In_69);
or U3603 (N_3603,In_1329,N_175);
and U3604 (N_3604,In_1536,N_76);
or U3605 (N_3605,N_318,In_345);
or U3606 (N_3606,N_1643,In_2815);
xnor U3607 (N_3607,N_872,N_748);
or U3608 (N_3608,In_3588,In_3736);
and U3609 (N_3609,In_1845,N_475);
xor U3610 (N_3610,N_1749,N_1798);
nand U3611 (N_3611,N_1917,N_1260);
nand U3612 (N_3612,In_1,In_4532);
nor U3613 (N_3613,In_4195,In_4966);
nand U3614 (N_3614,N_1180,N_1087);
or U3615 (N_3615,N_1134,In_3326);
nand U3616 (N_3616,N_1701,In_2650);
and U3617 (N_3617,N_1158,N_1755);
nand U3618 (N_3618,N_678,In_4478);
xor U3619 (N_3619,In_74,N_206);
nand U3620 (N_3620,N_319,N_1105);
xnor U3621 (N_3621,In_4017,N_885);
nand U3622 (N_3622,N_1061,N_394);
nor U3623 (N_3623,N_147,N_945);
nor U3624 (N_3624,N_1514,In_1944);
xnor U3625 (N_3625,N_1584,In_3313);
and U3626 (N_3626,N_30,In_762);
xnor U3627 (N_3627,N_2,In_3488);
xor U3628 (N_3628,N_358,In_3973);
nor U3629 (N_3629,N_1589,N_1840);
and U3630 (N_3630,N_1822,N_1184);
or U3631 (N_3631,In_4392,In_2642);
and U3632 (N_3632,N_1263,N_1830);
nand U3633 (N_3633,N_137,N_724);
xnor U3634 (N_3634,In_31,In_3088);
or U3635 (N_3635,N_1621,In_4124);
or U3636 (N_3636,N_1736,N_770);
xnor U3637 (N_3637,N_947,N_483);
and U3638 (N_3638,N_510,N_1635);
nand U3639 (N_3639,N_1268,N_1682);
nand U3640 (N_3640,N_1064,N_1865);
and U3641 (N_3641,N_1071,N_1927);
xnor U3642 (N_3642,N_348,N_1093);
nor U3643 (N_3643,N_1441,N_1613);
and U3644 (N_3644,N_1614,N_173);
nor U3645 (N_3645,N_1560,N_1363);
or U3646 (N_3646,N_1269,N_178);
or U3647 (N_3647,In_2535,In_3336);
and U3648 (N_3648,N_824,In_4467);
xnor U3649 (N_3649,In_2157,N_1586);
nand U3650 (N_3650,In_2629,N_240);
nand U3651 (N_3651,In_351,N_1413);
nor U3652 (N_3652,N_700,In_2188);
and U3653 (N_3653,N_1143,N_1091);
and U3654 (N_3654,N_388,In_4906);
or U3655 (N_3655,N_1484,N_1953);
xor U3656 (N_3656,In_3949,N_258);
or U3657 (N_3657,In_4262,N_121);
nor U3658 (N_3658,In_1740,N_694);
nand U3659 (N_3659,In_4706,N_1539);
nor U3660 (N_3660,N_220,N_239);
and U3661 (N_3661,N_1328,N_1272);
or U3662 (N_3662,N_1054,In_3477);
nor U3663 (N_3663,N_1329,N_1397);
or U3664 (N_3664,N_1735,N_925);
or U3665 (N_3665,N_789,N_1850);
nand U3666 (N_3666,In_2979,N_1402);
nand U3667 (N_3667,N_1990,N_56);
xor U3668 (N_3668,N_371,N_833);
nand U3669 (N_3669,N_226,N_371);
or U3670 (N_3670,N_1760,In_2535);
nor U3671 (N_3671,N_407,N_1716);
and U3672 (N_3672,N_1422,N_1498);
or U3673 (N_3673,N_691,N_1152);
xor U3674 (N_3674,N_958,N_1646);
nor U3675 (N_3675,In_479,N_590);
nor U3676 (N_3676,In_2616,N_1569);
or U3677 (N_3677,In_3855,N_526);
or U3678 (N_3678,N_1305,N_934);
nand U3679 (N_3679,N_1563,In_1792);
xnor U3680 (N_3680,N_1254,N_1807);
or U3681 (N_3681,In_4078,N_438);
and U3682 (N_3682,N_1288,In_610);
and U3683 (N_3683,In_1019,In_953);
and U3684 (N_3684,In_3294,In_3215);
and U3685 (N_3685,In_171,In_949);
nand U3686 (N_3686,N_429,In_4938);
nand U3687 (N_3687,N_340,N_1462);
nand U3688 (N_3688,In_2074,N_913);
xnor U3689 (N_3689,In_1093,N_196);
nand U3690 (N_3690,N_1326,N_1302);
or U3691 (N_3691,In_1933,N_1992);
or U3692 (N_3692,N_628,In_2088);
xor U3693 (N_3693,N_1115,In_3096);
and U3694 (N_3694,In_2088,N_1337);
or U3695 (N_3695,In_813,In_3738);
or U3696 (N_3696,N_1519,In_1241);
nor U3697 (N_3697,N_1474,N_422);
xor U3698 (N_3698,In_1023,N_421);
and U3699 (N_3699,N_1558,N_1679);
nor U3700 (N_3700,N_714,N_250);
nor U3701 (N_3701,In_2916,N_559);
nand U3702 (N_3702,N_141,N_1059);
xnor U3703 (N_3703,N_237,In_1675);
or U3704 (N_3704,N_161,In_2640);
and U3705 (N_3705,N_1724,N_1687);
xnor U3706 (N_3706,N_1492,N_1411);
nand U3707 (N_3707,N_1302,In_4044);
nor U3708 (N_3708,N_611,N_968);
and U3709 (N_3709,N_1858,In_2059);
or U3710 (N_3710,N_847,In_4439);
nand U3711 (N_3711,N_332,N_1306);
nor U3712 (N_3712,In_4004,In_4042);
xnor U3713 (N_3713,N_1770,N_1051);
nor U3714 (N_3714,In_3482,N_1070);
and U3715 (N_3715,N_1995,In_4849);
xor U3716 (N_3716,N_401,In_703);
xnor U3717 (N_3717,N_178,N_587);
xor U3718 (N_3718,N_1577,In_2446);
and U3719 (N_3719,In_3855,In_2113);
xor U3720 (N_3720,N_858,N_1157);
nand U3721 (N_3721,N_322,In_2727);
nand U3722 (N_3722,In_3420,N_8);
or U3723 (N_3723,N_1267,In_2979);
and U3724 (N_3724,In_1786,In_2988);
or U3725 (N_3725,N_1964,N_1617);
nand U3726 (N_3726,N_1045,N_654);
nand U3727 (N_3727,N_1463,In_4901);
or U3728 (N_3728,N_1243,In_4628);
nand U3729 (N_3729,N_1557,N_646);
xor U3730 (N_3730,In_354,N_611);
xnor U3731 (N_3731,N_1868,N_700);
nand U3732 (N_3732,In_2170,N_689);
nand U3733 (N_3733,In_1593,N_159);
xor U3734 (N_3734,N_347,N_247);
or U3735 (N_3735,In_2359,In_3334);
xor U3736 (N_3736,In_412,N_1395);
nand U3737 (N_3737,N_555,N_1335);
or U3738 (N_3738,N_803,N_1733);
and U3739 (N_3739,In_1461,N_327);
xor U3740 (N_3740,N_1394,In_4330);
nand U3741 (N_3741,N_95,N_1395);
xor U3742 (N_3742,In_2731,In_3272);
and U3743 (N_3743,In_3034,N_1477);
or U3744 (N_3744,N_1036,N_1621);
nor U3745 (N_3745,N_1184,N_942);
and U3746 (N_3746,N_216,In_3404);
or U3747 (N_3747,N_971,N_246);
nor U3748 (N_3748,N_1655,N_678);
xor U3749 (N_3749,N_354,In_2629);
nor U3750 (N_3750,N_1248,In_0);
nand U3751 (N_3751,N_1496,N_782);
and U3752 (N_3752,N_997,In_3383);
and U3753 (N_3753,In_2665,N_1704);
xnor U3754 (N_3754,In_3686,N_1162);
xor U3755 (N_3755,In_977,In_4927);
or U3756 (N_3756,N_206,N_1103);
or U3757 (N_3757,In_3602,In_1208);
or U3758 (N_3758,N_317,N_1741);
xor U3759 (N_3759,In_813,N_768);
xor U3760 (N_3760,N_772,N_139);
xnor U3761 (N_3761,N_705,N_258);
nand U3762 (N_3762,In_2642,N_77);
nor U3763 (N_3763,N_579,N_659);
nor U3764 (N_3764,N_100,N_346);
and U3765 (N_3765,In_4787,In_1792);
nor U3766 (N_3766,In_4844,N_174);
and U3767 (N_3767,N_1502,N_1247);
or U3768 (N_3768,In_4995,In_202);
xor U3769 (N_3769,N_1449,N_802);
and U3770 (N_3770,N_868,In_1208);
or U3771 (N_3771,N_1756,In_4618);
xnor U3772 (N_3772,N_1305,N_1416);
and U3773 (N_3773,N_988,N_1036);
nand U3774 (N_3774,In_3990,In_800);
and U3775 (N_3775,N_880,In_4937);
and U3776 (N_3776,N_587,N_1503);
xor U3777 (N_3777,N_336,N_1088);
nor U3778 (N_3778,In_2111,N_84);
or U3779 (N_3779,N_1610,In_2273);
nand U3780 (N_3780,N_429,N_1479);
or U3781 (N_3781,In_4718,N_1236);
nand U3782 (N_3782,N_1707,N_1693);
nand U3783 (N_3783,N_1787,N_1980);
or U3784 (N_3784,In_4627,N_722);
and U3785 (N_3785,In_562,N_805);
xnor U3786 (N_3786,N_1721,In_2779);
and U3787 (N_3787,N_956,In_4018);
xor U3788 (N_3788,In_2702,N_795);
xnor U3789 (N_3789,N_1101,N_880);
xnor U3790 (N_3790,N_688,N_790);
and U3791 (N_3791,N_84,N_1596);
nand U3792 (N_3792,N_1116,N_1513);
nand U3793 (N_3793,N_244,N_1126);
and U3794 (N_3794,N_1039,N_420);
xnor U3795 (N_3795,In_4556,N_1497);
nand U3796 (N_3796,In_1955,N_1845);
xnor U3797 (N_3797,N_1455,N_581);
nor U3798 (N_3798,N_972,N_986);
nor U3799 (N_3799,N_1753,N_237);
xnor U3800 (N_3800,N_1747,In_4439);
or U3801 (N_3801,N_1198,In_1972);
nand U3802 (N_3802,N_259,In_2644);
nand U3803 (N_3803,In_620,In_3187);
or U3804 (N_3804,In_1093,N_1233);
or U3805 (N_3805,N_1102,N_745);
and U3806 (N_3806,N_369,N_794);
nand U3807 (N_3807,N_225,In_873);
nor U3808 (N_3808,N_6,In_4690);
nor U3809 (N_3809,In_3825,N_971);
or U3810 (N_3810,In_4598,N_1288);
or U3811 (N_3811,N_850,In_4571);
xnor U3812 (N_3812,N_790,In_1195);
xor U3813 (N_3813,In_1939,N_119);
or U3814 (N_3814,N_892,In_2049);
nand U3815 (N_3815,N_1354,N_1776);
nor U3816 (N_3816,N_981,N_1605);
and U3817 (N_3817,N_1431,In_3209);
nor U3818 (N_3818,N_1152,N_1748);
xor U3819 (N_3819,N_1733,N_1172);
and U3820 (N_3820,In_2379,In_4316);
and U3821 (N_3821,In_2170,In_3612);
or U3822 (N_3822,N_1212,N_979);
or U3823 (N_3823,In_2273,In_2434);
and U3824 (N_3824,N_1397,N_35);
nand U3825 (N_3825,In_1917,N_1715);
xnor U3826 (N_3826,N_1286,N_1668);
nor U3827 (N_3827,N_1421,N_153);
nand U3828 (N_3828,N_283,N_37);
and U3829 (N_3829,N_607,In_1536);
and U3830 (N_3830,N_1499,In_443);
nor U3831 (N_3831,In_3248,N_1507);
xnor U3832 (N_3832,In_3074,In_3778);
nand U3833 (N_3833,In_3133,N_1626);
and U3834 (N_3834,N_635,N_354);
nand U3835 (N_3835,In_4044,In_1087);
xnor U3836 (N_3836,N_680,N_588);
xor U3837 (N_3837,N_1398,N_1692);
nor U3838 (N_3838,N_99,In_4686);
nand U3839 (N_3839,N_129,In_4237);
or U3840 (N_3840,N_1164,In_3514);
xnor U3841 (N_3841,In_4281,N_1848);
or U3842 (N_3842,N_1807,In_550);
or U3843 (N_3843,In_1854,N_459);
nand U3844 (N_3844,In_2306,N_1065);
nand U3845 (N_3845,N_1337,N_890);
nand U3846 (N_3846,N_1970,N_491);
xnor U3847 (N_3847,In_155,In_1661);
nor U3848 (N_3848,In_2616,N_1998);
and U3849 (N_3849,N_197,N_92);
nand U3850 (N_3850,N_1011,N_467);
and U3851 (N_3851,In_1658,N_1642);
or U3852 (N_3852,In_780,N_1646);
nand U3853 (N_3853,N_167,N_1548);
nor U3854 (N_3854,N_558,N_1686);
nor U3855 (N_3855,N_868,N_1878);
nand U3856 (N_3856,N_1381,N_899);
nor U3857 (N_3857,In_3612,N_1292);
nor U3858 (N_3858,In_3663,N_1546);
and U3859 (N_3859,N_1596,N_921);
nor U3860 (N_3860,In_1372,N_1781);
xor U3861 (N_3861,In_1765,N_1541);
and U3862 (N_3862,In_4068,N_370);
xnor U3863 (N_3863,N_70,N_1357);
xnor U3864 (N_3864,N_1947,N_109);
xor U3865 (N_3865,N_1044,In_4222);
xnor U3866 (N_3866,In_185,N_1223);
and U3867 (N_3867,In_3124,N_731);
or U3868 (N_3868,In_863,In_3609);
xnor U3869 (N_3869,N_113,N_412);
xor U3870 (N_3870,N_782,N_295);
nand U3871 (N_3871,In_3437,N_390);
xnor U3872 (N_3872,N_647,N_1780);
and U3873 (N_3873,N_1391,In_2991);
nor U3874 (N_3874,N_1396,N_1771);
nor U3875 (N_3875,N_1660,N_1171);
xnor U3876 (N_3876,N_230,In_479);
nor U3877 (N_3877,In_1446,N_475);
nor U3878 (N_3878,In_4439,In_3933);
or U3879 (N_3879,N_1130,N_580);
or U3880 (N_3880,N_353,N_999);
nor U3881 (N_3881,In_4054,In_627);
xnor U3882 (N_3882,N_1209,N_776);
nand U3883 (N_3883,In_1118,N_909);
xor U3884 (N_3884,N_1083,N_692);
and U3885 (N_3885,N_1115,N_745);
or U3886 (N_3886,In_550,In_4347);
nor U3887 (N_3887,N_141,N_1986);
xor U3888 (N_3888,N_1755,N_679);
or U3889 (N_3889,In_3215,N_1172);
or U3890 (N_3890,N_206,N_1123);
nor U3891 (N_3891,N_1464,N_703);
or U3892 (N_3892,In_3210,N_1261);
xor U3893 (N_3893,In_2088,N_844);
xnor U3894 (N_3894,In_936,N_1382);
nand U3895 (N_3895,N_1802,N_1097);
or U3896 (N_3896,In_1676,In_504);
nand U3897 (N_3897,N_1140,N_709);
and U3898 (N_3898,In_4331,N_1948);
nand U3899 (N_3899,N_33,In_1659);
and U3900 (N_3900,N_1165,N_519);
and U3901 (N_3901,N_143,N_1054);
xnor U3902 (N_3902,N_1291,In_2647);
or U3903 (N_3903,N_1340,N_1604);
nor U3904 (N_3904,In_2846,N_681);
or U3905 (N_3905,N_374,N_76);
nand U3906 (N_3906,N_626,N_996);
or U3907 (N_3907,In_996,N_511);
nor U3908 (N_3908,N_1172,In_4200);
or U3909 (N_3909,N_1089,N_1633);
xnor U3910 (N_3910,In_3149,N_1219);
and U3911 (N_3911,N_1431,N_580);
nor U3912 (N_3912,N_1733,In_4305);
xor U3913 (N_3913,In_2859,N_242);
nand U3914 (N_3914,N_1620,N_1301);
or U3915 (N_3915,In_3001,In_2651);
nand U3916 (N_3916,In_1572,In_2719);
nor U3917 (N_3917,In_858,N_987);
xnor U3918 (N_3918,N_6,In_1606);
or U3919 (N_3919,N_594,N_640);
nand U3920 (N_3920,In_2509,In_2859);
or U3921 (N_3921,In_4719,N_1848);
xor U3922 (N_3922,In_3018,N_781);
nand U3923 (N_3923,In_4365,N_174);
nor U3924 (N_3924,In_374,N_1388);
nand U3925 (N_3925,N_755,N_535);
nand U3926 (N_3926,In_1951,In_670);
nand U3927 (N_3927,In_4707,N_469);
nand U3928 (N_3928,In_4626,N_341);
xor U3929 (N_3929,In_1847,N_1878);
xnor U3930 (N_3930,N_1943,N_714);
xnor U3931 (N_3931,N_24,N_676);
nor U3932 (N_3932,N_1728,N_579);
or U3933 (N_3933,N_815,In_648);
nor U3934 (N_3934,N_174,In_4623);
nor U3935 (N_3935,In_1457,N_1465);
nor U3936 (N_3936,N_377,N_1074);
and U3937 (N_3937,N_705,N_477);
xor U3938 (N_3938,N_428,N_1115);
and U3939 (N_3939,In_4571,In_647);
xor U3940 (N_3940,In_194,N_549);
xor U3941 (N_3941,In_4542,N_1123);
and U3942 (N_3942,In_2292,N_1359);
nor U3943 (N_3943,N_537,In_414);
nor U3944 (N_3944,N_1753,In_3350);
nand U3945 (N_3945,N_1505,N_988);
or U3946 (N_3946,In_2533,N_1165);
xnor U3947 (N_3947,N_227,N_1575);
nor U3948 (N_3948,N_77,N_592);
and U3949 (N_3949,N_1392,In_2920);
and U3950 (N_3950,In_2298,In_465);
and U3951 (N_3951,N_1088,In_2939);
and U3952 (N_3952,N_951,N_577);
nor U3953 (N_3953,N_1784,N_1988);
and U3954 (N_3954,In_1452,N_1275);
nor U3955 (N_3955,In_3096,N_1756);
nor U3956 (N_3956,N_1393,In_2335);
nor U3957 (N_3957,N_546,In_4702);
nand U3958 (N_3958,N_1808,N_1891);
and U3959 (N_3959,In_1091,N_482);
nor U3960 (N_3960,N_1494,N_689);
and U3961 (N_3961,N_463,N_1498);
xor U3962 (N_3962,N_1785,N_608);
or U3963 (N_3963,N_1375,N_530);
and U3964 (N_3964,N_22,N_1006);
or U3965 (N_3965,In_2500,N_1194);
nand U3966 (N_3966,In_2508,In_4233);
xnor U3967 (N_3967,In_2165,N_579);
and U3968 (N_3968,N_130,N_1184);
nand U3969 (N_3969,N_659,In_1546);
nor U3970 (N_3970,N_1082,N_1652);
and U3971 (N_3971,N_802,N_1918);
and U3972 (N_3972,N_874,In_351);
and U3973 (N_3973,In_3843,N_1301);
xor U3974 (N_3974,In_2849,N_243);
nor U3975 (N_3975,In_885,N_948);
and U3976 (N_3976,N_313,In_3840);
or U3977 (N_3977,In_1972,N_233);
xnor U3978 (N_3978,N_849,In_4978);
nor U3979 (N_3979,N_1570,In_3411);
xor U3980 (N_3980,In_2138,N_1897);
nand U3981 (N_3981,N_561,N_161);
nand U3982 (N_3982,N_313,N_1799);
xnor U3983 (N_3983,N_1443,N_1323);
and U3984 (N_3984,N_1789,N_1250);
xnor U3985 (N_3985,In_4097,N_259);
nand U3986 (N_3986,In_3253,N_845);
and U3987 (N_3987,N_1188,In_2410);
xnor U3988 (N_3988,In_4233,In_790);
nand U3989 (N_3989,In_581,In_4636);
xor U3990 (N_3990,N_1691,N_298);
nor U3991 (N_3991,N_1947,N_505);
xnor U3992 (N_3992,N_648,In_1019);
or U3993 (N_3993,In_171,In_132);
nand U3994 (N_3994,In_4901,N_66);
or U3995 (N_3995,N_29,In_2428);
nand U3996 (N_3996,In_3249,N_575);
xor U3997 (N_3997,N_1846,In_4818);
or U3998 (N_3998,N_47,N_650);
xnor U3999 (N_3999,N_842,In_4474);
nor U4000 (N_4000,N_2654,N_2977);
nand U4001 (N_4001,N_3312,N_2154);
nand U4002 (N_4002,N_3670,N_3615);
and U4003 (N_4003,N_3474,N_3100);
nor U4004 (N_4004,N_3604,N_3983);
or U4005 (N_4005,N_3215,N_2723);
or U4006 (N_4006,N_2372,N_3045);
nor U4007 (N_4007,N_3674,N_2906);
or U4008 (N_4008,N_3007,N_3158);
nor U4009 (N_4009,N_2568,N_2134);
and U4010 (N_4010,N_2000,N_3816);
and U4011 (N_4011,N_2132,N_3694);
and U4012 (N_4012,N_2042,N_3430);
nor U4013 (N_4013,N_2533,N_2358);
xor U4014 (N_4014,N_3176,N_2005);
xor U4015 (N_4015,N_3463,N_3705);
xnor U4016 (N_4016,N_2843,N_2991);
nand U4017 (N_4017,N_2752,N_3721);
nor U4018 (N_4018,N_2657,N_2873);
or U4019 (N_4019,N_3610,N_3370);
nor U4020 (N_4020,N_3563,N_3508);
and U4021 (N_4021,N_2253,N_2043);
or U4022 (N_4022,N_2213,N_3427);
nand U4023 (N_4023,N_2607,N_2879);
nand U4024 (N_4024,N_3881,N_3682);
and U4025 (N_4025,N_3667,N_2835);
nand U4026 (N_4026,N_2016,N_3933);
or U4027 (N_4027,N_2363,N_3889);
or U4028 (N_4028,N_2829,N_2224);
nor U4029 (N_4029,N_3124,N_2422);
nor U4030 (N_4030,N_3236,N_3573);
nand U4031 (N_4031,N_3336,N_3260);
xor U4032 (N_4032,N_3286,N_2150);
xor U4033 (N_4033,N_2694,N_3301);
xor U4034 (N_4034,N_2442,N_2608);
nand U4035 (N_4035,N_3338,N_3028);
or U4036 (N_4036,N_3685,N_2440);
nand U4037 (N_4037,N_3525,N_3869);
or U4038 (N_4038,N_2047,N_3255);
nand U4039 (N_4039,N_3310,N_2823);
nor U4040 (N_4040,N_3838,N_3799);
and U4041 (N_4041,N_2973,N_2765);
or U4042 (N_4042,N_3015,N_2252);
nand U4043 (N_4043,N_3003,N_3837);
or U4044 (N_4044,N_2196,N_2280);
nand U4045 (N_4045,N_3473,N_3104);
or U4046 (N_4046,N_2255,N_2472);
nor U4047 (N_4047,N_2920,N_2040);
xnor U4048 (N_4048,N_3687,N_2511);
nor U4049 (N_4049,N_2563,N_3668);
nand U4050 (N_4050,N_2424,N_3600);
nor U4051 (N_4051,N_3303,N_3153);
xnor U4052 (N_4052,N_2335,N_3232);
xor U4053 (N_4053,N_2082,N_3396);
xnor U4054 (N_4054,N_2094,N_2558);
nand U4055 (N_4055,N_3186,N_2177);
or U4056 (N_4056,N_2448,N_3718);
nor U4057 (N_4057,N_2902,N_3541);
nor U4058 (N_4058,N_3460,N_3531);
or U4059 (N_4059,N_2249,N_3561);
nand U4060 (N_4060,N_2749,N_2797);
xor U4061 (N_4061,N_2205,N_3331);
nand U4062 (N_4062,N_3676,N_2439);
or U4063 (N_4063,N_2529,N_2460);
nand U4064 (N_4064,N_3137,N_2528);
nand U4065 (N_4065,N_3918,N_2199);
or U4066 (N_4066,N_2524,N_3784);
nand U4067 (N_4067,N_3022,N_2161);
nor U4068 (N_4068,N_2599,N_3327);
and U4069 (N_4069,N_3097,N_2293);
nand U4070 (N_4070,N_2854,N_2167);
nor U4071 (N_4071,N_2171,N_3647);
or U4072 (N_4072,N_2716,N_3517);
xnor U4073 (N_4073,N_3098,N_2832);
nand U4074 (N_4074,N_2061,N_3996);
nand U4075 (N_4075,N_3597,N_3879);
xor U4076 (N_4076,N_3434,N_3841);
nor U4077 (N_4077,N_2767,N_2002);
nand U4078 (N_4078,N_2126,N_3916);
and U4079 (N_4079,N_3972,N_3042);
xor U4080 (N_4080,N_3311,N_3535);
and U4081 (N_4081,N_2294,N_3502);
nor U4082 (N_4082,N_3295,N_3318);
or U4083 (N_4083,N_2600,N_2410);
or U4084 (N_4084,N_2411,N_3372);
nand U4085 (N_4085,N_3570,N_3367);
or U4086 (N_4086,N_3131,N_2690);
nor U4087 (N_4087,N_3533,N_3469);
nor U4088 (N_4088,N_2951,N_3776);
nor U4089 (N_4089,N_2302,N_2284);
nand U4090 (N_4090,N_2142,N_2223);
nand U4091 (N_4091,N_3840,N_2022);
nand U4092 (N_4092,N_2332,N_3140);
nor U4093 (N_4093,N_2816,N_2130);
or U4094 (N_4094,N_3998,N_2646);
nor U4095 (N_4095,N_3689,N_2643);
and U4096 (N_4096,N_2935,N_3126);
nand U4097 (N_4097,N_3806,N_2905);
or U4098 (N_4098,N_2513,N_3686);
nand U4099 (N_4099,N_2421,N_3965);
xnor U4100 (N_4100,N_2926,N_3834);
and U4101 (N_4101,N_2236,N_3757);
nand U4102 (N_4102,N_2446,N_2779);
and U4103 (N_4103,N_2259,N_3872);
nor U4104 (N_4104,N_2079,N_3649);
xnor U4105 (N_4105,N_3530,N_2331);
nand U4106 (N_4106,N_2403,N_3700);
or U4107 (N_4107,N_3760,N_2455);
nor U4108 (N_4108,N_2578,N_2503);
or U4109 (N_4109,N_3431,N_2846);
xor U4110 (N_4110,N_3946,N_2112);
xor U4111 (N_4111,N_3424,N_3302);
or U4112 (N_4112,N_3103,N_2048);
and U4113 (N_4113,N_3221,N_2370);
and U4114 (N_4114,N_3985,N_3127);
xor U4115 (N_4115,N_2787,N_3076);
nor U4116 (N_4116,N_2995,N_3004);
nor U4117 (N_4117,N_2809,N_2173);
or U4118 (N_4118,N_2349,N_3165);
nor U4119 (N_4119,N_3617,N_3388);
or U4120 (N_4120,N_2831,N_2174);
nand U4121 (N_4121,N_2939,N_3375);
or U4122 (N_4122,N_2728,N_3909);
and U4123 (N_4123,N_3267,N_3052);
xor U4124 (N_4124,N_2894,N_3954);
nor U4125 (N_4125,N_3160,N_3216);
nand U4126 (N_4126,N_2093,N_3328);
xnor U4127 (N_4127,N_2508,N_3017);
nor U4128 (N_4128,N_3523,N_2532);
and U4129 (N_4129,N_3788,N_3629);
or U4130 (N_4130,N_2998,N_3264);
xnor U4131 (N_4131,N_2605,N_3813);
and U4132 (N_4132,N_3989,N_3758);
nand U4133 (N_4133,N_2869,N_2390);
or U4134 (N_4134,N_2592,N_3596);
nor U4135 (N_4135,N_3555,N_3402);
nor U4136 (N_4136,N_2121,N_2191);
xor U4137 (N_4137,N_3280,N_2827);
and U4138 (N_4138,N_3270,N_3334);
and U4139 (N_4139,N_3032,N_3298);
xor U4140 (N_4140,N_2006,N_2451);
nand U4141 (N_4141,N_3391,N_3284);
and U4142 (N_4142,N_3754,N_3478);
nand U4143 (N_4143,N_2652,N_2110);
nand U4144 (N_4144,N_2023,N_2516);
nand U4145 (N_4145,N_3102,N_2137);
nand U4146 (N_4146,N_3661,N_2409);
and U4147 (N_4147,N_2287,N_2651);
nand U4148 (N_4148,N_2189,N_3060);
or U4149 (N_4149,N_2758,N_2378);
nand U4150 (N_4150,N_2609,N_2864);
nand U4151 (N_4151,N_2026,N_2891);
xor U4152 (N_4152,N_3575,N_3392);
or U4153 (N_4153,N_3703,N_2895);
nor U4154 (N_4154,N_2678,N_2470);
nand U4155 (N_4155,N_3217,N_2207);
and U4156 (N_4156,N_3458,N_2176);
nor U4157 (N_4157,N_3121,N_3254);
and U4158 (N_4158,N_3969,N_3352);
and U4159 (N_4159,N_2925,N_3404);
xor U4160 (N_4160,N_3543,N_2394);
or U4161 (N_4161,N_3428,N_2887);
or U4162 (N_4162,N_3401,N_2180);
xor U4163 (N_4163,N_3932,N_2763);
and U4164 (N_4164,N_3651,N_2840);
nand U4165 (N_4165,N_3400,N_3897);
nor U4166 (N_4166,N_2083,N_2203);
nor U4167 (N_4167,N_3603,N_2882);
and U4168 (N_4168,N_3901,N_3155);
xor U4169 (N_4169,N_2541,N_3500);
nor U4170 (N_4170,N_2086,N_3751);
nand U4171 (N_4171,N_2943,N_2281);
and U4172 (N_4172,N_3586,N_3992);
and U4173 (N_4173,N_3742,N_2826);
nand U4174 (N_4174,N_3557,N_2756);
nor U4175 (N_4175,N_2957,N_2586);
nand U4176 (N_4176,N_3315,N_3956);
xnor U4177 (N_4177,N_2352,N_3622);
or U4178 (N_4178,N_3783,N_2750);
or U4179 (N_4179,N_3537,N_3021);
xnor U4180 (N_4180,N_2710,N_3406);
and U4181 (N_4181,N_2932,N_3511);
nand U4182 (N_4182,N_2796,N_2534);
nor U4183 (N_4183,N_3099,N_2860);
nor U4184 (N_4184,N_3238,N_3962);
nand U4185 (N_4185,N_3510,N_2789);
and U4186 (N_4186,N_3836,N_3867);
xnor U4187 (N_4187,N_3815,N_3810);
nand U4188 (N_4188,N_2668,N_2052);
xor U4189 (N_4189,N_3566,N_3387);
nor U4190 (N_4190,N_3114,N_3189);
xnor U4191 (N_4191,N_2170,N_2851);
or U4192 (N_4192,N_2389,N_3562);
or U4193 (N_4193,N_2509,N_2703);
nand U4194 (N_4194,N_3496,N_3393);
nand U4195 (N_4195,N_3039,N_2837);
or U4196 (N_4196,N_2613,N_2172);
nand U4197 (N_4197,N_3968,N_3823);
or U4198 (N_4198,N_2665,N_3150);
xnor U4199 (N_4199,N_3398,N_3206);
nand U4200 (N_4200,N_3486,N_3964);
nand U4201 (N_4201,N_2221,N_2368);
and U4202 (N_4202,N_3178,N_2072);
and U4203 (N_4203,N_2077,N_2581);
and U4204 (N_4204,N_3467,N_2536);
or U4205 (N_4205,N_2429,N_3066);
or U4206 (N_4206,N_3378,N_3877);
or U4207 (N_4207,N_2037,N_3316);
or U4208 (N_4208,N_2053,N_2098);
or U4209 (N_4209,N_2493,N_3110);
nor U4210 (N_4210,N_2341,N_2618);
xnor U4211 (N_4211,N_2232,N_3413);
and U4212 (N_4212,N_3792,N_3067);
xor U4213 (N_4213,N_3084,N_3196);
xor U4214 (N_4214,N_3012,N_2660);
nor U4215 (N_4215,N_3138,N_2515);
nor U4216 (N_4216,N_2096,N_2233);
nor U4217 (N_4217,N_3927,N_2111);
nor U4218 (N_4218,N_3513,N_2814);
or U4219 (N_4219,N_2308,N_3584);
nor U4220 (N_4220,N_3937,N_2834);
xnor U4221 (N_4221,N_3288,N_3569);
and U4222 (N_4222,N_2548,N_2744);
or U4223 (N_4223,N_3276,N_2616);
and U4224 (N_4224,N_3726,N_3053);
xor U4225 (N_4225,N_2867,N_2244);
or U4226 (N_4226,N_3187,N_2518);
and U4227 (N_4227,N_3735,N_3619);
xnor U4228 (N_4228,N_3296,N_2215);
nand U4229 (N_4229,N_2907,N_3846);
and U4230 (N_4230,N_2531,N_2754);
xnor U4231 (N_4231,N_2383,N_2899);
xnor U4232 (N_4232,N_2916,N_3292);
or U4233 (N_4233,N_2702,N_3395);
or U4234 (N_4234,N_2418,N_2123);
and U4235 (N_4235,N_3179,N_2011);
or U4236 (N_4236,N_3529,N_2799);
nand U4237 (N_4237,N_2987,N_2041);
nand U4238 (N_4238,N_2550,N_3704);
nor U4239 (N_4239,N_2245,N_2769);
and U4240 (N_4240,N_3074,N_2165);
nor U4241 (N_4241,N_3174,N_3157);
or U4242 (N_4242,N_2343,N_2482);
and U4243 (N_4243,N_3545,N_2007);
nor U4244 (N_4244,N_3766,N_3987);
nand U4245 (N_4245,N_2676,N_3118);
nand U4246 (N_4246,N_2947,N_3034);
and U4247 (N_4247,N_3148,N_3663);
xnor U4248 (N_4248,N_2025,N_2718);
nor U4249 (N_4249,N_3811,N_2068);
and U4250 (N_4250,N_2514,N_3536);
nand U4251 (N_4251,N_2241,N_2641);
or U4252 (N_4252,N_3866,N_3873);
xnor U4253 (N_4253,N_3170,N_3677);
nor U4254 (N_4254,N_3928,N_3835);
nand U4255 (N_4255,N_2419,N_3963);
nor U4256 (N_4256,N_2050,N_3914);
and U4257 (N_4257,N_3480,N_2046);
nand U4258 (N_4258,N_3068,N_2539);
nor U4259 (N_4259,N_3579,N_3379);
nor U4260 (N_4260,N_2024,N_2594);
and U4261 (N_4261,N_2670,N_3779);
nand U4262 (N_4262,N_2788,N_3361);
xor U4263 (N_4263,N_2922,N_3452);
nand U4264 (N_4264,N_3226,N_2512);
and U4265 (N_4265,N_3040,N_3958);
nand U4266 (N_4266,N_3441,N_2521);
or U4267 (N_4267,N_3457,N_3602);
and U4268 (N_4268,N_2152,N_2468);
and U4269 (N_4269,N_3414,N_3553);
or U4270 (N_4270,N_2066,N_2450);
nor U4271 (N_4271,N_3229,N_3159);
nand U4272 (N_4272,N_2675,N_3135);
xor U4273 (N_4273,N_2724,N_2801);
and U4274 (N_4274,N_3773,N_2103);
nor U4275 (N_4275,N_2538,N_2742);
and U4276 (N_4276,N_3059,N_3408);
or U4277 (N_4277,N_3304,N_3297);
xor U4278 (N_4278,N_2510,N_2226);
xor U4279 (N_4279,N_3652,N_2264);
or U4280 (N_4280,N_2507,N_2642);
and U4281 (N_4281,N_2457,N_3384);
or U4282 (N_4282,N_3656,N_2069);
xnor U4283 (N_4283,N_2525,N_2178);
xnor U4284 (N_4284,N_2163,N_2612);
nor U4285 (N_4285,N_2139,N_3803);
and U4286 (N_4286,N_2903,N_2453);
nand U4287 (N_4287,N_2382,N_2685);
and U4288 (N_4288,N_2473,N_3505);
nor U4289 (N_4289,N_3058,N_3141);
and U4290 (N_4290,N_3724,N_2737);
xnor U4291 (N_4291,N_2212,N_3540);
nand U4292 (N_4292,N_3167,N_2380);
and U4293 (N_4293,N_3306,N_2481);
or U4294 (N_4294,N_2279,N_3854);
nor U4295 (N_4295,N_3262,N_2117);
nand U4296 (N_4296,N_3000,N_3990);
or U4297 (N_4297,N_2062,N_2108);
nand U4298 (N_4298,N_3344,N_3415);
or U4299 (N_4299,N_3797,N_2547);
or U4300 (N_4300,N_2099,N_2780);
nand U4301 (N_4301,N_2753,N_2362);
nor U4302 (N_4302,N_2156,N_2311);
or U4303 (N_4303,N_3382,N_3432);
nand U4304 (N_4304,N_3542,N_3849);
nand U4305 (N_4305,N_3934,N_2119);
nand U4306 (N_4306,N_2963,N_2129);
or U4307 (N_4307,N_2603,N_3234);
nor U4308 (N_4308,N_2396,N_3199);
and U4309 (N_4309,N_2949,N_2102);
nor U4310 (N_4310,N_3719,N_3504);
nor U4311 (N_4311,N_3623,N_3678);
and U4312 (N_4312,N_2719,N_3714);
nand U4313 (N_4313,N_3935,N_2771);
nor U4314 (N_4314,N_3082,N_2461);
and U4315 (N_4315,N_3429,N_2088);
or U4316 (N_4316,N_2234,N_2138);
and U4317 (N_4317,N_3892,N_2530);
nor U4318 (N_4318,N_3061,N_2218);
nand U4319 (N_4319,N_2970,N_2036);
or U4320 (N_4320,N_3534,N_3886);
nand U4321 (N_4321,N_2008,N_2373);
or U4322 (N_4322,N_3509,N_3787);
nand U4323 (N_4323,N_2804,N_2722);
xnor U4324 (N_4324,N_2115,N_3321);
or U4325 (N_4325,N_3043,N_3056);
xnor U4326 (N_4326,N_3208,N_3911);
or U4327 (N_4327,N_3466,N_2790);
and U4328 (N_4328,N_3633,N_3494);
nand U4329 (N_4329,N_3743,N_2059);
or U4330 (N_4330,N_2051,N_2638);
nand U4331 (N_4331,N_2464,N_3885);
nor U4332 (N_4332,N_2385,N_3723);
or U4333 (N_4333,N_2397,N_3612);
and U4334 (N_4334,N_3926,N_2499);
nor U4335 (N_4335,N_2549,N_3746);
nand U4336 (N_4336,N_2113,N_2168);
and U4337 (N_4337,N_2746,N_2961);
or U4338 (N_4338,N_2818,N_3961);
xnor U4339 (N_4339,N_3922,N_2198);
and U4340 (N_4340,N_2865,N_3411);
nor U4341 (N_4341,N_2462,N_3679);
xnor U4342 (N_4342,N_3499,N_3636);
or U4343 (N_4343,N_2348,N_2222);
nor U4344 (N_4344,N_2713,N_3775);
nand U4345 (N_4345,N_3246,N_3093);
nor U4346 (N_4346,N_3330,N_2375);
xor U4347 (N_4347,N_2900,N_3078);
and U4348 (N_4348,N_2700,N_2821);
nor U4349 (N_4349,N_3213,N_2587);
xnor U4350 (N_4350,N_2242,N_3732);
nor U4351 (N_4351,N_2291,N_2169);
xnor U4352 (N_4352,N_3745,N_2185);
or U4353 (N_4353,N_2488,N_3878);
nor U4354 (N_4354,N_2369,N_3089);
nand U4355 (N_4355,N_2452,N_3339);
xnor U4356 (N_4356,N_2565,N_2795);
nand U4357 (N_4357,N_2246,N_3606);
xnor U4358 (N_4358,N_3168,N_2803);
xnor U4359 (N_4359,N_3607,N_3852);
nor U4360 (N_4360,N_3699,N_2420);
or U4361 (N_4361,N_3701,N_3894);
nand U4362 (N_4362,N_3422,N_2334);
nor U4363 (N_4363,N_2144,N_3626);
and U4364 (N_4364,N_3483,N_3193);
or U4365 (N_4365,N_2915,N_3580);
xor U4366 (N_4366,N_3472,N_2190);
and U4367 (N_4367,N_3461,N_3861);
xnor U4368 (N_4368,N_3695,N_3278);
nor U4369 (N_4369,N_3948,N_3605);
xnor U4370 (N_4370,N_2553,N_2064);
nor U4371 (N_4371,N_3717,N_2273);
nor U4372 (N_4372,N_2009,N_3549);
or U4373 (N_4373,N_2393,N_3591);
xnor U4374 (N_4374,N_2761,N_3681);
xor U4375 (N_4375,N_2105,N_2251);
xor U4376 (N_4376,N_2354,N_2625);
and U4377 (N_4377,N_2444,N_2564);
and U4378 (N_4378,N_3405,N_3993);
nor U4379 (N_4379,N_3036,N_3203);
nand U4380 (N_4380,N_3675,N_3786);
and U4381 (N_4381,N_2543,N_2433);
nor U4382 (N_4382,N_2181,N_3738);
nor U4383 (N_4383,N_2910,N_2732);
nor U4384 (N_4384,N_3495,N_3433);
or U4385 (N_4385,N_2381,N_2076);
nand U4386 (N_4386,N_2884,N_2590);
nand U4387 (N_4387,N_3149,N_3123);
or U4388 (N_4388,N_2931,N_2591);
nand U4389 (N_4389,N_2347,N_2576);
nor U4390 (N_4390,N_3484,N_2658);
xor U4391 (N_4391,N_2175,N_2313);
xnor U4392 (N_4392,N_2365,N_3490);
or U4393 (N_4393,N_2239,N_2684);
or U4394 (N_4394,N_3639,N_2885);
nor U4395 (N_4395,N_3645,N_3613);
xnor U4396 (N_4396,N_3005,N_3556);
nor U4397 (N_4397,N_3368,N_2817);
xor U4398 (N_4398,N_2540,N_3666);
nor U4399 (N_4399,N_2946,N_2351);
xor U4400 (N_4400,N_2345,N_2184);
or U4401 (N_4401,N_2208,N_2248);
and U4402 (N_4402,N_2376,N_3275);
nand U4403 (N_4403,N_3120,N_3539);
or U4404 (N_4404,N_2933,N_2104);
or U4405 (N_4405,N_2889,N_3857);
and U4406 (N_4406,N_3876,N_2357);
or U4407 (N_4407,N_2193,N_3895);
nand U4408 (N_4408,N_3527,N_3250);
nor U4409 (N_4409,N_3271,N_2621);
xnor U4410 (N_4410,N_3654,N_3506);
nand U4411 (N_4411,N_3048,N_3741);
nand U4412 (N_4412,N_2140,N_3163);
nand U4413 (N_4413,N_3581,N_2400);
xnor U4414 (N_4414,N_3664,N_2990);
and U4415 (N_4415,N_3062,N_3353);
or U4416 (N_4416,N_2489,N_3212);
or U4417 (N_4417,N_2467,N_2339);
nand U4418 (N_4418,N_2116,N_2941);
nand U4419 (N_4419,N_2633,N_2655);
nand U4420 (N_4420,N_2686,N_2209);
or U4421 (N_4421,N_3180,N_2782);
xor U4422 (N_4422,N_3294,N_3354);
nand U4423 (N_4423,N_3641,N_2325);
and U4424 (N_4424,N_3790,N_3905);
nand U4425 (N_4425,N_3266,N_2555);
and U4426 (N_4426,N_2322,N_3269);
and U4427 (N_4427,N_2984,N_2361);
or U4428 (N_4428,N_3913,N_3978);
nand U4429 (N_4429,N_3439,N_2778);
xor U4430 (N_4430,N_2537,N_3013);
xnor U4431 (N_4431,N_3655,N_2960);
or U4432 (N_4432,N_2741,N_2261);
xor U4433 (N_4433,N_3514,N_2477);
and U4434 (N_4434,N_2055,N_2135);
nand U4435 (N_4435,N_2101,N_3038);
nand U4436 (N_4436,N_3863,N_2927);
xor U4437 (N_4437,N_3026,N_3493);
nor U4438 (N_4438,N_3018,N_2704);
nor U4439 (N_4439,N_3410,N_3739);
nor U4440 (N_4440,N_2263,N_2972);
nor U4441 (N_4441,N_3839,N_3988);
nand U4442 (N_4442,N_2691,N_2425);
or U4443 (N_4443,N_3436,N_2274);
xor U4444 (N_4444,N_2890,N_3397);
and U4445 (N_4445,N_3862,N_2542);
nand U4446 (N_4446,N_3448,N_2109);
nand U4447 (N_4447,N_3921,N_3554);
xor U4448 (N_4448,N_3290,N_3628);
and U4449 (N_4449,N_2974,N_2692);
and U4450 (N_4450,N_2794,N_2388);
nor U4451 (N_4451,N_3577,N_2614);
or U4452 (N_4452,N_3244,N_2876);
and U4453 (N_4453,N_2214,N_3202);
and U4454 (N_4454,N_2644,N_2211);
or U4455 (N_4455,N_2635,N_2342);
nand U4456 (N_4456,N_2045,N_3955);
or U4457 (N_4457,N_3172,N_3241);
or U4458 (N_4458,N_3750,N_3309);
or U4459 (N_4459,N_2930,N_2768);
or U4460 (N_4460,N_2909,N_3008);
nor U4461 (N_4461,N_3594,N_2063);
xnor U4462 (N_4462,N_3357,N_3890);
nor U4463 (N_4463,N_3403,N_2777);
nand U4464 (N_4464,N_2559,N_2838);
xor U4465 (N_4465,N_3497,N_3971);
and U4466 (N_4466,N_3171,N_3571);
xnor U4467 (N_4467,N_3332,N_3548);
xnor U4468 (N_4468,N_3512,N_2001);
xnor U4469 (N_4469,N_2852,N_3377);
xor U4470 (N_4470,N_3169,N_2430);
nor U4471 (N_4471,N_2812,N_2019);
and U4472 (N_4472,N_3143,N_2791);
nor U4473 (N_4473,N_3273,N_3808);
xor U4474 (N_4474,N_2798,N_2551);
and U4475 (N_4475,N_3821,N_2377);
xor U4476 (N_4476,N_3374,N_2060);
nor U4477 (N_4477,N_2427,N_2632);
and U4478 (N_4478,N_2924,N_3325);
nor U4479 (N_4479,N_3347,N_2863);
nor U4480 (N_4480,N_2476,N_3669);
nand U4481 (N_4481,N_3830,N_2828);
or U4482 (N_4482,N_3091,N_2384);
nor U4483 (N_4483,N_3322,N_2288);
or U4484 (N_4484,N_2556,N_2398);
and U4485 (N_4485,N_3842,N_2575);
xnor U4486 (N_4486,N_2321,N_2483);
xnor U4487 (N_4487,N_3106,N_2344);
and U4488 (N_4488,N_2875,N_3945);
nor U4489 (N_4489,N_3907,N_3247);
nor U4490 (N_4490,N_2441,N_2602);
and U4491 (N_4491,N_2028,N_3481);
nor U4492 (N_4492,N_2095,N_2087);
xor U4493 (N_4493,N_3634,N_3552);
nand U4494 (N_4494,N_2959,N_2844);
and U4495 (N_4495,N_3477,N_3740);
nor U4496 (N_4496,N_2664,N_2604);
nor U4497 (N_4497,N_2029,N_3319);
and U4498 (N_4498,N_3708,N_3200);
xnor U4499 (N_4499,N_3888,N_2672);
xor U4500 (N_4500,N_3030,N_2136);
xnor U4501 (N_4501,N_2751,N_3692);
and U4502 (N_4502,N_2770,N_2486);
nand U4503 (N_4503,N_2387,N_2883);
nand U4504 (N_4504,N_2364,N_3590);
nand U4505 (N_4505,N_3770,N_2426);
nor U4506 (N_4506,N_3774,N_3129);
xor U4507 (N_4507,N_3939,N_3248);
or U4508 (N_4508,N_2725,N_3936);
nor U4509 (N_4509,N_3417,N_3489);
xor U4510 (N_4510,N_3930,N_2494);
nor U4511 (N_4511,N_2738,N_3219);
nor U4512 (N_4512,N_2650,N_3642);
or U4513 (N_4513,N_3999,N_2501);
nand U4514 (N_4514,N_2519,N_2412);
nand U4515 (N_4515,N_2622,N_3583);
or U4516 (N_4516,N_2997,N_2289);
nand U4517 (N_4517,N_2333,N_2897);
nor U4518 (N_4518,N_3230,N_2012);
or U4519 (N_4519,N_2912,N_3109);
and U4520 (N_4520,N_2159,N_3501);
or U4521 (N_4521,N_3025,N_2228);
nor U4522 (N_4522,N_3997,N_3363);
xor U4523 (N_4523,N_2458,N_3782);
nand U4524 (N_4524,N_3265,N_3329);
or U4525 (N_4525,N_2454,N_3585);
and U4526 (N_4526,N_2893,N_3348);
xor U4527 (N_4527,N_3285,N_3145);
nand U4528 (N_4528,N_3112,N_3228);
nand U4529 (N_4529,N_3360,N_2407);
or U4530 (N_4530,N_2148,N_2597);
nand U4531 (N_4531,N_3454,N_3435);
nand U4532 (N_4532,N_2975,N_2092);
nand U4533 (N_4533,N_3730,N_3092);
nor U4534 (N_4534,N_3680,N_3528);
or U4535 (N_4535,N_3049,N_3672);
and U4536 (N_4536,N_2696,N_2449);
xor U4537 (N_4537,N_3188,N_3618);
or U4538 (N_4538,N_2731,N_2588);
nand U4539 (N_4539,N_2661,N_3173);
nand U4540 (N_4540,N_3002,N_3812);
and U4541 (N_4541,N_2100,N_3064);
xnor U4542 (N_4542,N_3952,N_2904);
nand U4543 (N_4543,N_3252,N_3399);
nand U4544 (N_4544,N_3683,N_3749);
xnor U4545 (N_4545,N_3507,N_2316);
nor U4546 (N_4546,N_2300,N_2557);
or U4547 (N_4547,N_2219,N_3698);
nand U4548 (N_4548,N_3546,N_2734);
nand U4549 (N_4549,N_2114,N_2089);
xor U4550 (N_4550,N_2438,N_2629);
xnor U4551 (N_4551,N_2118,N_2766);
and U4552 (N_4552,N_3027,N_2631);
nand U4553 (N_4553,N_2416,N_3132);
nand U4554 (N_4554,N_2182,N_2526);
nor U4555 (N_4555,N_3204,N_2067);
nor U4556 (N_4556,N_3598,N_2697);
xnor U4557 (N_4557,N_2162,N_2404);
nor U4558 (N_4558,N_3748,N_2853);
xor U4559 (N_4559,N_2120,N_2978);
nor U4560 (N_4560,N_3083,N_2923);
and U4561 (N_4561,N_3720,N_3957);
xnor U4562 (N_4562,N_2706,N_2445);
xnor U4563 (N_4563,N_3055,N_2034);
and U4564 (N_4564,N_3065,N_3035);
nor U4565 (N_4565,N_2431,N_2892);
nand U4566 (N_4566,N_2994,N_2004);
xor U4567 (N_4567,N_2671,N_2535);
or U4568 (N_4568,N_2955,N_3938);
xnor U4569 (N_4569,N_2679,N_3595);
nand U4570 (N_4570,N_3919,N_2478);
xor U4571 (N_4571,N_3638,N_2554);
or U4572 (N_4572,N_3565,N_3272);
nor U4573 (N_4573,N_2337,N_3482);
nand U4574 (N_4574,N_2392,N_3342);
nor U4575 (N_4575,N_3016,N_2669);
xor U4576 (N_4576,N_2183,N_3421);
xor U4577 (N_4577,N_2802,N_2969);
and U4578 (N_4578,N_3896,N_3182);
nor U4579 (N_4579,N_2201,N_2775);
nand U4580 (N_4580,N_2149,N_3195);
and U4581 (N_4581,N_3258,N_2628);
xnor U4582 (N_4582,N_3376,N_2545);
and U4583 (N_4583,N_3744,N_2320);
or U4584 (N_4584,N_3593,N_3462);
or U4585 (N_4585,N_2262,N_2841);
nand U4586 (N_4586,N_3868,N_2032);
nor U4587 (N_4587,N_3568,N_3665);
xnor U4588 (N_4588,N_2656,N_3800);
and U4589 (N_4589,N_2286,N_2074);
nand U4590 (N_4590,N_3931,N_3259);
nor U4591 (N_4591,N_2634,N_3524);
or U4592 (N_4592,N_2459,N_2391);
or U4593 (N_4593,N_3383,N_3305);
xor U4594 (N_4594,N_3809,N_2265);
xnor U4595 (N_4595,N_2755,N_3381);
nor U4596 (N_4596,N_2953,N_2128);
and U4597 (N_4597,N_2940,N_3054);
and U4598 (N_4598,N_2805,N_3712);
nand U4599 (N_4599,N_2463,N_2146);
and U4600 (N_4600,N_2680,N_2921);
xnor U4601 (N_4601,N_2405,N_2709);
xor U4602 (N_4602,N_3449,N_2496);
nor U4603 (N_4603,N_3802,N_3156);
or U4604 (N_4604,N_3753,N_2570);
nand U4605 (N_4605,N_2056,N_2465);
nand U4606 (N_4606,N_3818,N_3785);
or U4607 (N_4607,N_3161,N_3822);
and U4608 (N_4608,N_2996,N_2626);
and U4609 (N_4609,N_3242,N_2272);
and U4610 (N_4610,N_2582,N_2985);
nand U4611 (N_4611,N_2944,N_3558);
or U4612 (N_4612,N_2304,N_2317);
nor U4613 (N_4613,N_2667,N_3950);
nor U4614 (N_4614,N_3438,N_2663);
or U4615 (N_4615,N_3152,N_2648);
and U4616 (N_4616,N_2645,N_3237);
or U4617 (N_4617,N_2436,N_2266);
nand U4618 (N_4618,N_3476,N_2282);
nand U4619 (N_4619,N_3105,N_2329);
or U4620 (N_4620,N_3047,N_3116);
xor U4621 (N_4621,N_3346,N_3807);
and U4622 (N_4622,N_3702,N_2874);
nand U4623 (N_4623,N_3653,N_2982);
xor U4624 (N_4624,N_3487,N_2275);
and U4625 (N_4625,N_2014,N_2886);
and U4626 (N_4626,N_2808,N_3673);
nand U4627 (N_4627,N_3940,N_2229);
or U4628 (N_4628,N_3906,N_2839);
or U4629 (N_4629,N_2033,N_2367);
xnor U4630 (N_4630,N_2466,N_3077);
or U4631 (N_4631,N_2911,N_3826);
xnor U4632 (N_4632,N_3728,N_3337);
nor U4633 (N_4633,N_2027,N_2620);
xor U4634 (N_4634,N_2267,N_2845);
or U4635 (N_4635,N_3870,N_3974);
xor U4636 (N_4636,N_3804,N_3609);
xor U4637 (N_4637,N_2967,N_3207);
or U4638 (N_4638,N_3780,N_3859);
nand U4639 (N_4639,N_3589,N_3817);
nor U4640 (N_4640,N_3865,N_2993);
nor U4641 (N_4641,N_2585,N_2571);
or U4642 (N_4642,N_2500,N_2965);
nor U4643 (N_4643,N_3194,N_2240);
or U4644 (N_4644,N_3847,N_3991);
nor U4645 (N_4645,N_2131,N_2980);
nand U4646 (N_4646,N_2402,N_2729);
or U4647 (N_4647,N_3139,N_3759);
xor U4648 (N_4648,N_3086,N_2566);
xor U4649 (N_4649,N_3908,N_3883);
or U4650 (N_4650,N_2938,N_3011);
nand U4651 (N_4651,N_2714,N_3085);
xor U4652 (N_4652,N_3544,N_3224);
xor U4653 (N_4653,N_2552,N_2764);
xor U4654 (N_4654,N_3416,N_3671);
nor U4655 (N_4655,N_2659,N_2793);
or U4656 (N_4656,N_3136,N_3335);
and U4657 (N_4657,N_3162,N_3041);
or U4658 (N_4658,N_2480,N_3833);
and U4659 (N_4659,N_2247,N_2647);
nor U4660 (N_4660,N_2862,N_2399);
and U4661 (N_4661,N_3268,N_2127);
or U4662 (N_4662,N_2071,N_3240);
or U4663 (N_4663,N_3825,N_2340);
xor U4664 (N_4664,N_2784,N_2250);
or U4665 (N_4665,N_2054,N_2231);
or U4666 (N_4666,N_2210,N_3736);
and U4667 (N_4667,N_2235,N_3166);
xnor U4668 (N_4668,N_2623,N_2155);
xnor U4669 (N_4669,N_2810,N_2151);
nor U4670 (N_4670,N_3796,N_2021);
nor U4671 (N_4671,N_3350,N_3475);
xnor U4672 (N_4672,N_2206,N_2683);
xnor U4673 (N_4673,N_2983,N_3616);
and U4674 (N_4674,N_3443,N_3635);
or U4675 (N_4675,N_3426,N_3079);
nand U4676 (N_4676,N_2822,N_3063);
or U4677 (N_4677,N_3437,N_2868);
and U4678 (N_4678,N_3516,N_3731);
xnor U4679 (N_4679,N_2836,N_3684);
nand U4680 (N_4680,N_3197,N_3177);
xnor U4681 (N_4681,N_3640,N_2580);
nand U4682 (N_4682,N_2490,N_3643);
xor U4683 (N_4683,N_3094,N_2619);
nor U4684 (N_4684,N_2330,N_2505);
and U4685 (N_4685,N_3364,N_2666);
nor U4686 (N_4686,N_3960,N_3853);
and U4687 (N_4687,N_2057,N_3115);
and U4688 (N_4688,N_3944,N_3324);
and U4689 (N_4689,N_2701,N_2277);
and U4690 (N_4690,N_3175,N_3282);
xnor U4691 (N_4691,N_3729,N_2687);
or U4692 (N_4692,N_3756,N_3824);
or U4693 (N_4693,N_2825,N_3887);
nand U4694 (N_4694,N_2065,N_3394);
or U4695 (N_4695,N_3631,N_2217);
or U4696 (N_4696,N_2187,N_2640);
nand U4697 (N_4697,N_3072,N_2073);
and U4698 (N_4698,N_3560,N_3884);
nand U4699 (N_4699,N_3769,N_2649);
xor U4700 (N_4700,N_3491,N_3794);
or U4701 (N_4701,N_3929,N_3767);
or U4702 (N_4702,N_3874,N_2447);
xnor U4703 (N_4703,N_2039,N_2192);
nand U4704 (N_4704,N_2268,N_2842);
xor U4705 (N_4705,N_2085,N_2319);
xnor U4706 (N_4706,N_2356,N_2598);
or U4707 (N_4707,N_2018,N_3690);
and U4708 (N_4708,N_2200,N_3088);
or U4709 (N_4709,N_2958,N_3380);
and U4710 (N_4710,N_2674,N_3696);
and U4711 (N_4711,N_3198,N_3185);
nor U4712 (N_4712,N_2583,N_3220);
nor U4713 (N_4713,N_2739,N_3341);
nor U4714 (N_4714,N_3146,N_3941);
nor U4715 (N_4715,N_3468,N_2830);
nor U4716 (N_4716,N_2299,N_3761);
and U4717 (N_4717,N_2456,N_3253);
xor U4718 (N_4718,N_2318,N_2374);
nand U4719 (N_4719,N_2964,N_3033);
or U4720 (N_4720,N_3624,N_2495);
nand U4721 (N_4721,N_3805,N_2708);
nor U4722 (N_4722,N_3716,N_3087);
xor U4723 (N_4723,N_3819,N_3009);
and U4724 (N_4724,N_2479,N_2355);
nand U4725 (N_4725,N_2971,N_2914);
nor U4726 (N_4726,N_3459,N_3828);
nor U4727 (N_4727,N_3080,N_3791);
nand U4728 (N_4728,N_3407,N_3359);
nand U4729 (N_4729,N_2471,N_2371);
nand U4730 (N_4730,N_3233,N_3455);
nand U4731 (N_4731,N_2871,N_2015);
nand U4732 (N_4732,N_2800,N_3995);
and U4733 (N_4733,N_2237,N_3650);
xor U4734 (N_4734,N_2760,N_3071);
nand U4735 (N_4735,N_2270,N_2908);
and U4736 (N_4736,N_3953,N_2188);
or U4737 (N_4737,N_2035,N_3801);
and U4738 (N_4738,N_2258,N_2950);
xnor U4739 (N_4739,N_3706,N_3864);
xor U4740 (N_4740,N_3725,N_2715);
and U4741 (N_4741,N_2745,N_3688);
nand U4742 (N_4742,N_2013,N_3521);
nand U4743 (N_4743,N_2157,N_3313);
xor U4744 (N_4744,N_2981,N_2569);
nor U4745 (N_4745,N_3850,N_2928);
nand U4746 (N_4746,N_2593,N_2194);
and U4747 (N_4747,N_3925,N_2336);
nor U4748 (N_4748,N_3444,N_2107);
or U4749 (N_4749,N_2058,N_3979);
nor U4750 (N_4750,N_3442,N_2145);
nand U4751 (N_4751,N_3772,N_2968);
xnor U4752 (N_4752,N_2937,N_3893);
nor U4753 (N_4753,N_2820,N_3632);
or U4754 (N_4754,N_3522,N_2888);
nor U4755 (N_4755,N_3777,N_2179);
or U4756 (N_4756,N_3291,N_3902);
nor U4757 (N_4757,N_3113,N_2824);
xor U4758 (N_4758,N_3820,N_2727);
nand U4759 (N_4759,N_2870,N_3201);
xnor U4760 (N_4760,N_2254,N_3592);
xor U4761 (N_4761,N_3747,N_2003);
nand U4762 (N_4762,N_2491,N_3470);
nand U4763 (N_4763,N_2819,N_3119);
nor U4764 (N_4764,N_2278,N_2918);
nor U4765 (N_4765,N_3358,N_3323);
xor U4766 (N_4766,N_3386,N_2673);
xor U4767 (N_4767,N_3658,N_3620);
nor U4768 (N_4768,N_2785,N_3898);
xor U4769 (N_4769,N_3707,N_3423);
nor U4770 (N_4770,N_3257,N_2502);
nor U4771 (N_4771,N_2297,N_3856);
nand U4772 (N_4772,N_3293,N_3320);
or U4773 (N_4773,N_3691,N_3418);
or U4774 (N_4774,N_2807,N_2522);
nand U4775 (N_4775,N_3567,N_2090);
nand U4776 (N_4776,N_3218,N_2919);
or U4777 (N_4777,N_3515,N_2757);
and U4778 (N_4778,N_2084,N_2589);
nor U4779 (N_4779,N_2220,N_3019);
and U4780 (N_4780,N_2730,N_2901);
xnor U4781 (N_4781,N_2081,N_3637);
nand U4782 (N_4782,N_3069,N_2896);
nor U4783 (N_4783,N_2269,N_2681);
nor U4784 (N_4784,N_3981,N_2283);
nand U4785 (N_4785,N_2527,N_3831);
nor U4786 (N_4786,N_3882,N_3184);
and U4787 (N_4787,N_3147,N_3644);
and U4788 (N_4788,N_2164,N_3287);
nor U4789 (N_4789,N_3860,N_2806);
or U4790 (N_4790,N_2562,N_2271);
nor U4791 (N_4791,N_3793,N_3343);
xnor U4792 (N_4792,N_2080,N_2075);
and U4793 (N_4793,N_3660,N_2406);
nand U4794 (N_4794,N_2606,N_2573);
nor U4795 (N_4795,N_3975,N_2366);
and U4796 (N_4796,N_2707,N_3465);
or U4797 (N_4797,N_2952,N_3814);
and U4798 (N_4798,N_3389,N_3243);
nand U4799 (N_4799,N_2498,N_3755);
xor U4800 (N_4800,N_3037,N_3648);
or U4801 (N_4801,N_3715,N_3662);
xor U4802 (N_4802,N_2567,N_2296);
nand U4803 (N_4803,N_2601,N_3845);
or U4804 (N_4804,N_3281,N_2546);
nor U4805 (N_4805,N_2721,N_2848);
nor U4806 (N_4806,N_3559,N_2303);
and U4807 (N_4807,N_2520,N_2492);
or U4808 (N_4808,N_3959,N_3345);
nor U4809 (N_4809,N_2740,N_3789);
and U4810 (N_4810,N_2662,N_2811);
and U4811 (N_4811,N_3574,N_2160);
and U4812 (N_4812,N_2857,N_3125);
or U4813 (N_4813,N_3190,N_2423);
nand U4814 (N_4814,N_3709,N_3154);
and U4815 (N_4815,N_3970,N_3299);
nor U4816 (N_4816,N_3029,N_3711);
xnor U4817 (N_4817,N_2966,N_3924);
and U4818 (N_4818,N_2762,N_2849);
nor U4819 (N_4819,N_3044,N_3317);
or U4820 (N_4820,N_2636,N_2295);
nand U4821 (N_4821,N_2204,N_3915);
nor U4822 (N_4822,N_2125,N_2504);
and U4823 (N_4823,N_2202,N_3231);
nand U4824 (N_4824,N_3440,N_3976);
nand U4825 (N_4825,N_2359,N_2748);
and U4826 (N_4826,N_2484,N_2166);
nor U4827 (N_4827,N_2030,N_2786);
xnor U4828 (N_4828,N_3899,N_3263);
nor U4829 (N_4829,N_2736,N_3453);
or U4830 (N_4830,N_3073,N_2743);
and U4831 (N_4831,N_2913,N_3277);
or U4832 (N_4832,N_2350,N_2773);
or U4833 (N_4833,N_3737,N_3625);
nand U4834 (N_4834,N_2637,N_2195);
or U4835 (N_4835,N_3947,N_3710);
nand U4836 (N_4836,N_2759,N_3485);
nor U4837 (N_4837,N_2353,N_3464);
nor U4838 (N_4838,N_3134,N_2298);
and U4839 (N_4839,N_2326,N_3447);
and U4840 (N_4840,N_3130,N_3239);
nand U4841 (N_4841,N_2850,N_2310);
xnor U4842 (N_4842,N_3122,N_2948);
and U4843 (N_4843,N_3456,N_3977);
xor U4844 (N_4844,N_2485,N_3734);
or U4845 (N_4845,N_2256,N_2677);
or U4846 (N_4846,N_2813,N_3657);
nor U4847 (N_4847,N_2772,N_2312);
xor U4848 (N_4848,N_2639,N_2610);
and U4849 (N_4849,N_2954,N_2106);
nand U4850 (N_4850,N_2230,N_2833);
and U4851 (N_4851,N_2315,N_2305);
or U4852 (N_4852,N_3621,N_3183);
or U4853 (N_4853,N_3046,N_3843);
nand U4854 (N_4854,N_3051,N_2717);
or U4855 (N_4855,N_2976,N_3599);
nand U4856 (N_4856,N_3564,N_3910);
or U4857 (N_4857,N_3697,N_2861);
or U4858 (N_4858,N_3614,N_3001);
or U4859 (N_4859,N_3300,N_3451);
xnor U4860 (N_4860,N_2415,N_2747);
or U4861 (N_4861,N_3369,N_3526);
and U4862 (N_4862,N_3659,N_3763);
and U4863 (N_4863,N_2227,N_3307);
nor U4864 (N_4864,N_2044,N_3117);
xnor U4865 (N_4865,N_2097,N_3880);
or U4866 (N_4866,N_2934,N_2611);
nand U4867 (N_4867,N_3986,N_3848);
or U4868 (N_4868,N_2487,N_2574);
and U4869 (N_4869,N_3980,N_2523);
or U4870 (N_4870,N_3778,N_3450);
and U4871 (N_4871,N_3627,N_3075);
or U4872 (N_4872,N_2699,N_2945);
xnor U4873 (N_4873,N_3020,N_2561);
nand U4874 (N_4874,N_2881,N_3191);
nand U4875 (N_4875,N_3727,N_3050);
nor U4876 (N_4876,N_2401,N_3951);
nand U4877 (N_4877,N_2158,N_2783);
nand U4878 (N_4878,N_3479,N_3781);
nor U4879 (N_4879,N_2010,N_3151);
nand U4880 (N_4880,N_2847,N_2705);
and U4881 (N_4881,N_2630,N_2314);
or U4882 (N_4882,N_2624,N_3984);
and U4883 (N_4883,N_2497,N_3920);
or U4884 (N_4884,N_3762,N_3014);
nand U4885 (N_4885,N_3587,N_3764);
xnor U4886 (N_4886,N_2328,N_3425);
nor U4887 (N_4887,N_3289,N_3576);
nand U4888 (N_4888,N_3795,N_3355);
xor U4889 (N_4889,N_2858,N_2124);
or U4890 (N_4890,N_3142,N_3409);
and U4891 (N_4891,N_2225,N_3733);
xnor U4892 (N_4892,N_2346,N_2017);
nor U4893 (N_4893,N_2443,N_2859);
xnor U4894 (N_4894,N_3274,N_3608);
nor U4895 (N_4895,N_3518,N_3752);
nand U4896 (N_4896,N_3851,N_3349);
or U4897 (N_4897,N_3765,N_2992);
nand U4898 (N_4898,N_3108,N_2292);
or U4899 (N_4899,N_3235,N_2877);
or U4900 (N_4900,N_3949,N_3023);
nor U4901 (N_4901,N_3832,N_3031);
xor U4902 (N_4902,N_3192,N_3006);
or U4903 (N_4903,N_2049,N_2216);
xor U4904 (N_4904,N_2872,N_2474);
nor U4905 (N_4905,N_3611,N_2327);
or U4906 (N_4906,N_3798,N_2720);
or U4907 (N_4907,N_3256,N_3283);
nand U4908 (N_4908,N_2942,N_3520);
nand U4909 (N_4909,N_3551,N_3722);
nand U4910 (N_4910,N_3858,N_3326);
nand U4911 (N_4911,N_3471,N_2475);
nor U4912 (N_4912,N_2544,N_2695);
and U4913 (N_4913,N_3601,N_3855);
xor U4914 (N_4914,N_2428,N_2413);
and U4915 (N_4915,N_3912,N_2437);
nand U4916 (N_4916,N_2584,N_3973);
nor U4917 (N_4917,N_2956,N_2698);
or U4918 (N_4918,N_3214,N_3111);
nand U4919 (N_4919,N_2309,N_3373);
nand U4920 (N_4920,N_3446,N_2379);
and U4921 (N_4921,N_3492,N_3827);
xor U4922 (N_4922,N_2020,N_3340);
nand U4923 (N_4923,N_3095,N_3519);
and U4924 (N_4924,N_2962,N_2866);
nor U4925 (N_4925,N_3181,N_3871);
and U4926 (N_4926,N_3829,N_2323);
xnor U4927 (N_4927,N_2435,N_2290);
xor U4928 (N_4928,N_3646,N_3227);
nor U4929 (N_4929,N_3875,N_3128);
nor U4930 (N_4930,N_3923,N_3308);
and U4931 (N_4931,N_2577,N_2979);
nand U4932 (N_4932,N_2386,N_2735);
and U4933 (N_4933,N_3024,N_2693);
nand U4934 (N_4934,N_3365,N_2615);
nor U4935 (N_4935,N_2653,N_3503);
and U4936 (N_4936,N_3538,N_3982);
or U4937 (N_4937,N_3356,N_2133);
nand U4938 (N_4938,N_2238,N_2776);
or U4939 (N_4939,N_2469,N_3222);
nor U4940 (N_4940,N_2338,N_3070);
nor U4941 (N_4941,N_3942,N_3385);
xnor U4942 (N_4942,N_3420,N_2260);
or U4943 (N_4943,N_3488,N_2078);
nand U4944 (N_4944,N_2153,N_3900);
or U4945 (N_4945,N_2408,N_2091);
nand U4946 (N_4946,N_2560,N_2792);
and U4947 (N_4947,N_3205,N_2596);
nand U4948 (N_4948,N_3693,N_2147);
xor U4949 (N_4949,N_2989,N_3390);
or U4950 (N_4950,N_3366,N_3419);
or U4951 (N_4951,N_2917,N_2733);
or U4952 (N_4952,N_3768,N_3578);
nor U4953 (N_4953,N_2988,N_3844);
nor U4954 (N_4954,N_2432,N_3994);
or U4955 (N_4955,N_3412,N_3245);
nand U4956 (N_4956,N_3550,N_3445);
nor U4957 (N_4957,N_3223,N_2579);
or U4958 (N_4958,N_2880,N_2434);
or U4959 (N_4959,N_2878,N_2517);
nand U4960 (N_4960,N_2572,N_3279);
nand U4961 (N_4961,N_3891,N_3211);
xor U4962 (N_4962,N_2276,N_2781);
nand U4963 (N_4963,N_3133,N_3362);
nor U4964 (N_4964,N_2031,N_2712);
or U4965 (N_4965,N_3532,N_3010);
nor U4966 (N_4966,N_2417,N_2257);
xor U4967 (N_4967,N_2855,N_2324);
xor U4968 (N_4968,N_3588,N_2414);
nor U4969 (N_4969,N_2595,N_3713);
nand U4970 (N_4970,N_3057,N_2285);
nand U4971 (N_4971,N_2143,N_3966);
nand U4972 (N_4972,N_3251,N_2856);
and U4973 (N_4973,N_3314,N_2197);
or U4974 (N_4974,N_2307,N_3090);
nand U4975 (N_4975,N_3582,N_2936);
or U4976 (N_4976,N_3904,N_3164);
xor U4977 (N_4977,N_3209,N_3351);
or U4978 (N_4978,N_3917,N_2306);
or U4979 (N_4979,N_2506,N_3967);
xor U4980 (N_4980,N_2627,N_2141);
nor U4981 (N_4981,N_3081,N_2038);
nor U4982 (N_4982,N_3771,N_3107);
xor U4983 (N_4983,N_2711,N_2999);
or U4984 (N_4984,N_2243,N_2301);
nor U4985 (N_4985,N_2122,N_2898);
nand U4986 (N_4986,N_3498,N_3101);
or U4987 (N_4987,N_3261,N_3572);
nor U4988 (N_4988,N_2726,N_2688);
nor U4989 (N_4989,N_2360,N_2682);
or U4990 (N_4990,N_3547,N_3333);
and U4991 (N_4991,N_3943,N_3210);
xor U4992 (N_4992,N_3144,N_2070);
and U4993 (N_4993,N_2186,N_3096);
or U4994 (N_4994,N_2774,N_3630);
nor U4995 (N_4995,N_3225,N_2986);
or U4996 (N_4996,N_2395,N_2815);
nand U4997 (N_4997,N_2689,N_3371);
or U4998 (N_4998,N_3903,N_2617);
and U4999 (N_4999,N_3249,N_2929);
nor U5000 (N_5000,N_2359,N_3502);
or U5001 (N_5001,N_3324,N_3798);
nand U5002 (N_5002,N_3901,N_3151);
or U5003 (N_5003,N_3656,N_3883);
xor U5004 (N_5004,N_2197,N_3561);
or U5005 (N_5005,N_2721,N_3759);
or U5006 (N_5006,N_3674,N_3069);
xnor U5007 (N_5007,N_3850,N_3980);
nand U5008 (N_5008,N_2517,N_3357);
nand U5009 (N_5009,N_2779,N_3994);
and U5010 (N_5010,N_2544,N_3403);
or U5011 (N_5011,N_2682,N_3840);
xor U5012 (N_5012,N_2208,N_3407);
nand U5013 (N_5013,N_2446,N_3868);
nor U5014 (N_5014,N_3656,N_3592);
nor U5015 (N_5015,N_3814,N_3838);
xor U5016 (N_5016,N_3726,N_3699);
or U5017 (N_5017,N_3440,N_2847);
nand U5018 (N_5018,N_2976,N_2014);
nor U5019 (N_5019,N_2989,N_3639);
nand U5020 (N_5020,N_2080,N_3490);
nor U5021 (N_5021,N_2977,N_2615);
nor U5022 (N_5022,N_3507,N_2524);
nor U5023 (N_5023,N_3032,N_3490);
and U5024 (N_5024,N_3699,N_2170);
nand U5025 (N_5025,N_2186,N_3830);
nand U5026 (N_5026,N_2024,N_3015);
or U5027 (N_5027,N_2701,N_2243);
or U5028 (N_5028,N_3088,N_3981);
and U5029 (N_5029,N_3535,N_3926);
nor U5030 (N_5030,N_3532,N_2769);
nor U5031 (N_5031,N_3834,N_3156);
nand U5032 (N_5032,N_3472,N_3568);
xnor U5033 (N_5033,N_3203,N_2597);
and U5034 (N_5034,N_3013,N_3380);
or U5035 (N_5035,N_3049,N_3566);
xnor U5036 (N_5036,N_2544,N_3833);
nor U5037 (N_5037,N_2637,N_2971);
and U5038 (N_5038,N_3911,N_3870);
or U5039 (N_5039,N_3785,N_3781);
nand U5040 (N_5040,N_3459,N_2857);
and U5041 (N_5041,N_2360,N_3763);
or U5042 (N_5042,N_3425,N_3659);
nor U5043 (N_5043,N_3314,N_2846);
xor U5044 (N_5044,N_2813,N_3460);
nand U5045 (N_5045,N_2648,N_3037);
and U5046 (N_5046,N_2900,N_2144);
nor U5047 (N_5047,N_3314,N_2400);
xnor U5048 (N_5048,N_2611,N_3754);
or U5049 (N_5049,N_3177,N_3632);
nand U5050 (N_5050,N_2580,N_2780);
xnor U5051 (N_5051,N_3013,N_2834);
and U5052 (N_5052,N_2110,N_2562);
nand U5053 (N_5053,N_2132,N_3312);
or U5054 (N_5054,N_2548,N_3164);
xnor U5055 (N_5055,N_3085,N_2646);
and U5056 (N_5056,N_2553,N_3447);
or U5057 (N_5057,N_2995,N_2210);
nand U5058 (N_5058,N_2257,N_2817);
nand U5059 (N_5059,N_3076,N_3106);
and U5060 (N_5060,N_3462,N_2329);
nand U5061 (N_5061,N_3273,N_2059);
or U5062 (N_5062,N_3488,N_2896);
and U5063 (N_5063,N_2623,N_2323);
nor U5064 (N_5064,N_3527,N_2771);
or U5065 (N_5065,N_3951,N_3062);
xor U5066 (N_5066,N_2924,N_3485);
nor U5067 (N_5067,N_3388,N_3352);
nand U5068 (N_5068,N_2887,N_2039);
xnor U5069 (N_5069,N_2022,N_2573);
nand U5070 (N_5070,N_2390,N_2240);
or U5071 (N_5071,N_2121,N_3483);
nor U5072 (N_5072,N_3491,N_2177);
xor U5073 (N_5073,N_3832,N_3953);
nor U5074 (N_5074,N_3188,N_2578);
or U5075 (N_5075,N_2920,N_2930);
and U5076 (N_5076,N_3044,N_3738);
or U5077 (N_5077,N_3007,N_3748);
or U5078 (N_5078,N_2633,N_3006);
or U5079 (N_5079,N_2968,N_2258);
xor U5080 (N_5080,N_2385,N_3188);
nand U5081 (N_5081,N_3905,N_3379);
or U5082 (N_5082,N_3222,N_3924);
and U5083 (N_5083,N_3001,N_3196);
nor U5084 (N_5084,N_2951,N_3534);
or U5085 (N_5085,N_3288,N_3200);
nand U5086 (N_5086,N_2532,N_3106);
or U5087 (N_5087,N_2190,N_3623);
nand U5088 (N_5088,N_3065,N_3013);
nor U5089 (N_5089,N_2352,N_3797);
or U5090 (N_5090,N_2789,N_2123);
or U5091 (N_5091,N_3184,N_2193);
nor U5092 (N_5092,N_3863,N_2629);
and U5093 (N_5093,N_2939,N_2037);
nand U5094 (N_5094,N_3961,N_2934);
xnor U5095 (N_5095,N_3810,N_2181);
nor U5096 (N_5096,N_3192,N_2266);
nand U5097 (N_5097,N_3102,N_3123);
or U5098 (N_5098,N_3958,N_2423);
or U5099 (N_5099,N_2629,N_3285);
or U5100 (N_5100,N_2970,N_2891);
xor U5101 (N_5101,N_2901,N_3798);
nor U5102 (N_5102,N_3290,N_3843);
xor U5103 (N_5103,N_3084,N_3371);
and U5104 (N_5104,N_3184,N_2095);
xor U5105 (N_5105,N_2320,N_2565);
xor U5106 (N_5106,N_2892,N_2091);
or U5107 (N_5107,N_2121,N_2227);
xnor U5108 (N_5108,N_2949,N_2833);
nor U5109 (N_5109,N_2547,N_3965);
nand U5110 (N_5110,N_2849,N_3738);
nand U5111 (N_5111,N_2058,N_2856);
nor U5112 (N_5112,N_2691,N_3024);
xor U5113 (N_5113,N_2333,N_2677);
or U5114 (N_5114,N_3507,N_2945);
nor U5115 (N_5115,N_3026,N_2470);
nor U5116 (N_5116,N_2850,N_2647);
nor U5117 (N_5117,N_2904,N_2706);
nor U5118 (N_5118,N_3645,N_3572);
or U5119 (N_5119,N_3876,N_3967);
nor U5120 (N_5120,N_3596,N_2874);
or U5121 (N_5121,N_3528,N_3056);
or U5122 (N_5122,N_2527,N_3926);
nand U5123 (N_5123,N_3354,N_3349);
or U5124 (N_5124,N_2020,N_3060);
and U5125 (N_5125,N_2953,N_2081);
or U5126 (N_5126,N_3151,N_2310);
and U5127 (N_5127,N_3299,N_2116);
and U5128 (N_5128,N_2652,N_3570);
xor U5129 (N_5129,N_2834,N_2890);
nor U5130 (N_5130,N_2984,N_3273);
and U5131 (N_5131,N_2071,N_2012);
and U5132 (N_5132,N_2659,N_2151);
nand U5133 (N_5133,N_3606,N_2137);
nand U5134 (N_5134,N_2676,N_2621);
nor U5135 (N_5135,N_3771,N_3811);
or U5136 (N_5136,N_3227,N_3670);
and U5137 (N_5137,N_3277,N_2116);
nor U5138 (N_5138,N_3417,N_2938);
and U5139 (N_5139,N_2976,N_2362);
xor U5140 (N_5140,N_2422,N_2735);
nand U5141 (N_5141,N_3403,N_2956);
xnor U5142 (N_5142,N_3023,N_2970);
nor U5143 (N_5143,N_2473,N_3864);
nand U5144 (N_5144,N_2645,N_2271);
xnor U5145 (N_5145,N_3643,N_3086);
xnor U5146 (N_5146,N_2582,N_2337);
or U5147 (N_5147,N_3896,N_2104);
nand U5148 (N_5148,N_2660,N_2143);
xnor U5149 (N_5149,N_3583,N_3680);
xnor U5150 (N_5150,N_3039,N_3302);
nand U5151 (N_5151,N_3597,N_2398);
or U5152 (N_5152,N_3764,N_3958);
nand U5153 (N_5153,N_2548,N_2137);
or U5154 (N_5154,N_3390,N_3795);
or U5155 (N_5155,N_3985,N_2178);
nor U5156 (N_5156,N_3038,N_2287);
nor U5157 (N_5157,N_2322,N_3941);
nor U5158 (N_5158,N_3769,N_3215);
or U5159 (N_5159,N_2881,N_2015);
or U5160 (N_5160,N_3389,N_2834);
nor U5161 (N_5161,N_2929,N_3351);
nor U5162 (N_5162,N_2163,N_3224);
and U5163 (N_5163,N_3082,N_2041);
and U5164 (N_5164,N_3180,N_2010);
nor U5165 (N_5165,N_2666,N_3186);
nor U5166 (N_5166,N_3023,N_2294);
nor U5167 (N_5167,N_2690,N_2604);
xor U5168 (N_5168,N_3907,N_2375);
nor U5169 (N_5169,N_3694,N_2908);
nand U5170 (N_5170,N_3522,N_3133);
or U5171 (N_5171,N_2303,N_2309);
nor U5172 (N_5172,N_2715,N_2471);
xor U5173 (N_5173,N_2394,N_3315);
nand U5174 (N_5174,N_2674,N_3812);
and U5175 (N_5175,N_2275,N_3083);
or U5176 (N_5176,N_3324,N_2266);
or U5177 (N_5177,N_3638,N_3165);
nor U5178 (N_5178,N_2515,N_3655);
xnor U5179 (N_5179,N_2005,N_3669);
and U5180 (N_5180,N_3048,N_2967);
and U5181 (N_5181,N_2372,N_2641);
or U5182 (N_5182,N_2287,N_2492);
nand U5183 (N_5183,N_2188,N_3302);
or U5184 (N_5184,N_3288,N_2808);
nor U5185 (N_5185,N_2314,N_2549);
nand U5186 (N_5186,N_2754,N_3177);
and U5187 (N_5187,N_3546,N_2813);
nor U5188 (N_5188,N_3381,N_2993);
or U5189 (N_5189,N_3362,N_2345);
or U5190 (N_5190,N_3949,N_3488);
or U5191 (N_5191,N_3184,N_3933);
nand U5192 (N_5192,N_3479,N_3604);
and U5193 (N_5193,N_2352,N_2760);
or U5194 (N_5194,N_3006,N_3132);
or U5195 (N_5195,N_2010,N_3024);
or U5196 (N_5196,N_2812,N_2907);
and U5197 (N_5197,N_2418,N_2832);
and U5198 (N_5198,N_2644,N_3616);
nor U5199 (N_5199,N_2012,N_2047);
and U5200 (N_5200,N_2070,N_3462);
xnor U5201 (N_5201,N_2234,N_3289);
and U5202 (N_5202,N_2242,N_2957);
xnor U5203 (N_5203,N_2299,N_3007);
or U5204 (N_5204,N_2655,N_2007);
and U5205 (N_5205,N_3518,N_3432);
nand U5206 (N_5206,N_3325,N_3741);
nand U5207 (N_5207,N_2496,N_2614);
xnor U5208 (N_5208,N_3324,N_2849);
or U5209 (N_5209,N_2950,N_2756);
nand U5210 (N_5210,N_3587,N_3958);
or U5211 (N_5211,N_2367,N_2451);
nor U5212 (N_5212,N_3890,N_3451);
and U5213 (N_5213,N_3661,N_2604);
and U5214 (N_5214,N_3445,N_3740);
xnor U5215 (N_5215,N_3907,N_3940);
and U5216 (N_5216,N_3480,N_2962);
nand U5217 (N_5217,N_2454,N_2786);
nand U5218 (N_5218,N_2157,N_3633);
and U5219 (N_5219,N_2256,N_2213);
nor U5220 (N_5220,N_2264,N_2420);
nor U5221 (N_5221,N_2676,N_3063);
nand U5222 (N_5222,N_3544,N_3145);
xor U5223 (N_5223,N_2031,N_3844);
xor U5224 (N_5224,N_3201,N_2464);
nand U5225 (N_5225,N_2479,N_3950);
and U5226 (N_5226,N_2320,N_3569);
nand U5227 (N_5227,N_2820,N_2718);
nor U5228 (N_5228,N_2978,N_3660);
nor U5229 (N_5229,N_3797,N_2600);
or U5230 (N_5230,N_2827,N_2071);
or U5231 (N_5231,N_3601,N_3810);
nand U5232 (N_5232,N_2694,N_2007);
and U5233 (N_5233,N_3644,N_2318);
nand U5234 (N_5234,N_3185,N_2271);
xnor U5235 (N_5235,N_2802,N_2399);
nor U5236 (N_5236,N_3664,N_2035);
and U5237 (N_5237,N_3374,N_3946);
or U5238 (N_5238,N_2484,N_3084);
nor U5239 (N_5239,N_3761,N_3648);
or U5240 (N_5240,N_2972,N_2055);
and U5241 (N_5241,N_3063,N_2254);
or U5242 (N_5242,N_3043,N_2583);
xor U5243 (N_5243,N_3407,N_2207);
nand U5244 (N_5244,N_2411,N_2791);
nand U5245 (N_5245,N_2014,N_3761);
or U5246 (N_5246,N_3901,N_2267);
and U5247 (N_5247,N_2805,N_2957);
nor U5248 (N_5248,N_3720,N_3471);
xnor U5249 (N_5249,N_3408,N_2442);
nor U5250 (N_5250,N_2945,N_3757);
nor U5251 (N_5251,N_2869,N_3833);
xnor U5252 (N_5252,N_3886,N_3499);
or U5253 (N_5253,N_3801,N_2479);
or U5254 (N_5254,N_3541,N_2959);
or U5255 (N_5255,N_2182,N_3770);
and U5256 (N_5256,N_2817,N_3234);
nor U5257 (N_5257,N_2717,N_2426);
xor U5258 (N_5258,N_2358,N_2043);
nand U5259 (N_5259,N_2788,N_3034);
nand U5260 (N_5260,N_3465,N_3450);
nor U5261 (N_5261,N_2649,N_3556);
and U5262 (N_5262,N_3169,N_2528);
and U5263 (N_5263,N_3294,N_3181);
nand U5264 (N_5264,N_3389,N_3357);
nand U5265 (N_5265,N_3768,N_2921);
xor U5266 (N_5266,N_3463,N_3380);
and U5267 (N_5267,N_3571,N_3418);
or U5268 (N_5268,N_3435,N_3159);
and U5269 (N_5269,N_3363,N_3877);
xnor U5270 (N_5270,N_3884,N_3017);
xnor U5271 (N_5271,N_3700,N_2293);
or U5272 (N_5272,N_2213,N_2559);
or U5273 (N_5273,N_2961,N_2258);
xnor U5274 (N_5274,N_3084,N_3551);
nand U5275 (N_5275,N_2449,N_3218);
xor U5276 (N_5276,N_2445,N_2232);
or U5277 (N_5277,N_3697,N_2278);
or U5278 (N_5278,N_2797,N_3161);
nand U5279 (N_5279,N_3388,N_2271);
nand U5280 (N_5280,N_3344,N_3420);
or U5281 (N_5281,N_3347,N_3510);
and U5282 (N_5282,N_2490,N_3665);
and U5283 (N_5283,N_3583,N_2251);
or U5284 (N_5284,N_3551,N_2066);
and U5285 (N_5285,N_2405,N_3422);
or U5286 (N_5286,N_2524,N_2938);
or U5287 (N_5287,N_3338,N_3931);
nand U5288 (N_5288,N_2163,N_3675);
nor U5289 (N_5289,N_2466,N_3544);
or U5290 (N_5290,N_2374,N_2774);
and U5291 (N_5291,N_3662,N_2693);
xor U5292 (N_5292,N_2849,N_2046);
xor U5293 (N_5293,N_3337,N_3924);
or U5294 (N_5294,N_2595,N_3327);
nand U5295 (N_5295,N_2116,N_2942);
nor U5296 (N_5296,N_2774,N_3044);
xor U5297 (N_5297,N_3253,N_2574);
nor U5298 (N_5298,N_2241,N_2276);
or U5299 (N_5299,N_3313,N_3227);
or U5300 (N_5300,N_3990,N_3629);
nand U5301 (N_5301,N_3203,N_3657);
xnor U5302 (N_5302,N_3055,N_3368);
and U5303 (N_5303,N_3256,N_2923);
xnor U5304 (N_5304,N_2075,N_3375);
and U5305 (N_5305,N_2341,N_3982);
nand U5306 (N_5306,N_3832,N_3743);
nand U5307 (N_5307,N_2967,N_3597);
nand U5308 (N_5308,N_3100,N_2355);
or U5309 (N_5309,N_2677,N_3787);
nor U5310 (N_5310,N_3061,N_2274);
nand U5311 (N_5311,N_2126,N_2381);
xor U5312 (N_5312,N_3861,N_3938);
xor U5313 (N_5313,N_3306,N_3918);
and U5314 (N_5314,N_2945,N_3358);
and U5315 (N_5315,N_2078,N_2621);
or U5316 (N_5316,N_3903,N_3325);
or U5317 (N_5317,N_2117,N_3982);
xor U5318 (N_5318,N_3311,N_3383);
or U5319 (N_5319,N_2281,N_2534);
or U5320 (N_5320,N_2869,N_2122);
or U5321 (N_5321,N_3591,N_2675);
and U5322 (N_5322,N_3785,N_2465);
or U5323 (N_5323,N_3916,N_2665);
and U5324 (N_5324,N_2318,N_3256);
or U5325 (N_5325,N_2271,N_3290);
nor U5326 (N_5326,N_2402,N_2658);
or U5327 (N_5327,N_2451,N_3046);
or U5328 (N_5328,N_2386,N_2009);
and U5329 (N_5329,N_3088,N_2958);
and U5330 (N_5330,N_3792,N_3467);
nand U5331 (N_5331,N_3459,N_2008);
nand U5332 (N_5332,N_2521,N_2717);
nand U5333 (N_5333,N_2237,N_3728);
and U5334 (N_5334,N_3201,N_2207);
nor U5335 (N_5335,N_3437,N_3823);
or U5336 (N_5336,N_2919,N_3131);
and U5337 (N_5337,N_2947,N_3581);
nor U5338 (N_5338,N_2677,N_2952);
nor U5339 (N_5339,N_3199,N_2720);
nor U5340 (N_5340,N_3338,N_2598);
or U5341 (N_5341,N_3212,N_2290);
xnor U5342 (N_5342,N_3100,N_3435);
nand U5343 (N_5343,N_2812,N_3602);
or U5344 (N_5344,N_2162,N_3884);
or U5345 (N_5345,N_3843,N_3696);
nand U5346 (N_5346,N_3217,N_2131);
nor U5347 (N_5347,N_2500,N_3032);
and U5348 (N_5348,N_3070,N_3410);
nor U5349 (N_5349,N_2939,N_2138);
or U5350 (N_5350,N_3471,N_2687);
and U5351 (N_5351,N_3843,N_3826);
nand U5352 (N_5352,N_2789,N_2645);
nand U5353 (N_5353,N_2274,N_3701);
or U5354 (N_5354,N_3680,N_3979);
or U5355 (N_5355,N_3183,N_3948);
nor U5356 (N_5356,N_3812,N_2714);
nand U5357 (N_5357,N_2131,N_3111);
nor U5358 (N_5358,N_2992,N_2030);
and U5359 (N_5359,N_3944,N_3261);
nor U5360 (N_5360,N_2029,N_3605);
or U5361 (N_5361,N_2785,N_3670);
nor U5362 (N_5362,N_2663,N_3542);
xnor U5363 (N_5363,N_3784,N_3642);
nand U5364 (N_5364,N_3622,N_3901);
xnor U5365 (N_5365,N_3621,N_3826);
xor U5366 (N_5366,N_3320,N_2125);
or U5367 (N_5367,N_2677,N_2154);
nor U5368 (N_5368,N_3583,N_3505);
and U5369 (N_5369,N_3849,N_3638);
and U5370 (N_5370,N_2425,N_3123);
nor U5371 (N_5371,N_3534,N_3491);
and U5372 (N_5372,N_2566,N_3466);
nor U5373 (N_5373,N_3079,N_2226);
and U5374 (N_5374,N_3264,N_2705);
nor U5375 (N_5375,N_3897,N_3918);
nand U5376 (N_5376,N_2371,N_2339);
and U5377 (N_5377,N_3090,N_3054);
nand U5378 (N_5378,N_2302,N_3431);
or U5379 (N_5379,N_2320,N_2573);
nand U5380 (N_5380,N_3028,N_3902);
nor U5381 (N_5381,N_2353,N_3141);
or U5382 (N_5382,N_3317,N_3153);
and U5383 (N_5383,N_2066,N_2976);
or U5384 (N_5384,N_2477,N_3463);
nand U5385 (N_5385,N_3712,N_3767);
nor U5386 (N_5386,N_2946,N_2409);
xnor U5387 (N_5387,N_2825,N_3465);
nand U5388 (N_5388,N_3068,N_3435);
nor U5389 (N_5389,N_2671,N_3987);
xor U5390 (N_5390,N_2092,N_3762);
nor U5391 (N_5391,N_2319,N_3626);
or U5392 (N_5392,N_3008,N_3006);
or U5393 (N_5393,N_3088,N_2745);
nor U5394 (N_5394,N_3748,N_2239);
or U5395 (N_5395,N_3982,N_3357);
xor U5396 (N_5396,N_3958,N_3202);
or U5397 (N_5397,N_2461,N_3059);
or U5398 (N_5398,N_2929,N_2679);
and U5399 (N_5399,N_3979,N_3612);
nor U5400 (N_5400,N_2848,N_2056);
and U5401 (N_5401,N_3371,N_2826);
xor U5402 (N_5402,N_2085,N_3004);
xor U5403 (N_5403,N_2654,N_2433);
nor U5404 (N_5404,N_2204,N_3194);
nand U5405 (N_5405,N_2445,N_3764);
or U5406 (N_5406,N_2137,N_2090);
or U5407 (N_5407,N_2872,N_2879);
or U5408 (N_5408,N_3184,N_2292);
or U5409 (N_5409,N_3092,N_2509);
and U5410 (N_5410,N_3683,N_3865);
nor U5411 (N_5411,N_2110,N_3993);
nor U5412 (N_5412,N_3764,N_3517);
nor U5413 (N_5413,N_3409,N_3060);
or U5414 (N_5414,N_3493,N_2396);
or U5415 (N_5415,N_2029,N_3110);
nand U5416 (N_5416,N_3490,N_2952);
nor U5417 (N_5417,N_3184,N_2315);
and U5418 (N_5418,N_2037,N_2388);
and U5419 (N_5419,N_3005,N_2182);
or U5420 (N_5420,N_3168,N_2186);
and U5421 (N_5421,N_3906,N_2941);
nor U5422 (N_5422,N_2242,N_2088);
nand U5423 (N_5423,N_3981,N_2825);
or U5424 (N_5424,N_2497,N_3811);
or U5425 (N_5425,N_3049,N_3011);
nand U5426 (N_5426,N_3636,N_2363);
or U5427 (N_5427,N_3208,N_3841);
xnor U5428 (N_5428,N_3754,N_3719);
nand U5429 (N_5429,N_3894,N_3331);
xor U5430 (N_5430,N_3779,N_2165);
xnor U5431 (N_5431,N_2325,N_3439);
nor U5432 (N_5432,N_2419,N_2112);
nor U5433 (N_5433,N_3799,N_3532);
nand U5434 (N_5434,N_2501,N_3140);
and U5435 (N_5435,N_2030,N_3904);
or U5436 (N_5436,N_2311,N_2730);
xnor U5437 (N_5437,N_3680,N_3064);
or U5438 (N_5438,N_3846,N_2894);
or U5439 (N_5439,N_2220,N_3320);
and U5440 (N_5440,N_3873,N_3218);
nand U5441 (N_5441,N_3462,N_3976);
nor U5442 (N_5442,N_3640,N_3765);
nor U5443 (N_5443,N_3710,N_2207);
and U5444 (N_5444,N_3755,N_2212);
nor U5445 (N_5445,N_3905,N_3931);
nor U5446 (N_5446,N_3287,N_2338);
xnor U5447 (N_5447,N_2185,N_2525);
nor U5448 (N_5448,N_3661,N_3796);
nor U5449 (N_5449,N_2653,N_2446);
nor U5450 (N_5450,N_3094,N_2212);
xor U5451 (N_5451,N_2096,N_3799);
and U5452 (N_5452,N_3585,N_2884);
or U5453 (N_5453,N_3970,N_3873);
xor U5454 (N_5454,N_3855,N_3368);
nor U5455 (N_5455,N_2632,N_2470);
nor U5456 (N_5456,N_2632,N_3942);
nand U5457 (N_5457,N_2909,N_2958);
nor U5458 (N_5458,N_3701,N_3288);
xor U5459 (N_5459,N_2547,N_2669);
nor U5460 (N_5460,N_2524,N_3988);
or U5461 (N_5461,N_3871,N_3761);
nor U5462 (N_5462,N_3468,N_3594);
xnor U5463 (N_5463,N_3400,N_2448);
or U5464 (N_5464,N_3888,N_3272);
nand U5465 (N_5465,N_2415,N_2069);
nor U5466 (N_5466,N_3008,N_2017);
xnor U5467 (N_5467,N_2303,N_3829);
nor U5468 (N_5468,N_3458,N_3676);
nor U5469 (N_5469,N_2932,N_3232);
nor U5470 (N_5470,N_2680,N_2971);
xnor U5471 (N_5471,N_3358,N_2506);
nand U5472 (N_5472,N_2909,N_2315);
nand U5473 (N_5473,N_3280,N_3316);
nand U5474 (N_5474,N_2825,N_3364);
nor U5475 (N_5475,N_3409,N_3642);
nor U5476 (N_5476,N_2075,N_3827);
xnor U5477 (N_5477,N_3930,N_3276);
nand U5478 (N_5478,N_3983,N_3241);
and U5479 (N_5479,N_3108,N_2046);
xnor U5480 (N_5480,N_3199,N_2370);
xnor U5481 (N_5481,N_3988,N_3180);
nor U5482 (N_5482,N_3445,N_2555);
nor U5483 (N_5483,N_2888,N_3132);
nand U5484 (N_5484,N_2698,N_2513);
xnor U5485 (N_5485,N_2245,N_2859);
and U5486 (N_5486,N_3161,N_3813);
xnor U5487 (N_5487,N_2431,N_3909);
and U5488 (N_5488,N_3762,N_3013);
or U5489 (N_5489,N_3221,N_3372);
nand U5490 (N_5490,N_2375,N_2253);
nand U5491 (N_5491,N_2634,N_2506);
nand U5492 (N_5492,N_2765,N_2035);
or U5493 (N_5493,N_3720,N_2392);
or U5494 (N_5494,N_3922,N_2833);
and U5495 (N_5495,N_2839,N_2778);
nand U5496 (N_5496,N_2520,N_2590);
or U5497 (N_5497,N_2858,N_3040);
and U5498 (N_5498,N_3989,N_2478);
xor U5499 (N_5499,N_3874,N_3796);
nor U5500 (N_5500,N_2276,N_2777);
nand U5501 (N_5501,N_2489,N_3733);
or U5502 (N_5502,N_3876,N_2246);
nor U5503 (N_5503,N_2991,N_2195);
xor U5504 (N_5504,N_2590,N_2803);
and U5505 (N_5505,N_2472,N_2585);
nand U5506 (N_5506,N_3334,N_3148);
and U5507 (N_5507,N_2788,N_2880);
nor U5508 (N_5508,N_3534,N_2947);
or U5509 (N_5509,N_3555,N_2595);
or U5510 (N_5510,N_2260,N_3448);
or U5511 (N_5511,N_3498,N_3751);
nor U5512 (N_5512,N_3091,N_3048);
nor U5513 (N_5513,N_2058,N_2125);
nand U5514 (N_5514,N_3785,N_2747);
nand U5515 (N_5515,N_2020,N_2995);
nand U5516 (N_5516,N_2038,N_2507);
xor U5517 (N_5517,N_3683,N_3470);
nor U5518 (N_5518,N_3029,N_3134);
xnor U5519 (N_5519,N_2956,N_3427);
nor U5520 (N_5520,N_3736,N_3576);
nand U5521 (N_5521,N_2523,N_3448);
or U5522 (N_5522,N_2767,N_3923);
nor U5523 (N_5523,N_3336,N_2524);
nor U5524 (N_5524,N_2087,N_2570);
and U5525 (N_5525,N_3618,N_2720);
and U5526 (N_5526,N_3259,N_2477);
nand U5527 (N_5527,N_2095,N_3146);
and U5528 (N_5528,N_3176,N_2573);
or U5529 (N_5529,N_3154,N_3810);
nand U5530 (N_5530,N_3574,N_3001);
and U5531 (N_5531,N_3779,N_3737);
or U5532 (N_5532,N_3751,N_2168);
or U5533 (N_5533,N_2787,N_3426);
and U5534 (N_5534,N_2742,N_2635);
nand U5535 (N_5535,N_3489,N_2088);
or U5536 (N_5536,N_3602,N_3550);
and U5537 (N_5537,N_3904,N_2072);
or U5538 (N_5538,N_2923,N_2702);
or U5539 (N_5539,N_2013,N_2683);
nand U5540 (N_5540,N_2914,N_3200);
nor U5541 (N_5541,N_3014,N_3371);
nand U5542 (N_5542,N_2119,N_2124);
or U5543 (N_5543,N_3737,N_3040);
nand U5544 (N_5544,N_3468,N_2847);
or U5545 (N_5545,N_3512,N_2446);
xnor U5546 (N_5546,N_2417,N_3951);
nor U5547 (N_5547,N_2998,N_3118);
xnor U5548 (N_5548,N_3434,N_2126);
xor U5549 (N_5549,N_3649,N_3121);
nor U5550 (N_5550,N_3068,N_2622);
nor U5551 (N_5551,N_2439,N_2028);
and U5552 (N_5552,N_2086,N_2384);
or U5553 (N_5553,N_3817,N_2125);
or U5554 (N_5554,N_2258,N_2213);
nand U5555 (N_5555,N_2937,N_2984);
nand U5556 (N_5556,N_3592,N_2169);
nor U5557 (N_5557,N_3834,N_3479);
nand U5558 (N_5558,N_3335,N_2496);
or U5559 (N_5559,N_3757,N_2202);
xor U5560 (N_5560,N_2786,N_2764);
and U5561 (N_5561,N_3455,N_2794);
xor U5562 (N_5562,N_3172,N_2865);
or U5563 (N_5563,N_2794,N_2467);
and U5564 (N_5564,N_3031,N_2007);
or U5565 (N_5565,N_3433,N_3878);
or U5566 (N_5566,N_2237,N_3897);
xnor U5567 (N_5567,N_3148,N_2957);
or U5568 (N_5568,N_2107,N_3782);
nand U5569 (N_5569,N_2585,N_2527);
nand U5570 (N_5570,N_3737,N_3072);
xnor U5571 (N_5571,N_3582,N_2685);
xor U5572 (N_5572,N_3793,N_3084);
nand U5573 (N_5573,N_3231,N_2376);
or U5574 (N_5574,N_3490,N_2521);
nand U5575 (N_5575,N_3001,N_3408);
xnor U5576 (N_5576,N_3022,N_3899);
xnor U5577 (N_5577,N_2516,N_3615);
or U5578 (N_5578,N_3166,N_2666);
or U5579 (N_5579,N_3671,N_3830);
or U5580 (N_5580,N_2854,N_2306);
xor U5581 (N_5581,N_3454,N_2513);
nand U5582 (N_5582,N_2445,N_2225);
or U5583 (N_5583,N_3602,N_2967);
nand U5584 (N_5584,N_3239,N_2318);
and U5585 (N_5585,N_3308,N_3939);
or U5586 (N_5586,N_3386,N_2137);
xnor U5587 (N_5587,N_2201,N_3755);
xor U5588 (N_5588,N_3983,N_2237);
nand U5589 (N_5589,N_2194,N_2957);
nand U5590 (N_5590,N_3028,N_2282);
or U5591 (N_5591,N_2118,N_3493);
and U5592 (N_5592,N_3370,N_2506);
or U5593 (N_5593,N_2388,N_2352);
nor U5594 (N_5594,N_3371,N_2547);
or U5595 (N_5595,N_2523,N_2964);
nand U5596 (N_5596,N_2954,N_2413);
or U5597 (N_5597,N_2289,N_2284);
and U5598 (N_5598,N_3239,N_3816);
nand U5599 (N_5599,N_3242,N_3397);
nand U5600 (N_5600,N_2651,N_2608);
nand U5601 (N_5601,N_2265,N_2154);
nand U5602 (N_5602,N_3785,N_3724);
and U5603 (N_5603,N_3828,N_3693);
xnor U5604 (N_5604,N_2398,N_2669);
and U5605 (N_5605,N_3545,N_3463);
or U5606 (N_5606,N_2678,N_3404);
nand U5607 (N_5607,N_3459,N_2651);
xnor U5608 (N_5608,N_2240,N_3842);
nor U5609 (N_5609,N_3551,N_3307);
xnor U5610 (N_5610,N_3782,N_2295);
and U5611 (N_5611,N_2548,N_3698);
and U5612 (N_5612,N_2931,N_3591);
xor U5613 (N_5613,N_2689,N_2707);
nand U5614 (N_5614,N_2121,N_2166);
nand U5615 (N_5615,N_3227,N_2774);
nor U5616 (N_5616,N_3332,N_3132);
or U5617 (N_5617,N_3502,N_3284);
nor U5618 (N_5618,N_3141,N_2079);
xor U5619 (N_5619,N_2485,N_2282);
and U5620 (N_5620,N_3224,N_3310);
or U5621 (N_5621,N_2323,N_2562);
or U5622 (N_5622,N_3944,N_2223);
nor U5623 (N_5623,N_3970,N_2733);
nand U5624 (N_5624,N_3128,N_2127);
nand U5625 (N_5625,N_3147,N_2089);
xor U5626 (N_5626,N_3934,N_2168);
xnor U5627 (N_5627,N_3716,N_3437);
nand U5628 (N_5628,N_2393,N_2225);
or U5629 (N_5629,N_2614,N_2133);
nand U5630 (N_5630,N_2003,N_3738);
nand U5631 (N_5631,N_3694,N_3171);
nor U5632 (N_5632,N_3347,N_2069);
xor U5633 (N_5633,N_2486,N_3576);
or U5634 (N_5634,N_2343,N_2082);
or U5635 (N_5635,N_3642,N_3231);
nor U5636 (N_5636,N_2115,N_2964);
nand U5637 (N_5637,N_3472,N_3125);
nor U5638 (N_5638,N_2081,N_3444);
nand U5639 (N_5639,N_3301,N_2625);
or U5640 (N_5640,N_3740,N_2745);
and U5641 (N_5641,N_2260,N_3178);
xor U5642 (N_5642,N_3042,N_3442);
and U5643 (N_5643,N_2985,N_3398);
nor U5644 (N_5644,N_3286,N_2495);
nand U5645 (N_5645,N_3558,N_3506);
nor U5646 (N_5646,N_3524,N_3556);
nand U5647 (N_5647,N_2135,N_3784);
xnor U5648 (N_5648,N_2025,N_2948);
nor U5649 (N_5649,N_3455,N_3786);
xnor U5650 (N_5650,N_3902,N_3686);
or U5651 (N_5651,N_3491,N_2531);
or U5652 (N_5652,N_2920,N_3928);
and U5653 (N_5653,N_2920,N_2531);
nor U5654 (N_5654,N_2609,N_2061);
and U5655 (N_5655,N_3799,N_2463);
xor U5656 (N_5656,N_3555,N_3910);
and U5657 (N_5657,N_3829,N_2487);
nor U5658 (N_5658,N_3122,N_2057);
or U5659 (N_5659,N_2921,N_3232);
or U5660 (N_5660,N_2179,N_2238);
xnor U5661 (N_5661,N_3100,N_2036);
or U5662 (N_5662,N_2201,N_3359);
and U5663 (N_5663,N_2232,N_2375);
or U5664 (N_5664,N_2180,N_3834);
nand U5665 (N_5665,N_3689,N_2380);
xnor U5666 (N_5666,N_3344,N_2785);
and U5667 (N_5667,N_3775,N_3719);
or U5668 (N_5668,N_3778,N_3087);
nor U5669 (N_5669,N_3648,N_2141);
nand U5670 (N_5670,N_3591,N_3534);
or U5671 (N_5671,N_2668,N_3945);
xor U5672 (N_5672,N_3477,N_2033);
nor U5673 (N_5673,N_3572,N_2447);
nand U5674 (N_5674,N_2757,N_2201);
xor U5675 (N_5675,N_3480,N_3929);
nor U5676 (N_5676,N_3121,N_2152);
nand U5677 (N_5677,N_3376,N_2443);
xor U5678 (N_5678,N_3571,N_2472);
nand U5679 (N_5679,N_3161,N_3461);
and U5680 (N_5680,N_3806,N_2276);
and U5681 (N_5681,N_2590,N_2613);
nand U5682 (N_5682,N_3477,N_2403);
nand U5683 (N_5683,N_3190,N_2919);
or U5684 (N_5684,N_2698,N_3206);
nor U5685 (N_5685,N_3504,N_2019);
xnor U5686 (N_5686,N_2719,N_2124);
and U5687 (N_5687,N_3874,N_2702);
and U5688 (N_5688,N_2770,N_3791);
or U5689 (N_5689,N_2030,N_3447);
or U5690 (N_5690,N_2951,N_2198);
nand U5691 (N_5691,N_2718,N_3232);
nor U5692 (N_5692,N_3343,N_2055);
and U5693 (N_5693,N_2633,N_3771);
xor U5694 (N_5694,N_2647,N_2686);
nand U5695 (N_5695,N_3235,N_2259);
and U5696 (N_5696,N_2949,N_3699);
nand U5697 (N_5697,N_3040,N_3772);
and U5698 (N_5698,N_2234,N_3940);
or U5699 (N_5699,N_3768,N_3684);
xor U5700 (N_5700,N_3363,N_2346);
nor U5701 (N_5701,N_3668,N_3637);
nand U5702 (N_5702,N_2358,N_3220);
and U5703 (N_5703,N_2782,N_3436);
xnor U5704 (N_5704,N_2310,N_3153);
xnor U5705 (N_5705,N_3412,N_2996);
and U5706 (N_5706,N_2343,N_3816);
xnor U5707 (N_5707,N_2193,N_3053);
and U5708 (N_5708,N_2782,N_2984);
xnor U5709 (N_5709,N_3213,N_3549);
and U5710 (N_5710,N_2168,N_2322);
nor U5711 (N_5711,N_3711,N_3040);
and U5712 (N_5712,N_2707,N_3458);
nand U5713 (N_5713,N_3277,N_2791);
nand U5714 (N_5714,N_3664,N_3772);
and U5715 (N_5715,N_3047,N_3447);
xor U5716 (N_5716,N_3947,N_3908);
xor U5717 (N_5717,N_3811,N_2595);
nor U5718 (N_5718,N_3843,N_2141);
and U5719 (N_5719,N_2698,N_2254);
xor U5720 (N_5720,N_3349,N_2954);
xnor U5721 (N_5721,N_2218,N_2055);
nor U5722 (N_5722,N_3821,N_2401);
nand U5723 (N_5723,N_2283,N_3819);
and U5724 (N_5724,N_3094,N_2015);
xor U5725 (N_5725,N_3713,N_2829);
nand U5726 (N_5726,N_3381,N_2221);
and U5727 (N_5727,N_3359,N_2554);
nand U5728 (N_5728,N_3326,N_2154);
or U5729 (N_5729,N_3930,N_3158);
nand U5730 (N_5730,N_3586,N_3242);
nor U5731 (N_5731,N_3658,N_3843);
or U5732 (N_5732,N_2535,N_2054);
or U5733 (N_5733,N_3146,N_2530);
xor U5734 (N_5734,N_2863,N_3330);
nor U5735 (N_5735,N_2695,N_2572);
or U5736 (N_5736,N_3268,N_3680);
or U5737 (N_5737,N_2675,N_2175);
nand U5738 (N_5738,N_3896,N_2090);
nor U5739 (N_5739,N_2632,N_2832);
and U5740 (N_5740,N_3712,N_2451);
and U5741 (N_5741,N_3107,N_3499);
xnor U5742 (N_5742,N_3565,N_2610);
nor U5743 (N_5743,N_3923,N_3924);
or U5744 (N_5744,N_3802,N_3623);
xnor U5745 (N_5745,N_3058,N_3148);
or U5746 (N_5746,N_2140,N_3484);
nand U5747 (N_5747,N_3995,N_2952);
nand U5748 (N_5748,N_3917,N_3213);
xor U5749 (N_5749,N_3104,N_2538);
and U5750 (N_5750,N_3675,N_3347);
and U5751 (N_5751,N_3274,N_2286);
nor U5752 (N_5752,N_3385,N_2690);
nor U5753 (N_5753,N_2270,N_2754);
nand U5754 (N_5754,N_3602,N_2393);
nor U5755 (N_5755,N_2803,N_2862);
or U5756 (N_5756,N_3365,N_3862);
or U5757 (N_5757,N_2216,N_3543);
nand U5758 (N_5758,N_3320,N_3669);
xor U5759 (N_5759,N_3436,N_3380);
and U5760 (N_5760,N_2501,N_2623);
or U5761 (N_5761,N_2338,N_2374);
or U5762 (N_5762,N_2199,N_2763);
nand U5763 (N_5763,N_2786,N_3233);
and U5764 (N_5764,N_2884,N_3354);
and U5765 (N_5765,N_3963,N_2138);
nor U5766 (N_5766,N_2401,N_2570);
nor U5767 (N_5767,N_2780,N_3254);
nand U5768 (N_5768,N_2897,N_2167);
nand U5769 (N_5769,N_2602,N_2277);
xnor U5770 (N_5770,N_2941,N_3932);
or U5771 (N_5771,N_3338,N_2050);
nand U5772 (N_5772,N_3941,N_3824);
nor U5773 (N_5773,N_3985,N_3340);
xor U5774 (N_5774,N_3066,N_3248);
or U5775 (N_5775,N_2604,N_2454);
nand U5776 (N_5776,N_3701,N_3898);
and U5777 (N_5777,N_2615,N_2244);
and U5778 (N_5778,N_2068,N_3821);
and U5779 (N_5779,N_2298,N_2630);
and U5780 (N_5780,N_3978,N_3954);
and U5781 (N_5781,N_2761,N_2011);
or U5782 (N_5782,N_3597,N_3931);
xor U5783 (N_5783,N_3274,N_3132);
nor U5784 (N_5784,N_2779,N_2137);
xor U5785 (N_5785,N_2507,N_2665);
xnor U5786 (N_5786,N_2062,N_3570);
xor U5787 (N_5787,N_2175,N_2648);
xnor U5788 (N_5788,N_2315,N_2106);
nor U5789 (N_5789,N_3879,N_2471);
and U5790 (N_5790,N_2695,N_2915);
xor U5791 (N_5791,N_2445,N_3049);
xnor U5792 (N_5792,N_3200,N_3266);
or U5793 (N_5793,N_2487,N_2741);
or U5794 (N_5794,N_2580,N_2363);
and U5795 (N_5795,N_3991,N_2245);
or U5796 (N_5796,N_2279,N_2899);
or U5797 (N_5797,N_2845,N_3123);
or U5798 (N_5798,N_2200,N_3206);
and U5799 (N_5799,N_3393,N_3132);
or U5800 (N_5800,N_3898,N_2792);
nor U5801 (N_5801,N_2466,N_3045);
xor U5802 (N_5802,N_2030,N_3244);
nand U5803 (N_5803,N_2643,N_3169);
xnor U5804 (N_5804,N_2559,N_3848);
nor U5805 (N_5805,N_3159,N_3887);
and U5806 (N_5806,N_2165,N_3056);
or U5807 (N_5807,N_2874,N_2101);
and U5808 (N_5808,N_3672,N_2775);
nor U5809 (N_5809,N_3146,N_2944);
nor U5810 (N_5810,N_2677,N_2068);
nor U5811 (N_5811,N_3820,N_3668);
xor U5812 (N_5812,N_3168,N_3772);
nor U5813 (N_5813,N_3592,N_2435);
nand U5814 (N_5814,N_2876,N_2720);
xor U5815 (N_5815,N_3738,N_3074);
or U5816 (N_5816,N_2934,N_2459);
xor U5817 (N_5817,N_3979,N_2558);
nor U5818 (N_5818,N_3533,N_3568);
xor U5819 (N_5819,N_2023,N_2897);
nand U5820 (N_5820,N_3316,N_2894);
or U5821 (N_5821,N_2182,N_3976);
nor U5822 (N_5822,N_3960,N_2677);
and U5823 (N_5823,N_3290,N_3181);
and U5824 (N_5824,N_2069,N_2983);
or U5825 (N_5825,N_3556,N_2917);
or U5826 (N_5826,N_3255,N_2987);
xnor U5827 (N_5827,N_2955,N_2794);
nor U5828 (N_5828,N_2292,N_2225);
nand U5829 (N_5829,N_2843,N_2445);
xor U5830 (N_5830,N_2070,N_2528);
nand U5831 (N_5831,N_3135,N_2272);
or U5832 (N_5832,N_2633,N_2207);
nand U5833 (N_5833,N_2370,N_3610);
nand U5834 (N_5834,N_2224,N_3870);
xor U5835 (N_5835,N_3203,N_2984);
xor U5836 (N_5836,N_2027,N_3021);
xnor U5837 (N_5837,N_3786,N_3761);
nor U5838 (N_5838,N_2314,N_3691);
and U5839 (N_5839,N_2877,N_2235);
nor U5840 (N_5840,N_2993,N_3301);
or U5841 (N_5841,N_3304,N_2420);
xnor U5842 (N_5842,N_3961,N_3955);
and U5843 (N_5843,N_3330,N_2459);
and U5844 (N_5844,N_3343,N_2818);
nor U5845 (N_5845,N_3215,N_2905);
or U5846 (N_5846,N_2488,N_2669);
nor U5847 (N_5847,N_3871,N_3558);
or U5848 (N_5848,N_2700,N_3251);
nor U5849 (N_5849,N_2469,N_3741);
nor U5850 (N_5850,N_2996,N_2981);
or U5851 (N_5851,N_3108,N_3278);
xor U5852 (N_5852,N_3494,N_2027);
or U5853 (N_5853,N_2545,N_2196);
or U5854 (N_5854,N_3912,N_3290);
or U5855 (N_5855,N_3305,N_2358);
or U5856 (N_5856,N_3560,N_2032);
nor U5857 (N_5857,N_3310,N_3902);
nor U5858 (N_5858,N_2521,N_2379);
nor U5859 (N_5859,N_2690,N_3825);
xnor U5860 (N_5860,N_3045,N_3925);
and U5861 (N_5861,N_3315,N_2633);
nor U5862 (N_5862,N_3089,N_3449);
nand U5863 (N_5863,N_3991,N_2677);
or U5864 (N_5864,N_2913,N_3831);
nand U5865 (N_5865,N_3655,N_3424);
xnor U5866 (N_5866,N_2242,N_2319);
nand U5867 (N_5867,N_3964,N_2285);
nor U5868 (N_5868,N_2405,N_2986);
xnor U5869 (N_5869,N_2223,N_3590);
xor U5870 (N_5870,N_3922,N_3485);
and U5871 (N_5871,N_3353,N_3182);
nand U5872 (N_5872,N_2743,N_2955);
nand U5873 (N_5873,N_3577,N_2138);
nor U5874 (N_5874,N_3579,N_3271);
and U5875 (N_5875,N_2034,N_2548);
and U5876 (N_5876,N_3605,N_3028);
nand U5877 (N_5877,N_2286,N_3980);
xnor U5878 (N_5878,N_3935,N_3003);
xnor U5879 (N_5879,N_3730,N_3446);
nor U5880 (N_5880,N_2594,N_3055);
nor U5881 (N_5881,N_3613,N_3998);
and U5882 (N_5882,N_2815,N_3072);
xor U5883 (N_5883,N_2776,N_3810);
nor U5884 (N_5884,N_3790,N_3875);
or U5885 (N_5885,N_3942,N_3871);
and U5886 (N_5886,N_3126,N_3911);
xor U5887 (N_5887,N_3998,N_3221);
xnor U5888 (N_5888,N_3561,N_3044);
and U5889 (N_5889,N_3429,N_2686);
nor U5890 (N_5890,N_3038,N_2642);
nand U5891 (N_5891,N_3277,N_2977);
nand U5892 (N_5892,N_2376,N_2214);
xnor U5893 (N_5893,N_2047,N_3082);
nand U5894 (N_5894,N_2453,N_2832);
or U5895 (N_5895,N_2416,N_2587);
nor U5896 (N_5896,N_2817,N_2069);
nand U5897 (N_5897,N_3309,N_2283);
nand U5898 (N_5898,N_2682,N_2304);
and U5899 (N_5899,N_2816,N_2444);
xor U5900 (N_5900,N_3832,N_2606);
nor U5901 (N_5901,N_2862,N_3318);
xor U5902 (N_5902,N_3015,N_3393);
nor U5903 (N_5903,N_2524,N_3920);
nor U5904 (N_5904,N_2250,N_2073);
and U5905 (N_5905,N_3783,N_3177);
nor U5906 (N_5906,N_2098,N_3030);
nor U5907 (N_5907,N_2573,N_3680);
nor U5908 (N_5908,N_2758,N_2077);
xnor U5909 (N_5909,N_2588,N_2215);
nor U5910 (N_5910,N_2304,N_2769);
and U5911 (N_5911,N_3667,N_2779);
and U5912 (N_5912,N_2390,N_2039);
nand U5913 (N_5913,N_3425,N_2221);
nand U5914 (N_5914,N_2587,N_2807);
or U5915 (N_5915,N_3031,N_3046);
xor U5916 (N_5916,N_2885,N_3659);
nor U5917 (N_5917,N_2815,N_3114);
xnor U5918 (N_5918,N_3586,N_2345);
and U5919 (N_5919,N_3901,N_3480);
xor U5920 (N_5920,N_2046,N_3574);
nand U5921 (N_5921,N_2549,N_2807);
nor U5922 (N_5922,N_3774,N_2438);
or U5923 (N_5923,N_3059,N_2957);
nor U5924 (N_5924,N_3072,N_2742);
or U5925 (N_5925,N_3441,N_3525);
nor U5926 (N_5926,N_3503,N_3771);
and U5927 (N_5927,N_2500,N_2540);
xor U5928 (N_5928,N_2117,N_2948);
and U5929 (N_5929,N_3324,N_3392);
nor U5930 (N_5930,N_2443,N_3319);
xor U5931 (N_5931,N_3834,N_2467);
xnor U5932 (N_5932,N_2772,N_3340);
nand U5933 (N_5933,N_2481,N_2629);
nand U5934 (N_5934,N_3430,N_2342);
and U5935 (N_5935,N_3047,N_3170);
xor U5936 (N_5936,N_2009,N_3473);
nor U5937 (N_5937,N_2779,N_2799);
and U5938 (N_5938,N_3342,N_3566);
or U5939 (N_5939,N_2313,N_3191);
nor U5940 (N_5940,N_3181,N_2776);
xor U5941 (N_5941,N_2048,N_2514);
and U5942 (N_5942,N_3201,N_3587);
xor U5943 (N_5943,N_2558,N_2830);
or U5944 (N_5944,N_2640,N_2484);
and U5945 (N_5945,N_3882,N_3455);
or U5946 (N_5946,N_2888,N_3022);
nand U5947 (N_5947,N_2984,N_3806);
xnor U5948 (N_5948,N_3643,N_2197);
xnor U5949 (N_5949,N_3077,N_3753);
xnor U5950 (N_5950,N_2722,N_2207);
xor U5951 (N_5951,N_2824,N_3616);
xnor U5952 (N_5952,N_3037,N_2283);
nand U5953 (N_5953,N_2388,N_2699);
and U5954 (N_5954,N_2151,N_2683);
and U5955 (N_5955,N_2556,N_2498);
or U5956 (N_5956,N_2746,N_3069);
xor U5957 (N_5957,N_3797,N_3067);
nor U5958 (N_5958,N_3022,N_3788);
and U5959 (N_5959,N_2269,N_3093);
or U5960 (N_5960,N_3617,N_3900);
nor U5961 (N_5961,N_2498,N_3108);
or U5962 (N_5962,N_2015,N_3247);
or U5963 (N_5963,N_2990,N_2511);
and U5964 (N_5964,N_2405,N_3541);
nor U5965 (N_5965,N_3393,N_2609);
or U5966 (N_5966,N_3414,N_2451);
nand U5967 (N_5967,N_3350,N_3460);
nor U5968 (N_5968,N_2025,N_3125);
and U5969 (N_5969,N_2783,N_2491);
xnor U5970 (N_5970,N_2357,N_3050);
and U5971 (N_5971,N_3192,N_2204);
nand U5972 (N_5972,N_2733,N_2194);
nor U5973 (N_5973,N_2533,N_3537);
or U5974 (N_5974,N_3125,N_2444);
and U5975 (N_5975,N_3370,N_2504);
or U5976 (N_5976,N_2690,N_3315);
nor U5977 (N_5977,N_2220,N_3400);
nor U5978 (N_5978,N_3398,N_3152);
xnor U5979 (N_5979,N_3048,N_2585);
xnor U5980 (N_5980,N_3955,N_3219);
and U5981 (N_5981,N_2606,N_2805);
and U5982 (N_5982,N_3569,N_3807);
xor U5983 (N_5983,N_3002,N_3877);
or U5984 (N_5984,N_3556,N_3520);
nor U5985 (N_5985,N_3239,N_2767);
xnor U5986 (N_5986,N_2608,N_3287);
nand U5987 (N_5987,N_2773,N_3088);
or U5988 (N_5988,N_2447,N_2444);
or U5989 (N_5989,N_2504,N_3569);
nand U5990 (N_5990,N_2998,N_3510);
xor U5991 (N_5991,N_2252,N_2130);
and U5992 (N_5992,N_3411,N_2000);
xnor U5993 (N_5993,N_3774,N_3150);
nand U5994 (N_5994,N_3698,N_3957);
nand U5995 (N_5995,N_2165,N_3519);
nand U5996 (N_5996,N_2638,N_3118);
nand U5997 (N_5997,N_2248,N_3432);
xnor U5998 (N_5998,N_2403,N_2327);
and U5999 (N_5999,N_3829,N_3229);
or U6000 (N_6000,N_5353,N_4990);
and U6001 (N_6001,N_4543,N_4946);
nor U6002 (N_6002,N_4933,N_4937);
or U6003 (N_6003,N_5699,N_5230);
nand U6004 (N_6004,N_4723,N_5479);
nand U6005 (N_6005,N_5847,N_4101);
nor U6006 (N_6006,N_4998,N_4696);
xor U6007 (N_6007,N_5131,N_4500);
xor U6008 (N_6008,N_5133,N_5826);
or U6009 (N_6009,N_5053,N_5561);
or U6010 (N_6010,N_4014,N_5812);
or U6011 (N_6011,N_5491,N_4005);
and U6012 (N_6012,N_4330,N_4428);
nor U6013 (N_6013,N_5168,N_4994);
or U6014 (N_6014,N_4917,N_4496);
and U6015 (N_6015,N_4032,N_4605);
nand U6016 (N_6016,N_4580,N_5486);
nand U6017 (N_6017,N_4073,N_5770);
and U6018 (N_6018,N_4858,N_4286);
and U6019 (N_6019,N_4690,N_4854);
nor U6020 (N_6020,N_5104,N_4702);
nor U6021 (N_6021,N_5748,N_5458);
nand U6022 (N_6022,N_5388,N_5063);
and U6023 (N_6023,N_4754,N_4042);
nand U6024 (N_6024,N_4852,N_4873);
xnor U6025 (N_6025,N_4640,N_5554);
and U6026 (N_6026,N_4148,N_4145);
nor U6027 (N_6027,N_4920,N_4447);
and U6028 (N_6028,N_4810,N_5771);
nor U6029 (N_6029,N_5326,N_4621);
or U6030 (N_6030,N_4597,N_4179);
or U6031 (N_6031,N_5312,N_5420);
nand U6032 (N_6032,N_4840,N_4289);
nand U6033 (N_6033,N_4913,N_4611);
nand U6034 (N_6034,N_5006,N_5531);
nor U6035 (N_6035,N_4384,N_5153);
nand U6036 (N_6036,N_4468,N_4086);
or U6037 (N_6037,N_5315,N_4189);
or U6038 (N_6038,N_5490,N_4398);
nand U6039 (N_6039,N_4035,N_5615);
or U6040 (N_6040,N_5555,N_5546);
and U6041 (N_6041,N_4066,N_5782);
or U6042 (N_6042,N_4886,N_5805);
xnor U6043 (N_6043,N_4107,N_4195);
nor U6044 (N_6044,N_4400,N_5648);
xnor U6045 (N_6045,N_5606,N_5525);
nor U6046 (N_6046,N_5849,N_5470);
xnor U6047 (N_6047,N_5138,N_4471);
xnor U6048 (N_6048,N_5210,N_5824);
and U6049 (N_6049,N_5270,N_4351);
nor U6050 (N_6050,N_4362,N_4747);
or U6051 (N_6051,N_4105,N_5079);
nand U6052 (N_6052,N_5054,N_5686);
xor U6053 (N_6053,N_4647,N_4223);
nor U6054 (N_6054,N_5533,N_5366);
and U6055 (N_6055,N_4487,N_5495);
xor U6056 (N_6056,N_5099,N_5905);
and U6057 (N_6057,N_5499,N_4415);
xnor U6058 (N_6058,N_5779,N_5067);
xnor U6059 (N_6059,N_4836,N_4764);
or U6060 (N_6060,N_5948,N_5136);
and U6061 (N_6061,N_4536,N_4555);
nor U6062 (N_6062,N_5220,N_4569);
or U6063 (N_6063,N_5384,N_4650);
or U6064 (N_6064,N_5897,N_4359);
or U6065 (N_6065,N_5840,N_5218);
or U6066 (N_6066,N_4341,N_4448);
or U6067 (N_6067,N_4720,N_5511);
nand U6068 (N_6068,N_4094,N_4576);
and U6069 (N_6069,N_4401,N_4615);
and U6070 (N_6070,N_4164,N_5758);
and U6071 (N_6071,N_5471,N_5888);
or U6072 (N_6072,N_5266,N_5576);
nor U6073 (N_6073,N_5708,N_4649);
nor U6074 (N_6074,N_4343,N_4509);
xnor U6075 (N_6075,N_4224,N_4114);
or U6076 (N_6076,N_4349,N_4001);
xnor U6077 (N_6077,N_5057,N_4502);
and U6078 (N_6078,N_4860,N_5354);
nor U6079 (N_6079,N_4353,N_4914);
and U6080 (N_6080,N_5636,N_5478);
and U6081 (N_6081,N_5919,N_4390);
xor U6082 (N_6082,N_5653,N_5788);
xnor U6083 (N_6083,N_4602,N_5151);
nand U6084 (N_6084,N_5375,N_5473);
and U6085 (N_6085,N_4078,N_5338);
nand U6086 (N_6086,N_5268,N_4648);
and U6087 (N_6087,N_5090,N_4182);
nor U6088 (N_6088,N_5144,N_4120);
and U6089 (N_6089,N_5907,N_4756);
nor U6090 (N_6090,N_5065,N_5221);
or U6091 (N_6091,N_4187,N_5896);
or U6092 (N_6092,N_5706,N_5660);
nand U6093 (N_6093,N_4516,N_4089);
xor U6094 (N_6094,N_5007,N_5272);
nand U6095 (N_6095,N_5629,N_5405);
and U6096 (N_6096,N_4628,N_4241);
nor U6097 (N_6097,N_5581,N_4667);
nand U6098 (N_6098,N_5768,N_4897);
or U6099 (N_6099,N_4916,N_5833);
nand U6100 (N_6100,N_5031,N_5619);
nand U6101 (N_6101,N_4176,N_4675);
and U6102 (N_6102,N_4177,N_5997);
xnor U6103 (N_6103,N_5317,N_4772);
and U6104 (N_6104,N_5194,N_5383);
and U6105 (N_6105,N_5801,N_4358);
or U6106 (N_6106,N_4503,N_4497);
nand U6107 (N_6107,N_4910,N_5687);
nor U6108 (N_6108,N_5627,N_4950);
xnor U6109 (N_6109,N_5593,N_5475);
xnor U6110 (N_6110,N_4738,N_4634);
nand U6111 (N_6111,N_5208,N_4807);
xnor U6112 (N_6112,N_4581,N_5774);
or U6113 (N_6113,N_4967,N_4713);
or U6114 (N_6114,N_4318,N_5372);
nand U6115 (N_6115,N_5158,N_4760);
nor U6116 (N_6116,N_4368,N_4593);
nor U6117 (N_6117,N_5407,N_4282);
nand U6118 (N_6118,N_4725,N_5392);
xnor U6119 (N_6119,N_5460,N_4135);
and U6120 (N_6120,N_5953,N_4494);
or U6121 (N_6121,N_5841,N_4534);
xnor U6122 (N_6122,N_5042,N_4595);
and U6123 (N_6123,N_5258,N_5890);
xnor U6124 (N_6124,N_5584,N_4076);
or U6125 (N_6125,N_5331,N_4273);
xor U6126 (N_6126,N_5111,N_4780);
xnor U6127 (N_6127,N_4201,N_5431);
nand U6128 (N_6128,N_4952,N_4252);
and U6129 (N_6129,N_4827,N_5966);
nor U6130 (N_6130,N_4969,N_5021);
nand U6131 (N_6131,N_4226,N_4488);
nand U6132 (N_6132,N_5514,N_4731);
xor U6133 (N_6133,N_5709,N_5704);
and U6134 (N_6134,N_5624,N_5886);
or U6135 (N_6135,N_5573,N_5229);
or U6136 (N_6136,N_4656,N_5149);
xnor U6137 (N_6137,N_5910,N_4557);
nor U6138 (N_6138,N_4792,N_4459);
or U6139 (N_6139,N_4927,N_4470);
and U6140 (N_6140,N_4165,N_4207);
xnor U6141 (N_6141,N_5736,N_5175);
nor U6142 (N_6142,N_4213,N_5303);
xor U6143 (N_6143,N_4857,N_5887);
or U6144 (N_6144,N_4370,N_4681);
or U6145 (N_6145,N_4413,N_5726);
nor U6146 (N_6146,N_5677,N_4638);
nor U6147 (N_6147,N_5797,N_5493);
nor U6148 (N_6148,N_5050,N_4833);
xor U6149 (N_6149,N_5510,N_4092);
nand U6150 (N_6150,N_4402,N_5901);
xnor U6151 (N_6151,N_4717,N_5800);
and U6152 (N_6152,N_5459,N_5682);
nand U6153 (N_6153,N_5981,N_5189);
or U6154 (N_6154,N_5792,N_4715);
and U6155 (N_6155,N_5160,N_5364);
and U6156 (N_6156,N_4976,N_4924);
xor U6157 (N_6157,N_4708,N_5608);
nor U6158 (N_6158,N_5535,N_5938);
or U6159 (N_6159,N_4169,N_4229);
or U6160 (N_6160,N_4452,N_5185);
and U6161 (N_6161,N_5643,N_4083);
nand U6162 (N_6162,N_5976,N_5003);
nand U6163 (N_6163,N_4185,N_4275);
and U6164 (N_6164,N_4124,N_4054);
nor U6165 (N_6165,N_4624,N_4737);
nand U6166 (N_6166,N_4668,N_4683);
xor U6167 (N_6167,N_4588,N_4830);
or U6168 (N_6168,N_5062,N_5080);
nand U6169 (N_6169,N_5305,N_5601);
xor U6170 (N_6170,N_4344,N_5162);
or U6171 (N_6171,N_5716,N_5568);
and U6172 (N_6172,N_5813,N_5061);
xnor U6173 (N_6173,N_4440,N_4791);
and U6174 (N_6174,N_4865,N_5698);
xnor U6175 (N_6175,N_5645,N_4257);
and U6176 (N_6176,N_5191,N_4877);
nor U6177 (N_6177,N_4811,N_5735);
nand U6178 (N_6178,N_5879,N_4979);
xor U6179 (N_6179,N_5323,N_4197);
and U6180 (N_6180,N_5836,N_4255);
nor U6181 (N_6181,N_4556,N_4531);
or U6182 (N_6182,N_5279,N_5937);
or U6183 (N_6183,N_5052,N_4396);
nor U6184 (N_6184,N_5588,N_5763);
or U6185 (N_6185,N_5492,N_5900);
xnor U6186 (N_6186,N_4377,N_5227);
or U6187 (N_6187,N_4117,N_4333);
xnor U6188 (N_6188,N_4878,N_5424);
nor U6189 (N_6189,N_4080,N_5505);
nor U6190 (N_6190,N_4485,N_5127);
nand U6191 (N_6191,N_5330,N_4016);
nor U6192 (N_6192,N_4512,N_5286);
or U6193 (N_6193,N_5283,N_5846);
nor U6194 (N_6194,N_5806,N_4298);
or U6195 (N_6195,N_5607,N_5569);
nor U6196 (N_6196,N_4206,N_5742);
or U6197 (N_6197,N_4566,N_4309);
and U6198 (N_6198,N_5030,N_4064);
nor U6199 (N_6199,N_5026,N_4112);
nor U6200 (N_6200,N_4160,N_4748);
and U6201 (N_6201,N_4700,N_4726);
or U6202 (N_6202,N_5260,N_4855);
nand U6203 (N_6203,N_5710,N_5853);
and U6204 (N_6204,N_4276,N_4711);
and U6205 (N_6205,N_4590,N_5579);
nor U6206 (N_6206,N_5999,N_4002);
nor U6207 (N_6207,N_4239,N_5074);
and U6208 (N_6208,N_5044,N_4366);
nand U6209 (N_6209,N_5835,N_4443);
and U6210 (N_6210,N_5603,N_4859);
nand U6211 (N_6211,N_5688,N_5228);
or U6212 (N_6212,N_5411,N_4460);
nor U6213 (N_6213,N_5254,N_4520);
and U6214 (N_6214,N_4710,N_5327);
and U6215 (N_6215,N_4012,N_4321);
nor U6216 (N_6216,N_5832,N_5845);
and U6217 (N_6217,N_5920,N_5998);
nand U6218 (N_6218,N_5134,N_4481);
nor U6219 (N_6219,N_4641,N_5250);
nand U6220 (N_6220,N_4272,N_5440);
or U6221 (N_6221,N_4437,N_5929);
xor U6222 (N_6222,N_5963,N_5059);
or U6223 (N_6223,N_5817,N_4332);
nor U6224 (N_6224,N_4584,N_5213);
xnor U6225 (N_6225,N_4819,N_5591);
xor U6226 (N_6226,N_4184,N_5772);
or U6227 (N_6227,N_4123,N_5516);
and U6228 (N_6228,N_4564,N_4911);
nor U6229 (N_6229,N_4354,N_5413);
nand U6230 (N_6230,N_4074,N_5098);
xor U6231 (N_6231,N_4313,N_5039);
nand U6232 (N_6232,N_5542,N_4813);
or U6233 (N_6233,N_5173,N_4941);
and U6234 (N_6234,N_5683,N_4698);
nor U6235 (N_6235,N_4997,N_5638);
nor U6236 (N_6236,N_4155,N_5680);
and U6237 (N_6237,N_4655,N_5344);
or U6238 (N_6238,N_4242,N_5773);
nand U6239 (N_6239,N_4186,N_4826);
or U6240 (N_6240,N_4922,N_4104);
xor U6241 (N_6241,N_5930,N_4323);
nand U6242 (N_6242,N_4316,N_5496);
xnor U6243 (N_6243,N_4974,N_4767);
and U6244 (N_6244,N_4191,N_5081);
nor U6245 (N_6245,N_5744,N_4430);
or U6246 (N_6246,N_5859,N_5156);
xor U6247 (N_6247,N_5519,N_4525);
and U6248 (N_6248,N_5426,N_4750);
or U6249 (N_6249,N_4706,N_5861);
nor U6250 (N_6250,N_4909,N_5345);
xor U6251 (N_6251,N_4434,N_4126);
xnor U6252 (N_6252,N_4142,N_5640);
xnor U6253 (N_6253,N_4539,N_4306);
and U6254 (N_6254,N_5357,N_4567);
and U6255 (N_6255,N_4181,N_5750);
nor U6256 (N_6256,N_4968,N_4227);
nand U6257 (N_6257,N_5321,N_5784);
xor U6258 (N_6258,N_5666,N_5425);
xnor U6259 (N_6259,N_4834,N_5702);
nor U6260 (N_6260,N_4339,N_5301);
nand U6261 (N_6261,N_4194,N_5298);
or U6262 (N_6262,N_5862,N_5926);
nand U6263 (N_6263,N_4336,N_4793);
and U6264 (N_6264,N_4815,N_5646);
or U6265 (N_6265,N_4847,N_4929);
and U6266 (N_6266,N_5015,N_5122);
nor U6267 (N_6267,N_4371,N_5055);
nor U6268 (N_6268,N_5786,N_4270);
xnor U6269 (N_6269,N_5180,N_4600);
or U6270 (N_6270,N_4015,N_4719);
nand U6271 (N_6271,N_5667,N_4975);
nor U6272 (N_6272,N_4109,N_4778);
xor U6273 (N_6273,N_5237,N_4940);
xor U6274 (N_6274,N_5913,N_5439);
nand U6275 (N_6275,N_4279,N_4458);
nand U6276 (N_6276,N_5393,N_4730);
nor U6277 (N_6277,N_4131,N_4904);
nand U6278 (N_6278,N_5723,N_5794);
nor U6279 (N_6279,N_4510,N_5793);
nand U6280 (N_6280,N_5572,N_5285);
nor U6281 (N_6281,N_5759,N_5373);
or U6282 (N_6282,N_5060,N_5116);
and U6283 (N_6283,N_5123,N_5087);
xor U6284 (N_6284,N_5170,N_5165);
and U6285 (N_6285,N_4800,N_5662);
or U6286 (N_6286,N_5022,N_4570);
nand U6287 (N_6287,N_4938,N_5565);
xor U6288 (N_6288,N_4444,N_5322);
nor U6289 (N_6289,N_4880,N_5537);
nor U6290 (N_6290,N_5802,N_5939);
and U6291 (N_6291,N_4085,N_5091);
xnor U6292 (N_6292,N_4703,N_4561);
nor U6293 (N_6293,N_5147,N_5583);
or U6294 (N_6294,N_5747,N_4954);
nand U6295 (N_6295,N_4571,N_5520);
or U6296 (N_6296,N_4307,N_4820);
nor U6297 (N_6297,N_5314,N_5140);
and U6298 (N_6298,N_5261,N_5540);
xnor U6299 (N_6299,N_4315,N_4274);
nor U6300 (N_6300,N_4449,N_5130);
and U6301 (N_6301,N_4939,N_5614);
and U6302 (N_6302,N_4423,N_4193);
or U6303 (N_6303,N_5652,N_4716);
nand U6304 (N_6304,N_4971,N_4832);
and U6305 (N_6305,N_4118,N_5013);
or U6306 (N_6306,N_5946,N_4781);
xor U6307 (N_6307,N_4410,N_4809);
and U6308 (N_6308,N_5329,N_4232);
or U6309 (N_6309,N_5755,N_4484);
or U6310 (N_6310,N_4517,N_4742);
and U6311 (N_6311,N_4258,N_4028);
nor U6312 (N_6312,N_4798,N_4823);
xor U6313 (N_6313,N_4388,N_4299);
or U6314 (N_6314,N_5951,N_4003);
nand U6315 (N_6315,N_4486,N_5417);
and U6316 (N_6316,N_4314,N_4235);
nand U6317 (N_6317,N_5611,N_4613);
nand U6318 (N_6318,N_4023,N_4524);
xor U6319 (N_6319,N_4345,N_5635);
or U6320 (N_6320,N_5334,N_5455);
xor U6321 (N_6321,N_4373,N_4743);
nor U6322 (N_6322,N_5668,N_5198);
nor U6323 (N_6323,N_5066,N_5560);
nor U6324 (N_6324,N_5828,N_4856);
and U6325 (N_6325,N_4757,N_5255);
or U6326 (N_6326,N_4870,N_4669);
nor U6327 (N_6327,N_5665,N_5796);
nor U6328 (N_6328,N_4499,N_5441);
xnor U6329 (N_6329,N_4987,N_4728);
and U6330 (N_6330,N_5863,N_4558);
nand U6331 (N_6331,N_4672,N_5501);
and U6332 (N_6332,N_4381,N_5857);
xnor U6333 (N_6333,N_5368,N_5647);
xor U6334 (N_6334,N_5864,N_4753);
nand U6335 (N_6335,N_5429,N_5017);
and U6336 (N_6336,N_5957,N_5422);
nand U6337 (N_6337,N_4596,N_5713);
nor U6338 (N_6338,N_4659,N_5450);
nor U6339 (N_6339,N_5819,N_5192);
nor U6340 (N_6340,N_4661,N_4419);
nand U6341 (N_6341,N_4689,N_4046);
or U6342 (N_6342,N_5989,N_4462);
xor U6343 (N_6343,N_4346,N_5274);
xnor U6344 (N_6344,N_5076,N_5644);
nand U6345 (N_6345,N_4053,N_5086);
nor U6346 (N_6346,N_5454,N_4755);
xor U6347 (N_6347,N_5848,N_5075);
nor U6348 (N_6348,N_5179,N_5115);
xnor U6349 (N_6349,N_4612,N_5503);
or U6350 (N_6350,N_4495,N_4418);
nand U6351 (N_6351,N_4765,N_4412);
nand U6352 (N_6352,N_5476,N_4945);
nor U6353 (N_6353,N_5316,N_5226);
and U6354 (N_6354,N_4347,N_5558);
nand U6355 (N_6355,N_4477,N_4125);
nand U6356 (N_6356,N_4718,N_5690);
and U6357 (N_6357,N_5442,N_5547);
nand U6358 (N_6358,N_5852,N_4296);
nor U6359 (N_6359,N_4523,N_5186);
nor U6360 (N_6360,N_4773,N_4542);
nand U6361 (N_6361,N_5814,N_5933);
or U6362 (N_6362,N_4721,N_5958);
nor U6363 (N_6363,N_4797,N_4029);
nand U6364 (N_6364,N_4565,N_4949);
nand U6365 (N_6365,N_4901,N_4008);
xor U6366 (N_6366,N_4483,N_5893);
or U6367 (N_6367,N_5245,N_4021);
nand U6368 (N_6368,N_5599,N_4635);
xor U6369 (N_6369,N_5892,N_5273);
nor U6370 (N_6370,N_5409,N_4249);
nor U6371 (N_6371,N_5906,N_5700);
and U6372 (N_6372,N_5985,N_4744);
nor U6373 (N_6373,N_4674,N_4845);
and U6374 (N_6374,N_5685,N_4006);
nand U6375 (N_6375,N_5679,N_4694);
nor U6376 (N_6376,N_4930,N_5674);
nand U6377 (N_6377,N_4287,N_5775);
nor U6378 (N_6378,N_4283,N_4657);
and U6379 (N_6379,N_4127,N_5359);
xnor U6380 (N_6380,N_5453,N_4426);
nor U6381 (N_6381,N_4662,N_5928);
and U6382 (N_6382,N_5243,N_5717);
or U6383 (N_6383,N_4592,N_5877);
nand U6384 (N_6384,N_5033,N_5159);
or U6385 (N_6385,N_4876,N_5046);
nand U6386 (N_6386,N_4693,N_5415);
nand U6387 (N_6387,N_5880,N_5382);
nor U6388 (N_6388,N_4060,N_4093);
nor U6389 (N_6389,N_4899,N_4095);
nand U6390 (N_6390,N_4508,N_5304);
and U6391 (N_6391,N_4055,N_5798);
nand U6392 (N_6392,N_4884,N_4424);
or U6393 (N_6393,N_4892,N_5038);
nor U6394 (N_6394,N_4266,N_4931);
or U6395 (N_6395,N_5288,N_4106);
nor U6396 (N_6396,N_5068,N_5350);
and U6397 (N_6397,N_5870,N_5727);
nand U6398 (N_6398,N_5625,N_5232);
and U6399 (N_6399,N_5843,N_4958);
xnor U6400 (N_6400,N_4658,N_5231);
nand U6401 (N_6401,N_5000,N_4153);
and U6402 (N_6402,N_5975,N_4944);
or U6403 (N_6403,N_4137,N_4705);
xor U6404 (N_6404,N_4671,N_4311);
or U6405 (N_6405,N_4453,N_4769);
and U6406 (N_6406,N_5952,N_5306);
nand U6407 (N_6407,N_5672,N_5477);
nand U6408 (N_6408,N_5355,N_5837);
or U6409 (N_6409,N_4156,N_4775);
nand U6410 (N_6410,N_4614,N_4507);
or U6411 (N_6411,N_5823,N_4215);
and U6412 (N_6412,N_5696,N_5869);
nand U6413 (N_6413,N_5497,N_4217);
and U6414 (N_6414,N_4328,N_4943);
or U6415 (N_6415,N_4240,N_5737);
or U6416 (N_6416,N_5214,N_5597);
and U6417 (N_6417,N_4983,N_5570);
nor U6418 (N_6418,N_5803,N_4806);
nor U6419 (N_6419,N_4573,N_4000);
xnor U6420 (N_6420,N_5012,N_5464);
and U6421 (N_6421,N_4464,N_5148);
and U6422 (N_6422,N_4547,N_5113);
nor U6423 (N_6423,N_5663,N_4977);
nand U6424 (N_6424,N_4271,N_5223);
nand U6425 (N_6425,N_4896,N_5918);
nor U6426 (N_6426,N_4526,N_4455);
or U6427 (N_6427,N_4161,N_4546);
nor U6428 (N_6428,N_5348,N_4680);
xnor U6429 (N_6429,N_5203,N_4335);
or U6430 (N_6430,N_4660,N_5567);
nor U6431 (N_6431,N_5522,N_4166);
nand U6432 (N_6432,N_4626,N_5083);
xnor U6433 (N_6433,N_5965,N_4350);
or U6434 (N_6434,N_5810,N_4212);
and U6435 (N_6435,N_5362,N_5871);
or U6436 (N_6436,N_5856,N_5552);
nand U6437 (N_6437,N_5942,N_4849);
and U6438 (N_6438,N_4456,N_5152);
xor U6439 (N_6439,N_4491,N_5831);
or U6440 (N_6440,N_5884,N_4972);
nor U6441 (N_6441,N_5557,N_4218);
and U6442 (N_6442,N_5071,N_4637);
nor U6443 (N_6443,N_5340,N_4727);
or U6444 (N_6444,N_5724,N_5387);
xnor U6445 (N_6445,N_4399,N_5137);
nor U6446 (N_6446,N_4466,N_5633);
nand U6447 (N_6447,N_4956,N_5002);
or U6448 (N_6448,N_5527,N_4794);
nor U6449 (N_6449,N_5275,N_5177);
nor U6450 (N_6450,N_4248,N_4281);
xnor U6451 (N_6451,N_5851,N_5436);
xnor U6452 (N_6452,N_4905,N_4018);
xor U6453 (N_6453,N_4643,N_5551);
nor U6454 (N_6454,N_4790,N_5927);
xnor U6455 (N_6455,N_4139,N_5754);
and U6456 (N_6456,N_5947,N_5371);
or U6457 (N_6457,N_4267,N_4084);
nor U6458 (N_6458,N_4246,N_4233);
or U6459 (N_6459,N_5733,N_5419);
xnor U6460 (N_6460,N_5449,N_5743);
or U6461 (N_6461,N_4277,N_5019);
xnor U6462 (N_6462,N_5932,N_4540);
and U6463 (N_6463,N_4397,N_5783);
or U6464 (N_6464,N_5307,N_4872);
xor U6465 (N_6465,N_5563,N_4686);
nor U6466 (N_6466,N_5815,N_5728);
nor U6467 (N_6467,N_4045,N_4438);
or U6468 (N_6468,N_4928,N_4688);
or U6469 (N_6469,N_5457,N_4642);
xnor U6470 (N_6470,N_5539,N_4416);
xnor U6471 (N_6471,N_4868,N_4532);
nand U6472 (N_6472,N_4871,N_4818);
nand U6473 (N_6473,N_4995,N_4630);
nand U6474 (N_6474,N_4219,N_5903);
xnor U6475 (N_6475,N_5167,N_4947);
xor U6476 (N_6476,N_5882,N_5534);
nor U6477 (N_6477,N_5181,N_4162);
xor U6478 (N_6478,N_4036,N_5135);
nor U6479 (N_6479,N_5923,N_4704);
or U6480 (N_6480,N_4964,N_4966);
or U6481 (N_6481,N_4620,N_5294);
nor U6482 (N_6482,N_4091,N_5705);
nor U6483 (N_6483,N_5760,N_4250);
nor U6484 (N_6484,N_4766,N_5617);
or U6485 (N_6485,N_5990,N_5820);
and U6486 (N_6486,N_4712,N_5487);
xnor U6487 (N_6487,N_4861,N_4665);
nor U6488 (N_6488,N_4202,N_4171);
xnor U6489 (N_6489,N_4692,N_4454);
and U6490 (N_6490,N_5598,N_5515);
and U6491 (N_6491,N_5657,N_4041);
xor U6492 (N_6492,N_4549,N_5049);
or U6493 (N_6493,N_4110,N_4088);
or U6494 (N_6494,N_4034,N_5566);
nand U6495 (N_6495,N_4514,N_4408);
xnor U6496 (N_6496,N_5023,N_5944);
nand U6497 (N_6497,N_4312,N_5146);
nor U6498 (N_6498,N_4993,N_5289);
xor U6499 (N_6499,N_4821,N_4493);
and U6500 (N_6500,N_4887,N_4926);
nand U6501 (N_6501,N_4942,N_5623);
and U6502 (N_6502,N_5973,N_4450);
nor U6503 (N_6503,N_5577,N_5311);
xor U6504 (N_6504,N_5675,N_5452);
nor U6505 (N_6505,N_4157,N_4480);
nor U6506 (N_6506,N_5504,N_4379);
or U6507 (N_6507,N_5589,N_5414);
and U6508 (N_6508,N_5585,N_5078);
nor U6509 (N_6509,N_5196,N_5960);
and U6510 (N_6510,N_4141,N_4603);
nor U6511 (N_6511,N_4752,N_5512);
xor U6512 (N_6512,N_5445,N_5889);
nand U6513 (N_6513,N_5058,N_4801);
nand U6514 (N_6514,N_5269,N_4303);
nand U6515 (N_6515,N_4869,N_5749);
xor U6516 (N_6516,N_4327,N_5883);
xor U6517 (N_6517,N_5300,N_4251);
xor U6518 (N_6518,N_5549,N_5402);
or U6519 (N_6519,N_4779,N_4687);
or U6520 (N_6520,N_4382,N_5873);
xnor U6521 (N_6521,N_5866,N_4147);
xor U6522 (N_6522,N_4724,N_5632);
xnor U6523 (N_6523,N_5481,N_4051);
nor U6524 (N_6524,N_4133,N_5163);
nand U6525 (N_6525,N_4898,N_5885);
xnor U6526 (N_6526,N_5894,N_5001);
and U6527 (N_6527,N_4208,N_5313);
nand U6528 (N_6528,N_5084,N_5988);
and U6529 (N_6529,N_5474,N_5265);
nor U6530 (N_6530,N_5154,N_5949);
or U6531 (N_6531,N_5290,N_4190);
nor U6532 (N_6532,N_4039,N_4519);
nand U6533 (N_6533,N_4069,N_4770);
nor U6534 (N_6534,N_4915,N_5169);
nand U6535 (N_6535,N_5924,N_4150);
and U6536 (N_6536,N_5207,N_5374);
nand U6537 (N_6537,N_5982,N_5281);
and U6538 (N_6538,N_4632,N_4268);
xnor U6539 (N_6539,N_4985,N_5484);
or U6540 (N_6540,N_4623,N_4888);
nand U6541 (N_6541,N_5746,N_4163);
nor U6542 (N_6542,N_5738,N_5132);
and U6543 (N_6543,N_4010,N_5241);
and U6544 (N_6544,N_5526,N_5112);
or U6545 (N_6545,N_5881,N_5047);
and U6546 (N_6546,N_4269,N_4572);
nor U6547 (N_6547,N_5139,N_4594);
or U6548 (N_6548,N_5124,N_5661);
xnor U6549 (N_6549,N_5034,N_5968);
xor U6550 (N_6550,N_5757,N_5073);
xnor U6551 (N_6551,N_4619,N_5020);
or U6552 (N_6552,N_5187,N_5876);
nand U6553 (N_6553,N_5277,N_4553);
or U6554 (N_6554,N_4639,N_4260);
nand U6555 (N_6555,N_5339,N_4552);
and U6556 (N_6556,N_4759,N_4537);
or U6557 (N_6557,N_5120,N_5586);
nor U6558 (N_6558,N_5955,N_5463);
nor U6559 (N_6559,N_4828,N_4262);
nand U6560 (N_6560,N_5945,N_5764);
xor U6561 (N_6561,N_4749,N_4951);
xnor U6562 (N_6562,N_4607,N_4294);
xor U6563 (N_6563,N_5018,N_4441);
or U6564 (N_6564,N_5753,N_5631);
xor U6565 (N_6565,N_4253,N_5070);
and U6566 (N_6566,N_5821,N_5390);
nand U6567 (N_6567,N_5681,N_5358);
nor U6568 (N_6568,N_4038,N_5695);
nor U6569 (N_6569,N_5781,N_4103);
nor U6570 (N_6570,N_4900,N_5891);
or U6571 (N_6571,N_4387,N_5751);
nor U6572 (N_6572,N_5200,N_4875);
and U6573 (N_6573,N_4234,N_4442);
xor U6574 (N_6574,N_5541,N_4636);
nand U6575 (N_6575,N_4825,N_5010);
nand U6576 (N_6576,N_4254,N_5011);
nand U6577 (N_6577,N_4682,N_4203);
and U6578 (N_6578,N_4152,N_4411);
and U6579 (N_6579,N_4850,N_4374);
nand U6580 (N_6580,N_4172,N_4098);
nor U6581 (N_6581,N_4265,N_4782);
or U6582 (N_6582,N_5992,N_5712);
or U6583 (N_6583,N_4340,N_4919);
nor U6584 (N_6584,N_5253,N_5027);
xnor U6585 (N_6585,N_4629,N_5105);
and U6586 (N_6586,N_5095,N_5795);
xor U6587 (N_6587,N_5618,N_4992);
nor U6588 (N_6588,N_4545,N_5502);
nand U6589 (N_6589,N_5430,N_4158);
nand U6590 (N_6590,N_4071,N_4563);
and U6591 (N_6591,N_5829,N_5335);
xor U6592 (N_6592,N_5145,N_5293);
nor U6593 (N_6593,N_5498,N_4541);
nor U6594 (N_6594,N_5333,N_5908);
and U6595 (N_6595,N_5834,N_4652);
and U6596 (N_6596,N_5962,N_5217);
and U6597 (N_6597,N_5969,N_5816);
nor U6598 (N_6598,N_5718,N_5064);
xnor U6599 (N_6599,N_5400,N_4367);
or U6600 (N_6600,N_4885,N_5443);
xor U6601 (N_6601,N_5142,N_5921);
or U6602 (N_6602,N_4902,N_4864);
nand U6603 (N_6603,N_5418,N_4835);
xnor U6604 (N_6604,N_4457,N_5378);
nand U6605 (N_6605,N_4027,N_4799);
nor U6606 (N_6606,N_5909,N_5488);
or U6607 (N_6607,N_4013,N_5671);
nand U6608 (N_6608,N_5872,N_5435);
or U6609 (N_6609,N_5637,N_4548);
and U6610 (N_6610,N_4599,N_4331);
xnor U6611 (N_6611,N_4099,N_5045);
and U6612 (N_6612,N_4288,N_5818);
or U6613 (N_6613,N_5532,N_5320);
and U6614 (N_6614,N_4739,N_4445);
and U6615 (N_6615,N_4421,N_5655);
or U6616 (N_6616,N_5240,N_5518);
or U6617 (N_6617,N_4862,N_4129);
or U6618 (N_6618,N_5991,N_4204);
nor U6619 (N_6619,N_4986,N_4957);
and U6620 (N_6620,N_5467,N_5182);
nor U6621 (N_6621,N_4653,N_5844);
nor U6622 (N_6622,N_5363,N_4210);
and U6623 (N_6623,N_5117,N_5398);
or U6624 (N_6624,N_5389,N_5209);
and U6625 (N_6625,N_4867,N_5711);
nand U6626 (N_6626,N_4812,N_5267);
nor U6627 (N_6627,N_4802,N_4465);
xor U6628 (N_6628,N_4116,N_4079);
nand U6629 (N_6629,N_4735,N_4435);
nand U6630 (N_6630,N_4132,N_4645);
or U6631 (N_6631,N_5256,N_4263);
nand U6632 (N_6632,N_5244,N_5257);
or U6633 (N_6633,N_5296,N_5291);
nand U6634 (N_6634,N_4965,N_4225);
and U6635 (N_6635,N_5689,N_4808);
and U6636 (N_6636,N_4057,N_5590);
or U6637 (N_6637,N_4280,N_4691);
and U6638 (N_6638,N_4577,N_4087);
nor U6639 (N_6639,N_4676,N_5219);
and U6640 (N_6640,N_4231,N_4722);
nor U6641 (N_6641,N_5238,N_5205);
nand U6642 (N_6642,N_4200,N_5352);
or U6643 (N_6643,N_5143,N_4505);
or U6644 (N_6644,N_4030,N_4290);
and U6645 (N_6645,N_5360,N_5069);
nand U6646 (N_6646,N_4617,N_5215);
nand U6647 (N_6647,N_5456,N_4259);
and U6648 (N_6648,N_5808,N_5654);
or U6649 (N_6649,N_5048,N_5935);
and U6650 (N_6650,N_5094,N_4199);
nor U6651 (N_6651,N_4360,N_4734);
xnor U6652 (N_6652,N_5336,N_5934);
and U6653 (N_6653,N_5842,N_4325);
and U6654 (N_6654,N_4244,N_5157);
and U6655 (N_6655,N_5550,N_4461);
nor U6656 (N_6656,N_5649,N_5089);
and U6657 (N_6657,N_5204,N_4222);
xnor U6658 (N_6658,N_4154,N_4999);
nand U6659 (N_6659,N_4559,N_5610);
xnor U6660 (N_6660,N_4839,N_4238);
nand U6661 (N_6661,N_4511,N_5943);
nand U6662 (N_6662,N_4173,N_4026);
or U6663 (N_6663,N_5658,N_4096);
nor U6664 (N_6664,N_5234,N_5613);
xnor U6665 (N_6665,N_4891,N_5964);
and U6666 (N_6666,N_4774,N_4304);
and U6667 (N_6667,N_4198,N_4378);
and U6668 (N_6668,N_4319,N_4420);
or U6669 (N_6669,N_4236,N_5102);
and U6670 (N_6670,N_5308,N_4970);
nor U6671 (N_6671,N_4352,N_5485);
and U6672 (N_6672,N_5656,N_4052);
and U6673 (N_6673,N_5101,N_4518);
or U6674 (N_6674,N_4044,N_5318);
nor U6675 (N_6675,N_5741,N_5121);
and U6676 (N_6676,N_5437,N_4535);
nor U6677 (N_6677,N_5150,N_5029);
or U6678 (N_6678,N_5468,N_5097);
xor U6679 (N_6679,N_5839,N_4009);
xor U6680 (N_6680,N_4527,N_5941);
nor U6681 (N_6681,N_5508,N_5199);
xnor U6682 (N_6682,N_4521,N_5571);
and U6683 (N_6683,N_4824,N_5129);
nor U6684 (N_6684,N_4663,N_4934);
nand U6685 (N_6685,N_4533,N_5292);
xnor U6686 (N_6686,N_5521,N_4697);
nand U6687 (N_6687,N_5595,N_4538);
nand U6688 (N_6688,N_4081,N_5838);
nand U6689 (N_6689,N_4804,N_5448);
nand U6690 (N_6690,N_5472,N_4771);
nor U6691 (N_6691,N_5280,N_5513);
nand U6692 (N_6692,N_4334,N_5251);
or U6693 (N_6693,N_4608,N_4019);
and U6694 (N_6694,N_5931,N_4805);
nand U6695 (N_6695,N_5423,N_5216);
nand U6696 (N_6696,N_4385,N_4490);
xnor U6697 (N_6697,N_5427,N_4589);
and U6698 (N_6698,N_4243,N_5404);
nand U6699 (N_6699,N_4167,N_4988);
xor U6700 (N_6700,N_5902,N_5107);
xor U6701 (N_6701,N_5103,N_4404);
xor U6702 (N_6702,N_4893,N_5341);
nor U6703 (N_6703,N_4431,N_5830);
nand U6704 (N_6704,N_4784,N_5582);
xor U6705 (N_6705,N_5166,N_5536);
nand U6706 (N_6706,N_5155,N_4844);
nand U6707 (N_6707,N_5622,N_5451);
nor U6708 (N_6708,N_5401,N_4136);
nand U6709 (N_6709,N_5394,N_4554);
or U6710 (N_6710,N_4326,N_4077);
nor U6711 (N_6711,N_4146,N_5004);
xor U6712 (N_6712,N_5016,N_4439);
xnor U6713 (N_6713,N_5119,N_4245);
nand U6714 (N_6714,N_4618,N_5282);
or U6715 (N_6715,N_5925,N_5174);
xor U6716 (N_6716,N_4033,N_4405);
and U6717 (N_6717,N_4796,N_4031);
and U6718 (N_6718,N_5391,N_5295);
or U6719 (N_6719,N_4587,N_4407);
nor U6720 (N_6720,N_5195,N_5956);
nand U6721 (N_6721,N_5789,N_4881);
nand U6722 (N_6722,N_4814,N_4786);
and U6723 (N_6723,N_4903,N_5114);
xor U6724 (N_6724,N_5904,N_4740);
or U6725 (N_6725,N_5641,N_4478);
or U6726 (N_6726,N_5403,N_5264);
or U6727 (N_6727,N_4787,N_4357);
xor U6728 (N_6728,N_5630,N_5574);
or U6729 (N_6729,N_4961,N_5164);
xnor U6730 (N_6730,N_4575,N_4059);
xnor U6731 (N_6731,N_5692,N_4701);
nor U6732 (N_6732,N_4768,N_4004);
nand U6733 (N_6733,N_5684,N_5993);
nand U6734 (N_6734,N_4022,N_5523);
and U6735 (N_6735,N_5776,N_5118);
nor U6736 (N_6736,N_5005,N_5088);
nor U6737 (N_6737,N_5299,N_5380);
or U6738 (N_6738,N_4989,N_4376);
and U6739 (N_6739,N_4302,N_5730);
and U6740 (N_6740,N_5025,N_4380);
nand U6741 (N_6741,N_4838,N_5791);
xor U6742 (N_6742,N_4732,N_4846);
or U6743 (N_6743,N_5056,N_4670);
xor U6744 (N_6744,N_4578,N_5379);
xor U6745 (N_6745,N_4677,N_4606);
and U6746 (N_6746,N_4816,N_4586);
or U6747 (N_6747,N_4361,N_4981);
or U6748 (N_6748,N_4475,N_5978);
or U6749 (N_6749,N_5346,N_4568);
nor U6750 (N_6750,N_5212,N_4843);
or U6751 (N_6751,N_4317,N_5556);
nor U6752 (N_6752,N_4196,N_5950);
nor U6753 (N_6753,N_5276,N_5302);
and U6754 (N_6754,N_4921,N_4322);
nand U6755 (N_6755,N_5412,N_4451);
and U6756 (N_6756,N_4646,N_5875);
xor U6757 (N_6757,N_5252,N_5670);
xor U6758 (N_6758,N_4935,N_5085);
xor U6759 (N_6759,N_5483,N_4394);
and U6760 (N_6760,N_4895,N_4406);
or U6761 (N_6761,N_4072,N_4417);
or U6762 (N_6762,N_4261,N_4386);
xnor U6763 (N_6763,N_4375,N_5489);
nand U6764 (N_6764,N_5804,N_5287);
or U6765 (N_6765,N_5126,N_4501);
and U6766 (N_6766,N_5434,N_5971);
xor U6767 (N_6767,N_5769,N_4409);
and U6768 (N_6768,N_5691,N_5161);
or U6769 (N_6769,N_4119,N_4100);
nand U6770 (N_6770,N_5715,N_4528);
nor U6771 (N_6771,N_4789,N_4183);
xnor U6772 (N_6772,N_4908,N_4097);
xnor U6773 (N_6773,N_5093,N_5242);
and U6774 (N_6774,N_5224,N_4923);
xor U6775 (N_6775,N_4389,N_5043);
xor U6776 (N_6776,N_5082,N_4329);
nand U6777 (N_6777,N_4230,N_4297);
nor U6778 (N_6778,N_4714,N_5036);
nand U6779 (N_6779,N_5202,N_5529);
and U6780 (N_6780,N_4037,N_5278);
and U6781 (N_6781,N_5995,N_4425);
or U6782 (N_6782,N_4372,N_5178);
nand U6783 (N_6783,N_4436,N_4889);
or U6784 (N_6784,N_5983,N_5850);
nand U6785 (N_6785,N_4342,N_5507);
and U6786 (N_6786,N_4433,N_5416);
or U6787 (N_6787,N_5506,N_5959);
or U6788 (N_6788,N_5235,N_5790);
xnor U6789 (N_6789,N_4625,N_5543);
and U6790 (N_6790,N_4122,N_4338);
xnor U6791 (N_6791,N_4803,N_4392);
nor U6792 (N_6792,N_4666,N_4130);
xor U6793 (N_6793,N_5729,N_4973);
xor U6794 (N_6794,N_4963,N_5697);
and U6795 (N_6795,N_4962,N_4040);
or U6796 (N_6796,N_5369,N_4068);
nor U6797 (N_6797,N_5421,N_5399);
and U6798 (N_6798,N_4627,N_4469);
nor U6799 (N_6799,N_4777,N_5720);
nand U6800 (N_6800,N_5538,N_4984);
nor U6801 (N_6801,N_5184,N_4707);
nand U6802 (N_6802,N_5297,N_4365);
or U6803 (N_6803,N_5605,N_5347);
or U6804 (N_6804,N_4758,N_5722);
and U6805 (N_6805,N_5096,N_4337);
nand U6806 (N_6806,N_5509,N_4403);
xnor U6807 (N_6807,N_4912,N_4102);
xnor U6808 (N_6808,N_5032,N_4143);
or U6809 (N_6809,N_4853,N_4292);
or U6810 (N_6810,N_4414,N_5954);
nand U6811 (N_6811,N_4295,N_5024);
or U6812 (N_6812,N_5319,N_5878);
or U6813 (N_6813,N_4980,N_5259);
or U6814 (N_6814,N_5385,N_4111);
xnor U6815 (N_6815,N_5482,N_5128);
or U6816 (N_6816,N_4644,N_5865);
nand U6817 (N_6817,N_4383,N_5141);
nand U6818 (N_6818,N_4180,N_5461);
nand U6819 (N_6819,N_4616,N_4121);
xnor U6820 (N_6820,N_4978,N_4285);
xor U6821 (N_6821,N_5703,N_5899);
and U6822 (N_6822,N_4622,N_5309);
nand U6823 (N_6823,N_4544,N_4948);
nor U6824 (N_6824,N_4363,N_4684);
and U6825 (N_6825,N_5912,N_4209);
or U6826 (N_6826,N_4879,N_4829);
xor U6827 (N_6827,N_5673,N_4489);
xor U6828 (N_6828,N_5201,N_4678);
nand U6829 (N_6829,N_5092,N_5028);
nand U6830 (N_6830,N_4991,N_4221);
xnor U6831 (N_6831,N_4393,N_5349);
and U6832 (N_6832,N_5365,N_4651);
nor U6833 (N_6833,N_5386,N_5530);
xnor U6834 (N_6834,N_4560,N_5524);
xor U6835 (N_6835,N_5197,N_4128);
nand U6836 (N_6836,N_4498,N_5756);
nand U6837 (N_6837,N_5994,N_5898);
and U6838 (N_6838,N_5446,N_5246);
nor U6839 (N_6839,N_5171,N_5807);
or U6840 (N_6840,N_5406,N_4591);
nor U6841 (N_6841,N_4115,N_5621);
and U6842 (N_6842,N_5037,N_5108);
nand U6843 (N_6843,N_5620,N_4551);
and U6844 (N_6844,N_4953,N_5528);
nand U6845 (N_6845,N_5225,N_5517);
nand U6846 (N_6846,N_5765,N_4709);
nor U6847 (N_6847,N_4056,N_4348);
nor U6848 (N_6848,N_4174,N_5592);
or U6849 (N_6849,N_5767,N_4175);
nor U6850 (N_6850,N_5193,N_5972);
nand U6851 (N_6851,N_5077,N_4515);
xnor U6852 (N_6852,N_4134,N_5263);
nor U6853 (N_6853,N_5752,N_5262);
xnor U6854 (N_6854,N_4982,N_5936);
or U6855 (N_6855,N_5874,N_5970);
nor U6856 (N_6856,N_4763,N_5721);
nand U6857 (N_6857,N_4310,N_5634);
xor U6858 (N_6858,N_5825,N_4149);
nand U6859 (N_6859,N_4291,N_5051);
nor U6860 (N_6860,N_4293,N_4324);
xor U6861 (N_6861,N_5110,N_5236);
and U6862 (N_6862,N_4391,N_5780);
and U6863 (N_6863,N_4831,N_5396);
and U6864 (N_6864,N_5109,N_5701);
nor U6865 (N_6865,N_5190,N_4467);
and U6866 (N_6866,N_5587,N_5100);
and U6867 (N_6867,N_4479,N_5676);
and U6868 (N_6868,N_5408,N_5922);
nor U6869 (N_6869,N_5854,N_4932);
nor U6870 (N_6870,N_4474,N_5745);
or U6871 (N_6871,N_5562,N_5996);
nor U6872 (N_6872,N_5432,N_5249);
nor U6873 (N_6873,N_5580,N_4476);
nand U6874 (N_6874,N_4320,N_5469);
and U6875 (N_6875,N_4506,N_5987);
and U6876 (N_6876,N_4851,N_5725);
or U6877 (N_6877,N_5247,N_5609);
xor U6878 (N_6878,N_4138,N_5626);
nor U6879 (N_6879,N_5858,N_4151);
nand U6880 (N_6880,N_4492,N_5855);
nor U6881 (N_6881,N_5284,N_4745);
xor U6882 (N_6882,N_5466,N_5410);
and U6883 (N_6883,N_4783,N_5984);
nand U6884 (N_6884,N_5732,N_4308);
nand U6885 (N_6885,N_5361,N_4061);
and U6886 (N_6886,N_4216,N_4733);
nor U6887 (N_6887,N_4062,N_4047);
and U6888 (N_6888,N_4140,N_5009);
or U6889 (N_6889,N_4918,N_5324);
xnor U6890 (N_6890,N_5041,N_4049);
xnor U6891 (N_6891,N_4841,N_5916);
nor U6892 (N_6892,N_4761,N_5480);
or U6893 (N_6893,N_4609,N_5381);
nand U6894 (N_6894,N_4070,N_5979);
nor U6895 (N_6895,N_4228,N_5822);
or U6896 (N_6896,N_4067,N_4482);
or U6897 (N_6897,N_5351,N_4736);
and U6898 (N_6898,N_5370,N_5659);
nand U6899 (N_6899,N_5271,N_5600);
nor U6900 (N_6900,N_4695,N_5980);
and U6901 (N_6901,N_5553,N_5544);
nand U6902 (N_6902,N_4504,N_4822);
xor U6903 (N_6903,N_4936,N_5602);
and U6904 (N_6904,N_4598,N_5125);
nand U6905 (N_6905,N_4795,N_5248);
nand U6906 (N_6906,N_5465,N_4866);
nand U6907 (N_6907,N_4817,N_5895);
nand U6908 (N_6908,N_4048,N_4159);
xor U6909 (N_6909,N_4024,N_5612);
or U6910 (N_6910,N_5867,N_4305);
nand U6911 (N_6911,N_4007,N_4178);
and U6912 (N_6912,N_4075,N_4090);
nand U6913 (N_6913,N_5343,N_4220);
xnor U6914 (N_6914,N_4785,N_5206);
or U6915 (N_6915,N_4925,N_5739);
or U6916 (N_6916,N_4604,N_5766);
or U6917 (N_6917,N_5714,N_5438);
xnor U6918 (N_6918,N_4996,N_4395);
nand U6919 (N_6919,N_4679,N_4529);
or U6920 (N_6920,N_4113,N_5211);
xor U6921 (N_6921,N_5596,N_4205);
or U6922 (N_6922,N_5014,N_4762);
nor U6923 (N_6923,N_4063,N_4890);
or U6924 (N_6924,N_4574,N_4065);
and U6925 (N_6925,N_4960,N_5967);
xor U6926 (N_6926,N_4776,N_4673);
and U6927 (N_6927,N_4247,N_4082);
or U6928 (N_6928,N_4050,N_4170);
xor U6929 (N_6929,N_5325,N_5707);
or U6930 (N_6930,N_4429,N_4256);
nor U6931 (N_6931,N_4585,N_5651);
and U6932 (N_6932,N_4729,N_5977);
xnor U6933 (N_6933,N_4369,N_4472);
xnor U6934 (N_6934,N_5183,N_4446);
or U6935 (N_6935,N_5545,N_5762);
nor U6936 (N_6936,N_4364,N_5719);
and U6937 (N_6937,N_5310,N_5222);
nor U6938 (N_6938,N_4214,N_5669);
nor U6939 (N_6939,N_4432,N_4874);
nand U6940 (N_6940,N_5740,N_4356);
xnor U6941 (N_6941,N_5008,N_4550);
xor U6942 (N_6942,N_5639,N_5961);
or U6943 (N_6943,N_4188,N_4043);
or U6944 (N_6944,N_5860,N_5035);
and U6945 (N_6945,N_4582,N_4631);
or U6946 (N_6946,N_5548,N_4264);
and U6947 (N_6947,N_4601,N_4583);
xor U6948 (N_6948,N_4863,N_4017);
or U6949 (N_6949,N_5734,N_4746);
xnor U6950 (N_6950,N_5176,N_4906);
nor U6951 (N_6951,N_5678,N_4633);
or U6952 (N_6952,N_4355,N_5664);
and U6953 (N_6953,N_4522,N_5575);
or U6954 (N_6954,N_5693,N_4422);
nand U6955 (N_6955,N_5367,N_4300);
nor U6956 (N_6956,N_4955,N_4664);
nor U6957 (N_6957,N_4788,N_4513);
nand U6958 (N_6958,N_4278,N_4741);
nand U6959 (N_6959,N_5337,N_5785);
nand U6960 (N_6960,N_5914,N_5559);
nand U6961 (N_6961,N_5172,N_5494);
xor U6962 (N_6962,N_5915,N_5428);
or U6963 (N_6963,N_5462,N_5040);
xnor U6964 (N_6964,N_5809,N_5787);
xnor U6965 (N_6965,N_4211,N_4848);
nand U6966 (N_6966,N_5447,N_4699);
and U6967 (N_6967,N_5628,N_4907);
or U6968 (N_6968,N_4192,N_4654);
and U6969 (N_6969,N_5433,N_5731);
nand U6970 (N_6970,N_4427,N_4011);
or U6971 (N_6971,N_5827,N_4685);
xnor U6972 (N_6972,N_5233,N_5940);
nand U6973 (N_6973,N_5444,N_5578);
nor U6974 (N_6974,N_4168,N_4473);
or U6975 (N_6975,N_4882,N_5106);
xor U6976 (N_6976,N_4058,N_5188);
and U6977 (N_6977,N_4530,N_5778);
or U6978 (N_6978,N_5377,N_4144);
and U6979 (N_6979,N_4463,N_4883);
or U6980 (N_6980,N_4959,N_5397);
nand U6981 (N_6981,N_5395,N_5642);
nand U6982 (N_6982,N_4108,N_4020);
nor U6983 (N_6983,N_5500,N_4837);
nor U6984 (N_6984,N_4284,N_5604);
and U6985 (N_6985,N_5761,N_5376);
nor U6986 (N_6986,N_5332,N_5777);
nor U6987 (N_6987,N_5342,N_4751);
and U6988 (N_6988,N_5911,N_5811);
xnor U6989 (N_6989,N_5917,N_5564);
xor U6990 (N_6990,N_4894,N_4237);
and U6991 (N_6991,N_5650,N_5356);
nor U6992 (N_6992,N_5868,N_4562);
xor U6993 (N_6993,N_5974,N_5072);
and U6994 (N_6994,N_4842,N_4301);
nor U6995 (N_6995,N_5328,N_5986);
or U6996 (N_6996,N_4579,N_4610);
or U6997 (N_6997,N_5694,N_4025);
and U6998 (N_6998,N_5799,N_5239);
xor U6999 (N_6999,N_5616,N_5594);
nand U7000 (N_7000,N_5776,N_5528);
nor U7001 (N_7001,N_5959,N_4134);
nor U7002 (N_7002,N_4558,N_5004);
nor U7003 (N_7003,N_5730,N_4715);
nor U7004 (N_7004,N_5660,N_4268);
and U7005 (N_7005,N_4089,N_5872);
nor U7006 (N_7006,N_4354,N_5650);
or U7007 (N_7007,N_5128,N_5305);
nor U7008 (N_7008,N_4981,N_5551);
and U7009 (N_7009,N_4670,N_5385);
nor U7010 (N_7010,N_5111,N_4920);
nand U7011 (N_7011,N_4582,N_5901);
nand U7012 (N_7012,N_5598,N_4939);
nand U7013 (N_7013,N_5482,N_5811);
nor U7014 (N_7014,N_5420,N_4896);
xor U7015 (N_7015,N_4502,N_5510);
and U7016 (N_7016,N_5334,N_5710);
xor U7017 (N_7017,N_5777,N_4930);
nor U7018 (N_7018,N_4898,N_4471);
nor U7019 (N_7019,N_5938,N_4598);
nand U7020 (N_7020,N_5447,N_4628);
and U7021 (N_7021,N_4915,N_4265);
xor U7022 (N_7022,N_4282,N_4986);
nand U7023 (N_7023,N_5293,N_4399);
xor U7024 (N_7024,N_5431,N_4306);
nor U7025 (N_7025,N_4369,N_5936);
or U7026 (N_7026,N_5727,N_5075);
nand U7027 (N_7027,N_5176,N_4311);
nand U7028 (N_7028,N_5953,N_4899);
or U7029 (N_7029,N_4264,N_4335);
nand U7030 (N_7030,N_4683,N_5052);
nand U7031 (N_7031,N_5122,N_5469);
xnor U7032 (N_7032,N_5249,N_4546);
nor U7033 (N_7033,N_4778,N_5827);
and U7034 (N_7034,N_5320,N_5080);
and U7035 (N_7035,N_5737,N_5994);
and U7036 (N_7036,N_5872,N_4266);
nand U7037 (N_7037,N_4533,N_4564);
xor U7038 (N_7038,N_4873,N_5332);
or U7039 (N_7039,N_5903,N_4906);
xnor U7040 (N_7040,N_4386,N_4091);
nand U7041 (N_7041,N_5248,N_5608);
nor U7042 (N_7042,N_5610,N_4165);
nor U7043 (N_7043,N_5877,N_4150);
nand U7044 (N_7044,N_4206,N_4010);
xor U7045 (N_7045,N_4625,N_5113);
nand U7046 (N_7046,N_5671,N_4694);
nand U7047 (N_7047,N_4207,N_4964);
or U7048 (N_7048,N_4188,N_4920);
nor U7049 (N_7049,N_4382,N_5569);
and U7050 (N_7050,N_4641,N_5309);
xnor U7051 (N_7051,N_4868,N_5831);
or U7052 (N_7052,N_5756,N_4388);
and U7053 (N_7053,N_4020,N_5702);
and U7054 (N_7054,N_5116,N_4309);
xor U7055 (N_7055,N_5438,N_4066);
or U7056 (N_7056,N_5078,N_5933);
xnor U7057 (N_7057,N_5853,N_5673);
nor U7058 (N_7058,N_4833,N_5901);
and U7059 (N_7059,N_4011,N_4042);
or U7060 (N_7060,N_5619,N_5539);
or U7061 (N_7061,N_4813,N_4258);
and U7062 (N_7062,N_5217,N_4550);
xor U7063 (N_7063,N_4112,N_4309);
or U7064 (N_7064,N_5513,N_5039);
and U7065 (N_7065,N_4352,N_4881);
nand U7066 (N_7066,N_4673,N_5975);
or U7067 (N_7067,N_4893,N_4178);
nor U7068 (N_7068,N_4366,N_5236);
xnor U7069 (N_7069,N_5274,N_5794);
nand U7070 (N_7070,N_4900,N_4846);
and U7071 (N_7071,N_5187,N_5884);
nor U7072 (N_7072,N_4570,N_5690);
nor U7073 (N_7073,N_4707,N_4152);
or U7074 (N_7074,N_5981,N_5305);
nand U7075 (N_7075,N_4953,N_5097);
nand U7076 (N_7076,N_5969,N_5274);
or U7077 (N_7077,N_5213,N_5340);
nor U7078 (N_7078,N_5952,N_5545);
xor U7079 (N_7079,N_4794,N_4760);
xnor U7080 (N_7080,N_5894,N_5366);
or U7081 (N_7081,N_5558,N_4462);
xor U7082 (N_7082,N_4683,N_4094);
nand U7083 (N_7083,N_5085,N_4972);
nand U7084 (N_7084,N_5996,N_4472);
or U7085 (N_7085,N_4233,N_5060);
xnor U7086 (N_7086,N_5749,N_4995);
xor U7087 (N_7087,N_4781,N_5963);
nand U7088 (N_7088,N_5500,N_5792);
nor U7089 (N_7089,N_5109,N_4778);
xnor U7090 (N_7090,N_5097,N_5160);
or U7091 (N_7091,N_5132,N_5687);
nand U7092 (N_7092,N_4291,N_5841);
xor U7093 (N_7093,N_4749,N_4239);
nor U7094 (N_7094,N_5198,N_4274);
or U7095 (N_7095,N_4734,N_5676);
or U7096 (N_7096,N_4437,N_4065);
nor U7097 (N_7097,N_4031,N_5504);
nor U7098 (N_7098,N_4220,N_4552);
nand U7099 (N_7099,N_4104,N_4723);
and U7100 (N_7100,N_4978,N_5764);
nor U7101 (N_7101,N_5604,N_4920);
nand U7102 (N_7102,N_4504,N_5049);
xnor U7103 (N_7103,N_5198,N_5511);
and U7104 (N_7104,N_5250,N_4104);
or U7105 (N_7105,N_4711,N_4853);
nor U7106 (N_7106,N_5315,N_5669);
and U7107 (N_7107,N_5707,N_4092);
nand U7108 (N_7108,N_4845,N_5139);
nor U7109 (N_7109,N_4892,N_5318);
xor U7110 (N_7110,N_4643,N_4595);
nand U7111 (N_7111,N_4263,N_5759);
nand U7112 (N_7112,N_4158,N_4077);
or U7113 (N_7113,N_5712,N_5321);
nand U7114 (N_7114,N_4949,N_4006);
nor U7115 (N_7115,N_4697,N_5978);
nor U7116 (N_7116,N_4111,N_5189);
xor U7117 (N_7117,N_5095,N_5011);
or U7118 (N_7118,N_4295,N_5213);
and U7119 (N_7119,N_4114,N_5234);
nor U7120 (N_7120,N_4087,N_4038);
or U7121 (N_7121,N_4786,N_4209);
nand U7122 (N_7122,N_5378,N_5253);
nand U7123 (N_7123,N_5067,N_5439);
and U7124 (N_7124,N_4685,N_4385);
nand U7125 (N_7125,N_5246,N_4741);
or U7126 (N_7126,N_4047,N_5024);
nor U7127 (N_7127,N_5902,N_4834);
nand U7128 (N_7128,N_4965,N_5762);
or U7129 (N_7129,N_5745,N_5550);
or U7130 (N_7130,N_5819,N_5034);
nor U7131 (N_7131,N_5032,N_5390);
or U7132 (N_7132,N_5168,N_4918);
and U7133 (N_7133,N_5066,N_4194);
xor U7134 (N_7134,N_4661,N_4859);
xor U7135 (N_7135,N_4563,N_5355);
nor U7136 (N_7136,N_4523,N_5209);
or U7137 (N_7137,N_4025,N_5173);
and U7138 (N_7138,N_5217,N_4733);
nand U7139 (N_7139,N_4244,N_4329);
nand U7140 (N_7140,N_4196,N_5151);
and U7141 (N_7141,N_4908,N_4948);
nor U7142 (N_7142,N_4105,N_5303);
nor U7143 (N_7143,N_4003,N_4961);
xor U7144 (N_7144,N_5287,N_5781);
nor U7145 (N_7145,N_4764,N_4970);
nor U7146 (N_7146,N_4167,N_4273);
or U7147 (N_7147,N_4743,N_4872);
nor U7148 (N_7148,N_4008,N_5553);
and U7149 (N_7149,N_5413,N_5341);
and U7150 (N_7150,N_4878,N_4469);
or U7151 (N_7151,N_4679,N_5798);
nor U7152 (N_7152,N_4872,N_4356);
xor U7153 (N_7153,N_4438,N_4359);
or U7154 (N_7154,N_4525,N_4604);
or U7155 (N_7155,N_4297,N_4324);
or U7156 (N_7156,N_4925,N_5480);
xnor U7157 (N_7157,N_5710,N_4283);
xor U7158 (N_7158,N_4900,N_4531);
xnor U7159 (N_7159,N_4652,N_5266);
and U7160 (N_7160,N_5846,N_5005);
or U7161 (N_7161,N_5927,N_5596);
nand U7162 (N_7162,N_5471,N_4436);
nor U7163 (N_7163,N_4843,N_4677);
nand U7164 (N_7164,N_4437,N_5815);
or U7165 (N_7165,N_4519,N_5916);
nor U7166 (N_7166,N_4373,N_4768);
nand U7167 (N_7167,N_5908,N_4082);
nor U7168 (N_7168,N_5423,N_5837);
and U7169 (N_7169,N_5009,N_4432);
nand U7170 (N_7170,N_5341,N_5471);
nand U7171 (N_7171,N_5453,N_4061);
and U7172 (N_7172,N_4400,N_5820);
and U7173 (N_7173,N_5645,N_5985);
nand U7174 (N_7174,N_4918,N_5108);
nor U7175 (N_7175,N_4781,N_5153);
or U7176 (N_7176,N_4364,N_5922);
xnor U7177 (N_7177,N_4888,N_4655);
nor U7178 (N_7178,N_4172,N_5770);
nor U7179 (N_7179,N_4183,N_5538);
nor U7180 (N_7180,N_5545,N_5276);
nand U7181 (N_7181,N_4723,N_5481);
nand U7182 (N_7182,N_4784,N_5292);
and U7183 (N_7183,N_4710,N_5856);
nand U7184 (N_7184,N_4207,N_5466);
xnor U7185 (N_7185,N_5377,N_5910);
or U7186 (N_7186,N_4716,N_4055);
nand U7187 (N_7187,N_4747,N_5641);
nor U7188 (N_7188,N_5324,N_4358);
nor U7189 (N_7189,N_5287,N_5511);
and U7190 (N_7190,N_5474,N_5894);
xnor U7191 (N_7191,N_5026,N_5600);
nor U7192 (N_7192,N_5106,N_5868);
or U7193 (N_7193,N_5332,N_4176);
and U7194 (N_7194,N_5603,N_4386);
nand U7195 (N_7195,N_4942,N_4360);
xnor U7196 (N_7196,N_5173,N_4410);
nand U7197 (N_7197,N_4433,N_5539);
or U7198 (N_7198,N_5277,N_5283);
nand U7199 (N_7199,N_5763,N_5934);
xor U7200 (N_7200,N_4410,N_5137);
or U7201 (N_7201,N_5988,N_5548);
nand U7202 (N_7202,N_5793,N_5310);
and U7203 (N_7203,N_4654,N_5375);
nand U7204 (N_7204,N_4071,N_4949);
or U7205 (N_7205,N_5687,N_5623);
xor U7206 (N_7206,N_4539,N_4344);
xor U7207 (N_7207,N_5205,N_4583);
xor U7208 (N_7208,N_5943,N_4599);
and U7209 (N_7209,N_5889,N_4949);
nor U7210 (N_7210,N_5588,N_4331);
xor U7211 (N_7211,N_5585,N_4172);
xnor U7212 (N_7212,N_5113,N_5384);
nand U7213 (N_7213,N_4020,N_5021);
or U7214 (N_7214,N_4782,N_5459);
or U7215 (N_7215,N_4305,N_4536);
nand U7216 (N_7216,N_5901,N_5460);
nand U7217 (N_7217,N_5403,N_4750);
nand U7218 (N_7218,N_4281,N_4410);
or U7219 (N_7219,N_5527,N_4574);
and U7220 (N_7220,N_4719,N_4916);
nor U7221 (N_7221,N_5848,N_4320);
nand U7222 (N_7222,N_4768,N_5991);
or U7223 (N_7223,N_5960,N_5041);
nor U7224 (N_7224,N_5867,N_4102);
or U7225 (N_7225,N_4593,N_4569);
or U7226 (N_7226,N_4543,N_5373);
and U7227 (N_7227,N_4730,N_4027);
and U7228 (N_7228,N_5410,N_5272);
nor U7229 (N_7229,N_5385,N_4831);
nand U7230 (N_7230,N_5870,N_5320);
or U7231 (N_7231,N_4503,N_5057);
nor U7232 (N_7232,N_5454,N_5040);
nand U7233 (N_7233,N_5218,N_4685);
or U7234 (N_7234,N_4120,N_5945);
xnor U7235 (N_7235,N_4960,N_4976);
or U7236 (N_7236,N_5877,N_4145);
or U7237 (N_7237,N_5732,N_5467);
or U7238 (N_7238,N_5281,N_4209);
nand U7239 (N_7239,N_5545,N_5029);
and U7240 (N_7240,N_4688,N_4570);
and U7241 (N_7241,N_5799,N_4953);
or U7242 (N_7242,N_4722,N_5134);
xnor U7243 (N_7243,N_5317,N_4280);
nand U7244 (N_7244,N_5137,N_4379);
and U7245 (N_7245,N_5599,N_4521);
or U7246 (N_7246,N_5188,N_4555);
nand U7247 (N_7247,N_4098,N_4615);
nand U7248 (N_7248,N_5010,N_5377);
nand U7249 (N_7249,N_4703,N_5670);
nor U7250 (N_7250,N_4407,N_5520);
and U7251 (N_7251,N_4295,N_5825);
xnor U7252 (N_7252,N_4754,N_5836);
xnor U7253 (N_7253,N_5914,N_5334);
xnor U7254 (N_7254,N_4149,N_5212);
xnor U7255 (N_7255,N_5911,N_4136);
nand U7256 (N_7256,N_4443,N_5290);
or U7257 (N_7257,N_5092,N_4556);
nand U7258 (N_7258,N_4340,N_4713);
nand U7259 (N_7259,N_5414,N_4648);
nand U7260 (N_7260,N_5576,N_4095);
and U7261 (N_7261,N_4982,N_5379);
xor U7262 (N_7262,N_5073,N_5080);
or U7263 (N_7263,N_5812,N_5423);
and U7264 (N_7264,N_5466,N_4017);
xor U7265 (N_7265,N_4457,N_4603);
nor U7266 (N_7266,N_5407,N_4601);
nand U7267 (N_7267,N_5728,N_4489);
or U7268 (N_7268,N_5925,N_5513);
nand U7269 (N_7269,N_4190,N_4827);
xnor U7270 (N_7270,N_5785,N_4064);
nor U7271 (N_7271,N_4599,N_5713);
nor U7272 (N_7272,N_4477,N_4017);
xnor U7273 (N_7273,N_5540,N_5025);
or U7274 (N_7274,N_4296,N_4644);
nor U7275 (N_7275,N_4355,N_5231);
nor U7276 (N_7276,N_5298,N_4621);
or U7277 (N_7277,N_4624,N_4994);
or U7278 (N_7278,N_4031,N_4564);
and U7279 (N_7279,N_4685,N_5412);
or U7280 (N_7280,N_5606,N_4170);
xor U7281 (N_7281,N_5617,N_4528);
or U7282 (N_7282,N_5608,N_5452);
or U7283 (N_7283,N_5604,N_5145);
xnor U7284 (N_7284,N_4655,N_5935);
or U7285 (N_7285,N_4318,N_4686);
or U7286 (N_7286,N_4172,N_5587);
nand U7287 (N_7287,N_4003,N_5172);
nand U7288 (N_7288,N_5889,N_5594);
and U7289 (N_7289,N_4457,N_5395);
nor U7290 (N_7290,N_5240,N_4814);
nand U7291 (N_7291,N_4857,N_5225);
nor U7292 (N_7292,N_5105,N_5543);
nor U7293 (N_7293,N_5024,N_5036);
and U7294 (N_7294,N_4948,N_4319);
xnor U7295 (N_7295,N_4802,N_5114);
xor U7296 (N_7296,N_4590,N_5563);
and U7297 (N_7297,N_4547,N_5915);
nor U7298 (N_7298,N_5895,N_5707);
or U7299 (N_7299,N_4588,N_5476);
nor U7300 (N_7300,N_4242,N_5701);
xor U7301 (N_7301,N_5920,N_4174);
or U7302 (N_7302,N_5329,N_5189);
nand U7303 (N_7303,N_4076,N_4921);
nand U7304 (N_7304,N_5031,N_4215);
xnor U7305 (N_7305,N_5782,N_4024);
nand U7306 (N_7306,N_5049,N_4122);
or U7307 (N_7307,N_4135,N_5266);
or U7308 (N_7308,N_5156,N_5261);
nor U7309 (N_7309,N_5565,N_4568);
or U7310 (N_7310,N_5231,N_5874);
nor U7311 (N_7311,N_4373,N_5459);
xnor U7312 (N_7312,N_5311,N_4742);
nor U7313 (N_7313,N_5589,N_5769);
or U7314 (N_7314,N_5656,N_5826);
nand U7315 (N_7315,N_4264,N_5073);
xnor U7316 (N_7316,N_4484,N_4024);
xor U7317 (N_7317,N_5649,N_4184);
nor U7318 (N_7318,N_5173,N_4848);
and U7319 (N_7319,N_5923,N_4349);
or U7320 (N_7320,N_4015,N_4091);
xnor U7321 (N_7321,N_5604,N_4238);
xor U7322 (N_7322,N_5867,N_4303);
or U7323 (N_7323,N_5953,N_5714);
nand U7324 (N_7324,N_5626,N_5669);
nand U7325 (N_7325,N_4700,N_4953);
nor U7326 (N_7326,N_5000,N_4938);
xor U7327 (N_7327,N_5355,N_4281);
nand U7328 (N_7328,N_5206,N_5184);
nand U7329 (N_7329,N_5468,N_4596);
and U7330 (N_7330,N_5247,N_5642);
xnor U7331 (N_7331,N_5779,N_5735);
nor U7332 (N_7332,N_4612,N_5997);
nand U7333 (N_7333,N_4193,N_5341);
or U7334 (N_7334,N_4302,N_5841);
or U7335 (N_7335,N_4136,N_5865);
nor U7336 (N_7336,N_5385,N_4042);
xnor U7337 (N_7337,N_5510,N_5873);
nor U7338 (N_7338,N_4440,N_4187);
nor U7339 (N_7339,N_5329,N_4240);
and U7340 (N_7340,N_4353,N_5191);
nor U7341 (N_7341,N_5749,N_4547);
nand U7342 (N_7342,N_5229,N_4670);
xor U7343 (N_7343,N_5298,N_4025);
and U7344 (N_7344,N_5715,N_5258);
xnor U7345 (N_7345,N_5128,N_5693);
xor U7346 (N_7346,N_4210,N_4573);
nor U7347 (N_7347,N_5289,N_5802);
xnor U7348 (N_7348,N_5372,N_4053);
or U7349 (N_7349,N_4989,N_4393);
xnor U7350 (N_7350,N_4480,N_4595);
or U7351 (N_7351,N_4133,N_5453);
nor U7352 (N_7352,N_4518,N_4523);
nor U7353 (N_7353,N_5643,N_5226);
or U7354 (N_7354,N_5186,N_5966);
nor U7355 (N_7355,N_5958,N_4390);
nand U7356 (N_7356,N_4613,N_4365);
nor U7357 (N_7357,N_4050,N_4237);
xor U7358 (N_7358,N_4111,N_5480);
and U7359 (N_7359,N_4361,N_4876);
or U7360 (N_7360,N_5109,N_4370);
and U7361 (N_7361,N_4901,N_5982);
nand U7362 (N_7362,N_5246,N_4441);
xnor U7363 (N_7363,N_5670,N_4327);
xnor U7364 (N_7364,N_4108,N_4728);
or U7365 (N_7365,N_4515,N_4900);
nand U7366 (N_7366,N_4869,N_4635);
and U7367 (N_7367,N_5476,N_5311);
or U7368 (N_7368,N_5973,N_5712);
nand U7369 (N_7369,N_4720,N_4064);
nand U7370 (N_7370,N_5894,N_5454);
or U7371 (N_7371,N_5210,N_5444);
or U7372 (N_7372,N_5268,N_5730);
xor U7373 (N_7373,N_5639,N_4145);
nand U7374 (N_7374,N_4596,N_4209);
and U7375 (N_7375,N_5260,N_5198);
xor U7376 (N_7376,N_5431,N_5982);
xnor U7377 (N_7377,N_4562,N_4577);
nor U7378 (N_7378,N_5676,N_5019);
nor U7379 (N_7379,N_5405,N_5577);
xnor U7380 (N_7380,N_5545,N_4736);
nor U7381 (N_7381,N_4856,N_5927);
and U7382 (N_7382,N_5890,N_4863);
or U7383 (N_7383,N_5069,N_4345);
and U7384 (N_7384,N_4842,N_5709);
xor U7385 (N_7385,N_5102,N_4133);
nand U7386 (N_7386,N_5841,N_4124);
xnor U7387 (N_7387,N_4190,N_4660);
and U7388 (N_7388,N_5447,N_4348);
or U7389 (N_7389,N_4775,N_4428);
or U7390 (N_7390,N_4376,N_5893);
xor U7391 (N_7391,N_4875,N_4016);
or U7392 (N_7392,N_5805,N_5692);
nor U7393 (N_7393,N_5585,N_4173);
or U7394 (N_7394,N_5540,N_4877);
or U7395 (N_7395,N_4775,N_4562);
or U7396 (N_7396,N_5429,N_5301);
or U7397 (N_7397,N_4488,N_5977);
and U7398 (N_7398,N_4821,N_5003);
or U7399 (N_7399,N_4860,N_5223);
nor U7400 (N_7400,N_4247,N_5238);
xnor U7401 (N_7401,N_4285,N_5124);
xor U7402 (N_7402,N_5189,N_5394);
or U7403 (N_7403,N_5046,N_5084);
and U7404 (N_7404,N_4077,N_5869);
nor U7405 (N_7405,N_4087,N_4547);
nor U7406 (N_7406,N_5696,N_4018);
xnor U7407 (N_7407,N_5649,N_4224);
nor U7408 (N_7408,N_5314,N_5333);
or U7409 (N_7409,N_4730,N_5363);
nand U7410 (N_7410,N_4005,N_5753);
xnor U7411 (N_7411,N_5439,N_4419);
nand U7412 (N_7412,N_4594,N_4444);
xnor U7413 (N_7413,N_4819,N_5181);
or U7414 (N_7414,N_4071,N_5139);
or U7415 (N_7415,N_4362,N_4082);
and U7416 (N_7416,N_4956,N_4740);
nand U7417 (N_7417,N_5880,N_5097);
xor U7418 (N_7418,N_5846,N_4422);
or U7419 (N_7419,N_5956,N_4015);
nor U7420 (N_7420,N_5648,N_4753);
nand U7421 (N_7421,N_5592,N_4112);
nor U7422 (N_7422,N_5557,N_4849);
or U7423 (N_7423,N_5402,N_4688);
and U7424 (N_7424,N_5309,N_4167);
xnor U7425 (N_7425,N_5324,N_5095);
xnor U7426 (N_7426,N_4540,N_4173);
nand U7427 (N_7427,N_4567,N_5428);
or U7428 (N_7428,N_4668,N_4335);
and U7429 (N_7429,N_4589,N_5203);
nor U7430 (N_7430,N_4374,N_4567);
xor U7431 (N_7431,N_5612,N_5050);
nor U7432 (N_7432,N_4631,N_4139);
or U7433 (N_7433,N_5006,N_5869);
and U7434 (N_7434,N_4421,N_5565);
and U7435 (N_7435,N_5226,N_4341);
nor U7436 (N_7436,N_4643,N_5660);
or U7437 (N_7437,N_4712,N_4480);
and U7438 (N_7438,N_5690,N_4678);
or U7439 (N_7439,N_4067,N_4877);
xnor U7440 (N_7440,N_5598,N_5821);
or U7441 (N_7441,N_4027,N_4866);
nand U7442 (N_7442,N_4176,N_5275);
xor U7443 (N_7443,N_4641,N_4698);
and U7444 (N_7444,N_4866,N_5688);
nor U7445 (N_7445,N_4363,N_5037);
nor U7446 (N_7446,N_5390,N_5601);
nor U7447 (N_7447,N_4949,N_4925);
nand U7448 (N_7448,N_4345,N_5281);
nor U7449 (N_7449,N_5302,N_5067);
or U7450 (N_7450,N_5348,N_5158);
nand U7451 (N_7451,N_4192,N_5109);
nand U7452 (N_7452,N_5580,N_4050);
xnor U7453 (N_7453,N_4502,N_4217);
nor U7454 (N_7454,N_4464,N_5459);
and U7455 (N_7455,N_4011,N_4975);
or U7456 (N_7456,N_5807,N_4068);
nand U7457 (N_7457,N_5422,N_5203);
nor U7458 (N_7458,N_4820,N_5025);
and U7459 (N_7459,N_4822,N_5339);
and U7460 (N_7460,N_4203,N_4957);
nor U7461 (N_7461,N_4228,N_4345);
nor U7462 (N_7462,N_4434,N_4384);
nor U7463 (N_7463,N_5744,N_4063);
xnor U7464 (N_7464,N_5041,N_5277);
or U7465 (N_7465,N_5171,N_5501);
or U7466 (N_7466,N_4076,N_5379);
nand U7467 (N_7467,N_4368,N_5698);
or U7468 (N_7468,N_5028,N_4970);
and U7469 (N_7469,N_4121,N_5510);
or U7470 (N_7470,N_4117,N_5423);
xor U7471 (N_7471,N_5246,N_5496);
and U7472 (N_7472,N_4942,N_5117);
nand U7473 (N_7473,N_4230,N_4565);
or U7474 (N_7474,N_4022,N_4083);
nand U7475 (N_7475,N_4025,N_5183);
nand U7476 (N_7476,N_5057,N_5924);
or U7477 (N_7477,N_4760,N_5847);
or U7478 (N_7478,N_4997,N_4971);
nand U7479 (N_7479,N_4128,N_5274);
and U7480 (N_7480,N_4348,N_4185);
nand U7481 (N_7481,N_4554,N_4545);
and U7482 (N_7482,N_4565,N_4988);
and U7483 (N_7483,N_5633,N_5551);
and U7484 (N_7484,N_4423,N_5817);
and U7485 (N_7485,N_4326,N_5495);
xor U7486 (N_7486,N_5149,N_5854);
and U7487 (N_7487,N_5094,N_4609);
or U7488 (N_7488,N_4279,N_5768);
xnor U7489 (N_7489,N_5792,N_4514);
nor U7490 (N_7490,N_5703,N_4907);
and U7491 (N_7491,N_5550,N_4453);
nand U7492 (N_7492,N_4910,N_4228);
nand U7493 (N_7493,N_4126,N_4659);
nor U7494 (N_7494,N_5213,N_5713);
and U7495 (N_7495,N_4548,N_4903);
or U7496 (N_7496,N_4232,N_5016);
xor U7497 (N_7497,N_5539,N_4306);
or U7498 (N_7498,N_4397,N_4538);
or U7499 (N_7499,N_4645,N_5864);
xnor U7500 (N_7500,N_5323,N_4672);
and U7501 (N_7501,N_5016,N_4683);
nor U7502 (N_7502,N_5140,N_4925);
xor U7503 (N_7503,N_5801,N_5300);
or U7504 (N_7504,N_5778,N_5326);
xor U7505 (N_7505,N_4150,N_5665);
or U7506 (N_7506,N_5847,N_4775);
nand U7507 (N_7507,N_4129,N_4993);
xor U7508 (N_7508,N_5557,N_4969);
and U7509 (N_7509,N_5639,N_4970);
nand U7510 (N_7510,N_4413,N_4128);
or U7511 (N_7511,N_4873,N_5881);
nor U7512 (N_7512,N_4446,N_5515);
and U7513 (N_7513,N_4569,N_5187);
nand U7514 (N_7514,N_4693,N_5676);
xor U7515 (N_7515,N_5520,N_4664);
xor U7516 (N_7516,N_4760,N_5712);
or U7517 (N_7517,N_4473,N_4557);
xor U7518 (N_7518,N_4849,N_5269);
and U7519 (N_7519,N_4612,N_5254);
or U7520 (N_7520,N_5759,N_4770);
nor U7521 (N_7521,N_5734,N_4732);
xnor U7522 (N_7522,N_4955,N_5090);
nor U7523 (N_7523,N_4865,N_4015);
nor U7524 (N_7524,N_5404,N_4454);
and U7525 (N_7525,N_5393,N_5350);
or U7526 (N_7526,N_5765,N_5127);
xor U7527 (N_7527,N_5508,N_4316);
nand U7528 (N_7528,N_4878,N_4865);
nand U7529 (N_7529,N_5259,N_4563);
xnor U7530 (N_7530,N_4157,N_4674);
nor U7531 (N_7531,N_4910,N_4567);
or U7532 (N_7532,N_5943,N_5175);
nand U7533 (N_7533,N_5863,N_5184);
xor U7534 (N_7534,N_5227,N_4230);
nor U7535 (N_7535,N_4851,N_5185);
and U7536 (N_7536,N_5695,N_5255);
or U7537 (N_7537,N_4986,N_4151);
nand U7538 (N_7538,N_5323,N_4552);
nand U7539 (N_7539,N_4045,N_5495);
nand U7540 (N_7540,N_5519,N_5344);
and U7541 (N_7541,N_4290,N_5172);
nand U7542 (N_7542,N_4184,N_5515);
xor U7543 (N_7543,N_4403,N_4140);
nand U7544 (N_7544,N_5585,N_5875);
nor U7545 (N_7545,N_4688,N_4746);
nand U7546 (N_7546,N_5746,N_4862);
or U7547 (N_7547,N_5168,N_4558);
or U7548 (N_7548,N_5138,N_4753);
and U7549 (N_7549,N_4784,N_4984);
nor U7550 (N_7550,N_4393,N_4907);
or U7551 (N_7551,N_4553,N_5932);
nand U7552 (N_7552,N_5578,N_4094);
nor U7553 (N_7553,N_4779,N_4816);
and U7554 (N_7554,N_5218,N_5720);
and U7555 (N_7555,N_4414,N_5614);
nor U7556 (N_7556,N_4139,N_4301);
nand U7557 (N_7557,N_5545,N_4318);
nor U7558 (N_7558,N_5273,N_4477);
nand U7559 (N_7559,N_5694,N_4134);
and U7560 (N_7560,N_4209,N_5081);
or U7561 (N_7561,N_4081,N_5326);
nand U7562 (N_7562,N_5582,N_5824);
and U7563 (N_7563,N_5466,N_5238);
xnor U7564 (N_7564,N_4653,N_4345);
nand U7565 (N_7565,N_5943,N_5672);
nor U7566 (N_7566,N_5757,N_5670);
or U7567 (N_7567,N_4421,N_5527);
nor U7568 (N_7568,N_5608,N_4171);
nor U7569 (N_7569,N_5428,N_5381);
nand U7570 (N_7570,N_5355,N_5288);
xor U7571 (N_7571,N_4158,N_4317);
or U7572 (N_7572,N_5143,N_5987);
nor U7573 (N_7573,N_5075,N_4183);
and U7574 (N_7574,N_4847,N_4623);
nand U7575 (N_7575,N_4965,N_5978);
and U7576 (N_7576,N_5928,N_4467);
and U7577 (N_7577,N_4170,N_4910);
or U7578 (N_7578,N_5664,N_5582);
and U7579 (N_7579,N_4406,N_4613);
and U7580 (N_7580,N_5144,N_5153);
xor U7581 (N_7581,N_5234,N_5971);
and U7582 (N_7582,N_4121,N_4786);
nor U7583 (N_7583,N_4279,N_5594);
xnor U7584 (N_7584,N_4871,N_5148);
and U7585 (N_7585,N_5021,N_5409);
or U7586 (N_7586,N_5781,N_4083);
nor U7587 (N_7587,N_5987,N_4387);
nand U7588 (N_7588,N_4700,N_5873);
or U7589 (N_7589,N_5915,N_5305);
nand U7590 (N_7590,N_4484,N_5119);
xnor U7591 (N_7591,N_5995,N_5819);
or U7592 (N_7592,N_5381,N_5095);
nand U7593 (N_7593,N_5550,N_5653);
xnor U7594 (N_7594,N_5527,N_5351);
and U7595 (N_7595,N_4162,N_4233);
nand U7596 (N_7596,N_4129,N_4642);
nor U7597 (N_7597,N_4528,N_4826);
nand U7598 (N_7598,N_5715,N_4566);
and U7599 (N_7599,N_4358,N_4243);
and U7600 (N_7600,N_5176,N_5262);
or U7601 (N_7601,N_5120,N_4527);
or U7602 (N_7602,N_4700,N_4024);
nand U7603 (N_7603,N_5956,N_4907);
xnor U7604 (N_7604,N_5442,N_4198);
and U7605 (N_7605,N_5796,N_5272);
and U7606 (N_7606,N_4252,N_5224);
xnor U7607 (N_7607,N_5479,N_5101);
xnor U7608 (N_7608,N_4469,N_5010);
or U7609 (N_7609,N_4262,N_4727);
and U7610 (N_7610,N_4996,N_5415);
nand U7611 (N_7611,N_5825,N_5778);
nor U7612 (N_7612,N_5462,N_4820);
and U7613 (N_7613,N_4234,N_5331);
or U7614 (N_7614,N_5154,N_5651);
nor U7615 (N_7615,N_4321,N_5979);
and U7616 (N_7616,N_4663,N_4233);
xnor U7617 (N_7617,N_4499,N_4823);
or U7618 (N_7618,N_5499,N_4451);
nand U7619 (N_7619,N_4391,N_5720);
xnor U7620 (N_7620,N_4100,N_4168);
and U7621 (N_7621,N_4225,N_4592);
xnor U7622 (N_7622,N_5228,N_4098);
nor U7623 (N_7623,N_4641,N_5654);
xor U7624 (N_7624,N_5084,N_4831);
and U7625 (N_7625,N_5535,N_4995);
nor U7626 (N_7626,N_5559,N_4380);
nor U7627 (N_7627,N_4537,N_5286);
and U7628 (N_7628,N_4628,N_5196);
or U7629 (N_7629,N_4882,N_4973);
or U7630 (N_7630,N_5272,N_5798);
xor U7631 (N_7631,N_4249,N_5629);
or U7632 (N_7632,N_5744,N_5107);
nor U7633 (N_7633,N_5078,N_4250);
xnor U7634 (N_7634,N_4324,N_5982);
and U7635 (N_7635,N_5433,N_5843);
xnor U7636 (N_7636,N_5143,N_4263);
nand U7637 (N_7637,N_4131,N_5321);
or U7638 (N_7638,N_5074,N_4892);
xor U7639 (N_7639,N_5178,N_4982);
nand U7640 (N_7640,N_4499,N_4992);
nor U7641 (N_7641,N_4817,N_4915);
nand U7642 (N_7642,N_4011,N_5645);
xor U7643 (N_7643,N_4607,N_5469);
xnor U7644 (N_7644,N_4003,N_5675);
nor U7645 (N_7645,N_4074,N_4120);
or U7646 (N_7646,N_4872,N_5952);
xnor U7647 (N_7647,N_4629,N_5349);
and U7648 (N_7648,N_5787,N_4976);
nand U7649 (N_7649,N_5355,N_5368);
nor U7650 (N_7650,N_4448,N_5876);
or U7651 (N_7651,N_5058,N_5642);
xnor U7652 (N_7652,N_5544,N_4193);
nor U7653 (N_7653,N_4614,N_5219);
or U7654 (N_7654,N_4151,N_4200);
or U7655 (N_7655,N_5348,N_4100);
or U7656 (N_7656,N_5103,N_4099);
xor U7657 (N_7657,N_4131,N_5217);
nor U7658 (N_7658,N_5618,N_4926);
or U7659 (N_7659,N_4646,N_5155);
nand U7660 (N_7660,N_4820,N_4297);
xnor U7661 (N_7661,N_4601,N_5767);
xnor U7662 (N_7662,N_4826,N_5350);
and U7663 (N_7663,N_5475,N_4184);
xor U7664 (N_7664,N_5174,N_4758);
and U7665 (N_7665,N_4326,N_4098);
or U7666 (N_7666,N_4036,N_5240);
nor U7667 (N_7667,N_4614,N_4029);
nor U7668 (N_7668,N_4636,N_4185);
nor U7669 (N_7669,N_4233,N_5358);
nor U7670 (N_7670,N_5405,N_4277);
nand U7671 (N_7671,N_4557,N_4181);
or U7672 (N_7672,N_5658,N_4856);
xnor U7673 (N_7673,N_4621,N_4005);
xnor U7674 (N_7674,N_5893,N_4398);
and U7675 (N_7675,N_5978,N_4258);
nor U7676 (N_7676,N_4537,N_4309);
nand U7677 (N_7677,N_4920,N_4955);
nand U7678 (N_7678,N_5302,N_5648);
xnor U7679 (N_7679,N_5338,N_4805);
and U7680 (N_7680,N_5678,N_4844);
or U7681 (N_7681,N_5716,N_5779);
or U7682 (N_7682,N_5601,N_4055);
nand U7683 (N_7683,N_5597,N_5913);
nor U7684 (N_7684,N_5303,N_4315);
or U7685 (N_7685,N_4397,N_4141);
nor U7686 (N_7686,N_4680,N_5933);
or U7687 (N_7687,N_4021,N_5291);
xor U7688 (N_7688,N_5788,N_4008);
nor U7689 (N_7689,N_5533,N_4241);
nand U7690 (N_7690,N_4620,N_5258);
or U7691 (N_7691,N_4082,N_5829);
xnor U7692 (N_7692,N_5925,N_5199);
and U7693 (N_7693,N_5022,N_4211);
and U7694 (N_7694,N_5375,N_4645);
nor U7695 (N_7695,N_5606,N_5623);
nand U7696 (N_7696,N_4353,N_5022);
and U7697 (N_7697,N_5790,N_5362);
nor U7698 (N_7698,N_4407,N_5483);
or U7699 (N_7699,N_5947,N_4992);
or U7700 (N_7700,N_4769,N_5487);
or U7701 (N_7701,N_5970,N_5650);
xor U7702 (N_7702,N_4700,N_4337);
or U7703 (N_7703,N_4292,N_4261);
nor U7704 (N_7704,N_5404,N_4571);
nand U7705 (N_7705,N_5901,N_5763);
or U7706 (N_7706,N_5109,N_5511);
or U7707 (N_7707,N_5561,N_5189);
xnor U7708 (N_7708,N_4663,N_5685);
nor U7709 (N_7709,N_4309,N_5411);
nand U7710 (N_7710,N_5363,N_5617);
and U7711 (N_7711,N_4301,N_4268);
xor U7712 (N_7712,N_4348,N_5418);
or U7713 (N_7713,N_5934,N_4762);
xnor U7714 (N_7714,N_4866,N_5011);
nand U7715 (N_7715,N_5702,N_4855);
xor U7716 (N_7716,N_4902,N_4566);
and U7717 (N_7717,N_4618,N_4413);
xor U7718 (N_7718,N_4036,N_5224);
xnor U7719 (N_7719,N_5171,N_5088);
and U7720 (N_7720,N_4815,N_4669);
and U7721 (N_7721,N_5160,N_4863);
nor U7722 (N_7722,N_5354,N_5469);
xnor U7723 (N_7723,N_5155,N_5708);
nand U7724 (N_7724,N_4000,N_4876);
nor U7725 (N_7725,N_5706,N_5105);
and U7726 (N_7726,N_5746,N_5132);
or U7727 (N_7727,N_4711,N_4152);
and U7728 (N_7728,N_4756,N_4047);
nand U7729 (N_7729,N_5740,N_5406);
xnor U7730 (N_7730,N_4694,N_4278);
xor U7731 (N_7731,N_5049,N_4625);
nand U7732 (N_7732,N_4324,N_4820);
and U7733 (N_7733,N_4291,N_5748);
or U7734 (N_7734,N_5883,N_4309);
or U7735 (N_7735,N_5200,N_4012);
or U7736 (N_7736,N_5628,N_4103);
or U7737 (N_7737,N_4428,N_4197);
nor U7738 (N_7738,N_4677,N_5737);
and U7739 (N_7739,N_5474,N_4192);
nand U7740 (N_7740,N_4761,N_5127);
xor U7741 (N_7741,N_4336,N_4096);
nand U7742 (N_7742,N_4669,N_4905);
nand U7743 (N_7743,N_5354,N_4752);
nand U7744 (N_7744,N_4610,N_4336);
or U7745 (N_7745,N_4318,N_5475);
xor U7746 (N_7746,N_5854,N_4958);
or U7747 (N_7747,N_5246,N_5448);
nand U7748 (N_7748,N_4624,N_4997);
and U7749 (N_7749,N_4062,N_5516);
or U7750 (N_7750,N_4938,N_4599);
nor U7751 (N_7751,N_4549,N_5289);
nand U7752 (N_7752,N_4496,N_4062);
xnor U7753 (N_7753,N_5456,N_4812);
and U7754 (N_7754,N_4642,N_4149);
and U7755 (N_7755,N_5301,N_4977);
and U7756 (N_7756,N_4607,N_4153);
nor U7757 (N_7757,N_5277,N_5949);
xnor U7758 (N_7758,N_4876,N_4472);
or U7759 (N_7759,N_4902,N_5164);
xor U7760 (N_7760,N_4169,N_5948);
or U7761 (N_7761,N_5258,N_5504);
nor U7762 (N_7762,N_5412,N_4406);
and U7763 (N_7763,N_4194,N_4176);
or U7764 (N_7764,N_4553,N_5537);
xor U7765 (N_7765,N_4706,N_4177);
xor U7766 (N_7766,N_5375,N_5956);
nor U7767 (N_7767,N_5588,N_4131);
and U7768 (N_7768,N_5057,N_4404);
nand U7769 (N_7769,N_4965,N_5975);
xnor U7770 (N_7770,N_4808,N_5110);
xnor U7771 (N_7771,N_4627,N_5359);
or U7772 (N_7772,N_5589,N_5439);
nand U7773 (N_7773,N_4984,N_4134);
nor U7774 (N_7774,N_5284,N_5296);
and U7775 (N_7775,N_4308,N_4695);
nand U7776 (N_7776,N_4882,N_4161);
and U7777 (N_7777,N_5918,N_4762);
nand U7778 (N_7778,N_4357,N_5775);
xnor U7779 (N_7779,N_5727,N_5427);
and U7780 (N_7780,N_4595,N_4501);
or U7781 (N_7781,N_4009,N_5034);
nor U7782 (N_7782,N_4957,N_4537);
nand U7783 (N_7783,N_4271,N_4129);
nor U7784 (N_7784,N_5585,N_5744);
and U7785 (N_7785,N_5145,N_5737);
or U7786 (N_7786,N_5889,N_5296);
or U7787 (N_7787,N_4305,N_4539);
or U7788 (N_7788,N_5924,N_4653);
nor U7789 (N_7789,N_4037,N_4693);
xor U7790 (N_7790,N_4018,N_4984);
and U7791 (N_7791,N_4252,N_5167);
nor U7792 (N_7792,N_4028,N_4023);
xor U7793 (N_7793,N_4038,N_4345);
and U7794 (N_7794,N_4778,N_4165);
and U7795 (N_7795,N_5499,N_5294);
nand U7796 (N_7796,N_5345,N_5056);
nor U7797 (N_7797,N_5057,N_5890);
nand U7798 (N_7798,N_4460,N_5291);
or U7799 (N_7799,N_4538,N_4734);
nor U7800 (N_7800,N_5065,N_5512);
xor U7801 (N_7801,N_4527,N_4167);
nor U7802 (N_7802,N_4366,N_4879);
xnor U7803 (N_7803,N_4783,N_5734);
and U7804 (N_7804,N_5717,N_4182);
xnor U7805 (N_7805,N_5941,N_4606);
or U7806 (N_7806,N_4162,N_4977);
and U7807 (N_7807,N_4195,N_5161);
or U7808 (N_7808,N_4148,N_4168);
nand U7809 (N_7809,N_5103,N_4886);
and U7810 (N_7810,N_4396,N_5765);
nand U7811 (N_7811,N_4964,N_5689);
nor U7812 (N_7812,N_4858,N_4352);
nand U7813 (N_7813,N_4374,N_5354);
nand U7814 (N_7814,N_5585,N_5685);
xor U7815 (N_7815,N_4505,N_5118);
nor U7816 (N_7816,N_4002,N_5001);
nor U7817 (N_7817,N_4381,N_5343);
xor U7818 (N_7818,N_5367,N_5633);
and U7819 (N_7819,N_4471,N_5013);
nand U7820 (N_7820,N_4179,N_4238);
nand U7821 (N_7821,N_5036,N_5137);
and U7822 (N_7822,N_5291,N_5616);
nand U7823 (N_7823,N_5847,N_5292);
and U7824 (N_7824,N_5163,N_4071);
nor U7825 (N_7825,N_4865,N_4381);
nor U7826 (N_7826,N_4993,N_4922);
nor U7827 (N_7827,N_4196,N_5317);
and U7828 (N_7828,N_4100,N_5377);
nand U7829 (N_7829,N_4856,N_4311);
or U7830 (N_7830,N_5577,N_5836);
and U7831 (N_7831,N_5439,N_4636);
nand U7832 (N_7832,N_4373,N_4179);
or U7833 (N_7833,N_4207,N_4078);
nand U7834 (N_7834,N_4015,N_5218);
nor U7835 (N_7835,N_5087,N_5404);
xor U7836 (N_7836,N_4716,N_5709);
or U7837 (N_7837,N_4567,N_4341);
xor U7838 (N_7838,N_5150,N_4817);
and U7839 (N_7839,N_5430,N_4592);
nand U7840 (N_7840,N_4733,N_4914);
nor U7841 (N_7841,N_5663,N_4445);
or U7842 (N_7842,N_5320,N_5254);
xnor U7843 (N_7843,N_5321,N_5252);
and U7844 (N_7844,N_5748,N_4331);
nand U7845 (N_7845,N_4871,N_4260);
nor U7846 (N_7846,N_4887,N_4337);
nor U7847 (N_7847,N_5548,N_4699);
or U7848 (N_7848,N_4109,N_5436);
or U7849 (N_7849,N_5582,N_4764);
xor U7850 (N_7850,N_5638,N_4405);
and U7851 (N_7851,N_4872,N_5425);
or U7852 (N_7852,N_5705,N_4856);
and U7853 (N_7853,N_4477,N_4967);
and U7854 (N_7854,N_4142,N_4935);
nor U7855 (N_7855,N_4091,N_5868);
and U7856 (N_7856,N_5805,N_5250);
nor U7857 (N_7857,N_5360,N_5231);
and U7858 (N_7858,N_4259,N_5334);
nor U7859 (N_7859,N_5188,N_5887);
nor U7860 (N_7860,N_4343,N_5588);
or U7861 (N_7861,N_5868,N_4121);
or U7862 (N_7862,N_5723,N_5427);
xor U7863 (N_7863,N_4041,N_4504);
xor U7864 (N_7864,N_5305,N_5517);
nand U7865 (N_7865,N_5556,N_5261);
xnor U7866 (N_7866,N_4955,N_5959);
nand U7867 (N_7867,N_4044,N_4301);
or U7868 (N_7868,N_5709,N_5505);
nand U7869 (N_7869,N_5015,N_4336);
or U7870 (N_7870,N_5778,N_5999);
nand U7871 (N_7871,N_5391,N_5505);
nor U7872 (N_7872,N_4527,N_4064);
xnor U7873 (N_7873,N_5351,N_5003);
nand U7874 (N_7874,N_4662,N_4585);
and U7875 (N_7875,N_5945,N_4728);
and U7876 (N_7876,N_4868,N_5536);
and U7877 (N_7877,N_4440,N_5379);
or U7878 (N_7878,N_4145,N_5904);
or U7879 (N_7879,N_4486,N_5036);
and U7880 (N_7880,N_5915,N_5838);
and U7881 (N_7881,N_4647,N_4626);
nand U7882 (N_7882,N_4221,N_5355);
xnor U7883 (N_7883,N_4927,N_4923);
xor U7884 (N_7884,N_4175,N_4521);
nor U7885 (N_7885,N_5456,N_4599);
nand U7886 (N_7886,N_5397,N_5094);
and U7887 (N_7887,N_4717,N_5516);
or U7888 (N_7888,N_4726,N_4882);
and U7889 (N_7889,N_4162,N_4085);
or U7890 (N_7890,N_5022,N_4203);
or U7891 (N_7891,N_4603,N_5607);
or U7892 (N_7892,N_5143,N_5906);
and U7893 (N_7893,N_5949,N_4352);
nor U7894 (N_7894,N_4167,N_4041);
nand U7895 (N_7895,N_4713,N_5963);
xor U7896 (N_7896,N_4270,N_4195);
nand U7897 (N_7897,N_4375,N_4361);
nand U7898 (N_7898,N_5135,N_5948);
nand U7899 (N_7899,N_4803,N_5905);
and U7900 (N_7900,N_4474,N_4018);
and U7901 (N_7901,N_4383,N_5733);
and U7902 (N_7902,N_5420,N_5880);
or U7903 (N_7903,N_4033,N_5310);
and U7904 (N_7904,N_5017,N_5095);
xnor U7905 (N_7905,N_4984,N_5087);
nand U7906 (N_7906,N_4137,N_4349);
xnor U7907 (N_7907,N_4522,N_5612);
nand U7908 (N_7908,N_5358,N_5748);
or U7909 (N_7909,N_5142,N_4971);
nand U7910 (N_7910,N_4949,N_4409);
nand U7911 (N_7911,N_4550,N_4730);
xnor U7912 (N_7912,N_5128,N_4916);
nand U7913 (N_7913,N_5295,N_5419);
nand U7914 (N_7914,N_5469,N_5332);
or U7915 (N_7915,N_5349,N_4049);
nor U7916 (N_7916,N_4360,N_4584);
and U7917 (N_7917,N_4039,N_5790);
nor U7918 (N_7918,N_4903,N_5882);
xnor U7919 (N_7919,N_4706,N_5084);
nor U7920 (N_7920,N_5209,N_5639);
nand U7921 (N_7921,N_5908,N_5886);
and U7922 (N_7922,N_5566,N_4059);
nor U7923 (N_7923,N_5559,N_4212);
xor U7924 (N_7924,N_4091,N_5470);
and U7925 (N_7925,N_4960,N_4231);
or U7926 (N_7926,N_4124,N_4908);
or U7927 (N_7927,N_4826,N_4863);
or U7928 (N_7928,N_4353,N_5739);
and U7929 (N_7929,N_5643,N_5417);
nand U7930 (N_7930,N_4375,N_4236);
or U7931 (N_7931,N_4485,N_5391);
or U7932 (N_7932,N_4268,N_4620);
xor U7933 (N_7933,N_4244,N_4460);
nor U7934 (N_7934,N_4247,N_5558);
nand U7935 (N_7935,N_4971,N_5590);
nand U7936 (N_7936,N_5307,N_5822);
and U7937 (N_7937,N_4660,N_5807);
and U7938 (N_7938,N_4947,N_4416);
and U7939 (N_7939,N_5167,N_5014);
or U7940 (N_7940,N_4209,N_4677);
nor U7941 (N_7941,N_4766,N_4401);
xor U7942 (N_7942,N_5058,N_5555);
nand U7943 (N_7943,N_4851,N_5211);
nor U7944 (N_7944,N_5030,N_5778);
xnor U7945 (N_7945,N_5425,N_5186);
or U7946 (N_7946,N_4665,N_5260);
nand U7947 (N_7947,N_4966,N_4670);
or U7948 (N_7948,N_4735,N_5665);
or U7949 (N_7949,N_4186,N_4811);
xor U7950 (N_7950,N_5571,N_5342);
nor U7951 (N_7951,N_5340,N_5069);
nand U7952 (N_7952,N_4573,N_4401);
and U7953 (N_7953,N_4975,N_4504);
nor U7954 (N_7954,N_4436,N_5500);
xor U7955 (N_7955,N_5038,N_5843);
nor U7956 (N_7956,N_4862,N_5813);
and U7957 (N_7957,N_4308,N_5656);
and U7958 (N_7958,N_4886,N_4748);
nor U7959 (N_7959,N_4084,N_5105);
nand U7960 (N_7960,N_5145,N_4395);
or U7961 (N_7961,N_4059,N_5267);
xnor U7962 (N_7962,N_4869,N_5890);
nor U7963 (N_7963,N_4824,N_5746);
nor U7964 (N_7964,N_5105,N_4042);
and U7965 (N_7965,N_4650,N_5559);
and U7966 (N_7966,N_5900,N_4957);
xnor U7967 (N_7967,N_5269,N_4038);
nand U7968 (N_7968,N_4893,N_4895);
and U7969 (N_7969,N_4608,N_4845);
and U7970 (N_7970,N_5975,N_5009);
and U7971 (N_7971,N_4194,N_5823);
xnor U7972 (N_7972,N_4828,N_5006);
nor U7973 (N_7973,N_5838,N_5742);
nor U7974 (N_7974,N_5433,N_4266);
xnor U7975 (N_7975,N_5073,N_5004);
xnor U7976 (N_7976,N_4484,N_4193);
xor U7977 (N_7977,N_5287,N_4400);
xor U7978 (N_7978,N_4521,N_4287);
nand U7979 (N_7979,N_5752,N_4888);
xor U7980 (N_7980,N_4503,N_5378);
and U7981 (N_7981,N_4867,N_4248);
or U7982 (N_7982,N_4102,N_5768);
or U7983 (N_7983,N_4022,N_4371);
or U7984 (N_7984,N_5373,N_5855);
xnor U7985 (N_7985,N_4244,N_4042);
and U7986 (N_7986,N_4138,N_5565);
and U7987 (N_7987,N_5560,N_5997);
nand U7988 (N_7988,N_4772,N_5584);
and U7989 (N_7989,N_4494,N_5795);
nor U7990 (N_7990,N_4992,N_5422);
or U7991 (N_7991,N_5749,N_4797);
and U7992 (N_7992,N_5814,N_5651);
nand U7993 (N_7993,N_5634,N_4554);
and U7994 (N_7994,N_5268,N_5789);
nand U7995 (N_7995,N_5066,N_5385);
nand U7996 (N_7996,N_4307,N_5270);
or U7997 (N_7997,N_5521,N_5099);
or U7998 (N_7998,N_4960,N_4689);
and U7999 (N_7999,N_5577,N_4333);
xnor U8000 (N_8000,N_7740,N_6352);
and U8001 (N_8001,N_6271,N_7648);
or U8002 (N_8002,N_6050,N_7510);
or U8003 (N_8003,N_6110,N_7078);
nand U8004 (N_8004,N_7706,N_6964);
or U8005 (N_8005,N_6917,N_7048);
nand U8006 (N_8006,N_7286,N_7214);
xor U8007 (N_8007,N_7958,N_6792);
nand U8008 (N_8008,N_6475,N_6389);
and U8009 (N_8009,N_6859,N_7416);
nand U8010 (N_8010,N_7255,N_6405);
or U8011 (N_8011,N_6032,N_6830);
nand U8012 (N_8012,N_6738,N_7871);
and U8013 (N_8013,N_6321,N_7972);
xnor U8014 (N_8014,N_7542,N_6610);
and U8015 (N_8015,N_6960,N_6320);
or U8016 (N_8016,N_7637,N_7716);
nor U8017 (N_8017,N_7742,N_7237);
and U8018 (N_8018,N_6106,N_6282);
xor U8019 (N_8019,N_7195,N_7913);
nand U8020 (N_8020,N_7628,N_6024);
xor U8021 (N_8021,N_6929,N_7643);
or U8022 (N_8022,N_7312,N_6556);
nor U8023 (N_8023,N_7157,N_6111);
nand U8024 (N_8024,N_7346,N_6460);
xor U8025 (N_8025,N_6971,N_6477);
xor U8026 (N_8026,N_6086,N_7406);
nor U8027 (N_8027,N_7508,N_7095);
or U8028 (N_8028,N_7762,N_7124);
or U8029 (N_8029,N_6848,N_7390);
xnor U8030 (N_8030,N_6711,N_7401);
and U8031 (N_8031,N_6627,N_6347);
and U8032 (N_8032,N_6443,N_6979);
nand U8033 (N_8033,N_7501,N_6870);
nor U8034 (N_8034,N_6723,N_6666);
xor U8035 (N_8035,N_7528,N_6289);
xnor U8036 (N_8036,N_6537,N_7968);
or U8037 (N_8037,N_7348,N_7884);
xor U8038 (N_8038,N_7333,N_6868);
or U8039 (N_8039,N_7307,N_6961);
nand U8040 (N_8040,N_7512,N_6297);
xor U8041 (N_8041,N_7503,N_6363);
and U8042 (N_8042,N_6850,N_6747);
xnor U8043 (N_8043,N_6863,N_7232);
xor U8044 (N_8044,N_7155,N_7571);
or U8045 (N_8045,N_7424,N_6126);
and U8046 (N_8046,N_6878,N_6004);
nand U8047 (N_8047,N_6467,N_6586);
and U8048 (N_8048,N_6327,N_7365);
nand U8049 (N_8049,N_7407,N_6206);
or U8050 (N_8050,N_6055,N_6770);
nor U8051 (N_8051,N_7259,N_6398);
xor U8052 (N_8052,N_6708,N_6171);
and U8053 (N_8053,N_7771,N_6632);
or U8054 (N_8054,N_6031,N_7785);
nor U8055 (N_8055,N_7100,N_7970);
or U8056 (N_8056,N_7960,N_6644);
nand U8057 (N_8057,N_6757,N_7544);
or U8058 (N_8058,N_7736,N_7163);
or U8059 (N_8059,N_7376,N_7747);
nand U8060 (N_8060,N_7351,N_7246);
nor U8061 (N_8061,N_6845,N_7844);
nand U8062 (N_8062,N_7437,N_7493);
nor U8063 (N_8063,N_6115,N_7897);
nand U8064 (N_8064,N_7760,N_7241);
and U8065 (N_8065,N_6535,N_7971);
or U8066 (N_8066,N_7654,N_6502);
and U8067 (N_8067,N_6232,N_7103);
nor U8068 (N_8068,N_6240,N_7277);
nor U8069 (N_8069,N_6052,N_7197);
nand U8070 (N_8070,N_6790,N_7222);
or U8071 (N_8071,N_7064,N_6325);
xor U8072 (N_8072,N_7506,N_6874);
and U8073 (N_8073,N_6436,N_6296);
xnor U8074 (N_8074,N_7854,N_7610);
and U8075 (N_8075,N_7561,N_7011);
xnor U8076 (N_8076,N_7344,N_7082);
and U8077 (N_8077,N_6680,N_6408);
or U8078 (N_8078,N_6020,N_7946);
or U8079 (N_8079,N_6500,N_7725);
nor U8080 (N_8080,N_7577,N_6761);
nand U8081 (N_8081,N_6508,N_7388);
nand U8082 (N_8082,N_7253,N_6675);
xor U8083 (N_8083,N_6784,N_6943);
nand U8084 (N_8084,N_7692,N_6259);
and U8085 (N_8085,N_6479,N_7696);
and U8086 (N_8086,N_7768,N_6862);
or U8087 (N_8087,N_7172,N_7961);
nand U8088 (N_8088,N_6151,N_7670);
nor U8089 (N_8089,N_6950,N_6821);
nand U8090 (N_8090,N_6470,N_6759);
nor U8091 (N_8091,N_7459,N_6065);
xor U8092 (N_8092,N_6310,N_6753);
and U8093 (N_8093,N_7184,N_7447);
nand U8094 (N_8094,N_7896,N_7888);
nand U8095 (N_8095,N_6957,N_6384);
and U8096 (N_8096,N_6989,N_6194);
nor U8097 (N_8097,N_7051,N_6141);
xnor U8098 (N_8098,N_7220,N_7339);
nand U8099 (N_8099,N_7022,N_6841);
nand U8100 (N_8100,N_6308,N_6605);
nor U8101 (N_8101,N_7759,N_7835);
nor U8102 (N_8102,N_7616,N_7474);
nor U8103 (N_8103,N_7243,N_7038);
and U8104 (N_8104,N_7533,N_6112);
nor U8105 (N_8105,N_7426,N_6887);
xor U8106 (N_8106,N_7781,N_6737);
and U8107 (N_8107,N_7594,N_7532);
and U8108 (N_8108,N_6923,N_7429);
nand U8109 (N_8109,N_6563,N_6026);
nand U8110 (N_8110,N_7353,N_7583);
and U8111 (N_8111,N_7994,N_6358);
and U8112 (N_8112,N_7983,N_7120);
or U8113 (N_8113,N_7012,N_6455);
nor U8114 (N_8114,N_7289,N_7721);
xor U8115 (N_8115,N_6699,N_6542);
nor U8116 (N_8116,N_7701,N_7436);
and U8117 (N_8117,N_6499,N_6814);
nor U8118 (N_8118,N_6498,N_6655);
nand U8119 (N_8119,N_6799,N_6402);
and U8120 (N_8120,N_6865,N_7359);
nor U8121 (N_8121,N_7470,N_7797);
nand U8122 (N_8122,N_6385,N_6672);
nor U8123 (N_8123,N_6671,N_7130);
xnor U8124 (N_8124,N_6169,N_6785);
xor U8125 (N_8125,N_7402,N_6158);
xnor U8126 (N_8126,N_6999,N_7977);
xor U8127 (N_8127,N_6349,N_7749);
nand U8128 (N_8128,N_7223,N_7743);
and U8129 (N_8129,N_7770,N_6013);
nand U8130 (N_8130,N_7644,N_7445);
and U8131 (N_8131,N_7154,N_6987);
nand U8132 (N_8132,N_7591,N_6447);
and U8133 (N_8133,N_6184,N_6825);
nor U8134 (N_8134,N_7182,N_6375);
xor U8135 (N_8135,N_6290,N_6202);
or U8136 (N_8136,N_7438,N_7336);
nand U8137 (N_8137,N_6210,N_7595);
nand U8138 (N_8138,N_7341,N_6886);
and U8139 (N_8139,N_6018,N_7240);
and U8140 (N_8140,N_6278,N_6426);
nor U8141 (N_8141,N_7627,N_7687);
nor U8142 (N_8142,N_7020,N_7855);
nor U8143 (N_8143,N_7774,N_6397);
and U8144 (N_8144,N_6133,N_7794);
or U8145 (N_8145,N_7008,N_7966);
xnor U8146 (N_8146,N_7384,N_7442);
xnor U8147 (N_8147,N_6913,N_7722);
xor U8148 (N_8148,N_7802,N_7865);
nand U8149 (N_8149,N_6485,N_7773);
or U8150 (N_8150,N_7305,N_7181);
nor U8151 (N_8151,N_7763,N_6474);
and U8152 (N_8152,N_6764,N_7929);
nand U8153 (N_8153,N_6557,N_6372);
and U8154 (N_8154,N_7803,N_6947);
nand U8155 (N_8155,N_6403,N_6687);
nor U8156 (N_8156,N_6673,N_6459);
nand U8157 (N_8157,N_6142,N_7735);
and U8158 (N_8158,N_6645,N_6953);
and U8159 (N_8159,N_7073,N_6554);
and U8160 (N_8160,N_6619,N_7449);
or U8161 (N_8161,N_6730,N_6382);
or U8162 (N_8162,N_6073,N_7058);
xnor U8163 (N_8163,N_6251,N_7114);
nor U8164 (N_8164,N_7981,N_7631);
and U8165 (N_8165,N_7717,N_7988);
nor U8166 (N_8166,N_7828,N_6506);
nand U8167 (N_8167,N_6057,N_6201);
nor U8168 (N_8168,N_6659,N_7371);
nand U8169 (N_8169,N_7541,N_6734);
nor U8170 (N_8170,N_7748,N_7582);
and U8171 (N_8171,N_7822,N_6951);
or U8172 (N_8172,N_6736,N_6551);
nor U8173 (N_8173,N_7604,N_6583);
nor U8174 (N_8174,N_7974,N_6488);
nor U8175 (N_8175,N_6762,N_7420);
nand U8176 (N_8176,N_6279,N_6016);
or U8177 (N_8177,N_6955,N_6660);
or U8178 (N_8178,N_6587,N_7059);
xnor U8179 (N_8179,N_6524,N_7366);
or U8180 (N_8180,N_6180,N_6882);
xor U8181 (N_8181,N_7584,N_6079);
and U8182 (N_8182,N_7909,N_6203);
nand U8183 (N_8183,N_7187,N_6003);
or U8184 (N_8184,N_7985,N_7554);
xor U8185 (N_8185,N_7505,N_7302);
nor U8186 (N_8186,N_6027,N_6724);
xnor U8187 (N_8187,N_6684,N_6341);
nor U8188 (N_8188,N_7036,N_6530);
nor U8189 (N_8189,N_6714,N_6435);
xnor U8190 (N_8190,N_7391,N_7309);
nand U8191 (N_8191,N_6264,N_6433);
nand U8192 (N_8192,N_7709,N_7301);
nand U8193 (N_8193,N_7826,N_7964);
or U8194 (N_8194,N_6849,N_7373);
xnor U8195 (N_8195,N_6776,N_7818);
nor U8196 (N_8196,N_7870,N_7024);
xor U8197 (N_8197,N_6803,N_6513);
and U8198 (N_8198,N_6649,N_7236);
nand U8199 (N_8199,N_7492,N_6829);
nand U8200 (N_8200,N_6975,N_6316);
nand U8201 (N_8201,N_6442,N_7546);
xnor U8202 (N_8202,N_6466,N_7500);
nor U8203 (N_8203,N_7832,N_7094);
xnor U8204 (N_8204,N_7882,N_7144);
or U8205 (N_8205,N_7112,N_7230);
xor U8206 (N_8206,N_6471,N_7685);
nand U8207 (N_8207,N_7601,N_7110);
and U8208 (N_8208,N_7694,N_6005);
nor U8209 (N_8209,N_6454,N_7142);
nand U8210 (N_8210,N_7663,N_6159);
and U8211 (N_8211,N_7469,N_7495);
nor U8212 (N_8212,N_7667,N_6797);
nor U8213 (N_8213,N_7535,N_7620);
xnor U8214 (N_8214,N_6072,N_7317);
nor U8215 (N_8215,N_7250,N_7349);
and U8216 (N_8216,N_6992,N_7991);
nor U8217 (N_8217,N_6033,N_7521);
nor U8218 (N_8218,N_7488,N_6120);
xnor U8219 (N_8219,N_7937,N_7887);
and U8220 (N_8220,N_7191,N_7903);
nor U8221 (N_8221,N_7940,N_7810);
nor U8222 (N_8222,N_7816,N_6885);
or U8223 (N_8223,N_7815,N_6766);
or U8224 (N_8224,N_7350,N_7096);
nor U8225 (N_8225,N_6553,N_6162);
nand U8226 (N_8226,N_7238,N_6407);
nand U8227 (N_8227,N_7283,N_6892);
and U8228 (N_8228,N_7446,N_7821);
xor U8229 (N_8229,N_6096,N_7545);
nand U8230 (N_8230,N_6225,N_6128);
nor U8231 (N_8231,N_6369,N_7558);
xor U8232 (N_8232,N_7877,N_6928);
or U8233 (N_8233,N_7476,N_6547);
and U8234 (N_8234,N_7607,N_7872);
and U8235 (N_8235,N_6360,N_6959);
nor U8236 (N_8236,N_6620,N_7889);
nor U8237 (N_8237,N_7379,N_6107);
xor U8238 (N_8238,N_6097,N_7672);
xor U8239 (N_8239,N_7265,N_6365);
nor U8240 (N_8240,N_7261,N_6323);
nand U8241 (N_8241,N_6175,N_7829);
and U8242 (N_8242,N_7761,N_6525);
xor U8243 (N_8243,N_7710,N_7704);
nor U8244 (N_8244,N_6836,N_7150);
and U8245 (N_8245,N_7143,N_7751);
xor U8246 (N_8246,N_6438,N_7173);
xnor U8247 (N_8247,N_7868,N_7450);
or U8248 (N_8248,N_6905,N_7915);
nor U8249 (N_8249,N_6326,N_6574);
or U8250 (N_8250,N_6359,N_7820);
nor U8251 (N_8251,N_7664,N_6200);
or U8252 (N_8252,N_7718,N_6920);
and U8253 (N_8253,N_7389,N_6420);
xor U8254 (N_8254,N_7262,N_6896);
nand U8255 (N_8255,N_7080,N_6064);
nor U8256 (N_8256,N_7603,N_7953);
or U8257 (N_8257,N_7473,N_7562);
nor U8258 (N_8258,N_6085,N_6504);
nor U8259 (N_8259,N_6116,N_6395);
nand U8260 (N_8260,N_7592,N_7586);
nand U8261 (N_8261,N_6108,N_7196);
and U8262 (N_8262,N_6639,N_7380);
xnor U8263 (N_8263,N_7395,N_7726);
and U8264 (N_8264,N_6676,N_6795);
xor U8265 (N_8265,N_6516,N_7757);
and U8266 (N_8266,N_7817,N_6897);
xnor U8267 (N_8267,N_6001,N_6678);
xor U8268 (N_8268,N_6510,N_6457);
xnor U8269 (N_8269,N_6994,N_6253);
nand U8270 (N_8270,N_7779,N_6315);
or U8271 (N_8271,N_6722,N_6067);
and U8272 (N_8272,N_7671,N_7529);
and U8273 (N_8273,N_7254,N_6414);
nor U8274 (N_8274,N_6854,N_7444);
nand U8275 (N_8275,N_6130,N_6851);
and U8276 (N_8276,N_6099,N_7606);
nand U8277 (N_8277,N_7568,N_7626);
and U8278 (N_8278,N_7923,N_6152);
and U8279 (N_8279,N_7408,N_6198);
nand U8280 (N_8280,N_7860,N_6332);
nor U8281 (N_8281,N_7753,N_6230);
or U8282 (N_8282,N_7634,N_7484);
xnor U8283 (N_8283,N_6331,N_6589);
xnor U8284 (N_8284,N_7224,N_7908);
and U8285 (N_8285,N_7543,N_7364);
xor U8286 (N_8286,N_7853,N_6842);
or U8287 (N_8287,N_6793,N_7400);
nand U8288 (N_8288,N_6534,N_7252);
and U8289 (N_8289,N_7686,N_7233);
or U8290 (N_8290,N_6658,N_7976);
xor U8291 (N_8291,N_7314,N_6638);
or U8292 (N_8292,N_7405,N_6935);
or U8293 (N_8293,N_7192,N_7126);
nor U8294 (N_8294,N_7840,N_7665);
nor U8295 (N_8295,N_7830,N_6280);
and U8296 (N_8296,N_7920,N_6137);
or U8297 (N_8297,N_7471,N_6294);
and U8298 (N_8298,N_7662,N_7030);
nor U8299 (N_8299,N_6756,N_7153);
xnor U8300 (N_8300,N_7332,N_6239);
or U8301 (N_8301,N_6117,N_7814);
nand U8302 (N_8302,N_6394,N_6755);
or U8303 (N_8303,N_6520,N_7356);
nor U8304 (N_8304,N_6195,N_6374);
and U8305 (N_8305,N_6741,N_7813);
nor U8306 (N_8306,N_6453,N_6937);
xnor U8307 (N_8307,N_6906,N_7969);
nor U8308 (N_8308,N_6314,N_6689);
nand U8309 (N_8309,N_6324,N_7042);
nand U8310 (N_8310,N_7691,N_6211);
xor U8311 (N_8311,N_6787,N_6575);
xor U8312 (N_8312,N_7750,N_7002);
nor U8313 (N_8313,N_6875,N_6135);
or U8314 (N_8314,N_6894,N_7919);
or U8315 (N_8315,N_7018,N_7019);
and U8316 (N_8316,N_7918,N_7394);
xor U8317 (N_8317,N_7699,N_7481);
or U8318 (N_8318,N_6009,N_6266);
or U8319 (N_8319,N_6468,N_6462);
and U8320 (N_8320,N_7282,N_6765);
nand U8321 (N_8321,N_7147,N_7180);
and U8322 (N_8322,N_6100,N_6691);
xnor U8323 (N_8323,N_7303,N_7202);
or U8324 (N_8324,N_6172,N_6679);
nand U8325 (N_8325,N_6725,N_7737);
or U8326 (N_8326,N_7891,N_6512);
nand U8327 (N_8327,N_7905,N_7319);
nand U8328 (N_8328,N_7652,N_6348);
nand U8329 (N_8329,N_7066,N_6908);
and U8330 (N_8330,N_7386,N_6340);
xor U8331 (N_8331,N_6933,N_6188);
xor U8332 (N_8332,N_6091,N_7403);
and U8333 (N_8333,N_6503,N_7827);
or U8334 (N_8334,N_6484,N_7653);
nor U8335 (N_8335,N_6731,N_7331);
nor U8336 (N_8336,N_6643,N_6872);
nor U8337 (N_8337,N_6631,N_7496);
nand U8338 (N_8338,N_6548,N_6647);
or U8339 (N_8339,N_6307,N_7987);
nand U8340 (N_8340,N_7839,N_7858);
nor U8341 (N_8341,N_7183,N_7084);
xnor U8342 (N_8342,N_6599,N_6998);
nand U8343 (N_8343,N_7873,N_7363);
nor U8344 (N_8344,N_6312,N_7378);
nand U8345 (N_8345,N_6518,N_7724);
xnor U8346 (N_8346,N_6584,N_7057);
or U8347 (N_8347,N_6606,N_7178);
or U8348 (N_8348,N_6342,N_7475);
nand U8349 (N_8349,N_6921,N_7498);
nand U8350 (N_8350,N_7169,N_6925);
or U8351 (N_8351,N_7907,N_6489);
xor U8352 (N_8352,N_6982,N_6411);
or U8353 (N_8353,N_7419,N_6607);
nor U8354 (N_8354,N_6629,N_6010);
and U8355 (N_8355,N_7553,N_6160);
nor U8356 (N_8356,N_7306,N_7605);
or U8357 (N_8357,N_6428,N_7863);
nand U8358 (N_8358,N_6061,N_6059);
nand U8359 (N_8359,N_7451,N_7825);
xor U8360 (N_8360,N_6977,N_6995);
nand U8361 (N_8361,N_6451,N_7000);
and U8362 (N_8362,N_7808,N_6573);
or U8363 (N_8363,N_6161,N_6648);
nor U8364 (N_8364,N_6060,N_6427);
nor U8365 (N_8365,N_6749,N_6336);
or U8366 (N_8366,N_7198,N_7372);
or U8367 (N_8367,N_6751,N_6809);
nor U8368 (N_8368,N_6746,N_6881);
nor U8369 (N_8369,N_7354,N_7101);
and U8370 (N_8370,N_7478,N_7249);
nand U8371 (N_8371,N_7128,N_6011);
or U8372 (N_8372,N_6155,N_6798);
nor U8373 (N_8373,N_7792,N_6245);
and U8374 (N_8374,N_6772,N_6740);
nand U8375 (N_8375,N_6274,N_6864);
nand U8376 (N_8376,N_6909,N_6227);
nand U8377 (N_8377,N_6568,N_7515);
and U8378 (N_8378,N_6527,N_7675);
xnor U8379 (N_8379,N_6805,N_6378);
nor U8380 (N_8380,N_7567,N_6983);
and U8381 (N_8381,N_6248,N_7795);
xnor U8382 (N_8382,N_7279,N_6140);
nor U8383 (N_8383,N_7487,N_6663);
nor U8384 (N_8384,N_6536,N_7092);
xor U8385 (N_8385,N_6837,N_6727);
and U8386 (N_8386,N_7219,N_7458);
nand U8387 (N_8387,N_7911,N_7931);
or U8388 (N_8388,N_7593,N_7764);
nand U8389 (N_8389,N_7581,N_7275);
nor U8390 (N_8390,N_7382,N_7656);
nand U8391 (N_8391,N_7945,N_7185);
nand U8392 (N_8392,N_6424,N_7215);
and U8393 (N_8393,N_6828,N_7035);
and U8394 (N_8394,N_7936,N_7732);
nor U8395 (N_8395,N_7479,N_7801);
nand U8396 (N_8396,N_7557,N_7385);
and U8397 (N_8397,N_7875,N_6368);
xor U8398 (N_8398,N_6039,N_6063);
nand U8399 (N_8399,N_6721,N_6415);
nand U8400 (N_8400,N_6818,N_7170);
and U8401 (N_8401,N_6856,N_6241);
or U8402 (N_8402,N_7922,N_6540);
nor U8403 (N_8403,N_7646,N_7878);
and U8404 (N_8404,N_6208,N_6807);
nand U8405 (N_8405,N_7097,N_7069);
nor U8406 (N_8406,N_7127,N_6042);
xnor U8407 (N_8407,N_6739,N_7811);
or U8408 (N_8408,N_6523,N_6123);
or U8409 (N_8409,N_6509,N_7697);
or U8410 (N_8410,N_7149,N_7746);
or U8411 (N_8411,N_7315,N_6700);
nand U8412 (N_8412,N_7428,N_7037);
nand U8413 (N_8413,N_6430,N_7580);
nand U8414 (N_8414,N_7688,N_7893);
and U8415 (N_8415,N_7158,N_6356);
nand U8416 (N_8416,N_7962,N_7461);
xnor U8417 (N_8417,N_6019,N_7235);
or U8418 (N_8418,N_6002,N_7910);
and U8419 (N_8419,N_7398,N_6329);
and U8420 (N_8420,N_7338,N_7116);
nand U8421 (N_8421,N_6150,N_6339);
xor U8422 (N_8422,N_6613,N_6461);
nor U8423 (N_8423,N_6616,N_6493);
or U8424 (N_8424,N_7041,N_7951);
or U8425 (N_8425,N_6726,N_6800);
and U8426 (N_8426,N_7006,N_7269);
nor U8427 (N_8427,N_6284,N_6577);
nand U8428 (N_8428,N_7993,N_7098);
nor U8429 (N_8429,N_7745,N_6432);
or U8430 (N_8430,N_7015,N_7793);
and U8431 (N_8431,N_6177,N_6665);
nand U8432 (N_8432,N_7530,N_6936);
xnor U8433 (N_8433,N_6838,N_7523);
nor U8434 (N_8434,N_7714,N_7619);
and U8435 (N_8435,N_6735,N_6446);
nor U8436 (N_8436,N_6246,N_7174);
or U8437 (N_8437,N_6233,N_7355);
and U8438 (N_8438,N_6379,N_7713);
and U8439 (N_8439,N_6907,N_6924);
nor U8440 (N_8440,N_6263,N_7085);
or U8441 (N_8441,N_6634,N_6662);
xnor U8442 (N_8442,N_6434,N_7052);
or U8443 (N_8443,N_7293,N_6565);
and U8444 (N_8444,N_7838,N_7809);
xnor U8445 (N_8445,N_6552,N_7071);
nor U8446 (N_8446,N_7491,N_6601);
nand U8447 (N_8447,N_6945,N_6852);
and U8448 (N_8448,N_7831,N_7517);
and U8449 (N_8449,N_7739,N_7590);
xnor U8450 (N_8450,N_7404,N_6322);
nor U8451 (N_8451,N_7899,N_6891);
xnor U8452 (N_8452,N_6113,N_6058);
nand U8453 (N_8453,N_6633,N_6831);
and U8454 (N_8454,N_7062,N_6694);
nand U8455 (N_8455,N_6173,N_7520);
nor U8456 (N_8456,N_6304,N_6603);
nor U8457 (N_8457,N_6581,N_7755);
or U8458 (N_8458,N_6636,N_6223);
nor U8459 (N_8459,N_6667,N_6265);
xnor U8460 (N_8460,N_6781,N_6683);
nand U8461 (N_8461,N_7531,N_6078);
nor U8462 (N_8462,N_6733,N_7957);
and U8463 (N_8463,N_6533,N_6546);
nand U8464 (N_8464,N_6301,N_6926);
nand U8465 (N_8465,N_6715,N_7703);
nor U8466 (N_8466,N_6853,N_7635);
or U8467 (N_8467,N_7477,N_6914);
nor U8468 (N_8468,N_7859,N_6791);
and U8469 (N_8469,N_6915,N_6939);
and U8470 (N_8470,N_6710,N_6650);
xor U8471 (N_8471,N_7556,N_7145);
nand U8472 (N_8472,N_7565,N_7466);
xnor U8473 (N_8473,N_6495,N_7707);
nand U8474 (N_8474,N_6070,N_6661);
and U8475 (N_8475,N_7924,N_6048);
or U8476 (N_8476,N_6823,N_7621);
xnor U8477 (N_8477,N_7290,N_7758);
nand U8478 (N_8478,N_6769,N_7190);
xnor U8479 (N_8479,N_7399,N_6835);
nor U8480 (N_8480,N_6732,N_6306);
or U8481 (N_8481,N_6178,N_7370);
and U8482 (N_8482,N_6092,N_6147);
and U8483 (N_8483,N_7211,N_7454);
and U8484 (N_8484,N_7998,N_6229);
and U8485 (N_8485,N_7847,N_7087);
or U8486 (N_8486,N_7851,N_6285);
xnor U8487 (N_8487,N_7693,N_6614);
nor U8488 (N_8488,N_6529,N_6025);
or U8489 (N_8489,N_6558,N_6387);
and U8490 (N_8490,N_7368,N_6640);
nand U8491 (N_8491,N_6651,N_6932);
and U8492 (N_8492,N_6981,N_6624);
nor U8493 (N_8493,N_7549,N_7787);
xnor U8494 (N_8494,N_6228,N_6934);
nand U8495 (N_8495,N_7677,N_6621);
nor U8496 (N_8496,N_7700,N_6305);
xor U8497 (N_8497,N_7415,N_6090);
and U8498 (N_8498,N_6431,N_6441);
nand U8499 (N_8499,N_6812,N_6539);
and U8500 (N_8500,N_7330,N_7141);
nor U8501 (N_8501,N_7719,N_7723);
nand U8502 (N_8502,N_7752,N_6641);
or U8503 (N_8503,N_7658,N_6164);
or U8504 (N_8504,N_7999,N_7090);
or U8505 (N_8505,N_7979,N_7106);
nor U8506 (N_8506,N_6094,N_6617);
or U8507 (N_8507,N_6393,N_7228);
or U8508 (N_8508,N_6890,N_7016);
nand U8509 (N_8509,N_7705,N_6464);
nand U8510 (N_8510,N_6388,N_7266);
or U8511 (N_8511,N_7956,N_6416);
nor U8512 (N_8512,N_6879,N_7025);
or U8513 (N_8513,N_7698,N_6993);
nand U8514 (N_8514,N_7291,N_6144);
and U8515 (N_8515,N_6867,N_7189);
nand U8516 (N_8516,N_6952,N_6528);
nand U8517 (N_8517,N_7866,N_7845);
nor U8518 (N_8518,N_7932,N_7633);
and U8519 (N_8519,N_7421,N_6973);
or U8520 (N_8520,N_7328,N_7433);
nor U8521 (N_8521,N_6703,N_6463);
nor U8522 (N_8522,N_7796,N_6292);
or U8523 (N_8523,N_6390,N_7849);
nor U8524 (N_8524,N_6138,N_6802);
and U8525 (N_8525,N_7525,N_7930);
or U8526 (N_8526,N_6077,N_6256);
or U8527 (N_8527,N_6082,N_6129);
nor U8528 (N_8528,N_7712,N_6709);
and U8529 (N_8529,N_7857,N_7263);
nor U8530 (N_8530,N_7782,N_6317);
or U8531 (N_8531,N_7507,N_6986);
nor U8532 (N_8532,N_6866,N_7137);
nand U8533 (N_8533,N_6743,N_6948);
or U8534 (N_8534,N_6777,N_6779);
or U8535 (N_8535,N_7618,N_7131);
and U8536 (N_8536,N_7093,N_7852);
nor U8537 (N_8537,N_6215,N_7369);
or U8538 (N_8538,N_7744,N_7200);
nor U8539 (N_8539,N_7435,N_6801);
xnor U8540 (N_8540,N_7367,N_7362);
nor U8541 (N_8541,N_6399,N_6693);
nor U8542 (N_8542,N_7898,N_6148);
nand U8543 (N_8543,N_7014,N_6084);
nor U8544 (N_8544,N_6889,N_6839);
xnor U8545 (N_8545,N_7702,N_6071);
nor U8546 (N_8546,N_6771,N_7115);
xnor U8547 (N_8547,N_6521,N_7798);
nor U8548 (N_8548,N_7657,N_7996);
and U8549 (N_8549,N_7902,N_7602);
or U8550 (N_8550,N_7452,N_7916);
xor U8551 (N_8551,N_7661,N_7609);
nor U8552 (N_8552,N_6083,N_7334);
xor U8553 (N_8553,N_6205,N_7926);
nor U8554 (N_8554,N_7159,N_7357);
and U8555 (N_8555,N_7070,N_7026);
nand U8556 (N_8556,N_6105,N_7728);
and U8557 (N_8557,N_6181,N_7343);
nor U8558 (N_8558,N_7846,N_7617);
xor U8559 (N_8559,N_7140,N_7519);
or U8560 (N_8560,N_6602,N_7807);
xnor U8561 (N_8561,N_7050,N_7273);
xor U8562 (N_8562,N_6718,N_6218);
and U8563 (N_8563,N_6361,N_6486);
nand U8564 (N_8564,N_6623,N_7848);
and U8565 (N_8565,N_6043,N_6775);
xnor U8566 (N_8566,N_7463,N_7177);
nand U8567 (N_8567,N_6409,N_6517);
nor U8568 (N_8568,N_6255,N_7088);
nor U8569 (N_8569,N_7598,N_6444);
or U8570 (N_8570,N_7392,N_6910);
nand U8571 (N_8571,N_7612,N_7731);
xnor U8572 (N_8572,N_7374,N_7324);
and U8573 (N_8573,N_6187,N_6247);
nand U8574 (N_8574,N_6046,N_7053);
nand U8575 (N_8575,N_6417,N_6783);
nor U8576 (N_8576,N_6422,N_7624);
xnor U8577 (N_8577,N_7242,N_7063);
xnor U8578 (N_8578,N_7280,N_6491);
and U8579 (N_8579,N_6174,N_6822);
nor U8580 (N_8580,N_7417,N_7431);
xnor U8581 (N_8581,N_6668,N_6592);
and U8582 (N_8582,N_6258,N_7711);
nor U8583 (N_8583,N_7780,N_7292);
and U8584 (N_8584,N_7199,N_6847);
nor U8585 (N_8585,N_6635,N_7494);
xor U8586 (N_8586,N_6189,N_6963);
xor U8587 (N_8587,N_7944,N_6139);
xnor U8588 (N_8588,N_7342,N_6656);
nor U8589 (N_8589,N_6037,N_6237);
nor U8590 (N_8590,N_7669,N_6418);
nor U8591 (N_8591,N_6600,N_6269);
and U8592 (N_8592,N_6238,N_6996);
nor U8593 (N_8593,N_7720,N_7497);
xnor U8594 (N_8594,N_7335,N_7117);
nor U8595 (N_8595,N_7683,N_6114);
xnor U8596 (N_8596,N_7203,N_7049);
or U8597 (N_8597,N_7276,N_6482);
xor U8598 (N_8598,N_7133,N_7917);
and U8599 (N_8599,N_7287,N_7432);
nor U8600 (N_8600,N_7514,N_6819);
and U8601 (N_8601,N_6012,N_7695);
and U8602 (N_8602,N_6125,N_7666);
nor U8603 (N_8603,N_6705,N_7004);
or U8604 (N_8604,N_6334,N_7105);
nor U8605 (N_8605,N_6901,N_7067);
nor U8606 (N_8606,N_7194,N_7833);
nor U8607 (N_8607,N_7056,N_7457);
nand U8608 (N_8608,N_7756,N_6413);
and U8609 (N_8609,N_7322,N_6978);
nor U8610 (N_8610,N_6226,N_7730);
nand U8611 (N_8611,N_6191,N_6811);
nor U8612 (N_8612,N_6054,N_7842);
nor U8613 (N_8613,N_7448,N_7358);
and U8614 (N_8614,N_6944,N_6681);
or U8615 (N_8615,N_7864,N_7193);
or U8616 (N_8616,N_6806,N_6450);
xor U8617 (N_8617,N_6904,N_7104);
and U8618 (N_8618,N_6653,N_6146);
or U8619 (N_8619,N_7651,N_6492);
xor U8620 (N_8620,N_7805,N_7485);
nor U8621 (N_8621,N_6044,N_7861);
or U8622 (N_8622,N_7572,N_7823);
or U8623 (N_8623,N_7212,N_6871);
nor U8624 (N_8624,N_7927,N_7630);
nand U8625 (N_8625,N_6121,N_6873);
and U8626 (N_8626,N_6350,N_7099);
or U8627 (N_8627,N_7947,N_6118);
xnor U8628 (N_8628,N_7086,N_7352);
nor U8629 (N_8629,N_6927,N_7862);
nand U8630 (N_8630,N_7260,N_7361);
nor U8631 (N_8631,N_7921,N_6391);
and U8632 (N_8632,N_7285,N_6222);
nor U8633 (N_8633,N_7272,N_6938);
xnor U8634 (N_8634,N_6804,N_7121);
and U8635 (N_8635,N_7513,N_7791);
and U8636 (N_8636,N_7122,N_6337);
nand U8637 (N_8637,N_7281,N_6355);
and U8638 (N_8638,N_7423,N_6036);
or U8639 (N_8639,N_7576,N_7892);
or U8640 (N_8640,N_6041,N_7005);
or U8641 (N_8641,N_7638,N_7480);
nor U8642 (N_8642,N_7679,N_7347);
nand U8643 (N_8643,N_6021,N_7650);
nand U8644 (N_8644,N_7992,N_6931);
nand U8645 (N_8645,N_6367,N_7534);
xor U8646 (N_8646,N_6028,N_6490);
xnor U8647 (N_8647,N_7589,N_7790);
or U8648 (N_8648,N_7869,N_7856);
nand U8649 (N_8649,N_7271,N_6089);
or U8650 (N_8650,N_6930,N_6224);
and U8651 (N_8651,N_6465,N_6918);
or U8652 (N_8652,N_6344,N_7234);
nand U8653 (N_8653,N_6754,N_6040);
and U8654 (N_8654,N_7453,N_7055);
and U8655 (N_8655,N_6131,N_7337);
nor U8656 (N_8656,N_6949,N_6682);
xor U8657 (N_8657,N_6750,N_6940);
xor U8658 (N_8658,N_6768,N_7566);
nor U8659 (N_8659,N_7152,N_7901);
and U8660 (N_8660,N_6748,N_6127);
nor U8661 (N_8661,N_7984,N_7570);
nor U8662 (N_8662,N_7550,N_6550);
xnor U8663 (N_8663,N_6439,N_6701);
and U8664 (N_8664,N_7188,N_6782);
xor U8665 (N_8665,N_6778,N_6965);
nor U8666 (N_8666,N_7778,N_6309);
and U8667 (N_8667,N_6015,N_6351);
xnor U8668 (N_8668,N_6007,N_6899);
and U8669 (N_8669,N_7660,N_6883);
or U8670 (N_8670,N_6302,N_6216);
nand U8671 (N_8671,N_6313,N_7054);
nor U8672 (N_8672,N_7935,N_6345);
nand U8673 (N_8673,N_6287,N_6445);
and U8674 (N_8674,N_7614,N_7880);
xor U8675 (N_8675,N_6448,N_6810);
xnor U8676 (N_8676,N_7486,N_6585);
and U8677 (N_8677,N_6697,N_7850);
nand U8678 (N_8678,N_6591,N_6192);
or U8679 (N_8679,N_6834,N_7949);
xnor U8680 (N_8680,N_7075,N_7995);
xor U8681 (N_8681,N_7033,N_7772);
nor U8682 (N_8682,N_7540,N_6531);
xnor U8683 (N_8683,N_6252,N_6532);
or U8684 (N_8684,N_6242,N_6075);
nand U8685 (N_8685,N_7229,N_6145);
or U8686 (N_8686,N_6991,N_7765);
or U8687 (N_8687,N_6622,N_6149);
nand U8688 (N_8688,N_7575,N_7555);
xnor U8689 (N_8689,N_7608,N_7060);
or U8690 (N_8690,N_7874,N_7323);
xor U8691 (N_8691,N_7548,N_6990);
nor U8692 (N_8692,N_7629,N_7539);
xor U8693 (N_8693,N_6234,N_6354);
nand U8694 (N_8694,N_6877,N_6707);
nand U8695 (N_8695,N_7107,N_7091);
nand U8696 (N_8696,N_7411,N_7490);
or U8697 (N_8697,N_6642,N_7257);
nand U8698 (N_8698,N_6396,N_7560);
xnor U8699 (N_8699,N_6832,N_6400);
xnor U8700 (N_8700,N_7166,N_7296);
or U8701 (N_8701,N_7834,N_7216);
nor U8702 (N_8702,N_6576,N_6386);
nor U8703 (N_8703,N_6056,N_6199);
or U8704 (N_8704,N_6880,N_6410);
or U8705 (N_8705,N_7270,N_6712);
xnor U8706 (N_8706,N_7640,N_6646);
or U8707 (N_8707,N_7034,N_6157);
and U8708 (N_8708,N_7786,N_6022);
xor U8709 (N_8709,N_6596,N_7221);
or U8710 (N_8710,N_7072,N_7489);
nand U8711 (N_8711,N_7077,N_7151);
or U8712 (N_8712,N_6562,N_6008);
nor U8713 (N_8713,N_6366,N_6519);
xnor U8714 (N_8714,N_6888,N_7176);
nand U8715 (N_8715,N_7676,N_7146);
nand U8716 (N_8716,N_7321,N_6244);
xnor U8717 (N_8717,N_6066,N_6167);
xnor U8718 (N_8718,N_6373,N_6068);
nand U8719 (N_8719,N_7538,N_7645);
xnor U8720 (N_8720,N_6295,N_6153);
nor U8721 (N_8721,N_6579,N_7767);
nand U8722 (N_8722,N_6293,N_6154);
nand U8723 (N_8723,N_6514,N_7673);
and U8724 (N_8724,N_7439,N_7298);
nor U8725 (N_8725,N_7375,N_6401);
nand U8726 (N_8726,N_6197,N_6846);
or U8727 (N_8727,N_6545,N_6267);
xnor U8728 (N_8728,N_7278,N_6168);
xnor U8729 (N_8729,N_6984,N_7329);
nand U8730 (N_8730,N_6855,N_6900);
xnor U8731 (N_8731,N_6919,N_7600);
or U8732 (N_8732,N_7574,N_7649);
or U8733 (N_8733,N_6688,N_7074);
nor U8734 (N_8734,N_6858,N_6702);
and U8735 (N_8735,N_6903,N_6692);
or U8736 (N_8736,N_7027,N_6132);
nor U8737 (N_8737,N_6298,N_6911);
xor U8738 (N_8738,N_6962,N_6170);
xnor U8739 (N_8739,N_6549,N_7413);
nand U8740 (N_8740,N_6095,N_7162);
and U8741 (N_8741,N_7678,N_7209);
nand U8742 (N_8742,N_6333,N_7247);
nand U8743 (N_8743,N_6559,N_7208);
nand U8744 (N_8744,N_6392,N_6893);
nand U8745 (N_8745,N_6214,N_7295);
and U8746 (N_8746,N_6235,N_7990);
xor U8747 (N_8747,N_7611,N_7047);
xnor U8748 (N_8748,N_6515,N_7081);
xnor U8749 (N_8749,N_7955,N_7527);
or U8750 (N_8750,N_6544,N_7914);
or U8751 (N_8751,N_6729,N_6567);
or U8752 (N_8752,N_7410,N_7537);
nor U8753 (N_8753,N_7186,N_7659);
xnor U8754 (N_8754,N_7596,N_7207);
and U8755 (N_8755,N_6136,N_6053);
and U8756 (N_8756,N_7689,N_7879);
and U8757 (N_8757,N_6690,N_6824);
or U8758 (N_8758,N_7284,N_7733);
xor U8759 (N_8759,N_6213,N_7418);
or U8760 (N_8760,N_7325,N_6186);
and U8761 (N_8761,N_7113,N_7599);
nand U8762 (N_8762,N_7136,N_6404);
and U8763 (N_8763,N_7109,N_6541);
xor U8764 (N_8764,N_7377,N_7387);
xnor U8765 (N_8765,N_7942,N_6966);
or U8766 (N_8766,N_6590,N_7682);
nand U8767 (N_8767,N_6406,N_7516);
nand U8768 (N_8768,N_6674,N_6098);
nand U8769 (N_8769,N_6319,N_6311);
nand U8770 (N_8770,N_7010,N_6686);
nand U8771 (N_8771,N_7904,N_6449);
xor U8772 (N_8772,N_7409,N_6364);
and U8773 (N_8773,N_6972,N_7775);
and U8774 (N_8774,N_7129,N_7134);
xnor U8775 (N_8775,N_6419,N_7119);
and U8776 (N_8776,N_7304,N_7824);
and U8777 (N_8777,N_6481,N_6608);
nor U8778 (N_8778,N_6538,N_6190);
and U8779 (N_8779,N_6997,N_7641);
or U8780 (N_8780,N_6288,N_7690);
nand U8781 (N_8781,N_6270,N_7210);
and U8782 (N_8782,N_7132,N_6716);
nor U8783 (N_8783,N_6182,N_7552);
xor U8784 (N_8784,N_6974,N_7061);
or U8785 (N_8785,N_6261,N_7161);
nor U8786 (N_8786,N_6456,N_7462);
nor U8787 (N_8787,N_6380,N_6335);
nand U8788 (N_8788,N_6330,N_7680);
nor U8789 (N_8789,N_6429,N_7467);
or U8790 (N_8790,N_7681,N_6505);
nand U8791 (N_8791,N_6049,N_6902);
xnor U8792 (N_8792,N_6122,N_7727);
xnor U8793 (N_8793,N_6912,N_7789);
nor U8794 (N_8794,N_6522,N_7434);
nand U8795 (N_8795,N_7766,N_7708);
and U8796 (N_8796,N_7948,N_7715);
nand U8797 (N_8797,N_6827,N_6156);
nor U8798 (N_8798,N_6717,N_7258);
or U8799 (N_8799,N_6817,N_6511);
nor U8800 (N_8800,N_6728,N_6371);
nor U8801 (N_8801,N_6968,N_7511);
nor U8802 (N_8802,N_6630,N_7003);
and U8803 (N_8803,N_7569,N_7340);
or U8804 (N_8804,N_7288,N_6604);
or U8805 (N_8805,N_6954,N_7943);
nor U8806 (N_8806,N_6744,N_6101);
nor U8807 (N_8807,N_6794,N_7310);
xor U8808 (N_8808,N_6593,N_6555);
nand U8809 (N_8809,N_6272,N_6813);
or U8810 (N_8810,N_7065,N_6970);
nand U8811 (N_8811,N_7441,N_7928);
and U8812 (N_8812,N_7499,N_6250);
nand U8813 (N_8813,N_7615,N_6268);
nand U8814 (N_8814,N_6277,N_7308);
and U8815 (N_8815,N_7895,N_7783);
xnor U8816 (N_8816,N_7967,N_6569);
nand U8817 (N_8817,N_6685,N_7204);
or U8818 (N_8818,N_7784,N_7213);
nor U8819 (N_8819,N_7941,N_7939);
xnor U8820 (N_8820,N_7579,N_6487);
or U8821 (N_8821,N_6260,N_7965);
or U8822 (N_8822,N_6501,N_6494);
and U8823 (N_8823,N_7164,N_7179);
or U8824 (N_8824,N_6976,N_7837);
and U8825 (N_8825,N_7950,N_6221);
or U8826 (N_8826,N_7934,N_7980);
and U8827 (N_8827,N_7244,N_7118);
nor U8828 (N_8828,N_6185,N_6412);
nand U8829 (N_8829,N_6062,N_6507);
or U8830 (N_8830,N_7973,N_6069);
nand U8831 (N_8831,N_7647,N_7455);
xnor U8832 (N_8832,N_7320,N_6212);
or U8833 (N_8833,N_7788,N_7954);
xnor U8834 (N_8834,N_7925,N_6196);
xor U8835 (N_8835,N_6109,N_7046);
nand U8836 (N_8836,N_6219,N_6249);
and U8837 (N_8837,N_6257,N_6283);
or U8838 (N_8838,N_6916,N_7381);
nor U8839 (N_8839,N_6526,N_7427);
nor U8840 (N_8840,N_6452,N_6808);
and U8841 (N_8841,N_7952,N_6571);
xnor U8842 (N_8842,N_6788,N_7536);
or U8843 (N_8843,N_7264,N_7068);
and U8844 (N_8844,N_6102,N_6045);
nand U8845 (N_8845,N_6473,N_7738);
and U8846 (N_8846,N_6786,N_7029);
and U8847 (N_8847,N_6376,N_7502);
or U8848 (N_8848,N_6163,N_6843);
and U8849 (N_8849,N_7585,N_7300);
nor U8850 (N_8850,N_7089,N_6437);
xnor U8851 (N_8851,N_6698,N_7684);
and U8852 (N_8852,N_7776,N_6611);
nor U8853 (N_8853,N_6695,N_7267);
or U8854 (N_8854,N_6262,N_6217);
nand U8855 (N_8855,N_6119,N_7430);
or U8856 (N_8856,N_6840,N_6826);
xor U8857 (N_8857,N_6104,N_7079);
and U8858 (N_8858,N_6988,N_7397);
or U8859 (N_8859,N_7165,N_6876);
or U8860 (N_8860,N_6483,N_7039);
xor U8861 (N_8861,N_6243,N_6047);
nand U8862 (N_8862,N_6051,N_6669);
xnor U8863 (N_8863,N_6478,N_7563);
nor U8864 (N_8864,N_6017,N_7360);
and U8865 (N_8865,N_6652,N_7894);
nand U8866 (N_8866,N_7881,N_7465);
nor U8867 (N_8867,N_7412,N_7245);
and U8868 (N_8868,N_6713,N_6615);
or U8869 (N_8869,N_7456,N_6625);
and U8870 (N_8870,N_7636,N_7256);
nand U8871 (N_8871,N_6561,N_6637);
nand U8872 (N_8872,N_6014,N_7890);
xor U8873 (N_8873,N_7933,N_7959);
or U8874 (N_8874,N_6745,N_7819);
xor U8875 (N_8875,N_7040,N_6343);
nor U8876 (N_8876,N_6833,N_7800);
nand U8877 (N_8877,N_6566,N_6143);
or U8878 (N_8878,N_7674,N_6318);
xor U8879 (N_8879,N_7963,N_6472);
nand U8880 (N_8880,N_6980,N_7883);
or U8881 (N_8881,N_7227,N_7125);
xnor U8882 (N_8882,N_7668,N_6597);
or U8883 (N_8883,N_6844,N_6273);
or U8884 (N_8884,N_7912,N_7804);
and U8885 (N_8885,N_6124,N_7226);
xnor U8886 (N_8886,N_7123,N_7045);
nor U8887 (N_8887,N_6476,N_6594);
and U8888 (N_8888,N_7460,N_6338);
or U8889 (N_8889,N_6328,N_7425);
or U8890 (N_8890,N_7031,N_6654);
nand U8891 (N_8891,N_7547,N_6942);
nor U8892 (N_8892,N_6572,N_6496);
nand U8893 (N_8893,N_6560,N_6183);
or U8894 (N_8894,N_6922,N_6134);
or U8895 (N_8895,N_7518,N_7841);
nor U8896 (N_8896,N_7345,N_7326);
nor U8897 (N_8897,N_6789,N_6275);
and U8898 (N_8898,N_7013,N_6000);
and U8899 (N_8899,N_7139,N_6956);
xnor U8900 (N_8900,N_6440,N_7217);
nand U8901 (N_8901,N_7806,N_7906);
nor U8902 (N_8902,N_7613,N_7588);
nand U8903 (N_8903,N_7171,N_6609);
nand U8904 (N_8904,N_7311,N_6670);
xor U8905 (N_8905,N_6898,N_6236);
xor U8906 (N_8906,N_7482,N_6093);
or U8907 (N_8907,N_7225,N_6946);
nand U8908 (N_8908,N_7876,N_6497);
nand U8909 (N_8909,N_6696,N_6780);
nor U8910 (N_8910,N_6582,N_6254);
nand U8911 (N_8911,N_7622,N_6276);
nand U8912 (N_8912,N_7551,N_7978);
or U8913 (N_8913,N_6626,N_6742);
nand U8914 (N_8914,N_6664,N_6034);
and U8915 (N_8915,N_7205,N_7986);
or U8916 (N_8916,N_6030,N_6861);
nand U8917 (N_8917,N_6421,N_6773);
xnor U8918 (N_8918,N_7483,N_6598);
xnor U8919 (N_8919,N_7564,N_7989);
or U8920 (N_8920,N_6204,N_6383);
xor U8921 (N_8921,N_7138,N_7472);
or U8922 (N_8922,N_7587,N_6719);
and U8923 (N_8923,N_6720,N_6578);
xor U8924 (N_8924,N_6362,N_6618);
nand U8925 (N_8925,N_7001,N_6767);
nor U8926 (N_8926,N_6570,N_7639);
and U8927 (N_8927,N_7867,N_7997);
nor U8928 (N_8928,N_7777,N_6752);
nor U8929 (N_8929,N_7023,N_7009);
and U8930 (N_8930,N_7729,N_6353);
nor U8931 (N_8931,N_7468,N_6035);
nor U8932 (N_8932,N_6816,N_6941);
xnor U8933 (N_8933,N_6884,N_7218);
xor U8934 (N_8934,N_6704,N_6469);
nand U8935 (N_8935,N_6303,N_7975);
nand U8936 (N_8936,N_6967,N_7422);
nor U8937 (N_8937,N_6760,N_6088);
nor U8938 (N_8938,N_7297,N_6038);
or U8939 (N_8939,N_7043,N_7597);
and U8940 (N_8940,N_6820,N_6895);
nand U8941 (N_8941,N_6796,N_7524);
and U8942 (N_8942,N_7522,N_6758);
nor U8943 (N_8943,N_6209,N_7274);
nand U8944 (N_8944,N_7007,N_6291);
nor U8945 (N_8945,N_7982,N_6628);
and U8946 (N_8946,N_7156,N_6774);
nor U8947 (N_8947,N_6023,N_6543);
nand U8948 (N_8948,N_7316,N_7843);
nand U8949 (N_8949,N_6029,N_7623);
nand U8950 (N_8950,N_6231,N_6869);
nand U8951 (N_8951,N_7111,N_7021);
nor U8952 (N_8952,N_7414,N_6006);
nor U8953 (N_8953,N_7239,N_6103);
nand U8954 (N_8954,N_6706,N_7017);
nor U8955 (N_8955,N_6193,N_6176);
or U8956 (N_8956,N_6969,N_6763);
or U8957 (N_8957,N_6588,N_7509);
and U8958 (N_8958,N_6677,N_7299);
nor U8959 (N_8959,N_7559,N_7754);
or U8960 (N_8960,N_6580,N_7741);
and U8961 (N_8961,N_7885,N_7248);
nor U8962 (N_8962,N_7076,N_7578);
xnor U8963 (N_8963,N_6286,N_7504);
xnor U8964 (N_8964,N_7167,N_7168);
nor U8965 (N_8965,N_6377,N_7799);
nor U8966 (N_8966,N_7836,N_7655);
nand U8967 (N_8967,N_6179,N_7175);
nand U8968 (N_8968,N_7812,N_6857);
or U8969 (N_8969,N_6958,N_6346);
xnor U8970 (N_8970,N_6423,N_6564);
xnor U8971 (N_8971,N_7526,N_6480);
nor U8972 (N_8972,N_7083,N_7251);
xor U8973 (N_8973,N_7642,N_7573);
xor U8974 (N_8974,N_7886,N_6080);
or U8975 (N_8975,N_7108,N_6166);
and U8976 (N_8976,N_7135,N_6207);
or U8977 (N_8977,N_7044,N_7327);
or U8978 (N_8978,N_7294,N_6985);
nand U8979 (N_8979,N_6299,N_6357);
xnor U8980 (N_8980,N_7938,N_7318);
or U8981 (N_8981,N_7206,N_7231);
nand U8982 (N_8982,N_6458,N_6657);
and U8983 (N_8983,N_6595,N_6076);
or U8984 (N_8984,N_6815,N_6281);
or U8985 (N_8985,N_7464,N_6087);
or U8986 (N_8986,N_6425,N_7383);
nor U8987 (N_8987,N_6860,N_6370);
or U8988 (N_8988,N_7900,N_7443);
nand U8989 (N_8989,N_7028,N_7313);
nand U8990 (N_8990,N_7102,N_7148);
xnor U8991 (N_8991,N_7393,N_6381);
xor U8992 (N_8992,N_6300,N_6165);
and U8993 (N_8993,N_7160,N_7032);
or U8994 (N_8994,N_7769,N_7632);
nand U8995 (N_8995,N_7440,N_7268);
nor U8996 (N_8996,N_6081,N_7734);
or U8997 (N_8997,N_6612,N_6074);
nor U8998 (N_8998,N_7625,N_7396);
and U8999 (N_8999,N_7201,N_6220);
and U9000 (N_9000,N_7078,N_7950);
nor U9001 (N_9001,N_7877,N_6009);
or U9002 (N_9002,N_7193,N_6695);
nor U9003 (N_9003,N_7986,N_6928);
xnor U9004 (N_9004,N_6463,N_7286);
nor U9005 (N_9005,N_6491,N_6333);
nand U9006 (N_9006,N_7399,N_7775);
or U9007 (N_9007,N_6549,N_6389);
or U9008 (N_9008,N_7547,N_7970);
or U9009 (N_9009,N_6021,N_6390);
xnor U9010 (N_9010,N_6657,N_6957);
xor U9011 (N_9011,N_6023,N_6521);
xnor U9012 (N_9012,N_7576,N_7763);
and U9013 (N_9013,N_7449,N_6701);
xor U9014 (N_9014,N_7440,N_7912);
or U9015 (N_9015,N_7035,N_6562);
nor U9016 (N_9016,N_7979,N_6168);
or U9017 (N_9017,N_6917,N_7812);
nor U9018 (N_9018,N_7606,N_6413);
xor U9019 (N_9019,N_6756,N_7966);
and U9020 (N_9020,N_7248,N_7089);
xor U9021 (N_9021,N_7609,N_6123);
nand U9022 (N_9022,N_7378,N_7223);
or U9023 (N_9023,N_6211,N_7616);
or U9024 (N_9024,N_7990,N_7094);
xor U9025 (N_9025,N_6328,N_6468);
nor U9026 (N_9026,N_7616,N_7054);
nor U9027 (N_9027,N_7846,N_6927);
xnor U9028 (N_9028,N_6751,N_7868);
or U9029 (N_9029,N_6981,N_7262);
and U9030 (N_9030,N_7985,N_6290);
xnor U9031 (N_9031,N_7772,N_6176);
nor U9032 (N_9032,N_6168,N_7636);
nor U9033 (N_9033,N_7762,N_7213);
or U9034 (N_9034,N_6214,N_7108);
or U9035 (N_9035,N_7094,N_6180);
and U9036 (N_9036,N_6127,N_7267);
xnor U9037 (N_9037,N_6381,N_7976);
and U9038 (N_9038,N_6493,N_6658);
and U9039 (N_9039,N_7030,N_7506);
xor U9040 (N_9040,N_6352,N_7272);
or U9041 (N_9041,N_7046,N_7255);
xor U9042 (N_9042,N_7632,N_6769);
xor U9043 (N_9043,N_6334,N_7614);
nand U9044 (N_9044,N_6680,N_7675);
and U9045 (N_9045,N_7413,N_7822);
nand U9046 (N_9046,N_7777,N_7474);
xor U9047 (N_9047,N_6341,N_6170);
or U9048 (N_9048,N_7756,N_7764);
or U9049 (N_9049,N_7795,N_7522);
xnor U9050 (N_9050,N_7192,N_7854);
and U9051 (N_9051,N_7944,N_6018);
nor U9052 (N_9052,N_6320,N_7448);
nand U9053 (N_9053,N_6949,N_7060);
or U9054 (N_9054,N_6976,N_7054);
xor U9055 (N_9055,N_6674,N_7463);
or U9056 (N_9056,N_6771,N_7052);
and U9057 (N_9057,N_7385,N_7640);
nor U9058 (N_9058,N_7806,N_6119);
xnor U9059 (N_9059,N_7185,N_6812);
nand U9060 (N_9060,N_7265,N_7457);
or U9061 (N_9061,N_7448,N_6432);
and U9062 (N_9062,N_6205,N_6976);
nor U9063 (N_9063,N_7570,N_6111);
nand U9064 (N_9064,N_7074,N_6982);
xnor U9065 (N_9065,N_7701,N_7614);
or U9066 (N_9066,N_6455,N_6458);
nand U9067 (N_9067,N_7766,N_6947);
nor U9068 (N_9068,N_7841,N_7123);
and U9069 (N_9069,N_6610,N_6476);
nor U9070 (N_9070,N_6722,N_6621);
nand U9071 (N_9071,N_6851,N_7218);
xnor U9072 (N_9072,N_6710,N_7873);
or U9073 (N_9073,N_6209,N_7024);
nor U9074 (N_9074,N_7130,N_7102);
xor U9075 (N_9075,N_6508,N_6390);
and U9076 (N_9076,N_7853,N_7687);
nand U9077 (N_9077,N_6824,N_7903);
and U9078 (N_9078,N_7439,N_7320);
or U9079 (N_9079,N_6399,N_7913);
or U9080 (N_9080,N_7689,N_7974);
nand U9081 (N_9081,N_6204,N_7241);
nor U9082 (N_9082,N_6866,N_7576);
nor U9083 (N_9083,N_6163,N_6370);
xor U9084 (N_9084,N_7319,N_7583);
and U9085 (N_9085,N_6077,N_6168);
nor U9086 (N_9086,N_6556,N_7808);
or U9087 (N_9087,N_7614,N_7096);
xnor U9088 (N_9088,N_7107,N_6863);
nand U9089 (N_9089,N_7146,N_7137);
or U9090 (N_9090,N_7052,N_6383);
nor U9091 (N_9091,N_6722,N_6412);
or U9092 (N_9092,N_6354,N_7989);
nand U9093 (N_9093,N_6798,N_6806);
or U9094 (N_9094,N_6068,N_6746);
or U9095 (N_9095,N_6205,N_6332);
and U9096 (N_9096,N_6859,N_6739);
or U9097 (N_9097,N_6759,N_7180);
or U9098 (N_9098,N_6449,N_6393);
or U9099 (N_9099,N_6365,N_7084);
xnor U9100 (N_9100,N_6130,N_7521);
and U9101 (N_9101,N_6024,N_6047);
or U9102 (N_9102,N_6354,N_7598);
xnor U9103 (N_9103,N_7267,N_6125);
nand U9104 (N_9104,N_6310,N_7171);
nand U9105 (N_9105,N_6269,N_7127);
nor U9106 (N_9106,N_6219,N_6522);
or U9107 (N_9107,N_6475,N_7925);
nor U9108 (N_9108,N_6732,N_7746);
or U9109 (N_9109,N_7724,N_7463);
nand U9110 (N_9110,N_7501,N_6558);
xor U9111 (N_9111,N_6603,N_7605);
xnor U9112 (N_9112,N_6934,N_7623);
nor U9113 (N_9113,N_7973,N_6302);
xor U9114 (N_9114,N_6671,N_6398);
nor U9115 (N_9115,N_7909,N_6416);
and U9116 (N_9116,N_7749,N_7563);
nand U9117 (N_9117,N_7896,N_6104);
or U9118 (N_9118,N_7984,N_7030);
xnor U9119 (N_9119,N_6664,N_6868);
or U9120 (N_9120,N_7888,N_7246);
and U9121 (N_9121,N_7138,N_6521);
xor U9122 (N_9122,N_7341,N_6902);
or U9123 (N_9123,N_7873,N_7768);
nand U9124 (N_9124,N_6026,N_7962);
and U9125 (N_9125,N_7270,N_6836);
nand U9126 (N_9126,N_6970,N_6089);
and U9127 (N_9127,N_6395,N_7682);
nand U9128 (N_9128,N_7837,N_7251);
and U9129 (N_9129,N_6998,N_7960);
nand U9130 (N_9130,N_7624,N_6997);
xnor U9131 (N_9131,N_7921,N_7177);
xnor U9132 (N_9132,N_7509,N_6742);
and U9133 (N_9133,N_7585,N_6163);
or U9134 (N_9134,N_7039,N_7165);
and U9135 (N_9135,N_7287,N_6004);
or U9136 (N_9136,N_7672,N_7996);
or U9137 (N_9137,N_6269,N_7983);
nor U9138 (N_9138,N_7500,N_7988);
or U9139 (N_9139,N_6273,N_7356);
nor U9140 (N_9140,N_7446,N_6183);
and U9141 (N_9141,N_6993,N_6407);
xnor U9142 (N_9142,N_7903,N_7265);
xor U9143 (N_9143,N_6975,N_7765);
xor U9144 (N_9144,N_6832,N_7797);
nand U9145 (N_9145,N_6357,N_7074);
and U9146 (N_9146,N_6163,N_6406);
and U9147 (N_9147,N_6674,N_7968);
and U9148 (N_9148,N_6758,N_6485);
and U9149 (N_9149,N_6718,N_6203);
nor U9150 (N_9150,N_7379,N_6679);
nand U9151 (N_9151,N_7394,N_6275);
and U9152 (N_9152,N_6318,N_7037);
or U9153 (N_9153,N_7095,N_6925);
or U9154 (N_9154,N_6192,N_7407);
nand U9155 (N_9155,N_6491,N_7949);
and U9156 (N_9156,N_7942,N_6491);
or U9157 (N_9157,N_7881,N_6422);
nor U9158 (N_9158,N_6547,N_7433);
xor U9159 (N_9159,N_6291,N_6158);
xor U9160 (N_9160,N_7335,N_7951);
nor U9161 (N_9161,N_6684,N_7876);
and U9162 (N_9162,N_6053,N_6238);
xor U9163 (N_9163,N_6572,N_6699);
xnor U9164 (N_9164,N_6616,N_6125);
xnor U9165 (N_9165,N_7173,N_7607);
nor U9166 (N_9166,N_7201,N_7531);
nand U9167 (N_9167,N_6305,N_7105);
xnor U9168 (N_9168,N_6854,N_6574);
and U9169 (N_9169,N_7736,N_7414);
nand U9170 (N_9170,N_6712,N_7652);
xor U9171 (N_9171,N_7824,N_7855);
or U9172 (N_9172,N_6972,N_7299);
or U9173 (N_9173,N_6112,N_6039);
nor U9174 (N_9174,N_6467,N_6793);
nand U9175 (N_9175,N_7173,N_6038);
nand U9176 (N_9176,N_6993,N_7401);
xor U9177 (N_9177,N_6640,N_7223);
or U9178 (N_9178,N_7431,N_7383);
xor U9179 (N_9179,N_7864,N_7589);
and U9180 (N_9180,N_6205,N_7313);
nor U9181 (N_9181,N_6878,N_7586);
xnor U9182 (N_9182,N_7112,N_7582);
and U9183 (N_9183,N_6113,N_7313);
or U9184 (N_9184,N_7687,N_6421);
and U9185 (N_9185,N_7524,N_7784);
nor U9186 (N_9186,N_7506,N_6744);
xor U9187 (N_9187,N_7282,N_6566);
nor U9188 (N_9188,N_6124,N_7539);
nand U9189 (N_9189,N_6649,N_6529);
and U9190 (N_9190,N_7203,N_6056);
nand U9191 (N_9191,N_7738,N_7791);
nand U9192 (N_9192,N_6525,N_7089);
xor U9193 (N_9193,N_6919,N_6801);
nor U9194 (N_9194,N_6784,N_6010);
nand U9195 (N_9195,N_7011,N_7252);
or U9196 (N_9196,N_6853,N_7942);
and U9197 (N_9197,N_6505,N_6467);
xor U9198 (N_9198,N_6674,N_6356);
or U9199 (N_9199,N_6549,N_7364);
nand U9200 (N_9200,N_7794,N_7992);
nand U9201 (N_9201,N_7685,N_6521);
xor U9202 (N_9202,N_6439,N_7482);
or U9203 (N_9203,N_6280,N_6076);
nand U9204 (N_9204,N_7420,N_6720);
and U9205 (N_9205,N_7035,N_7019);
and U9206 (N_9206,N_6653,N_7648);
or U9207 (N_9207,N_7683,N_6832);
or U9208 (N_9208,N_7995,N_7799);
nor U9209 (N_9209,N_6512,N_6679);
and U9210 (N_9210,N_7195,N_7945);
nand U9211 (N_9211,N_7488,N_6520);
nand U9212 (N_9212,N_7016,N_6893);
and U9213 (N_9213,N_7557,N_7291);
and U9214 (N_9214,N_7757,N_7669);
xor U9215 (N_9215,N_6467,N_6226);
nand U9216 (N_9216,N_7101,N_6360);
nand U9217 (N_9217,N_6905,N_6909);
and U9218 (N_9218,N_6354,N_7182);
and U9219 (N_9219,N_6830,N_6234);
xnor U9220 (N_9220,N_7314,N_7088);
and U9221 (N_9221,N_7638,N_6220);
and U9222 (N_9222,N_6137,N_7480);
nor U9223 (N_9223,N_7265,N_7156);
nor U9224 (N_9224,N_7307,N_6913);
or U9225 (N_9225,N_7724,N_6283);
xnor U9226 (N_9226,N_7178,N_7109);
xor U9227 (N_9227,N_6818,N_6404);
or U9228 (N_9228,N_6761,N_7975);
or U9229 (N_9229,N_7869,N_6611);
nand U9230 (N_9230,N_7867,N_6081);
xnor U9231 (N_9231,N_6173,N_7947);
or U9232 (N_9232,N_6473,N_6990);
nand U9233 (N_9233,N_6377,N_7760);
nand U9234 (N_9234,N_6156,N_7890);
nor U9235 (N_9235,N_6884,N_6627);
or U9236 (N_9236,N_7765,N_6293);
nor U9237 (N_9237,N_6099,N_7741);
xnor U9238 (N_9238,N_6027,N_7774);
xnor U9239 (N_9239,N_6032,N_6686);
nand U9240 (N_9240,N_7044,N_6215);
or U9241 (N_9241,N_6459,N_6581);
and U9242 (N_9242,N_6544,N_7676);
or U9243 (N_9243,N_6244,N_7580);
nor U9244 (N_9244,N_7064,N_7208);
nor U9245 (N_9245,N_6106,N_6558);
nor U9246 (N_9246,N_7056,N_6871);
or U9247 (N_9247,N_6868,N_6950);
and U9248 (N_9248,N_7902,N_7159);
or U9249 (N_9249,N_7707,N_7354);
and U9250 (N_9250,N_6126,N_7263);
or U9251 (N_9251,N_7159,N_7061);
nand U9252 (N_9252,N_7548,N_7050);
nor U9253 (N_9253,N_7861,N_7495);
nor U9254 (N_9254,N_7873,N_7854);
and U9255 (N_9255,N_6142,N_7866);
or U9256 (N_9256,N_7179,N_6201);
and U9257 (N_9257,N_7373,N_7452);
nor U9258 (N_9258,N_7847,N_6020);
or U9259 (N_9259,N_7524,N_7564);
nand U9260 (N_9260,N_6616,N_6040);
nand U9261 (N_9261,N_7390,N_7611);
and U9262 (N_9262,N_7398,N_7761);
xnor U9263 (N_9263,N_7289,N_7114);
nand U9264 (N_9264,N_6582,N_6649);
and U9265 (N_9265,N_6340,N_6613);
nand U9266 (N_9266,N_7951,N_7888);
xnor U9267 (N_9267,N_7416,N_7983);
or U9268 (N_9268,N_7373,N_7701);
nor U9269 (N_9269,N_7747,N_7725);
xor U9270 (N_9270,N_6780,N_6765);
nor U9271 (N_9271,N_7037,N_6600);
and U9272 (N_9272,N_7711,N_6614);
nor U9273 (N_9273,N_7139,N_6119);
xnor U9274 (N_9274,N_7591,N_7058);
and U9275 (N_9275,N_7314,N_7560);
xnor U9276 (N_9276,N_6986,N_6448);
xnor U9277 (N_9277,N_6086,N_7114);
nand U9278 (N_9278,N_7453,N_6887);
or U9279 (N_9279,N_6071,N_7290);
nor U9280 (N_9280,N_6232,N_6827);
nor U9281 (N_9281,N_6092,N_7411);
or U9282 (N_9282,N_6090,N_7752);
and U9283 (N_9283,N_6482,N_7739);
nor U9284 (N_9284,N_7907,N_7240);
xor U9285 (N_9285,N_6391,N_7214);
and U9286 (N_9286,N_7822,N_7974);
nor U9287 (N_9287,N_6718,N_7627);
or U9288 (N_9288,N_7532,N_7925);
or U9289 (N_9289,N_7324,N_7202);
xor U9290 (N_9290,N_6622,N_6312);
and U9291 (N_9291,N_7740,N_6108);
xnor U9292 (N_9292,N_6414,N_6456);
nand U9293 (N_9293,N_6417,N_6747);
nand U9294 (N_9294,N_7713,N_7402);
and U9295 (N_9295,N_6124,N_7983);
nor U9296 (N_9296,N_7938,N_6701);
and U9297 (N_9297,N_7433,N_7040);
xor U9298 (N_9298,N_6794,N_7554);
or U9299 (N_9299,N_6284,N_6614);
nand U9300 (N_9300,N_7685,N_7504);
nand U9301 (N_9301,N_7633,N_6727);
and U9302 (N_9302,N_6205,N_6612);
or U9303 (N_9303,N_6224,N_6032);
or U9304 (N_9304,N_6541,N_7048);
nand U9305 (N_9305,N_7696,N_7919);
nand U9306 (N_9306,N_6648,N_7808);
and U9307 (N_9307,N_7170,N_6256);
or U9308 (N_9308,N_7978,N_6183);
xor U9309 (N_9309,N_7674,N_7135);
and U9310 (N_9310,N_6425,N_6870);
and U9311 (N_9311,N_7360,N_7058);
nand U9312 (N_9312,N_7556,N_6941);
and U9313 (N_9313,N_6807,N_6897);
or U9314 (N_9314,N_6055,N_6092);
xor U9315 (N_9315,N_6957,N_6372);
nor U9316 (N_9316,N_7916,N_6475);
nand U9317 (N_9317,N_6912,N_6406);
or U9318 (N_9318,N_6081,N_6755);
and U9319 (N_9319,N_6541,N_7378);
nor U9320 (N_9320,N_6551,N_7765);
or U9321 (N_9321,N_7254,N_7747);
or U9322 (N_9322,N_6395,N_6719);
and U9323 (N_9323,N_6941,N_7320);
or U9324 (N_9324,N_7283,N_6377);
xor U9325 (N_9325,N_6721,N_6926);
and U9326 (N_9326,N_6461,N_6370);
nor U9327 (N_9327,N_6540,N_7880);
xor U9328 (N_9328,N_7125,N_6513);
xor U9329 (N_9329,N_7694,N_6465);
or U9330 (N_9330,N_6069,N_7072);
nor U9331 (N_9331,N_7019,N_6565);
nor U9332 (N_9332,N_7088,N_6104);
and U9333 (N_9333,N_6590,N_7289);
and U9334 (N_9334,N_6250,N_7366);
and U9335 (N_9335,N_7197,N_6100);
nand U9336 (N_9336,N_7896,N_7201);
and U9337 (N_9337,N_6266,N_7254);
nor U9338 (N_9338,N_7341,N_7967);
nand U9339 (N_9339,N_7423,N_6693);
and U9340 (N_9340,N_6286,N_6411);
nand U9341 (N_9341,N_7712,N_7853);
nor U9342 (N_9342,N_6829,N_6455);
or U9343 (N_9343,N_7012,N_6625);
nor U9344 (N_9344,N_7757,N_6820);
nor U9345 (N_9345,N_7584,N_7382);
nand U9346 (N_9346,N_6706,N_6396);
xnor U9347 (N_9347,N_6138,N_6237);
or U9348 (N_9348,N_6444,N_7803);
nand U9349 (N_9349,N_7195,N_6230);
xnor U9350 (N_9350,N_7219,N_7794);
or U9351 (N_9351,N_6708,N_6560);
and U9352 (N_9352,N_7697,N_7497);
and U9353 (N_9353,N_7619,N_6923);
and U9354 (N_9354,N_7700,N_6652);
and U9355 (N_9355,N_6514,N_6878);
xnor U9356 (N_9356,N_6739,N_7011);
nor U9357 (N_9357,N_7425,N_6406);
nor U9358 (N_9358,N_7553,N_6056);
and U9359 (N_9359,N_6183,N_7778);
nor U9360 (N_9360,N_7018,N_6020);
xnor U9361 (N_9361,N_6457,N_6229);
and U9362 (N_9362,N_7953,N_6897);
xnor U9363 (N_9363,N_7324,N_6709);
nor U9364 (N_9364,N_6782,N_7241);
and U9365 (N_9365,N_6052,N_7783);
nand U9366 (N_9366,N_7414,N_7212);
or U9367 (N_9367,N_7699,N_7192);
nor U9368 (N_9368,N_6485,N_6134);
or U9369 (N_9369,N_7540,N_7489);
nand U9370 (N_9370,N_7921,N_7622);
nand U9371 (N_9371,N_6854,N_6933);
and U9372 (N_9372,N_7887,N_6428);
and U9373 (N_9373,N_6530,N_7512);
and U9374 (N_9374,N_7414,N_6248);
and U9375 (N_9375,N_6925,N_6364);
nand U9376 (N_9376,N_7833,N_6826);
xor U9377 (N_9377,N_6228,N_7359);
and U9378 (N_9378,N_7258,N_7750);
and U9379 (N_9379,N_7383,N_6295);
xor U9380 (N_9380,N_7394,N_6326);
nand U9381 (N_9381,N_7497,N_6547);
nor U9382 (N_9382,N_6833,N_6408);
xnor U9383 (N_9383,N_6069,N_7316);
or U9384 (N_9384,N_6996,N_6407);
xor U9385 (N_9385,N_6312,N_6130);
nor U9386 (N_9386,N_7065,N_7899);
and U9387 (N_9387,N_7644,N_6156);
xnor U9388 (N_9388,N_7585,N_6097);
xor U9389 (N_9389,N_7378,N_6559);
or U9390 (N_9390,N_6764,N_6480);
and U9391 (N_9391,N_6192,N_6790);
nor U9392 (N_9392,N_7036,N_6297);
or U9393 (N_9393,N_7018,N_7862);
and U9394 (N_9394,N_7869,N_6574);
or U9395 (N_9395,N_7663,N_7076);
or U9396 (N_9396,N_6244,N_6177);
nand U9397 (N_9397,N_6510,N_7004);
xnor U9398 (N_9398,N_6900,N_7397);
or U9399 (N_9399,N_6863,N_7744);
and U9400 (N_9400,N_7237,N_6018);
nand U9401 (N_9401,N_7844,N_7558);
nor U9402 (N_9402,N_6898,N_7288);
nand U9403 (N_9403,N_7640,N_6220);
nor U9404 (N_9404,N_6157,N_7511);
nand U9405 (N_9405,N_6435,N_6682);
nand U9406 (N_9406,N_7697,N_7902);
nor U9407 (N_9407,N_7114,N_7355);
nor U9408 (N_9408,N_7020,N_6914);
nor U9409 (N_9409,N_6360,N_6726);
or U9410 (N_9410,N_6226,N_6144);
nor U9411 (N_9411,N_7468,N_6136);
and U9412 (N_9412,N_7131,N_7758);
or U9413 (N_9413,N_6906,N_7073);
and U9414 (N_9414,N_6767,N_6010);
and U9415 (N_9415,N_6775,N_6286);
xor U9416 (N_9416,N_6198,N_6910);
and U9417 (N_9417,N_7281,N_6649);
nor U9418 (N_9418,N_6710,N_6095);
xor U9419 (N_9419,N_6751,N_7171);
nand U9420 (N_9420,N_7453,N_6102);
and U9421 (N_9421,N_6885,N_6469);
nor U9422 (N_9422,N_6939,N_6663);
or U9423 (N_9423,N_7383,N_7704);
nor U9424 (N_9424,N_6407,N_7177);
nor U9425 (N_9425,N_6228,N_6498);
nor U9426 (N_9426,N_6464,N_7348);
nand U9427 (N_9427,N_7715,N_7544);
and U9428 (N_9428,N_7303,N_6832);
nor U9429 (N_9429,N_6918,N_6649);
or U9430 (N_9430,N_7004,N_7632);
or U9431 (N_9431,N_6627,N_6988);
and U9432 (N_9432,N_6668,N_6017);
nand U9433 (N_9433,N_6756,N_7846);
nand U9434 (N_9434,N_6167,N_6996);
and U9435 (N_9435,N_7493,N_6437);
and U9436 (N_9436,N_6253,N_7834);
and U9437 (N_9437,N_6453,N_6920);
nand U9438 (N_9438,N_6749,N_6268);
nand U9439 (N_9439,N_6843,N_6275);
and U9440 (N_9440,N_6918,N_7278);
or U9441 (N_9441,N_6010,N_7629);
and U9442 (N_9442,N_7011,N_6079);
or U9443 (N_9443,N_7755,N_6984);
or U9444 (N_9444,N_7782,N_7391);
nand U9445 (N_9445,N_7514,N_7818);
nand U9446 (N_9446,N_7202,N_7623);
nand U9447 (N_9447,N_7569,N_7356);
xnor U9448 (N_9448,N_7515,N_6091);
or U9449 (N_9449,N_6338,N_6334);
and U9450 (N_9450,N_7532,N_6287);
or U9451 (N_9451,N_6027,N_7714);
xnor U9452 (N_9452,N_6974,N_7196);
or U9453 (N_9453,N_7571,N_6917);
xor U9454 (N_9454,N_6201,N_7225);
xor U9455 (N_9455,N_7352,N_6183);
xor U9456 (N_9456,N_7514,N_7580);
and U9457 (N_9457,N_7384,N_6835);
nor U9458 (N_9458,N_6346,N_6845);
nand U9459 (N_9459,N_7240,N_6532);
and U9460 (N_9460,N_6067,N_6314);
nand U9461 (N_9461,N_7491,N_6918);
xnor U9462 (N_9462,N_6022,N_6433);
and U9463 (N_9463,N_6496,N_7581);
xnor U9464 (N_9464,N_6590,N_6912);
and U9465 (N_9465,N_7473,N_6158);
xnor U9466 (N_9466,N_7196,N_6203);
xnor U9467 (N_9467,N_6456,N_6964);
nand U9468 (N_9468,N_7430,N_6568);
xor U9469 (N_9469,N_6779,N_6784);
xor U9470 (N_9470,N_7489,N_7532);
and U9471 (N_9471,N_6893,N_6133);
nor U9472 (N_9472,N_7544,N_7796);
nand U9473 (N_9473,N_6282,N_6782);
nand U9474 (N_9474,N_6430,N_7812);
nand U9475 (N_9475,N_6773,N_7953);
nand U9476 (N_9476,N_7482,N_7236);
and U9477 (N_9477,N_6488,N_7257);
or U9478 (N_9478,N_6363,N_6643);
or U9479 (N_9479,N_6100,N_7387);
and U9480 (N_9480,N_7718,N_6737);
xor U9481 (N_9481,N_6228,N_6064);
or U9482 (N_9482,N_6420,N_7008);
xor U9483 (N_9483,N_7283,N_7402);
and U9484 (N_9484,N_6767,N_7886);
xnor U9485 (N_9485,N_7331,N_7358);
xor U9486 (N_9486,N_7377,N_6204);
xor U9487 (N_9487,N_7187,N_6143);
and U9488 (N_9488,N_6955,N_6793);
and U9489 (N_9489,N_6452,N_7573);
or U9490 (N_9490,N_7915,N_7174);
or U9491 (N_9491,N_7425,N_7429);
nor U9492 (N_9492,N_6300,N_6570);
xor U9493 (N_9493,N_6651,N_6614);
or U9494 (N_9494,N_6493,N_6215);
nor U9495 (N_9495,N_7898,N_7847);
xnor U9496 (N_9496,N_7099,N_7073);
and U9497 (N_9497,N_7333,N_7195);
or U9498 (N_9498,N_7613,N_6748);
xnor U9499 (N_9499,N_7016,N_6442);
and U9500 (N_9500,N_6628,N_6292);
or U9501 (N_9501,N_7299,N_6428);
and U9502 (N_9502,N_6930,N_7948);
and U9503 (N_9503,N_7261,N_6749);
xor U9504 (N_9504,N_6844,N_7324);
or U9505 (N_9505,N_6968,N_7418);
and U9506 (N_9506,N_6064,N_7170);
nand U9507 (N_9507,N_6222,N_7320);
nor U9508 (N_9508,N_7040,N_6721);
nor U9509 (N_9509,N_7517,N_7863);
nor U9510 (N_9510,N_6743,N_7337);
xor U9511 (N_9511,N_7426,N_7443);
or U9512 (N_9512,N_6415,N_6160);
nor U9513 (N_9513,N_6048,N_6505);
and U9514 (N_9514,N_6811,N_6372);
and U9515 (N_9515,N_6510,N_7750);
nand U9516 (N_9516,N_7377,N_6998);
or U9517 (N_9517,N_7469,N_7200);
and U9518 (N_9518,N_7782,N_6835);
xor U9519 (N_9519,N_7464,N_7964);
and U9520 (N_9520,N_7113,N_6786);
nor U9521 (N_9521,N_6035,N_7772);
nor U9522 (N_9522,N_7166,N_6506);
or U9523 (N_9523,N_6702,N_7526);
nor U9524 (N_9524,N_6250,N_6386);
nand U9525 (N_9525,N_6352,N_7366);
nor U9526 (N_9526,N_7334,N_7097);
xor U9527 (N_9527,N_6689,N_7636);
xor U9528 (N_9528,N_7985,N_6713);
and U9529 (N_9529,N_6867,N_6730);
or U9530 (N_9530,N_7199,N_6976);
or U9531 (N_9531,N_7106,N_7679);
and U9532 (N_9532,N_6202,N_6360);
and U9533 (N_9533,N_7435,N_6685);
nor U9534 (N_9534,N_6230,N_7228);
nand U9535 (N_9535,N_6379,N_6181);
or U9536 (N_9536,N_6179,N_7687);
or U9537 (N_9537,N_7928,N_7973);
or U9538 (N_9538,N_7967,N_6277);
nand U9539 (N_9539,N_6193,N_6400);
or U9540 (N_9540,N_7997,N_7983);
xor U9541 (N_9541,N_6812,N_6035);
or U9542 (N_9542,N_7239,N_6600);
or U9543 (N_9543,N_7371,N_6999);
and U9544 (N_9544,N_6906,N_6377);
nor U9545 (N_9545,N_6089,N_7555);
or U9546 (N_9546,N_6221,N_6762);
and U9547 (N_9547,N_7299,N_7488);
xor U9548 (N_9548,N_6071,N_6572);
or U9549 (N_9549,N_6000,N_7570);
and U9550 (N_9550,N_6802,N_7732);
xnor U9551 (N_9551,N_6507,N_6958);
or U9552 (N_9552,N_6806,N_7807);
or U9553 (N_9553,N_6557,N_6605);
nor U9554 (N_9554,N_7520,N_7417);
or U9555 (N_9555,N_6069,N_7028);
and U9556 (N_9556,N_7031,N_6002);
or U9557 (N_9557,N_6970,N_7732);
and U9558 (N_9558,N_6875,N_6307);
and U9559 (N_9559,N_6805,N_7174);
nand U9560 (N_9560,N_7455,N_7703);
or U9561 (N_9561,N_6559,N_7481);
or U9562 (N_9562,N_6048,N_6450);
and U9563 (N_9563,N_6350,N_7555);
or U9564 (N_9564,N_6834,N_7382);
and U9565 (N_9565,N_7128,N_7516);
nand U9566 (N_9566,N_6953,N_6042);
and U9567 (N_9567,N_6808,N_6702);
xor U9568 (N_9568,N_6176,N_6240);
nor U9569 (N_9569,N_7626,N_7312);
or U9570 (N_9570,N_6136,N_7475);
nor U9571 (N_9571,N_7487,N_7302);
xor U9572 (N_9572,N_6912,N_6154);
nor U9573 (N_9573,N_6974,N_7083);
xor U9574 (N_9574,N_6792,N_6007);
nand U9575 (N_9575,N_7818,N_7991);
nor U9576 (N_9576,N_7078,N_7392);
and U9577 (N_9577,N_7144,N_7852);
nand U9578 (N_9578,N_7181,N_7485);
nand U9579 (N_9579,N_7776,N_7499);
nand U9580 (N_9580,N_6686,N_7343);
xnor U9581 (N_9581,N_6080,N_7396);
or U9582 (N_9582,N_6574,N_6924);
and U9583 (N_9583,N_7303,N_6294);
and U9584 (N_9584,N_6401,N_7978);
and U9585 (N_9585,N_6825,N_7499);
xor U9586 (N_9586,N_6066,N_7562);
xnor U9587 (N_9587,N_6300,N_7854);
and U9588 (N_9588,N_6110,N_7206);
and U9589 (N_9589,N_6126,N_7637);
nor U9590 (N_9590,N_7124,N_6555);
nand U9591 (N_9591,N_6831,N_6481);
or U9592 (N_9592,N_6726,N_6267);
and U9593 (N_9593,N_7465,N_7301);
nand U9594 (N_9594,N_7785,N_7029);
xor U9595 (N_9595,N_6123,N_7606);
or U9596 (N_9596,N_7101,N_7947);
or U9597 (N_9597,N_6355,N_7803);
xnor U9598 (N_9598,N_6493,N_7312);
nor U9599 (N_9599,N_6308,N_7653);
nand U9600 (N_9600,N_6029,N_6170);
xor U9601 (N_9601,N_7851,N_7332);
nand U9602 (N_9602,N_7076,N_6502);
xnor U9603 (N_9603,N_6853,N_6110);
nand U9604 (N_9604,N_6856,N_6330);
or U9605 (N_9605,N_7670,N_6109);
xor U9606 (N_9606,N_7134,N_6536);
nand U9607 (N_9607,N_7176,N_7777);
or U9608 (N_9608,N_7064,N_7786);
nand U9609 (N_9609,N_6446,N_7652);
and U9610 (N_9610,N_6715,N_7040);
nor U9611 (N_9611,N_6510,N_7774);
or U9612 (N_9612,N_6194,N_6996);
and U9613 (N_9613,N_7605,N_6866);
nand U9614 (N_9614,N_7829,N_7651);
or U9615 (N_9615,N_6256,N_6836);
xor U9616 (N_9616,N_6817,N_6497);
and U9617 (N_9617,N_6477,N_7184);
or U9618 (N_9618,N_7561,N_7786);
nand U9619 (N_9619,N_7687,N_7887);
nand U9620 (N_9620,N_7505,N_6800);
xor U9621 (N_9621,N_7210,N_7360);
and U9622 (N_9622,N_7588,N_7730);
and U9623 (N_9623,N_7648,N_6077);
or U9624 (N_9624,N_6144,N_6219);
nor U9625 (N_9625,N_7264,N_7197);
nor U9626 (N_9626,N_7334,N_7479);
nand U9627 (N_9627,N_6627,N_7823);
nand U9628 (N_9628,N_6970,N_6318);
nor U9629 (N_9629,N_7137,N_7992);
and U9630 (N_9630,N_7247,N_6352);
xnor U9631 (N_9631,N_7974,N_7715);
nor U9632 (N_9632,N_7252,N_7940);
nand U9633 (N_9633,N_7611,N_6753);
xor U9634 (N_9634,N_7752,N_7765);
xor U9635 (N_9635,N_7423,N_6300);
or U9636 (N_9636,N_7185,N_6027);
or U9637 (N_9637,N_6274,N_7433);
nor U9638 (N_9638,N_6642,N_6298);
nand U9639 (N_9639,N_6019,N_6552);
xnor U9640 (N_9640,N_7683,N_6293);
xor U9641 (N_9641,N_6101,N_6918);
or U9642 (N_9642,N_6950,N_6774);
xnor U9643 (N_9643,N_7659,N_6329);
and U9644 (N_9644,N_7643,N_7119);
and U9645 (N_9645,N_7587,N_6329);
nor U9646 (N_9646,N_6604,N_6393);
or U9647 (N_9647,N_7049,N_6705);
nor U9648 (N_9648,N_6852,N_6519);
or U9649 (N_9649,N_7534,N_7998);
or U9650 (N_9650,N_6642,N_6606);
nor U9651 (N_9651,N_7983,N_6893);
xor U9652 (N_9652,N_6425,N_7365);
and U9653 (N_9653,N_7367,N_6106);
and U9654 (N_9654,N_6122,N_6327);
or U9655 (N_9655,N_6590,N_6242);
nand U9656 (N_9656,N_7064,N_6718);
or U9657 (N_9657,N_7258,N_6867);
nand U9658 (N_9658,N_6228,N_6206);
nand U9659 (N_9659,N_6748,N_6664);
and U9660 (N_9660,N_7472,N_7366);
xnor U9661 (N_9661,N_7552,N_6951);
xnor U9662 (N_9662,N_6637,N_6615);
xnor U9663 (N_9663,N_7677,N_7615);
or U9664 (N_9664,N_7091,N_6895);
xor U9665 (N_9665,N_6043,N_7760);
and U9666 (N_9666,N_6964,N_7865);
nand U9667 (N_9667,N_6680,N_6309);
nand U9668 (N_9668,N_6503,N_6600);
nor U9669 (N_9669,N_7027,N_7986);
nor U9670 (N_9670,N_6561,N_7467);
xnor U9671 (N_9671,N_7820,N_6582);
nor U9672 (N_9672,N_6778,N_7309);
and U9673 (N_9673,N_6666,N_7618);
nand U9674 (N_9674,N_7582,N_7650);
xor U9675 (N_9675,N_7616,N_6660);
xor U9676 (N_9676,N_7662,N_6059);
xor U9677 (N_9677,N_6113,N_6864);
xnor U9678 (N_9678,N_6591,N_7679);
or U9679 (N_9679,N_6720,N_7711);
nand U9680 (N_9680,N_6191,N_6013);
nand U9681 (N_9681,N_6712,N_7332);
xnor U9682 (N_9682,N_6612,N_7386);
and U9683 (N_9683,N_7335,N_7850);
xor U9684 (N_9684,N_6097,N_6215);
or U9685 (N_9685,N_6363,N_6995);
xnor U9686 (N_9686,N_7105,N_7129);
and U9687 (N_9687,N_7894,N_7133);
xnor U9688 (N_9688,N_7958,N_7613);
nand U9689 (N_9689,N_6671,N_6196);
or U9690 (N_9690,N_6164,N_7368);
nor U9691 (N_9691,N_7874,N_6103);
nor U9692 (N_9692,N_6857,N_7866);
or U9693 (N_9693,N_6432,N_6501);
nand U9694 (N_9694,N_7600,N_7876);
xor U9695 (N_9695,N_7099,N_7709);
or U9696 (N_9696,N_6967,N_7297);
nor U9697 (N_9697,N_7757,N_7455);
nor U9698 (N_9698,N_6506,N_7061);
nor U9699 (N_9699,N_7926,N_7902);
or U9700 (N_9700,N_6936,N_6265);
nor U9701 (N_9701,N_7147,N_6168);
or U9702 (N_9702,N_7675,N_6840);
nor U9703 (N_9703,N_7251,N_6863);
or U9704 (N_9704,N_6535,N_6460);
or U9705 (N_9705,N_6337,N_7183);
and U9706 (N_9706,N_6377,N_6242);
nor U9707 (N_9707,N_7604,N_7829);
and U9708 (N_9708,N_7727,N_7349);
nor U9709 (N_9709,N_7266,N_6406);
and U9710 (N_9710,N_7646,N_6803);
or U9711 (N_9711,N_7777,N_6173);
nand U9712 (N_9712,N_7394,N_7314);
and U9713 (N_9713,N_6800,N_6085);
or U9714 (N_9714,N_7897,N_7140);
xnor U9715 (N_9715,N_7294,N_7845);
xnor U9716 (N_9716,N_7482,N_7242);
xor U9717 (N_9717,N_7509,N_7826);
and U9718 (N_9718,N_6493,N_7126);
or U9719 (N_9719,N_7117,N_6757);
nand U9720 (N_9720,N_6593,N_7899);
nor U9721 (N_9721,N_6608,N_7666);
and U9722 (N_9722,N_7111,N_7956);
xor U9723 (N_9723,N_7277,N_6891);
and U9724 (N_9724,N_6108,N_7088);
and U9725 (N_9725,N_6307,N_6287);
nor U9726 (N_9726,N_6169,N_7275);
nand U9727 (N_9727,N_6398,N_6598);
nand U9728 (N_9728,N_6641,N_6024);
nor U9729 (N_9729,N_7676,N_6534);
or U9730 (N_9730,N_6576,N_7030);
nor U9731 (N_9731,N_7496,N_7922);
and U9732 (N_9732,N_7877,N_7654);
xor U9733 (N_9733,N_6842,N_6740);
nor U9734 (N_9734,N_6690,N_7917);
nand U9735 (N_9735,N_7659,N_7581);
and U9736 (N_9736,N_6174,N_6764);
nor U9737 (N_9737,N_7112,N_7373);
or U9738 (N_9738,N_7658,N_6149);
xnor U9739 (N_9739,N_7445,N_6762);
nand U9740 (N_9740,N_7180,N_7380);
nand U9741 (N_9741,N_7345,N_7873);
nor U9742 (N_9742,N_6595,N_6403);
or U9743 (N_9743,N_7367,N_6929);
nor U9744 (N_9744,N_7605,N_6464);
and U9745 (N_9745,N_6855,N_7382);
nand U9746 (N_9746,N_7610,N_6257);
or U9747 (N_9747,N_6578,N_7105);
nor U9748 (N_9748,N_6641,N_7991);
and U9749 (N_9749,N_6207,N_7720);
xor U9750 (N_9750,N_7826,N_6080);
and U9751 (N_9751,N_6102,N_6957);
or U9752 (N_9752,N_7239,N_6723);
and U9753 (N_9753,N_7253,N_6723);
xnor U9754 (N_9754,N_7718,N_7076);
nand U9755 (N_9755,N_7489,N_6117);
nand U9756 (N_9756,N_7031,N_7515);
xnor U9757 (N_9757,N_7159,N_6466);
and U9758 (N_9758,N_6643,N_6889);
nand U9759 (N_9759,N_7380,N_7466);
and U9760 (N_9760,N_7848,N_6902);
nor U9761 (N_9761,N_6341,N_6378);
or U9762 (N_9762,N_6356,N_6691);
xor U9763 (N_9763,N_7639,N_6809);
nand U9764 (N_9764,N_7724,N_7076);
nand U9765 (N_9765,N_7986,N_6891);
nand U9766 (N_9766,N_7458,N_7844);
nand U9767 (N_9767,N_6992,N_6248);
nand U9768 (N_9768,N_7990,N_7376);
or U9769 (N_9769,N_7666,N_7004);
and U9770 (N_9770,N_6953,N_7211);
xor U9771 (N_9771,N_6536,N_6565);
xor U9772 (N_9772,N_6385,N_7229);
and U9773 (N_9773,N_7628,N_7453);
and U9774 (N_9774,N_6482,N_6007);
nor U9775 (N_9775,N_6912,N_7481);
xnor U9776 (N_9776,N_6074,N_7071);
and U9777 (N_9777,N_7533,N_7262);
or U9778 (N_9778,N_7136,N_7245);
and U9779 (N_9779,N_6400,N_7887);
nand U9780 (N_9780,N_6324,N_7652);
and U9781 (N_9781,N_7832,N_7935);
xnor U9782 (N_9782,N_7635,N_6201);
xor U9783 (N_9783,N_6802,N_7319);
or U9784 (N_9784,N_6627,N_7842);
nor U9785 (N_9785,N_6888,N_6284);
nor U9786 (N_9786,N_6736,N_6893);
xnor U9787 (N_9787,N_7271,N_6688);
or U9788 (N_9788,N_7832,N_7970);
and U9789 (N_9789,N_7386,N_7082);
nor U9790 (N_9790,N_7104,N_7970);
and U9791 (N_9791,N_7968,N_6643);
nand U9792 (N_9792,N_7889,N_7714);
and U9793 (N_9793,N_6981,N_6680);
nand U9794 (N_9794,N_6209,N_6781);
nand U9795 (N_9795,N_6046,N_6761);
and U9796 (N_9796,N_6936,N_6193);
or U9797 (N_9797,N_7170,N_6084);
xor U9798 (N_9798,N_7793,N_7370);
or U9799 (N_9799,N_6700,N_6135);
nor U9800 (N_9800,N_6413,N_6520);
nor U9801 (N_9801,N_6344,N_6556);
and U9802 (N_9802,N_7573,N_7351);
nor U9803 (N_9803,N_6690,N_7032);
or U9804 (N_9804,N_7542,N_6346);
or U9805 (N_9805,N_7871,N_7253);
xnor U9806 (N_9806,N_7769,N_7612);
nor U9807 (N_9807,N_7683,N_6537);
or U9808 (N_9808,N_6124,N_6840);
xnor U9809 (N_9809,N_7335,N_6464);
nand U9810 (N_9810,N_7335,N_6623);
or U9811 (N_9811,N_6440,N_6867);
or U9812 (N_9812,N_7663,N_7855);
nand U9813 (N_9813,N_7979,N_7149);
nand U9814 (N_9814,N_7734,N_6555);
xor U9815 (N_9815,N_6863,N_6063);
xor U9816 (N_9816,N_7621,N_6193);
or U9817 (N_9817,N_7817,N_6372);
xnor U9818 (N_9818,N_6953,N_7712);
xor U9819 (N_9819,N_7022,N_6153);
nand U9820 (N_9820,N_6096,N_6062);
and U9821 (N_9821,N_7678,N_7648);
or U9822 (N_9822,N_6582,N_7838);
nand U9823 (N_9823,N_6063,N_6744);
nand U9824 (N_9824,N_7403,N_7599);
nor U9825 (N_9825,N_7723,N_6468);
and U9826 (N_9826,N_6042,N_6163);
xnor U9827 (N_9827,N_6988,N_7611);
or U9828 (N_9828,N_7149,N_7119);
and U9829 (N_9829,N_6006,N_7881);
xor U9830 (N_9830,N_6163,N_6714);
and U9831 (N_9831,N_6660,N_6953);
or U9832 (N_9832,N_6319,N_6547);
or U9833 (N_9833,N_7714,N_6039);
xnor U9834 (N_9834,N_6907,N_6448);
nand U9835 (N_9835,N_7577,N_6753);
nor U9836 (N_9836,N_6632,N_7491);
and U9837 (N_9837,N_7974,N_6349);
xor U9838 (N_9838,N_6454,N_7354);
xnor U9839 (N_9839,N_7843,N_6803);
xor U9840 (N_9840,N_6478,N_7258);
nor U9841 (N_9841,N_7677,N_6361);
nand U9842 (N_9842,N_7642,N_6007);
nand U9843 (N_9843,N_6421,N_6134);
nor U9844 (N_9844,N_6131,N_6600);
xor U9845 (N_9845,N_6093,N_6428);
nor U9846 (N_9846,N_6286,N_6145);
and U9847 (N_9847,N_7828,N_7982);
and U9848 (N_9848,N_6781,N_7421);
nor U9849 (N_9849,N_7531,N_6103);
nor U9850 (N_9850,N_6889,N_7695);
nor U9851 (N_9851,N_7421,N_7955);
nand U9852 (N_9852,N_7061,N_6322);
nand U9853 (N_9853,N_7312,N_6997);
nand U9854 (N_9854,N_6130,N_7104);
and U9855 (N_9855,N_6964,N_7139);
nand U9856 (N_9856,N_7002,N_6263);
nand U9857 (N_9857,N_6769,N_6494);
and U9858 (N_9858,N_7346,N_6484);
nor U9859 (N_9859,N_6762,N_7843);
and U9860 (N_9860,N_7114,N_6679);
xor U9861 (N_9861,N_7677,N_7904);
nand U9862 (N_9862,N_6367,N_7721);
xnor U9863 (N_9863,N_6454,N_6128);
nand U9864 (N_9864,N_7723,N_6804);
xor U9865 (N_9865,N_7168,N_6155);
and U9866 (N_9866,N_6028,N_6763);
nand U9867 (N_9867,N_7976,N_6066);
xnor U9868 (N_9868,N_6701,N_7404);
or U9869 (N_9869,N_7569,N_7710);
nor U9870 (N_9870,N_6356,N_7452);
nor U9871 (N_9871,N_7747,N_6525);
xor U9872 (N_9872,N_6056,N_6279);
or U9873 (N_9873,N_7414,N_6907);
and U9874 (N_9874,N_6550,N_6800);
nor U9875 (N_9875,N_6482,N_7417);
nor U9876 (N_9876,N_7986,N_6993);
and U9877 (N_9877,N_7177,N_7135);
nor U9878 (N_9878,N_7965,N_6563);
nor U9879 (N_9879,N_7101,N_6641);
xor U9880 (N_9880,N_6977,N_7262);
or U9881 (N_9881,N_6284,N_6647);
nand U9882 (N_9882,N_7424,N_6143);
or U9883 (N_9883,N_6084,N_6534);
nor U9884 (N_9884,N_7826,N_6119);
nor U9885 (N_9885,N_6805,N_7902);
or U9886 (N_9886,N_6176,N_6954);
nand U9887 (N_9887,N_6794,N_7692);
or U9888 (N_9888,N_7804,N_6605);
xnor U9889 (N_9889,N_6649,N_6792);
nor U9890 (N_9890,N_7147,N_6932);
and U9891 (N_9891,N_7642,N_6610);
xnor U9892 (N_9892,N_6052,N_7727);
xnor U9893 (N_9893,N_7900,N_6431);
nor U9894 (N_9894,N_7164,N_6852);
and U9895 (N_9895,N_6050,N_7724);
xnor U9896 (N_9896,N_6309,N_7332);
nand U9897 (N_9897,N_6790,N_6752);
and U9898 (N_9898,N_7559,N_7913);
nand U9899 (N_9899,N_7980,N_7754);
and U9900 (N_9900,N_6672,N_6549);
nor U9901 (N_9901,N_6955,N_6822);
xor U9902 (N_9902,N_7183,N_6485);
and U9903 (N_9903,N_6058,N_7771);
or U9904 (N_9904,N_6572,N_6452);
nor U9905 (N_9905,N_7899,N_7619);
xor U9906 (N_9906,N_6535,N_7941);
or U9907 (N_9907,N_6477,N_6172);
nand U9908 (N_9908,N_6895,N_6210);
and U9909 (N_9909,N_6513,N_6771);
nand U9910 (N_9910,N_6581,N_6771);
nor U9911 (N_9911,N_7176,N_6593);
nor U9912 (N_9912,N_6137,N_6551);
and U9913 (N_9913,N_6233,N_6877);
or U9914 (N_9914,N_7776,N_6970);
nand U9915 (N_9915,N_6828,N_6515);
xor U9916 (N_9916,N_6677,N_6622);
xnor U9917 (N_9917,N_6502,N_6712);
or U9918 (N_9918,N_7669,N_6540);
or U9919 (N_9919,N_7323,N_7782);
nor U9920 (N_9920,N_6489,N_6688);
and U9921 (N_9921,N_7986,N_6368);
nand U9922 (N_9922,N_7968,N_6793);
nor U9923 (N_9923,N_6718,N_7569);
or U9924 (N_9924,N_6995,N_6127);
xor U9925 (N_9925,N_6611,N_6363);
and U9926 (N_9926,N_6832,N_7662);
nor U9927 (N_9927,N_6188,N_6354);
nor U9928 (N_9928,N_6659,N_6495);
xor U9929 (N_9929,N_6668,N_6475);
nor U9930 (N_9930,N_6919,N_6942);
xor U9931 (N_9931,N_6181,N_6380);
xor U9932 (N_9932,N_7255,N_6773);
xor U9933 (N_9933,N_7580,N_6832);
xnor U9934 (N_9934,N_7883,N_7384);
or U9935 (N_9935,N_6930,N_7897);
xor U9936 (N_9936,N_6117,N_7683);
nand U9937 (N_9937,N_7512,N_7150);
nor U9938 (N_9938,N_7235,N_6859);
nor U9939 (N_9939,N_6712,N_6693);
nand U9940 (N_9940,N_7605,N_6519);
or U9941 (N_9941,N_7459,N_7244);
nor U9942 (N_9942,N_7211,N_7024);
nand U9943 (N_9943,N_7007,N_6177);
or U9944 (N_9944,N_6589,N_7217);
and U9945 (N_9945,N_6836,N_6443);
nor U9946 (N_9946,N_6918,N_7318);
nor U9947 (N_9947,N_7251,N_6248);
nor U9948 (N_9948,N_6057,N_7136);
nand U9949 (N_9949,N_7048,N_6749);
and U9950 (N_9950,N_7294,N_7373);
xor U9951 (N_9951,N_7958,N_6247);
xnor U9952 (N_9952,N_7547,N_7872);
and U9953 (N_9953,N_6049,N_6600);
nand U9954 (N_9954,N_6020,N_6583);
xor U9955 (N_9955,N_7140,N_6635);
nor U9956 (N_9956,N_7464,N_6483);
xor U9957 (N_9957,N_7650,N_6082);
nor U9958 (N_9958,N_7119,N_7986);
xor U9959 (N_9959,N_6672,N_7231);
nor U9960 (N_9960,N_6354,N_6433);
or U9961 (N_9961,N_6201,N_6174);
xor U9962 (N_9962,N_7115,N_7428);
xnor U9963 (N_9963,N_7921,N_7229);
or U9964 (N_9964,N_7885,N_6160);
xor U9965 (N_9965,N_6038,N_7835);
and U9966 (N_9966,N_7152,N_7680);
xnor U9967 (N_9967,N_7624,N_6427);
nor U9968 (N_9968,N_6241,N_7769);
xor U9969 (N_9969,N_7912,N_6516);
or U9970 (N_9970,N_6087,N_7170);
and U9971 (N_9971,N_6420,N_7530);
and U9972 (N_9972,N_7004,N_6876);
and U9973 (N_9973,N_6254,N_6486);
xnor U9974 (N_9974,N_6718,N_6060);
or U9975 (N_9975,N_6207,N_6817);
nand U9976 (N_9976,N_7021,N_6667);
or U9977 (N_9977,N_6006,N_7315);
or U9978 (N_9978,N_7027,N_7821);
xnor U9979 (N_9979,N_6849,N_6710);
or U9980 (N_9980,N_7637,N_7316);
xnor U9981 (N_9981,N_7300,N_7508);
or U9982 (N_9982,N_6141,N_6397);
xor U9983 (N_9983,N_7113,N_7092);
xnor U9984 (N_9984,N_7890,N_6498);
or U9985 (N_9985,N_6209,N_7102);
or U9986 (N_9986,N_7600,N_7456);
xnor U9987 (N_9987,N_6755,N_7756);
xnor U9988 (N_9988,N_7449,N_7548);
nor U9989 (N_9989,N_7952,N_7443);
nand U9990 (N_9990,N_6354,N_7254);
xnor U9991 (N_9991,N_6612,N_7410);
nor U9992 (N_9992,N_6381,N_7244);
nand U9993 (N_9993,N_6978,N_6575);
nand U9994 (N_9994,N_6645,N_7020);
xnor U9995 (N_9995,N_6102,N_6152);
xnor U9996 (N_9996,N_7509,N_6733);
nand U9997 (N_9997,N_6476,N_6091);
or U9998 (N_9998,N_7740,N_7704);
or U9999 (N_9999,N_6497,N_7437);
xor U10000 (N_10000,N_8768,N_8070);
xnor U10001 (N_10001,N_9879,N_9436);
or U10002 (N_10002,N_9834,N_8061);
or U10003 (N_10003,N_8605,N_9959);
and U10004 (N_10004,N_8232,N_8996);
and U10005 (N_10005,N_9745,N_8690);
xor U10006 (N_10006,N_8796,N_8699);
or U10007 (N_10007,N_8964,N_9375);
and U10008 (N_10008,N_9165,N_8506);
nor U10009 (N_10009,N_8733,N_9659);
nor U10010 (N_10010,N_9036,N_9923);
or U10011 (N_10011,N_9449,N_9593);
or U10012 (N_10012,N_8821,N_9685);
nor U10013 (N_10013,N_8755,N_9163);
xor U10014 (N_10014,N_9836,N_8106);
nor U10015 (N_10015,N_9204,N_9250);
nor U10016 (N_10016,N_9133,N_9722);
xnor U10017 (N_10017,N_9690,N_9422);
or U10018 (N_10018,N_9240,N_9962);
nor U10019 (N_10019,N_8771,N_8075);
nand U10020 (N_10020,N_8382,N_8154);
and U10021 (N_10021,N_9904,N_9976);
nor U10022 (N_10022,N_8785,N_9175);
and U10023 (N_10023,N_9852,N_9022);
xor U10024 (N_10024,N_9403,N_8218);
nor U10025 (N_10025,N_8470,N_9103);
xnor U10026 (N_10026,N_8802,N_9000);
or U10027 (N_10027,N_8359,N_9694);
nand U10028 (N_10028,N_9629,N_8011);
and U10029 (N_10029,N_9054,N_9990);
nand U10030 (N_10030,N_9660,N_8779);
or U10031 (N_10031,N_8186,N_9965);
and U10032 (N_10032,N_9993,N_8419);
or U10033 (N_10033,N_9913,N_9195);
nand U10034 (N_10034,N_9364,N_8930);
and U10035 (N_10035,N_8910,N_8621);
nor U10036 (N_10036,N_9193,N_9982);
or U10037 (N_10037,N_8150,N_9570);
xnor U10038 (N_10038,N_9490,N_9257);
nand U10039 (N_10039,N_9017,N_9277);
or U10040 (N_10040,N_9853,N_8087);
xnor U10041 (N_10041,N_8704,N_9046);
or U10042 (N_10042,N_8635,N_8761);
xnor U10043 (N_10043,N_8980,N_9543);
and U10044 (N_10044,N_8467,N_8185);
nand U10045 (N_10045,N_9316,N_8228);
or U10046 (N_10046,N_8289,N_8847);
nand U10047 (N_10047,N_9339,N_9485);
and U10048 (N_10048,N_8326,N_8101);
xnor U10049 (N_10049,N_9977,N_9329);
and U10050 (N_10050,N_9956,N_9874);
xor U10051 (N_10051,N_9237,N_8933);
and U10052 (N_10052,N_9898,N_9026);
or U10053 (N_10053,N_8532,N_8428);
xnor U10054 (N_10054,N_9641,N_8788);
or U10055 (N_10055,N_9002,N_9215);
or U10056 (N_10056,N_9730,N_9806);
nor U10057 (N_10057,N_8845,N_8808);
or U10058 (N_10058,N_9692,N_9625);
nand U10059 (N_10059,N_9394,N_9970);
or U10060 (N_10060,N_8753,N_9628);
or U10061 (N_10061,N_8444,N_8257);
xor U10062 (N_10062,N_8970,N_9553);
and U10063 (N_10063,N_8581,N_8663);
nand U10064 (N_10064,N_9247,N_8725);
and U10065 (N_10065,N_9424,N_8880);
nor U10066 (N_10066,N_9487,N_8311);
nor U10067 (N_10067,N_9212,N_8914);
and U10068 (N_10068,N_9604,N_8861);
or U10069 (N_10069,N_9259,N_8034);
or U10070 (N_10070,N_9537,N_8905);
xnor U10071 (N_10071,N_9646,N_8738);
nand U10072 (N_10072,N_8668,N_9087);
nor U10073 (N_10073,N_9912,N_8637);
and U10074 (N_10074,N_9887,N_8521);
and U10075 (N_10075,N_9102,N_8938);
nand U10076 (N_10076,N_9926,N_8054);
or U10077 (N_10077,N_8867,N_8869);
and U10078 (N_10078,N_9337,N_9010);
and U10079 (N_10079,N_8751,N_9832);
xnor U10080 (N_10080,N_9032,N_9297);
nor U10081 (N_10081,N_8091,N_9275);
xnor U10082 (N_10082,N_9450,N_9704);
and U10083 (N_10083,N_9776,N_8547);
nand U10084 (N_10084,N_9517,N_9914);
or U10085 (N_10085,N_9860,N_9458);
and U10086 (N_10086,N_9236,N_9334);
xor U10087 (N_10087,N_9154,N_9991);
and U10088 (N_10088,N_9968,N_8292);
nor U10089 (N_10089,N_8344,N_9476);
and U10090 (N_10090,N_9348,N_8098);
nand U10091 (N_10091,N_9547,N_9693);
and U10092 (N_10092,N_8037,N_9995);
nand U10093 (N_10093,N_8279,N_8610);
nand U10094 (N_10094,N_9443,N_9217);
and U10095 (N_10095,N_8891,N_9492);
nor U10096 (N_10096,N_9619,N_8315);
xnor U10097 (N_10097,N_9018,N_9453);
nand U10098 (N_10098,N_9078,N_8717);
and U10099 (N_10099,N_9858,N_9960);
nand U10100 (N_10100,N_8597,N_9183);
xnor U10101 (N_10101,N_9735,N_8531);
and U10102 (N_10102,N_9510,N_9774);
and U10103 (N_10103,N_9624,N_8670);
nand U10104 (N_10104,N_8440,N_9918);
nor U10105 (N_10105,N_9409,N_8058);
and U10106 (N_10106,N_8176,N_8081);
xnor U10107 (N_10107,N_9708,N_9939);
xor U10108 (N_10108,N_9686,N_8072);
and U10109 (N_10109,N_8269,N_8687);
and U10110 (N_10110,N_9650,N_9354);
nor U10111 (N_10111,N_8692,N_9131);
or U10112 (N_10112,N_8060,N_9601);
xor U10113 (N_10113,N_9588,N_8373);
nand U10114 (N_10114,N_9933,N_8653);
or U10115 (N_10115,N_8607,N_9023);
nand U10116 (N_10116,N_8741,N_9664);
and U10117 (N_10117,N_9260,N_9321);
or U10118 (N_10118,N_9179,N_9115);
nor U10119 (N_10119,N_8294,N_9727);
and U10120 (N_10120,N_8418,N_8332);
or U10121 (N_10121,N_8795,N_8994);
or U10122 (N_10122,N_8556,N_8857);
or U10123 (N_10123,N_9372,N_8212);
and U10124 (N_10124,N_8416,N_8873);
or U10125 (N_10125,N_8934,N_8633);
nor U10126 (N_10126,N_9987,N_9396);
xnor U10127 (N_10127,N_9572,N_8383);
nand U10128 (N_10128,N_8133,N_9651);
and U10129 (N_10129,N_9435,N_8716);
nor U10130 (N_10130,N_9089,N_9592);
and U10131 (N_10131,N_9932,N_9839);
and U10132 (N_10132,N_8838,N_9800);
nand U10133 (N_10133,N_8609,N_9737);
nand U10134 (N_10134,N_8090,N_9139);
nor U10135 (N_10135,N_8507,N_9764);
nor U10136 (N_10136,N_9135,N_9438);
nand U10137 (N_10137,N_8756,N_8274);
xor U10138 (N_10138,N_9121,N_8837);
xnor U10139 (N_10139,N_8680,N_8846);
or U10140 (N_10140,N_8807,N_8196);
and U10141 (N_10141,N_8360,N_9966);
nand U10142 (N_10142,N_8799,N_8760);
nor U10143 (N_10143,N_8304,N_9526);
or U10144 (N_10144,N_9331,N_9917);
nand U10145 (N_10145,N_9057,N_8530);
and U10146 (N_10146,N_8153,N_9120);
and U10147 (N_10147,N_8801,N_9478);
nor U10148 (N_10148,N_8046,N_9752);
nand U10149 (N_10149,N_9811,N_9019);
xnor U10150 (N_10150,N_8365,N_9461);
nand U10151 (N_10151,N_8083,N_8248);
and U10152 (N_10152,N_8245,N_9793);
nor U10153 (N_10153,N_8131,N_9371);
nand U10154 (N_10154,N_9413,N_8517);
nor U10155 (N_10155,N_9091,N_8544);
nor U10156 (N_10156,N_8399,N_8481);
nor U10157 (N_10157,N_9299,N_9094);
or U10158 (N_10158,N_8225,N_9929);
nand U10159 (N_10159,N_9496,N_9431);
nand U10160 (N_10160,N_9227,N_8285);
xor U10161 (N_10161,N_9969,N_8335);
and U10162 (N_10162,N_9439,N_9361);
nor U10163 (N_10163,N_9639,N_9454);
xnor U10164 (N_10164,N_8975,N_9097);
and U10165 (N_10165,N_8527,N_8040);
nor U10166 (N_10166,N_8486,N_9278);
xnor U10167 (N_10167,N_9554,N_9666);
nand U10168 (N_10168,N_8921,N_9609);
nand U10169 (N_10169,N_8707,N_9981);
xnor U10170 (N_10170,N_9859,N_9840);
and U10171 (N_10171,N_9164,N_9480);
xor U10172 (N_10172,N_8255,N_8723);
or U10173 (N_10173,N_9290,N_9099);
nand U10174 (N_10174,N_9583,N_9368);
xnor U10175 (N_10175,N_9612,N_8791);
nand U10176 (N_10176,N_9908,N_8278);
or U10177 (N_10177,N_8667,N_8032);
xnor U10178 (N_10178,N_8631,N_8268);
or U10179 (N_10179,N_9238,N_9518);
nor U10180 (N_10180,N_8883,N_9497);
or U10181 (N_10181,N_9009,N_9079);
nand U10182 (N_10182,N_8906,N_9726);
or U10183 (N_10183,N_9746,N_8823);
nand U10184 (N_10184,N_9508,N_9614);
nor U10185 (N_10185,N_8282,N_8340);
nor U10186 (N_10186,N_8671,N_9446);
and U10187 (N_10187,N_8008,N_8525);
xor U10188 (N_10188,N_9479,N_8818);
nor U10189 (N_10189,N_8708,N_8949);
or U10190 (N_10190,N_9883,N_9491);
nor U10191 (N_10191,N_9167,N_8765);
nor U10192 (N_10192,N_9043,N_8743);
and U10193 (N_10193,N_9444,N_8432);
or U10194 (N_10194,N_8398,N_9066);
and U10195 (N_10195,N_8526,N_8446);
nor U10196 (N_10196,N_8678,N_8342);
nand U10197 (N_10197,N_8831,N_8998);
xor U10198 (N_10198,N_8264,N_9597);
or U10199 (N_10199,N_9129,N_8627);
or U10200 (N_10200,N_8497,N_9777);
nand U10201 (N_10201,N_9028,N_9613);
and U10202 (N_10202,N_9653,N_8135);
and U10203 (N_10203,N_9620,N_8961);
or U10204 (N_10204,N_8180,N_8164);
and U10205 (N_10205,N_8129,N_9642);
xnor U10206 (N_10206,N_9228,N_8580);
xor U10207 (N_10207,N_8728,N_9170);
xor U10208 (N_10208,N_8537,N_8896);
nand U10209 (N_10209,N_8959,N_9213);
xnor U10210 (N_10210,N_8149,N_9025);
and U10211 (N_10211,N_8660,N_8543);
xnor U10212 (N_10212,N_9332,N_9055);
nor U10213 (N_10213,N_9846,N_9723);
nor U10214 (N_10214,N_9804,N_8664);
xnor U10215 (N_10215,N_9447,N_9037);
and U10216 (N_10216,N_8026,N_8057);
or U10217 (N_10217,N_8734,N_8159);
or U10218 (N_10218,N_9781,N_8613);
and U10219 (N_10219,N_8510,N_9753);
or U10220 (N_10220,N_8381,N_8643);
or U10221 (N_10221,N_9562,N_9787);
or U10222 (N_10222,N_9468,N_9455);
xnor U10223 (N_10223,N_9732,N_9560);
xor U10224 (N_10224,N_9598,N_8448);
nand U10225 (N_10225,N_9638,N_8460);
xnor U10226 (N_10226,N_8015,N_9816);
nor U10227 (N_10227,N_9008,N_8296);
or U10228 (N_10228,N_8356,N_9633);
xnor U10229 (N_10229,N_8618,N_9313);
xor U10230 (N_10230,N_9113,N_8071);
or U10231 (N_10231,N_8115,N_8393);
nand U10232 (N_10232,N_8952,N_8059);
nor U10233 (N_10233,N_9505,N_9005);
nor U10234 (N_10234,N_8346,N_9684);
or U10235 (N_10235,N_9599,N_9239);
and U10236 (N_10236,N_9482,N_9280);
and U10237 (N_10237,N_8895,N_8038);
or U10238 (N_10238,N_8407,N_8236);
xnor U10239 (N_10239,N_9367,N_8983);
nand U10240 (N_10240,N_8216,N_9166);
and U10241 (N_10241,N_9876,N_9184);
and U10242 (N_10242,N_9922,N_9092);
nand U10243 (N_10243,N_9532,N_9397);
and U10244 (N_10244,N_9360,N_8794);
nand U10245 (N_10245,N_9825,N_8465);
nand U10246 (N_10246,N_8999,N_8447);
and U10247 (N_10247,N_8151,N_8960);
nand U10248 (N_10248,N_9739,N_8214);
nor U10249 (N_10249,N_8140,N_9952);
and U10250 (N_10250,N_9483,N_8554);
xor U10251 (N_10251,N_8834,N_9034);
nand U10252 (N_10252,N_9178,N_9390);
or U10253 (N_10253,N_8612,N_9622);
nand U10254 (N_10254,N_9682,N_9441);
and U10255 (N_10255,N_9581,N_9556);
nor U10256 (N_10256,N_8764,N_9665);
nand U10257 (N_10257,N_8806,N_9210);
nor U10258 (N_10258,N_8413,N_9500);
nor U10259 (N_10259,N_9181,N_8065);
or U10260 (N_10260,N_9862,N_8384);
xor U10261 (N_10261,N_9549,N_9267);
xnor U10262 (N_10262,N_8495,N_9644);
nor U10263 (N_10263,N_8191,N_8367);
xor U10264 (N_10264,N_9504,N_8334);
and U10265 (N_10265,N_9885,N_9366);
xnor U10266 (N_10266,N_8966,N_8193);
xor U10267 (N_10267,N_8265,N_9958);
nor U10268 (N_10268,N_8247,N_8155);
and U10269 (N_10269,N_8870,N_8804);
or U10270 (N_10270,N_9200,N_8957);
xnor U10271 (N_10271,N_8860,N_8024);
xor U10272 (N_10272,N_8144,N_9927);
or U10273 (N_10273,N_9370,N_8665);
nor U10274 (N_10274,N_9052,N_8809);
and U10275 (N_10275,N_8939,N_8752);
nand U10276 (N_10276,N_8173,N_9673);
nor U10277 (N_10277,N_9153,N_8235);
and U10278 (N_10278,N_8324,N_8479);
xor U10279 (N_10279,N_9743,N_9851);
or U10280 (N_10280,N_8887,N_9391);
or U10281 (N_10281,N_8001,N_8591);
or U10282 (N_10282,N_9616,N_9668);
nor U10283 (N_10283,N_8630,N_9437);
xnor U10284 (N_10284,N_9080,N_9663);
or U10285 (N_10285,N_9232,N_8230);
nand U10286 (N_10286,N_9871,N_8069);
nor U10287 (N_10287,N_8995,N_9320);
and U10288 (N_10288,N_9417,N_9911);
and U10289 (N_10289,N_8240,N_9314);
xor U10290 (N_10290,N_8586,N_9868);
xor U10291 (N_10291,N_9784,N_9655);
nor U10292 (N_10292,N_9070,N_9477);
and U10293 (N_10293,N_9930,N_8339);
and U10294 (N_10294,N_9670,N_9657);
nand U10295 (N_10295,N_8589,N_9798);
or U10296 (N_10296,N_9067,N_8199);
xor U10297 (N_10297,N_9039,N_8003);
or U10298 (N_10298,N_8063,N_8619);
nand U10299 (N_10299,N_8826,N_8392);
xor U10300 (N_10300,N_8498,N_9288);
or U10301 (N_10301,N_9654,N_8112);
nand U10302 (N_10302,N_8251,N_9740);
and U10303 (N_10303,N_9548,N_9276);
xor U10304 (N_10304,N_8829,N_9600);
nand U10305 (N_10305,N_8175,N_9835);
nor U10306 (N_10306,N_9919,N_8714);
xnor U10307 (N_10307,N_8014,N_8650);
or U10308 (N_10308,N_9219,N_8575);
and U10309 (N_10309,N_8572,N_9293);
xor U10310 (N_10310,N_8417,N_8878);
xnor U10311 (N_10311,N_9140,N_8594);
nand U10312 (N_10312,N_8574,N_9707);
nor U10313 (N_10313,N_8441,N_9738);
nand U10314 (N_10314,N_8721,N_9627);
or U10315 (N_10315,N_8951,N_9234);
xor U10316 (N_10316,N_8920,N_9187);
and U10317 (N_10317,N_9697,N_8390);
nor U10318 (N_10318,N_8863,N_8489);
and U10319 (N_10319,N_9233,N_9808);
xnor U10320 (N_10320,N_9744,N_8080);
nand U10321 (N_10321,N_9985,N_8555);
nor U10322 (N_10322,N_9263,N_9117);
nand U10323 (N_10323,N_9160,N_9757);
or U10324 (N_10324,N_8041,N_9950);
nand U10325 (N_10325,N_8512,N_9141);
xnor U10326 (N_10326,N_9235,N_8732);
or U10327 (N_10327,N_9821,N_9538);
nand U10328 (N_10328,N_8466,N_9452);
nand U10329 (N_10329,N_8227,N_9177);
and U10330 (N_10330,N_8234,N_9013);
nor U10331 (N_10331,N_8542,N_9778);
or U10332 (N_10332,N_9635,N_8852);
or U10333 (N_10333,N_9016,N_9829);
xnor U10334 (N_10334,N_8972,N_9395);
or U10335 (N_10335,N_8825,N_9512);
and U10336 (N_10336,N_9751,N_8726);
or U10337 (N_10337,N_9696,N_8992);
xnor U10338 (N_10338,N_9376,N_9782);
xnor U10339 (N_10339,N_8425,N_9486);
nand U10340 (N_10340,N_8253,N_8792);
nand U10341 (N_10341,N_9311,N_8188);
and U10342 (N_10342,N_9369,N_8520);
nand U10343 (N_10343,N_8669,N_8473);
or U10344 (N_10344,N_9405,N_9145);
or U10345 (N_10345,N_8888,N_9683);
nand U10346 (N_10346,N_8666,N_9856);
xor U10347 (N_10347,N_8443,N_8207);
or U10348 (N_10348,N_9291,N_9794);
xor U10349 (N_10349,N_9151,N_9729);
nand U10350 (N_10350,N_9414,N_9051);
nand U10351 (N_10351,N_9813,N_9564);
and U10352 (N_10352,N_8926,N_8408);
nand U10353 (N_10353,N_9185,N_8181);
xor U10354 (N_10354,N_8757,N_8864);
and U10355 (N_10355,N_9596,N_8267);
or U10356 (N_10356,N_9065,N_9587);
xnor U10357 (N_10357,N_8195,N_8431);
and U10358 (N_10358,N_8590,N_9035);
or U10359 (N_10359,N_8104,N_8222);
or U10360 (N_10360,N_9189,N_8701);
nor U10361 (N_10361,N_8929,N_8731);
nand U10362 (N_10362,N_9605,N_9652);
nor U10363 (N_10363,N_8099,N_8299);
and U10364 (N_10364,N_8436,N_9999);
or U10365 (N_10365,N_9569,N_8674);
xnor U10366 (N_10366,N_8522,N_9317);
nor U10367 (N_10367,N_8076,N_9946);
nor U10368 (N_10368,N_9105,N_8389);
nand U10369 (N_10369,N_9506,N_9042);
or U10370 (N_10370,N_9411,N_8501);
nand U10371 (N_10371,N_9779,N_8463);
or U10372 (N_10372,N_8657,N_9373);
and U10373 (N_10373,N_9473,N_9818);
nand U10374 (N_10374,N_8803,N_8620);
or U10375 (N_10375,N_8836,N_8318);
and U10376 (N_10376,N_8737,N_8711);
or U10377 (N_10377,N_9146,N_8048);
or U10378 (N_10378,N_9341,N_9632);
nand U10379 (N_10379,N_8096,N_9425);
nand U10380 (N_10380,N_8640,N_8491);
nor U10381 (N_10381,N_8215,N_9713);
xnor U10382 (N_10382,N_8100,N_8971);
nor U10383 (N_10383,N_8210,N_9585);
and U10384 (N_10384,N_8685,N_8366);
nor U10385 (N_10385,N_8056,N_8923);
xnor U10386 (N_10386,N_9756,N_8200);
and U10387 (N_10387,N_9662,N_8017);
nor U10388 (N_10388,N_8426,N_8897);
and U10389 (N_10389,N_8851,N_8976);
nor U10390 (N_10390,N_8492,N_8592);
nor U10391 (N_10391,N_9284,N_9229);
xnor U10392 (N_10392,N_9571,N_8258);
nand U10393 (N_10393,N_9083,N_8696);
and U10394 (N_10394,N_8524,N_8908);
or U10395 (N_10395,N_9617,N_9350);
nand U10396 (N_10396,N_9152,N_8156);
or U10397 (N_10397,N_8505,N_8508);
nor U10398 (N_10398,N_9566,N_8604);
xnor U10399 (N_10399,N_9792,N_9182);
and U10400 (N_10400,N_9827,N_9241);
nand U10401 (N_10401,N_8954,N_9509);
xor U10402 (N_10402,N_8277,N_9807);
xor U10403 (N_10403,N_8793,N_8546);
xor U10404 (N_10404,N_9706,N_9203);
xor U10405 (N_10405,N_9724,N_8509);
nand U10406 (N_10406,N_8774,N_9867);
nand U10407 (N_10407,N_8045,N_9503);
and U10408 (N_10408,N_8031,N_9081);
and U10409 (N_10409,N_8169,N_8325);
or U10410 (N_10410,N_9516,N_9637);
and U10411 (N_10411,N_9199,N_9897);
nor U10412 (N_10412,N_9671,N_9830);
xor U10413 (N_10413,N_8433,N_9649);
xnor U10414 (N_10414,N_9064,N_8239);
nand U10415 (N_10415,N_8455,N_9426);
and U10416 (N_10416,N_9700,N_8474);
nor U10417 (N_10417,N_8719,N_9389);
nand U10418 (N_10418,N_8749,N_8744);
xor U10419 (N_10419,N_9355,N_9429);
nor U10420 (N_10420,N_8357,N_9824);
and U10421 (N_10421,N_8217,N_8480);
and U10422 (N_10422,N_8535,N_8601);
xnor U10423 (N_10423,N_9901,N_8903);
xnor U10424 (N_10424,N_9661,N_9006);
or U10425 (N_10425,N_8437,N_8515);
nand U10426 (N_10426,N_9356,N_9298);
nor U10427 (N_10427,N_8892,N_9305);
nand U10428 (N_10428,N_9074,N_8623);
nand U10429 (N_10429,N_8167,N_8927);
nor U10430 (N_10430,N_9495,N_8379);
and U10431 (N_10431,N_8940,N_8567);
or U10432 (N_10432,N_8622,N_8879);
or U10433 (N_10433,N_9607,N_8783);
or U10434 (N_10434,N_9957,N_9399);
nand U10435 (N_10435,N_9838,N_8445);
or U10436 (N_10436,N_9961,N_9550);
nand U10437 (N_10437,N_8720,N_9269);
xor U10438 (N_10438,N_8588,N_9225);
xor U10439 (N_10439,N_9979,N_8835);
nor U10440 (N_10440,N_8904,N_8396);
nor U10441 (N_10441,N_9534,N_8848);
and U10442 (N_10442,N_8249,N_9150);
xnor U10443 (N_10443,N_9988,N_8261);
and U10444 (N_10444,N_8922,N_9699);
xor U10445 (N_10445,N_9725,N_9271);
and U10446 (N_10446,N_9983,N_9775);
nand U10447 (N_10447,N_9925,N_8308);
xor U10448 (N_10448,N_8937,N_9410);
nor U10449 (N_10449,N_8982,N_8137);
and U10450 (N_10450,N_8912,N_9942);
nor U10451 (N_10451,N_9168,N_8502);
and U10452 (N_10452,N_9875,N_9172);
and U10453 (N_10453,N_9645,N_8868);
xnor U10454 (N_10454,N_8010,N_9680);
nand U10455 (N_10455,N_9940,N_8706);
nor U10456 (N_10456,N_9902,N_9771);
xnor U10457 (N_10457,N_8615,N_9198);
nand U10458 (N_10458,N_8965,N_8602);
nor U10459 (N_10459,N_9760,N_9058);
or U10460 (N_10460,N_9507,N_8850);
and U10461 (N_10461,N_8241,N_8557);
xnor U10462 (N_10462,N_9462,N_9938);
nor U10463 (N_10463,N_9056,N_9432);
nor U10464 (N_10464,N_9815,N_8679);
and U10465 (N_10465,N_8184,N_8244);
nand U10466 (N_10466,N_9289,N_8288);
nand U10467 (N_10467,N_8715,N_8004);
nand U10468 (N_10468,N_9324,N_8351);
xor U10469 (N_10469,N_8727,N_9114);
nor U10470 (N_10470,N_9471,N_9796);
nand U10471 (N_10471,N_9124,N_9963);
nor U10472 (N_10472,N_9197,N_8276);
nor U10473 (N_10473,N_9786,N_9921);
or U10474 (N_10474,N_8259,N_9845);
nand U10475 (N_10475,N_8962,N_8088);
and U10476 (N_10476,N_8742,N_9501);
xnor U10477 (N_10477,N_8842,N_8682);
and U10478 (N_10478,N_9457,N_9591);
nand U10479 (N_10479,N_9423,N_9681);
or U10480 (N_10480,N_8559,N_8166);
nand U10481 (N_10481,N_9877,N_9279);
nor U10482 (N_10482,N_9679,N_9021);
xor U10483 (N_10483,N_9134,N_9270);
xor U10484 (N_10484,N_9944,N_8528);
or U10485 (N_10485,N_8499,N_9866);
xor U10486 (N_10486,N_8973,N_9935);
or U10487 (N_10487,N_8658,N_8673);
nor U10488 (N_10488,N_8798,N_9418);
xnor U10489 (N_10489,N_8513,N_9676);
nor U10490 (N_10490,N_8415,N_9116);
nor U10491 (N_10491,N_8608,N_8275);
nor U10492 (N_10492,N_9286,N_8121);
nor U10493 (N_10493,N_8931,N_8483);
or U10494 (N_10494,N_9865,N_8363);
and U10495 (N_10495,N_8073,N_9967);
or U10496 (N_10496,N_8206,N_8358);
xnor U10497 (N_10497,N_8958,N_8298);
nor U10498 (N_10498,N_8283,N_9630);
xnor U10499 (N_10499,N_8917,N_8012);
nor U10500 (N_10500,N_9173,N_9861);
or U10501 (N_10501,N_8691,N_9323);
nor U10502 (N_10502,N_8172,N_8503);
nor U10503 (N_10503,N_9015,N_9315);
or U10504 (N_10504,N_8077,N_8986);
or U10505 (N_10505,N_8617,N_9608);
xor U10506 (N_10506,N_8766,N_8313);
and U10507 (N_10507,N_9513,N_9978);
and U10508 (N_10508,N_9848,N_8577);
or U10509 (N_10509,N_9304,N_9767);
nand U10510 (N_10510,N_8238,N_8307);
nand U10511 (N_10511,N_8456,N_8700);
nor U10512 (N_10512,N_9736,N_8220);
and U10513 (N_10513,N_9850,N_9442);
xor U10514 (N_10514,N_8595,N_8411);
or U10515 (N_10515,N_8890,N_9325);
and U10516 (N_10516,N_8790,N_9949);
nor U10517 (N_10517,N_9849,N_9206);
nor U10518 (N_10518,N_8943,N_9750);
xnor U10519 (N_10519,N_8321,N_8082);
or U10520 (N_10520,N_8394,N_9205);
and U10521 (N_10521,N_8772,N_9906);
nor U10522 (N_10522,N_9169,N_8936);
or U10523 (N_10523,N_8147,N_8451);
and U10524 (N_10524,N_8093,N_9469);
and U10525 (N_10525,N_8472,N_9086);
nor U10526 (N_10526,N_9803,N_9493);
or U10527 (N_10527,N_8642,N_8518);
xor U10528 (N_10528,N_8143,N_9196);
or U10529 (N_10529,N_8600,N_9899);
and U10530 (N_10530,N_9053,N_9741);
nor U10531 (N_10531,N_9123,N_9085);
and U10532 (N_10532,N_9253,N_8141);
and U10533 (N_10533,N_9365,N_8585);
or U10534 (N_10534,N_8388,N_9201);
and U10535 (N_10535,N_8849,N_8049);
nand U10536 (N_10536,N_9675,N_8784);
and U10537 (N_10537,N_8712,N_8944);
or U10538 (N_10538,N_9243,N_9310);
nand U10539 (N_10539,N_9420,N_9326);
nand U10540 (N_10540,N_9770,N_8333);
xor U10541 (N_10541,N_9953,N_9698);
nor U10542 (N_10542,N_8881,N_8331);
xor U10543 (N_10543,N_8163,N_8578);
nor U10544 (N_10544,N_9451,N_9590);
xor U10545 (N_10545,N_8898,N_8409);
and U10546 (N_10546,N_8780,N_9111);
nor U10547 (N_10547,N_9256,N_8647);
nand U10548 (N_10548,N_8815,N_9156);
or U10549 (N_10549,N_8029,N_8387);
xnor U10550 (N_10550,N_9347,N_8945);
xor U10551 (N_10551,N_8858,N_9755);
xor U10552 (N_10552,N_8349,N_8649);
and U10553 (N_10553,N_9068,N_9359);
nand U10554 (N_10554,N_9194,N_9717);
nand U10555 (N_10555,N_8280,N_9656);
nor U10556 (N_10556,N_9520,N_8006);
xor U10557 (N_10557,N_8086,N_9272);
nor U10558 (N_10558,N_8187,N_9847);
and U10559 (N_10559,N_9309,N_9344);
and U10560 (N_10560,N_8770,N_8924);
and U10561 (N_10561,N_9448,N_9631);
nor U10562 (N_10562,N_8582,N_9514);
and U10563 (N_10563,N_9546,N_8052);
nor U10564 (N_10564,N_8735,N_9658);
xor U10565 (N_10565,N_8656,N_9208);
or U10566 (N_10566,N_8639,N_8400);
nand U10567 (N_10567,N_8092,N_9768);
nand U10568 (N_10568,N_8552,N_8859);
xnor U10569 (N_10569,N_8893,N_9882);
xor U10570 (N_10570,N_8564,N_9349);
and U10571 (N_10571,N_9301,N_8266);
and U10572 (N_10572,N_9951,N_9004);
xnor U10573 (N_10573,N_8533,N_8830);
nand U10574 (N_10574,N_9873,N_8989);
nand U10575 (N_10575,N_8224,N_9388);
or U10576 (N_10576,N_8571,N_8993);
and U10577 (N_10577,N_8616,N_8452);
xor U10578 (N_10578,N_8900,N_8102);
nor U10579 (N_10579,N_9430,N_9363);
nor U10580 (N_10580,N_9801,N_9383);
xnor U10581 (N_10581,N_8345,N_8301);
or U10582 (N_10582,N_8110,N_8205);
nor U10583 (N_10583,N_9033,N_9252);
nand U10584 (N_10584,N_9362,N_9997);
nor U10585 (N_10585,N_8877,N_9328);
or U10586 (N_10586,N_9720,N_9082);
or U10587 (N_10587,N_9254,N_8722);
or U10588 (N_10588,N_8781,N_9749);
nor U10589 (N_10589,N_9580,N_9440);
and U10590 (N_10590,N_8157,N_8984);
xnor U10591 (N_10591,N_8705,N_8841);
nand U10592 (N_10592,N_9467,N_9602);
nor U10593 (N_10593,N_9351,N_8271);
xor U10594 (N_10594,N_8569,N_9230);
nand U10595 (N_10595,N_8353,N_8907);
nor U10596 (N_10596,N_8762,N_9157);
and U10597 (N_10597,N_9207,N_8380);
or U10598 (N_10598,N_8855,N_8250);
nor U10599 (N_10599,N_9242,N_9176);
nand U10600 (N_10600,N_8684,N_8314);
and U10601 (N_10601,N_8464,N_8134);
xor U10602 (N_10602,N_9523,N_9947);
nor U10603 (N_10603,N_9907,N_8323);
xnor U10604 (N_10604,N_8758,N_9780);
or U10605 (N_10605,N_9382,N_9881);
or U10606 (N_10606,N_8688,N_8485);
nand U10607 (N_10607,N_9251,N_8988);
xnor U10608 (N_10608,N_9937,N_8634);
nand U10609 (N_10609,N_9460,N_9144);
or U10610 (N_10610,N_9626,N_8844);
and U10611 (N_10611,N_9828,N_9542);
or U10612 (N_10612,N_9529,N_9606);
xor U10613 (N_10613,N_9812,N_9007);
nand U10614 (N_10614,N_9011,N_9636);
nor U10615 (N_10615,N_9059,N_8606);
or U10616 (N_10616,N_8659,N_8773);
nand U10617 (N_10617,N_8085,N_8754);
and U10618 (N_10618,N_9531,N_8068);
nor U10619 (N_10619,N_9048,N_8391);
or U10620 (N_10620,N_9943,N_9790);
nor U10621 (N_10621,N_8461,N_8347);
xor U10622 (N_10622,N_8925,N_9728);
nand U10623 (N_10623,N_8127,N_8476);
nand U10624 (N_10624,N_9174,N_9889);
xor U10625 (N_10625,N_9702,N_8871);
or U10626 (N_10626,N_8745,N_8422);
nand U10627 (N_10627,N_8786,N_9202);
xor U10628 (N_10628,N_8405,N_9255);
xnor U10629 (N_10629,N_8062,N_9336);
nor U10630 (N_10630,N_8703,N_9406);
nor U10631 (N_10631,N_9319,N_8328);
or U10632 (N_10632,N_8401,N_8894);
nor U10633 (N_10633,N_9799,N_8435);
nor U10634 (N_10634,N_9511,N_9330);
nand U10635 (N_10635,N_9691,N_8231);
xor U10636 (N_10636,N_9470,N_8429);
or U10637 (N_10637,N_9061,N_8739);
and U10638 (N_10638,N_8337,N_8805);
nor U10639 (N_10639,N_8759,N_8968);
or U10640 (N_10640,N_8284,N_9719);
nor U10641 (N_10641,N_8675,N_8302);
or U10642 (N_10642,N_8570,N_8430);
xnor U10643 (N_10643,N_9714,N_9826);
nor U10644 (N_10644,N_8079,N_9648);
nand U10645 (N_10645,N_9248,N_8662);
or U10646 (N_10646,N_9262,N_8882);
and U10647 (N_10647,N_9345,N_8827);
nand U10648 (N_10648,N_9107,N_9119);
nor U10649 (N_10649,N_8097,N_8563);
and U10650 (N_10650,N_9100,N_9773);
or U10651 (N_10651,N_9421,N_9211);
nand U10652 (N_10652,N_9936,N_9924);
or U10653 (N_10653,N_8978,N_8018);
and U10654 (N_10654,N_8953,N_8950);
and U10655 (N_10655,N_8913,N_9073);
nand U10656 (N_10656,N_8022,N_9831);
xor U10657 (N_10657,N_8915,N_9191);
or U10658 (N_10658,N_9896,N_8475);
nor U10659 (N_10659,N_8661,N_9992);
and U10660 (N_10660,N_9783,N_8462);
and U10661 (N_10661,N_8516,N_9063);
nor U10662 (N_10662,N_8641,N_8587);
xnor U10663 (N_10663,N_9575,N_8854);
xor U10664 (N_10664,N_9687,N_9484);
xnor U10665 (N_10665,N_9731,N_8545);
and U10666 (N_10666,N_9433,N_8377);
xor U10667 (N_10667,N_8021,N_8254);
or U10668 (N_10668,N_8406,N_9891);
nor U10669 (N_10669,N_9306,N_9049);
xor U10670 (N_10670,N_9075,N_9335);
and U10671 (N_10671,N_8439,N_9577);
or U10672 (N_10672,N_9093,N_9069);
and U10673 (N_10673,N_9975,N_8044);
or U10674 (N_10674,N_8484,N_9147);
or U10675 (N_10675,N_8111,N_8122);
or U10676 (N_10676,N_9302,N_9584);
and U10677 (N_10677,N_8824,N_8094);
or U10678 (N_10678,N_9855,N_8372);
xor U10679 (N_10679,N_9711,N_9380);
or U10680 (N_10680,N_9809,N_9221);
nand U10681 (N_10681,N_8103,N_8107);
nor U10682 (N_10682,N_8074,N_8016);
xnor U10683 (N_10683,N_9088,N_9322);
and U10684 (N_10684,N_9888,N_9819);
xor U10685 (N_10685,N_8865,N_9029);
nor U10686 (N_10686,N_8487,N_8902);
and U10687 (N_10687,N_8202,N_9127);
nand U10688 (N_10688,N_8028,N_8260);
xnor U10689 (N_10689,N_8190,N_8330);
xnor U10690 (N_10690,N_8899,N_8534);
nand U10691 (N_10691,N_9945,N_8350);
nor U10692 (N_10692,N_8974,N_9558);
or U10693 (N_10693,N_8009,N_9281);
nand U10694 (N_10694,N_8991,N_9695);
nand U10695 (N_10695,N_9716,N_8948);
xor U10696 (N_10696,N_8730,N_9374);
or U10697 (N_10697,N_9986,N_9231);
xnor U10698 (N_10698,N_8599,N_9031);
or U10699 (N_10699,N_8946,N_9718);
nor U10700 (N_10700,N_9710,N_8775);
nand U10701 (N_10701,N_8192,N_8822);
nor U10702 (N_10702,N_8120,N_8209);
or U10703 (N_10703,N_8148,N_8593);
nand U10704 (N_10704,N_8303,N_8158);
and U10705 (N_10705,N_9072,N_8797);
nand U10706 (N_10706,N_9973,N_8125);
xor U10707 (N_10707,N_8477,N_9989);
xor U10708 (N_10708,N_8748,N_9869);
nand U10709 (N_10709,N_9712,N_8568);
xor U10710 (N_10710,N_8990,N_8584);
nand U10711 (N_10711,N_9109,N_9582);
nor U10712 (N_10712,N_8128,N_9101);
or U10713 (N_10713,N_8395,N_8320);
or U10714 (N_10714,N_8875,N_8449);
and U10715 (N_10715,N_8194,N_8306);
and U10716 (N_10716,N_8025,N_9535);
nor U10717 (N_10717,N_9721,N_8252);
xnor U10718 (N_10718,N_9474,N_8490);
and U10719 (N_10719,N_8402,N_9300);
nor U10720 (N_10720,N_9733,N_8471);
or U10721 (N_10721,N_9402,N_9296);
and U10722 (N_10722,N_9579,N_8197);
or U10723 (N_10723,N_8565,N_9878);
xor U10724 (N_10724,N_9766,N_8636);
nor U10725 (N_10725,N_8352,N_9038);
and U10726 (N_10726,N_9864,N_8262);
xnor U10727 (N_10727,N_8450,N_8229);
nand U10728 (N_10728,N_8204,N_9915);
or U10729 (N_10729,N_8124,N_8343);
nand U10730 (N_10730,N_8198,N_9138);
nor U10731 (N_10731,N_9903,N_8625);
or U10732 (N_10732,N_8290,N_8702);
and U10733 (N_10733,N_9338,N_8763);
xnor U10734 (N_10734,N_8105,N_8213);
nor U10735 (N_10735,N_9971,N_8309);
or U10736 (N_10736,N_8322,N_9162);
nor U10737 (N_10737,N_8541,N_9012);
xnor U10738 (N_10738,N_9024,N_8457);
nor U10739 (N_10739,N_8030,N_9761);
or U10740 (N_10740,N_9618,N_8560);
and U10741 (N_10741,N_8412,N_9343);
or U10742 (N_10742,N_9041,N_9561);
xor U10743 (N_10743,N_8272,N_8116);
nand U10744 (N_10744,N_9464,N_8853);
xor U10745 (N_10745,N_8182,N_8536);
nor U10746 (N_10746,N_8270,N_9295);
or U10747 (N_10747,N_9427,N_8139);
xnor U10748 (N_10748,N_9472,N_9994);
nor U10749 (N_10749,N_9084,N_8540);
xnor U10750 (N_10750,N_8312,N_9261);
or U10751 (N_10751,N_8548,N_8787);
nor U10752 (N_10752,N_9401,N_8740);
nand U10753 (N_10753,N_8812,N_8233);
and U10754 (N_10754,N_9465,N_9647);
nor U10755 (N_10755,N_9294,N_9841);
and U10756 (N_10756,N_8281,N_9216);
nand U10757 (N_10757,N_8942,N_9672);
nor U10758 (N_10758,N_9377,N_9171);
and U10759 (N_10759,N_9573,N_8603);
xor U10760 (N_10760,N_9122,N_9916);
nand U10761 (N_10761,N_8171,N_8713);
nor U10762 (N_10762,N_9705,N_8956);
nor U10763 (N_10763,N_9398,N_9905);
xor U10764 (N_10764,N_8697,N_8000);
nand U10765 (N_10765,N_9540,N_8504);
xnor U10766 (N_10766,N_9498,N_8042);
and U10767 (N_10767,N_8297,N_9245);
and U10768 (N_10768,N_8551,N_9734);
xnor U10769 (N_10769,N_8885,N_8468);
xnor U10770 (N_10770,N_9307,N_8237);
nor U10771 (N_10771,N_9096,N_9623);
nand U10772 (N_10772,N_9791,N_9090);
or U10773 (N_10773,N_8529,N_9400);
nand U10774 (N_10774,N_8397,N_8500);
xor U10775 (N_10775,N_8242,N_9844);
nand U10776 (N_10776,N_9747,N_9077);
or U10777 (N_10777,N_8496,N_8438);
nor U10778 (N_10778,N_9488,N_8810);
xnor U10779 (N_10779,N_9459,N_8420);
or U10780 (N_10780,N_8036,N_8138);
xor U10781 (N_10781,N_9226,N_8368);
nor U10782 (N_10782,N_8341,N_8628);
and U10783 (N_10783,N_9342,N_9062);
nor U10784 (N_10784,N_8626,N_9863);
nand U10785 (N_10785,N_8911,N_8047);
xnor U10786 (N_10786,N_9128,N_9837);
or U10787 (N_10787,N_8095,N_9567);
and U10788 (N_10788,N_8423,N_9785);
nand U10789 (N_10789,N_8813,N_9475);
or U10790 (N_10790,N_9428,N_8969);
nor U10791 (N_10791,N_9098,N_8614);
nand U10792 (N_10792,N_9308,N_8538);
or U10793 (N_10793,N_8375,N_9404);
nand U10794 (N_10794,N_8203,N_9353);
xnor U10795 (N_10795,N_8573,N_8549);
xor U10796 (N_10796,N_9810,N_8403);
and U10797 (N_10797,N_9759,N_9667);
nor U10798 (N_10798,N_8655,N_8364);
nor U10799 (N_10799,N_9980,N_8651);
nor U10800 (N_10800,N_9136,N_9378);
or U10801 (N_10801,N_9186,N_8055);
or U10802 (N_10802,N_8839,N_8039);
and U10803 (N_10803,N_9519,N_8488);
or U10804 (N_10804,N_8583,N_9246);
nand U10805 (N_10805,N_9340,N_9886);
nand U10806 (N_10806,N_9218,N_8689);
nand U10807 (N_10807,N_9762,N_8511);
and U10808 (N_10808,N_9358,N_8576);
nand U10809 (N_10809,N_9499,N_9110);
nor U10810 (N_10810,N_8729,N_8632);
and U10811 (N_10811,N_9273,N_9814);
nand U10812 (N_10812,N_8694,N_8424);
nand U10813 (N_10813,N_8305,N_9333);
or U10814 (N_10814,N_9594,N_8355);
xor U10815 (N_10815,N_8084,N_9494);
nand U10816 (N_10816,N_8109,N_8371);
nand U10817 (N_10817,N_9984,N_8114);
or U10818 (N_10818,N_8050,N_8310);
xor U10819 (N_10819,N_9407,N_8919);
or U10820 (N_10820,N_8550,N_8291);
nand U10821 (N_10821,N_9565,N_9589);
nor U10822 (N_10822,N_9106,N_8819);
xor U10823 (N_10823,N_9709,N_8002);
nor U10824 (N_10824,N_8007,N_8648);
xnor U10825 (N_10825,N_8300,N_9408);
and U10826 (N_10826,N_8750,N_8977);
nor U10827 (N_10827,N_9071,N_8005);
or U10828 (N_10828,N_9379,N_9689);
nor U10829 (N_10829,N_9703,N_9595);
nor U10830 (N_10830,N_8293,N_9327);
or U10831 (N_10831,N_9528,N_9223);
and U10832 (N_10832,N_9857,N_8833);
and U10833 (N_10833,N_9769,N_9112);
nor U10834 (N_10834,N_9895,N_9393);
xnor U10835 (N_10835,N_9892,N_9948);
nor U10836 (N_10836,N_9795,N_9920);
or U10837 (N_10837,N_8693,N_9674);
nor U10838 (N_10838,N_9155,N_9539);
nor U10839 (N_10839,N_8035,N_9972);
or U10840 (N_10840,N_8329,N_8404);
xnor U10841 (N_10841,N_8427,N_9880);
nand U10842 (N_10842,N_8033,N_8816);
xor U10843 (N_10843,N_9318,N_9765);
xor U10844 (N_10844,N_8889,N_8113);
nor U10845 (N_10845,N_9544,N_9563);
nand U10846 (N_10846,N_9014,N_8624);
nor U10847 (N_10847,N_9854,N_9149);
and U10848 (N_10848,N_8361,N_9264);
nor U10849 (N_10849,N_9557,N_9677);
and U10850 (N_10850,N_9634,N_9559);
and U10851 (N_10851,N_8672,N_8414);
and U10852 (N_10852,N_8168,N_9872);
and U10853 (N_10853,N_8918,N_8814);
xnor U10854 (N_10854,N_8828,N_8747);
and U10855 (N_10855,N_8295,N_9522);
or U10856 (N_10856,N_9541,N_9108);
nand U10857 (N_10857,N_8458,N_8362);
nor U10858 (N_10858,N_8469,N_8916);
and U10859 (N_10859,N_8767,N_8287);
nor U10860 (N_10860,N_9050,N_9412);
xnor U10861 (N_10861,N_9466,N_9249);
nand U10862 (N_10862,N_8638,N_8064);
nor U10863 (N_10863,N_8800,N_8776);
nor U10864 (N_10864,N_9931,N_8027);
nor U10865 (N_10865,N_8119,N_9220);
xnor U10866 (N_10866,N_8843,N_8023);
nor U10867 (N_10867,N_9287,N_9578);
nor U10868 (N_10868,N_8872,N_9533);
nor U10869 (N_10869,N_9044,N_8442);
and U10870 (N_10870,N_9434,N_9258);
xnor U10871 (N_10871,N_9386,N_8686);
and U10872 (N_10872,N_8170,N_9574);
nor U10873 (N_10873,N_9268,N_8645);
nand U10874 (N_10874,N_8327,N_9669);
and U10875 (N_10875,N_8683,N_9003);
nand U10876 (N_10876,N_8778,N_8317);
or U10877 (N_10877,N_9955,N_9282);
nand U10878 (N_10878,N_8598,N_9159);
nor U10879 (N_10879,N_9104,N_9481);
xor U10880 (N_10880,N_9047,N_8183);
xor U10881 (N_10881,N_8160,N_8263);
nor U10882 (N_10882,N_9974,N_8817);
xor U10883 (N_10883,N_8179,N_9463);
and U10884 (N_10884,N_9894,N_9678);
xor U10885 (N_10885,N_9244,N_9521);
and U10886 (N_10886,N_8862,N_9188);
or U10887 (N_10887,N_8840,N_9040);
and U10888 (N_10888,N_9802,N_8316);
or U10889 (N_10889,N_8053,N_9833);
or U10890 (N_10890,N_8219,N_8553);
nor U10891 (N_10891,N_9772,N_9283);
or U10892 (N_10892,N_9419,N_8126);
nand U10893 (N_10893,N_9615,N_8376);
xnor U10894 (N_10894,N_8676,N_8201);
nand U10895 (N_10895,N_8286,N_9214);
nand U10896 (N_10896,N_8243,N_8354);
xor U10897 (N_10897,N_8142,N_8928);
xor U10898 (N_10898,N_9551,N_8256);
nand U10899 (N_10899,N_9688,N_9842);
or U10900 (N_10900,N_8947,N_8777);
nand U10901 (N_10901,N_9909,N_8646);
or U10902 (N_10902,N_9893,N_8876);
nand U10903 (N_10903,N_9143,N_9964);
nor U10904 (N_10904,N_8177,N_9928);
or U10905 (N_10905,N_8374,N_8226);
and U10906 (N_10906,N_8386,N_9701);
and U10907 (N_10907,N_9118,N_8561);
nand U10908 (N_10908,N_9020,N_9076);
nand U10909 (N_10909,N_8019,N_9890);
xor U10910 (N_10910,N_9515,N_8493);
or U10911 (N_10911,N_8178,N_9027);
nor U10912 (N_10912,N_9346,N_8886);
and U10913 (N_10913,N_8108,N_9456);
and U10914 (N_10914,N_9555,N_9303);
nand U10915 (N_10915,N_9789,N_8558);
or U10916 (N_10916,N_8136,N_9357);
nand U10917 (N_10917,N_8695,N_8161);
nand U10918 (N_10918,N_9445,N_9820);
or U10919 (N_10919,N_8874,N_8596);
xnor U10920 (N_10920,N_8746,N_9552);
and U10921 (N_10921,N_9823,N_8677);
and U10922 (N_10922,N_9568,N_8043);
nor U10923 (N_10923,N_8724,N_9385);
xor U10924 (N_10924,N_8410,N_9640);
or U10925 (N_10925,N_8385,N_9742);
nor U10926 (N_10926,N_9158,N_9192);
and U10927 (N_10927,N_9610,N_9934);
xnor U10928 (N_10928,N_9996,N_9611);
or U10929 (N_10929,N_8579,N_9822);
nor U10930 (N_10930,N_8652,N_9312);
nor U10931 (N_10931,N_8820,N_8421);
xnor U10932 (N_10932,N_8981,N_9224);
nor U10933 (N_10933,N_8901,N_8152);
nand U10934 (N_10934,N_8709,N_8013);
or U10935 (N_10935,N_8478,N_9415);
or U10936 (N_10936,N_9222,N_8866);
nand U10937 (N_10937,N_8146,N_8519);
xnor U10938 (N_10938,N_9001,N_8979);
or U10939 (N_10939,N_8348,N_8020);
or U10940 (N_10940,N_9763,N_8123);
xor U10941 (N_10941,N_8130,N_9797);
nor U10942 (N_10942,N_9754,N_8165);
nor U10943 (N_10943,N_9137,N_8736);
nor U10944 (N_10944,N_8434,N_8319);
or U10945 (N_10945,N_9180,N_9060);
nand U10946 (N_10946,N_9545,N_8985);
nor U10947 (N_10947,N_8909,N_9758);
or U10948 (N_10948,N_9586,N_8459);
xnor U10949 (N_10949,N_8145,N_8789);
nor U10950 (N_10950,N_9530,N_8629);
nor U10951 (N_10951,N_9621,N_9954);
or U10952 (N_10952,N_9125,N_9817);
nor U10953 (N_10953,N_9266,N_8967);
xor U10954 (N_10954,N_8644,N_8189);
and U10955 (N_10955,N_8769,N_9142);
xnor U10956 (N_10956,N_8482,N_8067);
xnor U10957 (N_10957,N_8174,N_8514);
nand U10958 (N_10958,N_8955,N_8221);
nand U10959 (N_10959,N_8370,N_9265);
and U10960 (N_10960,N_9045,N_8566);
and U10961 (N_10961,N_8453,N_8963);
xnor U10962 (N_10962,N_9190,N_9502);
xnor U10963 (N_10963,N_8078,N_8832);
nor U10964 (N_10964,N_9748,N_9384);
or U10965 (N_10965,N_8941,N_8494);
nor U10966 (N_10966,N_8935,N_8884);
and U10967 (N_10967,N_8539,N_9132);
xnor U10968 (N_10968,N_8611,N_8932);
or U10969 (N_10969,N_8369,N_8273);
nand U10970 (N_10970,N_9910,N_8223);
or U10971 (N_10971,N_9030,N_9381);
nand U10972 (N_10972,N_8987,N_8454);
nor U10973 (N_10973,N_9524,N_9843);
and U10974 (N_10974,N_9900,N_8117);
xnor U10975 (N_10975,N_9643,N_9274);
or U10976 (N_10976,N_9576,N_9884);
or U10977 (N_10977,N_9527,N_8523);
nor U10978 (N_10978,N_9805,N_9525);
nor U10979 (N_10979,N_8208,N_8338);
xnor U10980 (N_10980,N_8118,N_8811);
and U10981 (N_10981,N_9126,N_8710);
or U10982 (N_10982,N_9130,N_9387);
nor U10983 (N_10983,N_8132,N_8681);
nor U10984 (N_10984,N_8162,N_8782);
xnor U10985 (N_10985,N_8066,N_9941);
nor U10986 (N_10986,N_9352,N_9998);
nand U10987 (N_10987,N_9148,N_8336);
nand U10988 (N_10988,N_9489,N_9416);
and U10989 (N_10989,N_9209,N_8698);
nand U10990 (N_10990,N_9095,N_8856);
and U10991 (N_10991,N_8089,N_8378);
nand U10992 (N_10992,N_8997,N_9161);
and U10993 (N_10993,N_9788,N_9715);
nor U10994 (N_10994,N_8051,N_9285);
and U10995 (N_10995,N_8718,N_9536);
or U10996 (N_10996,N_8211,N_9870);
xnor U10997 (N_10997,N_9603,N_9392);
or U10998 (N_10998,N_8562,N_9292);
xor U10999 (N_10999,N_8654,N_8246);
and U11000 (N_11000,N_9755,N_9863);
and U11001 (N_11001,N_8618,N_9248);
nor U11002 (N_11002,N_8828,N_8132);
or U11003 (N_11003,N_9126,N_9650);
nand U11004 (N_11004,N_8171,N_9399);
nand U11005 (N_11005,N_9337,N_8201);
xnor U11006 (N_11006,N_8869,N_8462);
nand U11007 (N_11007,N_8534,N_8561);
and U11008 (N_11008,N_8943,N_8870);
nand U11009 (N_11009,N_9607,N_8170);
nand U11010 (N_11010,N_9757,N_9607);
and U11011 (N_11011,N_9687,N_9173);
nor U11012 (N_11012,N_8010,N_9699);
or U11013 (N_11013,N_9888,N_9220);
or U11014 (N_11014,N_8096,N_9465);
xnor U11015 (N_11015,N_9967,N_8468);
nor U11016 (N_11016,N_8512,N_8926);
nor U11017 (N_11017,N_9559,N_8437);
nand U11018 (N_11018,N_9712,N_9046);
xnor U11019 (N_11019,N_9931,N_8351);
or U11020 (N_11020,N_9732,N_8350);
nand U11021 (N_11021,N_9187,N_8189);
nand U11022 (N_11022,N_8881,N_9603);
xnor U11023 (N_11023,N_8386,N_9915);
nor U11024 (N_11024,N_8102,N_8296);
xnor U11025 (N_11025,N_8925,N_8356);
xnor U11026 (N_11026,N_8109,N_8042);
xnor U11027 (N_11027,N_9098,N_9965);
xnor U11028 (N_11028,N_8981,N_9193);
nor U11029 (N_11029,N_8981,N_8141);
nor U11030 (N_11030,N_8745,N_9094);
xnor U11031 (N_11031,N_9481,N_8592);
nor U11032 (N_11032,N_8078,N_8169);
or U11033 (N_11033,N_9298,N_8613);
nand U11034 (N_11034,N_8375,N_8917);
nor U11035 (N_11035,N_8980,N_9695);
nor U11036 (N_11036,N_9245,N_9480);
nand U11037 (N_11037,N_9176,N_8625);
or U11038 (N_11038,N_9509,N_8397);
nand U11039 (N_11039,N_8815,N_8887);
or U11040 (N_11040,N_9007,N_8919);
xor U11041 (N_11041,N_8421,N_9582);
or U11042 (N_11042,N_9742,N_8412);
and U11043 (N_11043,N_9305,N_9439);
nor U11044 (N_11044,N_9124,N_8075);
nand U11045 (N_11045,N_8037,N_9162);
and U11046 (N_11046,N_9066,N_9279);
nand U11047 (N_11047,N_9939,N_8915);
or U11048 (N_11048,N_9164,N_9158);
or U11049 (N_11049,N_8522,N_9870);
and U11050 (N_11050,N_9061,N_9020);
and U11051 (N_11051,N_9119,N_9039);
nor U11052 (N_11052,N_8013,N_8706);
nor U11053 (N_11053,N_9865,N_9248);
nor U11054 (N_11054,N_9654,N_9504);
xor U11055 (N_11055,N_8930,N_8888);
or U11056 (N_11056,N_8297,N_8191);
xor U11057 (N_11057,N_8284,N_9248);
and U11058 (N_11058,N_9882,N_8278);
or U11059 (N_11059,N_8867,N_9837);
nor U11060 (N_11060,N_9434,N_9544);
xor U11061 (N_11061,N_9660,N_9990);
nor U11062 (N_11062,N_8265,N_9598);
nor U11063 (N_11063,N_8912,N_8020);
and U11064 (N_11064,N_8873,N_8024);
nor U11065 (N_11065,N_9676,N_8039);
and U11066 (N_11066,N_9093,N_9260);
and U11067 (N_11067,N_8101,N_9748);
nand U11068 (N_11068,N_9613,N_9265);
xor U11069 (N_11069,N_9263,N_9549);
xnor U11070 (N_11070,N_9357,N_9010);
nor U11071 (N_11071,N_8910,N_9962);
and U11072 (N_11072,N_8569,N_8562);
or U11073 (N_11073,N_8344,N_9967);
xor U11074 (N_11074,N_9399,N_8176);
nand U11075 (N_11075,N_8833,N_9411);
nor U11076 (N_11076,N_9052,N_8406);
nand U11077 (N_11077,N_9076,N_8969);
nor U11078 (N_11078,N_9307,N_8475);
and U11079 (N_11079,N_8337,N_9468);
and U11080 (N_11080,N_8175,N_8505);
or U11081 (N_11081,N_8931,N_9356);
nand U11082 (N_11082,N_9574,N_8173);
nand U11083 (N_11083,N_9819,N_8250);
xor U11084 (N_11084,N_8111,N_9282);
nor U11085 (N_11085,N_8373,N_8419);
nor U11086 (N_11086,N_9999,N_8191);
nor U11087 (N_11087,N_8447,N_8176);
nor U11088 (N_11088,N_8845,N_9359);
nand U11089 (N_11089,N_8486,N_8163);
xor U11090 (N_11090,N_8457,N_8556);
nor U11091 (N_11091,N_8856,N_8683);
and U11092 (N_11092,N_9783,N_8701);
nor U11093 (N_11093,N_9709,N_8397);
or U11094 (N_11094,N_9766,N_9209);
xor U11095 (N_11095,N_9439,N_8852);
or U11096 (N_11096,N_8910,N_9216);
nand U11097 (N_11097,N_9649,N_9909);
or U11098 (N_11098,N_8906,N_8532);
nand U11099 (N_11099,N_9171,N_8975);
nor U11100 (N_11100,N_8354,N_9769);
and U11101 (N_11101,N_9279,N_9963);
nor U11102 (N_11102,N_9627,N_8070);
nand U11103 (N_11103,N_8256,N_9806);
or U11104 (N_11104,N_9668,N_9265);
and U11105 (N_11105,N_9404,N_9959);
or U11106 (N_11106,N_8072,N_9561);
nand U11107 (N_11107,N_8719,N_9477);
xnor U11108 (N_11108,N_9137,N_8108);
nand U11109 (N_11109,N_9008,N_8004);
or U11110 (N_11110,N_8474,N_8075);
nor U11111 (N_11111,N_9688,N_8894);
nor U11112 (N_11112,N_8325,N_9279);
or U11113 (N_11113,N_8533,N_9760);
nor U11114 (N_11114,N_9973,N_8098);
nand U11115 (N_11115,N_8324,N_9983);
and U11116 (N_11116,N_8873,N_9813);
nand U11117 (N_11117,N_8486,N_8799);
xor U11118 (N_11118,N_9525,N_9911);
and U11119 (N_11119,N_8269,N_9610);
nor U11120 (N_11120,N_9961,N_9113);
xor U11121 (N_11121,N_8281,N_8398);
and U11122 (N_11122,N_9926,N_9371);
nand U11123 (N_11123,N_9071,N_9513);
xor U11124 (N_11124,N_9489,N_8146);
and U11125 (N_11125,N_9076,N_9490);
and U11126 (N_11126,N_9905,N_9863);
nand U11127 (N_11127,N_8074,N_8417);
xnor U11128 (N_11128,N_9803,N_9773);
xnor U11129 (N_11129,N_9423,N_9389);
or U11130 (N_11130,N_8982,N_9073);
nor U11131 (N_11131,N_8603,N_9135);
nand U11132 (N_11132,N_8367,N_9315);
and U11133 (N_11133,N_9664,N_9551);
and U11134 (N_11134,N_8057,N_8722);
nor U11135 (N_11135,N_8033,N_8424);
xnor U11136 (N_11136,N_9801,N_9989);
nand U11137 (N_11137,N_9227,N_8225);
or U11138 (N_11138,N_8920,N_8720);
nand U11139 (N_11139,N_9909,N_8467);
or U11140 (N_11140,N_8279,N_8406);
xor U11141 (N_11141,N_9119,N_8704);
nor U11142 (N_11142,N_9290,N_9134);
and U11143 (N_11143,N_9967,N_8068);
and U11144 (N_11144,N_9842,N_8520);
and U11145 (N_11145,N_8950,N_9080);
xnor U11146 (N_11146,N_8150,N_8803);
or U11147 (N_11147,N_8119,N_8676);
nand U11148 (N_11148,N_9337,N_8697);
and U11149 (N_11149,N_8090,N_9523);
xnor U11150 (N_11150,N_9059,N_8839);
and U11151 (N_11151,N_8706,N_8650);
or U11152 (N_11152,N_9969,N_8916);
xor U11153 (N_11153,N_9556,N_8989);
nand U11154 (N_11154,N_9122,N_8226);
nor U11155 (N_11155,N_9686,N_9446);
nor U11156 (N_11156,N_9461,N_8692);
or U11157 (N_11157,N_8374,N_9748);
nor U11158 (N_11158,N_8206,N_8642);
or U11159 (N_11159,N_9265,N_9634);
nor U11160 (N_11160,N_9412,N_8432);
nor U11161 (N_11161,N_8315,N_8658);
nor U11162 (N_11162,N_8560,N_8433);
nor U11163 (N_11163,N_8718,N_8169);
xor U11164 (N_11164,N_9362,N_8215);
or U11165 (N_11165,N_8958,N_9600);
nor U11166 (N_11166,N_8466,N_8112);
and U11167 (N_11167,N_9478,N_9597);
xnor U11168 (N_11168,N_8581,N_9231);
nand U11169 (N_11169,N_9866,N_9033);
and U11170 (N_11170,N_9828,N_8073);
and U11171 (N_11171,N_9089,N_9428);
nand U11172 (N_11172,N_8571,N_8496);
or U11173 (N_11173,N_8638,N_9636);
and U11174 (N_11174,N_9956,N_8287);
and U11175 (N_11175,N_9532,N_8751);
nor U11176 (N_11176,N_9382,N_8076);
or U11177 (N_11177,N_8172,N_8296);
and U11178 (N_11178,N_8177,N_9079);
and U11179 (N_11179,N_9767,N_9928);
nor U11180 (N_11180,N_8318,N_9833);
nand U11181 (N_11181,N_8703,N_8466);
xor U11182 (N_11182,N_8083,N_9028);
xnor U11183 (N_11183,N_9543,N_8333);
nand U11184 (N_11184,N_8012,N_9912);
nand U11185 (N_11185,N_9422,N_8155);
xor U11186 (N_11186,N_8780,N_9987);
or U11187 (N_11187,N_9384,N_9293);
nand U11188 (N_11188,N_9204,N_8634);
xor U11189 (N_11189,N_8816,N_9445);
nand U11190 (N_11190,N_9095,N_8794);
nand U11191 (N_11191,N_9118,N_9240);
nand U11192 (N_11192,N_8054,N_8076);
or U11193 (N_11193,N_9048,N_9500);
and U11194 (N_11194,N_8611,N_8418);
or U11195 (N_11195,N_9836,N_9402);
or U11196 (N_11196,N_9653,N_9854);
xnor U11197 (N_11197,N_9298,N_9976);
xnor U11198 (N_11198,N_9242,N_8291);
or U11199 (N_11199,N_8253,N_9238);
nor U11200 (N_11200,N_8131,N_8428);
and U11201 (N_11201,N_8993,N_8219);
or U11202 (N_11202,N_9044,N_8381);
nand U11203 (N_11203,N_9777,N_9290);
nor U11204 (N_11204,N_9166,N_8804);
xor U11205 (N_11205,N_9603,N_8464);
or U11206 (N_11206,N_8517,N_8936);
or U11207 (N_11207,N_8617,N_9594);
xor U11208 (N_11208,N_9068,N_9896);
or U11209 (N_11209,N_8809,N_8161);
nand U11210 (N_11210,N_9937,N_9744);
xnor U11211 (N_11211,N_9866,N_9929);
nor U11212 (N_11212,N_9473,N_8778);
xnor U11213 (N_11213,N_8386,N_9719);
xor U11214 (N_11214,N_8509,N_9391);
and U11215 (N_11215,N_8343,N_9415);
or U11216 (N_11216,N_8397,N_9243);
nand U11217 (N_11217,N_8177,N_9890);
or U11218 (N_11218,N_8802,N_9296);
and U11219 (N_11219,N_9800,N_8748);
nand U11220 (N_11220,N_8695,N_8095);
xnor U11221 (N_11221,N_8481,N_9675);
xnor U11222 (N_11222,N_9371,N_8595);
or U11223 (N_11223,N_8411,N_9918);
xnor U11224 (N_11224,N_8057,N_8337);
xnor U11225 (N_11225,N_8461,N_8610);
or U11226 (N_11226,N_9549,N_9827);
and U11227 (N_11227,N_8337,N_9203);
nor U11228 (N_11228,N_9340,N_9993);
nand U11229 (N_11229,N_8671,N_8780);
nor U11230 (N_11230,N_9959,N_9669);
nand U11231 (N_11231,N_9586,N_9966);
nand U11232 (N_11232,N_8939,N_8421);
and U11233 (N_11233,N_8205,N_8219);
or U11234 (N_11234,N_9099,N_8436);
and U11235 (N_11235,N_8090,N_8145);
nand U11236 (N_11236,N_8247,N_9537);
xnor U11237 (N_11237,N_9232,N_8481);
xnor U11238 (N_11238,N_8968,N_9891);
xnor U11239 (N_11239,N_8830,N_8825);
nor U11240 (N_11240,N_8197,N_8079);
and U11241 (N_11241,N_9518,N_9559);
nor U11242 (N_11242,N_8660,N_8355);
nand U11243 (N_11243,N_8285,N_8278);
or U11244 (N_11244,N_8722,N_8319);
and U11245 (N_11245,N_8481,N_8188);
and U11246 (N_11246,N_9062,N_8664);
nor U11247 (N_11247,N_9360,N_9488);
xnor U11248 (N_11248,N_8085,N_9970);
nor U11249 (N_11249,N_9218,N_8254);
nor U11250 (N_11250,N_9195,N_8727);
nand U11251 (N_11251,N_9666,N_9522);
nor U11252 (N_11252,N_9544,N_8716);
nor U11253 (N_11253,N_8934,N_8006);
or U11254 (N_11254,N_9690,N_8040);
and U11255 (N_11255,N_9642,N_9386);
nor U11256 (N_11256,N_8636,N_8089);
and U11257 (N_11257,N_8650,N_9006);
nand U11258 (N_11258,N_8027,N_8887);
nand U11259 (N_11259,N_8952,N_8106);
xnor U11260 (N_11260,N_9434,N_9194);
nand U11261 (N_11261,N_8712,N_9965);
xnor U11262 (N_11262,N_8091,N_8914);
nand U11263 (N_11263,N_9853,N_9652);
and U11264 (N_11264,N_9050,N_9553);
nor U11265 (N_11265,N_9409,N_9844);
and U11266 (N_11266,N_9058,N_9159);
nand U11267 (N_11267,N_9269,N_8194);
xor U11268 (N_11268,N_9889,N_9198);
xnor U11269 (N_11269,N_8308,N_8226);
xor U11270 (N_11270,N_8852,N_9975);
nor U11271 (N_11271,N_9210,N_9455);
nand U11272 (N_11272,N_8894,N_9095);
and U11273 (N_11273,N_9889,N_9030);
nand U11274 (N_11274,N_9221,N_9803);
and U11275 (N_11275,N_9865,N_8534);
or U11276 (N_11276,N_9235,N_9132);
and U11277 (N_11277,N_9145,N_8957);
and U11278 (N_11278,N_8118,N_8923);
and U11279 (N_11279,N_8097,N_8930);
or U11280 (N_11280,N_9592,N_9193);
xnor U11281 (N_11281,N_9035,N_9956);
xor U11282 (N_11282,N_8046,N_8865);
nor U11283 (N_11283,N_8942,N_9493);
xor U11284 (N_11284,N_8300,N_9690);
and U11285 (N_11285,N_8976,N_8839);
nand U11286 (N_11286,N_9500,N_9240);
xor U11287 (N_11287,N_9651,N_9057);
and U11288 (N_11288,N_8149,N_9703);
xor U11289 (N_11289,N_8151,N_8306);
nor U11290 (N_11290,N_9946,N_9107);
and U11291 (N_11291,N_9218,N_8701);
or U11292 (N_11292,N_9564,N_9003);
nor U11293 (N_11293,N_8201,N_8092);
nand U11294 (N_11294,N_9711,N_9644);
nor U11295 (N_11295,N_9975,N_9268);
xnor U11296 (N_11296,N_9854,N_9148);
nand U11297 (N_11297,N_9110,N_9422);
nand U11298 (N_11298,N_9293,N_9300);
and U11299 (N_11299,N_9181,N_9942);
xor U11300 (N_11300,N_9002,N_8374);
or U11301 (N_11301,N_9371,N_8047);
xor U11302 (N_11302,N_9820,N_8660);
nand U11303 (N_11303,N_9741,N_9029);
xor U11304 (N_11304,N_8935,N_8291);
nor U11305 (N_11305,N_8614,N_9018);
and U11306 (N_11306,N_8965,N_8198);
xor U11307 (N_11307,N_8069,N_9260);
or U11308 (N_11308,N_8333,N_9560);
nor U11309 (N_11309,N_9037,N_9404);
xor U11310 (N_11310,N_8256,N_8905);
or U11311 (N_11311,N_8151,N_8435);
and U11312 (N_11312,N_9782,N_9352);
nor U11313 (N_11313,N_9224,N_8596);
xnor U11314 (N_11314,N_8817,N_8783);
or U11315 (N_11315,N_8066,N_8341);
and U11316 (N_11316,N_9849,N_9249);
nor U11317 (N_11317,N_8391,N_8079);
or U11318 (N_11318,N_8685,N_9456);
nand U11319 (N_11319,N_8056,N_8524);
nand U11320 (N_11320,N_8119,N_8960);
and U11321 (N_11321,N_9132,N_8395);
nand U11322 (N_11322,N_8851,N_9950);
or U11323 (N_11323,N_8511,N_8442);
nor U11324 (N_11324,N_9511,N_8526);
and U11325 (N_11325,N_8185,N_8659);
nand U11326 (N_11326,N_8900,N_8780);
or U11327 (N_11327,N_9528,N_8979);
xor U11328 (N_11328,N_8377,N_9282);
nor U11329 (N_11329,N_8784,N_8185);
xnor U11330 (N_11330,N_8578,N_9429);
nand U11331 (N_11331,N_8909,N_8565);
and U11332 (N_11332,N_9542,N_9868);
nor U11333 (N_11333,N_8273,N_8315);
nand U11334 (N_11334,N_9364,N_8918);
nand U11335 (N_11335,N_9376,N_9726);
nor U11336 (N_11336,N_9157,N_9621);
and U11337 (N_11337,N_8819,N_8097);
xor U11338 (N_11338,N_8586,N_9672);
xor U11339 (N_11339,N_8562,N_8582);
or U11340 (N_11340,N_8476,N_8954);
nor U11341 (N_11341,N_8843,N_9504);
nor U11342 (N_11342,N_9267,N_8322);
or U11343 (N_11343,N_9009,N_9808);
or U11344 (N_11344,N_8607,N_8400);
nor U11345 (N_11345,N_9369,N_8743);
or U11346 (N_11346,N_8955,N_8654);
and U11347 (N_11347,N_9830,N_8161);
nor U11348 (N_11348,N_9436,N_9338);
xor U11349 (N_11349,N_9867,N_9485);
xor U11350 (N_11350,N_8834,N_8580);
nand U11351 (N_11351,N_8565,N_9109);
nor U11352 (N_11352,N_8525,N_9151);
nor U11353 (N_11353,N_9952,N_9626);
xor U11354 (N_11354,N_8135,N_8504);
xor U11355 (N_11355,N_8506,N_9283);
or U11356 (N_11356,N_9017,N_9907);
xnor U11357 (N_11357,N_9932,N_8731);
xor U11358 (N_11358,N_9063,N_9036);
or U11359 (N_11359,N_9797,N_9548);
or U11360 (N_11360,N_9393,N_9357);
or U11361 (N_11361,N_8086,N_9286);
xor U11362 (N_11362,N_9036,N_9566);
xor U11363 (N_11363,N_9458,N_8222);
xor U11364 (N_11364,N_9510,N_9377);
xnor U11365 (N_11365,N_8645,N_8981);
and U11366 (N_11366,N_9586,N_8520);
nor U11367 (N_11367,N_9514,N_8117);
xnor U11368 (N_11368,N_9479,N_8377);
or U11369 (N_11369,N_8188,N_9212);
xor U11370 (N_11370,N_9086,N_8707);
or U11371 (N_11371,N_8727,N_8556);
xnor U11372 (N_11372,N_9305,N_9986);
xor U11373 (N_11373,N_9928,N_8411);
and U11374 (N_11374,N_9311,N_9373);
nand U11375 (N_11375,N_9730,N_8459);
xnor U11376 (N_11376,N_9266,N_8289);
or U11377 (N_11377,N_8880,N_9035);
xnor U11378 (N_11378,N_8551,N_8029);
or U11379 (N_11379,N_8242,N_8881);
or U11380 (N_11380,N_8025,N_9158);
xnor U11381 (N_11381,N_9850,N_8795);
nor U11382 (N_11382,N_9299,N_9052);
nor U11383 (N_11383,N_9600,N_9963);
nor U11384 (N_11384,N_8903,N_9707);
xnor U11385 (N_11385,N_9115,N_8779);
nand U11386 (N_11386,N_9841,N_8089);
or U11387 (N_11387,N_8030,N_8607);
or U11388 (N_11388,N_8116,N_8593);
or U11389 (N_11389,N_8349,N_8241);
nor U11390 (N_11390,N_8106,N_9228);
and U11391 (N_11391,N_8998,N_8999);
xnor U11392 (N_11392,N_8829,N_9682);
or U11393 (N_11393,N_8180,N_9055);
and U11394 (N_11394,N_9816,N_8880);
or U11395 (N_11395,N_8342,N_8492);
nor U11396 (N_11396,N_9214,N_9118);
and U11397 (N_11397,N_9481,N_9484);
xor U11398 (N_11398,N_9921,N_9813);
or U11399 (N_11399,N_9697,N_8555);
and U11400 (N_11400,N_8465,N_8504);
nand U11401 (N_11401,N_8003,N_9145);
xnor U11402 (N_11402,N_8120,N_8028);
and U11403 (N_11403,N_8689,N_8717);
nor U11404 (N_11404,N_9122,N_8075);
xor U11405 (N_11405,N_9694,N_9933);
and U11406 (N_11406,N_9391,N_9619);
or U11407 (N_11407,N_8994,N_8749);
or U11408 (N_11408,N_8403,N_8675);
and U11409 (N_11409,N_9454,N_9676);
and U11410 (N_11410,N_9160,N_9303);
and U11411 (N_11411,N_9964,N_8864);
or U11412 (N_11412,N_8619,N_9924);
nand U11413 (N_11413,N_9409,N_9800);
and U11414 (N_11414,N_8633,N_9272);
or U11415 (N_11415,N_8802,N_8997);
or U11416 (N_11416,N_8097,N_9584);
xnor U11417 (N_11417,N_8844,N_8171);
nand U11418 (N_11418,N_8865,N_8482);
nor U11419 (N_11419,N_8587,N_8969);
or U11420 (N_11420,N_9815,N_8454);
or U11421 (N_11421,N_9761,N_9560);
and U11422 (N_11422,N_8521,N_9811);
xor U11423 (N_11423,N_8341,N_9291);
nand U11424 (N_11424,N_9210,N_9200);
nor U11425 (N_11425,N_8981,N_9452);
nand U11426 (N_11426,N_9723,N_8037);
nand U11427 (N_11427,N_8309,N_8081);
xnor U11428 (N_11428,N_9883,N_8006);
nand U11429 (N_11429,N_8308,N_9938);
nand U11430 (N_11430,N_8494,N_8609);
or U11431 (N_11431,N_9986,N_9517);
and U11432 (N_11432,N_8330,N_9620);
or U11433 (N_11433,N_9666,N_8625);
xnor U11434 (N_11434,N_8191,N_9132);
nand U11435 (N_11435,N_9509,N_9423);
nor U11436 (N_11436,N_8036,N_9175);
or U11437 (N_11437,N_8773,N_8969);
xnor U11438 (N_11438,N_9973,N_8438);
nor U11439 (N_11439,N_9588,N_8706);
nor U11440 (N_11440,N_9379,N_9834);
and U11441 (N_11441,N_9394,N_8230);
nor U11442 (N_11442,N_9672,N_8173);
nor U11443 (N_11443,N_9951,N_8619);
and U11444 (N_11444,N_9658,N_8775);
xnor U11445 (N_11445,N_8203,N_9268);
nand U11446 (N_11446,N_8362,N_9130);
or U11447 (N_11447,N_8407,N_9178);
nor U11448 (N_11448,N_8737,N_8561);
or U11449 (N_11449,N_9950,N_8768);
and U11450 (N_11450,N_8545,N_8779);
and U11451 (N_11451,N_8439,N_9508);
or U11452 (N_11452,N_8587,N_9919);
xor U11453 (N_11453,N_9251,N_8799);
nor U11454 (N_11454,N_8759,N_9157);
or U11455 (N_11455,N_9307,N_8231);
nand U11456 (N_11456,N_8358,N_9230);
nand U11457 (N_11457,N_9657,N_8844);
xnor U11458 (N_11458,N_8854,N_8178);
or U11459 (N_11459,N_8480,N_9890);
or U11460 (N_11460,N_8982,N_9894);
xor U11461 (N_11461,N_9497,N_8765);
xor U11462 (N_11462,N_8405,N_8721);
xnor U11463 (N_11463,N_9280,N_9424);
nor U11464 (N_11464,N_9629,N_9994);
nor U11465 (N_11465,N_8137,N_8450);
or U11466 (N_11466,N_9439,N_9507);
or U11467 (N_11467,N_9878,N_8277);
and U11468 (N_11468,N_9752,N_9142);
and U11469 (N_11469,N_8006,N_9866);
nand U11470 (N_11470,N_8068,N_9642);
and U11471 (N_11471,N_9416,N_8550);
nand U11472 (N_11472,N_9671,N_8832);
and U11473 (N_11473,N_8232,N_9778);
xor U11474 (N_11474,N_9996,N_8262);
nand U11475 (N_11475,N_9321,N_8051);
nor U11476 (N_11476,N_9786,N_8510);
xnor U11477 (N_11477,N_9583,N_8155);
nand U11478 (N_11478,N_8412,N_8815);
xor U11479 (N_11479,N_9506,N_8496);
and U11480 (N_11480,N_9052,N_9984);
and U11481 (N_11481,N_8165,N_9976);
or U11482 (N_11482,N_8410,N_9131);
and U11483 (N_11483,N_8386,N_8835);
nand U11484 (N_11484,N_9184,N_9520);
xor U11485 (N_11485,N_9444,N_9218);
xnor U11486 (N_11486,N_8609,N_8449);
nor U11487 (N_11487,N_9178,N_9728);
xor U11488 (N_11488,N_9611,N_8817);
xor U11489 (N_11489,N_9445,N_9884);
and U11490 (N_11490,N_9718,N_8148);
nand U11491 (N_11491,N_8690,N_8996);
and U11492 (N_11492,N_8999,N_9230);
or U11493 (N_11493,N_8086,N_9410);
nor U11494 (N_11494,N_8028,N_9738);
nor U11495 (N_11495,N_9174,N_9711);
or U11496 (N_11496,N_9269,N_9264);
and U11497 (N_11497,N_8875,N_8839);
and U11498 (N_11498,N_9387,N_8667);
xnor U11499 (N_11499,N_8587,N_9754);
nand U11500 (N_11500,N_8633,N_9975);
nor U11501 (N_11501,N_8719,N_8777);
or U11502 (N_11502,N_9989,N_8752);
nand U11503 (N_11503,N_9911,N_9563);
or U11504 (N_11504,N_8550,N_9736);
or U11505 (N_11505,N_9670,N_9918);
xor U11506 (N_11506,N_9735,N_8016);
and U11507 (N_11507,N_9175,N_8243);
nand U11508 (N_11508,N_9711,N_8246);
and U11509 (N_11509,N_9010,N_9681);
or U11510 (N_11510,N_8331,N_8833);
nor U11511 (N_11511,N_8117,N_9353);
or U11512 (N_11512,N_9186,N_8720);
nand U11513 (N_11513,N_9360,N_9007);
and U11514 (N_11514,N_9707,N_8517);
and U11515 (N_11515,N_8392,N_8137);
xor U11516 (N_11516,N_8311,N_9341);
nor U11517 (N_11517,N_9123,N_8053);
xnor U11518 (N_11518,N_9696,N_9978);
and U11519 (N_11519,N_9946,N_8377);
nor U11520 (N_11520,N_8545,N_9875);
or U11521 (N_11521,N_8358,N_8621);
or U11522 (N_11522,N_9949,N_8937);
nor U11523 (N_11523,N_8267,N_9752);
or U11524 (N_11524,N_9915,N_9792);
and U11525 (N_11525,N_8520,N_9950);
or U11526 (N_11526,N_9179,N_9172);
nand U11527 (N_11527,N_8075,N_8402);
nor U11528 (N_11528,N_8109,N_8323);
nand U11529 (N_11529,N_9745,N_9591);
and U11530 (N_11530,N_9894,N_8787);
and U11531 (N_11531,N_8321,N_8481);
or U11532 (N_11532,N_9020,N_9855);
nor U11533 (N_11533,N_9761,N_8327);
nor U11534 (N_11534,N_8526,N_9467);
xnor U11535 (N_11535,N_8142,N_8573);
and U11536 (N_11536,N_9591,N_8472);
and U11537 (N_11537,N_8018,N_9977);
and U11538 (N_11538,N_9638,N_8797);
xnor U11539 (N_11539,N_9035,N_9561);
or U11540 (N_11540,N_9240,N_9625);
and U11541 (N_11541,N_9856,N_9736);
and U11542 (N_11542,N_9712,N_8157);
nand U11543 (N_11543,N_9660,N_8305);
xor U11544 (N_11544,N_8477,N_9803);
nand U11545 (N_11545,N_9387,N_9956);
or U11546 (N_11546,N_9985,N_8003);
nand U11547 (N_11547,N_9350,N_8070);
nor U11548 (N_11548,N_8014,N_8207);
and U11549 (N_11549,N_8174,N_9721);
and U11550 (N_11550,N_8869,N_9465);
xnor U11551 (N_11551,N_9450,N_9934);
nand U11552 (N_11552,N_9396,N_8039);
nor U11553 (N_11553,N_9711,N_8506);
and U11554 (N_11554,N_8219,N_8487);
or U11555 (N_11555,N_9350,N_9030);
xor U11556 (N_11556,N_8568,N_9769);
xor U11557 (N_11557,N_9899,N_9910);
and U11558 (N_11558,N_8188,N_9455);
or U11559 (N_11559,N_9744,N_8349);
xnor U11560 (N_11560,N_8712,N_9722);
and U11561 (N_11561,N_9132,N_9895);
or U11562 (N_11562,N_8081,N_9671);
nand U11563 (N_11563,N_9131,N_8619);
nor U11564 (N_11564,N_8247,N_9776);
or U11565 (N_11565,N_9530,N_9209);
xnor U11566 (N_11566,N_9165,N_9105);
and U11567 (N_11567,N_8791,N_8710);
nor U11568 (N_11568,N_9072,N_8294);
nor U11569 (N_11569,N_9328,N_8170);
nand U11570 (N_11570,N_8027,N_9346);
xor U11571 (N_11571,N_8943,N_9959);
nand U11572 (N_11572,N_8575,N_8138);
or U11573 (N_11573,N_9318,N_9313);
or U11574 (N_11574,N_9981,N_9806);
xor U11575 (N_11575,N_8441,N_9362);
nor U11576 (N_11576,N_8940,N_9685);
nor U11577 (N_11577,N_9809,N_9185);
nor U11578 (N_11578,N_9572,N_8194);
or U11579 (N_11579,N_9270,N_9561);
nand U11580 (N_11580,N_9596,N_9414);
or U11581 (N_11581,N_9640,N_9858);
xnor U11582 (N_11582,N_8101,N_8764);
or U11583 (N_11583,N_9559,N_8166);
nand U11584 (N_11584,N_8127,N_8595);
and U11585 (N_11585,N_9735,N_8410);
and U11586 (N_11586,N_8956,N_8322);
nor U11587 (N_11587,N_9179,N_8599);
xor U11588 (N_11588,N_8946,N_8436);
or U11589 (N_11589,N_9663,N_8031);
or U11590 (N_11590,N_9418,N_9158);
nand U11591 (N_11591,N_9502,N_8762);
nor U11592 (N_11592,N_9369,N_9861);
nor U11593 (N_11593,N_8886,N_9386);
or U11594 (N_11594,N_9922,N_9171);
nand U11595 (N_11595,N_9259,N_9903);
xor U11596 (N_11596,N_9465,N_8314);
xnor U11597 (N_11597,N_9164,N_9905);
xnor U11598 (N_11598,N_9147,N_8045);
and U11599 (N_11599,N_8698,N_9289);
nor U11600 (N_11600,N_9894,N_9145);
or U11601 (N_11601,N_9913,N_9020);
nor U11602 (N_11602,N_9226,N_8506);
xor U11603 (N_11603,N_9537,N_9859);
nand U11604 (N_11604,N_8379,N_9938);
and U11605 (N_11605,N_9968,N_8853);
nand U11606 (N_11606,N_8840,N_8895);
xnor U11607 (N_11607,N_9205,N_8704);
xor U11608 (N_11608,N_9876,N_9882);
nor U11609 (N_11609,N_9641,N_8602);
nor U11610 (N_11610,N_8177,N_9218);
and U11611 (N_11611,N_9936,N_9051);
or U11612 (N_11612,N_8685,N_9417);
and U11613 (N_11613,N_8915,N_8354);
xnor U11614 (N_11614,N_8553,N_9610);
and U11615 (N_11615,N_8069,N_8368);
or U11616 (N_11616,N_8529,N_9518);
and U11617 (N_11617,N_8755,N_9178);
nand U11618 (N_11618,N_8716,N_9450);
nand U11619 (N_11619,N_9589,N_8003);
and U11620 (N_11620,N_8061,N_9885);
and U11621 (N_11621,N_9535,N_8280);
xnor U11622 (N_11622,N_9262,N_9711);
nor U11623 (N_11623,N_9196,N_8880);
xnor U11624 (N_11624,N_9854,N_8020);
or U11625 (N_11625,N_8174,N_9344);
or U11626 (N_11626,N_8342,N_9978);
nand U11627 (N_11627,N_8675,N_9242);
and U11628 (N_11628,N_9811,N_9096);
or U11629 (N_11629,N_9757,N_8787);
or U11630 (N_11630,N_8919,N_9986);
and U11631 (N_11631,N_8069,N_8093);
nand U11632 (N_11632,N_9950,N_9434);
or U11633 (N_11633,N_9881,N_8962);
nor U11634 (N_11634,N_8946,N_8642);
and U11635 (N_11635,N_8578,N_8177);
and U11636 (N_11636,N_8537,N_9620);
or U11637 (N_11637,N_9884,N_8567);
and U11638 (N_11638,N_8066,N_8310);
nand U11639 (N_11639,N_8024,N_9761);
xor U11640 (N_11640,N_8039,N_8464);
nor U11641 (N_11641,N_8602,N_8084);
and U11642 (N_11642,N_9835,N_9104);
and U11643 (N_11643,N_8366,N_8510);
nand U11644 (N_11644,N_9173,N_8181);
and U11645 (N_11645,N_8714,N_9055);
nand U11646 (N_11646,N_8040,N_8213);
xor U11647 (N_11647,N_8939,N_9657);
or U11648 (N_11648,N_8275,N_8027);
xor U11649 (N_11649,N_8878,N_9890);
nor U11650 (N_11650,N_9104,N_8749);
and U11651 (N_11651,N_8555,N_8946);
nand U11652 (N_11652,N_9760,N_9825);
or U11653 (N_11653,N_9968,N_9502);
nand U11654 (N_11654,N_8700,N_8735);
or U11655 (N_11655,N_9162,N_9415);
xor U11656 (N_11656,N_9404,N_9243);
and U11657 (N_11657,N_8186,N_9134);
xnor U11658 (N_11658,N_8488,N_9255);
or U11659 (N_11659,N_8787,N_9778);
and U11660 (N_11660,N_8548,N_9212);
and U11661 (N_11661,N_8112,N_9503);
nor U11662 (N_11662,N_8164,N_9971);
or U11663 (N_11663,N_8727,N_8764);
nand U11664 (N_11664,N_9049,N_8483);
or U11665 (N_11665,N_9073,N_8210);
nor U11666 (N_11666,N_8094,N_8735);
or U11667 (N_11667,N_8664,N_9803);
or U11668 (N_11668,N_9482,N_9838);
nand U11669 (N_11669,N_8152,N_9825);
and U11670 (N_11670,N_8457,N_8608);
nand U11671 (N_11671,N_9597,N_8953);
and U11672 (N_11672,N_9884,N_9928);
and U11673 (N_11673,N_8663,N_9476);
or U11674 (N_11674,N_8873,N_9026);
and U11675 (N_11675,N_8746,N_8433);
nor U11676 (N_11676,N_9347,N_9783);
xor U11677 (N_11677,N_8150,N_9948);
nor U11678 (N_11678,N_9659,N_9018);
and U11679 (N_11679,N_9825,N_8438);
xor U11680 (N_11680,N_9466,N_9213);
nor U11681 (N_11681,N_8355,N_8348);
xnor U11682 (N_11682,N_9846,N_8074);
xor U11683 (N_11683,N_9031,N_8606);
or U11684 (N_11684,N_9914,N_9778);
nor U11685 (N_11685,N_9251,N_8449);
and U11686 (N_11686,N_9665,N_9550);
and U11687 (N_11687,N_8903,N_8620);
and U11688 (N_11688,N_9533,N_8261);
nand U11689 (N_11689,N_8836,N_8855);
nand U11690 (N_11690,N_8333,N_8343);
or U11691 (N_11691,N_9331,N_9636);
nand U11692 (N_11692,N_8255,N_9081);
nor U11693 (N_11693,N_9850,N_9829);
xor U11694 (N_11694,N_8213,N_9327);
nor U11695 (N_11695,N_8468,N_9850);
and U11696 (N_11696,N_9119,N_9532);
nor U11697 (N_11697,N_9832,N_8415);
or U11698 (N_11698,N_8958,N_8801);
nor U11699 (N_11699,N_8813,N_9307);
or U11700 (N_11700,N_9504,N_9014);
nor U11701 (N_11701,N_8118,N_8837);
xnor U11702 (N_11702,N_8677,N_8968);
or U11703 (N_11703,N_9321,N_8347);
or U11704 (N_11704,N_9465,N_9858);
xnor U11705 (N_11705,N_8684,N_8324);
nand U11706 (N_11706,N_9805,N_8826);
and U11707 (N_11707,N_9582,N_8094);
and U11708 (N_11708,N_8582,N_9634);
or U11709 (N_11709,N_8387,N_8404);
nor U11710 (N_11710,N_8651,N_8063);
or U11711 (N_11711,N_9910,N_9254);
and U11712 (N_11712,N_9760,N_9377);
nor U11713 (N_11713,N_9026,N_9291);
nand U11714 (N_11714,N_8256,N_9066);
nand U11715 (N_11715,N_8464,N_9608);
nand U11716 (N_11716,N_9766,N_8892);
or U11717 (N_11717,N_9500,N_9637);
nand U11718 (N_11718,N_8180,N_9495);
and U11719 (N_11719,N_8941,N_8786);
xnor U11720 (N_11720,N_9267,N_9968);
nand U11721 (N_11721,N_9175,N_8366);
xnor U11722 (N_11722,N_9948,N_8738);
or U11723 (N_11723,N_8703,N_8454);
xnor U11724 (N_11724,N_9433,N_8253);
and U11725 (N_11725,N_9560,N_9523);
xnor U11726 (N_11726,N_9124,N_8133);
xor U11727 (N_11727,N_8080,N_9573);
or U11728 (N_11728,N_8498,N_9306);
nor U11729 (N_11729,N_8865,N_9055);
xor U11730 (N_11730,N_9935,N_9397);
xnor U11731 (N_11731,N_9705,N_9799);
xor U11732 (N_11732,N_8609,N_8948);
and U11733 (N_11733,N_9118,N_8834);
nand U11734 (N_11734,N_8432,N_8460);
nand U11735 (N_11735,N_8278,N_9845);
and U11736 (N_11736,N_9436,N_9570);
nand U11737 (N_11737,N_8099,N_9024);
nor U11738 (N_11738,N_8513,N_9580);
nand U11739 (N_11739,N_8831,N_8478);
nand U11740 (N_11740,N_8030,N_9079);
or U11741 (N_11741,N_9248,N_8023);
xnor U11742 (N_11742,N_9336,N_9101);
nor U11743 (N_11743,N_8965,N_8819);
and U11744 (N_11744,N_8791,N_8444);
or U11745 (N_11745,N_9333,N_8377);
and U11746 (N_11746,N_9261,N_8071);
nand U11747 (N_11747,N_9454,N_9256);
and U11748 (N_11748,N_8138,N_8509);
and U11749 (N_11749,N_9471,N_8039);
xnor U11750 (N_11750,N_9338,N_9448);
and U11751 (N_11751,N_8601,N_9425);
and U11752 (N_11752,N_9339,N_8655);
and U11753 (N_11753,N_8960,N_8044);
and U11754 (N_11754,N_9945,N_8649);
nand U11755 (N_11755,N_9995,N_9541);
and U11756 (N_11756,N_8451,N_8352);
nor U11757 (N_11757,N_8723,N_8217);
nand U11758 (N_11758,N_8109,N_8345);
nor U11759 (N_11759,N_8222,N_8021);
or U11760 (N_11760,N_9595,N_8297);
and U11761 (N_11761,N_8287,N_9006);
and U11762 (N_11762,N_9508,N_9126);
and U11763 (N_11763,N_9783,N_8134);
or U11764 (N_11764,N_8902,N_9089);
and U11765 (N_11765,N_9588,N_8066);
nand U11766 (N_11766,N_9323,N_9952);
nor U11767 (N_11767,N_8400,N_8796);
nor U11768 (N_11768,N_8762,N_9393);
and U11769 (N_11769,N_8115,N_9395);
nand U11770 (N_11770,N_9565,N_8862);
and U11771 (N_11771,N_9234,N_8765);
xnor U11772 (N_11772,N_8964,N_9435);
and U11773 (N_11773,N_9389,N_9397);
and U11774 (N_11774,N_8819,N_9489);
xnor U11775 (N_11775,N_8618,N_9978);
and U11776 (N_11776,N_8916,N_8255);
xor U11777 (N_11777,N_9127,N_8762);
and U11778 (N_11778,N_8140,N_8946);
or U11779 (N_11779,N_8085,N_9930);
xor U11780 (N_11780,N_8250,N_8453);
nand U11781 (N_11781,N_8664,N_8081);
and U11782 (N_11782,N_9125,N_8866);
nor U11783 (N_11783,N_8101,N_9907);
or U11784 (N_11784,N_9771,N_9045);
and U11785 (N_11785,N_8308,N_8033);
and U11786 (N_11786,N_8609,N_8893);
and U11787 (N_11787,N_8973,N_8829);
and U11788 (N_11788,N_9162,N_8231);
nand U11789 (N_11789,N_8862,N_8067);
and U11790 (N_11790,N_9605,N_9945);
xor U11791 (N_11791,N_9824,N_9198);
or U11792 (N_11792,N_8313,N_9048);
or U11793 (N_11793,N_8417,N_9709);
and U11794 (N_11794,N_9445,N_8977);
xor U11795 (N_11795,N_8177,N_9502);
and U11796 (N_11796,N_9483,N_8258);
xnor U11797 (N_11797,N_9666,N_9831);
nor U11798 (N_11798,N_9265,N_9339);
or U11799 (N_11799,N_9684,N_8436);
nand U11800 (N_11800,N_9760,N_9227);
xnor U11801 (N_11801,N_9263,N_9374);
and U11802 (N_11802,N_8901,N_9804);
nand U11803 (N_11803,N_9745,N_9751);
xor U11804 (N_11804,N_8037,N_9627);
nand U11805 (N_11805,N_8485,N_8150);
nand U11806 (N_11806,N_8043,N_9831);
xor U11807 (N_11807,N_8941,N_8100);
and U11808 (N_11808,N_9732,N_8317);
xor U11809 (N_11809,N_9073,N_8872);
and U11810 (N_11810,N_9255,N_9189);
and U11811 (N_11811,N_8645,N_8699);
nor U11812 (N_11812,N_8331,N_8551);
and U11813 (N_11813,N_9138,N_9080);
or U11814 (N_11814,N_8411,N_8131);
and U11815 (N_11815,N_8179,N_9673);
nor U11816 (N_11816,N_9693,N_9493);
and U11817 (N_11817,N_8992,N_8560);
or U11818 (N_11818,N_8571,N_8956);
nand U11819 (N_11819,N_8208,N_9346);
nand U11820 (N_11820,N_8938,N_8186);
or U11821 (N_11821,N_9367,N_9487);
and U11822 (N_11822,N_8288,N_9701);
nor U11823 (N_11823,N_8021,N_8305);
nand U11824 (N_11824,N_8689,N_8762);
xnor U11825 (N_11825,N_9702,N_8064);
xor U11826 (N_11826,N_8024,N_9407);
xor U11827 (N_11827,N_9380,N_9962);
and U11828 (N_11828,N_9515,N_9734);
xor U11829 (N_11829,N_9877,N_9958);
xnor U11830 (N_11830,N_9461,N_8341);
nor U11831 (N_11831,N_9920,N_8136);
nand U11832 (N_11832,N_8236,N_9424);
and U11833 (N_11833,N_9374,N_9220);
nor U11834 (N_11834,N_8704,N_8526);
xor U11835 (N_11835,N_8486,N_8171);
nand U11836 (N_11836,N_9790,N_9413);
or U11837 (N_11837,N_9484,N_8798);
xnor U11838 (N_11838,N_8614,N_9943);
xor U11839 (N_11839,N_9978,N_9662);
nand U11840 (N_11840,N_9143,N_9382);
nand U11841 (N_11841,N_8103,N_8628);
nand U11842 (N_11842,N_8311,N_8931);
nand U11843 (N_11843,N_9563,N_9195);
nor U11844 (N_11844,N_9192,N_8645);
xnor U11845 (N_11845,N_8609,N_9065);
nor U11846 (N_11846,N_9524,N_8636);
nand U11847 (N_11847,N_8681,N_9413);
nor U11848 (N_11848,N_8059,N_9967);
nor U11849 (N_11849,N_8767,N_8311);
and U11850 (N_11850,N_9074,N_9446);
nor U11851 (N_11851,N_9282,N_8618);
or U11852 (N_11852,N_8130,N_9121);
nor U11853 (N_11853,N_8826,N_9717);
nand U11854 (N_11854,N_8355,N_9808);
nand U11855 (N_11855,N_9500,N_8991);
nor U11856 (N_11856,N_8667,N_9570);
nor U11857 (N_11857,N_8696,N_8793);
xnor U11858 (N_11858,N_8578,N_8584);
nand U11859 (N_11859,N_8662,N_9706);
and U11860 (N_11860,N_9980,N_9433);
or U11861 (N_11861,N_9989,N_9505);
nor U11862 (N_11862,N_9550,N_8197);
or U11863 (N_11863,N_9055,N_9789);
nand U11864 (N_11864,N_9398,N_9022);
and U11865 (N_11865,N_8767,N_9385);
and U11866 (N_11866,N_8925,N_8045);
or U11867 (N_11867,N_8595,N_9718);
xor U11868 (N_11868,N_9521,N_8045);
or U11869 (N_11869,N_8512,N_9309);
and U11870 (N_11870,N_8540,N_9982);
nor U11871 (N_11871,N_9429,N_9904);
nor U11872 (N_11872,N_8286,N_9060);
nand U11873 (N_11873,N_9259,N_9178);
or U11874 (N_11874,N_8811,N_9237);
nor U11875 (N_11875,N_9421,N_9129);
and U11876 (N_11876,N_8437,N_9474);
xor U11877 (N_11877,N_9892,N_8546);
or U11878 (N_11878,N_9085,N_8751);
or U11879 (N_11879,N_8296,N_8748);
and U11880 (N_11880,N_8673,N_8651);
xnor U11881 (N_11881,N_9308,N_9638);
nand U11882 (N_11882,N_8848,N_9309);
nand U11883 (N_11883,N_9064,N_9118);
xnor U11884 (N_11884,N_8209,N_8825);
and U11885 (N_11885,N_8894,N_9847);
nor U11886 (N_11886,N_8055,N_8223);
nand U11887 (N_11887,N_9671,N_8754);
xnor U11888 (N_11888,N_9992,N_8172);
and U11889 (N_11889,N_8787,N_8583);
or U11890 (N_11890,N_8243,N_9502);
xnor U11891 (N_11891,N_8903,N_9895);
nor U11892 (N_11892,N_9098,N_8987);
xor U11893 (N_11893,N_8459,N_8336);
xor U11894 (N_11894,N_8167,N_9559);
xor U11895 (N_11895,N_8413,N_9701);
nand U11896 (N_11896,N_8377,N_8534);
nand U11897 (N_11897,N_8445,N_9877);
and U11898 (N_11898,N_8896,N_9826);
and U11899 (N_11899,N_8932,N_9429);
or U11900 (N_11900,N_8476,N_9711);
or U11901 (N_11901,N_8570,N_8874);
nand U11902 (N_11902,N_8044,N_8229);
nand U11903 (N_11903,N_9601,N_8015);
and U11904 (N_11904,N_8191,N_8536);
or U11905 (N_11905,N_8457,N_9600);
nor U11906 (N_11906,N_8127,N_9188);
nor U11907 (N_11907,N_8249,N_8723);
and U11908 (N_11908,N_9710,N_9137);
or U11909 (N_11909,N_9474,N_9608);
or U11910 (N_11910,N_8960,N_9915);
and U11911 (N_11911,N_9441,N_8205);
nand U11912 (N_11912,N_9515,N_8936);
or U11913 (N_11913,N_9792,N_8493);
nor U11914 (N_11914,N_9515,N_8902);
nand U11915 (N_11915,N_8590,N_8753);
or U11916 (N_11916,N_8259,N_9789);
and U11917 (N_11917,N_8373,N_9066);
and U11918 (N_11918,N_9215,N_9305);
nor U11919 (N_11919,N_8479,N_8086);
or U11920 (N_11920,N_9489,N_9486);
and U11921 (N_11921,N_8991,N_9581);
nand U11922 (N_11922,N_8624,N_9834);
nand U11923 (N_11923,N_9106,N_9912);
and U11924 (N_11924,N_8617,N_8620);
and U11925 (N_11925,N_9664,N_9295);
nor U11926 (N_11926,N_9811,N_8291);
nand U11927 (N_11927,N_9357,N_8387);
xnor U11928 (N_11928,N_8724,N_9230);
and U11929 (N_11929,N_9400,N_8550);
nor U11930 (N_11930,N_8929,N_8009);
nand U11931 (N_11931,N_8589,N_8415);
or U11932 (N_11932,N_9346,N_8345);
or U11933 (N_11933,N_8228,N_8278);
nor U11934 (N_11934,N_9702,N_9058);
and U11935 (N_11935,N_8156,N_9369);
nand U11936 (N_11936,N_9318,N_8485);
nand U11937 (N_11937,N_8031,N_9167);
and U11938 (N_11938,N_9360,N_9684);
nor U11939 (N_11939,N_9983,N_9715);
nor U11940 (N_11940,N_9792,N_8647);
and U11941 (N_11941,N_9146,N_9022);
xor U11942 (N_11942,N_8190,N_9298);
or U11943 (N_11943,N_9917,N_8237);
xor U11944 (N_11944,N_8687,N_9166);
or U11945 (N_11945,N_8815,N_9146);
and U11946 (N_11946,N_8044,N_8971);
nor U11947 (N_11947,N_8078,N_8802);
xor U11948 (N_11948,N_9553,N_9839);
xor U11949 (N_11949,N_8290,N_8199);
xor U11950 (N_11950,N_8923,N_9802);
nor U11951 (N_11951,N_8773,N_9256);
nor U11952 (N_11952,N_9069,N_8357);
nand U11953 (N_11953,N_8378,N_8165);
nand U11954 (N_11954,N_8076,N_9515);
nor U11955 (N_11955,N_9101,N_9064);
nor U11956 (N_11956,N_8171,N_9715);
or U11957 (N_11957,N_8326,N_8371);
nand U11958 (N_11958,N_9662,N_8101);
nand U11959 (N_11959,N_9139,N_9875);
xnor U11960 (N_11960,N_8961,N_8331);
or U11961 (N_11961,N_9350,N_8672);
and U11962 (N_11962,N_8974,N_9187);
nand U11963 (N_11963,N_9639,N_8685);
nor U11964 (N_11964,N_9729,N_9563);
and U11965 (N_11965,N_8438,N_8782);
nand U11966 (N_11966,N_8357,N_8420);
nor U11967 (N_11967,N_9103,N_9483);
nand U11968 (N_11968,N_8130,N_8234);
nand U11969 (N_11969,N_8133,N_9634);
xor U11970 (N_11970,N_9385,N_9455);
and U11971 (N_11971,N_9736,N_8830);
and U11972 (N_11972,N_8008,N_8789);
and U11973 (N_11973,N_9939,N_8385);
nor U11974 (N_11974,N_8841,N_9794);
and U11975 (N_11975,N_8546,N_9363);
nand U11976 (N_11976,N_8509,N_9677);
nor U11977 (N_11977,N_9351,N_9805);
xor U11978 (N_11978,N_9405,N_8451);
and U11979 (N_11979,N_9471,N_9655);
or U11980 (N_11980,N_8056,N_9845);
nand U11981 (N_11981,N_9306,N_9896);
nand U11982 (N_11982,N_9548,N_9467);
xor U11983 (N_11983,N_9681,N_8221);
nor U11984 (N_11984,N_8355,N_9590);
and U11985 (N_11985,N_9246,N_8763);
nand U11986 (N_11986,N_9291,N_8249);
and U11987 (N_11987,N_8908,N_8657);
xnor U11988 (N_11988,N_8686,N_8647);
xor U11989 (N_11989,N_8289,N_8756);
or U11990 (N_11990,N_8914,N_8970);
nand U11991 (N_11991,N_9731,N_9494);
or U11992 (N_11992,N_8946,N_8038);
nor U11993 (N_11993,N_9461,N_9118);
xnor U11994 (N_11994,N_8169,N_8306);
and U11995 (N_11995,N_8961,N_8426);
and U11996 (N_11996,N_9574,N_8989);
nand U11997 (N_11997,N_9245,N_8399);
or U11998 (N_11998,N_9263,N_8050);
nor U11999 (N_11999,N_8401,N_8530);
and U12000 (N_12000,N_11496,N_10121);
nand U12001 (N_12001,N_11017,N_10776);
and U12002 (N_12002,N_11736,N_10645);
or U12003 (N_12003,N_10949,N_11554);
nand U12004 (N_12004,N_10283,N_11688);
nand U12005 (N_12005,N_11150,N_10331);
and U12006 (N_12006,N_10246,N_10008);
xnor U12007 (N_12007,N_10365,N_10132);
nand U12008 (N_12008,N_11747,N_11205);
or U12009 (N_12009,N_10047,N_10168);
nor U12010 (N_12010,N_10934,N_10466);
xor U12011 (N_12011,N_10295,N_11035);
and U12012 (N_12012,N_11248,N_10455);
nand U12013 (N_12013,N_11225,N_11516);
nand U12014 (N_12014,N_10083,N_10723);
and U12015 (N_12015,N_10255,N_10686);
nor U12016 (N_12016,N_10948,N_11731);
or U12017 (N_12017,N_11710,N_10313);
and U12018 (N_12018,N_11379,N_11139);
or U12019 (N_12019,N_10933,N_10731);
nor U12020 (N_12020,N_11473,N_11758);
nor U12021 (N_12021,N_11675,N_11897);
xor U12022 (N_12022,N_10427,N_10034);
xor U12023 (N_12023,N_11174,N_11885);
xor U12024 (N_12024,N_11657,N_11370);
xnor U12025 (N_12025,N_11653,N_10183);
nor U12026 (N_12026,N_11495,N_11330);
and U12027 (N_12027,N_10995,N_10451);
or U12028 (N_12028,N_11314,N_10982);
nor U12029 (N_12029,N_11721,N_11494);
and U12030 (N_12030,N_10742,N_10227);
nand U12031 (N_12031,N_10738,N_11700);
and U12032 (N_12032,N_10299,N_11147);
or U12033 (N_12033,N_10517,N_11222);
nand U12034 (N_12034,N_10219,N_10072);
xnor U12035 (N_12035,N_10156,N_11451);
xor U12036 (N_12036,N_11179,N_11790);
and U12037 (N_12037,N_10878,N_11734);
nor U12038 (N_12038,N_10523,N_11566);
xor U12039 (N_12039,N_11301,N_11963);
nand U12040 (N_12040,N_11097,N_10813);
nand U12041 (N_12041,N_10476,N_11486);
xnor U12042 (N_12042,N_10820,N_11198);
and U12043 (N_12043,N_10358,N_10234);
nor U12044 (N_12044,N_11047,N_10847);
or U12045 (N_12045,N_10157,N_11601);
and U12046 (N_12046,N_10791,N_11841);
nand U12047 (N_12047,N_11580,N_10543);
nor U12048 (N_12048,N_11055,N_11338);
and U12049 (N_12049,N_11378,N_11285);
nor U12050 (N_12050,N_11238,N_11944);
nor U12051 (N_12051,N_10558,N_10929);
or U12052 (N_12052,N_10879,N_11218);
nand U12053 (N_12053,N_10470,N_11418);
or U12054 (N_12054,N_10081,N_11470);
nand U12055 (N_12055,N_10725,N_10074);
and U12056 (N_12056,N_10672,N_11712);
xnor U12057 (N_12057,N_11530,N_11114);
or U12058 (N_12058,N_10651,N_10733);
or U12059 (N_12059,N_10740,N_11864);
or U12060 (N_12060,N_10592,N_10479);
or U12061 (N_12061,N_11011,N_11899);
and U12062 (N_12062,N_11938,N_10010);
or U12063 (N_12063,N_11627,N_11837);
xor U12064 (N_12064,N_11973,N_11110);
xnor U12065 (N_12065,N_11412,N_11748);
xor U12066 (N_12066,N_10102,N_10556);
or U12067 (N_12067,N_10239,N_11089);
nor U12068 (N_12068,N_10508,N_11974);
nor U12069 (N_12069,N_10262,N_10411);
nor U12070 (N_12070,N_10642,N_10610);
and U12071 (N_12071,N_10320,N_11191);
and U12072 (N_12072,N_10636,N_11664);
nand U12073 (N_12073,N_10369,N_10175);
or U12074 (N_12074,N_10093,N_10668);
and U12075 (N_12075,N_11215,N_11127);
nand U12076 (N_12076,N_11927,N_10771);
xnor U12077 (N_12077,N_10352,N_10326);
nand U12078 (N_12078,N_11517,N_10000);
or U12079 (N_12079,N_11299,N_10045);
or U12080 (N_12080,N_11970,N_10433);
or U12081 (N_12081,N_11019,N_10419);
xnor U12082 (N_12082,N_10542,N_10106);
and U12083 (N_12083,N_10525,N_10452);
and U12084 (N_12084,N_11672,N_10113);
or U12085 (N_12085,N_11779,N_11087);
nand U12086 (N_12086,N_10026,N_11062);
nor U12087 (N_12087,N_10584,N_10531);
xor U12088 (N_12088,N_11625,N_10781);
nand U12089 (N_12089,N_10908,N_11702);
nor U12090 (N_12090,N_10648,N_10235);
nor U12091 (N_12091,N_10973,N_10565);
nand U12092 (N_12092,N_10893,N_10250);
and U12093 (N_12093,N_11171,N_11236);
or U12094 (N_12094,N_10504,N_11323);
nand U12095 (N_12095,N_11775,N_10602);
or U12096 (N_12096,N_10465,N_11667);
or U12097 (N_12097,N_10983,N_10752);
or U12098 (N_12098,N_10744,N_11784);
or U12099 (N_12099,N_10799,N_10915);
and U12100 (N_12100,N_11124,N_11083);
xor U12101 (N_12101,N_10817,N_11057);
nor U12102 (N_12102,N_10387,N_11768);
and U12103 (N_12103,N_11134,N_11297);
and U12104 (N_12104,N_11620,N_10085);
nand U12105 (N_12105,N_10244,N_11003);
and U12106 (N_12106,N_11827,N_10654);
xnor U12107 (N_12107,N_11777,N_10319);
xor U12108 (N_12108,N_10092,N_10344);
or U12109 (N_12109,N_11529,N_11234);
nand U12110 (N_12110,N_10756,N_11789);
nand U12111 (N_12111,N_10800,N_10539);
and U12112 (N_12112,N_11377,N_11628);
nor U12113 (N_12113,N_10345,N_11698);
or U12114 (N_12114,N_10545,N_11820);
and U12115 (N_12115,N_11293,N_11302);
or U12116 (N_12116,N_10335,N_11046);
xnor U12117 (N_12117,N_10696,N_11797);
xor U12118 (N_12118,N_10154,N_11891);
xnor U12119 (N_12119,N_11512,N_10328);
or U12120 (N_12120,N_10620,N_11051);
nand U12121 (N_12121,N_11884,N_11771);
and U12122 (N_12122,N_11984,N_10261);
and U12123 (N_12123,N_11261,N_10519);
nor U12124 (N_12124,N_11681,N_10056);
nor U12125 (N_12125,N_10841,N_10827);
or U12126 (N_12126,N_10152,N_10797);
or U12127 (N_12127,N_11332,N_11943);
or U12128 (N_12128,N_10371,N_10206);
xnor U12129 (N_12129,N_10058,N_10544);
nor U12130 (N_12130,N_11070,N_10515);
or U12131 (N_12131,N_11934,N_11611);
xnor U12132 (N_12132,N_11893,N_10861);
nand U12133 (N_12133,N_10057,N_10416);
nor U12134 (N_12134,N_10943,N_10643);
or U12135 (N_12135,N_10898,N_11983);
and U12136 (N_12136,N_10916,N_11699);
or U12137 (N_12137,N_10380,N_11277);
and U12138 (N_12138,N_11705,N_10571);
nand U12139 (N_12139,N_10919,N_10681);
or U12140 (N_12140,N_10198,N_11822);
xnor U12141 (N_12141,N_10376,N_11922);
nand U12142 (N_12142,N_10562,N_11869);
and U12143 (N_12143,N_11437,N_10670);
xor U12144 (N_12144,N_11313,N_11912);
nor U12145 (N_12145,N_10022,N_10133);
xnor U12146 (N_12146,N_11816,N_10798);
xor U12147 (N_12147,N_11276,N_11235);
and U12148 (N_12148,N_11880,N_10253);
and U12149 (N_12149,N_11388,N_11879);
or U12150 (N_12150,N_10862,N_10505);
xnor U12151 (N_12151,N_11868,N_10391);
and U12152 (N_12152,N_10128,N_10942);
or U12153 (N_12153,N_11108,N_10324);
xor U12154 (N_12154,N_10139,N_10086);
xnor U12155 (N_12155,N_10635,N_10432);
xnor U12156 (N_12156,N_10134,N_11803);
nand U12157 (N_12157,N_11872,N_11862);
nand U12158 (N_12158,N_10702,N_10502);
nor U12159 (N_12159,N_11630,N_11142);
nand U12160 (N_12160,N_11320,N_10518);
or U12161 (N_12161,N_11976,N_11654);
nand U12162 (N_12162,N_11077,N_11440);
and U12163 (N_12163,N_10378,N_11300);
and U12164 (N_12164,N_10209,N_10019);
and U12165 (N_12165,N_10413,N_11600);
and U12166 (N_12166,N_10900,N_11507);
nor U12167 (N_12167,N_10027,N_10207);
or U12168 (N_12168,N_11552,N_10099);
xor U12169 (N_12169,N_10520,N_10260);
nand U12170 (N_12170,N_11241,N_11761);
or U12171 (N_12171,N_11200,N_10578);
nor U12172 (N_12172,N_10596,N_10464);
and U12173 (N_12173,N_11204,N_10437);
and U12174 (N_12174,N_10016,N_10809);
nand U12175 (N_12175,N_11324,N_10698);
and U12176 (N_12176,N_11282,N_10035);
nand U12177 (N_12177,N_10541,N_11560);
xnor U12178 (N_12178,N_11279,N_11365);
nor U12179 (N_12179,N_11084,N_11123);
nor U12180 (N_12180,N_10223,N_11247);
nor U12181 (N_12181,N_10480,N_10341);
xor U12182 (N_12182,N_10783,N_10856);
and U12183 (N_12183,N_11564,N_10585);
nor U12184 (N_12184,N_11254,N_11481);
nand U12185 (N_12185,N_10888,N_10624);
and U12186 (N_12186,N_10422,N_10501);
xor U12187 (N_12187,N_10325,N_10766);
and U12188 (N_12188,N_10481,N_10489);
or U12189 (N_12189,N_10754,N_11082);
and U12190 (N_12190,N_11656,N_11099);
nor U12191 (N_12191,N_10037,N_11319);
xnor U12192 (N_12192,N_10986,N_10251);
xor U12193 (N_12193,N_11359,N_10751);
xnor U12194 (N_12194,N_10281,N_10876);
nand U12195 (N_12195,N_10402,N_10755);
xnor U12196 (N_12196,N_11619,N_11545);
xnor U12197 (N_12197,N_11304,N_10494);
or U12198 (N_12198,N_11170,N_11430);
nor U12199 (N_12199,N_10077,N_11343);
or U12200 (N_12200,N_11770,N_10843);
nor U12201 (N_12201,N_10023,N_10839);
and U12202 (N_12202,N_11211,N_11745);
or U12203 (N_12203,N_10289,N_11188);
nand U12204 (N_12204,N_10675,N_10445);
and U12205 (N_12205,N_10721,N_10231);
or U12206 (N_12206,N_10779,N_11358);
and U12207 (N_12207,N_10469,N_11068);
nor U12208 (N_12208,N_10393,N_11229);
nand U12209 (N_12209,N_11483,N_10184);
xnor U12210 (N_12210,N_11231,N_10478);
and U12211 (N_12211,N_11895,N_10832);
nor U12212 (N_12212,N_10745,N_10316);
nand U12213 (N_12213,N_10414,N_10288);
or U12214 (N_12214,N_11570,N_11383);
nand U12215 (N_12215,N_11535,N_11800);
nor U12216 (N_12216,N_10248,N_10739);
nor U12217 (N_12217,N_10887,N_11547);
and U12218 (N_12218,N_11206,N_10060);
and U12219 (N_12219,N_11067,N_10718);
nor U12220 (N_12220,N_10366,N_11273);
nand U12221 (N_12221,N_10905,N_11441);
or U12222 (N_12222,N_11726,N_11327);
xnor U12223 (N_12223,N_10979,N_11208);
xor U12224 (N_12224,N_10614,N_10155);
or U12225 (N_12225,N_10130,N_10397);
nor U12226 (N_12226,N_10275,N_11485);
nand U12227 (N_12227,N_10096,N_10497);
xnor U12228 (N_12228,N_10838,N_11531);
or U12229 (N_12229,N_10243,N_11998);
xnor U12230 (N_12230,N_10950,N_10138);
or U12231 (N_12231,N_11143,N_10191);
xnor U12232 (N_12232,N_11265,N_11130);
xor U12233 (N_12233,N_10323,N_10720);
or U12234 (N_12234,N_10103,N_11643);
nor U12235 (N_12235,N_10506,N_10753);
and U12236 (N_12236,N_11166,N_10978);
and U12237 (N_12237,N_11793,N_11366);
and U12238 (N_12238,N_10707,N_11116);
nor U12239 (N_12239,N_11344,N_10070);
and U12240 (N_12240,N_11730,N_11380);
nor U12241 (N_12241,N_10747,N_11281);
nor U12242 (N_12242,N_11972,N_10017);
nand U12243 (N_12243,N_10488,N_10549);
nor U12244 (N_12244,N_10974,N_10059);
xnor U12245 (N_12245,N_10492,N_10186);
nor U12246 (N_12246,N_10098,N_10994);
and U12247 (N_12247,N_10265,N_11598);
nor U12248 (N_12248,N_11095,N_11584);
xor U12249 (N_12249,N_10473,N_10100);
and U12250 (N_12250,N_11565,N_10105);
nor U12251 (N_12251,N_11334,N_10609);
and U12252 (N_12252,N_10457,N_11137);
nand U12253 (N_12253,N_10560,N_10435);
or U12254 (N_12254,N_11054,N_10914);
or U12255 (N_12255,N_11615,N_11802);
and U12256 (N_12256,N_10090,N_11508);
nor U12257 (N_12257,N_10200,N_11840);
nand U12258 (N_12258,N_11583,N_11394);
xor U12259 (N_12259,N_10342,N_11439);
and U12260 (N_12260,N_10412,N_10632);
or U12261 (N_12261,N_11053,N_11423);
nor U12262 (N_12262,N_10372,N_11932);
nor U12263 (N_12263,N_10811,N_11165);
xor U12264 (N_12264,N_10507,N_10247);
and U12265 (N_12265,N_10471,N_10762);
nand U12266 (N_12266,N_10171,N_10151);
or U12267 (N_12267,N_10068,N_10013);
nand U12268 (N_12268,N_10496,N_11772);
nor U12269 (N_12269,N_11157,N_10758);
nand U12270 (N_12270,N_11997,N_10415);
nor U12271 (N_12271,N_11275,N_11691);
nand U12272 (N_12272,N_10693,N_11420);
and U12273 (N_12273,N_11689,N_11367);
and U12274 (N_12274,N_11650,N_11538);
or U12275 (N_12275,N_11160,N_10095);
or U12276 (N_12276,N_11468,N_11262);
xor U12277 (N_12277,N_10237,N_11597);
nor U12278 (N_12278,N_11833,N_10303);
and U12279 (N_12279,N_10990,N_11574);
nor U12280 (N_12280,N_11638,N_11471);
nor U12281 (N_12281,N_11287,N_11969);
nor U12282 (N_12282,N_10462,N_11634);
or U12283 (N_12283,N_11350,N_11939);
nand U12284 (N_12284,N_11866,N_11957);
or U12285 (N_12285,N_10736,N_11582);
nand U12286 (N_12286,N_10947,N_11050);
nand U12287 (N_12287,N_10315,N_11295);
and U12288 (N_12288,N_10761,N_10317);
nand U12289 (N_12289,N_11227,N_10953);
xor U12290 (N_12290,N_10347,N_10939);
xor U12291 (N_12291,N_11284,N_10678);
or U12292 (N_12292,N_11318,N_11846);
nand U12293 (N_12293,N_11829,N_10835);
or U12294 (N_12294,N_11834,N_11852);
nand U12295 (N_12295,N_10576,N_11558);
nor U12296 (N_12296,N_11577,N_10423);
nand U12297 (N_12297,N_11467,N_10015);
or U12298 (N_12298,N_11990,N_10612);
nor U12299 (N_12299,N_10968,N_11203);
nand U12300 (N_12300,N_10004,N_11255);
xor U12301 (N_12301,N_10167,N_11416);
nand U12302 (N_12302,N_10854,N_11025);
xnor U12303 (N_12303,N_10886,N_11946);
and U12304 (N_12304,N_11106,N_10153);
or U12305 (N_12305,N_11080,N_11120);
and U12306 (N_12306,N_10824,N_10062);
nor U12307 (N_12307,N_11090,N_10927);
nand U12308 (N_12308,N_11931,N_10814);
nor U12309 (N_12309,N_11901,N_11052);
xor U12310 (N_12310,N_10012,N_11920);
or U12311 (N_12311,N_11523,N_10495);
xor U12312 (N_12312,N_11482,N_10181);
xor U12313 (N_12313,N_11493,N_11707);
and U12314 (N_12314,N_11626,N_10160);
and U12315 (N_12315,N_11743,N_10382);
and U12316 (N_12316,N_11609,N_10454);
nor U12317 (N_12317,N_10192,N_11991);
and U12318 (N_12318,N_10630,N_10601);
or U12319 (N_12319,N_10003,N_11075);
nand U12320 (N_12320,N_10212,N_11005);
nand U12321 (N_12321,N_11246,N_11873);
nor U12322 (N_12322,N_11823,N_10952);
nand U12323 (N_12323,N_10055,N_11417);
nor U12324 (N_12324,N_10821,N_11819);
and U12325 (N_12325,N_11477,N_10180);
and U12326 (N_12326,N_11103,N_11399);
nor U12327 (N_12327,N_10463,N_11724);
or U12328 (N_12328,N_10694,N_10374);
and U12329 (N_12329,N_11520,N_11867);
xnor U12330 (N_12330,N_10503,N_10407);
nor U12331 (N_12331,N_11753,N_11854);
or U12332 (N_12332,N_11043,N_10579);
nand U12333 (N_12333,N_11593,N_10373);
nor U12334 (N_12334,N_11904,N_11181);
nor U12335 (N_12335,N_10379,N_11333);
or U12336 (N_12336,N_10595,N_10390);
or U12337 (N_12337,N_11786,N_11469);
nand U12338 (N_12338,N_10785,N_10524);
and U12339 (N_12339,N_10395,N_10703);
nand U12340 (N_12340,N_10384,N_11817);
or U12341 (N_12341,N_11444,N_10748);
or U12342 (N_12342,N_10597,N_10906);
nand U12343 (N_12343,N_10605,N_10795);
or U12344 (N_12344,N_11413,N_10803);
nor U12345 (N_12345,N_10907,N_10705);
xor U12346 (N_12346,N_11875,N_11881);
nor U12347 (N_12347,N_10177,N_10587);
and U12348 (N_12348,N_10955,N_11385);
and U12349 (N_12349,N_11660,N_11402);
nand U12350 (N_12350,N_11812,N_11400);
nor U12351 (N_12351,N_11311,N_10129);
nand U12352 (N_12352,N_11038,N_10743);
xor U12353 (N_12353,N_11996,N_11453);
nand U12354 (N_12354,N_10339,N_10891);
xor U12355 (N_12355,N_11329,N_10400);
xor U12356 (N_12356,N_10730,N_11129);
xor U12357 (N_12357,N_10697,N_10306);
or U12358 (N_12358,N_11898,N_11941);
xnor U12359 (N_12359,N_10853,N_11924);
xor U12360 (N_12360,N_11141,N_10903);
or U12361 (N_12361,N_10930,N_10359);
nor U12362 (N_12362,N_11576,N_10849);
or U12363 (N_12363,N_10071,N_11253);
xor U12364 (N_12364,N_11387,N_11762);
or U12365 (N_12365,N_11550,N_11410);
nand U12366 (N_12366,N_10774,N_10552);
xor U12367 (N_12367,N_11785,N_11268);
xnor U12368 (N_12368,N_10759,N_11602);
and U12369 (N_12369,N_10162,N_11590);
xor U12370 (N_12370,N_10041,N_11733);
nand U12371 (N_12371,N_11781,N_11892);
xnor U12372 (N_12372,N_10161,N_11364);
nor U12373 (N_12373,N_11454,N_10428);
and U12374 (N_12374,N_11878,N_10144);
or U12375 (N_12375,N_10511,N_10176);
or U12376 (N_12376,N_11649,N_11940);
nand U12377 (N_12377,N_11795,N_11355);
nor U12378 (N_12378,N_11201,N_10540);
nor U12379 (N_12379,N_11925,N_11648);
and U12380 (N_12380,N_10336,N_11936);
nand U12381 (N_12381,N_11621,N_11543);
and U12382 (N_12382,N_10330,N_10954);
xor U12383 (N_12383,N_10691,N_11407);
nor U12384 (N_12384,N_11216,N_10591);
or U12385 (N_12385,N_10033,N_11573);
xnor U12386 (N_12386,N_11631,N_11419);
or U12387 (N_12387,N_10126,N_11349);
or U12388 (N_12388,N_10131,N_10700);
nor U12389 (N_12389,N_11286,N_10357);
nor U12390 (N_12390,N_10220,N_10305);
or U12391 (N_12391,N_11435,N_11040);
nor U12392 (N_12392,N_10362,N_10877);
or U12393 (N_12393,N_10810,N_11069);
nor U12394 (N_12394,N_11256,N_11985);
nand U12395 (N_12395,N_11168,N_11156);
nand U12396 (N_12396,N_10701,N_10166);
and U12397 (N_12397,N_10282,N_11118);
nor U12398 (N_12398,N_11346,N_10398);
nand U12399 (N_12399,N_10259,N_10992);
nand U12400 (N_12400,N_11890,N_11369);
or U12401 (N_12401,N_11677,N_11220);
and U12402 (N_12402,N_11128,N_10936);
and U12403 (N_12403,N_10286,N_10406);
xor U12404 (N_12404,N_10490,N_11223);
nor U12405 (N_12405,N_11684,N_11661);
or U12406 (N_12406,N_11680,N_11928);
nor U12407 (N_12407,N_10485,N_11371);
xnor U12408 (N_12408,N_10021,N_10439);
or U12409 (N_12409,N_11942,N_10680);
nand U12410 (N_12410,N_10536,N_10044);
nor U12411 (N_12411,N_10287,N_10815);
and U12412 (N_12412,N_11559,N_11161);
nand U12413 (N_12413,N_11632,N_10768);
or U12414 (N_12414,N_10859,N_10321);
and U12415 (N_12415,N_10882,N_10829);
xor U12416 (N_12416,N_10392,N_10493);
nor U12417 (N_12417,N_10637,N_10179);
nor U12418 (N_12418,N_11618,N_11339);
or U12419 (N_12419,N_10538,N_10770);
nor U12420 (N_12420,N_10461,N_10388);
nand U12421 (N_12421,N_10460,N_11751);
xor U12422 (N_12422,N_11152,N_10818);
or U12423 (N_12423,N_11818,N_11678);
and U12424 (N_12424,N_11154,N_11945);
xor U12425 (N_12425,N_10078,N_10989);
nand U12426 (N_12426,N_10961,N_11796);
or U12427 (N_12427,N_11671,N_11135);
and U12428 (N_12428,N_10205,N_10356);
nand U12429 (N_12429,N_11760,N_11877);
nand U12430 (N_12430,N_11125,N_11948);
nand U12431 (N_12431,N_11331,N_11317);
nor U12432 (N_12432,N_11528,N_11766);
nand U12433 (N_12433,N_11752,N_10007);
xnor U12434 (N_12434,N_10884,N_10006);
or U12435 (N_12435,N_11251,N_10441);
nor U12436 (N_12436,N_10036,N_10634);
nor U12437 (N_12437,N_11361,N_10896);
or U12438 (N_12438,N_10069,N_11352);
nand U12439 (N_12439,N_11424,N_11177);
nand U12440 (N_12440,N_11289,N_11288);
and U12441 (N_12441,N_11792,N_11446);
and U12442 (N_12442,N_11905,N_10683);
and U12443 (N_12443,N_11858,N_10959);
and U12444 (N_12444,N_10598,N_11567);
or U12445 (N_12445,N_11192,N_11722);
xnor U12446 (N_12446,N_10657,N_10364);
and U12447 (N_12447,N_11431,N_10079);
xnor U12448 (N_12448,N_11561,N_11719);
or U12449 (N_12449,N_11432,N_10890);
or U12450 (N_12450,N_11373,N_11956);
or U12451 (N_12451,N_10593,N_11836);
xor U12452 (N_12452,N_10474,N_11258);
nand U12453 (N_12453,N_10355,N_11754);
or U12454 (N_12454,N_10726,N_11968);
nand U12455 (N_12455,N_10728,N_11666);
nand U12456 (N_12456,N_11132,N_11799);
nor U12457 (N_12457,N_10271,N_11756);
or U12458 (N_12458,N_10440,N_10145);
nand U12459 (N_12459,N_11805,N_11159);
and U12460 (N_12460,N_11591,N_11544);
nor U12461 (N_12461,N_11024,N_10851);
nor U12462 (N_12462,N_11902,N_11079);
nand U12463 (N_12463,N_10381,N_10941);
or U12464 (N_12464,N_10073,N_10921);
and U12465 (N_12465,N_10049,N_11325);
nor U12466 (N_12466,N_11961,N_11967);
nor U12467 (N_12467,N_11259,N_11740);
or U12468 (N_12468,N_11636,N_11221);
xor U12469 (N_12469,N_10199,N_10669);
and U12470 (N_12470,N_11727,N_10977);
xor U12471 (N_12471,N_11032,N_10667);
nor U12472 (N_12472,N_10616,N_10945);
or U12473 (N_12473,N_11886,N_11042);
xnor U12474 (N_12474,N_10370,N_11614);
and U12475 (N_12475,N_11436,N_10279);
nor U12476 (N_12476,N_10285,N_11900);
nor U12477 (N_12477,N_10864,N_11140);
and U12478 (N_12478,N_11534,N_10737);
nand U12479 (N_12479,N_10573,N_10750);
xor U12480 (N_12480,N_11316,N_11662);
xor U12481 (N_12481,N_11683,N_10692);
xnor U12482 (N_12482,N_11540,N_10443);
nand U12483 (N_12483,N_11490,N_10677);
nor U12484 (N_12484,N_10603,N_11401);
nand U12485 (N_12485,N_11633,N_11310);
xnor U12486 (N_12486,N_11291,N_11230);
or U12487 (N_12487,N_10812,N_11189);
nor U12488 (N_12488,N_10899,N_11954);
nor U12489 (N_12489,N_10169,N_10837);
and U12490 (N_12490,N_10928,N_10091);
and U12491 (N_12491,N_11744,N_10984);
or U12492 (N_12492,N_10165,N_11674);
and U12493 (N_12493,N_10482,N_11233);
xor U12494 (N_12494,N_10238,N_10293);
nor U12495 (N_12495,N_11594,N_11870);
nand U12496 (N_12496,N_10658,N_11298);
xnor U12497 (N_12497,N_11510,N_11315);
nor U12498 (N_12498,N_11060,N_10028);
nand U12499 (N_12499,N_10120,N_11839);
nor U12500 (N_12500,N_11696,N_11151);
nor U12501 (N_12501,N_10712,N_10108);
and U12502 (N_12502,N_10242,N_10002);
and U12503 (N_12503,N_11850,N_11308);
nand U12504 (N_12504,N_11586,N_10170);
and U12505 (N_12505,N_10064,N_10604);
xnor U12506 (N_12506,N_11514,N_10794);
and U12507 (N_12507,N_10163,N_10229);
nand U12508 (N_12508,N_11176,N_11981);
xor U12509 (N_12509,N_11894,N_10580);
xor U12510 (N_12510,N_10218,N_11686);
xnor U12511 (N_12511,N_10240,N_11016);
nor U12512 (N_12512,N_10566,N_10548);
nand U12513 (N_12513,N_11755,N_11209);
and U12514 (N_12514,N_11646,N_10568);
nor U12515 (N_12515,N_11136,N_10546);
and U12516 (N_12516,N_11612,N_10586);
nand U12517 (N_12517,N_11018,N_10094);
xor U12518 (N_12518,N_10863,N_11764);
nand U12519 (N_12519,N_11153,N_10273);
and U12520 (N_12520,N_10918,N_11393);
xor U12521 (N_12521,N_11382,N_11085);
or U12522 (N_12522,N_10764,N_10836);
xor U12523 (N_12523,N_10032,N_11353);
nand U12524 (N_12524,N_10840,N_10567);
nand U12525 (N_12525,N_10575,N_10532);
xor U12526 (N_12526,N_10627,N_10985);
nand U12527 (N_12527,N_11475,N_10787);
xnor U12528 (N_12528,N_11427,N_11556);
nand U12529 (N_12529,N_11575,N_11146);
or U12530 (N_12530,N_10588,N_11742);
xnor U12531 (N_12531,N_11604,N_11414);
nor U12532 (N_12532,N_10582,N_11029);
nor U12533 (N_12533,N_10796,N_10221);
nor U12534 (N_12534,N_11526,N_10676);
and U12535 (N_12535,N_10926,N_10042);
nand U12536 (N_12536,N_11655,N_10872);
xnor U12537 (N_12537,N_11715,N_11728);
nand U12538 (N_12538,N_11266,N_11458);
and U12539 (N_12539,N_10444,N_10611);
nand U12540 (N_12540,N_11921,N_10555);
nand U12541 (N_12541,N_11511,N_11668);
nor U12542 (N_12542,N_11896,N_10822);
and U12543 (N_12543,N_10618,N_10115);
and U12544 (N_12544,N_11357,N_11955);
xor U12545 (N_12545,N_11623,N_11519);
nor U12546 (N_12546,N_11117,N_10722);
nor U12547 (N_12547,N_11704,N_11832);
nand U12548 (N_12548,N_10901,N_10641);
and U12549 (N_12549,N_11876,N_10332);
or U12550 (N_12550,N_11828,N_11086);
xor U12551 (N_12551,N_11257,N_11014);
or U12552 (N_12552,N_10581,N_11568);
nor U12553 (N_12553,N_11776,N_11104);
nor U12554 (N_12554,N_11616,N_11887);
nand U12555 (N_12555,N_11173,N_10228);
nand U12556 (N_12556,N_10656,N_10917);
xnor U12557 (N_12557,N_11456,N_10311);
xor U12558 (N_12558,N_10310,N_11548);
xnor U12559 (N_12559,N_10159,N_11536);
xnor U12560 (N_12560,N_10801,N_10991);
xnor U12561 (N_12561,N_11815,N_10819);
or U12562 (N_12562,N_11452,N_10011);
and U12563 (N_12563,N_11049,N_11384);
xor U12564 (N_12564,N_10865,N_11404);
xnor U12565 (N_12565,N_10429,N_11509);
and U12566 (N_12566,N_11263,N_10458);
and U12567 (N_12567,N_11853,N_11093);
and U12568 (N_12568,N_11903,N_10408);
nand U12569 (N_12569,N_11368,N_10043);
and U12570 (N_12570,N_10114,N_10561);
or U12571 (N_12571,N_10421,N_10276);
or U12572 (N_12572,N_11290,N_10732);
and U12573 (N_12573,N_10763,N_10972);
or U12574 (N_12574,N_10383,N_10867);
nand U12575 (N_12575,N_10902,N_11947);
or U12576 (N_12576,N_10354,N_11787);
nand U12577 (N_12577,N_10997,N_10401);
nor U12578 (N_12578,N_10909,N_11008);
or U12579 (N_12579,N_11659,N_11340);
or U12580 (N_12580,N_11542,N_11336);
or U12581 (N_12581,N_11163,N_10389);
nand U12582 (N_12582,N_11562,N_11065);
and U12583 (N_12583,N_11860,N_11381);
nor U12584 (N_12584,N_11194,N_11524);
nor U12585 (N_12585,N_11022,N_11838);
or U12586 (N_12586,N_11532,N_11305);
xor U12587 (N_12587,N_11605,N_11950);
and U12588 (N_12588,N_10533,N_11466);
and U12589 (N_12589,N_11100,N_10574);
and U12590 (N_12590,N_11498,N_11463);
or U12591 (N_12591,N_11824,N_11571);
nor U12592 (N_12592,N_10148,N_11765);
or U12593 (N_12593,N_11960,N_10993);
or U12594 (N_12594,N_11212,N_11443);
or U12595 (N_12595,N_10266,N_11987);
nor U12596 (N_12596,N_11389,N_10267);
nand U12597 (N_12597,N_11464,N_11971);
nand U12598 (N_12598,N_10377,N_11488);
nor U12599 (N_12599,N_10600,N_11500);
and U12600 (N_12600,N_10405,N_10263);
xor U12601 (N_12601,N_11557,N_10420);
xnor U12602 (N_12602,N_11629,N_10119);
nor U12603 (N_12603,N_11061,N_10149);
and U12604 (N_12604,N_11861,N_11798);
and U12605 (N_12605,N_10040,N_10475);
nor U12606 (N_12606,N_11809,N_11994);
and U12607 (N_12607,N_11682,N_11979);
nand U12608 (N_12608,N_11916,N_11250);
nor U12609 (N_12609,N_11502,N_11999);
and U12610 (N_12610,N_11309,N_11092);
nand U12611 (N_12611,N_11138,N_11652);
or U12612 (N_12612,N_11907,N_11294);
nor U12613 (N_12613,N_11169,N_10833);
xnor U12614 (N_12614,N_11269,N_11026);
nor U12615 (N_12615,N_10112,N_10301);
xnor U12616 (N_12616,N_11553,N_11716);
nor U12617 (N_12617,N_10146,N_10946);
xor U12618 (N_12618,N_10140,N_10619);
nor U12619 (N_12619,N_11848,N_10024);
and U12620 (N_12620,N_11739,N_10509);
or U12621 (N_12621,N_10883,N_10430);
xor U12622 (N_12622,N_10178,N_11709);
xor U12623 (N_12623,N_11773,N_11073);
or U12624 (N_12624,N_11953,N_11603);
xnor U12625 (N_12625,N_10987,N_10866);
and U12626 (N_12626,N_10975,N_11148);
nor U12627 (N_12627,N_11006,N_10786);
and U12628 (N_12628,N_10980,N_10333);
nand U12629 (N_12629,N_10711,N_11292);
or U12630 (N_12630,N_10889,N_11362);
or U12631 (N_12631,N_11952,N_10922);
xor U12632 (N_12632,N_11405,N_10844);
nor U12633 (N_12633,N_11923,N_11476);
and U12634 (N_12634,N_10367,N_11386);
xnor U12635 (N_12635,N_10477,N_11267);
and U12636 (N_12636,N_11578,N_11391);
nand U12637 (N_12637,N_11606,N_10804);
xnor U12638 (N_12638,N_11889,N_11096);
nand U12639 (N_12639,N_10174,N_10158);
and U12640 (N_12640,N_10188,N_10409);
xnor U12641 (N_12641,N_11541,N_11930);
nand U12642 (N_12642,N_10638,N_11064);
xnor U12643 (N_12643,N_11162,N_10793);
nand U12644 (N_12644,N_11312,N_11849);
nand U12645 (N_12645,N_10526,N_10468);
and U12646 (N_12646,N_10690,N_10510);
nor U12647 (N_12647,N_11645,N_10280);
xnor U12648 (N_12648,N_11992,N_11851);
xor U12649 (N_12649,N_10816,N_11926);
and U12650 (N_12650,N_11207,N_11409);
or U12651 (N_12651,N_10304,N_11487);
xor U12652 (N_12652,N_10009,N_10932);
nand U12653 (N_12653,N_10554,N_10190);
nand U12654 (N_12654,N_11757,N_10005);
nand U12655 (N_12655,N_11306,N_11909);
nor U12656 (N_12656,N_11537,N_10806);
or U12657 (N_12657,N_10410,N_11396);
nand U12658 (N_12658,N_10453,N_10349);
nand U12659 (N_12659,N_10665,N_10396);
nor U12660 (N_12660,N_10775,N_10647);
or U12661 (N_12661,N_10291,N_11749);
or U12662 (N_12662,N_10594,N_10590);
and U12663 (N_12663,N_10117,N_10957);
xor U12664 (N_12664,N_11098,N_11112);
and U12665 (N_12665,N_10960,N_11489);
nor U12666 (N_12666,N_10109,N_11088);
and U12667 (N_12667,N_11651,N_10258);
or U12668 (N_12668,N_10136,N_11158);
or U12669 (N_12669,N_10300,N_11581);
or U12670 (N_12670,N_11474,N_10014);
and U12671 (N_12671,N_11720,N_11694);
and U12672 (N_12672,N_10296,N_11101);
and U12673 (N_12673,N_10713,N_11746);
and U12674 (N_12674,N_11037,N_10399);
nand U12675 (N_12675,N_11326,N_10147);
nand U12676 (N_12676,N_10644,N_11272);
nand U12677 (N_12677,N_10424,N_10216);
and U12678 (N_12678,N_10920,N_11533);
nor U12679 (N_12679,N_11501,N_10082);
or U12680 (N_12680,N_11513,N_11723);
and U12681 (N_12681,N_11213,N_11503);
nor U12682 (N_12682,N_10570,N_11460);
nand U12683 (N_12683,N_10852,N_10530);
or U12684 (N_12684,N_11351,N_10196);
or U12685 (N_12685,N_11044,N_11865);
nor U12686 (N_12686,N_10075,N_11484);
nor U12687 (N_12687,N_10988,N_11644);
and U12688 (N_12688,N_11041,N_10487);
nor U12689 (N_12689,N_11001,N_11966);
or U12690 (N_12690,N_10757,N_10360);
nand U12691 (N_12691,N_10236,N_11610);
nand U12692 (N_12692,N_10516,N_10857);
and U12693 (N_12693,N_10629,N_11428);
and U12694 (N_12694,N_11750,N_10249);
nor U12695 (N_12695,N_10706,N_11525);
and U12696 (N_12696,N_11479,N_10735);
nor U12697 (N_12697,N_11429,N_10790);
or U12698 (N_12698,N_10046,N_11738);
nor U12699 (N_12699,N_10001,N_10628);
and U12700 (N_12700,N_10719,N_10871);
nand U12701 (N_12701,N_11808,N_11010);
nor U12702 (N_12702,N_11081,N_11640);
or U12703 (N_12703,N_10135,N_11763);
xor U12704 (N_12704,N_10189,N_11121);
nor U12705 (N_12705,N_11518,N_10150);
and U12706 (N_12706,N_10141,N_10684);
xnor U12707 (N_12707,N_10270,N_11197);
nand U12708 (N_12708,N_10873,N_11226);
nor U12709 (N_12709,N_10970,N_11185);
or U12710 (N_12710,N_10038,N_10222);
or U12711 (N_12711,N_10264,N_10449);
and U12712 (N_12712,N_10823,N_11982);
nor U12713 (N_12713,N_10417,N_11144);
xnor U12714 (N_12714,N_11271,N_10870);
or U12715 (N_12715,N_11579,N_10621);
nand U12716 (N_12716,N_11813,N_10724);
nor U12717 (N_12717,N_11522,N_10272);
and U12718 (N_12718,N_10976,N_11977);
nand U12719 (N_12719,N_11769,N_10767);
xor U12720 (N_12720,N_10913,N_11814);
nor U12721 (N_12721,N_10855,N_10456);
xor U12722 (N_12722,N_10557,N_11863);
nand U12723 (N_12723,N_10780,N_11398);
nor U12724 (N_12724,N_11240,N_11422);
nand U12725 (N_12725,N_10535,N_11497);
or U12726 (N_12726,N_10912,N_10769);
xor U12727 (N_12727,N_10459,N_11988);
xnor U12728 (N_12728,N_11455,N_10937);
and U12729 (N_12729,N_11933,N_10777);
or U12730 (N_12730,N_10309,N_11549);
or U12731 (N_12731,N_10051,N_11403);
and U12732 (N_12732,N_11411,N_11472);
nor U12733 (N_12733,N_11811,N_11434);
xnor U12734 (N_12734,N_10749,N_10252);
nor U12735 (N_12735,N_10963,N_11767);
xnor U12736 (N_12736,N_11551,N_10981);
or U12737 (N_12737,N_10613,N_10290);
and U12738 (N_12738,N_10564,N_11874);
nor U12739 (N_12739,N_10848,N_11199);
and U12740 (N_12740,N_10084,N_11937);
xnor U12741 (N_12741,N_10699,N_11167);
nor U12742 (N_12742,N_11149,N_11951);
or U12743 (N_12743,N_11421,N_10938);
and U12744 (N_12744,N_11855,N_10842);
and U12745 (N_12745,N_11569,N_11461);
and U12746 (N_12746,N_11214,N_11478);
nor U12747 (N_12747,N_11342,N_11202);
and U12748 (N_12748,N_10302,N_10053);
nand U12749 (N_12749,N_10962,N_11066);
or U12750 (N_12750,N_11539,N_11732);
or U12751 (N_12751,N_11395,N_10350);
xor U12752 (N_12752,N_11036,N_10127);
or U12753 (N_12753,N_11009,N_10868);
nand U12754 (N_12754,N_10521,N_11347);
nand U12755 (N_12755,N_10143,N_11810);
or U12756 (N_12756,N_10760,N_11457);
nor U12757 (N_12757,N_10765,N_11637);
nor U12758 (N_12758,N_10679,N_11015);
nand U12759 (N_12759,N_10164,N_10208);
or U12760 (N_12760,N_11989,N_11122);
or U12761 (N_12761,N_10825,N_11844);
or U12762 (N_12762,N_11109,N_11245);
or U12763 (N_12763,N_11871,N_10631);
nand U12764 (N_12764,N_10226,N_11690);
xor U12765 (N_12765,N_10363,N_11910);
nor U12766 (N_12766,N_10241,N_11426);
or U12767 (N_12767,N_11718,N_11354);
nand U12768 (N_12768,N_10203,N_11119);
nand U12769 (N_12769,N_11296,N_11433);
xnor U12770 (N_12770,N_11759,N_11774);
xor U12771 (N_12771,N_10622,N_11692);
nor U12772 (N_12772,N_10467,N_10187);
xnor U12773 (N_12773,N_11842,N_10671);
xor U12774 (N_12774,N_10746,N_11164);
nor U12775 (N_12775,N_10874,N_11670);
xor U12776 (N_12776,N_11447,N_11000);
or U12777 (N_12777,N_10931,N_11959);
nand U12778 (N_12778,N_10828,N_10277);
nor U12779 (N_12779,N_11232,N_10500);
or U12780 (N_12780,N_11845,N_11505);
or U12781 (N_12781,N_10101,N_11701);
nor U12782 (N_12782,N_11450,N_10689);
nor U12783 (N_12783,N_11617,N_10880);
nand U12784 (N_12784,N_10104,N_10895);
nor U12785 (N_12785,N_10534,N_11491);
nor U12786 (N_12786,N_11023,N_11059);
xor U12787 (N_12787,N_10527,N_11406);
xnor U12788 (N_12788,N_11045,N_10805);
xor U12789 (N_12789,N_11835,N_10308);
or U12790 (N_12790,N_11094,N_10322);
xor U12791 (N_12791,N_10649,N_11335);
and U12792 (N_12792,N_10716,N_11918);
nand U12793 (N_12793,N_11669,N_10018);
or U12794 (N_12794,N_11438,N_10788);
nand U12795 (N_12795,N_11182,N_11328);
or U12796 (N_12796,N_11074,N_11964);
and U12797 (N_12797,N_10881,N_11527);
xnor U12798 (N_12798,N_10687,N_10673);
nor U12799 (N_12799,N_10563,N_10834);
nor U12800 (N_12800,N_10340,N_10625);
xnor U12801 (N_12801,N_10646,N_10067);
and U12802 (N_12802,N_11826,N_10846);
or U12803 (N_12803,N_11252,N_11480);
nor U12804 (N_12804,N_10537,N_10965);
nor U12805 (N_12805,N_10025,N_10385);
xnor U12806 (N_12806,N_10193,N_10662);
nand U12807 (N_12807,N_10802,N_11007);
xor U12808 (N_12808,N_10967,N_11847);
xnor U12809 (N_12809,N_11914,N_11186);
nand U12810 (N_12810,N_10529,N_10063);
nor U12811 (N_12811,N_11183,N_11178);
nand U12812 (N_12812,N_11243,N_10201);
nor U12813 (N_12813,N_11929,N_11190);
or U12814 (N_12814,N_10029,N_10784);
and U12815 (N_12815,N_10923,N_11679);
nand U12816 (N_12816,N_10808,N_11280);
xor U12817 (N_12817,N_11172,N_11219);
and U12818 (N_12818,N_11242,N_10338);
and U12819 (N_12819,N_11706,N_10050);
nor U12820 (N_12820,N_10483,N_11415);
nor U12821 (N_12821,N_10123,N_11917);
and U12822 (N_12822,N_11260,N_10569);
or U12823 (N_12823,N_10403,N_11676);
nand U12824 (N_12824,N_11599,N_11806);
nand U12825 (N_12825,N_11307,N_10348);
and U12826 (N_12826,N_10269,N_11546);
xnor U12827 (N_12827,N_11072,N_10297);
or U12828 (N_12828,N_10971,N_10110);
nand U12829 (N_12829,N_11596,N_10312);
xor U12830 (N_12830,N_10617,N_10327);
and U12831 (N_12831,N_11975,N_10826);
nand U12832 (N_12832,N_10709,N_10257);
nor U12833 (N_12833,N_10076,N_11608);
nor U12834 (N_12834,N_11465,N_11224);
or U12835 (N_12835,N_10661,N_11210);
nor U12836 (N_12836,N_10727,N_10268);
nor U12837 (N_12837,N_11442,N_10118);
and U12838 (N_12838,N_11695,N_11239);
xnor U12839 (N_12839,N_10892,N_10232);
and U12840 (N_12840,N_10446,N_10185);
nor U12841 (N_12841,N_11521,N_11587);
nand U12842 (N_12842,N_11033,N_11588);
and U12843 (N_12843,N_10142,N_11857);
nor U12844 (N_12844,N_11397,N_11004);
xnor U12845 (N_12845,N_11217,N_10773);
xnor U12846 (N_12846,N_11237,N_10172);
xor U12847 (N_12847,N_11270,N_10020);
nor U12848 (N_12848,N_10663,N_10789);
nand U12849 (N_12849,N_11058,N_10860);
or U12850 (N_12850,N_11345,N_11445);
nor U12851 (N_12851,N_11283,N_10664);
xnor U12852 (N_12852,N_10894,N_11729);
nand U12853 (N_12853,N_11801,N_11725);
nor U12854 (N_12854,N_10080,N_11831);
xnor U12855 (N_12855,N_11425,N_10450);
nor U12856 (N_12856,N_11978,N_11980);
nand U12857 (N_12857,N_11360,N_10202);
xnor U12858 (N_12858,N_11031,N_11737);
xnor U12859 (N_12859,N_11078,N_10910);
xor U12860 (N_12860,N_10875,N_11303);
nor U12861 (N_12861,N_10958,N_11807);
and U12862 (N_12862,N_11021,N_10294);
nor U12863 (N_12863,N_11449,N_10211);
and U12864 (N_12864,N_11589,N_10885);
nand U12865 (N_12865,N_11107,N_11337);
or U12866 (N_12866,N_11012,N_10298);
nor U12867 (N_12867,N_10375,N_10717);
or U12868 (N_12868,N_10329,N_10653);
xnor U12869 (N_12869,N_10685,N_10404);
xor U12870 (N_12870,N_10194,N_10039);
nor U12871 (N_12871,N_11830,N_11131);
nor U12872 (N_12872,N_10448,N_11791);
nor U12873 (N_12873,N_10845,N_11647);
and U12874 (N_12874,N_10031,N_10897);
nand U12875 (N_12875,N_11113,N_10589);
and U12876 (N_12876,N_11030,N_10650);
and U12877 (N_12877,N_11911,N_10434);
nor U12878 (N_12878,N_10830,N_10137);
nand U12879 (N_12879,N_11687,N_10274);
xnor U12880 (N_12880,N_10666,N_11635);
or U12881 (N_12881,N_10215,N_11321);
or U12882 (N_12882,N_11372,N_11585);
xnor U12883 (N_12883,N_11322,N_10572);
xnor U12884 (N_12884,N_11115,N_10708);
xnor U12885 (N_12885,N_11613,N_11708);
nand U12886 (N_12886,N_11735,N_10512);
and U12887 (N_12887,N_11563,N_11392);
and U12888 (N_12888,N_10583,N_10951);
xor U12889 (N_12889,N_10284,N_10964);
or U12890 (N_12890,N_10858,N_11348);
nor U12891 (N_12891,N_10436,N_10394);
nand U12892 (N_12892,N_11375,N_11821);
and U12893 (N_12893,N_10772,N_10626);
and U12894 (N_12894,N_11071,N_11506);
nand U12895 (N_12895,N_11794,N_11962);
or U12896 (N_12896,N_10442,N_10368);
xor U12897 (N_12897,N_10484,N_10307);
xor U12898 (N_12898,N_10431,N_11804);
nand U12899 (N_12899,N_11882,N_11515);
or U12900 (N_12900,N_11693,N_10343);
xnor U12901 (N_12901,N_11105,N_11091);
and U12902 (N_12902,N_10337,N_10869);
nand U12903 (N_12903,N_11782,N_10606);
xnor U12904 (N_12904,N_10522,N_11145);
and U12905 (N_12905,N_11264,N_11703);
or U12906 (N_12906,N_10418,N_10924);
nor U12907 (N_12907,N_10956,N_10245);
nand U12908 (N_12908,N_10599,N_11843);
nand U12909 (N_12909,N_10778,N_10052);
nor U12910 (N_12910,N_10659,N_11658);
xor U12911 (N_12911,N_11126,N_11028);
nor U12912 (N_12912,N_10969,N_10447);
nor U12913 (N_12913,N_10925,N_10710);
or U12914 (N_12914,N_10499,N_10087);
nand U12915 (N_12915,N_11995,N_10125);
and U12916 (N_12916,N_10528,N_10030);
xnor U12917 (N_12917,N_11663,N_10633);
nor U12918 (N_12918,N_11187,N_10729);
nand U12919 (N_12919,N_11949,N_10807);
and U12920 (N_12920,N_11492,N_10346);
nand U12921 (N_12921,N_11039,N_10230);
xor U12922 (N_12922,N_10491,N_10214);
nor U12923 (N_12923,N_11624,N_11825);
and U12924 (N_12924,N_10351,N_10682);
and U12925 (N_12925,N_11448,N_11883);
xnor U12926 (N_12926,N_11915,N_10559);
and U12927 (N_12927,N_11390,N_10498);
xor U12928 (N_12928,N_10608,N_11741);
xor U12929 (N_12929,N_10688,N_10426);
or U12930 (N_12930,N_11783,N_11642);
nor U12931 (N_12931,N_10998,N_10213);
xnor U12932 (N_12932,N_10577,N_10182);
nor U12933 (N_12933,N_10911,N_10550);
nand U12934 (N_12934,N_10054,N_10122);
xnor U12935 (N_12935,N_10425,N_10066);
nand U12936 (N_12936,N_11133,N_11697);
and U12937 (N_12937,N_11102,N_10935);
xor U12938 (N_12938,N_10553,N_11592);
nor U12939 (N_12939,N_10831,N_10551);
nand U12940 (N_12940,N_10640,N_10225);
nand U12941 (N_12941,N_11607,N_10999);
nand U12942 (N_12942,N_11572,N_10486);
or U12943 (N_12943,N_11462,N_10996);
nor U12944 (N_12944,N_11376,N_10353);
nand U12945 (N_12945,N_11228,N_11180);
nor U12946 (N_12946,N_11965,N_10116);
or U12947 (N_12947,N_10652,N_10097);
nor U12948 (N_12948,N_11856,N_11063);
nor U12949 (N_12949,N_11919,N_10623);
xnor U12950 (N_12950,N_11958,N_10210);
xnor U12951 (N_12951,N_10256,N_10966);
xnor U12952 (N_12952,N_11780,N_11639);
xor U12953 (N_12953,N_10639,N_11184);
nor U12954 (N_12954,N_10655,N_11935);
nand U12955 (N_12955,N_11356,N_11685);
or U12956 (N_12956,N_11499,N_11027);
and U12957 (N_12957,N_10715,N_10204);
xnor U12958 (N_12958,N_11056,N_10195);
and U12959 (N_12959,N_11048,N_10278);
xor U12960 (N_12960,N_10107,N_11986);
nor U12961 (N_12961,N_10940,N_11341);
nand U12962 (N_12962,N_10514,N_10217);
or U12963 (N_12963,N_10472,N_10111);
nand U12964 (N_12964,N_11908,N_11195);
nand U12965 (N_12965,N_10089,N_11665);
or U12966 (N_12966,N_10792,N_10607);
and U12967 (N_12967,N_11717,N_10233);
or U12968 (N_12968,N_11193,N_10318);
xor U12969 (N_12969,N_10292,N_10513);
nand U12970 (N_12970,N_10386,N_11788);
xnor U12971 (N_12971,N_10254,N_10065);
or U12972 (N_12972,N_10438,N_10197);
nor U12973 (N_12973,N_11408,N_11363);
nor U12974 (N_12974,N_10314,N_11888);
nand U12975 (N_12975,N_11714,N_11778);
or U12976 (N_12976,N_11155,N_10660);
xnor U12977 (N_12977,N_11076,N_10944);
nor U12978 (N_12978,N_10061,N_11002);
and U12979 (N_12979,N_11555,N_10615);
nor U12980 (N_12980,N_10850,N_10048);
and U12981 (N_12981,N_10782,N_11906);
and U12982 (N_12982,N_11711,N_11020);
or U12983 (N_12983,N_10704,N_11278);
and U12984 (N_12984,N_10334,N_11244);
nand U12985 (N_12985,N_11249,N_11859);
nand U12986 (N_12986,N_11196,N_10734);
xor U12987 (N_12987,N_10741,N_10173);
nor U12988 (N_12988,N_11673,N_10224);
nor U12989 (N_12989,N_10904,N_10124);
or U12990 (N_12990,N_10361,N_11595);
nand U12991 (N_12991,N_11111,N_11274);
or U12992 (N_12992,N_11713,N_11993);
nand U12993 (N_12993,N_11013,N_10695);
nor U12994 (N_12994,N_11459,N_11504);
xnor U12995 (N_12995,N_10674,N_11175);
or U12996 (N_12996,N_10714,N_10547);
nand U12997 (N_12997,N_11374,N_11913);
xor U12998 (N_12998,N_11622,N_11641);
xor U12999 (N_12999,N_11034,N_10088);
nand U13000 (N_13000,N_10193,N_10370);
or U13001 (N_13001,N_11854,N_11716);
nand U13002 (N_13002,N_11018,N_11203);
and U13003 (N_13003,N_11598,N_10999);
and U13004 (N_13004,N_10838,N_10953);
nor U13005 (N_13005,N_10928,N_11074);
or U13006 (N_13006,N_11441,N_10332);
nor U13007 (N_13007,N_11262,N_11736);
and U13008 (N_13008,N_11907,N_10800);
and U13009 (N_13009,N_11165,N_10448);
nand U13010 (N_13010,N_10762,N_10227);
nor U13011 (N_13011,N_11151,N_11789);
or U13012 (N_13012,N_11335,N_11656);
or U13013 (N_13013,N_11814,N_11414);
and U13014 (N_13014,N_10204,N_10961);
or U13015 (N_13015,N_10803,N_10883);
or U13016 (N_13016,N_10330,N_10410);
nor U13017 (N_13017,N_11612,N_11293);
or U13018 (N_13018,N_11142,N_11389);
or U13019 (N_13019,N_10034,N_11900);
xnor U13020 (N_13020,N_10349,N_11132);
nor U13021 (N_13021,N_10522,N_10155);
nor U13022 (N_13022,N_10455,N_11897);
xnor U13023 (N_13023,N_10381,N_10259);
and U13024 (N_13024,N_11828,N_11431);
nor U13025 (N_13025,N_10742,N_10518);
and U13026 (N_13026,N_10340,N_11095);
nor U13027 (N_13027,N_10225,N_11851);
nor U13028 (N_13028,N_10472,N_10627);
or U13029 (N_13029,N_10051,N_10934);
xnor U13030 (N_13030,N_10724,N_10770);
and U13031 (N_13031,N_11553,N_10630);
and U13032 (N_13032,N_10716,N_11141);
or U13033 (N_13033,N_10853,N_11042);
nand U13034 (N_13034,N_10212,N_11707);
or U13035 (N_13035,N_10531,N_10731);
nor U13036 (N_13036,N_11256,N_11167);
xnor U13037 (N_13037,N_10671,N_10166);
nand U13038 (N_13038,N_10984,N_10914);
or U13039 (N_13039,N_10644,N_11817);
or U13040 (N_13040,N_11920,N_10542);
nand U13041 (N_13041,N_11863,N_10514);
xor U13042 (N_13042,N_10158,N_10871);
or U13043 (N_13043,N_11277,N_11964);
nor U13044 (N_13044,N_11103,N_10719);
xor U13045 (N_13045,N_11806,N_10732);
nand U13046 (N_13046,N_10060,N_11093);
nand U13047 (N_13047,N_10066,N_11304);
xor U13048 (N_13048,N_10284,N_11056);
xor U13049 (N_13049,N_11754,N_11470);
nor U13050 (N_13050,N_11348,N_10203);
nor U13051 (N_13051,N_11087,N_10046);
nand U13052 (N_13052,N_10647,N_11526);
nor U13053 (N_13053,N_10624,N_10936);
nor U13054 (N_13054,N_11125,N_10111);
and U13055 (N_13055,N_10759,N_11925);
nor U13056 (N_13056,N_10158,N_11355);
nor U13057 (N_13057,N_11224,N_10325);
and U13058 (N_13058,N_10146,N_11871);
nor U13059 (N_13059,N_10792,N_11087);
or U13060 (N_13060,N_11611,N_10196);
nand U13061 (N_13061,N_10613,N_11480);
xnor U13062 (N_13062,N_11969,N_10205);
or U13063 (N_13063,N_10661,N_10321);
or U13064 (N_13064,N_11452,N_11567);
or U13065 (N_13065,N_11030,N_11888);
xnor U13066 (N_13066,N_11182,N_10507);
nor U13067 (N_13067,N_10627,N_10872);
xnor U13068 (N_13068,N_11205,N_10029);
nand U13069 (N_13069,N_10053,N_11129);
nor U13070 (N_13070,N_10251,N_11556);
nor U13071 (N_13071,N_10669,N_11591);
nand U13072 (N_13072,N_11254,N_11922);
or U13073 (N_13073,N_11213,N_11403);
nor U13074 (N_13074,N_10141,N_11306);
nor U13075 (N_13075,N_10852,N_11638);
or U13076 (N_13076,N_11145,N_11798);
nor U13077 (N_13077,N_11511,N_10424);
and U13078 (N_13078,N_10159,N_11521);
nand U13079 (N_13079,N_11725,N_10107);
nor U13080 (N_13080,N_10491,N_11385);
and U13081 (N_13081,N_10417,N_10932);
nor U13082 (N_13082,N_11774,N_10322);
nand U13083 (N_13083,N_11448,N_10117);
nand U13084 (N_13084,N_10668,N_10809);
xnor U13085 (N_13085,N_11734,N_10230);
or U13086 (N_13086,N_11530,N_11347);
or U13087 (N_13087,N_11195,N_10805);
nand U13088 (N_13088,N_10942,N_11446);
nor U13089 (N_13089,N_10341,N_10901);
or U13090 (N_13090,N_11454,N_11196);
nand U13091 (N_13091,N_11936,N_11073);
and U13092 (N_13092,N_11439,N_11319);
and U13093 (N_13093,N_10052,N_11418);
and U13094 (N_13094,N_10117,N_11983);
nor U13095 (N_13095,N_10685,N_10550);
nand U13096 (N_13096,N_11075,N_11938);
nand U13097 (N_13097,N_10728,N_11272);
nor U13098 (N_13098,N_11896,N_10799);
or U13099 (N_13099,N_11930,N_10132);
nand U13100 (N_13100,N_10490,N_11937);
and U13101 (N_13101,N_11562,N_11697);
and U13102 (N_13102,N_10277,N_10916);
nor U13103 (N_13103,N_10124,N_11917);
xnor U13104 (N_13104,N_11992,N_11493);
xnor U13105 (N_13105,N_10193,N_11038);
or U13106 (N_13106,N_11148,N_10790);
or U13107 (N_13107,N_10075,N_11342);
or U13108 (N_13108,N_10963,N_11802);
or U13109 (N_13109,N_11839,N_10624);
and U13110 (N_13110,N_10741,N_10912);
or U13111 (N_13111,N_11280,N_10529);
and U13112 (N_13112,N_11456,N_11651);
nand U13113 (N_13113,N_10331,N_11151);
nor U13114 (N_13114,N_10814,N_11855);
xnor U13115 (N_13115,N_11340,N_10720);
or U13116 (N_13116,N_11764,N_10938);
xor U13117 (N_13117,N_10163,N_11083);
nand U13118 (N_13118,N_11387,N_10410);
or U13119 (N_13119,N_11570,N_11696);
and U13120 (N_13120,N_10567,N_10642);
and U13121 (N_13121,N_11130,N_10112);
and U13122 (N_13122,N_11288,N_11152);
and U13123 (N_13123,N_10401,N_10548);
nor U13124 (N_13124,N_10275,N_10911);
and U13125 (N_13125,N_11195,N_11132);
xor U13126 (N_13126,N_10574,N_11975);
nor U13127 (N_13127,N_11493,N_10723);
nand U13128 (N_13128,N_11981,N_11365);
nor U13129 (N_13129,N_10637,N_10864);
nand U13130 (N_13130,N_10613,N_11558);
or U13131 (N_13131,N_10376,N_11291);
and U13132 (N_13132,N_10633,N_10514);
and U13133 (N_13133,N_10481,N_11544);
nand U13134 (N_13134,N_10665,N_10353);
nand U13135 (N_13135,N_11291,N_11506);
and U13136 (N_13136,N_10522,N_10020);
and U13137 (N_13137,N_11811,N_11920);
xnor U13138 (N_13138,N_10720,N_10444);
nand U13139 (N_13139,N_10822,N_11676);
nand U13140 (N_13140,N_10347,N_10201);
nor U13141 (N_13141,N_11225,N_10546);
or U13142 (N_13142,N_10800,N_11243);
and U13143 (N_13143,N_10966,N_11820);
and U13144 (N_13144,N_10847,N_10762);
nor U13145 (N_13145,N_11562,N_11234);
nor U13146 (N_13146,N_10473,N_11734);
or U13147 (N_13147,N_11286,N_10109);
xnor U13148 (N_13148,N_11853,N_11828);
nor U13149 (N_13149,N_11583,N_11002);
and U13150 (N_13150,N_11594,N_11673);
or U13151 (N_13151,N_11275,N_11412);
xnor U13152 (N_13152,N_10638,N_11831);
nand U13153 (N_13153,N_10145,N_10591);
nand U13154 (N_13154,N_11384,N_10859);
nand U13155 (N_13155,N_11922,N_11445);
nor U13156 (N_13156,N_11056,N_11394);
xnor U13157 (N_13157,N_10501,N_11826);
nor U13158 (N_13158,N_10658,N_11991);
xor U13159 (N_13159,N_11286,N_10532);
nor U13160 (N_13160,N_10273,N_10432);
or U13161 (N_13161,N_10214,N_11002);
nand U13162 (N_13162,N_11811,N_10432);
xnor U13163 (N_13163,N_11045,N_10515);
nor U13164 (N_13164,N_11688,N_11106);
or U13165 (N_13165,N_10199,N_11741);
nand U13166 (N_13166,N_11743,N_10960);
or U13167 (N_13167,N_11019,N_10961);
xnor U13168 (N_13168,N_11728,N_11058);
nor U13169 (N_13169,N_10898,N_11865);
nor U13170 (N_13170,N_10109,N_10113);
xnor U13171 (N_13171,N_10646,N_10125);
xnor U13172 (N_13172,N_11388,N_11268);
and U13173 (N_13173,N_10717,N_11894);
and U13174 (N_13174,N_11469,N_10654);
or U13175 (N_13175,N_10536,N_10924);
xor U13176 (N_13176,N_10913,N_10513);
nand U13177 (N_13177,N_11367,N_10021);
xnor U13178 (N_13178,N_11061,N_10383);
nand U13179 (N_13179,N_11846,N_10704);
and U13180 (N_13180,N_11663,N_11355);
and U13181 (N_13181,N_11732,N_10369);
nor U13182 (N_13182,N_11828,N_11040);
xor U13183 (N_13183,N_10924,N_10046);
nand U13184 (N_13184,N_10592,N_10414);
nand U13185 (N_13185,N_11993,N_11108);
xor U13186 (N_13186,N_11677,N_10064);
or U13187 (N_13187,N_10625,N_11347);
and U13188 (N_13188,N_11456,N_11917);
nor U13189 (N_13189,N_11283,N_11671);
nand U13190 (N_13190,N_11184,N_10932);
xnor U13191 (N_13191,N_10321,N_10522);
or U13192 (N_13192,N_11705,N_11228);
xnor U13193 (N_13193,N_10911,N_11915);
or U13194 (N_13194,N_11102,N_11540);
or U13195 (N_13195,N_11057,N_11347);
or U13196 (N_13196,N_10846,N_11853);
nand U13197 (N_13197,N_10110,N_11039);
nor U13198 (N_13198,N_11518,N_10534);
or U13199 (N_13199,N_11075,N_11883);
and U13200 (N_13200,N_11064,N_11418);
or U13201 (N_13201,N_10484,N_10991);
xor U13202 (N_13202,N_10885,N_10273);
and U13203 (N_13203,N_11802,N_11832);
or U13204 (N_13204,N_11416,N_10550);
nand U13205 (N_13205,N_10884,N_10125);
nor U13206 (N_13206,N_10985,N_10987);
and U13207 (N_13207,N_10706,N_10459);
and U13208 (N_13208,N_10110,N_11131);
or U13209 (N_13209,N_11982,N_11515);
xor U13210 (N_13210,N_10324,N_11879);
nand U13211 (N_13211,N_11006,N_10489);
nand U13212 (N_13212,N_10783,N_11658);
nand U13213 (N_13213,N_10206,N_11469);
nand U13214 (N_13214,N_10541,N_10335);
or U13215 (N_13215,N_11613,N_10410);
nor U13216 (N_13216,N_10866,N_10264);
nand U13217 (N_13217,N_11753,N_10669);
nor U13218 (N_13218,N_10504,N_10436);
nor U13219 (N_13219,N_10020,N_11252);
nand U13220 (N_13220,N_11681,N_10505);
xor U13221 (N_13221,N_10964,N_10609);
nand U13222 (N_13222,N_11318,N_11884);
or U13223 (N_13223,N_10891,N_11591);
nand U13224 (N_13224,N_10142,N_10354);
nor U13225 (N_13225,N_10192,N_10240);
and U13226 (N_13226,N_11982,N_11846);
and U13227 (N_13227,N_11706,N_11707);
xor U13228 (N_13228,N_11944,N_10761);
nand U13229 (N_13229,N_11172,N_11022);
nand U13230 (N_13230,N_10801,N_10288);
nor U13231 (N_13231,N_11983,N_10310);
nor U13232 (N_13232,N_10868,N_11562);
xor U13233 (N_13233,N_11691,N_11041);
nor U13234 (N_13234,N_10264,N_11569);
or U13235 (N_13235,N_11089,N_10978);
or U13236 (N_13236,N_11860,N_11316);
nand U13237 (N_13237,N_10444,N_10261);
and U13238 (N_13238,N_10524,N_11963);
or U13239 (N_13239,N_11627,N_11900);
or U13240 (N_13240,N_11860,N_11840);
nor U13241 (N_13241,N_11441,N_11883);
nand U13242 (N_13242,N_11158,N_10350);
and U13243 (N_13243,N_10420,N_10450);
xor U13244 (N_13244,N_10858,N_11084);
xnor U13245 (N_13245,N_10848,N_10213);
or U13246 (N_13246,N_10143,N_10944);
nor U13247 (N_13247,N_10369,N_11431);
nand U13248 (N_13248,N_10796,N_10262);
nand U13249 (N_13249,N_11911,N_10314);
or U13250 (N_13250,N_10446,N_10531);
and U13251 (N_13251,N_10807,N_10861);
nand U13252 (N_13252,N_11045,N_11282);
xnor U13253 (N_13253,N_10982,N_11015);
xor U13254 (N_13254,N_11936,N_11597);
nor U13255 (N_13255,N_11670,N_10136);
or U13256 (N_13256,N_10824,N_10637);
nor U13257 (N_13257,N_11338,N_11850);
nor U13258 (N_13258,N_11329,N_11158);
or U13259 (N_13259,N_11204,N_11401);
or U13260 (N_13260,N_11433,N_11862);
nand U13261 (N_13261,N_11317,N_10150);
xnor U13262 (N_13262,N_11079,N_11191);
nand U13263 (N_13263,N_11122,N_11390);
nor U13264 (N_13264,N_10002,N_11212);
or U13265 (N_13265,N_10468,N_11852);
or U13266 (N_13266,N_10757,N_11854);
or U13267 (N_13267,N_11009,N_11167);
or U13268 (N_13268,N_10324,N_11740);
xor U13269 (N_13269,N_11154,N_10144);
and U13270 (N_13270,N_10494,N_10132);
xnor U13271 (N_13271,N_11227,N_10867);
and U13272 (N_13272,N_10929,N_10888);
and U13273 (N_13273,N_11155,N_10383);
xnor U13274 (N_13274,N_10510,N_11209);
nand U13275 (N_13275,N_10312,N_10933);
or U13276 (N_13276,N_10967,N_10505);
nand U13277 (N_13277,N_11873,N_11002);
or U13278 (N_13278,N_10852,N_11608);
and U13279 (N_13279,N_11231,N_10927);
or U13280 (N_13280,N_11247,N_10734);
xnor U13281 (N_13281,N_11958,N_11763);
xor U13282 (N_13282,N_11964,N_10463);
nor U13283 (N_13283,N_10795,N_10526);
nand U13284 (N_13284,N_11183,N_11256);
xnor U13285 (N_13285,N_10137,N_10560);
or U13286 (N_13286,N_10174,N_10123);
and U13287 (N_13287,N_11101,N_11888);
xnor U13288 (N_13288,N_11339,N_10024);
nor U13289 (N_13289,N_10163,N_10026);
nor U13290 (N_13290,N_10767,N_11934);
xnor U13291 (N_13291,N_11847,N_10119);
or U13292 (N_13292,N_10619,N_10076);
or U13293 (N_13293,N_10825,N_10787);
or U13294 (N_13294,N_11585,N_11017);
and U13295 (N_13295,N_10386,N_10972);
and U13296 (N_13296,N_11083,N_10445);
nor U13297 (N_13297,N_10194,N_10708);
nand U13298 (N_13298,N_10158,N_11174);
xnor U13299 (N_13299,N_11629,N_10986);
nand U13300 (N_13300,N_11685,N_10775);
and U13301 (N_13301,N_11634,N_10860);
nor U13302 (N_13302,N_11894,N_10941);
or U13303 (N_13303,N_11376,N_10782);
and U13304 (N_13304,N_10004,N_11729);
nand U13305 (N_13305,N_10008,N_10865);
and U13306 (N_13306,N_11141,N_10038);
nor U13307 (N_13307,N_11244,N_10183);
or U13308 (N_13308,N_10361,N_11810);
nor U13309 (N_13309,N_11103,N_11257);
nor U13310 (N_13310,N_10686,N_11178);
xor U13311 (N_13311,N_10813,N_11347);
or U13312 (N_13312,N_10097,N_11698);
xor U13313 (N_13313,N_11185,N_11521);
xnor U13314 (N_13314,N_10525,N_10303);
xor U13315 (N_13315,N_11665,N_11367);
or U13316 (N_13316,N_11587,N_11031);
nand U13317 (N_13317,N_11563,N_11041);
or U13318 (N_13318,N_10234,N_10880);
nor U13319 (N_13319,N_11459,N_10367);
nand U13320 (N_13320,N_10230,N_10846);
xnor U13321 (N_13321,N_10398,N_10059);
and U13322 (N_13322,N_10888,N_10205);
nand U13323 (N_13323,N_11533,N_11786);
nor U13324 (N_13324,N_11964,N_10510);
nor U13325 (N_13325,N_11872,N_10266);
nand U13326 (N_13326,N_11954,N_11012);
xor U13327 (N_13327,N_10445,N_10068);
nand U13328 (N_13328,N_10578,N_11731);
nor U13329 (N_13329,N_10469,N_11934);
nor U13330 (N_13330,N_10820,N_10195);
nor U13331 (N_13331,N_11860,N_11085);
xor U13332 (N_13332,N_10431,N_10900);
nand U13333 (N_13333,N_10426,N_11679);
and U13334 (N_13334,N_10139,N_11455);
or U13335 (N_13335,N_11850,N_11556);
nand U13336 (N_13336,N_11683,N_11979);
and U13337 (N_13337,N_11588,N_11196);
xnor U13338 (N_13338,N_11015,N_11881);
or U13339 (N_13339,N_10957,N_10784);
and U13340 (N_13340,N_11855,N_10138);
or U13341 (N_13341,N_11682,N_10947);
and U13342 (N_13342,N_10782,N_11230);
or U13343 (N_13343,N_11919,N_10948);
nor U13344 (N_13344,N_10500,N_10886);
and U13345 (N_13345,N_11403,N_11314);
xor U13346 (N_13346,N_11540,N_10176);
or U13347 (N_13347,N_11697,N_11112);
and U13348 (N_13348,N_11484,N_11430);
and U13349 (N_13349,N_11485,N_11700);
or U13350 (N_13350,N_11720,N_11506);
nor U13351 (N_13351,N_11342,N_10545);
nand U13352 (N_13352,N_11884,N_10910);
nand U13353 (N_13353,N_11819,N_10238);
nand U13354 (N_13354,N_10786,N_10274);
xnor U13355 (N_13355,N_10076,N_10766);
nand U13356 (N_13356,N_10168,N_10855);
and U13357 (N_13357,N_11655,N_10213);
and U13358 (N_13358,N_10448,N_11220);
nand U13359 (N_13359,N_11034,N_10735);
xnor U13360 (N_13360,N_11211,N_10191);
and U13361 (N_13361,N_10303,N_10427);
xnor U13362 (N_13362,N_11158,N_11755);
or U13363 (N_13363,N_10556,N_11881);
nand U13364 (N_13364,N_11755,N_11489);
xnor U13365 (N_13365,N_10091,N_11525);
xor U13366 (N_13366,N_10732,N_10625);
nand U13367 (N_13367,N_11858,N_11137);
and U13368 (N_13368,N_10827,N_10512);
xor U13369 (N_13369,N_10137,N_10430);
or U13370 (N_13370,N_11784,N_10330);
xor U13371 (N_13371,N_11389,N_10758);
xor U13372 (N_13372,N_10546,N_11699);
and U13373 (N_13373,N_11108,N_10297);
nor U13374 (N_13374,N_11683,N_10262);
and U13375 (N_13375,N_11697,N_10589);
nand U13376 (N_13376,N_10784,N_10425);
nor U13377 (N_13377,N_11790,N_11104);
nand U13378 (N_13378,N_10160,N_11576);
and U13379 (N_13379,N_11952,N_11761);
and U13380 (N_13380,N_11074,N_11211);
nand U13381 (N_13381,N_10640,N_11309);
and U13382 (N_13382,N_10225,N_10214);
nor U13383 (N_13383,N_10975,N_11850);
and U13384 (N_13384,N_10678,N_11907);
nor U13385 (N_13385,N_10151,N_11237);
and U13386 (N_13386,N_11581,N_11318);
nand U13387 (N_13387,N_10291,N_10426);
and U13388 (N_13388,N_11352,N_10557);
nand U13389 (N_13389,N_11109,N_10299);
nand U13390 (N_13390,N_10245,N_11915);
or U13391 (N_13391,N_10556,N_10852);
nand U13392 (N_13392,N_11567,N_11256);
nand U13393 (N_13393,N_10336,N_10747);
xor U13394 (N_13394,N_10182,N_10739);
or U13395 (N_13395,N_11261,N_10222);
or U13396 (N_13396,N_11636,N_10025);
and U13397 (N_13397,N_10457,N_11689);
nand U13398 (N_13398,N_10326,N_10339);
or U13399 (N_13399,N_11598,N_11512);
nor U13400 (N_13400,N_10639,N_11620);
and U13401 (N_13401,N_11694,N_11313);
and U13402 (N_13402,N_11907,N_10674);
nand U13403 (N_13403,N_11126,N_11654);
nor U13404 (N_13404,N_11394,N_10119);
and U13405 (N_13405,N_10097,N_10867);
or U13406 (N_13406,N_11211,N_10051);
and U13407 (N_13407,N_10400,N_11115);
or U13408 (N_13408,N_10800,N_10592);
xor U13409 (N_13409,N_10707,N_11128);
nand U13410 (N_13410,N_11168,N_10222);
or U13411 (N_13411,N_11719,N_10463);
nor U13412 (N_13412,N_11265,N_10743);
and U13413 (N_13413,N_10238,N_11062);
nor U13414 (N_13414,N_10188,N_11033);
xor U13415 (N_13415,N_11682,N_11459);
xnor U13416 (N_13416,N_10156,N_11942);
xnor U13417 (N_13417,N_10823,N_11301);
xor U13418 (N_13418,N_10314,N_10607);
or U13419 (N_13419,N_11337,N_11409);
and U13420 (N_13420,N_11021,N_10942);
or U13421 (N_13421,N_10370,N_11876);
nand U13422 (N_13422,N_11272,N_10381);
or U13423 (N_13423,N_10516,N_10634);
or U13424 (N_13424,N_11720,N_10488);
and U13425 (N_13425,N_11215,N_11445);
nand U13426 (N_13426,N_11354,N_11322);
and U13427 (N_13427,N_11003,N_10787);
xnor U13428 (N_13428,N_11267,N_10559);
and U13429 (N_13429,N_11782,N_10241);
xor U13430 (N_13430,N_11646,N_10043);
xnor U13431 (N_13431,N_11302,N_11305);
nand U13432 (N_13432,N_10575,N_10794);
nand U13433 (N_13433,N_10199,N_10489);
nand U13434 (N_13434,N_10916,N_11862);
or U13435 (N_13435,N_10508,N_10015);
xnor U13436 (N_13436,N_11138,N_10715);
or U13437 (N_13437,N_11060,N_11588);
and U13438 (N_13438,N_11212,N_11335);
and U13439 (N_13439,N_11298,N_10626);
or U13440 (N_13440,N_11829,N_11987);
nor U13441 (N_13441,N_10000,N_10262);
or U13442 (N_13442,N_10305,N_10710);
or U13443 (N_13443,N_11648,N_10654);
and U13444 (N_13444,N_11343,N_11783);
and U13445 (N_13445,N_10960,N_10041);
xor U13446 (N_13446,N_11737,N_10381);
or U13447 (N_13447,N_10795,N_11315);
nand U13448 (N_13448,N_10974,N_10507);
nor U13449 (N_13449,N_10882,N_10395);
xor U13450 (N_13450,N_10439,N_11305);
nand U13451 (N_13451,N_10925,N_10881);
and U13452 (N_13452,N_10420,N_10678);
nand U13453 (N_13453,N_11686,N_10989);
nand U13454 (N_13454,N_10594,N_10936);
and U13455 (N_13455,N_10672,N_11406);
nor U13456 (N_13456,N_11182,N_10319);
xor U13457 (N_13457,N_11779,N_11407);
or U13458 (N_13458,N_10896,N_10974);
and U13459 (N_13459,N_10102,N_10551);
xor U13460 (N_13460,N_11778,N_10722);
nand U13461 (N_13461,N_11450,N_10446);
nor U13462 (N_13462,N_11050,N_10191);
nor U13463 (N_13463,N_11338,N_11260);
and U13464 (N_13464,N_11091,N_11417);
nor U13465 (N_13465,N_10340,N_10194);
or U13466 (N_13466,N_10131,N_10529);
or U13467 (N_13467,N_11176,N_11469);
nand U13468 (N_13468,N_10721,N_10821);
or U13469 (N_13469,N_10866,N_10409);
nor U13470 (N_13470,N_10897,N_10183);
and U13471 (N_13471,N_10500,N_10547);
and U13472 (N_13472,N_10756,N_11276);
or U13473 (N_13473,N_10652,N_11720);
nor U13474 (N_13474,N_10713,N_10232);
and U13475 (N_13475,N_11245,N_10800);
and U13476 (N_13476,N_11480,N_11613);
xnor U13477 (N_13477,N_10236,N_11172);
nand U13478 (N_13478,N_10906,N_11487);
or U13479 (N_13479,N_10448,N_11036);
or U13480 (N_13480,N_11772,N_10073);
and U13481 (N_13481,N_10202,N_10042);
nor U13482 (N_13482,N_10306,N_11801);
xor U13483 (N_13483,N_10272,N_11300);
nor U13484 (N_13484,N_10322,N_10693);
nor U13485 (N_13485,N_11161,N_11257);
nor U13486 (N_13486,N_10745,N_11618);
nor U13487 (N_13487,N_11019,N_10485);
nor U13488 (N_13488,N_11854,N_11295);
nand U13489 (N_13489,N_11038,N_11506);
nor U13490 (N_13490,N_10033,N_10203);
and U13491 (N_13491,N_10602,N_10335);
nor U13492 (N_13492,N_11153,N_10100);
xnor U13493 (N_13493,N_11716,N_11902);
and U13494 (N_13494,N_10293,N_11567);
and U13495 (N_13495,N_11870,N_10830);
nand U13496 (N_13496,N_11430,N_11970);
nor U13497 (N_13497,N_11756,N_10813);
and U13498 (N_13498,N_11302,N_11814);
and U13499 (N_13499,N_10327,N_11602);
xnor U13500 (N_13500,N_10695,N_10849);
nor U13501 (N_13501,N_10667,N_10540);
nand U13502 (N_13502,N_11756,N_10301);
xor U13503 (N_13503,N_10604,N_11300);
nand U13504 (N_13504,N_11819,N_11228);
or U13505 (N_13505,N_11224,N_11062);
and U13506 (N_13506,N_10334,N_10082);
or U13507 (N_13507,N_10623,N_11975);
or U13508 (N_13508,N_11844,N_11662);
or U13509 (N_13509,N_11974,N_10544);
xor U13510 (N_13510,N_10772,N_10223);
xor U13511 (N_13511,N_11682,N_10711);
and U13512 (N_13512,N_10810,N_10376);
nor U13513 (N_13513,N_11319,N_11386);
and U13514 (N_13514,N_11496,N_10013);
xor U13515 (N_13515,N_11378,N_11787);
nor U13516 (N_13516,N_10291,N_10308);
nand U13517 (N_13517,N_10791,N_11330);
and U13518 (N_13518,N_10272,N_10490);
or U13519 (N_13519,N_10551,N_10990);
and U13520 (N_13520,N_11110,N_11224);
or U13521 (N_13521,N_11913,N_11124);
nand U13522 (N_13522,N_11998,N_11500);
xor U13523 (N_13523,N_10365,N_11127);
nor U13524 (N_13524,N_10979,N_10020);
xnor U13525 (N_13525,N_11009,N_10083);
nor U13526 (N_13526,N_10006,N_10956);
nand U13527 (N_13527,N_11926,N_10111);
xnor U13528 (N_13528,N_11356,N_10299);
and U13529 (N_13529,N_11602,N_11962);
nor U13530 (N_13530,N_11998,N_10945);
nor U13531 (N_13531,N_11885,N_11540);
or U13532 (N_13532,N_11223,N_11637);
or U13533 (N_13533,N_11951,N_11121);
or U13534 (N_13534,N_10904,N_10560);
or U13535 (N_13535,N_11872,N_11358);
xor U13536 (N_13536,N_11653,N_10881);
xnor U13537 (N_13537,N_11245,N_11533);
xnor U13538 (N_13538,N_11922,N_10246);
and U13539 (N_13539,N_10369,N_11553);
and U13540 (N_13540,N_10384,N_10841);
nand U13541 (N_13541,N_10643,N_10866);
nor U13542 (N_13542,N_10007,N_10611);
or U13543 (N_13543,N_11325,N_11405);
or U13544 (N_13544,N_11571,N_10627);
nor U13545 (N_13545,N_11055,N_10276);
or U13546 (N_13546,N_11216,N_10562);
nand U13547 (N_13547,N_11719,N_10444);
nand U13548 (N_13548,N_11388,N_11410);
nor U13549 (N_13549,N_10482,N_10869);
nor U13550 (N_13550,N_11153,N_10079);
nor U13551 (N_13551,N_11053,N_11342);
and U13552 (N_13552,N_11022,N_11245);
and U13553 (N_13553,N_11766,N_11445);
and U13554 (N_13554,N_11589,N_11123);
and U13555 (N_13555,N_10477,N_10188);
xnor U13556 (N_13556,N_11091,N_11107);
nand U13557 (N_13557,N_11881,N_11235);
and U13558 (N_13558,N_11693,N_10828);
nor U13559 (N_13559,N_11763,N_10127);
nor U13560 (N_13560,N_10903,N_11177);
nor U13561 (N_13561,N_10441,N_11499);
or U13562 (N_13562,N_11165,N_11657);
and U13563 (N_13563,N_10612,N_10471);
xnor U13564 (N_13564,N_10075,N_10671);
or U13565 (N_13565,N_11836,N_11642);
nand U13566 (N_13566,N_11189,N_10596);
nor U13567 (N_13567,N_10447,N_10808);
nor U13568 (N_13568,N_11155,N_11711);
nand U13569 (N_13569,N_11333,N_11221);
nor U13570 (N_13570,N_11888,N_11036);
xor U13571 (N_13571,N_10223,N_11428);
xor U13572 (N_13572,N_11995,N_10949);
xor U13573 (N_13573,N_11691,N_11229);
xnor U13574 (N_13574,N_10092,N_10732);
nand U13575 (N_13575,N_11526,N_10502);
and U13576 (N_13576,N_10818,N_11442);
xor U13577 (N_13577,N_10862,N_10323);
and U13578 (N_13578,N_11751,N_10199);
xor U13579 (N_13579,N_10014,N_11614);
or U13580 (N_13580,N_11942,N_10282);
or U13581 (N_13581,N_11032,N_10674);
nor U13582 (N_13582,N_11123,N_10473);
nor U13583 (N_13583,N_10534,N_11279);
xor U13584 (N_13584,N_11827,N_11929);
nor U13585 (N_13585,N_11025,N_10348);
and U13586 (N_13586,N_11424,N_11532);
xnor U13587 (N_13587,N_10309,N_10925);
or U13588 (N_13588,N_10677,N_11330);
and U13589 (N_13589,N_10997,N_10621);
and U13590 (N_13590,N_11303,N_10449);
nor U13591 (N_13591,N_10969,N_10088);
nor U13592 (N_13592,N_10772,N_10403);
and U13593 (N_13593,N_11362,N_10966);
or U13594 (N_13594,N_10745,N_11020);
xnor U13595 (N_13595,N_11570,N_11741);
nand U13596 (N_13596,N_10022,N_11530);
nor U13597 (N_13597,N_11516,N_11811);
xor U13598 (N_13598,N_11346,N_11997);
or U13599 (N_13599,N_11021,N_10814);
nand U13600 (N_13600,N_11618,N_11204);
nor U13601 (N_13601,N_11938,N_11861);
nand U13602 (N_13602,N_10264,N_10094);
xnor U13603 (N_13603,N_10130,N_10888);
nor U13604 (N_13604,N_11133,N_11248);
and U13605 (N_13605,N_10215,N_10445);
and U13606 (N_13606,N_11888,N_11445);
nor U13607 (N_13607,N_10748,N_10692);
nand U13608 (N_13608,N_10860,N_10343);
and U13609 (N_13609,N_11978,N_10102);
and U13610 (N_13610,N_10708,N_11223);
nor U13611 (N_13611,N_11016,N_10078);
or U13612 (N_13612,N_11947,N_10780);
or U13613 (N_13613,N_10851,N_11923);
or U13614 (N_13614,N_11587,N_10331);
nor U13615 (N_13615,N_11935,N_10653);
and U13616 (N_13616,N_11305,N_11015);
xnor U13617 (N_13617,N_11124,N_11990);
or U13618 (N_13618,N_11909,N_10361);
and U13619 (N_13619,N_11048,N_11015);
and U13620 (N_13620,N_10127,N_10641);
nand U13621 (N_13621,N_11875,N_10555);
xnor U13622 (N_13622,N_11138,N_11942);
or U13623 (N_13623,N_10040,N_10825);
nor U13624 (N_13624,N_10359,N_10215);
and U13625 (N_13625,N_11726,N_10223);
xnor U13626 (N_13626,N_10107,N_10947);
nor U13627 (N_13627,N_11475,N_10770);
xnor U13628 (N_13628,N_10280,N_11486);
or U13629 (N_13629,N_10468,N_11601);
xor U13630 (N_13630,N_11140,N_10339);
xnor U13631 (N_13631,N_10709,N_10276);
or U13632 (N_13632,N_10518,N_10838);
xor U13633 (N_13633,N_10914,N_10079);
or U13634 (N_13634,N_11771,N_11071);
nand U13635 (N_13635,N_11834,N_11234);
nand U13636 (N_13636,N_11720,N_11826);
nand U13637 (N_13637,N_11403,N_10245);
or U13638 (N_13638,N_11498,N_11039);
nor U13639 (N_13639,N_10283,N_10720);
xor U13640 (N_13640,N_11792,N_11420);
nor U13641 (N_13641,N_11300,N_11690);
and U13642 (N_13642,N_11366,N_11972);
or U13643 (N_13643,N_10304,N_10414);
and U13644 (N_13644,N_10724,N_11810);
nand U13645 (N_13645,N_11431,N_10038);
nand U13646 (N_13646,N_10257,N_11196);
xor U13647 (N_13647,N_10311,N_10604);
nor U13648 (N_13648,N_10787,N_11845);
xor U13649 (N_13649,N_11244,N_11628);
and U13650 (N_13650,N_11360,N_11417);
nand U13651 (N_13651,N_10785,N_11465);
nand U13652 (N_13652,N_10524,N_11084);
xor U13653 (N_13653,N_11518,N_10575);
nor U13654 (N_13654,N_11607,N_10138);
nand U13655 (N_13655,N_10695,N_11653);
nor U13656 (N_13656,N_11626,N_11863);
and U13657 (N_13657,N_10366,N_11966);
and U13658 (N_13658,N_10767,N_10609);
nand U13659 (N_13659,N_10879,N_11182);
xor U13660 (N_13660,N_11494,N_10155);
xor U13661 (N_13661,N_11298,N_11811);
nor U13662 (N_13662,N_10785,N_10854);
nor U13663 (N_13663,N_10250,N_11925);
nor U13664 (N_13664,N_11364,N_11864);
nor U13665 (N_13665,N_10453,N_10199);
nor U13666 (N_13666,N_10621,N_10242);
xnor U13667 (N_13667,N_11494,N_10906);
and U13668 (N_13668,N_10065,N_10450);
and U13669 (N_13669,N_10573,N_10858);
xor U13670 (N_13670,N_10357,N_10889);
or U13671 (N_13671,N_10999,N_10662);
xor U13672 (N_13672,N_11572,N_10648);
nor U13673 (N_13673,N_10951,N_10945);
and U13674 (N_13674,N_10835,N_10748);
xor U13675 (N_13675,N_10544,N_10988);
nand U13676 (N_13676,N_11482,N_10725);
or U13677 (N_13677,N_11114,N_10429);
nor U13678 (N_13678,N_11178,N_10826);
nor U13679 (N_13679,N_10902,N_11331);
xor U13680 (N_13680,N_10306,N_10394);
nor U13681 (N_13681,N_10979,N_11476);
and U13682 (N_13682,N_11575,N_10185);
nor U13683 (N_13683,N_11343,N_11821);
nor U13684 (N_13684,N_10898,N_11994);
xor U13685 (N_13685,N_10678,N_10156);
nand U13686 (N_13686,N_10654,N_10738);
nand U13687 (N_13687,N_10902,N_10615);
nand U13688 (N_13688,N_11979,N_10977);
or U13689 (N_13689,N_10119,N_11205);
xor U13690 (N_13690,N_11936,N_11718);
nor U13691 (N_13691,N_11177,N_10627);
or U13692 (N_13692,N_11398,N_11939);
xor U13693 (N_13693,N_10731,N_10167);
and U13694 (N_13694,N_11704,N_10822);
nand U13695 (N_13695,N_10327,N_11386);
and U13696 (N_13696,N_11908,N_10444);
nand U13697 (N_13697,N_10547,N_11573);
and U13698 (N_13698,N_11808,N_10287);
nor U13699 (N_13699,N_10650,N_11726);
xor U13700 (N_13700,N_10332,N_11024);
or U13701 (N_13701,N_10862,N_11310);
and U13702 (N_13702,N_11537,N_11212);
nor U13703 (N_13703,N_10584,N_10288);
and U13704 (N_13704,N_10524,N_11489);
nand U13705 (N_13705,N_11378,N_10394);
nor U13706 (N_13706,N_11670,N_11768);
and U13707 (N_13707,N_11663,N_10864);
or U13708 (N_13708,N_11578,N_10224);
and U13709 (N_13709,N_11142,N_10387);
and U13710 (N_13710,N_10298,N_11322);
and U13711 (N_13711,N_11319,N_10434);
xor U13712 (N_13712,N_11114,N_11536);
xnor U13713 (N_13713,N_10057,N_10881);
nor U13714 (N_13714,N_10348,N_11401);
xor U13715 (N_13715,N_11974,N_10803);
nor U13716 (N_13716,N_11858,N_10241);
nor U13717 (N_13717,N_11777,N_10884);
nand U13718 (N_13718,N_11475,N_10864);
and U13719 (N_13719,N_11792,N_11619);
and U13720 (N_13720,N_10066,N_11139);
and U13721 (N_13721,N_11019,N_11651);
nor U13722 (N_13722,N_11071,N_11851);
xor U13723 (N_13723,N_10274,N_11833);
nor U13724 (N_13724,N_11841,N_10350);
xnor U13725 (N_13725,N_10878,N_10693);
or U13726 (N_13726,N_11032,N_10757);
xnor U13727 (N_13727,N_10148,N_11301);
and U13728 (N_13728,N_10603,N_10100);
nor U13729 (N_13729,N_11531,N_11893);
xor U13730 (N_13730,N_10958,N_10027);
nand U13731 (N_13731,N_11771,N_11504);
and U13732 (N_13732,N_11129,N_11387);
nand U13733 (N_13733,N_11214,N_10572);
and U13734 (N_13734,N_10295,N_11064);
nand U13735 (N_13735,N_11587,N_10272);
xnor U13736 (N_13736,N_11625,N_11924);
and U13737 (N_13737,N_10357,N_11204);
nor U13738 (N_13738,N_10991,N_10955);
xnor U13739 (N_13739,N_10888,N_10481);
nand U13740 (N_13740,N_10721,N_11931);
or U13741 (N_13741,N_10777,N_10690);
xnor U13742 (N_13742,N_10932,N_10915);
nand U13743 (N_13743,N_10232,N_10346);
nand U13744 (N_13744,N_10366,N_10021);
or U13745 (N_13745,N_11554,N_10871);
and U13746 (N_13746,N_11190,N_11547);
nand U13747 (N_13747,N_11532,N_11158);
or U13748 (N_13748,N_10930,N_10745);
and U13749 (N_13749,N_11237,N_10499);
and U13750 (N_13750,N_10355,N_11602);
nand U13751 (N_13751,N_11140,N_10437);
nor U13752 (N_13752,N_11059,N_11530);
xor U13753 (N_13753,N_11976,N_11411);
or U13754 (N_13754,N_10794,N_11802);
and U13755 (N_13755,N_10716,N_10986);
xor U13756 (N_13756,N_11508,N_10176);
or U13757 (N_13757,N_11600,N_10025);
or U13758 (N_13758,N_10410,N_11928);
xnor U13759 (N_13759,N_10974,N_10919);
nor U13760 (N_13760,N_11149,N_11542);
xor U13761 (N_13761,N_10014,N_10027);
nor U13762 (N_13762,N_11512,N_10024);
xnor U13763 (N_13763,N_10767,N_11338);
xnor U13764 (N_13764,N_11200,N_11354);
nand U13765 (N_13765,N_10766,N_10892);
or U13766 (N_13766,N_11026,N_11170);
or U13767 (N_13767,N_11349,N_10427);
and U13768 (N_13768,N_10029,N_10625);
nand U13769 (N_13769,N_10349,N_11839);
and U13770 (N_13770,N_10050,N_10310);
xnor U13771 (N_13771,N_11902,N_10434);
or U13772 (N_13772,N_11411,N_11290);
or U13773 (N_13773,N_10246,N_11897);
nor U13774 (N_13774,N_11438,N_11152);
nand U13775 (N_13775,N_10762,N_11331);
or U13776 (N_13776,N_11456,N_11963);
xnor U13777 (N_13777,N_10764,N_10816);
and U13778 (N_13778,N_11656,N_10532);
or U13779 (N_13779,N_11681,N_10527);
and U13780 (N_13780,N_11462,N_10198);
or U13781 (N_13781,N_10214,N_10409);
nand U13782 (N_13782,N_10393,N_10774);
nor U13783 (N_13783,N_11991,N_11843);
and U13784 (N_13784,N_10467,N_11863);
nor U13785 (N_13785,N_10716,N_11153);
and U13786 (N_13786,N_11064,N_11668);
nand U13787 (N_13787,N_11928,N_11444);
nand U13788 (N_13788,N_11469,N_10005);
nor U13789 (N_13789,N_11168,N_11874);
nor U13790 (N_13790,N_10244,N_11953);
nand U13791 (N_13791,N_11729,N_11563);
nand U13792 (N_13792,N_10070,N_11550);
nor U13793 (N_13793,N_11844,N_11590);
or U13794 (N_13794,N_11224,N_11734);
or U13795 (N_13795,N_11729,N_11295);
and U13796 (N_13796,N_10998,N_11360);
or U13797 (N_13797,N_10370,N_11177);
xnor U13798 (N_13798,N_11087,N_11541);
and U13799 (N_13799,N_11177,N_11975);
and U13800 (N_13800,N_10059,N_10154);
nor U13801 (N_13801,N_10692,N_11747);
and U13802 (N_13802,N_11692,N_11803);
and U13803 (N_13803,N_11539,N_11608);
nor U13804 (N_13804,N_10711,N_10508);
or U13805 (N_13805,N_11186,N_11684);
or U13806 (N_13806,N_11256,N_11110);
or U13807 (N_13807,N_10780,N_10018);
nand U13808 (N_13808,N_11632,N_10913);
nor U13809 (N_13809,N_10617,N_11197);
xor U13810 (N_13810,N_11435,N_11497);
nor U13811 (N_13811,N_11198,N_10158);
or U13812 (N_13812,N_11703,N_10365);
or U13813 (N_13813,N_10902,N_10479);
and U13814 (N_13814,N_10484,N_10470);
xor U13815 (N_13815,N_10637,N_11331);
or U13816 (N_13816,N_11936,N_11852);
nand U13817 (N_13817,N_11631,N_10772);
nor U13818 (N_13818,N_11111,N_11663);
or U13819 (N_13819,N_11083,N_11098);
xor U13820 (N_13820,N_10833,N_11086);
xor U13821 (N_13821,N_10394,N_11173);
xnor U13822 (N_13822,N_11906,N_11903);
nand U13823 (N_13823,N_11339,N_10306);
xnor U13824 (N_13824,N_11817,N_10744);
and U13825 (N_13825,N_11701,N_11795);
nand U13826 (N_13826,N_10278,N_11838);
nand U13827 (N_13827,N_10591,N_11330);
nor U13828 (N_13828,N_11338,N_10215);
or U13829 (N_13829,N_11047,N_10637);
nand U13830 (N_13830,N_10845,N_10677);
or U13831 (N_13831,N_10543,N_10952);
nor U13832 (N_13832,N_10560,N_11298);
and U13833 (N_13833,N_11299,N_10563);
and U13834 (N_13834,N_11577,N_10576);
and U13835 (N_13835,N_10115,N_11938);
and U13836 (N_13836,N_11070,N_11111);
nor U13837 (N_13837,N_10818,N_11408);
nor U13838 (N_13838,N_10248,N_11745);
nand U13839 (N_13839,N_10551,N_10614);
or U13840 (N_13840,N_11001,N_10878);
and U13841 (N_13841,N_10799,N_10784);
and U13842 (N_13842,N_10189,N_11619);
nand U13843 (N_13843,N_10685,N_11389);
or U13844 (N_13844,N_10308,N_11277);
or U13845 (N_13845,N_10728,N_10189);
nand U13846 (N_13846,N_10095,N_10517);
nor U13847 (N_13847,N_10097,N_11178);
or U13848 (N_13848,N_10317,N_11293);
xor U13849 (N_13849,N_11681,N_11741);
and U13850 (N_13850,N_10842,N_11543);
or U13851 (N_13851,N_11108,N_11289);
xor U13852 (N_13852,N_10844,N_10189);
nand U13853 (N_13853,N_10016,N_10028);
xor U13854 (N_13854,N_11776,N_11659);
xnor U13855 (N_13855,N_10467,N_10298);
xnor U13856 (N_13856,N_10521,N_10633);
nand U13857 (N_13857,N_11971,N_10568);
nand U13858 (N_13858,N_11001,N_11567);
or U13859 (N_13859,N_11692,N_10963);
xnor U13860 (N_13860,N_10084,N_11384);
and U13861 (N_13861,N_10937,N_11673);
xor U13862 (N_13862,N_10086,N_11638);
nor U13863 (N_13863,N_11427,N_11691);
nor U13864 (N_13864,N_10957,N_11478);
xnor U13865 (N_13865,N_11591,N_11283);
nand U13866 (N_13866,N_10156,N_11940);
nand U13867 (N_13867,N_11470,N_10661);
xnor U13868 (N_13868,N_11317,N_10254);
or U13869 (N_13869,N_11137,N_11776);
or U13870 (N_13870,N_10171,N_10673);
nand U13871 (N_13871,N_10927,N_10773);
xor U13872 (N_13872,N_10487,N_10429);
xor U13873 (N_13873,N_11947,N_10602);
nor U13874 (N_13874,N_11455,N_10502);
and U13875 (N_13875,N_10658,N_10282);
or U13876 (N_13876,N_11226,N_11967);
nor U13877 (N_13877,N_11471,N_10616);
xnor U13878 (N_13878,N_11710,N_10071);
xnor U13879 (N_13879,N_10578,N_10940);
or U13880 (N_13880,N_11175,N_11352);
nor U13881 (N_13881,N_10365,N_11692);
xnor U13882 (N_13882,N_11064,N_11175);
and U13883 (N_13883,N_11974,N_11549);
nor U13884 (N_13884,N_11761,N_10114);
and U13885 (N_13885,N_11999,N_11538);
nand U13886 (N_13886,N_10837,N_10878);
nand U13887 (N_13887,N_11893,N_11769);
nand U13888 (N_13888,N_11660,N_11582);
nand U13889 (N_13889,N_11887,N_11665);
or U13890 (N_13890,N_10670,N_10138);
nand U13891 (N_13891,N_10164,N_11094);
and U13892 (N_13892,N_10318,N_11445);
nand U13893 (N_13893,N_10910,N_11763);
or U13894 (N_13894,N_11452,N_10409);
and U13895 (N_13895,N_10642,N_11111);
or U13896 (N_13896,N_10755,N_10255);
or U13897 (N_13897,N_10973,N_11965);
nor U13898 (N_13898,N_10834,N_10049);
nand U13899 (N_13899,N_11622,N_11649);
and U13900 (N_13900,N_11602,N_11650);
and U13901 (N_13901,N_11382,N_11058);
nand U13902 (N_13902,N_10292,N_10102);
and U13903 (N_13903,N_11678,N_11579);
nor U13904 (N_13904,N_11840,N_10106);
nand U13905 (N_13905,N_11514,N_10179);
xor U13906 (N_13906,N_10886,N_11602);
or U13907 (N_13907,N_11806,N_11023);
xor U13908 (N_13908,N_10138,N_11677);
xor U13909 (N_13909,N_11575,N_10641);
or U13910 (N_13910,N_10635,N_10315);
or U13911 (N_13911,N_11332,N_10717);
xnor U13912 (N_13912,N_11929,N_10619);
or U13913 (N_13913,N_11725,N_11559);
or U13914 (N_13914,N_11671,N_10597);
nand U13915 (N_13915,N_10313,N_11775);
xor U13916 (N_13916,N_10800,N_10293);
nand U13917 (N_13917,N_11657,N_10186);
xnor U13918 (N_13918,N_11872,N_10019);
or U13919 (N_13919,N_10052,N_10143);
or U13920 (N_13920,N_11112,N_10946);
or U13921 (N_13921,N_11698,N_10155);
or U13922 (N_13922,N_10450,N_11695);
xor U13923 (N_13923,N_10597,N_11804);
nor U13924 (N_13924,N_11893,N_11971);
nand U13925 (N_13925,N_10377,N_11110);
nand U13926 (N_13926,N_10411,N_10031);
xor U13927 (N_13927,N_11729,N_11474);
nand U13928 (N_13928,N_11653,N_10370);
nor U13929 (N_13929,N_11576,N_11090);
and U13930 (N_13930,N_11041,N_10119);
or U13931 (N_13931,N_11203,N_10268);
nand U13932 (N_13932,N_10144,N_11922);
xnor U13933 (N_13933,N_10479,N_10047);
nand U13934 (N_13934,N_10381,N_10590);
or U13935 (N_13935,N_11230,N_10628);
nor U13936 (N_13936,N_11515,N_11654);
and U13937 (N_13937,N_11711,N_10537);
and U13938 (N_13938,N_10764,N_11920);
xnor U13939 (N_13939,N_10065,N_11144);
nor U13940 (N_13940,N_11416,N_11802);
or U13941 (N_13941,N_11119,N_10832);
xor U13942 (N_13942,N_10631,N_11701);
and U13943 (N_13943,N_10993,N_10114);
and U13944 (N_13944,N_11527,N_10925);
or U13945 (N_13945,N_10288,N_10698);
nand U13946 (N_13946,N_11126,N_11990);
or U13947 (N_13947,N_11417,N_10507);
xor U13948 (N_13948,N_11635,N_11282);
nor U13949 (N_13949,N_11572,N_10910);
and U13950 (N_13950,N_10774,N_10112);
nand U13951 (N_13951,N_10531,N_11410);
and U13952 (N_13952,N_10065,N_10806);
nand U13953 (N_13953,N_11153,N_11084);
or U13954 (N_13954,N_10254,N_11498);
xnor U13955 (N_13955,N_11026,N_10907);
and U13956 (N_13956,N_10251,N_10053);
or U13957 (N_13957,N_10075,N_11893);
or U13958 (N_13958,N_11137,N_10668);
xor U13959 (N_13959,N_10123,N_11056);
and U13960 (N_13960,N_10660,N_10290);
or U13961 (N_13961,N_11172,N_10559);
or U13962 (N_13962,N_10246,N_11380);
nor U13963 (N_13963,N_10450,N_10468);
or U13964 (N_13964,N_11780,N_11601);
nor U13965 (N_13965,N_11159,N_11662);
xor U13966 (N_13966,N_11274,N_10362);
nor U13967 (N_13967,N_10907,N_10937);
xor U13968 (N_13968,N_10061,N_11209);
nand U13969 (N_13969,N_10837,N_10081);
and U13970 (N_13970,N_11077,N_10003);
nand U13971 (N_13971,N_10323,N_11648);
and U13972 (N_13972,N_11867,N_11528);
or U13973 (N_13973,N_10657,N_11775);
xor U13974 (N_13974,N_10672,N_10550);
nor U13975 (N_13975,N_10362,N_10215);
xor U13976 (N_13976,N_11051,N_11654);
nor U13977 (N_13977,N_11054,N_11406);
and U13978 (N_13978,N_10685,N_11595);
and U13979 (N_13979,N_11241,N_10761);
and U13980 (N_13980,N_11529,N_10967);
xor U13981 (N_13981,N_11326,N_10496);
or U13982 (N_13982,N_11500,N_10135);
and U13983 (N_13983,N_11074,N_11105);
or U13984 (N_13984,N_10927,N_10647);
nand U13985 (N_13985,N_11920,N_10857);
nand U13986 (N_13986,N_10343,N_11268);
and U13987 (N_13987,N_10868,N_10791);
nor U13988 (N_13988,N_10922,N_11042);
or U13989 (N_13989,N_11213,N_11312);
or U13990 (N_13990,N_10774,N_10925);
and U13991 (N_13991,N_10940,N_10989);
nand U13992 (N_13992,N_10927,N_11468);
nand U13993 (N_13993,N_11467,N_11614);
and U13994 (N_13994,N_10375,N_11926);
xnor U13995 (N_13995,N_10138,N_10360);
nand U13996 (N_13996,N_11659,N_11450);
and U13997 (N_13997,N_10270,N_10441);
or U13998 (N_13998,N_10951,N_11092);
xnor U13999 (N_13999,N_10458,N_10957);
nor U14000 (N_14000,N_12552,N_13170);
xor U14001 (N_14001,N_13627,N_13757);
xor U14002 (N_14002,N_13264,N_12027);
xor U14003 (N_14003,N_12082,N_12952);
nor U14004 (N_14004,N_12957,N_13218);
nor U14005 (N_14005,N_12854,N_13239);
or U14006 (N_14006,N_13310,N_13831);
nor U14007 (N_14007,N_12008,N_12569);
nand U14008 (N_14008,N_12137,N_12014);
xor U14009 (N_14009,N_12403,N_13197);
or U14010 (N_14010,N_12477,N_12271);
nor U14011 (N_14011,N_12523,N_12991);
or U14012 (N_14012,N_12761,N_13464);
nor U14013 (N_14013,N_12908,N_13625);
or U14014 (N_14014,N_12617,N_12055);
and U14015 (N_14015,N_12778,N_12184);
and U14016 (N_14016,N_13914,N_13832);
nor U14017 (N_14017,N_12006,N_12473);
and U14018 (N_14018,N_13650,N_13805);
nand U14019 (N_14019,N_13407,N_13613);
and U14020 (N_14020,N_13038,N_13255);
or U14021 (N_14021,N_13814,N_13516);
xnor U14022 (N_14022,N_13003,N_13350);
or U14023 (N_14023,N_12389,N_13697);
nand U14024 (N_14024,N_12507,N_13352);
or U14025 (N_14025,N_13668,N_13039);
xor U14026 (N_14026,N_12576,N_13940);
or U14027 (N_14027,N_13084,N_12423);
nor U14028 (N_14028,N_12465,N_13722);
xnor U14029 (N_14029,N_13124,N_13730);
and U14030 (N_14030,N_13287,N_13172);
nand U14031 (N_14031,N_13027,N_12983);
and U14032 (N_14032,N_12067,N_13185);
xor U14033 (N_14033,N_12489,N_13047);
nand U14034 (N_14034,N_13384,N_13813);
xor U14035 (N_14035,N_13385,N_13376);
and U14036 (N_14036,N_12881,N_12186);
nor U14037 (N_14037,N_12826,N_13508);
or U14038 (N_14038,N_12818,N_12589);
xnor U14039 (N_14039,N_12435,N_12764);
nand U14040 (N_14040,N_13900,N_12798);
or U14041 (N_14041,N_13041,N_12486);
and U14042 (N_14042,N_12412,N_13614);
nand U14043 (N_14043,N_13833,N_12438);
nor U14044 (N_14044,N_13546,N_13168);
and U14045 (N_14045,N_12825,N_13779);
xor U14046 (N_14046,N_12074,N_12125);
or U14047 (N_14047,N_13189,N_12660);
xnor U14048 (N_14048,N_12272,N_12227);
nand U14049 (N_14049,N_12765,N_12087);
and U14050 (N_14050,N_12513,N_13136);
xor U14051 (N_14051,N_13866,N_13817);
and U14052 (N_14052,N_13149,N_12872);
and U14053 (N_14053,N_13856,N_12926);
nand U14054 (N_14054,N_13563,N_12401);
nor U14055 (N_14055,N_12251,N_12340);
nor U14056 (N_14056,N_13782,N_12100);
and U14057 (N_14057,N_12607,N_13683);
nand U14058 (N_14058,N_13277,N_13420);
nand U14059 (N_14059,N_13556,N_13228);
or U14060 (N_14060,N_12715,N_13926);
nand U14061 (N_14061,N_12951,N_12758);
or U14062 (N_14062,N_12682,N_13447);
or U14063 (N_14063,N_12674,N_12322);
or U14064 (N_14064,N_12615,N_13765);
nand U14065 (N_14065,N_12167,N_12541);
nand U14066 (N_14066,N_12418,N_12638);
nand U14067 (N_14067,N_13799,N_12989);
nand U14068 (N_14068,N_12157,N_12153);
nor U14069 (N_14069,N_13225,N_13422);
nand U14070 (N_14070,N_12393,N_13959);
xor U14071 (N_14071,N_13899,N_13303);
xnor U14072 (N_14072,N_13834,N_12981);
and U14073 (N_14073,N_13864,N_12723);
xnor U14074 (N_14074,N_12813,N_12467);
nor U14075 (N_14075,N_13825,N_12429);
nand U14076 (N_14076,N_13948,N_13329);
and U14077 (N_14077,N_12487,N_13800);
xor U14078 (N_14078,N_13358,N_12613);
nand U14079 (N_14079,N_12211,N_12564);
and U14080 (N_14080,N_13934,N_13057);
nor U14081 (N_14081,N_12884,N_13048);
xor U14082 (N_14082,N_12388,N_12573);
and U14083 (N_14083,N_13776,N_12162);
xnor U14084 (N_14084,N_12649,N_13924);
or U14085 (N_14085,N_12598,N_13557);
and U14086 (N_14086,N_12852,N_12591);
nand U14087 (N_14087,N_13160,N_13028);
xor U14088 (N_14088,N_12833,N_12048);
and U14089 (N_14089,N_13290,N_13553);
nor U14090 (N_14090,N_12970,N_13411);
xnor U14091 (N_14091,N_13707,N_13970);
or U14092 (N_14092,N_12959,N_13706);
nand U14093 (N_14093,N_12858,N_12356);
xnor U14094 (N_14094,N_13473,N_12939);
nand U14095 (N_14095,N_12645,N_13316);
nand U14096 (N_14096,N_12695,N_13594);
nand U14097 (N_14097,N_13847,N_13762);
and U14098 (N_14098,N_13087,N_12492);
or U14099 (N_14099,N_13743,N_13714);
nand U14100 (N_14100,N_13001,N_12532);
nor U14101 (N_14101,N_13086,N_13885);
xnor U14102 (N_14102,N_13367,N_12640);
or U14103 (N_14103,N_13210,N_12352);
and U14104 (N_14104,N_12610,N_12309);
nand U14105 (N_14105,N_13512,N_12253);
nor U14106 (N_14106,N_13566,N_13345);
or U14107 (N_14107,N_13861,N_13661);
and U14108 (N_14108,N_13960,N_13285);
or U14109 (N_14109,N_12156,N_13092);
or U14110 (N_14110,N_13849,N_13259);
and U14111 (N_14111,N_12496,N_13432);
and U14112 (N_14112,N_12127,N_13102);
nor U14113 (N_14113,N_13209,N_12815);
and U14114 (N_14114,N_12205,N_12988);
nor U14115 (N_14115,N_13750,N_12197);
or U14116 (N_14116,N_12490,N_12809);
nor U14117 (N_14117,N_13907,N_13731);
nor U14118 (N_14118,N_12897,N_12353);
or U14119 (N_14119,N_13148,N_13443);
nand U14120 (N_14120,N_12287,N_13126);
nor U14121 (N_14121,N_13724,N_13437);
xnor U14122 (N_14122,N_12547,N_13488);
and U14123 (N_14123,N_13682,N_13314);
xnor U14124 (N_14124,N_12775,N_13659);
nand U14125 (N_14125,N_13903,N_13981);
nand U14126 (N_14126,N_12035,N_12779);
nor U14127 (N_14127,N_12023,N_12776);
nor U14128 (N_14128,N_12984,N_12871);
nand U14129 (N_14129,N_12044,N_13158);
or U14130 (N_14130,N_12215,N_12000);
nor U14131 (N_14131,N_13532,N_12196);
nor U14132 (N_14132,N_12380,N_12452);
and U14133 (N_14133,N_12670,N_13754);
nand U14134 (N_14134,N_12973,N_13195);
nor U14135 (N_14135,N_13562,N_12346);
xor U14136 (N_14136,N_13515,N_12129);
xor U14137 (N_14137,N_13662,N_12768);
nor U14138 (N_14138,N_13998,N_13536);
xnor U14139 (N_14139,N_13370,N_13029);
and U14140 (N_14140,N_12505,N_13693);
nand U14141 (N_14141,N_13151,N_13596);
and U14142 (N_14142,N_12150,N_13449);
nor U14143 (N_14143,N_12894,N_13675);
and U14144 (N_14144,N_13603,N_13558);
xor U14145 (N_14145,N_13424,N_13318);
nand U14146 (N_14146,N_12525,N_13839);
or U14147 (N_14147,N_12550,N_13169);
nor U14148 (N_14148,N_12834,N_13263);
nor U14149 (N_14149,N_12941,N_12241);
nand U14150 (N_14150,N_12923,N_13769);
or U14151 (N_14151,N_13579,N_13377);
or U14152 (N_14152,N_12737,N_12354);
xor U14153 (N_14153,N_12134,N_12965);
nand U14154 (N_14154,N_13090,N_13984);
nor U14155 (N_14155,N_12713,N_12302);
xnor U14156 (N_14156,N_13062,N_13685);
or U14157 (N_14157,N_12673,N_13327);
nand U14158 (N_14158,N_12792,N_12998);
nor U14159 (N_14159,N_13236,N_13269);
and U14160 (N_14160,N_12168,N_13286);
and U14161 (N_14161,N_12967,N_13340);
and U14162 (N_14162,N_12126,N_13241);
nor U14163 (N_14163,N_12371,N_13525);
and U14164 (N_14164,N_13419,N_12634);
nor U14165 (N_14165,N_13441,N_13810);
and U14166 (N_14166,N_13284,N_13275);
nor U14167 (N_14167,N_12447,N_13522);
or U14168 (N_14168,N_13671,N_13485);
or U14169 (N_14169,N_12138,N_13906);
nand U14170 (N_14170,N_13881,N_13231);
nand U14171 (N_14171,N_13143,N_12470);
nand U14172 (N_14172,N_13109,N_12052);
xor U14173 (N_14173,N_13439,N_12767);
and U14174 (N_14174,N_12880,N_12118);
nor U14175 (N_14175,N_12549,N_12231);
and U14176 (N_14176,N_13436,N_12772);
and U14177 (N_14177,N_12316,N_12260);
or U14178 (N_14178,N_13063,N_13595);
or U14179 (N_14179,N_13744,N_13409);
or U14180 (N_14180,N_13882,N_13787);
and U14181 (N_14181,N_12814,N_13359);
nand U14182 (N_14182,N_13876,N_12701);
nand U14183 (N_14183,N_12888,N_13381);
and U14184 (N_14184,N_13030,N_12278);
nand U14185 (N_14185,N_13695,N_13728);
xnor U14186 (N_14186,N_13932,N_13356);
xor U14187 (N_14187,N_13667,N_12643);
nand U14188 (N_14188,N_12618,N_13853);
nand U14189 (N_14189,N_13771,N_13949);
or U14190 (N_14190,N_13502,N_13735);
nand U14191 (N_14191,N_13745,N_13630);
nand U14192 (N_14192,N_12805,N_13624);
nor U14193 (N_14193,N_13016,N_13037);
xnor U14194 (N_14194,N_12104,N_13916);
xor U14195 (N_14195,N_12439,N_12720);
or U14196 (N_14196,N_13478,N_13105);
and U14197 (N_14197,N_13338,N_13248);
and U14198 (N_14198,N_12499,N_13908);
and U14199 (N_14199,N_13620,N_12568);
nand U14200 (N_14200,N_12786,N_13936);
or U14201 (N_14201,N_12783,N_13208);
and U14202 (N_14202,N_13397,N_12602);
nand U14203 (N_14203,N_12861,N_12306);
xnor U14204 (N_14204,N_13444,N_12180);
and U14205 (N_14205,N_13590,N_13953);
or U14206 (N_14206,N_13374,N_12025);
and U14207 (N_14207,N_13196,N_13199);
and U14208 (N_14208,N_13872,N_13360);
nand U14209 (N_14209,N_13403,N_12372);
and U14210 (N_14210,N_13788,N_13451);
nor U14211 (N_14211,N_13165,N_12046);
nor U14212 (N_14212,N_13206,N_13687);
xor U14213 (N_14213,N_13322,N_13234);
or U14214 (N_14214,N_12963,N_12259);
or U14215 (N_14215,N_13278,N_12053);
xor U14216 (N_14216,N_13379,N_12577);
or U14217 (N_14217,N_12413,N_13226);
nor U14218 (N_14218,N_12217,N_13487);
and U14219 (N_14219,N_12400,N_12324);
or U14220 (N_14220,N_13989,N_12169);
or U14221 (N_14221,N_13980,N_13611);
or U14222 (N_14222,N_12268,N_13660);
nor U14223 (N_14223,N_12837,N_12007);
and U14224 (N_14224,N_13055,N_13709);
xor U14225 (N_14225,N_12461,N_13104);
xor U14226 (N_14226,N_12684,N_13301);
or U14227 (N_14227,N_13729,N_12173);
xnor U14228 (N_14228,N_13162,N_13511);
and U14229 (N_14229,N_12191,N_12754);
xnor U14230 (N_14230,N_13673,N_13463);
nor U14231 (N_14231,N_13778,N_13163);
and U14232 (N_14232,N_12148,N_13884);
xnor U14233 (N_14233,N_13091,N_12734);
xor U14234 (N_14234,N_13095,N_13636);
nor U14235 (N_14235,N_13588,N_12635);
nor U14236 (N_14236,N_13362,N_13144);
xnor U14237 (N_14237,N_13755,N_12291);
or U14238 (N_14238,N_12182,N_12718);
and U14239 (N_14239,N_13442,N_13066);
or U14240 (N_14240,N_13843,N_12964);
or U14241 (N_14241,N_13772,N_13823);
and U14242 (N_14242,N_12277,N_13404);
nand U14243 (N_14243,N_13581,N_13475);
nand U14244 (N_14244,N_12990,N_12258);
xnor U14245 (N_14245,N_12844,N_12109);
nor U14246 (N_14246,N_13543,N_12903);
nand U14247 (N_14247,N_12263,N_13874);
nor U14248 (N_14248,N_12022,N_12870);
xnor U14249 (N_14249,N_13017,N_12992);
or U14250 (N_14250,N_13368,N_13184);
xor U14251 (N_14251,N_13628,N_13326);
or U14252 (N_14252,N_13455,N_13142);
xor U14253 (N_14253,N_13501,N_12338);
nor U14254 (N_14254,N_13305,N_13240);
and U14255 (N_14255,N_13547,N_12759);
nor U14256 (N_14256,N_13548,N_12476);
nor U14257 (N_14257,N_12917,N_13991);
nand U14258 (N_14258,N_13217,N_13387);
nor U14259 (N_14259,N_13559,N_13561);
nand U14260 (N_14260,N_12319,N_12960);
or U14261 (N_14261,N_12404,N_12948);
nor U14262 (N_14262,N_13068,N_12856);
nand U14263 (N_14263,N_12580,N_12039);
and U14264 (N_14264,N_13749,N_13117);
nand U14265 (N_14265,N_13680,N_13256);
xor U14266 (N_14266,N_13308,N_12971);
xnor U14267 (N_14267,N_12246,N_13394);
or U14268 (N_14268,N_13328,N_12632);
or U14269 (N_14269,N_12214,N_13279);
nor U14270 (N_14270,N_12471,N_13646);
and U14271 (N_14271,N_13270,N_12054);
nor U14272 (N_14272,N_12244,N_13032);
nor U14273 (N_14273,N_13760,N_12658);
and U14274 (N_14274,N_13111,N_12453);
and U14275 (N_14275,N_12079,N_13317);
nand U14276 (N_14276,N_13053,N_12112);
nor U14277 (N_14277,N_12807,N_12842);
nor U14278 (N_14278,N_12629,N_12620);
and U14279 (N_14279,N_13759,N_12974);
nand U14280 (N_14280,N_13229,N_12832);
nor U14281 (N_14281,N_13615,N_12245);
nor U14282 (N_14282,N_12528,N_12869);
xor U14283 (N_14283,N_12347,N_12364);
and U14284 (N_14284,N_12822,N_13012);
nor U14285 (N_14285,N_12510,N_12501);
nand U14286 (N_14286,N_12793,N_12683);
xnor U14287 (N_14287,N_13058,N_12828);
and U14288 (N_14288,N_12811,N_12284);
and U14289 (N_14289,N_12017,N_12124);
xor U14290 (N_14290,N_13325,N_12459);
nor U14291 (N_14291,N_12774,N_13577);
or U14292 (N_14292,N_13232,N_13933);
nand U14293 (N_14293,N_13167,N_13986);
or U14294 (N_14294,N_13828,N_12075);
or U14295 (N_14295,N_12266,N_12226);
nor U14296 (N_14296,N_12751,N_13097);
xor U14297 (N_14297,N_12582,N_13587);
and U14298 (N_14298,N_12120,N_12557);
xor U14299 (N_14299,N_13205,N_12804);
or U14300 (N_14300,N_12213,N_12599);
and U14301 (N_14301,N_12147,N_12097);
and U14302 (N_14302,N_13253,N_12175);
nor U14303 (N_14303,N_13602,N_13023);
nand U14304 (N_14304,N_13584,N_12614);
nor U14305 (N_14305,N_12891,N_12474);
nor U14306 (N_14306,N_13353,N_13664);
and U14307 (N_14307,N_12010,N_13835);
xnor U14308 (N_14308,N_12920,N_12940);
or U14309 (N_14309,N_12061,N_12427);
nand U14310 (N_14310,N_13483,N_12066);
nor U14311 (N_14311,N_13469,N_12788);
and U14312 (N_14312,N_13071,N_13271);
xnor U14313 (N_14313,N_12166,N_13837);
xnor U14314 (N_14314,N_13623,N_12114);
nand U14315 (N_14315,N_13541,N_12093);
nand U14316 (N_14316,N_12367,N_12623);
nand U14317 (N_14317,N_12399,N_12937);
nor U14318 (N_14318,N_12994,N_12575);
nor U14319 (N_14319,N_12567,N_13060);
or U14320 (N_14320,N_12454,N_12921);
and U14321 (N_14321,N_13493,N_13969);
xnor U14322 (N_14322,N_13796,N_13871);
or U14323 (N_14323,N_12616,N_13188);
and U14324 (N_14324,N_13074,N_13434);
nor U14325 (N_14325,N_12374,N_12101);
and U14326 (N_14326,N_13364,N_12236);
and U14327 (N_14327,N_13701,N_13155);
nor U14328 (N_14328,N_13296,N_13747);
or U14329 (N_14329,N_13190,N_12201);
nor U14330 (N_14330,N_13638,N_13334);
nand U14331 (N_14331,N_13363,N_12303);
or U14332 (N_14332,N_13951,N_12030);
nor U14333 (N_14333,N_12139,N_12254);
or U14334 (N_14334,N_12497,N_13486);
nor U14335 (N_14335,N_13246,N_12975);
and U14336 (N_14336,N_12502,N_12270);
and U14337 (N_14337,N_12841,N_13504);
xnor U14338 (N_14338,N_12285,N_12437);
or U14339 (N_14339,N_13178,N_13892);
nand U14340 (N_14340,N_12928,N_13272);
xor U14341 (N_14341,N_13617,N_13803);
and U14342 (N_14342,N_12526,N_12711);
nor U14343 (N_14343,N_12624,N_13101);
nor U14344 (N_14344,N_12790,N_12059);
or U14345 (N_14345,N_12076,N_12504);
and U14346 (N_14346,N_12890,N_12942);
xnor U14347 (N_14347,N_12410,N_13909);
nor U14348 (N_14348,N_13171,N_13224);
nor U14349 (N_14349,N_13950,N_12135);
and U14350 (N_14350,N_12119,N_13372);
and U14351 (N_14351,N_12220,N_12515);
nor U14352 (N_14352,N_13130,N_13077);
or U14353 (N_14353,N_13569,N_13637);
or U14354 (N_14354,N_12334,N_12795);
xor U14355 (N_14355,N_12181,N_13966);
nor U14356 (N_14356,N_12819,N_13069);
or U14357 (N_14357,N_12433,N_13021);
or U14358 (N_14358,N_13257,N_12242);
nor U14359 (N_14359,N_12081,N_13459);
nor U14360 (N_14360,N_12704,N_12559);
nand U14361 (N_14361,N_12801,N_13157);
or U14362 (N_14362,N_13869,N_12177);
nor U14363 (N_14363,N_12938,N_13396);
xor U14364 (N_14364,N_13173,N_12827);
nor U14365 (N_14365,N_12432,N_12899);
or U14366 (N_14366,N_13390,N_12846);
nand U14367 (N_14367,N_12351,N_12460);
and U14368 (N_14368,N_13816,N_12469);
and U14369 (N_14369,N_13770,N_13963);
xnor U14370 (N_14370,N_13156,N_13383);
xnor U14371 (N_14371,N_13652,N_12799);
or U14372 (N_14372,N_13705,N_12672);
nor U14373 (N_14373,N_13321,N_12700);
and U14374 (N_14374,N_12415,N_12847);
xor U14375 (N_14375,N_12015,N_12511);
nor U14376 (N_14376,N_13034,N_13774);
xnor U14377 (N_14377,N_13781,N_13079);
nand U14378 (N_14378,N_13470,N_12738);
and U14379 (N_14379,N_12276,N_13977);
or U14380 (N_14380,N_12561,N_12311);
xnor U14381 (N_14381,N_13975,N_12261);
or U14382 (N_14382,N_13260,N_12685);
nor U14383 (N_14383,N_12900,N_12019);
nor U14384 (N_14384,N_12444,N_13580);
or U14385 (N_14385,N_13369,N_13481);
nand U14386 (N_14386,N_12130,N_13235);
or U14387 (N_14387,N_13465,N_12609);
nand U14388 (N_14388,N_13115,N_12033);
nor U14389 (N_14389,N_12222,N_12235);
or U14390 (N_14390,N_12290,N_13653);
xor U14391 (N_14391,N_12892,N_13050);
nor U14392 (N_14392,N_12517,N_12556);
nor U14393 (N_14393,N_12578,N_12927);
xnor U14394 (N_14394,N_13937,N_12292);
xor U14395 (N_14395,N_13100,N_12202);
nor U14396 (N_14396,N_12835,N_12977);
xor U14397 (N_14397,N_13751,N_12655);
and U14398 (N_14398,N_13604,N_13212);
or U14399 (N_14399,N_12424,N_13133);
and U14400 (N_14400,N_13979,N_13306);
nand U14401 (N_14401,N_12387,N_12233);
or U14402 (N_14402,N_13457,N_13923);
nand U14403 (N_14403,N_12785,N_13642);
and U14404 (N_14404,N_12641,N_12536);
nor U14405 (N_14405,N_12457,N_12397);
nand U14406 (N_14406,N_13738,N_13333);
and U14407 (N_14407,N_13075,N_12028);
and U14408 (N_14408,N_12520,N_13015);
nor U14409 (N_14409,N_13621,N_12651);
or U14410 (N_14410,N_13393,N_12958);
nor U14411 (N_14411,N_12065,N_12430);
and U14412 (N_14412,N_12328,N_12539);
nand U14413 (N_14413,N_12375,N_13417);
or U14414 (N_14414,N_12425,N_13919);
and U14415 (N_14415,N_12771,N_12816);
nor U14416 (N_14416,N_13238,N_12255);
nand U14417 (N_14417,N_12836,N_12831);
xor U14418 (N_14418,N_13179,N_13445);
nor U14419 (N_14419,N_13448,N_13990);
or U14420 (N_14420,N_13768,N_12099);
nor U14421 (N_14421,N_12098,N_13987);
xnor U14422 (N_14422,N_13534,N_13798);
nand U14423 (N_14423,N_13051,N_13789);
nor U14424 (N_14424,N_13955,N_12090);
nand U14425 (N_14425,N_12151,N_12595);
and U14426 (N_14426,N_12553,N_12045);
or U14427 (N_14427,N_12727,N_12735);
or U14428 (N_14428,N_12566,N_12455);
nand U14429 (N_14429,N_12086,N_13361);
or U14430 (N_14430,N_13555,N_12931);
xnor U14431 (N_14431,N_13138,N_12882);
xnor U14432 (N_14432,N_12363,N_12360);
xnor U14433 (N_14433,N_12979,N_13116);
nand U14434 (N_14434,N_12083,N_13262);
or U14435 (N_14435,N_12449,N_12769);
nor U14436 (N_14436,N_13809,N_13720);
and U14437 (N_14437,N_12954,N_13471);
nand U14438 (N_14438,N_12376,N_12810);
xnor U14439 (N_14439,N_13399,N_12601);
and U14440 (N_14440,N_13480,N_12662);
and U14441 (N_14441,N_12312,N_12796);
xor U14442 (N_14442,N_12679,N_12336);
or U14443 (N_14443,N_13826,N_12648);
nand U14444 (N_14444,N_13453,N_12554);
nor U14445 (N_14445,N_12390,N_12043);
nor U14446 (N_14446,N_12203,N_13606);
xnor U14447 (N_14447,N_12442,N_13910);
or U14448 (N_14448,N_13514,N_12584);
and U14449 (N_14449,N_12228,N_12386);
nand U14450 (N_14450,N_13118,N_13713);
xor U14451 (N_14451,N_13461,N_13161);
xor U14452 (N_14452,N_13070,N_13088);
xor U14453 (N_14453,N_13568,N_12910);
nor U14454 (N_14454,N_13025,N_13806);
xnor U14455 (N_14455,N_13413,N_12369);
nand U14456 (N_14456,N_13593,N_12745);
or U14457 (N_14457,N_13635,N_13198);
xor U14458 (N_14458,N_13958,N_12678);
xor U14459 (N_14459,N_13406,N_12560);
and U14460 (N_14460,N_12806,N_13076);
nand U14461 (N_14461,N_12742,N_13295);
or U14462 (N_14462,N_13973,N_12358);
or U14463 (N_14463,N_12110,N_12611);
xor U14464 (N_14464,N_13474,N_13893);
xor U14465 (N_14465,N_12968,N_12495);
xor U14466 (N_14466,N_12705,N_12029);
or U14467 (N_14467,N_12298,N_12732);
or U14468 (N_14468,N_13812,N_12717);
nand U14469 (N_14469,N_13204,N_12187);
or U14470 (N_14470,N_13748,N_12961);
nor U14471 (N_14471,N_13865,N_13503);
nor U14472 (N_14472,N_13657,N_13222);
and U14473 (N_14473,N_12915,N_12391);
or U14474 (N_14474,N_12256,N_12762);
or U14475 (N_14475,N_12483,N_13967);
or U14476 (N_14476,N_13574,N_12283);
and U14477 (N_14477,N_13207,N_12335);
nor U14478 (N_14478,N_12456,N_13438);
or U14479 (N_14479,N_12875,N_12789);
nand U14480 (N_14480,N_13576,N_12172);
xor U14481 (N_14481,N_12144,N_12343);
and U14482 (N_14482,N_12192,N_12250);
nand U14483 (N_14483,N_13446,N_13862);
xor U14484 (N_14484,N_13402,N_12468);
and U14485 (N_14485,N_12216,N_12755);
xor U14486 (N_14486,N_12808,N_12596);
or U14487 (N_14487,N_13018,N_13802);
nor U14488 (N_14488,N_13734,N_13913);
xor U14489 (N_14489,N_13479,N_13073);
and U14490 (N_14490,N_13978,N_13227);
xnor U14491 (N_14491,N_13309,N_12026);
xnor U14492 (N_14492,N_12514,N_13656);
and U14493 (N_14493,N_13887,N_13388);
nand U14494 (N_14494,N_12855,N_12773);
or U14495 (N_14495,N_13996,N_12587);
or U14496 (N_14496,N_12031,N_13941);
nand U14497 (N_14497,N_13716,N_12563);
or U14498 (N_14498,N_13182,N_13678);
or U14499 (N_14499,N_12003,N_12555);
nor U14500 (N_14500,N_13992,N_12995);
or U14501 (N_14501,N_12543,N_13242);
or U14502 (N_14502,N_12896,N_12188);
xor U14503 (N_14503,N_12791,N_13009);
or U14504 (N_14504,N_13840,N_12190);
and U14505 (N_14505,N_12725,N_13676);
nand U14506 (N_14506,N_12094,N_13575);
or U14507 (N_14507,N_12441,N_13049);
xor U14508 (N_14508,N_12350,N_13103);
xnor U14509 (N_14509,N_12262,N_12274);
nor U14510 (N_14510,N_13431,N_13582);
nor U14511 (N_14511,N_12307,N_13120);
or U14512 (N_14512,N_12508,N_13727);
xnor U14513 (N_14513,N_13052,N_13067);
nor U14514 (N_14514,N_13993,N_13495);
xnor U14515 (N_14515,N_12491,N_12247);
xor U14516 (N_14516,N_13107,N_13761);
and U14517 (N_14517,N_13597,N_12056);
xor U14518 (N_14518,N_13551,N_13943);
or U14519 (N_14519,N_12264,N_12361);
nor U14520 (N_14520,N_12020,N_12102);
and U14521 (N_14521,N_12428,N_13690);
nor U14522 (N_14522,N_12451,N_13140);
or U14523 (N_14523,N_13509,N_13297);
nand U14524 (N_14524,N_13544,N_13154);
and U14525 (N_14525,N_13616,N_13550);
and U14526 (N_14526,N_13065,N_12434);
nand U14527 (N_14527,N_12506,N_12238);
and U14528 (N_14528,N_13392,N_13791);
nor U14529 (N_14529,N_12096,N_13570);
or U14530 (N_14530,N_13332,N_13790);
nor U14531 (N_14531,N_12295,N_13150);
or U14532 (N_14532,N_12657,N_12867);
nand U14533 (N_14533,N_12357,N_12402);
nand U14534 (N_14534,N_13000,N_12654);
or U14535 (N_14535,N_13530,N_13098);
nor U14536 (N_14536,N_12650,N_13921);
nor U14537 (N_14537,N_13875,N_12252);
nand U14538 (N_14538,N_13531,N_12699);
and U14539 (N_14539,N_12627,N_12680);
or U14540 (N_14540,N_12189,N_13010);
nor U14541 (N_14541,N_12161,N_13605);
or U14542 (N_14542,N_12812,N_12385);
nand U14543 (N_14543,N_13565,N_12529);
nand U14544 (N_14544,N_13742,N_12746);
or U14545 (N_14545,N_13648,N_13219);
xor U14546 (N_14546,N_13917,N_12605);
and U14547 (N_14547,N_12535,N_12710);
nand U14548 (N_14548,N_13007,N_13510);
and U14549 (N_14549,N_12122,N_13889);
xor U14550 (N_14550,N_13252,N_12071);
nand U14551 (N_14551,N_13035,N_13254);
and U14552 (N_14552,N_12996,N_13527);
nor U14553 (N_14553,N_13677,N_12011);
nand U14554 (N_14554,N_13026,N_13233);
or U14555 (N_14555,N_12558,N_13513);
and U14556 (N_14556,N_12675,N_12078);
or U14557 (N_14557,N_12666,N_12962);
nand U14558 (N_14558,N_12631,N_12411);
nand U14559 (N_14559,N_12207,N_13014);
and U14560 (N_14560,N_12321,N_12794);
nor U14561 (N_14561,N_12628,N_12916);
nor U14562 (N_14562,N_13410,N_12337);
nor U14563 (N_14563,N_13108,N_13780);
nor U14564 (N_14564,N_12275,N_13106);
nor U14565 (N_14565,N_12752,N_12730);
and U14566 (N_14566,N_12637,N_12689);
nor U14567 (N_14567,N_12608,N_13851);
nor U14568 (N_14568,N_13651,N_12953);
or U14569 (N_14569,N_12760,N_13398);
xor U14570 (N_14570,N_13243,N_12527);
nor U14571 (N_14571,N_12694,N_13521);
xor U14572 (N_14572,N_12933,N_12546);
nor U14573 (N_14573,N_12095,N_12945);
and U14574 (N_14574,N_13054,N_13666);
and U14575 (N_14575,N_13291,N_12229);
nand U14576 (N_14576,N_13824,N_13957);
or U14577 (N_14577,N_12712,N_13669);
nand U14578 (N_14578,N_13147,N_12289);
and U14579 (N_14579,N_13412,N_12091);
and U14580 (N_14580,N_13200,N_12034);
xnor U14581 (N_14581,N_13391,N_12571);
or U14582 (N_14582,N_13684,N_12873);
or U14583 (N_14583,N_13346,N_12070);
xor U14584 (N_14584,N_13462,N_12145);
or U14585 (N_14585,N_13099,N_12123);
xor U14586 (N_14586,N_12843,N_12946);
and U14587 (N_14587,N_12901,N_13647);
nor U14588 (N_14588,N_12817,N_12692);
or U14589 (N_14589,N_13783,N_12032);
or U14590 (N_14590,N_13911,N_12422);
xnor U14591 (N_14591,N_12696,N_12784);
nor U14592 (N_14592,N_12885,N_12594);
and U14593 (N_14593,N_13132,N_12728);
nand U14594 (N_14594,N_12905,N_12782);
and U14595 (N_14595,N_12077,N_12665);
or U14596 (N_14596,N_13968,N_13203);
or U14597 (N_14597,N_13583,N_13112);
nor U14598 (N_14598,N_12103,N_13641);
and U14599 (N_14599,N_12002,N_12348);
nand U14600 (N_14600,N_12562,N_12165);
or U14601 (N_14601,N_12279,N_12106);
and U14602 (N_14602,N_13526,N_13804);
nand U14603 (N_14603,N_13489,N_12540);
or U14604 (N_14604,N_12743,N_13859);
or U14605 (N_14605,N_12041,N_13268);
xnor U14606 (N_14606,N_12163,N_13421);
nor U14607 (N_14607,N_12886,N_12204);
and U14608 (N_14608,N_13719,N_13466);
nor U14609 (N_14609,N_13351,N_13046);
nand U14610 (N_14610,N_13873,N_13845);
xnor U14611 (N_14611,N_13922,N_13031);
and U14612 (N_14612,N_13961,N_13573);
and U14613 (N_14613,N_12749,N_13619);
nand U14614 (N_14614,N_13717,N_12141);
or U14615 (N_14615,N_12980,N_12341);
xnor U14616 (N_14616,N_12821,N_12777);
nand U14617 (N_14617,N_13607,N_12382);
or U14618 (N_14618,N_13533,N_12080);
xnor U14619 (N_14619,N_12845,N_12911);
or U14620 (N_14620,N_13213,N_13733);
or U14621 (N_14621,N_12440,N_13808);
or U14622 (N_14622,N_13183,N_12331);
and U14623 (N_14623,N_13373,N_13517);
nor U14624 (N_14624,N_12149,N_13863);
or U14625 (N_14625,N_13085,N_12223);
nand U14626 (N_14626,N_12748,N_13128);
nand U14627 (N_14627,N_13794,N_12320);
nor U14628 (N_14628,N_12866,N_13898);
nor U14629 (N_14629,N_13127,N_12972);
nor U14630 (N_14630,N_13786,N_13440);
and U14631 (N_14631,N_12409,N_12999);
xnor U14632 (N_14632,N_12781,N_13891);
nand U14633 (N_14633,N_13042,N_12326);
xnor U14634 (N_14634,N_12195,N_13221);
and U14635 (N_14635,N_12731,N_12132);
nand U14636 (N_14636,N_12060,N_12377);
nand U14637 (N_14637,N_13386,N_12907);
nor U14638 (N_14638,N_13612,N_13732);
xnor U14639 (N_14639,N_13591,N_13610);
or U14640 (N_14640,N_12626,N_13601);
xor U14641 (N_14641,N_13123,N_13758);
or U14642 (N_14642,N_12850,N_13216);
nor U14643 (N_14643,N_13793,N_12072);
nor U14644 (N_14644,N_13423,N_13496);
nor U14645 (N_14645,N_13467,N_12572);
nor U14646 (N_14646,N_12733,N_13930);
nand U14647 (N_14647,N_13726,N_12533);
nand U14648 (N_14648,N_12690,N_13545);
and U14649 (N_14649,N_12860,N_13852);
xor U14650 (N_14650,N_13918,N_12930);
xor U14651 (N_14651,N_12934,N_13059);
xnor U14652 (N_14652,N_13947,N_12542);
and U14653 (N_14653,N_13500,N_12824);
or U14654 (N_14654,N_13159,N_12273);
nor U14655 (N_14655,N_13299,N_13129);
xnor U14656 (N_14656,N_12703,N_13877);
nor U14657 (N_14657,N_12868,N_13846);
nand U14658 (N_14658,N_12327,N_13945);
nand U14659 (N_14659,N_12265,N_12639);
nand U14660 (N_14660,N_13288,N_13245);
xor U14661 (N_14661,N_12978,N_12493);
nor U14662 (N_14662,N_13266,N_13044);
and U14663 (N_14663,N_13304,N_12133);
xor U14664 (N_14664,N_13737,N_13223);
nand U14665 (N_14665,N_12416,N_12392);
xor U14666 (N_14666,N_13330,N_13905);
nand U14667 (N_14667,N_13335,N_13456);
or U14668 (N_14668,N_12741,N_12092);
or U14669 (N_14669,N_12661,N_12500);
nand U14670 (N_14670,N_13006,N_13838);
or U14671 (N_14671,N_13281,N_13498);
xor U14672 (N_14672,N_13460,N_13349);
nor U14673 (N_14673,N_13072,N_12987);
and U14674 (N_14674,N_12368,N_13307);
nand U14675 (N_14675,N_12359,N_13988);
nand U14676 (N_14676,N_12530,N_12448);
xnor U14677 (N_14677,N_13736,N_12301);
nand U14678 (N_14678,N_13371,N_13002);
and U14679 (N_14679,N_13649,N_12398);
xor U14680 (N_14680,N_12294,N_13848);
nor U14681 (N_14681,N_13946,N_13886);
or U14682 (N_14682,N_12068,N_12516);
or U14683 (N_14683,N_12947,N_12714);
and U14684 (N_14684,N_13819,N_12420);
or U14685 (N_14685,N_12859,N_12158);
and U14686 (N_14686,N_12479,N_13880);
xnor U14687 (N_14687,N_13686,N_13801);
nor U14688 (N_14688,N_13764,N_13187);
xnor U14689 (N_14689,N_13401,N_13337);
nor U14690 (N_14690,N_12756,N_13365);
nor U14691 (N_14691,N_12230,N_12706);
nor U14692 (N_14692,N_13965,N_13499);
or U14693 (N_14693,N_12421,N_13815);
nor U14694 (N_14694,N_13939,N_12653);
xor U14695 (N_14695,N_13629,N_13505);
nor U14696 (N_14696,N_13524,N_12944);
nand U14697 (N_14697,N_13249,N_13820);
nor U14698 (N_14698,N_12464,N_12200);
or U14699 (N_14699,N_13691,N_12909);
nor U14700 (N_14700,N_13347,N_12024);
nand U14701 (N_14701,N_13020,N_13490);
or U14702 (N_14702,N_13366,N_12450);
or U14703 (N_14703,N_13867,N_13339);
nor U14704 (N_14704,N_12373,N_12865);
nor U14705 (N_14705,N_13452,N_13643);
xnor U14706 (N_14706,N_12924,N_13740);
and U14707 (N_14707,N_13925,N_13137);
and U14708 (N_14708,N_12224,N_13131);
and U14709 (N_14709,N_13777,N_12823);
xnor U14710 (N_14710,N_13139,N_13520);
xnor U14711 (N_14711,N_12225,N_13818);
xnor U14712 (N_14712,N_13567,N_12113);
and U14713 (N_14713,N_13343,N_12396);
and U14714 (N_14714,N_13430,N_13357);
or U14715 (N_14715,N_13698,N_13191);
nand U14716 (N_14716,N_13718,N_13429);
nand U14717 (N_14717,N_12239,N_13174);
xor U14718 (N_14718,N_13681,N_13537);
and U14719 (N_14719,N_13425,N_12724);
nand U14720 (N_14720,N_12736,N_13592);
xor U14721 (N_14721,N_13497,N_13857);
nor U14722 (N_14722,N_12419,N_13599);
and U14723 (N_14723,N_12179,N_13696);
and U14724 (N_14724,N_12018,N_13145);
and U14725 (N_14725,N_12063,N_13858);
nor U14726 (N_14726,N_13096,N_13176);
nor U14727 (N_14727,N_12538,N_13302);
or U14728 (N_14728,N_12407,N_12709);
nor U14729 (N_14729,N_12379,N_13355);
xnor U14730 (N_14730,N_12604,N_12115);
or U14731 (N_14731,N_12592,N_12729);
xor U14732 (N_14732,N_13135,N_12370);
nor U14733 (N_14733,N_13011,N_13177);
nor U14734 (N_14734,N_13311,N_13983);
and U14735 (N_14735,N_13081,N_12164);
xor U14736 (N_14736,N_13879,N_13324);
and U14737 (N_14737,N_12583,N_12612);
nand U14738 (N_14738,N_13211,N_12128);
and U14739 (N_14739,N_12853,N_13854);
xor U14740 (N_14740,N_13665,N_12698);
or U14741 (N_14741,N_13146,N_13540);
and U14742 (N_14742,N_12719,N_12943);
nor U14743 (N_14743,N_12339,N_13655);
nand U14744 (N_14744,N_13855,N_12686);
nor U14745 (N_14745,N_12606,N_13842);
nor U14746 (N_14746,N_12524,N_13640);
xnor U14747 (N_14747,N_13708,N_12443);
nor U14748 (N_14748,N_12642,N_13894);
nor U14749 (N_14749,N_13632,N_12085);
nand U14750 (N_14750,N_13273,N_12208);
nor U14751 (N_14751,N_12004,N_12155);
and U14752 (N_14752,N_13089,N_12770);
nor U14753 (N_14753,N_12668,N_12062);
and U14754 (N_14754,N_13600,N_13523);
nand U14755 (N_14755,N_12257,N_12544);
nor U14756 (N_14756,N_12089,N_12013);
nor U14757 (N_14757,N_12021,N_12426);
nand U14758 (N_14758,N_13193,N_13114);
or U14759 (N_14759,N_13929,N_12722);
nor U14760 (N_14760,N_13699,N_12647);
xnor U14761 (N_14761,N_12621,N_13920);
xor U14762 (N_14762,N_13942,N_13416);
nand U14763 (N_14763,N_13375,N_13844);
nor U14764 (N_14764,N_13400,N_13040);
and U14765 (N_14765,N_12863,N_13122);
nand U14766 (N_14766,N_13689,N_13672);
nand U14767 (N_14767,N_12744,N_12198);
nand U14768 (N_14768,N_13395,N_13700);
or U14769 (N_14769,N_13415,N_12721);
nand U14770 (N_14770,N_13380,N_12919);
nand U14771 (N_14771,N_12982,N_12600);
or U14772 (N_14772,N_12408,N_13378);
xnor U14773 (N_14773,N_13300,N_13344);
or U14774 (N_14774,N_13045,N_12512);
and U14775 (N_14775,N_12669,N_12154);
nand U14776 (N_14776,N_12677,N_12879);
or U14777 (N_14777,N_13542,N_13639);
xor U14778 (N_14778,N_12038,N_12993);
nand U14779 (N_14779,N_13244,N_12234);
xnor U14780 (N_14780,N_12531,N_13472);
nor U14781 (N_14781,N_13141,N_13113);
nand U14782 (N_14782,N_12221,N_13538);
xor U14783 (N_14783,N_12193,N_12282);
nand U14784 (N_14784,N_12051,N_12838);
xnor U14785 (N_14785,N_13261,N_13585);
nor U14786 (N_14786,N_13093,N_12446);
nand U14787 (N_14787,N_13492,N_13830);
xor U14788 (N_14788,N_13679,N_12630);
nor U14789 (N_14789,N_13341,N_13702);
xnor U14790 (N_14790,N_13703,N_13897);
nor U14791 (N_14791,N_12088,N_12498);
and U14792 (N_14792,N_13283,N_13578);
nand U14793 (N_14793,N_12183,N_12750);
xor U14794 (N_14794,N_12484,N_12565);
nor U14795 (N_14795,N_13433,N_12297);
xnor U14796 (N_14796,N_13125,N_12864);
or U14797 (N_14797,N_13298,N_13294);
nor U14798 (N_14798,N_13121,N_13931);
nor U14799 (N_14799,N_12240,N_12545);
xnor U14800 (N_14800,N_12012,N_13535);
and U14801 (N_14801,N_13644,N_12478);
nor U14802 (N_14802,N_13293,N_13354);
nor U14803 (N_14803,N_12049,N_12955);
or U14804 (N_14804,N_13645,N_12603);
nand U14805 (N_14805,N_13928,N_13598);
nand U14806 (N_14806,N_13004,N_12797);
nor U14807 (N_14807,N_12210,N_12586);
and U14808 (N_14808,N_13944,N_12249);
or U14809 (N_14809,N_12697,N_12966);
nand U14810 (N_14810,N_13609,N_12199);
nor U14811 (N_14811,N_13094,N_13153);
nor U14812 (N_14812,N_13539,N_12016);
nor U14813 (N_14813,N_12308,N_12976);
or U14814 (N_14814,N_12480,N_13712);
xor U14815 (N_14815,N_12037,N_12330);
or U14816 (N_14816,N_13476,N_13739);
and U14817 (N_14817,N_12084,N_12688);
or U14818 (N_14818,N_13008,N_13752);
or U14819 (N_14819,N_13572,N_12757);
xnor U14820 (N_14820,N_12522,N_12105);
or U14821 (N_14821,N_13408,N_12325);
or U14822 (N_14822,N_12405,N_12518);
and U14823 (N_14823,N_12521,N_12581);
nor U14824 (N_14824,N_13552,N_12848);
or U14825 (N_14825,N_13323,N_13692);
and U14826 (N_14826,N_12763,N_13688);
nor U14827 (N_14827,N_12691,N_12243);
nand U14828 (N_14828,N_12194,N_12232);
nor U14829 (N_14829,N_12636,N_13971);
nand U14830 (N_14830,N_12839,N_12494);
and U14831 (N_14831,N_13152,N_12902);
and U14832 (N_14832,N_12579,N_13134);
nand U14833 (N_14833,N_12136,N_13468);
xnor U14834 (N_14834,N_13954,N_12001);
xor U14835 (N_14835,N_12333,N_12178);
nor U14836 (N_14836,N_12739,N_12986);
xor U14837 (N_14837,N_13994,N_12488);
or U14838 (N_14838,N_12288,N_13276);
nor U14839 (N_14839,N_13348,N_13860);
or U14840 (N_14840,N_12883,N_12671);
and U14841 (N_14841,N_13883,N_12570);
nand U14842 (N_14842,N_12935,N_12475);
and U14843 (N_14843,N_12466,N_12780);
nor U14844 (N_14844,N_12121,N_12889);
xor U14845 (N_14845,N_13938,N_13767);
nand U14846 (N_14846,N_12877,N_13711);
nor U14847 (N_14847,N_12830,N_12593);
nor U14848 (N_14848,N_13201,N_13753);
nor U14849 (N_14849,N_12707,N_12588);
nor U14850 (N_14850,N_13997,N_13715);
xor U14851 (N_14851,N_12548,N_12646);
nand U14852 (N_14852,N_12042,N_13878);
nand U14853 (N_14853,N_12218,N_13775);
and U14854 (N_14854,N_12857,N_13518);
nand U14855 (N_14855,N_13064,N_12969);
or U14856 (N_14856,N_12310,N_13654);
xnor U14857 (N_14857,N_12269,N_12887);
nor U14858 (N_14858,N_12436,N_12280);
nand U14859 (N_14859,N_12342,N_13721);
nor U14860 (N_14860,N_12005,N_13850);
nand U14861 (N_14861,N_13013,N_12140);
and U14862 (N_14862,N_12159,N_12057);
xor U14863 (N_14863,N_12997,N_13999);
nand U14864 (N_14864,N_12590,N_12914);
or U14865 (N_14865,N_13773,N_13811);
xnor U14866 (N_14866,N_13056,N_13792);
nand U14867 (N_14867,N_13704,N_12142);
and U14868 (N_14868,N_13312,N_12314);
and U14869 (N_14869,N_13895,N_13418);
xor U14870 (N_14870,N_13763,N_13618);
nand U14871 (N_14871,N_13078,N_13528);
and U14872 (N_14872,N_13870,N_12146);
nand U14873 (N_14873,N_13175,N_13082);
nand U14874 (N_14874,N_12219,N_12716);
and U14875 (N_14875,N_13785,N_12040);
and U14876 (N_14876,N_12659,N_13904);
or U14877 (N_14877,N_13292,N_12876);
nor U14878 (N_14878,N_13043,N_12212);
nor U14879 (N_14879,N_12414,N_12296);
xnor U14880 (N_14880,N_12073,N_13019);
or U14881 (N_14881,N_12574,N_13608);
and U14882 (N_14882,N_13477,N_13214);
xor U14883 (N_14883,N_12458,N_13435);
nor U14884 (N_14884,N_12293,N_13119);
nand U14885 (N_14885,N_12895,N_13723);
and U14886 (N_14886,N_13230,N_13974);
xor U14887 (N_14887,N_13428,N_13836);
or U14888 (N_14888,N_13902,N_13985);
nand U14889 (N_14889,N_13901,N_12383);
nand U14890 (N_14890,N_13571,N_13784);
xnor U14891 (N_14891,N_12619,N_12644);
nand U14892 (N_14892,N_13746,N_13265);
nand U14893 (N_14893,N_12597,N_12874);
or U14894 (N_14894,N_12131,N_13426);
nand U14895 (N_14895,N_13036,N_13586);
nor U14896 (N_14896,N_13663,N_12800);
and U14897 (N_14897,N_12787,N_12906);
or U14898 (N_14898,N_13110,N_13405);
nand U14899 (N_14899,N_13797,N_12585);
nor U14900 (N_14900,N_13482,N_12463);
and U14901 (N_14901,N_13956,N_12329);
nor U14902 (N_14902,N_13564,N_12766);
nor U14903 (N_14903,N_12956,N_12304);
xnor U14904 (N_14904,N_13829,N_13795);
xor U14905 (N_14905,N_13633,N_12503);
and U14906 (N_14906,N_12472,N_13506);
and U14907 (N_14907,N_12299,N_12950);
nor U14908 (N_14908,N_12726,N_12171);
xnor U14909 (N_14909,N_12174,N_12332);
xnor U14910 (N_14910,N_12176,N_13080);
xnor U14911 (N_14911,N_12534,N_13282);
xor U14912 (N_14912,N_13890,N_13710);
xnor U14913 (N_14913,N_13674,N_12445);
or U14914 (N_14914,N_12829,N_12384);
nor U14915 (N_14915,N_12300,N_13491);
or U14916 (N_14916,N_12932,N_13202);
nand U14917 (N_14917,N_13181,N_13454);
or U14918 (N_14918,N_12633,N_13237);
nand U14919 (N_14919,N_12305,N_12107);
and U14920 (N_14920,N_13220,N_13192);
and U14921 (N_14921,N_13927,N_12878);
nand U14922 (N_14922,N_13915,N_12318);
and U14923 (N_14923,N_13694,N_13756);
nand U14924 (N_14924,N_12362,N_12349);
or U14925 (N_14925,N_13194,N_12481);
or U14926 (N_14926,N_13962,N_12108);
or U14927 (N_14927,N_12898,N_13841);
nand U14928 (N_14928,N_13427,N_12753);
or U14929 (N_14929,N_13658,N_12344);
xor U14930 (N_14930,N_12509,N_12893);
or U14931 (N_14931,N_12922,N_12740);
nor U14932 (N_14932,N_13626,N_12313);
and U14933 (N_14933,N_13458,N_12009);
nand U14934 (N_14934,N_12925,N_13484);
and U14935 (N_14935,N_13868,N_13912);
nor U14936 (N_14936,N_12185,N_12918);
or U14937 (N_14937,N_12237,N_12851);
and U14938 (N_14938,N_12840,N_13166);
nand U14939 (N_14939,N_13450,N_12143);
nand U14940 (N_14940,N_12152,N_13251);
nor U14941 (N_14941,N_12687,N_13529);
and U14942 (N_14942,N_12395,N_12323);
xnor U14943 (N_14943,N_12664,N_13320);
nand U14944 (N_14944,N_13982,N_13589);
or U14945 (N_14945,N_12708,N_13896);
or U14946 (N_14946,N_13935,N_13519);
xnor U14947 (N_14947,N_12656,N_12663);
nand U14948 (N_14948,N_12366,N_13634);
and U14949 (N_14949,N_12117,N_13083);
nand U14950 (N_14950,N_12519,N_12209);
or U14951 (N_14951,N_12849,N_12681);
or U14952 (N_14952,N_12417,N_12431);
nor U14953 (N_14953,N_13827,N_13952);
nand U14954 (N_14954,N_12069,N_13888);
nand U14955 (N_14955,N_13280,N_12378);
and U14956 (N_14956,N_13964,N_12116);
nand U14957 (N_14957,N_12206,N_12345);
or U14958 (N_14958,N_13315,N_12050);
nand U14959 (N_14959,N_12820,N_12625);
or U14960 (N_14960,N_12315,N_12317);
nand U14961 (N_14961,N_13622,N_12064);
and U14962 (N_14962,N_13267,N_13554);
or U14963 (N_14963,N_13258,N_12462);
nor U14964 (N_14964,N_13215,N_12747);
nand U14965 (N_14965,N_13741,N_12803);
xnor U14966 (N_14966,N_13342,N_13336);
nor U14967 (N_14967,N_12985,N_13331);
nand U14968 (N_14968,N_13670,N_13494);
or U14969 (N_14969,N_13549,N_13180);
xnor U14970 (N_14970,N_12862,N_12652);
xnor U14971 (N_14971,N_12111,N_13766);
or U14972 (N_14972,N_12537,N_12551);
and U14973 (N_14973,N_12381,N_13274);
nand U14974 (N_14974,N_13382,N_12485);
or U14975 (N_14975,N_13821,N_13631);
nand U14976 (N_14976,N_13289,N_13164);
or U14977 (N_14977,N_12058,N_12949);
nand U14978 (N_14978,N_13005,N_13061);
nor U14979 (N_14979,N_12912,N_12482);
nand U14980 (N_14980,N_12281,N_12802);
nand U14981 (N_14981,N_13725,N_12693);
nor U14982 (N_14982,N_13972,N_12036);
nand U14983 (N_14983,N_13995,N_13807);
xor U14984 (N_14984,N_12622,N_12170);
nand U14985 (N_14985,N_12702,N_13319);
nor U14986 (N_14986,N_13022,N_12394);
or U14987 (N_14987,N_12929,N_13250);
or U14988 (N_14988,N_12676,N_13822);
and U14989 (N_14989,N_13247,N_13507);
and U14990 (N_14990,N_12267,N_13313);
xnor U14991 (N_14991,N_13976,N_12355);
nand U14992 (N_14992,N_13186,N_12913);
or U14993 (N_14993,N_12667,N_13024);
xor U14994 (N_14994,N_12904,N_12406);
nand U14995 (N_14995,N_13414,N_12160);
nor U14996 (N_14996,N_12047,N_13033);
nor U14997 (N_14997,N_12936,N_13389);
nor U14998 (N_14998,N_12248,N_13560);
nand U14999 (N_14999,N_12365,N_12286);
and U15000 (N_15000,N_12381,N_12736);
and U15001 (N_15001,N_13306,N_13927);
or U15002 (N_15002,N_12919,N_12268);
and U15003 (N_15003,N_13108,N_13192);
xnor U15004 (N_15004,N_13922,N_13072);
xor U15005 (N_15005,N_13849,N_13027);
xnor U15006 (N_15006,N_12482,N_13109);
and U15007 (N_15007,N_12796,N_12115);
nand U15008 (N_15008,N_13694,N_12460);
and U15009 (N_15009,N_12782,N_13371);
or U15010 (N_15010,N_13395,N_13261);
nor U15011 (N_15011,N_12417,N_12746);
nor U15012 (N_15012,N_12814,N_12967);
and U15013 (N_15013,N_12970,N_12784);
nand U15014 (N_15014,N_12499,N_13224);
or U15015 (N_15015,N_12033,N_13636);
or U15016 (N_15016,N_13076,N_13855);
xor U15017 (N_15017,N_12161,N_12255);
or U15018 (N_15018,N_13660,N_13282);
and U15019 (N_15019,N_12661,N_13190);
nor U15020 (N_15020,N_12700,N_13634);
nor U15021 (N_15021,N_13970,N_13621);
and U15022 (N_15022,N_13226,N_12209);
or U15023 (N_15023,N_12786,N_13610);
xor U15024 (N_15024,N_12266,N_13432);
nand U15025 (N_15025,N_13676,N_13609);
or U15026 (N_15026,N_12998,N_12901);
or U15027 (N_15027,N_12686,N_12712);
or U15028 (N_15028,N_13246,N_13933);
nand U15029 (N_15029,N_12506,N_12634);
nand U15030 (N_15030,N_13392,N_13999);
nor U15031 (N_15031,N_12501,N_12847);
nor U15032 (N_15032,N_12418,N_12833);
nand U15033 (N_15033,N_13260,N_13753);
xnor U15034 (N_15034,N_13997,N_13091);
or U15035 (N_15035,N_12721,N_12663);
or U15036 (N_15036,N_12806,N_13847);
and U15037 (N_15037,N_12367,N_12169);
and U15038 (N_15038,N_13949,N_12656);
or U15039 (N_15039,N_12696,N_13161);
nor U15040 (N_15040,N_12686,N_12583);
and U15041 (N_15041,N_12836,N_13338);
xor U15042 (N_15042,N_13592,N_13941);
nand U15043 (N_15043,N_12037,N_13413);
nor U15044 (N_15044,N_13154,N_12421);
xnor U15045 (N_15045,N_13959,N_12226);
and U15046 (N_15046,N_12421,N_13811);
nor U15047 (N_15047,N_13561,N_13769);
xor U15048 (N_15048,N_13985,N_13013);
xnor U15049 (N_15049,N_12765,N_12887);
and U15050 (N_15050,N_12849,N_13915);
nand U15051 (N_15051,N_13194,N_12937);
or U15052 (N_15052,N_13435,N_13414);
nor U15053 (N_15053,N_13628,N_13530);
nand U15054 (N_15054,N_13281,N_12239);
and U15055 (N_15055,N_12393,N_13975);
nor U15056 (N_15056,N_13028,N_13061);
nor U15057 (N_15057,N_12835,N_12814);
nand U15058 (N_15058,N_13263,N_12827);
nor U15059 (N_15059,N_12852,N_12487);
and U15060 (N_15060,N_12446,N_13209);
and U15061 (N_15061,N_13059,N_13165);
and U15062 (N_15062,N_12703,N_13889);
nor U15063 (N_15063,N_12297,N_13324);
xnor U15064 (N_15064,N_13160,N_12886);
nor U15065 (N_15065,N_13600,N_12278);
and U15066 (N_15066,N_13471,N_12373);
nand U15067 (N_15067,N_13104,N_13916);
and U15068 (N_15068,N_12659,N_13208);
nand U15069 (N_15069,N_12543,N_12044);
and U15070 (N_15070,N_12597,N_13598);
and U15071 (N_15071,N_12542,N_13673);
xnor U15072 (N_15072,N_13213,N_13294);
nor U15073 (N_15073,N_12718,N_13689);
xor U15074 (N_15074,N_12344,N_13082);
or U15075 (N_15075,N_13023,N_13742);
and U15076 (N_15076,N_12092,N_13661);
nand U15077 (N_15077,N_13351,N_13979);
nand U15078 (N_15078,N_12044,N_13343);
xor U15079 (N_15079,N_12115,N_13698);
nor U15080 (N_15080,N_13648,N_12116);
xor U15081 (N_15081,N_12901,N_12194);
nand U15082 (N_15082,N_12040,N_12340);
xnor U15083 (N_15083,N_12249,N_12537);
nand U15084 (N_15084,N_13951,N_13480);
nor U15085 (N_15085,N_12665,N_12063);
and U15086 (N_15086,N_13122,N_12735);
nand U15087 (N_15087,N_12130,N_12977);
nand U15088 (N_15088,N_12225,N_12682);
or U15089 (N_15089,N_13302,N_13009);
xor U15090 (N_15090,N_12530,N_12677);
or U15091 (N_15091,N_12881,N_13252);
nand U15092 (N_15092,N_13829,N_12989);
and U15093 (N_15093,N_12757,N_13422);
and U15094 (N_15094,N_12261,N_12195);
xnor U15095 (N_15095,N_12545,N_13924);
nand U15096 (N_15096,N_13523,N_12030);
or U15097 (N_15097,N_13168,N_12999);
or U15098 (N_15098,N_13238,N_12263);
nor U15099 (N_15099,N_12891,N_12480);
or U15100 (N_15100,N_12806,N_12926);
nor U15101 (N_15101,N_12032,N_13621);
nor U15102 (N_15102,N_13596,N_13299);
xor U15103 (N_15103,N_13923,N_12802);
nand U15104 (N_15104,N_13793,N_12640);
or U15105 (N_15105,N_13519,N_13022);
nand U15106 (N_15106,N_12516,N_13192);
and U15107 (N_15107,N_12255,N_13960);
or U15108 (N_15108,N_12742,N_13845);
nand U15109 (N_15109,N_13970,N_13706);
nand U15110 (N_15110,N_12681,N_13865);
or U15111 (N_15111,N_12454,N_13851);
nor U15112 (N_15112,N_12576,N_12580);
or U15113 (N_15113,N_13646,N_12629);
nand U15114 (N_15114,N_12366,N_13676);
xnor U15115 (N_15115,N_13448,N_12777);
nand U15116 (N_15116,N_13998,N_13496);
and U15117 (N_15117,N_12901,N_12506);
nand U15118 (N_15118,N_12745,N_12515);
xor U15119 (N_15119,N_13639,N_13934);
nor U15120 (N_15120,N_13750,N_13509);
nor U15121 (N_15121,N_12910,N_13262);
nor U15122 (N_15122,N_13712,N_12917);
or U15123 (N_15123,N_12114,N_12570);
nor U15124 (N_15124,N_12204,N_12442);
xnor U15125 (N_15125,N_13158,N_12532);
xor U15126 (N_15126,N_13313,N_13026);
nand U15127 (N_15127,N_13663,N_13058);
and U15128 (N_15128,N_13396,N_13477);
nand U15129 (N_15129,N_12699,N_13763);
xnor U15130 (N_15130,N_12533,N_12701);
or U15131 (N_15131,N_12807,N_12458);
nor U15132 (N_15132,N_13316,N_12411);
and U15133 (N_15133,N_12075,N_13339);
or U15134 (N_15134,N_13048,N_12355);
or U15135 (N_15135,N_13426,N_12097);
xnor U15136 (N_15136,N_13509,N_12167);
xnor U15137 (N_15137,N_12012,N_13879);
and U15138 (N_15138,N_13483,N_13306);
and U15139 (N_15139,N_13708,N_12039);
or U15140 (N_15140,N_13380,N_13456);
nand U15141 (N_15141,N_12330,N_12761);
and U15142 (N_15142,N_12470,N_12737);
nor U15143 (N_15143,N_13223,N_13218);
or U15144 (N_15144,N_12530,N_12727);
nand U15145 (N_15145,N_12128,N_12728);
xor U15146 (N_15146,N_13367,N_12604);
nand U15147 (N_15147,N_13053,N_12202);
xnor U15148 (N_15148,N_12400,N_13203);
nor U15149 (N_15149,N_13253,N_13726);
nor U15150 (N_15150,N_13905,N_12413);
nand U15151 (N_15151,N_13512,N_12057);
xnor U15152 (N_15152,N_13051,N_13004);
nor U15153 (N_15153,N_12805,N_13403);
xor U15154 (N_15154,N_12696,N_13049);
and U15155 (N_15155,N_13494,N_13056);
nand U15156 (N_15156,N_12221,N_12920);
nand U15157 (N_15157,N_12215,N_12633);
nor U15158 (N_15158,N_12234,N_13722);
or U15159 (N_15159,N_13376,N_12105);
nor U15160 (N_15160,N_12512,N_13303);
xnor U15161 (N_15161,N_13256,N_12751);
nand U15162 (N_15162,N_12754,N_13147);
xor U15163 (N_15163,N_13691,N_12140);
and U15164 (N_15164,N_13497,N_13285);
and U15165 (N_15165,N_13775,N_12303);
nand U15166 (N_15166,N_13713,N_13597);
or U15167 (N_15167,N_12340,N_12236);
and U15168 (N_15168,N_12596,N_13062);
xnor U15169 (N_15169,N_13679,N_12798);
xnor U15170 (N_15170,N_12950,N_13003);
and U15171 (N_15171,N_12237,N_12512);
xnor U15172 (N_15172,N_12838,N_13492);
nand U15173 (N_15173,N_13639,N_12441);
and U15174 (N_15174,N_12772,N_13985);
or U15175 (N_15175,N_13454,N_12794);
or U15176 (N_15176,N_12198,N_12679);
nand U15177 (N_15177,N_12427,N_12858);
or U15178 (N_15178,N_12496,N_13567);
and U15179 (N_15179,N_12055,N_12809);
and U15180 (N_15180,N_13797,N_12539);
nor U15181 (N_15181,N_13625,N_12133);
nand U15182 (N_15182,N_12840,N_13913);
and U15183 (N_15183,N_13067,N_13333);
nand U15184 (N_15184,N_12466,N_13874);
and U15185 (N_15185,N_13364,N_12724);
nor U15186 (N_15186,N_12599,N_12654);
or U15187 (N_15187,N_12255,N_13190);
or U15188 (N_15188,N_13954,N_12116);
xor U15189 (N_15189,N_13155,N_13603);
xnor U15190 (N_15190,N_12705,N_12115);
nand U15191 (N_15191,N_12526,N_13634);
and U15192 (N_15192,N_13439,N_13411);
and U15193 (N_15193,N_12232,N_13654);
nor U15194 (N_15194,N_12361,N_12181);
and U15195 (N_15195,N_13631,N_13935);
or U15196 (N_15196,N_13207,N_12118);
or U15197 (N_15197,N_12144,N_13688);
nor U15198 (N_15198,N_12333,N_12915);
xnor U15199 (N_15199,N_13702,N_13264);
or U15200 (N_15200,N_13048,N_13814);
nand U15201 (N_15201,N_12418,N_12769);
nor U15202 (N_15202,N_12594,N_12259);
xor U15203 (N_15203,N_12879,N_12693);
nor U15204 (N_15204,N_12172,N_12636);
and U15205 (N_15205,N_13355,N_13354);
nor U15206 (N_15206,N_13222,N_12380);
and U15207 (N_15207,N_13600,N_13853);
or U15208 (N_15208,N_13777,N_12370);
or U15209 (N_15209,N_13281,N_12223);
xor U15210 (N_15210,N_12426,N_13030);
nor U15211 (N_15211,N_12828,N_12002);
nor U15212 (N_15212,N_12463,N_12490);
nand U15213 (N_15213,N_13743,N_12966);
nand U15214 (N_15214,N_12993,N_12559);
xnor U15215 (N_15215,N_13662,N_13251);
and U15216 (N_15216,N_13360,N_13493);
and U15217 (N_15217,N_13693,N_13576);
nand U15218 (N_15218,N_13083,N_13110);
or U15219 (N_15219,N_13926,N_12586);
or U15220 (N_15220,N_12283,N_12670);
nor U15221 (N_15221,N_12563,N_12496);
and U15222 (N_15222,N_12604,N_13366);
and U15223 (N_15223,N_13230,N_13884);
or U15224 (N_15224,N_12857,N_12723);
or U15225 (N_15225,N_12422,N_13403);
xor U15226 (N_15226,N_12219,N_13136);
nand U15227 (N_15227,N_13531,N_13929);
xnor U15228 (N_15228,N_12261,N_12184);
xnor U15229 (N_15229,N_13841,N_13745);
or U15230 (N_15230,N_12581,N_13476);
xnor U15231 (N_15231,N_13802,N_12049);
nor U15232 (N_15232,N_12832,N_13794);
xnor U15233 (N_15233,N_12283,N_13810);
nor U15234 (N_15234,N_12001,N_13732);
nor U15235 (N_15235,N_13541,N_12379);
or U15236 (N_15236,N_12532,N_12413);
xnor U15237 (N_15237,N_13016,N_13771);
xor U15238 (N_15238,N_12686,N_13656);
xnor U15239 (N_15239,N_13441,N_12871);
nand U15240 (N_15240,N_12286,N_12535);
xor U15241 (N_15241,N_12815,N_12898);
and U15242 (N_15242,N_13410,N_12808);
nand U15243 (N_15243,N_12791,N_13791);
xor U15244 (N_15244,N_13769,N_13583);
nand U15245 (N_15245,N_12096,N_12514);
and U15246 (N_15246,N_13997,N_12075);
and U15247 (N_15247,N_13470,N_12108);
and U15248 (N_15248,N_13956,N_13729);
and U15249 (N_15249,N_12920,N_13101);
nor U15250 (N_15250,N_12375,N_12051);
and U15251 (N_15251,N_12261,N_12871);
nor U15252 (N_15252,N_13936,N_12353);
or U15253 (N_15253,N_13258,N_13719);
nor U15254 (N_15254,N_13314,N_12302);
and U15255 (N_15255,N_12943,N_13361);
nor U15256 (N_15256,N_12873,N_12039);
xor U15257 (N_15257,N_13803,N_13235);
nand U15258 (N_15258,N_13679,N_13317);
nor U15259 (N_15259,N_13649,N_12201);
and U15260 (N_15260,N_12286,N_12768);
nor U15261 (N_15261,N_13731,N_12124);
and U15262 (N_15262,N_12012,N_12895);
or U15263 (N_15263,N_12558,N_12340);
nand U15264 (N_15264,N_13416,N_12724);
or U15265 (N_15265,N_12361,N_12434);
nor U15266 (N_15266,N_12652,N_13344);
xor U15267 (N_15267,N_13993,N_13730);
nand U15268 (N_15268,N_13088,N_13281);
and U15269 (N_15269,N_13715,N_12195);
or U15270 (N_15270,N_12203,N_12861);
xor U15271 (N_15271,N_12774,N_12950);
nand U15272 (N_15272,N_13314,N_12478);
nand U15273 (N_15273,N_13219,N_12545);
nand U15274 (N_15274,N_12990,N_13348);
nand U15275 (N_15275,N_12478,N_12201);
nand U15276 (N_15276,N_13380,N_13881);
and U15277 (N_15277,N_13844,N_12908);
xnor U15278 (N_15278,N_12372,N_13768);
nor U15279 (N_15279,N_12054,N_13468);
nor U15280 (N_15280,N_13646,N_12565);
nand U15281 (N_15281,N_12119,N_12883);
xor U15282 (N_15282,N_13982,N_13469);
and U15283 (N_15283,N_13317,N_12519);
xnor U15284 (N_15284,N_12520,N_13355);
and U15285 (N_15285,N_12702,N_12555);
nand U15286 (N_15286,N_13258,N_12007);
or U15287 (N_15287,N_12211,N_12175);
or U15288 (N_15288,N_12296,N_13694);
and U15289 (N_15289,N_13970,N_12310);
nor U15290 (N_15290,N_12011,N_13081);
xnor U15291 (N_15291,N_13009,N_13347);
xor U15292 (N_15292,N_13789,N_13784);
or U15293 (N_15293,N_12365,N_13654);
or U15294 (N_15294,N_12872,N_13197);
nand U15295 (N_15295,N_13445,N_12302);
nand U15296 (N_15296,N_13225,N_13249);
nor U15297 (N_15297,N_12905,N_13827);
or U15298 (N_15298,N_13596,N_12994);
nand U15299 (N_15299,N_13896,N_13657);
nand U15300 (N_15300,N_13512,N_12905);
xnor U15301 (N_15301,N_12190,N_12295);
and U15302 (N_15302,N_13703,N_12476);
and U15303 (N_15303,N_13964,N_12763);
and U15304 (N_15304,N_12660,N_12142);
or U15305 (N_15305,N_12954,N_13983);
or U15306 (N_15306,N_12225,N_12893);
and U15307 (N_15307,N_13155,N_13628);
or U15308 (N_15308,N_13574,N_13358);
nand U15309 (N_15309,N_13161,N_13876);
nor U15310 (N_15310,N_12160,N_12695);
xor U15311 (N_15311,N_13999,N_12116);
xor U15312 (N_15312,N_13049,N_12883);
and U15313 (N_15313,N_13145,N_12560);
and U15314 (N_15314,N_12439,N_12960);
or U15315 (N_15315,N_12654,N_12303);
and U15316 (N_15316,N_12115,N_13942);
nand U15317 (N_15317,N_13615,N_12086);
nand U15318 (N_15318,N_12273,N_13942);
nand U15319 (N_15319,N_13070,N_12788);
xor U15320 (N_15320,N_13921,N_12747);
and U15321 (N_15321,N_12381,N_12030);
nor U15322 (N_15322,N_13393,N_13620);
nor U15323 (N_15323,N_12134,N_12996);
nor U15324 (N_15324,N_12107,N_13321);
xnor U15325 (N_15325,N_13073,N_13665);
and U15326 (N_15326,N_12275,N_13953);
xor U15327 (N_15327,N_13365,N_13234);
xor U15328 (N_15328,N_12942,N_12614);
xor U15329 (N_15329,N_13673,N_12906);
nand U15330 (N_15330,N_13998,N_12374);
and U15331 (N_15331,N_12195,N_13344);
xnor U15332 (N_15332,N_12827,N_12123);
and U15333 (N_15333,N_12720,N_13002);
nor U15334 (N_15334,N_13266,N_13918);
nand U15335 (N_15335,N_12818,N_12553);
nand U15336 (N_15336,N_13369,N_13729);
xor U15337 (N_15337,N_12384,N_12111);
xor U15338 (N_15338,N_12618,N_13720);
or U15339 (N_15339,N_12055,N_13751);
or U15340 (N_15340,N_13603,N_12392);
nor U15341 (N_15341,N_12772,N_13353);
or U15342 (N_15342,N_12707,N_13170);
xnor U15343 (N_15343,N_12500,N_13069);
nor U15344 (N_15344,N_13539,N_13160);
nand U15345 (N_15345,N_12822,N_12190);
nand U15346 (N_15346,N_13709,N_12701);
xor U15347 (N_15347,N_12119,N_12675);
xor U15348 (N_15348,N_13898,N_12352);
or U15349 (N_15349,N_13351,N_12862);
xnor U15350 (N_15350,N_13814,N_12416);
or U15351 (N_15351,N_12040,N_13169);
and U15352 (N_15352,N_13907,N_12194);
nor U15353 (N_15353,N_12666,N_12960);
or U15354 (N_15354,N_13530,N_12158);
nand U15355 (N_15355,N_12628,N_12997);
nand U15356 (N_15356,N_13304,N_13757);
nand U15357 (N_15357,N_13090,N_13036);
xnor U15358 (N_15358,N_13744,N_12755);
xor U15359 (N_15359,N_12765,N_13345);
nand U15360 (N_15360,N_12143,N_13023);
xor U15361 (N_15361,N_13831,N_13643);
xnor U15362 (N_15362,N_12902,N_13548);
or U15363 (N_15363,N_12949,N_13629);
nand U15364 (N_15364,N_13458,N_13975);
or U15365 (N_15365,N_12438,N_12843);
or U15366 (N_15366,N_12085,N_13418);
or U15367 (N_15367,N_12839,N_12057);
and U15368 (N_15368,N_12216,N_13396);
xor U15369 (N_15369,N_13657,N_12536);
nor U15370 (N_15370,N_12226,N_12838);
nand U15371 (N_15371,N_13967,N_13378);
or U15372 (N_15372,N_13423,N_13209);
xor U15373 (N_15373,N_13274,N_13514);
nor U15374 (N_15374,N_13574,N_12197);
nor U15375 (N_15375,N_12768,N_13780);
or U15376 (N_15376,N_12244,N_12507);
and U15377 (N_15377,N_13540,N_12814);
xnor U15378 (N_15378,N_12099,N_13037);
and U15379 (N_15379,N_13364,N_13148);
nor U15380 (N_15380,N_12923,N_13909);
xor U15381 (N_15381,N_12218,N_12957);
or U15382 (N_15382,N_12636,N_12078);
nand U15383 (N_15383,N_12167,N_12112);
or U15384 (N_15384,N_12164,N_12462);
nor U15385 (N_15385,N_13451,N_12033);
xnor U15386 (N_15386,N_13158,N_13579);
nor U15387 (N_15387,N_12699,N_12465);
and U15388 (N_15388,N_12490,N_12262);
xor U15389 (N_15389,N_12793,N_13166);
nand U15390 (N_15390,N_12036,N_12942);
nor U15391 (N_15391,N_12999,N_13128);
nor U15392 (N_15392,N_12144,N_12912);
xor U15393 (N_15393,N_13397,N_13325);
or U15394 (N_15394,N_13214,N_12907);
and U15395 (N_15395,N_12025,N_12420);
and U15396 (N_15396,N_13386,N_12106);
and U15397 (N_15397,N_12440,N_12958);
nand U15398 (N_15398,N_12801,N_12460);
nor U15399 (N_15399,N_12382,N_12558);
nor U15400 (N_15400,N_13516,N_13459);
and U15401 (N_15401,N_13545,N_13950);
or U15402 (N_15402,N_12425,N_13869);
and U15403 (N_15403,N_12269,N_12653);
and U15404 (N_15404,N_12690,N_13941);
xnor U15405 (N_15405,N_13354,N_12920);
nor U15406 (N_15406,N_12831,N_13740);
and U15407 (N_15407,N_13947,N_12509);
nor U15408 (N_15408,N_13139,N_13226);
or U15409 (N_15409,N_13384,N_13860);
xnor U15410 (N_15410,N_12740,N_13785);
nor U15411 (N_15411,N_13706,N_13967);
xor U15412 (N_15412,N_13072,N_12878);
nor U15413 (N_15413,N_13699,N_13172);
nand U15414 (N_15414,N_12799,N_13405);
nor U15415 (N_15415,N_12686,N_12258);
xnor U15416 (N_15416,N_13017,N_13415);
nor U15417 (N_15417,N_12532,N_12335);
or U15418 (N_15418,N_13465,N_13231);
xnor U15419 (N_15419,N_13494,N_12437);
and U15420 (N_15420,N_12152,N_12296);
nand U15421 (N_15421,N_12212,N_13530);
xor U15422 (N_15422,N_13914,N_13261);
nand U15423 (N_15423,N_12768,N_12244);
nand U15424 (N_15424,N_13988,N_13320);
nand U15425 (N_15425,N_12665,N_13318);
and U15426 (N_15426,N_12106,N_12013);
and U15427 (N_15427,N_12024,N_13157);
nor U15428 (N_15428,N_13037,N_13574);
and U15429 (N_15429,N_12175,N_12024);
nor U15430 (N_15430,N_13353,N_12936);
nand U15431 (N_15431,N_13006,N_12458);
or U15432 (N_15432,N_13861,N_13005);
or U15433 (N_15433,N_12291,N_12144);
nand U15434 (N_15434,N_12603,N_12922);
xnor U15435 (N_15435,N_13651,N_13917);
nor U15436 (N_15436,N_12082,N_13918);
or U15437 (N_15437,N_12575,N_12768);
or U15438 (N_15438,N_12792,N_12620);
and U15439 (N_15439,N_12709,N_12913);
or U15440 (N_15440,N_13608,N_13911);
xnor U15441 (N_15441,N_12980,N_12595);
and U15442 (N_15442,N_12062,N_13768);
xor U15443 (N_15443,N_12583,N_12534);
or U15444 (N_15444,N_13563,N_13212);
nand U15445 (N_15445,N_12905,N_13916);
nand U15446 (N_15446,N_12209,N_12367);
xnor U15447 (N_15447,N_12808,N_12343);
or U15448 (N_15448,N_12092,N_13673);
nor U15449 (N_15449,N_12451,N_12025);
and U15450 (N_15450,N_13130,N_13929);
nand U15451 (N_15451,N_12132,N_13065);
nor U15452 (N_15452,N_12943,N_13151);
xor U15453 (N_15453,N_13360,N_12671);
nor U15454 (N_15454,N_13649,N_12494);
nor U15455 (N_15455,N_12775,N_12644);
xnor U15456 (N_15456,N_13687,N_12867);
nor U15457 (N_15457,N_12106,N_13391);
xnor U15458 (N_15458,N_12589,N_12478);
nand U15459 (N_15459,N_12343,N_13250);
nor U15460 (N_15460,N_12254,N_12970);
xor U15461 (N_15461,N_12958,N_12952);
nor U15462 (N_15462,N_12689,N_13169);
or U15463 (N_15463,N_13670,N_12110);
and U15464 (N_15464,N_12574,N_12083);
and U15465 (N_15465,N_12267,N_13338);
nor U15466 (N_15466,N_12296,N_12047);
nand U15467 (N_15467,N_12713,N_12528);
and U15468 (N_15468,N_12223,N_13757);
nand U15469 (N_15469,N_13752,N_12677);
nor U15470 (N_15470,N_12579,N_13729);
or U15471 (N_15471,N_12890,N_12085);
nand U15472 (N_15472,N_12702,N_12787);
and U15473 (N_15473,N_13109,N_13315);
nor U15474 (N_15474,N_13570,N_13710);
or U15475 (N_15475,N_13069,N_12135);
nand U15476 (N_15476,N_13058,N_12104);
and U15477 (N_15477,N_12762,N_13664);
and U15478 (N_15478,N_13444,N_13386);
or U15479 (N_15479,N_13636,N_13911);
xnor U15480 (N_15480,N_12392,N_12337);
xor U15481 (N_15481,N_13343,N_12978);
xnor U15482 (N_15482,N_13705,N_12724);
nor U15483 (N_15483,N_12775,N_13348);
and U15484 (N_15484,N_13694,N_12775);
and U15485 (N_15485,N_13317,N_12660);
nand U15486 (N_15486,N_13995,N_12560);
xnor U15487 (N_15487,N_13320,N_12316);
or U15488 (N_15488,N_12940,N_13641);
and U15489 (N_15489,N_12956,N_13439);
and U15490 (N_15490,N_13864,N_13158);
and U15491 (N_15491,N_13483,N_12568);
or U15492 (N_15492,N_13130,N_12351);
and U15493 (N_15493,N_12717,N_13890);
nand U15494 (N_15494,N_13272,N_13674);
and U15495 (N_15495,N_12739,N_12437);
xor U15496 (N_15496,N_13469,N_12806);
and U15497 (N_15497,N_12163,N_12272);
nand U15498 (N_15498,N_13900,N_12783);
nand U15499 (N_15499,N_13821,N_12265);
nor U15500 (N_15500,N_13693,N_12453);
nand U15501 (N_15501,N_13134,N_12239);
nor U15502 (N_15502,N_12884,N_12223);
nand U15503 (N_15503,N_12010,N_12646);
and U15504 (N_15504,N_12308,N_12032);
and U15505 (N_15505,N_12895,N_13506);
or U15506 (N_15506,N_13354,N_13783);
nand U15507 (N_15507,N_12054,N_13372);
nor U15508 (N_15508,N_12456,N_13295);
nand U15509 (N_15509,N_13828,N_13222);
xor U15510 (N_15510,N_13272,N_13779);
xnor U15511 (N_15511,N_13002,N_13276);
nand U15512 (N_15512,N_12877,N_13627);
and U15513 (N_15513,N_12455,N_13977);
nand U15514 (N_15514,N_13636,N_13567);
and U15515 (N_15515,N_12925,N_12949);
xor U15516 (N_15516,N_12688,N_13631);
xor U15517 (N_15517,N_12352,N_13740);
xnor U15518 (N_15518,N_12381,N_12271);
nand U15519 (N_15519,N_13541,N_12245);
nor U15520 (N_15520,N_13911,N_13975);
nand U15521 (N_15521,N_13679,N_12817);
xor U15522 (N_15522,N_13073,N_13191);
and U15523 (N_15523,N_13342,N_13952);
nor U15524 (N_15524,N_13537,N_13610);
nand U15525 (N_15525,N_13135,N_12126);
and U15526 (N_15526,N_12433,N_13930);
and U15527 (N_15527,N_13405,N_12100);
or U15528 (N_15528,N_13619,N_12282);
nor U15529 (N_15529,N_12666,N_13907);
nand U15530 (N_15530,N_13125,N_12495);
or U15531 (N_15531,N_12989,N_13639);
nand U15532 (N_15532,N_12310,N_13437);
xor U15533 (N_15533,N_12852,N_12819);
nand U15534 (N_15534,N_12303,N_13071);
and U15535 (N_15535,N_12223,N_12315);
and U15536 (N_15536,N_13663,N_12911);
nand U15537 (N_15537,N_12267,N_13089);
or U15538 (N_15538,N_12913,N_13368);
and U15539 (N_15539,N_13938,N_13490);
nand U15540 (N_15540,N_13679,N_13594);
nor U15541 (N_15541,N_13512,N_12542);
nor U15542 (N_15542,N_12277,N_13885);
or U15543 (N_15543,N_13583,N_12588);
nor U15544 (N_15544,N_13488,N_12053);
or U15545 (N_15545,N_12175,N_12931);
nand U15546 (N_15546,N_12506,N_13847);
nor U15547 (N_15547,N_12850,N_12885);
xor U15548 (N_15548,N_12167,N_12286);
nor U15549 (N_15549,N_13054,N_12491);
and U15550 (N_15550,N_13113,N_12706);
xnor U15551 (N_15551,N_13531,N_12980);
xor U15552 (N_15552,N_13273,N_12110);
xnor U15553 (N_15553,N_13645,N_12476);
or U15554 (N_15554,N_13756,N_13052);
and U15555 (N_15555,N_13386,N_12233);
or U15556 (N_15556,N_13183,N_12057);
nand U15557 (N_15557,N_12903,N_12812);
nand U15558 (N_15558,N_13967,N_13539);
xor U15559 (N_15559,N_12874,N_12533);
xnor U15560 (N_15560,N_12555,N_12152);
nor U15561 (N_15561,N_12567,N_12590);
nor U15562 (N_15562,N_12142,N_12014);
and U15563 (N_15563,N_13015,N_12979);
nand U15564 (N_15564,N_12974,N_13379);
nor U15565 (N_15565,N_13380,N_13985);
or U15566 (N_15566,N_13952,N_13078);
nor U15567 (N_15567,N_13926,N_13728);
nor U15568 (N_15568,N_13405,N_12650);
nor U15569 (N_15569,N_13610,N_13776);
nand U15570 (N_15570,N_12870,N_12427);
nand U15571 (N_15571,N_13620,N_13855);
xor U15572 (N_15572,N_12591,N_12184);
nand U15573 (N_15573,N_12338,N_13658);
xnor U15574 (N_15574,N_13750,N_13407);
nor U15575 (N_15575,N_13435,N_13239);
or U15576 (N_15576,N_12937,N_12957);
and U15577 (N_15577,N_12645,N_13325);
and U15578 (N_15578,N_12746,N_12986);
or U15579 (N_15579,N_12655,N_13378);
nand U15580 (N_15580,N_13507,N_13343);
and U15581 (N_15581,N_12442,N_13468);
or U15582 (N_15582,N_12656,N_13361);
xnor U15583 (N_15583,N_12867,N_13353);
and U15584 (N_15584,N_13668,N_13819);
nand U15585 (N_15585,N_12337,N_13443);
xor U15586 (N_15586,N_13067,N_12581);
and U15587 (N_15587,N_12448,N_12666);
xor U15588 (N_15588,N_13074,N_12147);
and U15589 (N_15589,N_12810,N_12877);
and U15590 (N_15590,N_12902,N_13737);
xor U15591 (N_15591,N_12760,N_12289);
xnor U15592 (N_15592,N_13930,N_12671);
nand U15593 (N_15593,N_12366,N_13719);
nand U15594 (N_15594,N_13517,N_12052);
nor U15595 (N_15595,N_12469,N_12001);
or U15596 (N_15596,N_12496,N_12481);
nor U15597 (N_15597,N_12363,N_12386);
xor U15598 (N_15598,N_12818,N_12838);
nor U15599 (N_15599,N_12316,N_13227);
nor U15600 (N_15600,N_12214,N_13304);
nand U15601 (N_15601,N_13631,N_12758);
nand U15602 (N_15602,N_12305,N_12505);
nor U15603 (N_15603,N_13761,N_12925);
nor U15604 (N_15604,N_13009,N_13532);
nor U15605 (N_15605,N_13831,N_13468);
xnor U15606 (N_15606,N_12481,N_13899);
or U15607 (N_15607,N_12931,N_12283);
nor U15608 (N_15608,N_13847,N_12668);
and U15609 (N_15609,N_12504,N_12369);
nor U15610 (N_15610,N_13635,N_13787);
or U15611 (N_15611,N_13608,N_12741);
or U15612 (N_15612,N_12782,N_13414);
and U15613 (N_15613,N_12564,N_12752);
nor U15614 (N_15614,N_12582,N_12225);
xor U15615 (N_15615,N_13212,N_12277);
and U15616 (N_15616,N_12945,N_13788);
nand U15617 (N_15617,N_13758,N_13113);
xor U15618 (N_15618,N_13313,N_12731);
nand U15619 (N_15619,N_12454,N_12327);
and U15620 (N_15620,N_12751,N_13871);
nor U15621 (N_15621,N_12778,N_12861);
xor U15622 (N_15622,N_13029,N_12496);
xor U15623 (N_15623,N_12550,N_13531);
nand U15624 (N_15624,N_12059,N_13719);
or U15625 (N_15625,N_13693,N_12305);
and U15626 (N_15626,N_13625,N_12431);
and U15627 (N_15627,N_12452,N_12058);
nand U15628 (N_15628,N_13876,N_13482);
xnor U15629 (N_15629,N_13205,N_13069);
nor U15630 (N_15630,N_12749,N_12657);
and U15631 (N_15631,N_13865,N_13179);
or U15632 (N_15632,N_12208,N_13266);
or U15633 (N_15633,N_12834,N_13945);
nor U15634 (N_15634,N_13378,N_12593);
nor U15635 (N_15635,N_13602,N_13730);
nand U15636 (N_15636,N_12372,N_12971);
or U15637 (N_15637,N_12737,N_13436);
nor U15638 (N_15638,N_12561,N_12429);
or U15639 (N_15639,N_13004,N_12049);
nand U15640 (N_15640,N_13652,N_13207);
and U15641 (N_15641,N_13817,N_12809);
or U15642 (N_15642,N_13602,N_13308);
nor U15643 (N_15643,N_13559,N_13265);
and U15644 (N_15644,N_13022,N_12894);
or U15645 (N_15645,N_13248,N_12329);
and U15646 (N_15646,N_12100,N_12337);
nor U15647 (N_15647,N_13826,N_12139);
and U15648 (N_15648,N_13821,N_12781);
xor U15649 (N_15649,N_12059,N_13193);
nand U15650 (N_15650,N_13427,N_13702);
nor U15651 (N_15651,N_13886,N_12907);
nand U15652 (N_15652,N_12043,N_12228);
nor U15653 (N_15653,N_12528,N_13633);
or U15654 (N_15654,N_12324,N_12607);
or U15655 (N_15655,N_12244,N_13513);
nor U15656 (N_15656,N_12024,N_12050);
and U15657 (N_15657,N_13441,N_13160);
or U15658 (N_15658,N_13968,N_12097);
xor U15659 (N_15659,N_12706,N_12456);
nor U15660 (N_15660,N_12716,N_13388);
nand U15661 (N_15661,N_13422,N_13676);
nor U15662 (N_15662,N_13614,N_12464);
or U15663 (N_15663,N_12850,N_13070);
nand U15664 (N_15664,N_13553,N_13888);
or U15665 (N_15665,N_13596,N_12521);
nor U15666 (N_15666,N_13647,N_13249);
and U15667 (N_15667,N_13304,N_13964);
and U15668 (N_15668,N_12043,N_12204);
nor U15669 (N_15669,N_13873,N_13212);
nor U15670 (N_15670,N_13118,N_13041);
xnor U15671 (N_15671,N_12577,N_13547);
nand U15672 (N_15672,N_12332,N_12564);
nor U15673 (N_15673,N_12014,N_12068);
and U15674 (N_15674,N_12645,N_12581);
xor U15675 (N_15675,N_12020,N_13481);
and U15676 (N_15676,N_12258,N_12735);
or U15677 (N_15677,N_12186,N_13605);
nor U15678 (N_15678,N_13880,N_13684);
and U15679 (N_15679,N_13288,N_12097);
or U15680 (N_15680,N_12548,N_12961);
nand U15681 (N_15681,N_13336,N_12058);
and U15682 (N_15682,N_12885,N_12293);
or U15683 (N_15683,N_12885,N_13986);
and U15684 (N_15684,N_13460,N_13918);
and U15685 (N_15685,N_13276,N_12549);
or U15686 (N_15686,N_13830,N_13079);
nand U15687 (N_15687,N_12761,N_13254);
or U15688 (N_15688,N_13712,N_12671);
and U15689 (N_15689,N_12284,N_13082);
nand U15690 (N_15690,N_12439,N_12814);
and U15691 (N_15691,N_13491,N_13528);
xnor U15692 (N_15692,N_12983,N_12511);
nand U15693 (N_15693,N_13074,N_13467);
nor U15694 (N_15694,N_13210,N_13503);
nor U15695 (N_15695,N_13512,N_13474);
and U15696 (N_15696,N_12633,N_13067);
nor U15697 (N_15697,N_12013,N_13328);
or U15698 (N_15698,N_12963,N_13545);
xor U15699 (N_15699,N_12692,N_12967);
nor U15700 (N_15700,N_13693,N_13148);
nor U15701 (N_15701,N_13955,N_12970);
nand U15702 (N_15702,N_12756,N_13425);
or U15703 (N_15703,N_12827,N_13041);
xor U15704 (N_15704,N_12069,N_12622);
nand U15705 (N_15705,N_12178,N_12138);
nor U15706 (N_15706,N_13460,N_13183);
or U15707 (N_15707,N_13116,N_12690);
xor U15708 (N_15708,N_13777,N_13985);
or U15709 (N_15709,N_13395,N_13412);
nand U15710 (N_15710,N_12282,N_13453);
or U15711 (N_15711,N_12300,N_12856);
nand U15712 (N_15712,N_12649,N_12753);
xnor U15713 (N_15713,N_13978,N_13660);
nor U15714 (N_15714,N_12821,N_13547);
nand U15715 (N_15715,N_13036,N_13495);
nor U15716 (N_15716,N_13494,N_13813);
nand U15717 (N_15717,N_12184,N_12378);
and U15718 (N_15718,N_13235,N_12944);
or U15719 (N_15719,N_13952,N_13236);
nor U15720 (N_15720,N_12064,N_13757);
nand U15721 (N_15721,N_12228,N_12790);
and U15722 (N_15722,N_12047,N_13210);
and U15723 (N_15723,N_12390,N_13359);
nor U15724 (N_15724,N_13367,N_12064);
nor U15725 (N_15725,N_13250,N_12265);
xor U15726 (N_15726,N_13982,N_13132);
nand U15727 (N_15727,N_12707,N_13013);
nand U15728 (N_15728,N_13605,N_12018);
xor U15729 (N_15729,N_13011,N_13064);
nand U15730 (N_15730,N_13738,N_13397);
nand U15731 (N_15731,N_13829,N_13023);
nand U15732 (N_15732,N_13926,N_12387);
nor U15733 (N_15733,N_12430,N_13360);
nor U15734 (N_15734,N_13206,N_13321);
nand U15735 (N_15735,N_12636,N_12383);
xor U15736 (N_15736,N_13383,N_13195);
and U15737 (N_15737,N_12438,N_12230);
nor U15738 (N_15738,N_13057,N_13958);
or U15739 (N_15739,N_12853,N_12657);
nand U15740 (N_15740,N_12048,N_13439);
and U15741 (N_15741,N_12379,N_13043);
or U15742 (N_15742,N_13507,N_12214);
xor U15743 (N_15743,N_13177,N_13530);
and U15744 (N_15744,N_12622,N_13777);
and U15745 (N_15745,N_12997,N_12657);
or U15746 (N_15746,N_12650,N_13016);
nand U15747 (N_15747,N_13838,N_13984);
nor U15748 (N_15748,N_12936,N_13120);
and U15749 (N_15749,N_13074,N_12023);
xor U15750 (N_15750,N_13322,N_13290);
xnor U15751 (N_15751,N_13807,N_13668);
nand U15752 (N_15752,N_12997,N_12590);
or U15753 (N_15753,N_13786,N_12383);
nand U15754 (N_15754,N_13934,N_13880);
and U15755 (N_15755,N_12688,N_13804);
xor U15756 (N_15756,N_12875,N_12069);
or U15757 (N_15757,N_13010,N_13957);
and U15758 (N_15758,N_12799,N_13407);
nand U15759 (N_15759,N_13017,N_12476);
nand U15760 (N_15760,N_12393,N_12263);
or U15761 (N_15761,N_12173,N_12627);
or U15762 (N_15762,N_13801,N_12170);
nor U15763 (N_15763,N_13503,N_13677);
nor U15764 (N_15764,N_12551,N_12594);
nor U15765 (N_15765,N_12122,N_13339);
and U15766 (N_15766,N_12730,N_12948);
nor U15767 (N_15767,N_12122,N_12659);
nor U15768 (N_15768,N_13486,N_12645);
xor U15769 (N_15769,N_12647,N_12467);
and U15770 (N_15770,N_13885,N_12568);
nand U15771 (N_15771,N_13745,N_13725);
or U15772 (N_15772,N_12035,N_13044);
nand U15773 (N_15773,N_13259,N_13780);
nand U15774 (N_15774,N_13407,N_12490);
or U15775 (N_15775,N_12920,N_12339);
or U15776 (N_15776,N_13967,N_12330);
nand U15777 (N_15777,N_12609,N_13599);
nand U15778 (N_15778,N_12985,N_12430);
and U15779 (N_15779,N_13723,N_12679);
nor U15780 (N_15780,N_12207,N_12855);
or U15781 (N_15781,N_12958,N_13765);
nor U15782 (N_15782,N_12760,N_13393);
and U15783 (N_15783,N_13179,N_12190);
nand U15784 (N_15784,N_12829,N_12225);
xnor U15785 (N_15785,N_12063,N_13188);
nor U15786 (N_15786,N_13413,N_12944);
and U15787 (N_15787,N_12286,N_13829);
and U15788 (N_15788,N_12873,N_12546);
nor U15789 (N_15789,N_12282,N_13200);
nand U15790 (N_15790,N_13700,N_12994);
nand U15791 (N_15791,N_13310,N_13175);
xnor U15792 (N_15792,N_12032,N_12286);
nand U15793 (N_15793,N_12722,N_12822);
xor U15794 (N_15794,N_13685,N_13238);
nand U15795 (N_15795,N_12043,N_13274);
nand U15796 (N_15796,N_12458,N_12683);
or U15797 (N_15797,N_12484,N_12938);
or U15798 (N_15798,N_12886,N_13673);
and U15799 (N_15799,N_12502,N_13555);
and U15800 (N_15800,N_13423,N_12606);
nor U15801 (N_15801,N_12657,N_12656);
nand U15802 (N_15802,N_13675,N_13211);
nand U15803 (N_15803,N_12405,N_13350);
nor U15804 (N_15804,N_13540,N_12861);
nor U15805 (N_15805,N_13275,N_13642);
nand U15806 (N_15806,N_13955,N_13456);
nor U15807 (N_15807,N_13151,N_13513);
nand U15808 (N_15808,N_13392,N_13192);
and U15809 (N_15809,N_12416,N_12510);
xor U15810 (N_15810,N_12327,N_12906);
or U15811 (N_15811,N_13664,N_13240);
nand U15812 (N_15812,N_12009,N_13854);
and U15813 (N_15813,N_12243,N_12675);
nor U15814 (N_15814,N_12264,N_13732);
nor U15815 (N_15815,N_13771,N_13105);
nand U15816 (N_15816,N_13696,N_13078);
nor U15817 (N_15817,N_13923,N_13849);
or U15818 (N_15818,N_13533,N_13532);
xnor U15819 (N_15819,N_13183,N_12090);
nand U15820 (N_15820,N_13552,N_12297);
xor U15821 (N_15821,N_12631,N_12797);
or U15822 (N_15822,N_12619,N_12509);
xnor U15823 (N_15823,N_13868,N_13231);
xor U15824 (N_15824,N_12023,N_12574);
or U15825 (N_15825,N_12241,N_12525);
nor U15826 (N_15826,N_13252,N_13865);
or U15827 (N_15827,N_13965,N_13803);
and U15828 (N_15828,N_12201,N_12703);
nand U15829 (N_15829,N_12121,N_13390);
xor U15830 (N_15830,N_13767,N_13111);
or U15831 (N_15831,N_12977,N_13940);
nor U15832 (N_15832,N_13036,N_12714);
nand U15833 (N_15833,N_12586,N_13971);
nand U15834 (N_15834,N_12549,N_13612);
or U15835 (N_15835,N_13099,N_13540);
and U15836 (N_15836,N_13425,N_13980);
nor U15837 (N_15837,N_13405,N_12277);
and U15838 (N_15838,N_12953,N_12314);
or U15839 (N_15839,N_12195,N_12387);
nor U15840 (N_15840,N_13751,N_12218);
and U15841 (N_15841,N_12693,N_13687);
and U15842 (N_15842,N_13337,N_12019);
nand U15843 (N_15843,N_12581,N_12558);
and U15844 (N_15844,N_13754,N_13258);
xor U15845 (N_15845,N_13762,N_12517);
and U15846 (N_15846,N_12864,N_13577);
nand U15847 (N_15847,N_12790,N_13844);
or U15848 (N_15848,N_12756,N_12776);
nor U15849 (N_15849,N_12334,N_12625);
xor U15850 (N_15850,N_12932,N_12309);
nand U15851 (N_15851,N_12310,N_12275);
and U15852 (N_15852,N_12927,N_12964);
xnor U15853 (N_15853,N_12857,N_12517);
nor U15854 (N_15854,N_12420,N_12314);
nor U15855 (N_15855,N_13192,N_12703);
xnor U15856 (N_15856,N_12304,N_12535);
or U15857 (N_15857,N_13229,N_12263);
nand U15858 (N_15858,N_12209,N_12425);
xnor U15859 (N_15859,N_12953,N_13817);
nand U15860 (N_15860,N_13372,N_13203);
and U15861 (N_15861,N_13708,N_12249);
or U15862 (N_15862,N_12969,N_12083);
nor U15863 (N_15863,N_12453,N_12860);
or U15864 (N_15864,N_13654,N_13412);
xor U15865 (N_15865,N_12678,N_13375);
nor U15866 (N_15866,N_13194,N_13755);
xnor U15867 (N_15867,N_12886,N_13402);
and U15868 (N_15868,N_12261,N_12136);
xor U15869 (N_15869,N_12702,N_12562);
nor U15870 (N_15870,N_12217,N_12371);
nor U15871 (N_15871,N_12508,N_12450);
nor U15872 (N_15872,N_12904,N_13727);
and U15873 (N_15873,N_12515,N_12070);
or U15874 (N_15874,N_13396,N_12581);
xnor U15875 (N_15875,N_12950,N_13775);
nor U15876 (N_15876,N_12224,N_12064);
or U15877 (N_15877,N_13475,N_13440);
nand U15878 (N_15878,N_12813,N_12394);
or U15879 (N_15879,N_13233,N_13275);
and U15880 (N_15880,N_12396,N_12598);
nor U15881 (N_15881,N_13281,N_13532);
nor U15882 (N_15882,N_13292,N_13361);
and U15883 (N_15883,N_13727,N_13101);
nand U15884 (N_15884,N_12053,N_12344);
and U15885 (N_15885,N_12854,N_12918);
or U15886 (N_15886,N_13402,N_13945);
xnor U15887 (N_15887,N_13544,N_13710);
nand U15888 (N_15888,N_12610,N_13416);
nand U15889 (N_15889,N_12352,N_13136);
nand U15890 (N_15890,N_12682,N_13574);
nor U15891 (N_15891,N_13771,N_13712);
nand U15892 (N_15892,N_13619,N_12636);
xnor U15893 (N_15893,N_12122,N_13864);
nand U15894 (N_15894,N_13269,N_12008);
or U15895 (N_15895,N_13864,N_13308);
nand U15896 (N_15896,N_12918,N_12484);
nor U15897 (N_15897,N_12684,N_12021);
or U15898 (N_15898,N_12564,N_12864);
nor U15899 (N_15899,N_13134,N_13384);
nor U15900 (N_15900,N_13928,N_13848);
or U15901 (N_15901,N_12562,N_12430);
nand U15902 (N_15902,N_12081,N_13489);
xnor U15903 (N_15903,N_12615,N_13008);
nor U15904 (N_15904,N_13736,N_12328);
nor U15905 (N_15905,N_12263,N_13157);
and U15906 (N_15906,N_13118,N_12264);
or U15907 (N_15907,N_12935,N_12501);
nor U15908 (N_15908,N_13877,N_13651);
and U15909 (N_15909,N_12353,N_13014);
nor U15910 (N_15910,N_13386,N_13495);
and U15911 (N_15911,N_12535,N_12383);
nor U15912 (N_15912,N_13462,N_13883);
nor U15913 (N_15913,N_13827,N_12324);
nor U15914 (N_15914,N_12425,N_12303);
nor U15915 (N_15915,N_13443,N_13022);
and U15916 (N_15916,N_13049,N_12457);
or U15917 (N_15917,N_12192,N_12131);
nand U15918 (N_15918,N_13546,N_13725);
and U15919 (N_15919,N_12935,N_12898);
xor U15920 (N_15920,N_13989,N_12585);
and U15921 (N_15921,N_12558,N_12186);
and U15922 (N_15922,N_12136,N_13510);
or U15923 (N_15923,N_13014,N_13465);
nor U15924 (N_15924,N_13005,N_13312);
nand U15925 (N_15925,N_13404,N_12206);
nor U15926 (N_15926,N_13599,N_12102);
and U15927 (N_15927,N_13762,N_12082);
nand U15928 (N_15928,N_13129,N_13840);
xor U15929 (N_15929,N_12197,N_13805);
or U15930 (N_15930,N_13369,N_12701);
and U15931 (N_15931,N_13315,N_12309);
xor U15932 (N_15932,N_13831,N_12783);
nor U15933 (N_15933,N_13667,N_12368);
xor U15934 (N_15934,N_12500,N_12189);
or U15935 (N_15935,N_12235,N_12417);
nand U15936 (N_15936,N_12013,N_12941);
or U15937 (N_15937,N_13634,N_12240);
or U15938 (N_15938,N_12280,N_12814);
or U15939 (N_15939,N_13723,N_12105);
nand U15940 (N_15940,N_12348,N_13681);
or U15941 (N_15941,N_13220,N_12715);
nor U15942 (N_15942,N_12819,N_12662);
xor U15943 (N_15943,N_12137,N_13464);
and U15944 (N_15944,N_13790,N_13199);
xor U15945 (N_15945,N_12664,N_12035);
nor U15946 (N_15946,N_12500,N_12572);
or U15947 (N_15947,N_12153,N_13398);
nand U15948 (N_15948,N_12079,N_13245);
nor U15949 (N_15949,N_12495,N_12279);
nand U15950 (N_15950,N_13347,N_12819);
and U15951 (N_15951,N_12006,N_12341);
nor U15952 (N_15952,N_13812,N_13319);
xnor U15953 (N_15953,N_13849,N_12680);
nand U15954 (N_15954,N_12288,N_13654);
and U15955 (N_15955,N_12080,N_12675);
nand U15956 (N_15956,N_13712,N_13493);
nor U15957 (N_15957,N_12220,N_12877);
xor U15958 (N_15958,N_12823,N_13466);
nand U15959 (N_15959,N_13409,N_13813);
and U15960 (N_15960,N_12604,N_13257);
nor U15961 (N_15961,N_13586,N_13915);
or U15962 (N_15962,N_13915,N_12459);
nand U15963 (N_15963,N_12181,N_13879);
and U15964 (N_15964,N_13287,N_12525);
nor U15965 (N_15965,N_13276,N_13812);
or U15966 (N_15966,N_13686,N_13335);
xor U15967 (N_15967,N_12656,N_12728);
or U15968 (N_15968,N_13208,N_12403);
and U15969 (N_15969,N_12120,N_12787);
xnor U15970 (N_15970,N_13733,N_13378);
nor U15971 (N_15971,N_12228,N_12265);
or U15972 (N_15972,N_12853,N_12747);
xor U15973 (N_15973,N_12770,N_13760);
nand U15974 (N_15974,N_13846,N_13256);
nor U15975 (N_15975,N_12487,N_12878);
nand U15976 (N_15976,N_12014,N_13274);
xnor U15977 (N_15977,N_13687,N_13523);
nor U15978 (N_15978,N_13290,N_12769);
or U15979 (N_15979,N_13837,N_12327);
nor U15980 (N_15980,N_12774,N_12588);
or U15981 (N_15981,N_12971,N_12954);
or U15982 (N_15982,N_13405,N_13133);
nand U15983 (N_15983,N_13947,N_13272);
or U15984 (N_15984,N_13210,N_13505);
nand U15985 (N_15985,N_12589,N_12715);
and U15986 (N_15986,N_13442,N_13054);
nor U15987 (N_15987,N_12847,N_12575);
nor U15988 (N_15988,N_12118,N_12972);
nand U15989 (N_15989,N_13856,N_12803);
or U15990 (N_15990,N_13660,N_13006);
or U15991 (N_15991,N_13449,N_12080);
nor U15992 (N_15992,N_13741,N_12837);
and U15993 (N_15993,N_13575,N_12650);
xnor U15994 (N_15994,N_12994,N_13335);
nor U15995 (N_15995,N_12458,N_12009);
xor U15996 (N_15996,N_12383,N_13420);
xnor U15997 (N_15997,N_12819,N_13287);
nor U15998 (N_15998,N_13050,N_12116);
nand U15999 (N_15999,N_13384,N_12912);
or U16000 (N_16000,N_15618,N_14404);
nor U16001 (N_16001,N_15816,N_14772);
xnor U16002 (N_16002,N_14593,N_15567);
and U16003 (N_16003,N_14998,N_15543);
xor U16004 (N_16004,N_14101,N_14665);
nand U16005 (N_16005,N_15845,N_15891);
and U16006 (N_16006,N_14856,N_14103);
or U16007 (N_16007,N_14565,N_15938);
nand U16008 (N_16008,N_15827,N_14415);
nor U16009 (N_16009,N_14975,N_14810);
or U16010 (N_16010,N_14739,N_14821);
nand U16011 (N_16011,N_14852,N_15369);
nor U16012 (N_16012,N_15590,N_15706);
xnor U16013 (N_16013,N_15751,N_15526);
nand U16014 (N_16014,N_14115,N_15904);
nand U16015 (N_16015,N_15614,N_15785);
and U16016 (N_16016,N_15700,N_14639);
and U16017 (N_16017,N_14248,N_14498);
nor U16018 (N_16018,N_15948,N_15488);
and U16019 (N_16019,N_15296,N_15546);
nor U16020 (N_16020,N_15688,N_15886);
or U16021 (N_16021,N_15340,N_15789);
or U16022 (N_16022,N_15698,N_14876);
nand U16023 (N_16023,N_14267,N_14475);
xnor U16024 (N_16024,N_14082,N_14813);
nor U16025 (N_16025,N_14923,N_15986);
nand U16026 (N_16026,N_15790,N_14805);
and U16027 (N_16027,N_15941,N_14218);
nor U16028 (N_16028,N_14036,N_15737);
and U16029 (N_16029,N_14118,N_15588);
or U16030 (N_16030,N_15311,N_15875);
nand U16031 (N_16031,N_14793,N_15542);
and U16032 (N_16032,N_15987,N_14698);
or U16033 (N_16033,N_14357,N_14191);
or U16034 (N_16034,N_14410,N_15778);
and U16035 (N_16035,N_15067,N_14868);
or U16036 (N_16036,N_15158,N_14290);
xnor U16037 (N_16037,N_14866,N_14053);
or U16038 (N_16038,N_14936,N_14685);
nor U16039 (N_16039,N_15981,N_14968);
nand U16040 (N_16040,N_14459,N_15378);
and U16041 (N_16041,N_15834,N_14104);
nand U16042 (N_16042,N_14586,N_14594);
and U16043 (N_16043,N_15846,N_15723);
or U16044 (N_16044,N_15772,N_14519);
nand U16045 (N_16045,N_15294,N_14327);
nand U16046 (N_16046,N_15093,N_15727);
nor U16047 (N_16047,N_14385,N_15308);
nand U16048 (N_16048,N_14427,N_14478);
and U16049 (N_16049,N_14347,N_14567);
xor U16050 (N_16050,N_15556,N_14188);
nor U16051 (N_16051,N_15998,N_14880);
xor U16052 (N_16052,N_14642,N_14893);
or U16053 (N_16053,N_14530,N_15525);
and U16054 (N_16054,N_15092,N_15513);
or U16055 (N_16055,N_14303,N_14534);
nand U16056 (N_16056,N_14691,N_15157);
xnor U16057 (N_16057,N_14243,N_14570);
and U16058 (N_16058,N_15508,N_14881);
xor U16059 (N_16059,N_15693,N_14069);
or U16060 (N_16060,N_14786,N_14771);
or U16061 (N_16061,N_14169,N_15787);
nor U16062 (N_16062,N_15857,N_15582);
nand U16063 (N_16063,N_15667,N_15350);
xnor U16064 (N_16064,N_14662,N_14065);
or U16065 (N_16065,N_14807,N_14766);
xnor U16066 (N_16066,N_14367,N_14007);
and U16067 (N_16067,N_14251,N_15393);
nor U16068 (N_16068,N_14528,N_14734);
nand U16069 (N_16069,N_15195,N_15578);
xor U16070 (N_16070,N_14356,N_14401);
and U16071 (N_16071,N_14765,N_15042);
and U16072 (N_16072,N_15596,N_14254);
nand U16073 (N_16073,N_14215,N_15500);
xor U16074 (N_16074,N_15627,N_15359);
nand U16075 (N_16075,N_15775,N_15247);
nor U16076 (N_16076,N_15939,N_14536);
nand U16077 (N_16077,N_14063,N_14937);
nand U16078 (N_16078,N_15583,N_14195);
nor U16079 (N_16079,N_15759,N_14669);
xor U16080 (N_16080,N_15485,N_15664);
nand U16081 (N_16081,N_15849,N_15484);
and U16082 (N_16082,N_14078,N_14213);
or U16083 (N_16083,N_15019,N_14483);
nor U16084 (N_16084,N_15116,N_15553);
nand U16085 (N_16085,N_15464,N_14768);
or U16086 (N_16086,N_15275,N_15933);
nand U16087 (N_16087,N_15123,N_15000);
nor U16088 (N_16088,N_15741,N_15690);
and U16089 (N_16089,N_14462,N_14736);
and U16090 (N_16090,N_15906,N_14283);
xor U16091 (N_16091,N_14155,N_15397);
nor U16092 (N_16092,N_15476,N_15905);
and U16093 (N_16093,N_15370,N_14764);
or U16094 (N_16094,N_14173,N_14981);
nand U16095 (N_16095,N_14600,N_14130);
xor U16096 (N_16096,N_14783,N_15190);
xor U16097 (N_16097,N_14450,N_14754);
nor U16098 (N_16098,N_14321,N_14743);
xnor U16099 (N_16099,N_14549,N_14268);
nand U16100 (N_16100,N_15189,N_15745);
nor U16101 (N_16101,N_14770,N_14407);
or U16102 (N_16102,N_14910,N_15035);
nor U16103 (N_16103,N_15044,N_15844);
and U16104 (N_16104,N_15843,N_15911);
and U16105 (N_16105,N_15623,N_14080);
or U16106 (N_16106,N_15616,N_14884);
and U16107 (N_16107,N_15026,N_15233);
or U16108 (N_16108,N_15396,N_14819);
xnor U16109 (N_16109,N_14794,N_15868);
xor U16110 (N_16110,N_14216,N_14751);
or U16111 (N_16111,N_15991,N_15815);
and U16112 (N_16112,N_14129,N_15628);
xor U16113 (N_16113,N_15854,N_14343);
nand U16114 (N_16114,N_15413,N_15654);
and U16115 (N_16115,N_14220,N_15156);
xnor U16116 (N_16116,N_14317,N_15612);
nor U16117 (N_16117,N_14151,N_14399);
nor U16118 (N_16118,N_15557,N_15277);
nand U16119 (N_16119,N_15864,N_14087);
nand U16120 (N_16120,N_15070,N_14266);
or U16121 (N_16121,N_15381,N_14644);
or U16122 (N_16122,N_14707,N_14869);
nor U16123 (N_16123,N_14732,N_14603);
nand U16124 (N_16124,N_15328,N_15341);
and U16125 (N_16125,N_15115,N_15231);
nand U16126 (N_16126,N_14730,N_15848);
or U16127 (N_16127,N_15744,N_14311);
xor U16128 (N_16128,N_14544,N_15235);
and U16129 (N_16129,N_14481,N_14948);
nor U16130 (N_16130,N_14812,N_14919);
nand U16131 (N_16131,N_14066,N_14988);
nor U16132 (N_16132,N_14712,N_15021);
nand U16133 (N_16133,N_14822,N_15399);
and U16134 (N_16134,N_15504,N_15184);
and U16135 (N_16135,N_14389,N_15361);
nor U16136 (N_16136,N_15477,N_15808);
nand U16137 (N_16137,N_15368,N_15358);
nor U16138 (N_16138,N_15642,N_15168);
or U16139 (N_16139,N_15585,N_15382);
nand U16140 (N_16140,N_14461,N_14980);
nor U16141 (N_16141,N_14942,N_14500);
nor U16142 (N_16142,N_15315,N_14718);
nand U16143 (N_16143,N_15527,N_15813);
nor U16144 (N_16144,N_15427,N_14554);
and U16145 (N_16145,N_14895,N_14705);
xor U16146 (N_16146,N_15036,N_15022);
or U16147 (N_16147,N_15554,N_15602);
nor U16148 (N_16148,N_14967,N_14622);
nand U16149 (N_16149,N_14903,N_15204);
and U16150 (N_16150,N_15853,N_15812);
nor U16151 (N_16151,N_15877,N_15647);
nand U16152 (N_16152,N_14714,N_15946);
xnor U16153 (N_16153,N_15482,N_15901);
xnor U16154 (N_16154,N_15650,N_15803);
nand U16155 (N_16155,N_15112,N_15975);
or U16156 (N_16156,N_14201,N_15316);
nand U16157 (N_16157,N_15964,N_14380);
xor U16158 (N_16158,N_15979,N_14175);
and U16159 (N_16159,N_15739,N_15037);
nor U16160 (N_16160,N_15207,N_14741);
and U16161 (N_16161,N_15391,N_14829);
and U16162 (N_16162,N_15266,N_14274);
and U16163 (N_16163,N_15137,N_14862);
nor U16164 (N_16164,N_15564,N_14889);
nor U16165 (N_16165,N_14432,N_15593);
nand U16166 (N_16166,N_15101,N_15186);
nor U16167 (N_16167,N_15798,N_14933);
xor U16168 (N_16168,N_15704,N_15724);
and U16169 (N_16169,N_14178,N_14228);
xor U16170 (N_16170,N_15347,N_15534);
and U16171 (N_16171,N_14750,N_15434);
and U16172 (N_16172,N_14154,N_15185);
or U16173 (N_16173,N_14577,N_15565);
nor U16174 (N_16174,N_14495,N_15281);
nor U16175 (N_16175,N_14328,N_14072);
or U16176 (N_16176,N_15407,N_14106);
xor U16177 (N_16177,N_15383,N_15555);
nand U16178 (N_16178,N_15489,N_15071);
and U16179 (N_16179,N_14974,N_14767);
nor U16180 (N_16180,N_14197,N_14905);
nand U16181 (N_16181,N_15668,N_15379);
nor U16182 (N_16182,N_15620,N_14177);
nor U16183 (N_16183,N_15760,N_14985);
nor U16184 (N_16184,N_14443,N_15757);
nand U16185 (N_16185,N_14445,N_14575);
and U16186 (N_16186,N_15119,N_15129);
xor U16187 (N_16187,N_14476,N_14637);
and U16188 (N_16188,N_14150,N_15060);
nor U16189 (N_16189,N_15828,N_14945);
nand U16190 (N_16190,N_15100,N_14107);
or U16191 (N_16191,N_15097,N_14253);
nor U16192 (N_16192,N_15136,N_14326);
xor U16193 (N_16193,N_15122,N_15841);
or U16194 (N_16194,N_15175,N_14314);
nand U16195 (N_16195,N_15675,N_15142);
xnor U16196 (N_16196,N_14044,N_15882);
and U16197 (N_16197,N_15535,N_14011);
nor U16198 (N_16198,N_15963,N_14291);
and U16199 (N_16199,N_15989,N_15452);
and U16200 (N_16200,N_14791,N_15301);
or U16201 (N_16201,N_15162,N_14935);
and U16202 (N_16202,N_14913,N_14553);
or U16203 (N_16203,N_15514,N_15734);
or U16204 (N_16204,N_15694,N_14999);
nor U16205 (N_16205,N_15453,N_15012);
xor U16206 (N_16206,N_15171,N_15286);
or U16207 (N_16207,N_14433,N_15638);
nor U16208 (N_16208,N_14606,N_14839);
or U16209 (N_16209,N_15299,N_14378);
or U16210 (N_16210,N_14841,N_14735);
and U16211 (N_16211,N_14120,N_15742);
xor U16212 (N_16212,N_14275,N_15220);
or U16213 (N_16213,N_14752,N_15643);
or U16214 (N_16214,N_14789,N_15249);
nor U16215 (N_16215,N_14668,N_15120);
and U16216 (N_16216,N_15914,N_15290);
or U16217 (N_16217,N_15440,N_14288);
and U16218 (N_16218,N_14001,N_14131);
or U16219 (N_16219,N_15323,N_14260);
and U16220 (N_16220,N_14515,N_14806);
or U16221 (N_16221,N_14949,N_15715);
and U16222 (N_16222,N_14697,N_15591);
nor U16223 (N_16223,N_14894,N_15404);
and U16224 (N_16224,N_14664,N_14505);
nand U16225 (N_16225,N_14959,N_15151);
and U16226 (N_16226,N_14695,N_15897);
or U16227 (N_16227,N_14912,N_15716);
or U16228 (N_16228,N_15372,N_14004);
xor U16229 (N_16229,N_14047,N_14815);
or U16230 (N_16230,N_15641,N_15894);
xor U16231 (N_16231,N_15114,N_14859);
xor U16232 (N_16232,N_15264,N_14437);
nand U16233 (N_16233,N_14015,N_15697);
and U16234 (N_16234,N_14026,N_14121);
and U16235 (N_16235,N_14074,N_15385);
or U16236 (N_16236,N_15572,N_15260);
xnor U16237 (N_16237,N_15819,N_14111);
xnor U16238 (N_16238,N_14846,N_14997);
and U16239 (N_16239,N_15038,N_15059);
or U16240 (N_16240,N_14145,N_14143);
or U16241 (N_16241,N_15725,N_15245);
and U16242 (N_16242,N_15773,N_15273);
nand U16243 (N_16243,N_14406,N_15515);
xnor U16244 (N_16244,N_15839,N_15820);
nor U16245 (N_16245,N_14374,N_14711);
nand U16246 (N_16246,N_15199,N_14763);
and U16247 (N_16247,N_14064,N_15880);
nor U16248 (N_16248,N_15892,N_14079);
and U16249 (N_16249,N_14473,N_15153);
nand U16250 (N_16250,N_14636,N_14235);
nor U16251 (N_16251,N_14008,N_14715);
nand U16252 (N_16252,N_15083,N_15018);
nand U16253 (N_16253,N_14986,N_15943);
nand U16254 (N_16254,N_15467,N_15632);
nor U16255 (N_16255,N_14453,N_15659);
xnor U16256 (N_16256,N_14482,N_14262);
xnor U16257 (N_16257,N_15302,N_14511);
nor U16258 (N_16258,N_14616,N_15028);
or U16259 (N_16259,N_15133,N_14214);
nand U16260 (N_16260,N_14246,N_14513);
nand U16261 (N_16261,N_15931,N_14908);
nor U16262 (N_16262,N_15226,N_15146);
nand U16263 (N_16263,N_15858,N_15009);
or U16264 (N_16264,N_14413,N_15072);
nand U16265 (N_16265,N_15511,N_14496);
nor U16266 (N_16266,N_14068,N_14661);
or U16267 (N_16267,N_14397,N_14579);
or U16268 (N_16268,N_14133,N_15971);
nand U16269 (N_16269,N_15896,N_14409);
xor U16270 (N_16270,N_14452,N_14788);
and U16271 (N_16271,N_15814,N_14623);
or U16272 (N_16272,N_14993,N_14434);
nand U16273 (N_16273,N_14329,N_15164);
xor U16274 (N_16274,N_14323,N_15374);
or U16275 (N_16275,N_14860,N_15254);
nand U16276 (N_16276,N_15096,N_14541);
nand U16277 (N_16277,N_15961,N_15173);
nor U16278 (N_16278,N_14689,N_14117);
nand U16279 (N_16279,N_15597,N_15278);
and U16280 (N_16280,N_14164,N_15479);
or U16281 (N_16281,N_15522,N_15421);
xnor U16282 (N_16282,N_14010,N_15492);
nand U16283 (N_16283,N_14849,N_15962);
xor U16284 (N_16284,N_15767,N_14179);
and U16285 (N_16285,N_14836,N_14223);
xnor U16286 (N_16286,N_14635,N_15509);
nand U16287 (N_16287,N_15799,N_15624);
nor U16288 (N_16288,N_15353,N_15463);
and U16289 (N_16289,N_14414,N_15625);
xnor U16290 (N_16290,N_15159,N_15371);
or U16291 (N_16291,N_14672,N_14088);
nand U16292 (N_16292,N_15068,N_14900);
xnor U16293 (N_16293,N_15983,N_15405);
nor U16294 (N_16294,N_15373,N_15674);
xor U16295 (N_16295,N_14576,N_15054);
or U16296 (N_16296,N_14094,N_15292);
nand U16297 (N_16297,N_15430,N_15279);
xor U16298 (N_16298,N_15346,N_14073);
nor U16299 (N_16299,N_15900,N_15993);
or U16300 (N_16300,N_15563,N_15388);
and U16301 (N_16301,N_15005,N_15141);
and U16302 (N_16302,N_15013,N_15148);
and U16303 (N_16303,N_14281,N_14890);
xnor U16304 (N_16304,N_15539,N_14070);
or U16305 (N_16305,N_14146,N_15507);
nand U16306 (N_16306,N_15389,N_15763);
or U16307 (N_16307,N_14924,N_14817);
or U16308 (N_16308,N_14390,N_15058);
and U16309 (N_16309,N_14393,N_15280);
nand U16310 (N_16310,N_14950,N_14264);
nand U16311 (N_16311,N_15468,N_15995);
nor U16312 (N_16312,N_14899,N_14555);
and U16313 (N_16313,N_14052,N_14921);
nand U16314 (N_16314,N_15577,N_15147);
and U16315 (N_16315,N_14799,N_15793);
nor U16316 (N_16316,N_14420,N_14774);
nor U16317 (N_16317,N_15717,N_14388);
nor U16318 (N_16318,N_14350,N_14381);
xor U16319 (N_16319,N_14911,N_15826);
and U16320 (N_16320,N_15656,N_14244);
nand U16321 (N_16321,N_15663,N_14471);
and U16322 (N_16322,N_15465,N_14883);
nor U16323 (N_16323,N_15672,N_15551);
and U16324 (N_16324,N_15817,N_15532);
or U16325 (N_16325,N_14369,N_14673);
and U16326 (N_16326,N_14927,N_14640);
nand U16327 (N_16327,N_15291,N_15272);
and U16328 (N_16328,N_14840,N_14670);
or U16329 (N_16329,N_14828,N_14929);
nand U16330 (N_16330,N_15603,N_15924);
nand U16331 (N_16331,N_14435,N_15771);
and U16332 (N_16332,N_14067,N_14261);
xor U16333 (N_16333,N_14907,N_15615);
nand U16334 (N_16334,N_15258,N_14322);
nor U16335 (N_16335,N_14428,N_14493);
nor U16336 (N_16336,N_14863,N_15387);
nor U16337 (N_16337,N_15889,N_14609);
nand U16338 (N_16338,N_14250,N_15325);
and U16339 (N_16339,N_14124,N_15073);
or U16340 (N_16340,N_15053,N_15196);
xor U16341 (N_16341,N_14760,N_14688);
or U16342 (N_16342,N_15910,N_14231);
nand U16343 (N_16343,N_14904,N_14990);
nand U16344 (N_16344,N_15182,N_15985);
nand U16345 (N_16345,N_15738,N_15197);
nor U16346 (N_16346,N_15437,N_15940);
xnor U16347 (N_16347,N_14958,N_15458);
or U16348 (N_16348,N_14787,N_15203);
nand U16349 (N_16349,N_15351,N_15867);
or U16350 (N_16350,N_15214,N_15818);
or U16351 (N_16351,N_15211,N_15568);
xor U16352 (N_16352,N_15836,N_14558);
nand U16353 (N_16353,N_14604,N_14305);
xnor U16354 (N_16354,N_15970,N_14527);
nor U16355 (N_16355,N_15908,N_14503);
xor U16356 (N_16356,N_14324,N_14539);
nor U16357 (N_16357,N_15777,N_14611);
and U16358 (N_16358,N_15521,N_15598);
and U16359 (N_16359,N_14271,N_15749);
and U16360 (N_16360,N_15224,N_15860);
and U16361 (N_16361,N_14075,N_14973);
nand U16362 (N_16362,N_14666,N_14867);
and U16363 (N_16363,N_15866,N_14257);
nand U16364 (N_16364,N_14790,N_14396);
xor U16365 (N_16365,N_14897,N_14142);
and U16366 (N_16366,N_15640,N_14370);
or U16367 (N_16367,N_15746,N_14510);
xor U16368 (N_16368,N_15095,N_15890);
or U16369 (N_16369,N_14494,N_14674);
xnor U16370 (N_16370,N_15721,N_14280);
and U16371 (N_16371,N_15613,N_15718);
or U16372 (N_16372,N_15611,N_15055);
and U16373 (N_16373,N_15080,N_15735);
xnor U16374 (N_16374,N_14285,N_14134);
or U16375 (N_16375,N_15242,N_15478);
xor U16376 (N_16376,N_15363,N_14917);
xor U16377 (N_16377,N_15418,N_15960);
nand U16378 (N_16378,N_15893,N_14293);
xor U16379 (N_16379,N_15150,N_15781);
nand U16380 (N_16380,N_15110,N_15335);
and U16381 (N_16381,N_15105,N_14237);
and U16382 (N_16382,N_14458,N_15268);
xor U16383 (N_16383,N_15395,N_14012);
nor U16384 (N_16384,N_14831,N_14827);
and U16385 (N_16385,N_15743,N_14196);
xnor U16386 (N_16386,N_14330,N_14272);
nor U16387 (N_16387,N_14631,N_15671);
xnor U16388 (N_16388,N_15973,N_15592);
or U16389 (N_16389,N_14287,N_15855);
nand U16390 (N_16390,N_15409,N_15579);
xnor U16391 (N_16391,N_14242,N_14972);
xnor U16392 (N_16392,N_15202,N_14227);
or U16393 (N_16393,N_15135,N_15566);
xnor U16394 (N_16394,N_15431,N_15187);
or U16395 (N_16395,N_14308,N_14418);
xor U16396 (N_16396,N_14731,N_15248);
and U16397 (N_16397,N_15732,N_15861);
and U16398 (N_16398,N_15753,N_14844);
nand U16399 (N_16399,N_14375,N_14093);
or U16400 (N_16400,N_14159,N_14447);
xor U16401 (N_16401,N_15265,N_14795);
and U16402 (N_16402,N_15673,N_15040);
nand U16403 (N_16403,N_15322,N_15318);
or U16404 (N_16404,N_15108,N_15253);
nor U16405 (N_16405,N_15851,N_15102);
or U16406 (N_16406,N_14934,N_14132);
or U16407 (N_16407,N_15712,N_15008);
nand U16408 (N_16408,N_15953,N_14531);
and U16409 (N_16409,N_15017,N_14858);
and U16410 (N_16410,N_14028,N_15473);
or U16411 (N_16411,N_14671,N_15284);
and U16412 (N_16412,N_14190,N_15711);
nor U16413 (N_16413,N_14488,N_14708);
or U16414 (N_16414,N_15559,N_14588);
xnor U16415 (N_16415,N_15916,N_14372);
nor U16416 (N_16416,N_14803,N_14978);
or U16417 (N_16417,N_15143,N_14684);
or U16418 (N_16418,N_15402,N_14725);
or U16419 (N_16419,N_14710,N_14187);
xnor U16420 (N_16420,N_14773,N_15870);
or U16421 (N_16421,N_14032,N_14520);
nand U16422 (N_16422,N_14211,N_14572);
nand U16423 (N_16423,N_15837,N_14363);
xor U16424 (N_16424,N_14879,N_14229);
nor U16425 (N_16425,N_14584,N_15063);
xnor U16426 (N_16426,N_15685,N_14842);
or U16427 (N_16427,N_15917,N_15541);
or U16428 (N_16428,N_15954,N_15649);
xor U16429 (N_16429,N_15045,N_14125);
xnor U16430 (N_16430,N_15377,N_15394);
nand U16431 (N_16431,N_15531,N_15069);
and U16432 (N_16432,N_15586,N_14460);
nand U16433 (N_16433,N_14014,N_15776);
nor U16434 (N_16434,N_14769,N_15842);
nand U16435 (N_16435,N_14021,N_14762);
or U16436 (N_16436,N_14480,N_14338);
xnor U16437 (N_16437,N_14316,N_14048);
nand U16438 (N_16438,N_15425,N_15329);
nand U16439 (N_16439,N_15032,N_14901);
nand U16440 (N_16440,N_14171,N_14024);
and U16441 (N_16441,N_14147,N_14366);
or U16442 (N_16442,N_14502,N_14256);
nor U16443 (N_16443,N_14656,N_15832);
nor U16444 (N_16444,N_14564,N_14561);
nand U16445 (N_16445,N_14878,N_15401);
or U16446 (N_16446,N_14405,N_14587);
xnor U16447 (N_16447,N_14965,N_14027);
nand U16448 (N_16448,N_15885,N_15274);
nor U16449 (N_16449,N_14610,N_15747);
nor U16450 (N_16450,N_14626,N_15031);
nand U16451 (N_16451,N_14310,N_15215);
nand U16452 (N_16452,N_14874,N_14031);
and U16453 (N_16453,N_15289,N_14417);
xor U16454 (N_16454,N_14446,N_15726);
or U16455 (N_16455,N_14738,N_14960);
or U16456 (N_16456,N_15125,N_14699);
nand U16457 (N_16457,N_15634,N_14193);
xor U16458 (N_16458,N_15419,N_14776);
nand U16459 (N_16459,N_14941,N_14845);
nor U16460 (N_16460,N_15636,N_14848);
and U16461 (N_16461,N_15087,N_15172);
or U16462 (N_16462,N_14304,N_14144);
xor U16463 (N_16463,N_14277,N_15926);
or U16464 (N_16464,N_14189,N_15869);
xor U16465 (N_16465,N_14207,N_14747);
nor U16466 (N_16466,N_14158,N_15306);
and U16467 (N_16467,N_14373,N_15339);
nor U16468 (N_16468,N_14424,N_14233);
and U16469 (N_16469,N_14887,N_14816);
nand U16470 (N_16470,N_14161,N_15956);
xor U16471 (N_16471,N_15780,N_14922);
or U16472 (N_16472,N_14210,N_14952);
and U16473 (N_16473,N_14722,N_14368);
nand U16474 (N_16474,N_15439,N_14456);
nand U16475 (N_16475,N_15078,N_15337);
nand U16476 (N_16476,N_15495,N_15406);
and U16477 (N_16477,N_15004,N_15469);
xor U16478 (N_16478,N_14886,N_14782);
and U16479 (N_16479,N_15445,N_15109);
nor U16480 (N_16480,N_14025,N_15169);
xor U16481 (N_16481,N_14487,N_15560);
xnor U16482 (N_16482,N_14395,N_15165);
xor U16483 (N_16483,N_14112,N_15230);
nor U16484 (N_16484,N_15348,N_15392);
nor U16485 (N_16485,N_15208,N_15309);
nand U16486 (N_16486,N_14679,N_15608);
xnor U16487 (N_16487,N_15575,N_14463);
xor U16488 (N_16488,N_15902,N_14439);
nand U16489 (N_16489,N_15455,N_14537);
nand U16490 (N_16490,N_14550,N_14351);
or U16491 (N_16491,N_14020,N_15201);
or U16492 (N_16492,N_14690,N_14971);
and U16493 (N_16493,N_15034,N_15720);
nand U16494 (N_16494,N_14318,N_15587);
nor U16495 (N_16495,N_14721,N_14050);
or U16496 (N_16496,N_14002,N_15571);
xnor U16497 (N_16497,N_14995,N_14205);
nand U16498 (N_16498,N_14484,N_15517);
or U16499 (N_16499,N_14568,N_14116);
nor U16500 (N_16500,N_15084,N_15210);
or U16501 (N_16501,N_14043,N_14532);
and U16502 (N_16502,N_14258,N_14320);
or U16503 (N_16503,N_14953,N_14729);
nor U16504 (N_16504,N_14574,N_14966);
nand U16505 (N_16505,N_14226,N_14547);
and U16506 (N_16506,N_15574,N_14608);
xor U16507 (N_16507,N_14928,N_15255);
and U16508 (N_16508,N_15442,N_14961);
xnor U16509 (N_16509,N_15386,N_15124);
and U16510 (N_16510,N_15064,N_15212);
nor U16511 (N_16511,N_14440,N_15107);
nand U16512 (N_16512,N_15432,N_14601);
xnor U16513 (N_16513,N_15006,N_15225);
or U16514 (N_16514,N_14349,N_15326);
nand U16515 (N_16515,N_15804,N_14386);
nand U16516 (N_16516,N_14182,N_15498);
and U16517 (N_16517,N_14620,N_14379);
or U16518 (N_16518,N_15002,N_15736);
nor U16519 (N_16519,N_15501,N_15493);
and U16520 (N_16520,N_15251,N_15806);
xor U16521 (N_16521,N_14138,N_15528);
nand U16522 (N_16522,N_14221,N_15766);
nand U16523 (N_16523,N_15581,N_15365);
nand U16524 (N_16524,N_15246,N_15188);
or U16525 (N_16525,N_14703,N_14526);
xnor U16526 (N_16526,N_14954,N_15472);
nand U16527 (N_16527,N_14194,N_15191);
nand U16528 (N_16528,N_14516,N_14438);
and U16529 (N_16529,N_14464,N_14444);
or U16530 (N_16530,N_15285,N_15298);
nand U16531 (N_16531,N_14168,N_15356);
xnor U16532 (N_16532,N_14864,N_14548);
nor U16533 (N_16533,N_15502,N_14982);
or U16534 (N_16534,N_14140,N_14546);
nor U16535 (N_16535,N_15682,N_14423);
nor U16536 (N_16536,N_15888,N_14761);
or U16537 (N_16537,N_15106,N_15533);
or U16538 (N_16538,N_14371,N_15666);
xor U16539 (N_16539,N_14625,N_15786);
or U16540 (N_16540,N_14060,N_15118);
nand U16541 (N_16541,N_14384,N_14650);
nand U16542 (N_16542,N_15061,N_15410);
nor U16543 (N_16543,N_15444,N_15016);
nand U16544 (N_16544,N_15968,N_14556);
or U16545 (N_16545,N_14090,N_14391);
nand U16546 (N_16546,N_15213,N_14501);
nor U16547 (N_16547,N_14238,N_14259);
nor U16548 (N_16548,N_14830,N_14951);
nand U16549 (N_16549,N_14552,N_14888);
or U16550 (N_16550,N_14206,N_15241);
xor U16551 (N_16551,N_14092,N_14571);
xnor U16552 (N_16552,N_14595,N_14613);
and U16553 (N_16553,N_15921,N_14628);
nand U16554 (N_16554,N_15536,N_15994);
or U16555 (N_16555,N_14276,N_14529);
xnor U16556 (N_16556,N_15754,N_15139);
or U16557 (N_16557,N_14335,N_15179);
xnor U16558 (N_16558,N_15344,N_15283);
nor U16559 (N_16559,N_14156,N_15403);
nand U16560 (N_16560,N_14597,N_14126);
nand U16561 (N_16561,N_15307,N_15589);
nor U16562 (N_16562,N_14843,N_15460);
nand U16563 (N_16563,N_15011,N_14920);
and U16564 (N_16564,N_14346,N_15770);
nor U16565 (N_16565,N_15448,N_15181);
nor U16566 (N_16566,N_15205,N_15811);
nand U16567 (N_16567,N_15314,N_15046);
and U16568 (N_16568,N_15416,N_15113);
nor U16569 (N_16569,N_14524,N_15639);
or U16570 (N_16570,N_15048,N_15562);
xor U16571 (N_16571,N_15549,N_14914);
nand U16572 (N_16572,N_15244,N_14102);
or U16573 (N_16573,N_14153,N_14497);
and U16574 (N_16574,N_14013,N_14362);
xor U16575 (N_16575,N_14506,N_15878);
xnor U16576 (N_16576,N_14402,N_15701);
nor U16577 (N_16577,N_15788,N_15997);
nor U16578 (N_16578,N_15927,N_15606);
xor U16579 (N_16579,N_14838,N_15957);
and U16580 (N_16580,N_14748,N_14040);
and U16581 (N_16581,N_15163,N_14174);
nand U16582 (N_16582,N_15176,N_15007);
and U16583 (N_16583,N_14412,N_15680);
or U16584 (N_16584,N_14239,N_15872);
xnor U16585 (N_16585,N_15523,N_15177);
nand U16586 (N_16586,N_14465,N_14037);
xor U16587 (N_16587,N_14176,N_15695);
and U16588 (N_16588,N_14019,N_14165);
and U16589 (N_16589,N_15330,N_14542);
nand U16590 (N_16590,N_14098,N_14964);
or U16591 (N_16591,N_15267,N_15740);
or U16592 (N_16592,N_15600,N_14091);
and U16593 (N_16593,N_14331,N_14309);
nor U16594 (N_16594,N_14522,N_14742);
and U16595 (N_16595,N_14383,N_15833);
xnor U16596 (N_16596,N_14018,N_15300);
and U16597 (N_16597,N_15412,N_15333);
nor U16598 (N_16598,N_15219,N_15779);
nand U16599 (N_16599,N_14492,N_15584);
and U16600 (N_16600,N_14706,N_15081);
or U16601 (N_16601,N_15355,N_14931);
and U16602 (N_16602,N_15140,N_14660);
nor U16603 (N_16603,N_15681,N_15050);
nor U16604 (N_16604,N_14583,N_15376);
and U16605 (N_16605,N_15152,N_14940);
xor U16606 (N_16606,N_14749,N_15461);
nand U16607 (N_16607,N_14802,N_15756);
and U16608 (N_16608,N_15840,N_15617);
and U16609 (N_16609,N_14939,N_14702);
xnor U16610 (N_16610,N_14896,N_14779);
and U16611 (N_16611,N_14442,N_14619);
nor U16612 (N_16612,N_14781,N_15327);
nand U16613 (N_16613,N_14403,N_14162);
or U16614 (N_16614,N_15462,N_14596);
xor U16615 (N_16615,N_15138,N_14086);
or U16616 (N_16616,N_14591,N_15076);
nand U16617 (N_16617,N_14279,N_15988);
nor U16618 (N_16618,N_14157,N_15696);
nand U16619 (N_16619,N_14184,N_14255);
and U16620 (N_16620,N_14411,N_15051);
nor U16621 (N_16621,N_15699,N_15966);
xor U16622 (N_16622,N_14655,N_14185);
nor U16623 (N_16623,N_14930,N_14837);
nor U16624 (N_16624,N_15449,N_15569);
nand U16625 (N_16625,N_15722,N_15027);
or U16626 (N_16626,N_14166,N_15282);
nor U16627 (N_16627,N_15709,N_14061);
xor U16628 (N_16628,N_15692,N_14658);
and U16629 (N_16629,N_14302,N_14352);
xor U16630 (N_16630,N_15915,N_15240);
nand U16631 (N_16631,N_15835,N_14046);
nor U16632 (N_16632,N_14607,N_15678);
and U16633 (N_16633,N_15873,N_14716);
xor U16634 (N_16634,N_15033,N_15800);
nor U16635 (N_16635,N_15768,N_14376);
xor U16636 (N_16636,N_14649,N_14022);
or U16637 (N_16637,N_15573,N_15082);
nor U16638 (N_16638,N_15923,N_14489);
nand U16639 (N_16639,N_14408,N_15183);
xnor U16640 (N_16640,N_14835,N_15491);
nor U16641 (N_16641,N_15506,N_15967);
nor U16642 (N_16642,N_14857,N_15194);
nand U16643 (N_16643,N_15079,N_14263);
nor U16644 (N_16644,N_15558,N_15342);
and U16645 (N_16645,N_15919,N_15200);
or U16646 (N_16646,N_15198,N_14345);
xor U16647 (N_16647,N_15601,N_14006);
nand U16648 (N_16648,N_14578,N_14400);
or U16649 (N_16649,N_14332,N_14943);
nor U16650 (N_16650,N_15145,N_15216);
nand U16651 (N_16651,N_15922,N_14172);
or U16652 (N_16652,N_15937,N_15144);
and U16653 (N_16653,N_14089,N_14141);
and U16654 (N_16654,N_14701,N_15518);
or U16655 (N_16655,N_15545,N_14521);
nor U16656 (N_16656,N_15433,N_15451);
and U16657 (N_16657,N_14509,N_15415);
xor U16658 (N_16658,N_14353,N_14676);
or U16659 (N_16659,N_15099,N_14426);
nand U16660 (N_16660,N_15945,N_14682);
nor U16661 (N_16661,N_14605,N_14334);
and U16662 (N_16662,N_15687,N_14039);
or U16663 (N_16663,N_15662,N_15947);
nand U16664 (N_16664,N_14110,N_15503);
and U16665 (N_16665,N_14430,N_14016);
and U16666 (N_16666,N_15684,N_15952);
xor U16667 (N_16667,N_15426,N_14148);
nor U16668 (N_16668,N_14977,N_15446);
xor U16669 (N_16669,N_14289,N_14612);
nor U16670 (N_16670,N_14818,N_14203);
xnor U16671 (N_16671,N_14651,N_14947);
nor U16672 (N_16672,N_14240,N_15990);
or U16673 (N_16673,N_15646,N_15269);
and U16674 (N_16674,N_15429,N_15475);
xor U16675 (N_16675,N_14419,N_14633);
xnor U16676 (N_16676,N_15918,N_14009);
or U16677 (N_16677,N_14970,N_14431);
nand U16678 (N_16678,N_14833,N_14700);
nand U16679 (N_16679,N_14270,N_14209);
or U16680 (N_16680,N_14152,N_15810);
nand U16681 (N_16681,N_15935,N_15876);
xor U16682 (N_16682,N_14200,N_15170);
xor U16683 (N_16683,N_15982,N_15041);
and U16684 (N_16684,N_14652,N_15764);
nor U16685 (N_16685,N_14892,N_15512);
nor U16686 (N_16686,N_15336,N_15232);
nor U16687 (N_16687,N_15496,N_15056);
xor U16688 (N_16688,N_15487,N_14778);
and U16689 (N_16689,N_14269,N_14798);
and U16690 (N_16690,N_14361,N_14709);
xnor U16691 (N_16691,N_15263,N_15039);
xnor U16692 (N_16692,N_15955,N_14474);
nor U16693 (N_16693,N_14394,N_15570);
xor U16694 (N_16694,N_15436,N_14219);
nand U16695 (N_16695,N_14491,N_15821);
or U16696 (N_16696,N_14870,N_14186);
nor U16697 (N_16697,N_14167,N_14113);
xnor U16698 (N_16698,N_15605,N_15193);
nor U16699 (N_16699,N_15794,N_14560);
nand U16700 (N_16700,N_14508,N_15062);
xor U16701 (N_16701,N_14232,N_15237);
nor U16702 (N_16702,N_14946,N_15863);
and U16703 (N_16703,N_14128,N_14638);
nand U16704 (N_16704,N_15750,N_15802);
nor U16705 (N_16705,N_15091,N_14222);
xor U16706 (N_16706,N_14885,N_14265);
xnor U16707 (N_16707,N_15287,N_14085);
or U16708 (N_16708,N_15530,N_14615);
xor U16709 (N_16709,N_14657,N_15332);
nor U16710 (N_16710,N_15630,N_15631);
nand U16711 (N_16711,N_14045,N_14241);
nor U16712 (N_16712,N_14217,N_15801);
nor U16713 (N_16713,N_14717,N_14737);
or U16714 (N_16714,N_14925,N_14105);
nor U16715 (N_16715,N_15713,N_14871);
or U16716 (N_16716,N_14202,N_14540);
or U16717 (N_16717,N_15025,N_14545);
nand U16718 (N_16718,N_15653,N_14740);
nand U16719 (N_16719,N_14891,N_14023);
or U16720 (N_16720,N_15651,N_15400);
nand U16721 (N_16721,N_14421,N_15126);
and U16722 (N_16722,N_14518,N_14472);
nor U16723 (N_16723,N_14916,N_15676);
or U16724 (N_16724,N_15909,N_15748);
nor U16725 (N_16725,N_15090,N_14957);
nor U16726 (N_16726,N_15075,N_14127);
and U16727 (N_16727,N_14119,N_14704);
and U16728 (N_16728,N_15762,N_15829);
nand U16729 (N_16729,N_15576,N_14354);
or U16730 (N_16730,N_14029,N_14617);
xnor U16731 (N_16731,N_15879,N_15594);
nand U16732 (N_16732,N_15132,N_15227);
and U16733 (N_16733,N_15895,N_15949);
and U16734 (N_16734,N_15580,N_15980);
nand U16735 (N_16735,N_15544,N_14095);
or U16736 (N_16736,N_15474,N_14278);
or U16737 (N_16737,N_14035,N_14875);
nand U16738 (N_16738,N_15903,N_15658);
and U16739 (N_16739,N_14938,N_14713);
nor U16740 (N_16740,N_14429,N_14956);
nor U16741 (N_16741,N_14758,N_15086);
nand U16742 (N_16742,N_14784,N_15178);
and U16743 (N_16743,N_14249,N_14058);
nand U16744 (N_16744,N_15303,N_14543);
and U16745 (N_16745,N_14624,N_15470);
nand U16746 (N_16746,N_15486,N_15288);
nor U16747 (N_16747,N_15221,N_15057);
nor U16748 (N_16748,N_15677,N_15422);
or U16749 (N_16749,N_14825,N_15912);
nor U16750 (N_16750,N_15243,N_15271);
xor U16751 (N_16751,N_14470,N_15362);
nor U16752 (N_16752,N_15976,N_14198);
xnor U16753 (N_16753,N_14882,N_15209);
xnor U16754 (N_16754,N_15660,N_14630);
or U16755 (N_16755,N_14298,N_15629);
nand U16756 (N_16756,N_15497,N_15797);
nand U16757 (N_16757,N_15731,N_14096);
nand U16758 (N_16758,N_15505,N_15250);
and U16759 (N_16759,N_15599,N_15094);
nor U16760 (N_16760,N_15466,N_14654);
and U16761 (N_16761,N_14898,N_14873);
nand U16762 (N_16762,N_15089,N_15595);
or U16763 (N_16763,N_15217,N_14122);
or U16764 (N_16764,N_15852,N_15932);
or U16765 (N_16765,N_15364,N_14746);
or U16766 (N_16766,N_14592,N_14855);
nor U16767 (N_16767,N_15424,N_14598);
xor U16768 (N_16768,N_15884,N_14339);
nor U16769 (N_16769,N_15626,N_15343);
xnor U16770 (N_16770,N_15128,N_14114);
nor U16771 (N_16771,N_15149,N_14724);
or U16772 (N_16772,N_15331,N_15865);
nand U16773 (N_16773,N_14756,N_14017);
xnor U16774 (N_16774,N_15702,N_15066);
or U16775 (N_16775,N_14582,N_15238);
nand U16776 (N_16776,N_15360,N_15103);
xnor U16777 (N_16777,N_14467,N_15098);
nor U16778 (N_16778,N_14300,N_14034);
nor U16779 (N_16779,N_15236,N_14097);
or U16780 (N_16780,N_15375,N_15635);
or U16781 (N_16781,N_15805,N_15349);
nor U16782 (N_16782,N_14199,N_14811);
or U16783 (N_16783,N_15669,N_14932);
nor U16784 (N_16784,N_14780,N_15619);
nor U16785 (N_16785,N_15733,N_14944);
xor U16786 (N_16786,N_14507,N_15218);
or U16787 (N_16787,N_14183,N_14832);
nand U16788 (N_16788,N_15657,N_15085);
xor U16789 (N_16789,N_15450,N_15644);
or U16790 (N_16790,N_15420,N_15310);
nor U16791 (N_16791,N_14056,N_15354);
nand U16792 (N_16792,N_14580,N_14569);
nor U16793 (N_16793,N_14436,N_15357);
nand U16794 (N_16794,N_14360,N_14733);
or U16795 (N_16795,N_14525,N_15345);
or U16796 (N_16796,N_15665,N_14099);
or U16797 (N_16797,N_15154,N_15951);
nor U16798 (N_16798,N_14851,N_15689);
and U16799 (N_16799,N_14344,N_14566);
nand U16800 (N_16800,N_14225,N_14192);
xor U16801 (N_16801,N_14563,N_14861);
or U16802 (N_16802,N_14663,N_15499);
xnor U16803 (N_16803,N_14824,N_15252);
nor U16804 (N_16804,N_15438,N_15610);
nand U16805 (N_16805,N_14364,N_14000);
or U16806 (N_16806,N_14342,N_14077);
xor U16807 (N_16807,N_15223,N_14696);
and U16808 (N_16808,N_15297,N_14057);
nor U16809 (N_16809,N_14744,N_15510);
or U16810 (N_16810,N_14823,N_15974);
nand U16811 (N_16811,N_15708,N_14809);
and U16812 (N_16812,N_15705,N_14136);
nor U16813 (N_16813,N_15965,N_15719);
nand U16814 (N_16814,N_15752,N_14659);
xnor U16815 (N_16815,N_14041,N_14877);
and U16816 (N_16816,N_15417,N_15414);
nor U16817 (N_16817,N_14055,N_14297);
nor U16818 (N_16818,N_15683,N_15065);
or U16819 (N_16819,N_14359,N_15117);
or U16820 (N_16820,N_15622,N_14042);
nand U16821 (N_16821,N_14984,N_15338);
or U16822 (N_16822,N_14581,N_14441);
nand U16823 (N_16823,N_15913,N_15930);
and U16824 (N_16824,N_14170,N_15950);
or U16825 (N_16825,N_15457,N_14872);
and U16826 (N_16826,N_14559,N_14181);
xor U16827 (N_16827,N_14454,N_14059);
nor U16828 (N_16828,N_15774,N_15161);
xor U16829 (N_16829,N_14727,N_14759);
xnor U16830 (N_16830,N_14533,N_14753);
nand U16831 (N_16831,N_14348,N_14485);
nand U16832 (N_16832,N_14745,N_15648);
xor U16833 (N_16833,N_14051,N_14081);
nand U16834 (N_16834,N_15996,N_14589);
or U16835 (N_16835,N_14996,N_15174);
or U16836 (N_16836,N_14834,N_14030);
nor U16837 (N_16837,N_14681,N_15792);
xnor U16838 (N_16838,N_14377,N_14286);
or U16839 (N_16839,N_15334,N_14915);
or U16840 (N_16840,N_15850,N_14135);
nor U16841 (N_16841,N_14675,N_14512);
or U16842 (N_16842,N_14847,N_15256);
nand U16843 (N_16843,N_14785,N_15969);
and U16844 (N_16844,N_15447,N_14720);
nand U16845 (N_16845,N_14775,N_15023);
nor U16846 (N_16846,N_14994,N_15222);
xnor U16847 (N_16847,N_14645,N_14295);
xnor U16848 (N_16848,N_15293,N_14800);
nor U16849 (N_16849,N_15423,N_15537);
and U16850 (N_16850,N_15679,N_14902);
or U16851 (N_16851,N_15925,N_14797);
xnor U16852 (N_16852,N_14108,N_14909);
and U16853 (N_16853,N_14301,N_14755);
nor U16854 (N_16854,N_15192,N_15366);
or U16855 (N_16855,N_15552,N_14247);
nor U16856 (N_16856,N_14683,N_15992);
nor U16857 (N_16857,N_15261,N_15830);
or U16858 (N_16858,N_14340,N_15972);
nor U16859 (N_16859,N_15999,N_15928);
nor U16860 (N_16860,N_15714,N_14076);
or U16861 (N_16861,N_15131,N_15561);
nor U16862 (N_16862,N_15691,N_14149);
and U16863 (N_16863,N_14634,N_14273);
nand U16864 (N_16864,N_15077,N_14319);
and U16865 (N_16865,N_14850,N_15320);
nor U16866 (N_16866,N_14991,N_14160);
nor U16867 (N_16867,N_14230,N_15167);
and U16868 (N_16868,N_15783,N_14629);
and U16869 (N_16869,N_14425,N_14294);
nand U16870 (N_16870,N_15454,N_15324);
nor U16871 (N_16871,N_15621,N_14180);
and U16872 (N_16872,N_14337,N_15755);
nand U16873 (N_16873,N_14590,N_15847);
or U16874 (N_16874,N_14416,N_14667);
xor U16875 (N_16875,N_14003,N_14955);
or U16876 (N_16876,N_15239,N_14422);
nand U16877 (N_16877,N_14692,N_14336);
xor U16878 (N_16878,N_15874,N_14602);
and U16879 (N_16879,N_14678,N_14282);
nor U16880 (N_16880,N_14365,N_14854);
or U16881 (N_16881,N_15352,N_14477);
and U16882 (N_16882,N_14038,N_14962);
xnor U16883 (N_16883,N_15540,N_14792);
xor U16884 (N_16884,N_15319,N_15088);
and U16885 (N_16885,N_15538,N_14687);
nor U16886 (N_16886,N_15313,N_15765);
and U16887 (N_16887,N_15398,N_15390);
nor U16888 (N_16888,N_15807,N_15881);
nand U16889 (N_16889,N_15471,N_14804);
and U16890 (N_16890,N_14449,N_15276);
and U16891 (N_16891,N_15548,N_14826);
nand U16892 (N_16892,N_15978,N_14312);
xnor U16893 (N_16893,N_15047,N_14252);
or U16894 (N_16894,N_15121,N_14585);
nand U16895 (N_16895,N_14517,N_14504);
xnor U16896 (N_16896,N_15134,N_15270);
nand U16897 (N_16897,N_15871,N_15520);
or U16898 (N_16898,N_14100,N_14333);
and U16899 (N_16899,N_14514,N_15384);
nor U16900 (N_16900,N_15020,N_14208);
nand U16901 (N_16901,N_14468,N_15607);
and U16902 (N_16902,N_15831,N_15411);
or U16903 (N_16903,N_14728,N_14355);
nand U16904 (N_16904,N_15686,N_15609);
xnor U16905 (N_16905,N_15367,N_14455);
nand U16906 (N_16906,N_14490,N_15859);
nor U16907 (N_16907,N_14694,N_14062);
nand U16908 (N_16908,N_15321,N_14284);
or U16909 (N_16909,N_14814,N_14969);
xor U16910 (N_16910,N_14457,N_15959);
nor U16911 (N_16911,N_14680,N_14299);
nand U16912 (N_16912,N_14139,N_15825);
nand U16913 (N_16913,N_14358,N_15728);
xor U16914 (N_16914,N_14853,N_14296);
xnor U16915 (N_16915,N_14083,N_14926);
xnor U16916 (N_16916,N_15494,N_14479);
nor U16917 (N_16917,N_15480,N_15305);
or U16918 (N_16918,N_14315,N_14643);
and U16919 (N_16919,N_15958,N_15791);
and U16920 (N_16920,N_14719,N_14049);
or U16921 (N_16921,N_14387,N_14686);
nor U16922 (N_16922,N_15547,N_14341);
nand U16923 (N_16923,N_15637,N_15516);
nor U16924 (N_16924,N_15180,N_14538);
or U16925 (N_16925,N_15838,N_15130);
and U16926 (N_16926,N_14906,N_15441);
or U16927 (N_16927,N_15317,N_15784);
xor U16928 (N_16928,N_15529,N_14535);
nor U16929 (N_16929,N_14551,N_15052);
nand U16930 (N_16930,N_15887,N_15795);
and U16931 (N_16931,N_15758,N_15435);
and U16932 (N_16932,N_15257,N_14234);
xor U16933 (N_16933,N_14865,N_14292);
or U16934 (N_16934,N_15262,N_14918);
and U16935 (N_16935,N_14325,N_14033);
and U16936 (N_16936,N_14313,N_14627);
nand U16937 (N_16937,N_15024,N_14757);
nor U16938 (N_16938,N_15769,N_15661);
xnor U16939 (N_16939,N_15481,N_15703);
nor U16940 (N_16940,N_15524,N_14382);
or U16941 (N_16941,N_15899,N_15761);
nand U16942 (N_16942,N_14796,N_14071);
and U16943 (N_16943,N_15074,N_15160);
nor U16944 (N_16944,N_15633,N_14632);
or U16945 (N_16945,N_14306,N_14451);
and U16946 (N_16946,N_14976,N_15655);
nand U16947 (N_16947,N_15707,N_15408);
nor U16948 (N_16948,N_15942,N_15127);
nor U16949 (N_16949,N_14777,N_15824);
xnor U16950 (N_16950,N_15104,N_15234);
nand U16951 (N_16951,N_14466,N_14245);
nor U16952 (N_16952,N_15206,N_15155);
nand U16953 (N_16953,N_14726,N_14801);
xnor U16954 (N_16954,N_15823,N_15604);
or U16955 (N_16955,N_14212,N_14992);
and U16956 (N_16956,N_14307,N_15670);
and U16957 (N_16957,N_15490,N_14648);
xor U16958 (N_16958,N_14989,N_15934);
xor U16959 (N_16959,N_14054,N_15856);
nor U16960 (N_16960,N_14163,N_15862);
xnor U16961 (N_16961,N_14573,N_14523);
nor U16962 (N_16962,N_14693,N_15782);
or U16963 (N_16963,N_14005,N_14599);
nor U16964 (N_16964,N_14820,N_14677);
nand U16965 (N_16965,N_15883,N_15049);
nand U16966 (N_16966,N_14987,N_14236);
xnor U16967 (N_16967,N_15519,N_15029);
or U16968 (N_16968,N_15003,N_15010);
nand U16969 (N_16969,N_14123,N_15380);
and U16970 (N_16970,N_15229,N_15014);
nor U16971 (N_16971,N_15483,N_14224);
and U16972 (N_16972,N_14448,N_15456);
nand U16973 (N_16973,N_14614,N_15898);
nor U16974 (N_16974,N_15977,N_15907);
and U16975 (N_16975,N_15645,N_14618);
nor U16976 (N_16976,N_15015,N_15312);
or U16977 (N_16977,N_15001,N_15929);
or U16978 (N_16978,N_15295,N_14979);
and U16979 (N_16979,N_15550,N_15729);
and U16980 (N_16980,N_15730,N_15822);
nor U16981 (N_16981,N_15710,N_15796);
xor U16982 (N_16982,N_15304,N_14621);
nand U16983 (N_16983,N_15166,N_14723);
nor U16984 (N_16984,N_14557,N_14499);
nor U16985 (N_16985,N_14808,N_14084);
xnor U16986 (N_16986,N_14392,N_14562);
or U16987 (N_16987,N_14137,N_15944);
and U16988 (N_16988,N_14963,N_14204);
nand U16989 (N_16989,N_15259,N_15984);
and U16990 (N_16990,N_15459,N_14647);
and U16991 (N_16991,N_15652,N_14486);
nand U16992 (N_16992,N_15030,N_14398);
and U16993 (N_16993,N_14109,N_14641);
or U16994 (N_16994,N_15809,N_14646);
and U16995 (N_16995,N_15228,N_15428);
and U16996 (N_16996,N_15443,N_15043);
or U16997 (N_16997,N_14983,N_15936);
nand U16998 (N_16998,N_14653,N_15111);
nor U16999 (N_16999,N_14469,N_15920);
xnor U17000 (N_17000,N_14217,N_15376);
or U17001 (N_17001,N_14767,N_14126);
nor U17002 (N_17002,N_14627,N_15751);
and U17003 (N_17003,N_15791,N_15584);
and U17004 (N_17004,N_15560,N_14352);
nor U17005 (N_17005,N_14069,N_14983);
nor U17006 (N_17006,N_14070,N_15418);
xnor U17007 (N_17007,N_14870,N_15680);
and U17008 (N_17008,N_14197,N_14194);
or U17009 (N_17009,N_15106,N_14914);
nand U17010 (N_17010,N_15670,N_14897);
nor U17011 (N_17011,N_14627,N_14653);
and U17012 (N_17012,N_15221,N_14517);
and U17013 (N_17013,N_14762,N_15853);
xor U17014 (N_17014,N_14538,N_15419);
and U17015 (N_17015,N_14225,N_14252);
xor U17016 (N_17016,N_14620,N_15361);
and U17017 (N_17017,N_15101,N_14680);
or U17018 (N_17018,N_14790,N_14939);
nor U17019 (N_17019,N_15975,N_14120);
nor U17020 (N_17020,N_14356,N_15862);
nand U17021 (N_17021,N_15447,N_14405);
and U17022 (N_17022,N_14869,N_14790);
or U17023 (N_17023,N_15352,N_15748);
or U17024 (N_17024,N_14354,N_14919);
xnor U17025 (N_17025,N_15043,N_14245);
or U17026 (N_17026,N_14505,N_14051);
nand U17027 (N_17027,N_15903,N_14644);
xnor U17028 (N_17028,N_15202,N_14694);
xnor U17029 (N_17029,N_14930,N_14281);
and U17030 (N_17030,N_14389,N_15776);
or U17031 (N_17031,N_15895,N_14514);
or U17032 (N_17032,N_15879,N_15486);
xor U17033 (N_17033,N_15164,N_14068);
and U17034 (N_17034,N_15003,N_14545);
nand U17035 (N_17035,N_15367,N_15869);
xor U17036 (N_17036,N_14186,N_15411);
and U17037 (N_17037,N_15379,N_14293);
or U17038 (N_17038,N_15145,N_15421);
xor U17039 (N_17039,N_14609,N_14322);
nand U17040 (N_17040,N_14975,N_14718);
or U17041 (N_17041,N_14504,N_14970);
nor U17042 (N_17042,N_15745,N_15611);
nor U17043 (N_17043,N_15820,N_15445);
or U17044 (N_17044,N_14794,N_15706);
and U17045 (N_17045,N_15423,N_15011);
and U17046 (N_17046,N_15889,N_14895);
and U17047 (N_17047,N_15848,N_15722);
or U17048 (N_17048,N_15971,N_15042);
xor U17049 (N_17049,N_14076,N_14488);
and U17050 (N_17050,N_15509,N_14023);
nor U17051 (N_17051,N_14698,N_14146);
and U17052 (N_17052,N_15505,N_14229);
or U17053 (N_17053,N_15221,N_15157);
nor U17054 (N_17054,N_15244,N_15499);
nor U17055 (N_17055,N_15639,N_14493);
or U17056 (N_17056,N_14294,N_15372);
nand U17057 (N_17057,N_15318,N_15669);
and U17058 (N_17058,N_15801,N_15974);
nand U17059 (N_17059,N_14922,N_14685);
nor U17060 (N_17060,N_14427,N_15295);
or U17061 (N_17061,N_14002,N_14334);
and U17062 (N_17062,N_15219,N_14755);
and U17063 (N_17063,N_15837,N_15726);
nor U17064 (N_17064,N_15731,N_14624);
xor U17065 (N_17065,N_15831,N_14354);
nand U17066 (N_17066,N_15154,N_15519);
nand U17067 (N_17067,N_14778,N_15069);
and U17068 (N_17068,N_15836,N_14826);
xnor U17069 (N_17069,N_14564,N_15156);
nand U17070 (N_17070,N_14157,N_14165);
and U17071 (N_17071,N_15009,N_14269);
xor U17072 (N_17072,N_15169,N_15937);
and U17073 (N_17073,N_14439,N_15430);
xnor U17074 (N_17074,N_15470,N_14127);
nor U17075 (N_17075,N_14327,N_15321);
and U17076 (N_17076,N_15618,N_15127);
and U17077 (N_17077,N_15322,N_14123);
or U17078 (N_17078,N_15839,N_14456);
nor U17079 (N_17079,N_14121,N_15978);
and U17080 (N_17080,N_15523,N_15730);
or U17081 (N_17081,N_14210,N_15852);
nand U17082 (N_17082,N_15156,N_14129);
or U17083 (N_17083,N_15216,N_14625);
or U17084 (N_17084,N_15533,N_14069);
or U17085 (N_17085,N_14623,N_15795);
and U17086 (N_17086,N_14694,N_15320);
nand U17087 (N_17087,N_15563,N_14990);
xor U17088 (N_17088,N_14051,N_15024);
xor U17089 (N_17089,N_14733,N_15684);
and U17090 (N_17090,N_14499,N_15938);
xnor U17091 (N_17091,N_14727,N_15110);
nand U17092 (N_17092,N_14231,N_15343);
and U17093 (N_17093,N_14618,N_14802);
and U17094 (N_17094,N_14848,N_14910);
xnor U17095 (N_17095,N_15539,N_14498);
nor U17096 (N_17096,N_15182,N_14070);
and U17097 (N_17097,N_15764,N_15353);
nor U17098 (N_17098,N_14753,N_15557);
nor U17099 (N_17099,N_15493,N_14507);
or U17100 (N_17100,N_14094,N_15704);
xor U17101 (N_17101,N_14783,N_14628);
and U17102 (N_17102,N_14210,N_15168);
nand U17103 (N_17103,N_15651,N_15110);
or U17104 (N_17104,N_15962,N_15310);
and U17105 (N_17105,N_14951,N_14551);
xnor U17106 (N_17106,N_15582,N_15627);
xnor U17107 (N_17107,N_14027,N_15720);
nor U17108 (N_17108,N_15931,N_14123);
nor U17109 (N_17109,N_14942,N_15637);
nand U17110 (N_17110,N_14748,N_14740);
nand U17111 (N_17111,N_14084,N_14715);
and U17112 (N_17112,N_15083,N_15330);
xnor U17113 (N_17113,N_15735,N_14787);
or U17114 (N_17114,N_15450,N_14029);
nand U17115 (N_17115,N_14417,N_14857);
nor U17116 (N_17116,N_14100,N_14275);
or U17117 (N_17117,N_15152,N_15766);
nor U17118 (N_17118,N_15826,N_15320);
nor U17119 (N_17119,N_15771,N_14995);
nand U17120 (N_17120,N_14600,N_15756);
nand U17121 (N_17121,N_14120,N_14210);
nor U17122 (N_17122,N_15272,N_14602);
xor U17123 (N_17123,N_14137,N_14980);
xor U17124 (N_17124,N_15233,N_15623);
or U17125 (N_17125,N_15113,N_15924);
and U17126 (N_17126,N_14102,N_15110);
and U17127 (N_17127,N_15945,N_14616);
nand U17128 (N_17128,N_15001,N_14725);
xnor U17129 (N_17129,N_15426,N_14566);
nand U17130 (N_17130,N_15556,N_14613);
nand U17131 (N_17131,N_14815,N_15583);
nor U17132 (N_17132,N_15357,N_14413);
or U17133 (N_17133,N_15602,N_15116);
and U17134 (N_17134,N_15462,N_14786);
nand U17135 (N_17135,N_14495,N_15967);
or U17136 (N_17136,N_15115,N_15699);
nand U17137 (N_17137,N_14761,N_14240);
nand U17138 (N_17138,N_15368,N_14420);
xnor U17139 (N_17139,N_15956,N_15461);
nor U17140 (N_17140,N_15971,N_14994);
or U17141 (N_17141,N_15738,N_14832);
xnor U17142 (N_17142,N_15940,N_15030);
or U17143 (N_17143,N_14089,N_15721);
or U17144 (N_17144,N_14025,N_15858);
or U17145 (N_17145,N_14075,N_14555);
and U17146 (N_17146,N_14667,N_15483);
xnor U17147 (N_17147,N_14614,N_14286);
nor U17148 (N_17148,N_14531,N_14562);
or U17149 (N_17149,N_15718,N_15618);
nand U17150 (N_17150,N_14987,N_14739);
xor U17151 (N_17151,N_15907,N_14836);
and U17152 (N_17152,N_14830,N_15535);
nand U17153 (N_17153,N_15478,N_15078);
xnor U17154 (N_17154,N_15330,N_14706);
and U17155 (N_17155,N_14492,N_15034);
or U17156 (N_17156,N_15915,N_15415);
and U17157 (N_17157,N_15856,N_14321);
and U17158 (N_17158,N_15311,N_14714);
or U17159 (N_17159,N_15990,N_15147);
xnor U17160 (N_17160,N_15955,N_15747);
and U17161 (N_17161,N_14767,N_14699);
nand U17162 (N_17162,N_15375,N_15913);
and U17163 (N_17163,N_15289,N_14731);
nand U17164 (N_17164,N_15859,N_15654);
and U17165 (N_17165,N_15619,N_15840);
and U17166 (N_17166,N_15001,N_15215);
xor U17167 (N_17167,N_15220,N_15643);
nor U17168 (N_17168,N_14544,N_15109);
or U17169 (N_17169,N_14592,N_15274);
nand U17170 (N_17170,N_14152,N_14802);
and U17171 (N_17171,N_15144,N_14691);
nor U17172 (N_17172,N_15980,N_14389);
nand U17173 (N_17173,N_15800,N_15438);
nand U17174 (N_17174,N_15001,N_15220);
nand U17175 (N_17175,N_14293,N_15691);
and U17176 (N_17176,N_15443,N_15599);
xor U17177 (N_17177,N_15178,N_14284);
xnor U17178 (N_17178,N_14037,N_14521);
or U17179 (N_17179,N_15640,N_14481);
nor U17180 (N_17180,N_14736,N_14168);
nor U17181 (N_17181,N_15981,N_15856);
nand U17182 (N_17182,N_14449,N_14644);
or U17183 (N_17183,N_14911,N_15631);
xnor U17184 (N_17184,N_14404,N_14386);
xnor U17185 (N_17185,N_14552,N_14094);
or U17186 (N_17186,N_14241,N_14975);
and U17187 (N_17187,N_15209,N_15367);
nor U17188 (N_17188,N_15770,N_15585);
xnor U17189 (N_17189,N_15496,N_14591);
nor U17190 (N_17190,N_15234,N_14331);
or U17191 (N_17191,N_14326,N_14537);
and U17192 (N_17192,N_15282,N_15503);
or U17193 (N_17193,N_14224,N_14513);
nor U17194 (N_17194,N_15946,N_14481);
nor U17195 (N_17195,N_15858,N_14904);
nor U17196 (N_17196,N_15579,N_14332);
and U17197 (N_17197,N_15535,N_15789);
or U17198 (N_17198,N_15100,N_14343);
xnor U17199 (N_17199,N_14024,N_14255);
and U17200 (N_17200,N_14848,N_14147);
xnor U17201 (N_17201,N_14239,N_15274);
nor U17202 (N_17202,N_14038,N_14669);
xnor U17203 (N_17203,N_14255,N_15537);
nand U17204 (N_17204,N_14883,N_14590);
nand U17205 (N_17205,N_15040,N_15086);
nor U17206 (N_17206,N_14091,N_15406);
and U17207 (N_17207,N_14221,N_15180);
or U17208 (N_17208,N_14248,N_14626);
or U17209 (N_17209,N_14765,N_14085);
or U17210 (N_17210,N_15193,N_14007);
xnor U17211 (N_17211,N_14453,N_14326);
xnor U17212 (N_17212,N_14827,N_14102);
or U17213 (N_17213,N_14357,N_15864);
and U17214 (N_17214,N_14110,N_15026);
xnor U17215 (N_17215,N_14924,N_15406);
and U17216 (N_17216,N_14659,N_15155);
xor U17217 (N_17217,N_15650,N_14329);
or U17218 (N_17218,N_15495,N_15298);
nand U17219 (N_17219,N_14926,N_14946);
and U17220 (N_17220,N_15280,N_14104);
and U17221 (N_17221,N_14212,N_15329);
nand U17222 (N_17222,N_15451,N_14449);
and U17223 (N_17223,N_15721,N_15118);
and U17224 (N_17224,N_15194,N_14446);
and U17225 (N_17225,N_15310,N_14423);
and U17226 (N_17226,N_14216,N_14754);
nor U17227 (N_17227,N_14813,N_15039);
nand U17228 (N_17228,N_14158,N_14966);
xnor U17229 (N_17229,N_15373,N_14455);
and U17230 (N_17230,N_15740,N_15995);
or U17231 (N_17231,N_15983,N_15948);
xor U17232 (N_17232,N_15345,N_15182);
nor U17233 (N_17233,N_15492,N_14087);
xnor U17234 (N_17234,N_14146,N_15615);
xnor U17235 (N_17235,N_14391,N_14243);
or U17236 (N_17236,N_14504,N_15169);
nor U17237 (N_17237,N_14636,N_15236);
nand U17238 (N_17238,N_14541,N_15552);
and U17239 (N_17239,N_14297,N_15132);
and U17240 (N_17240,N_15694,N_14008);
nor U17241 (N_17241,N_14240,N_15698);
nor U17242 (N_17242,N_15983,N_15394);
or U17243 (N_17243,N_14133,N_15142);
xor U17244 (N_17244,N_14474,N_14111);
xor U17245 (N_17245,N_14426,N_14595);
and U17246 (N_17246,N_15770,N_14103);
xor U17247 (N_17247,N_14584,N_14419);
and U17248 (N_17248,N_14824,N_15635);
or U17249 (N_17249,N_15138,N_15260);
or U17250 (N_17250,N_15576,N_14706);
or U17251 (N_17251,N_14693,N_15960);
xnor U17252 (N_17252,N_14715,N_14258);
nor U17253 (N_17253,N_14648,N_14745);
nor U17254 (N_17254,N_15126,N_14867);
and U17255 (N_17255,N_14974,N_15474);
xnor U17256 (N_17256,N_14740,N_15549);
and U17257 (N_17257,N_15631,N_15860);
nand U17258 (N_17258,N_15148,N_15138);
xor U17259 (N_17259,N_14979,N_15887);
xor U17260 (N_17260,N_15523,N_15759);
and U17261 (N_17261,N_14637,N_14718);
nor U17262 (N_17262,N_14311,N_15497);
and U17263 (N_17263,N_15748,N_15094);
or U17264 (N_17264,N_14378,N_15828);
nor U17265 (N_17265,N_15168,N_14151);
xor U17266 (N_17266,N_15547,N_15787);
nor U17267 (N_17267,N_14990,N_14662);
nand U17268 (N_17268,N_15230,N_15777);
and U17269 (N_17269,N_15805,N_15422);
nor U17270 (N_17270,N_14046,N_14136);
xnor U17271 (N_17271,N_15756,N_14466);
nor U17272 (N_17272,N_14444,N_14253);
or U17273 (N_17273,N_15464,N_15307);
xnor U17274 (N_17274,N_14245,N_14942);
and U17275 (N_17275,N_15082,N_15658);
xor U17276 (N_17276,N_15465,N_14093);
xor U17277 (N_17277,N_14312,N_14665);
nor U17278 (N_17278,N_14352,N_15636);
or U17279 (N_17279,N_14354,N_15810);
nor U17280 (N_17280,N_14725,N_15212);
nand U17281 (N_17281,N_15687,N_15906);
nor U17282 (N_17282,N_14570,N_15674);
or U17283 (N_17283,N_14829,N_14167);
nand U17284 (N_17284,N_14217,N_14359);
and U17285 (N_17285,N_14988,N_15026);
or U17286 (N_17286,N_15565,N_14703);
or U17287 (N_17287,N_15464,N_14672);
nand U17288 (N_17288,N_15707,N_14834);
xnor U17289 (N_17289,N_14866,N_15052);
xor U17290 (N_17290,N_15659,N_15259);
nand U17291 (N_17291,N_15919,N_15175);
and U17292 (N_17292,N_15552,N_15832);
and U17293 (N_17293,N_14760,N_14577);
and U17294 (N_17294,N_14043,N_15890);
or U17295 (N_17295,N_14201,N_15604);
xor U17296 (N_17296,N_15889,N_14877);
and U17297 (N_17297,N_14741,N_15626);
xnor U17298 (N_17298,N_14838,N_15704);
nand U17299 (N_17299,N_14532,N_15031);
and U17300 (N_17300,N_14352,N_14376);
nand U17301 (N_17301,N_14082,N_15460);
and U17302 (N_17302,N_15510,N_15759);
xnor U17303 (N_17303,N_14615,N_15922);
xor U17304 (N_17304,N_14020,N_15223);
and U17305 (N_17305,N_15188,N_14490);
or U17306 (N_17306,N_14801,N_15620);
and U17307 (N_17307,N_14205,N_14795);
and U17308 (N_17308,N_14533,N_14398);
xnor U17309 (N_17309,N_14929,N_14968);
or U17310 (N_17310,N_15271,N_15617);
or U17311 (N_17311,N_15219,N_14588);
or U17312 (N_17312,N_15514,N_15519);
nor U17313 (N_17313,N_14101,N_15900);
and U17314 (N_17314,N_15886,N_14891);
or U17315 (N_17315,N_14620,N_14843);
nor U17316 (N_17316,N_15958,N_14723);
xnor U17317 (N_17317,N_14325,N_14790);
and U17318 (N_17318,N_15640,N_14193);
xor U17319 (N_17319,N_14916,N_14748);
nand U17320 (N_17320,N_14854,N_15501);
nor U17321 (N_17321,N_14334,N_14212);
nor U17322 (N_17322,N_15628,N_15884);
nor U17323 (N_17323,N_15896,N_15307);
xor U17324 (N_17324,N_14907,N_14116);
nand U17325 (N_17325,N_15132,N_14903);
and U17326 (N_17326,N_14610,N_15716);
nand U17327 (N_17327,N_15173,N_14099);
or U17328 (N_17328,N_15034,N_14805);
xor U17329 (N_17329,N_14619,N_14033);
nor U17330 (N_17330,N_15403,N_14962);
nor U17331 (N_17331,N_14882,N_14685);
nor U17332 (N_17332,N_15931,N_14917);
nand U17333 (N_17333,N_15056,N_15761);
or U17334 (N_17334,N_14085,N_15769);
and U17335 (N_17335,N_14540,N_15518);
nor U17336 (N_17336,N_15821,N_15332);
nor U17337 (N_17337,N_15003,N_14386);
nor U17338 (N_17338,N_14257,N_14246);
or U17339 (N_17339,N_15056,N_15827);
nand U17340 (N_17340,N_15489,N_14286);
and U17341 (N_17341,N_14022,N_14232);
nor U17342 (N_17342,N_15385,N_14190);
nor U17343 (N_17343,N_14493,N_15029);
and U17344 (N_17344,N_15504,N_14858);
and U17345 (N_17345,N_14318,N_14675);
xor U17346 (N_17346,N_14439,N_15941);
or U17347 (N_17347,N_15518,N_14820);
xnor U17348 (N_17348,N_15512,N_15881);
nor U17349 (N_17349,N_14946,N_15734);
nand U17350 (N_17350,N_14931,N_15393);
nand U17351 (N_17351,N_14208,N_15165);
xnor U17352 (N_17352,N_15635,N_15231);
or U17353 (N_17353,N_15323,N_15831);
nand U17354 (N_17354,N_14915,N_14808);
xor U17355 (N_17355,N_15024,N_14260);
xnor U17356 (N_17356,N_14879,N_15714);
or U17357 (N_17357,N_15912,N_14210);
xor U17358 (N_17358,N_14919,N_14548);
and U17359 (N_17359,N_15457,N_15433);
xor U17360 (N_17360,N_14947,N_15789);
or U17361 (N_17361,N_15198,N_15652);
and U17362 (N_17362,N_15826,N_15362);
xnor U17363 (N_17363,N_15120,N_14634);
xnor U17364 (N_17364,N_15356,N_15958);
xnor U17365 (N_17365,N_15329,N_14273);
or U17366 (N_17366,N_15288,N_15980);
and U17367 (N_17367,N_14665,N_14988);
or U17368 (N_17368,N_14624,N_14103);
or U17369 (N_17369,N_15877,N_14146);
and U17370 (N_17370,N_15375,N_14199);
nor U17371 (N_17371,N_14204,N_14905);
or U17372 (N_17372,N_14923,N_15670);
or U17373 (N_17373,N_15745,N_14032);
xnor U17374 (N_17374,N_15498,N_15968);
xnor U17375 (N_17375,N_15107,N_14547);
or U17376 (N_17376,N_15272,N_15238);
or U17377 (N_17377,N_14523,N_14019);
nand U17378 (N_17378,N_15298,N_14997);
xnor U17379 (N_17379,N_14186,N_14299);
and U17380 (N_17380,N_15064,N_14722);
xor U17381 (N_17381,N_14515,N_15899);
or U17382 (N_17382,N_14543,N_15240);
or U17383 (N_17383,N_15134,N_15009);
and U17384 (N_17384,N_15752,N_15933);
nand U17385 (N_17385,N_15043,N_15919);
nand U17386 (N_17386,N_15057,N_14944);
xor U17387 (N_17387,N_15564,N_15306);
xnor U17388 (N_17388,N_14037,N_15739);
nor U17389 (N_17389,N_14556,N_14451);
or U17390 (N_17390,N_14805,N_15702);
nor U17391 (N_17391,N_14801,N_15881);
and U17392 (N_17392,N_15677,N_14906);
or U17393 (N_17393,N_14603,N_14464);
xnor U17394 (N_17394,N_14073,N_14835);
and U17395 (N_17395,N_14765,N_15944);
or U17396 (N_17396,N_14817,N_14067);
or U17397 (N_17397,N_14041,N_14031);
and U17398 (N_17398,N_15175,N_14186);
and U17399 (N_17399,N_15119,N_14331);
nor U17400 (N_17400,N_14901,N_15252);
and U17401 (N_17401,N_14397,N_14156);
nand U17402 (N_17402,N_15278,N_14268);
xor U17403 (N_17403,N_15505,N_15884);
nor U17404 (N_17404,N_15658,N_15442);
nand U17405 (N_17405,N_15358,N_14417);
and U17406 (N_17406,N_14920,N_14179);
xor U17407 (N_17407,N_15725,N_15457);
xor U17408 (N_17408,N_15158,N_14066);
and U17409 (N_17409,N_15718,N_15063);
nor U17410 (N_17410,N_15031,N_15576);
nor U17411 (N_17411,N_14046,N_15563);
xor U17412 (N_17412,N_15469,N_15940);
nand U17413 (N_17413,N_15821,N_14608);
xor U17414 (N_17414,N_14908,N_15622);
nand U17415 (N_17415,N_14683,N_14977);
nand U17416 (N_17416,N_14095,N_14645);
and U17417 (N_17417,N_14795,N_14367);
xnor U17418 (N_17418,N_14355,N_15238);
and U17419 (N_17419,N_15428,N_14851);
or U17420 (N_17420,N_14236,N_15189);
xnor U17421 (N_17421,N_15505,N_14681);
and U17422 (N_17422,N_15182,N_15769);
and U17423 (N_17423,N_14157,N_15343);
nor U17424 (N_17424,N_14341,N_15831);
or U17425 (N_17425,N_15364,N_15485);
xor U17426 (N_17426,N_15492,N_14117);
nand U17427 (N_17427,N_14426,N_14641);
nand U17428 (N_17428,N_15941,N_15188);
nor U17429 (N_17429,N_14251,N_15244);
nand U17430 (N_17430,N_14654,N_15891);
nor U17431 (N_17431,N_14181,N_15216);
nor U17432 (N_17432,N_14227,N_15994);
and U17433 (N_17433,N_14169,N_14732);
nand U17434 (N_17434,N_14684,N_15695);
nand U17435 (N_17435,N_15510,N_14236);
nand U17436 (N_17436,N_14605,N_14187);
or U17437 (N_17437,N_15025,N_15666);
nand U17438 (N_17438,N_15126,N_14253);
nor U17439 (N_17439,N_14558,N_15015);
nor U17440 (N_17440,N_14438,N_15907);
xnor U17441 (N_17441,N_15778,N_14669);
or U17442 (N_17442,N_14639,N_15892);
nand U17443 (N_17443,N_14423,N_15100);
nand U17444 (N_17444,N_15116,N_14777);
nor U17445 (N_17445,N_14546,N_15059);
or U17446 (N_17446,N_14188,N_14005);
or U17447 (N_17447,N_15977,N_15518);
and U17448 (N_17448,N_15214,N_14520);
nor U17449 (N_17449,N_15896,N_15564);
and U17450 (N_17450,N_15831,N_15406);
nand U17451 (N_17451,N_15307,N_15836);
nor U17452 (N_17452,N_14009,N_15309);
nand U17453 (N_17453,N_14496,N_14823);
nand U17454 (N_17454,N_15529,N_14543);
and U17455 (N_17455,N_14844,N_14081);
and U17456 (N_17456,N_15930,N_14226);
nand U17457 (N_17457,N_15902,N_14402);
xnor U17458 (N_17458,N_14028,N_14925);
nand U17459 (N_17459,N_15817,N_14635);
nand U17460 (N_17460,N_14539,N_14844);
nand U17461 (N_17461,N_14858,N_15956);
nor U17462 (N_17462,N_14166,N_15318);
or U17463 (N_17463,N_14478,N_14411);
xnor U17464 (N_17464,N_14630,N_14406);
and U17465 (N_17465,N_15027,N_14385);
nand U17466 (N_17466,N_14155,N_14343);
nor U17467 (N_17467,N_14686,N_15069);
xnor U17468 (N_17468,N_14500,N_15820);
and U17469 (N_17469,N_14383,N_14729);
nor U17470 (N_17470,N_14500,N_14566);
nand U17471 (N_17471,N_14360,N_15563);
or U17472 (N_17472,N_15233,N_14886);
xnor U17473 (N_17473,N_14436,N_15671);
xor U17474 (N_17474,N_15118,N_14986);
xnor U17475 (N_17475,N_15127,N_14850);
xor U17476 (N_17476,N_15915,N_15347);
xor U17477 (N_17477,N_14963,N_15713);
and U17478 (N_17478,N_14448,N_15980);
or U17479 (N_17479,N_15990,N_15989);
xnor U17480 (N_17480,N_15884,N_14239);
or U17481 (N_17481,N_14505,N_14599);
nand U17482 (N_17482,N_15469,N_15150);
nand U17483 (N_17483,N_14320,N_14112);
or U17484 (N_17484,N_14325,N_14591);
nand U17485 (N_17485,N_15723,N_14994);
nand U17486 (N_17486,N_15094,N_14191);
xor U17487 (N_17487,N_15550,N_15377);
xnor U17488 (N_17488,N_15926,N_15582);
xor U17489 (N_17489,N_14879,N_14386);
nand U17490 (N_17490,N_15030,N_14447);
or U17491 (N_17491,N_15638,N_14321);
nor U17492 (N_17492,N_14946,N_14514);
and U17493 (N_17493,N_15817,N_15956);
xor U17494 (N_17494,N_14716,N_15567);
xor U17495 (N_17495,N_14305,N_15124);
or U17496 (N_17496,N_14420,N_15020);
xnor U17497 (N_17497,N_15769,N_14574);
and U17498 (N_17498,N_15684,N_15095);
and U17499 (N_17499,N_14958,N_15284);
nand U17500 (N_17500,N_15927,N_15141);
nand U17501 (N_17501,N_15803,N_14251);
xor U17502 (N_17502,N_14705,N_14894);
and U17503 (N_17503,N_15264,N_14011);
nor U17504 (N_17504,N_14674,N_15742);
xor U17505 (N_17505,N_14523,N_14608);
or U17506 (N_17506,N_15920,N_15253);
xor U17507 (N_17507,N_15645,N_14393);
and U17508 (N_17508,N_14125,N_15177);
xor U17509 (N_17509,N_14655,N_14739);
nand U17510 (N_17510,N_14226,N_14136);
and U17511 (N_17511,N_14865,N_14220);
nor U17512 (N_17512,N_14291,N_15250);
nor U17513 (N_17513,N_15551,N_14190);
xor U17514 (N_17514,N_15901,N_15600);
xnor U17515 (N_17515,N_14183,N_15525);
and U17516 (N_17516,N_14672,N_14174);
nor U17517 (N_17517,N_15074,N_14331);
or U17518 (N_17518,N_14973,N_15774);
or U17519 (N_17519,N_15318,N_14188);
xor U17520 (N_17520,N_14838,N_14033);
and U17521 (N_17521,N_15233,N_15699);
nand U17522 (N_17522,N_15204,N_15537);
xor U17523 (N_17523,N_15343,N_14814);
xnor U17524 (N_17524,N_15421,N_15116);
xnor U17525 (N_17525,N_14962,N_14879);
xor U17526 (N_17526,N_14175,N_14904);
xor U17527 (N_17527,N_15180,N_15085);
or U17528 (N_17528,N_15292,N_15820);
xnor U17529 (N_17529,N_15957,N_15621);
and U17530 (N_17530,N_15875,N_15590);
nor U17531 (N_17531,N_15253,N_14910);
nor U17532 (N_17532,N_15605,N_14570);
or U17533 (N_17533,N_15486,N_14848);
or U17534 (N_17534,N_14023,N_14077);
xnor U17535 (N_17535,N_15481,N_15443);
xnor U17536 (N_17536,N_14872,N_14828);
or U17537 (N_17537,N_15237,N_15433);
xor U17538 (N_17538,N_15008,N_15907);
and U17539 (N_17539,N_15100,N_14955);
nand U17540 (N_17540,N_15248,N_15848);
or U17541 (N_17541,N_15698,N_15177);
xor U17542 (N_17542,N_15681,N_15397);
nand U17543 (N_17543,N_14651,N_14874);
and U17544 (N_17544,N_14594,N_15596);
nor U17545 (N_17545,N_14618,N_14287);
xor U17546 (N_17546,N_14381,N_14139);
and U17547 (N_17547,N_15262,N_14806);
nor U17548 (N_17548,N_14422,N_14266);
nand U17549 (N_17549,N_14748,N_14620);
or U17550 (N_17550,N_15272,N_14619);
nand U17551 (N_17551,N_14807,N_15218);
and U17552 (N_17552,N_14226,N_15318);
nor U17553 (N_17553,N_14861,N_14206);
nor U17554 (N_17554,N_15408,N_15812);
nor U17555 (N_17555,N_14827,N_15828);
xor U17556 (N_17556,N_15145,N_14427);
nand U17557 (N_17557,N_15499,N_14267);
xor U17558 (N_17558,N_15666,N_15813);
nor U17559 (N_17559,N_15175,N_15089);
nand U17560 (N_17560,N_14295,N_15972);
or U17561 (N_17561,N_14125,N_14703);
and U17562 (N_17562,N_14971,N_14170);
or U17563 (N_17563,N_15757,N_15925);
and U17564 (N_17564,N_14020,N_14854);
and U17565 (N_17565,N_14363,N_15760);
and U17566 (N_17566,N_15906,N_15241);
xnor U17567 (N_17567,N_15404,N_15576);
or U17568 (N_17568,N_14283,N_14955);
nand U17569 (N_17569,N_15732,N_15928);
xor U17570 (N_17570,N_14770,N_15231);
nor U17571 (N_17571,N_14165,N_14941);
xor U17572 (N_17572,N_14055,N_15109);
or U17573 (N_17573,N_15819,N_15602);
or U17574 (N_17574,N_14488,N_15717);
nor U17575 (N_17575,N_15957,N_14665);
xor U17576 (N_17576,N_14043,N_15415);
nand U17577 (N_17577,N_15780,N_14253);
nand U17578 (N_17578,N_14483,N_15288);
nor U17579 (N_17579,N_15937,N_15195);
nand U17580 (N_17580,N_15941,N_14245);
or U17581 (N_17581,N_15501,N_15300);
or U17582 (N_17582,N_15564,N_14211);
or U17583 (N_17583,N_14392,N_14275);
nor U17584 (N_17584,N_14913,N_14977);
nor U17585 (N_17585,N_14309,N_15863);
nor U17586 (N_17586,N_15293,N_14885);
nor U17587 (N_17587,N_15722,N_14394);
or U17588 (N_17588,N_15299,N_14630);
xor U17589 (N_17589,N_14037,N_15805);
or U17590 (N_17590,N_15497,N_15791);
or U17591 (N_17591,N_15430,N_15211);
or U17592 (N_17592,N_14009,N_14970);
and U17593 (N_17593,N_15072,N_14942);
nor U17594 (N_17594,N_15690,N_15598);
or U17595 (N_17595,N_15606,N_15032);
and U17596 (N_17596,N_15053,N_15884);
xnor U17597 (N_17597,N_15275,N_15899);
nor U17598 (N_17598,N_14707,N_14496);
nand U17599 (N_17599,N_14994,N_15290);
nor U17600 (N_17600,N_14544,N_15737);
nand U17601 (N_17601,N_15179,N_15229);
and U17602 (N_17602,N_15248,N_15546);
nor U17603 (N_17603,N_15003,N_15291);
nor U17604 (N_17604,N_15109,N_14122);
and U17605 (N_17605,N_15418,N_14657);
xor U17606 (N_17606,N_14453,N_15059);
and U17607 (N_17607,N_14860,N_15603);
and U17608 (N_17608,N_15706,N_14800);
xor U17609 (N_17609,N_15674,N_14305);
xnor U17610 (N_17610,N_15865,N_15809);
nor U17611 (N_17611,N_14890,N_14326);
and U17612 (N_17612,N_15156,N_15741);
or U17613 (N_17613,N_15600,N_15956);
nor U17614 (N_17614,N_14348,N_14800);
nor U17615 (N_17615,N_14025,N_15101);
nor U17616 (N_17616,N_14094,N_14535);
or U17617 (N_17617,N_14193,N_15332);
xor U17618 (N_17618,N_15617,N_15167);
nor U17619 (N_17619,N_14023,N_14881);
xnor U17620 (N_17620,N_14910,N_15768);
and U17621 (N_17621,N_14055,N_15587);
xnor U17622 (N_17622,N_15231,N_14719);
nand U17623 (N_17623,N_15845,N_14011);
nor U17624 (N_17624,N_15975,N_15938);
or U17625 (N_17625,N_14127,N_15779);
nor U17626 (N_17626,N_15431,N_14615);
and U17627 (N_17627,N_15778,N_14275);
xor U17628 (N_17628,N_15928,N_14514);
nor U17629 (N_17629,N_15596,N_14264);
nand U17630 (N_17630,N_15699,N_14596);
and U17631 (N_17631,N_15133,N_15902);
and U17632 (N_17632,N_15970,N_14284);
or U17633 (N_17633,N_14601,N_14195);
and U17634 (N_17634,N_14093,N_14721);
nor U17635 (N_17635,N_14102,N_14931);
nor U17636 (N_17636,N_15879,N_14159);
and U17637 (N_17637,N_14155,N_15240);
and U17638 (N_17638,N_15463,N_14582);
or U17639 (N_17639,N_15948,N_15004);
nand U17640 (N_17640,N_14367,N_14136);
nand U17641 (N_17641,N_15273,N_14233);
xor U17642 (N_17642,N_14896,N_14083);
xor U17643 (N_17643,N_14645,N_14968);
nand U17644 (N_17644,N_15240,N_15997);
nand U17645 (N_17645,N_14502,N_14665);
nand U17646 (N_17646,N_15365,N_14926);
nand U17647 (N_17647,N_15666,N_14002);
and U17648 (N_17648,N_14383,N_14844);
xnor U17649 (N_17649,N_15912,N_15183);
or U17650 (N_17650,N_14753,N_15229);
and U17651 (N_17651,N_14343,N_15745);
nand U17652 (N_17652,N_14387,N_15090);
nand U17653 (N_17653,N_15806,N_15022);
and U17654 (N_17654,N_14687,N_15347);
nand U17655 (N_17655,N_15187,N_14272);
nor U17656 (N_17656,N_15224,N_15759);
and U17657 (N_17657,N_14558,N_15966);
nand U17658 (N_17658,N_15584,N_14150);
xnor U17659 (N_17659,N_14666,N_14001);
nand U17660 (N_17660,N_15739,N_14820);
xor U17661 (N_17661,N_15660,N_15386);
nand U17662 (N_17662,N_14138,N_15404);
and U17663 (N_17663,N_15278,N_15607);
or U17664 (N_17664,N_15290,N_14769);
nand U17665 (N_17665,N_15440,N_15184);
xor U17666 (N_17666,N_14433,N_15908);
nand U17667 (N_17667,N_15217,N_15232);
xor U17668 (N_17668,N_14860,N_15857);
nand U17669 (N_17669,N_15434,N_14468);
nand U17670 (N_17670,N_14836,N_14178);
and U17671 (N_17671,N_14195,N_15768);
nand U17672 (N_17672,N_14497,N_15892);
xor U17673 (N_17673,N_15213,N_14868);
nor U17674 (N_17674,N_14720,N_14004);
nor U17675 (N_17675,N_14652,N_15966);
nor U17676 (N_17676,N_15512,N_14524);
nand U17677 (N_17677,N_14130,N_14139);
and U17678 (N_17678,N_15684,N_15903);
or U17679 (N_17679,N_14272,N_14601);
nor U17680 (N_17680,N_15579,N_15620);
or U17681 (N_17681,N_14950,N_15632);
and U17682 (N_17682,N_15749,N_15032);
xor U17683 (N_17683,N_15308,N_14310);
and U17684 (N_17684,N_14334,N_15902);
or U17685 (N_17685,N_15738,N_15741);
nor U17686 (N_17686,N_14947,N_14355);
nand U17687 (N_17687,N_15881,N_15612);
nand U17688 (N_17688,N_14523,N_14815);
xor U17689 (N_17689,N_15784,N_15797);
nand U17690 (N_17690,N_14507,N_14528);
and U17691 (N_17691,N_15453,N_15652);
or U17692 (N_17692,N_14944,N_14295);
and U17693 (N_17693,N_14591,N_14989);
nand U17694 (N_17694,N_14358,N_14958);
or U17695 (N_17695,N_15830,N_15993);
or U17696 (N_17696,N_14083,N_14074);
xnor U17697 (N_17697,N_14256,N_14113);
nand U17698 (N_17698,N_15769,N_15321);
xor U17699 (N_17699,N_15191,N_15111);
xor U17700 (N_17700,N_14757,N_15285);
and U17701 (N_17701,N_14393,N_15012);
xor U17702 (N_17702,N_15948,N_15957);
nand U17703 (N_17703,N_15573,N_14868);
or U17704 (N_17704,N_15081,N_14074);
or U17705 (N_17705,N_15842,N_15082);
xor U17706 (N_17706,N_14763,N_15077);
nor U17707 (N_17707,N_15171,N_15347);
nand U17708 (N_17708,N_14297,N_15066);
or U17709 (N_17709,N_14332,N_14690);
xor U17710 (N_17710,N_14167,N_15759);
nor U17711 (N_17711,N_14648,N_15791);
nor U17712 (N_17712,N_15100,N_14997);
nor U17713 (N_17713,N_15488,N_14213);
nand U17714 (N_17714,N_15617,N_15691);
nand U17715 (N_17715,N_15421,N_14882);
nand U17716 (N_17716,N_15465,N_14612);
and U17717 (N_17717,N_15286,N_15226);
nand U17718 (N_17718,N_15909,N_15119);
or U17719 (N_17719,N_15354,N_14844);
and U17720 (N_17720,N_15716,N_14401);
or U17721 (N_17721,N_14408,N_15481);
xnor U17722 (N_17722,N_14913,N_14745);
nor U17723 (N_17723,N_15086,N_14571);
xnor U17724 (N_17724,N_14592,N_15259);
or U17725 (N_17725,N_15510,N_15194);
nor U17726 (N_17726,N_15283,N_14048);
xnor U17727 (N_17727,N_15049,N_15993);
xnor U17728 (N_17728,N_14799,N_14412);
or U17729 (N_17729,N_14327,N_15554);
nor U17730 (N_17730,N_15798,N_15443);
and U17731 (N_17731,N_14239,N_14738);
nand U17732 (N_17732,N_15377,N_14401);
and U17733 (N_17733,N_14391,N_14628);
or U17734 (N_17734,N_15782,N_15456);
or U17735 (N_17735,N_15338,N_15133);
and U17736 (N_17736,N_15617,N_15104);
and U17737 (N_17737,N_15000,N_15219);
nand U17738 (N_17738,N_14313,N_14409);
nand U17739 (N_17739,N_15947,N_15840);
and U17740 (N_17740,N_15002,N_14119);
and U17741 (N_17741,N_15302,N_15208);
and U17742 (N_17742,N_14210,N_14334);
nand U17743 (N_17743,N_15472,N_15926);
and U17744 (N_17744,N_14295,N_15969);
nor U17745 (N_17745,N_15479,N_14104);
xnor U17746 (N_17746,N_15691,N_14571);
xnor U17747 (N_17747,N_15278,N_14433);
nand U17748 (N_17748,N_14188,N_14426);
xor U17749 (N_17749,N_14197,N_15547);
and U17750 (N_17750,N_14059,N_14082);
nand U17751 (N_17751,N_14353,N_15672);
nor U17752 (N_17752,N_14479,N_14934);
or U17753 (N_17753,N_14212,N_15246);
and U17754 (N_17754,N_15014,N_14346);
nor U17755 (N_17755,N_14134,N_15635);
and U17756 (N_17756,N_14223,N_15703);
or U17757 (N_17757,N_15478,N_14891);
or U17758 (N_17758,N_15009,N_14298);
nand U17759 (N_17759,N_14980,N_14141);
or U17760 (N_17760,N_14198,N_14422);
and U17761 (N_17761,N_14154,N_15427);
nor U17762 (N_17762,N_14128,N_15099);
nand U17763 (N_17763,N_15201,N_15801);
xor U17764 (N_17764,N_14562,N_14199);
and U17765 (N_17765,N_15396,N_15530);
or U17766 (N_17766,N_15304,N_15862);
xnor U17767 (N_17767,N_14117,N_14138);
nor U17768 (N_17768,N_14877,N_15282);
nand U17769 (N_17769,N_14893,N_15561);
or U17770 (N_17770,N_14920,N_15451);
xor U17771 (N_17771,N_15739,N_15939);
or U17772 (N_17772,N_15035,N_14786);
nand U17773 (N_17773,N_14595,N_15145);
nor U17774 (N_17774,N_15931,N_15164);
xor U17775 (N_17775,N_14821,N_15125);
and U17776 (N_17776,N_15117,N_14453);
and U17777 (N_17777,N_14262,N_14121);
or U17778 (N_17778,N_14454,N_15599);
nor U17779 (N_17779,N_15559,N_14595);
nand U17780 (N_17780,N_15038,N_15866);
or U17781 (N_17781,N_15715,N_15424);
xor U17782 (N_17782,N_15151,N_15524);
or U17783 (N_17783,N_14029,N_14257);
xnor U17784 (N_17784,N_15693,N_15382);
nor U17785 (N_17785,N_15568,N_15209);
or U17786 (N_17786,N_14801,N_15589);
or U17787 (N_17787,N_14143,N_14285);
xor U17788 (N_17788,N_14910,N_15001);
and U17789 (N_17789,N_14053,N_14181);
or U17790 (N_17790,N_15770,N_14256);
xnor U17791 (N_17791,N_15415,N_14329);
or U17792 (N_17792,N_14375,N_15976);
and U17793 (N_17793,N_15914,N_14581);
and U17794 (N_17794,N_15182,N_15423);
nand U17795 (N_17795,N_15185,N_15462);
xnor U17796 (N_17796,N_14334,N_14972);
and U17797 (N_17797,N_15175,N_14890);
or U17798 (N_17798,N_15963,N_15355);
nor U17799 (N_17799,N_14083,N_15598);
xor U17800 (N_17800,N_15701,N_14692);
xor U17801 (N_17801,N_15196,N_15698);
or U17802 (N_17802,N_14051,N_14299);
and U17803 (N_17803,N_14731,N_15165);
nor U17804 (N_17804,N_14604,N_15940);
or U17805 (N_17805,N_15170,N_14772);
and U17806 (N_17806,N_14189,N_14795);
or U17807 (N_17807,N_14143,N_15906);
nand U17808 (N_17808,N_15245,N_14652);
nor U17809 (N_17809,N_15753,N_14845);
nand U17810 (N_17810,N_15449,N_14484);
xnor U17811 (N_17811,N_15599,N_14733);
xnor U17812 (N_17812,N_14507,N_15565);
nor U17813 (N_17813,N_14664,N_14693);
or U17814 (N_17814,N_14879,N_14198);
or U17815 (N_17815,N_15011,N_15119);
or U17816 (N_17816,N_14394,N_14349);
nor U17817 (N_17817,N_15528,N_15457);
and U17818 (N_17818,N_14794,N_14021);
xnor U17819 (N_17819,N_14507,N_14056);
nor U17820 (N_17820,N_15097,N_15937);
xor U17821 (N_17821,N_14549,N_14157);
xnor U17822 (N_17822,N_15183,N_15954);
xor U17823 (N_17823,N_14237,N_15661);
nor U17824 (N_17824,N_14042,N_14931);
nor U17825 (N_17825,N_14856,N_15860);
or U17826 (N_17826,N_15390,N_14274);
and U17827 (N_17827,N_15178,N_15285);
nand U17828 (N_17828,N_14441,N_15133);
xor U17829 (N_17829,N_14336,N_15933);
and U17830 (N_17830,N_14529,N_14825);
nand U17831 (N_17831,N_14013,N_14960);
and U17832 (N_17832,N_14844,N_14419);
or U17833 (N_17833,N_15008,N_15440);
and U17834 (N_17834,N_14501,N_15328);
and U17835 (N_17835,N_15854,N_14342);
or U17836 (N_17836,N_14095,N_15300);
nor U17837 (N_17837,N_15656,N_15239);
nand U17838 (N_17838,N_14283,N_15155);
and U17839 (N_17839,N_14394,N_14150);
xor U17840 (N_17840,N_14225,N_14810);
nor U17841 (N_17841,N_15456,N_14268);
and U17842 (N_17842,N_15111,N_14089);
or U17843 (N_17843,N_15452,N_15268);
nor U17844 (N_17844,N_15927,N_14938);
and U17845 (N_17845,N_14918,N_15197);
xnor U17846 (N_17846,N_15057,N_15620);
or U17847 (N_17847,N_15040,N_15166);
nor U17848 (N_17848,N_15414,N_15688);
nor U17849 (N_17849,N_14206,N_14176);
or U17850 (N_17850,N_15510,N_15437);
or U17851 (N_17851,N_15719,N_15051);
or U17852 (N_17852,N_14316,N_15090);
or U17853 (N_17853,N_14792,N_14622);
nor U17854 (N_17854,N_15085,N_15498);
and U17855 (N_17855,N_14460,N_15025);
nand U17856 (N_17856,N_15320,N_15214);
xor U17857 (N_17857,N_14583,N_14128);
xor U17858 (N_17858,N_14965,N_14087);
nand U17859 (N_17859,N_14459,N_14421);
xnor U17860 (N_17860,N_15522,N_15188);
and U17861 (N_17861,N_15707,N_14504);
nand U17862 (N_17862,N_14557,N_14843);
or U17863 (N_17863,N_15009,N_15264);
and U17864 (N_17864,N_15103,N_15261);
nand U17865 (N_17865,N_15520,N_14104);
or U17866 (N_17866,N_14818,N_15576);
or U17867 (N_17867,N_15305,N_15960);
or U17868 (N_17868,N_14999,N_14728);
and U17869 (N_17869,N_14661,N_14808);
and U17870 (N_17870,N_15949,N_15638);
nand U17871 (N_17871,N_14616,N_14014);
or U17872 (N_17872,N_14325,N_15570);
or U17873 (N_17873,N_14187,N_15802);
nor U17874 (N_17874,N_14957,N_14596);
or U17875 (N_17875,N_15365,N_15205);
xor U17876 (N_17876,N_14719,N_15932);
and U17877 (N_17877,N_14019,N_15108);
or U17878 (N_17878,N_14475,N_15924);
and U17879 (N_17879,N_14337,N_14642);
nor U17880 (N_17880,N_15813,N_15930);
or U17881 (N_17881,N_14088,N_15641);
nand U17882 (N_17882,N_14607,N_14686);
nand U17883 (N_17883,N_14688,N_15407);
xor U17884 (N_17884,N_15257,N_14734);
and U17885 (N_17885,N_14696,N_14153);
or U17886 (N_17886,N_15623,N_15073);
and U17887 (N_17887,N_14412,N_14990);
xnor U17888 (N_17888,N_14388,N_14635);
or U17889 (N_17889,N_15809,N_14556);
xor U17890 (N_17890,N_14601,N_14433);
and U17891 (N_17891,N_15811,N_15336);
xnor U17892 (N_17892,N_14915,N_15054);
or U17893 (N_17893,N_15711,N_15037);
nand U17894 (N_17894,N_14659,N_14373);
or U17895 (N_17895,N_14748,N_15830);
or U17896 (N_17896,N_14227,N_14254);
nor U17897 (N_17897,N_14765,N_14080);
nand U17898 (N_17898,N_15673,N_15436);
or U17899 (N_17899,N_14260,N_14107);
or U17900 (N_17900,N_15459,N_15234);
and U17901 (N_17901,N_14011,N_15966);
nand U17902 (N_17902,N_14594,N_15646);
nand U17903 (N_17903,N_14416,N_14758);
and U17904 (N_17904,N_15550,N_14542);
nor U17905 (N_17905,N_14067,N_14110);
nand U17906 (N_17906,N_15232,N_14760);
nand U17907 (N_17907,N_15017,N_15669);
nand U17908 (N_17908,N_14664,N_15274);
nor U17909 (N_17909,N_15550,N_14865);
xnor U17910 (N_17910,N_14032,N_14073);
xor U17911 (N_17911,N_15598,N_15766);
nor U17912 (N_17912,N_15570,N_15985);
nor U17913 (N_17913,N_15314,N_15921);
and U17914 (N_17914,N_15252,N_15702);
or U17915 (N_17915,N_14949,N_14489);
or U17916 (N_17916,N_15712,N_15887);
or U17917 (N_17917,N_14588,N_14310);
xor U17918 (N_17918,N_15766,N_15643);
or U17919 (N_17919,N_14831,N_15713);
and U17920 (N_17920,N_14160,N_15282);
nand U17921 (N_17921,N_14545,N_14643);
nor U17922 (N_17922,N_14365,N_14538);
or U17923 (N_17923,N_15733,N_15378);
and U17924 (N_17924,N_14180,N_14446);
xor U17925 (N_17925,N_14056,N_15416);
or U17926 (N_17926,N_15994,N_15073);
xnor U17927 (N_17927,N_14693,N_15216);
or U17928 (N_17928,N_14129,N_14582);
xnor U17929 (N_17929,N_14990,N_14138);
nand U17930 (N_17930,N_14711,N_14746);
xor U17931 (N_17931,N_14455,N_14908);
or U17932 (N_17932,N_15098,N_14909);
nor U17933 (N_17933,N_14084,N_14382);
xnor U17934 (N_17934,N_15134,N_15242);
and U17935 (N_17935,N_14954,N_14500);
nand U17936 (N_17936,N_15065,N_14780);
and U17937 (N_17937,N_15483,N_15400);
nand U17938 (N_17938,N_14180,N_15119);
nor U17939 (N_17939,N_15050,N_15211);
nor U17940 (N_17940,N_14376,N_15853);
nand U17941 (N_17941,N_15369,N_15307);
and U17942 (N_17942,N_15823,N_14314);
and U17943 (N_17943,N_14024,N_15817);
nand U17944 (N_17944,N_15049,N_15155);
and U17945 (N_17945,N_14075,N_15154);
and U17946 (N_17946,N_14300,N_14674);
or U17947 (N_17947,N_15119,N_15816);
and U17948 (N_17948,N_14428,N_15815);
nand U17949 (N_17949,N_14400,N_14643);
and U17950 (N_17950,N_15411,N_14389);
nand U17951 (N_17951,N_14357,N_14916);
nand U17952 (N_17952,N_14564,N_15281);
xnor U17953 (N_17953,N_14676,N_14971);
or U17954 (N_17954,N_14549,N_15549);
xnor U17955 (N_17955,N_14510,N_14178);
or U17956 (N_17956,N_15523,N_15267);
xor U17957 (N_17957,N_14718,N_15201);
nor U17958 (N_17958,N_14152,N_15596);
nor U17959 (N_17959,N_14392,N_15739);
xor U17960 (N_17960,N_15957,N_14028);
nor U17961 (N_17961,N_15837,N_15529);
or U17962 (N_17962,N_15494,N_15943);
nor U17963 (N_17963,N_15064,N_15948);
xor U17964 (N_17964,N_15045,N_14780);
nor U17965 (N_17965,N_15219,N_15446);
xor U17966 (N_17966,N_15149,N_14243);
and U17967 (N_17967,N_14556,N_15583);
xor U17968 (N_17968,N_15581,N_14953);
nand U17969 (N_17969,N_14679,N_15428);
or U17970 (N_17970,N_14442,N_15489);
nand U17971 (N_17971,N_15362,N_14970);
nor U17972 (N_17972,N_14524,N_14581);
nand U17973 (N_17973,N_14995,N_14906);
or U17974 (N_17974,N_15427,N_15886);
nor U17975 (N_17975,N_15677,N_15150);
or U17976 (N_17976,N_15570,N_15215);
and U17977 (N_17977,N_15325,N_15684);
nor U17978 (N_17978,N_15685,N_14395);
xor U17979 (N_17979,N_15024,N_14682);
and U17980 (N_17980,N_15849,N_15416);
xor U17981 (N_17981,N_14424,N_15528);
and U17982 (N_17982,N_15106,N_14241);
xor U17983 (N_17983,N_15530,N_15704);
xnor U17984 (N_17984,N_15888,N_15716);
xor U17985 (N_17985,N_14399,N_14039);
and U17986 (N_17986,N_15308,N_15864);
and U17987 (N_17987,N_15416,N_15498);
or U17988 (N_17988,N_14844,N_15049);
and U17989 (N_17989,N_14801,N_15062);
and U17990 (N_17990,N_14756,N_15232);
xor U17991 (N_17991,N_15666,N_14098);
or U17992 (N_17992,N_15653,N_14659);
nor U17993 (N_17993,N_15935,N_14488);
nor U17994 (N_17994,N_15547,N_14468);
xor U17995 (N_17995,N_15000,N_15212);
nand U17996 (N_17996,N_14227,N_14089);
nor U17997 (N_17997,N_14265,N_14387);
nand U17998 (N_17998,N_15938,N_15829);
or U17999 (N_17999,N_14701,N_14026);
nand U18000 (N_18000,N_17769,N_17593);
nand U18001 (N_18001,N_16209,N_16765);
or U18002 (N_18002,N_17151,N_16293);
nand U18003 (N_18003,N_16240,N_16020);
xor U18004 (N_18004,N_17740,N_17558);
nand U18005 (N_18005,N_16983,N_17312);
and U18006 (N_18006,N_17709,N_16460);
nand U18007 (N_18007,N_16528,N_17132);
xor U18008 (N_18008,N_16651,N_17400);
and U18009 (N_18009,N_16034,N_16173);
or U18010 (N_18010,N_17973,N_16878);
xor U18011 (N_18011,N_16971,N_16849);
or U18012 (N_18012,N_16814,N_17056);
or U18013 (N_18013,N_17430,N_16812);
and U18014 (N_18014,N_16492,N_17502);
xnor U18015 (N_18015,N_17107,N_16762);
nand U18016 (N_18016,N_17032,N_16349);
or U18017 (N_18017,N_16868,N_16246);
xor U18018 (N_18018,N_16415,N_17747);
nand U18019 (N_18019,N_17313,N_16106);
nor U18020 (N_18020,N_17315,N_17358);
and U18021 (N_18021,N_16411,N_16070);
or U18022 (N_18022,N_17858,N_17300);
nand U18023 (N_18023,N_16655,N_16316);
and U18024 (N_18024,N_17433,N_16829);
nor U18025 (N_18025,N_17701,N_17317);
nor U18026 (N_18026,N_17326,N_16869);
nor U18027 (N_18027,N_17954,N_17061);
nand U18028 (N_18028,N_17960,N_17970);
nand U18029 (N_18029,N_16413,N_16015);
xor U18030 (N_18030,N_16940,N_17240);
xnor U18031 (N_18031,N_17807,N_16251);
nand U18032 (N_18032,N_17945,N_17085);
nand U18033 (N_18033,N_16152,N_16953);
and U18034 (N_18034,N_16132,N_17283);
or U18035 (N_18035,N_17704,N_17310);
xor U18036 (N_18036,N_17956,N_17087);
or U18037 (N_18037,N_16027,N_17270);
nor U18038 (N_18038,N_16252,N_16111);
xor U18039 (N_18039,N_17182,N_17346);
or U18040 (N_18040,N_16479,N_17254);
and U18041 (N_18041,N_17154,N_16846);
and U18042 (N_18042,N_17103,N_16258);
nand U18043 (N_18043,N_16447,N_17206);
and U18044 (N_18044,N_17454,N_16353);
xor U18045 (N_18045,N_16158,N_17802);
nor U18046 (N_18046,N_17291,N_16683);
xnor U18047 (N_18047,N_16540,N_16225);
and U18048 (N_18048,N_17349,N_16203);
nor U18049 (N_18049,N_16457,N_17452);
nand U18050 (N_18050,N_16643,N_16134);
nand U18051 (N_18051,N_16295,N_17962);
and U18052 (N_18052,N_16872,N_16742);
and U18053 (N_18053,N_17810,N_17278);
and U18054 (N_18054,N_17217,N_17916);
or U18055 (N_18055,N_17840,N_17763);
nand U18056 (N_18056,N_16238,N_16630);
xnor U18057 (N_18057,N_16587,N_16636);
and U18058 (N_18058,N_17906,N_16698);
nand U18059 (N_18059,N_16109,N_17640);
and U18060 (N_18060,N_17901,N_16304);
nor U18061 (N_18061,N_17548,N_16740);
xor U18062 (N_18062,N_16004,N_17546);
nor U18063 (N_18063,N_16929,N_17775);
xnor U18064 (N_18064,N_16049,N_16091);
and U18065 (N_18065,N_17047,N_16767);
nor U18066 (N_18066,N_16571,N_16220);
xnor U18067 (N_18067,N_17095,N_17233);
or U18068 (N_18068,N_17086,N_16391);
or U18069 (N_18069,N_17332,N_17281);
and U18070 (N_18070,N_17881,N_17213);
xor U18071 (N_18071,N_16852,N_16544);
and U18072 (N_18072,N_16987,N_17849);
xnor U18073 (N_18073,N_17365,N_17311);
xnor U18074 (N_18074,N_16312,N_17439);
nand U18075 (N_18075,N_17808,N_17109);
or U18076 (N_18076,N_17083,N_17955);
nor U18077 (N_18077,N_16489,N_17417);
nand U18078 (N_18078,N_16164,N_17145);
nor U18079 (N_18079,N_17444,N_16517);
or U18080 (N_18080,N_17832,N_17553);
or U18081 (N_18081,N_17965,N_16486);
and U18082 (N_18082,N_16065,N_17494);
nand U18083 (N_18083,N_16261,N_16429);
or U18084 (N_18084,N_16546,N_17185);
and U18085 (N_18085,N_16501,N_17745);
nor U18086 (N_18086,N_16634,N_17748);
nor U18087 (N_18087,N_16563,N_16666);
nand U18088 (N_18088,N_17938,N_16461);
and U18089 (N_18089,N_16355,N_17484);
or U18090 (N_18090,N_17512,N_16827);
or U18091 (N_18091,N_17885,N_17790);
nor U18092 (N_18092,N_17379,N_17408);
or U18093 (N_18093,N_16318,N_16838);
nand U18094 (N_18094,N_17668,N_16837);
and U18095 (N_18095,N_16184,N_16670);
xor U18096 (N_18096,N_16508,N_16815);
nand U18097 (N_18097,N_17884,N_16017);
or U18098 (N_18098,N_17538,N_16752);
nor U18099 (N_18099,N_16310,N_17157);
xnor U18100 (N_18100,N_16061,N_17784);
nand U18101 (N_18101,N_17680,N_17274);
or U18102 (N_18102,N_16386,N_17943);
and U18103 (N_18103,N_17455,N_16340);
or U18104 (N_18104,N_16130,N_16319);
xor U18105 (N_18105,N_17035,N_17142);
or U18106 (N_18106,N_17895,N_16692);
nand U18107 (N_18107,N_17038,N_17075);
and U18108 (N_18108,N_16482,N_16298);
xor U18109 (N_18109,N_16821,N_17564);
and U18110 (N_18110,N_16466,N_17435);
and U18111 (N_18111,N_17860,N_16262);
and U18112 (N_18112,N_16373,N_16645);
nor U18113 (N_18113,N_16906,N_17952);
or U18114 (N_18114,N_17357,N_17575);
or U18115 (N_18115,N_16914,N_16671);
or U18116 (N_18116,N_17331,N_17819);
nor U18117 (N_18117,N_17366,N_16367);
or U18118 (N_18118,N_17856,N_17042);
or U18119 (N_18119,N_17027,N_16504);
xnor U18120 (N_18120,N_17999,N_16970);
nand U18121 (N_18121,N_16717,N_17496);
nor U18122 (N_18122,N_17987,N_16577);
or U18123 (N_18123,N_17200,N_17603);
and U18124 (N_18124,N_16819,N_17779);
or U18125 (N_18125,N_17486,N_17480);
or U18126 (N_18126,N_16343,N_16487);
nor U18127 (N_18127,N_17043,N_17355);
and U18128 (N_18128,N_16652,N_16522);
or U18129 (N_18129,N_16268,N_17762);
and U18130 (N_18130,N_17731,N_16398);
nand U18131 (N_18131,N_17950,N_17879);
and U18132 (N_18132,N_16001,N_16053);
nor U18133 (N_18133,N_16082,N_17186);
nand U18134 (N_18134,N_17729,N_16775);
nor U18135 (N_18135,N_16456,N_17631);
nand U18136 (N_18136,N_17215,N_16011);
and U18137 (N_18137,N_16993,N_17628);
nand U18138 (N_18138,N_16480,N_17882);
nand U18139 (N_18139,N_16472,N_17065);
nand U18140 (N_18140,N_17110,N_17339);
or U18141 (N_18141,N_17941,N_16513);
nand U18142 (N_18142,N_16916,N_16188);
and U18143 (N_18143,N_17117,N_17532);
or U18144 (N_18144,N_17738,N_17985);
and U18145 (N_18145,N_16875,N_16595);
or U18146 (N_18146,N_16687,N_17048);
xnor U18147 (N_18147,N_16650,N_17114);
or U18148 (N_18148,N_17483,N_16449);
nand U18149 (N_18149,N_17535,N_17523);
xnor U18150 (N_18150,N_16798,N_16206);
nor U18151 (N_18151,N_16503,N_16321);
and U18152 (N_18152,N_17464,N_17932);
and U18153 (N_18153,N_16073,N_16968);
nor U18154 (N_18154,N_16845,N_16085);
nor U18155 (N_18155,N_17539,N_17910);
or U18156 (N_18156,N_17124,N_16677);
xor U18157 (N_18157,N_17175,N_17244);
xor U18158 (N_18158,N_17000,N_17652);
and U18159 (N_18159,N_16409,N_16243);
nor U18160 (N_18160,N_17833,N_17012);
nor U18161 (N_18161,N_16700,N_16949);
nand U18162 (N_18162,N_17282,N_17466);
or U18163 (N_18163,N_17696,N_16756);
or U18164 (N_18164,N_17793,N_16191);
xnor U18165 (N_18165,N_17727,N_16214);
nand U18166 (N_18166,N_17074,N_17163);
nand U18167 (N_18167,N_17221,N_17304);
or U18168 (N_18168,N_16621,N_16344);
nand U18169 (N_18169,N_17398,N_17842);
xor U18170 (N_18170,N_17055,N_16640);
nor U18171 (N_18171,N_16789,N_17517);
and U18172 (N_18172,N_17482,N_16858);
nand U18173 (N_18173,N_16986,N_17610);
nor U18174 (N_18174,N_17015,N_17041);
xor U18175 (N_18175,N_17479,N_16769);
xor U18176 (N_18176,N_16974,N_16753);
xor U18177 (N_18177,N_17578,N_16359);
nand U18178 (N_18178,N_16143,N_17555);
or U18179 (N_18179,N_16614,N_17685);
nor U18180 (N_18180,N_16946,N_16113);
nor U18181 (N_18181,N_17150,N_17927);
and U18182 (N_18182,N_17638,N_16939);
and U18183 (N_18183,N_17725,N_17514);
and U18184 (N_18184,N_17227,N_16681);
xor U18185 (N_18185,N_17285,N_16913);
nor U18186 (N_18186,N_16750,N_16573);
or U18187 (N_18187,N_17886,N_17020);
nor U18188 (N_18188,N_17905,N_16785);
or U18189 (N_18189,N_17399,N_16684);
nor U18190 (N_18190,N_16463,N_17759);
xor U18191 (N_18191,N_17996,N_16952);
nor U18192 (N_18192,N_16446,N_16881);
nor U18193 (N_18193,N_16657,N_17294);
nor U18194 (N_18194,N_17926,N_17506);
and U18195 (N_18195,N_17783,N_16376);
nand U18196 (N_18196,N_17995,N_16779);
nand U18197 (N_18197,N_16305,N_17036);
nor U18198 (N_18198,N_17823,N_17198);
nand U18199 (N_18199,N_17653,N_17648);
xnor U18200 (N_18200,N_16580,N_16495);
nor U18201 (N_18201,N_16945,N_17467);
or U18202 (N_18202,N_17016,N_17633);
or U18203 (N_18203,N_17649,N_17991);
nor U18204 (N_18204,N_17112,N_17238);
nand U18205 (N_18205,N_16820,N_17395);
or U18206 (N_18206,N_17247,N_17156);
nor U18207 (N_18207,N_16934,N_16232);
nor U18208 (N_18208,N_17859,N_17976);
and U18209 (N_18209,N_17711,N_17513);
nand U18210 (N_18210,N_17409,N_17104);
and U18211 (N_18211,N_16112,N_17717);
and U18212 (N_18212,N_16836,N_17873);
and U18213 (N_18213,N_16537,N_17462);
and U18214 (N_18214,N_16094,N_17742);
nand U18215 (N_18215,N_17176,N_16688);
nand U18216 (N_18216,N_16417,N_16598);
or U18217 (N_18217,N_17908,N_17722);
nor U18218 (N_18218,N_16271,N_17583);
xor U18219 (N_18219,N_16464,N_16117);
nand U18220 (N_18220,N_16257,N_17251);
and U18221 (N_18221,N_16024,N_16961);
and U18222 (N_18222,N_17586,N_17557);
and U18223 (N_18223,N_17948,N_17867);
nor U18224 (N_18224,N_17090,N_17367);
or U18225 (N_18225,N_16506,N_17624);
and U18226 (N_18226,N_16626,N_17091);
nor U18227 (N_18227,N_17348,N_16327);
nor U18228 (N_18228,N_16610,N_17571);
or U18229 (N_18229,N_16227,N_16121);
nand U18230 (N_18230,N_17297,N_16424);
or U18231 (N_18231,N_16330,N_17771);
and U18232 (N_18232,N_17734,N_16625);
or U18233 (N_18233,N_16631,N_17359);
nor U18234 (N_18234,N_16364,N_16059);
nor U18235 (N_18235,N_17937,N_16994);
and U18236 (N_18236,N_17381,N_16891);
xor U18237 (N_18237,N_16808,N_16382);
and U18238 (N_18238,N_17724,N_16083);
or U18239 (N_18239,N_17096,N_17647);
xnor U18240 (N_18240,N_16129,N_17118);
nor U18241 (N_18241,N_16897,N_17449);
or U18242 (N_18242,N_16995,N_17865);
nor U18243 (N_18243,N_16156,N_17519);
or U18244 (N_18244,N_17997,N_16822);
xnor U18245 (N_18245,N_16910,N_16629);
nor U18246 (N_18246,N_16241,N_17106);
and U18247 (N_18247,N_17286,N_16354);
and U18248 (N_18248,N_17301,N_16427);
xor U18249 (N_18249,N_17947,N_16680);
and U18250 (N_18250,N_16476,N_17766);
xnor U18251 (N_18251,N_16541,N_17004);
nand U18252 (N_18252,N_16202,N_17595);
and U18253 (N_18253,N_17529,N_16281);
nor U18254 (N_18254,N_17299,N_17170);
xnor U18255 (N_18255,N_16781,N_17716);
or U18256 (N_18256,N_16028,N_16611);
and U18257 (N_18257,N_16925,N_17672);
xnor U18258 (N_18258,N_16992,N_17029);
nor U18259 (N_18259,N_16661,N_16695);
xnor U18260 (N_18260,N_17219,N_17728);
nor U18261 (N_18261,N_16467,N_17058);
or U18262 (N_18262,N_16641,N_16407);
and U18263 (N_18263,N_17656,N_17380);
or U18264 (N_18264,N_17429,N_17826);
xnor U18265 (N_18265,N_17388,N_16718);
nand U18266 (N_18266,N_17998,N_16600);
and U18267 (N_18267,N_16317,N_17582);
xor U18268 (N_18268,N_17646,N_17234);
nand U18269 (N_18269,N_17561,N_17149);
or U18270 (N_18270,N_17961,N_16632);
nor U18271 (N_18271,N_16419,N_17340);
nand U18272 (N_18272,N_17542,N_17116);
nand U18273 (N_18273,N_17168,N_17940);
or U18274 (N_18274,N_16441,N_17034);
or U18275 (N_18275,N_16628,N_17463);
nor U18276 (N_18276,N_17620,N_17302);
nor U18277 (N_18277,N_17416,N_16100);
xnor U18278 (N_18278,N_17053,N_16060);
nand U18279 (N_18279,N_16899,N_17959);
or U18280 (N_18280,N_16048,N_16301);
nand U18281 (N_18281,N_16704,N_17448);
or U18282 (N_18282,N_17585,N_16880);
or U18283 (N_18283,N_16841,N_16624);
nor U18284 (N_18284,N_16040,N_16644);
and U18285 (N_18285,N_16342,N_16269);
xor U18286 (N_18286,N_16991,N_16051);
xor U18287 (N_18287,N_17597,N_17713);
or U18288 (N_18288,N_17756,N_17081);
nand U18289 (N_18289,N_16850,N_16887);
and U18290 (N_18290,N_16337,N_17174);
or U18291 (N_18291,N_17147,N_16057);
or U18292 (N_18292,N_17017,N_17625);
nand U18293 (N_18293,N_17739,N_17663);
xnor U18294 (N_18294,N_17703,N_17815);
nand U18295 (N_18295,N_16603,N_17022);
or U18296 (N_18296,N_17014,N_16984);
xnor U18297 (N_18297,N_17457,N_17050);
or U18298 (N_18298,N_16564,N_16674);
or U18299 (N_18299,N_17394,N_17402);
and U18300 (N_18300,N_16155,N_16575);
or U18301 (N_18301,N_16380,N_17266);
and U18302 (N_18302,N_16216,N_17600);
nand U18303 (N_18303,N_17655,N_17073);
or U18304 (N_18304,N_17052,N_16557);
nand U18305 (N_18305,N_16902,N_16729);
and U18306 (N_18306,N_17627,N_17708);
or U18307 (N_18307,N_16263,N_16790);
nor U18308 (N_18308,N_16551,N_17851);
or U18309 (N_18309,N_16591,N_16041);
xnor U18310 (N_18310,N_16175,N_17431);
nand U18311 (N_18311,N_16068,N_16390);
nor U18312 (N_18312,N_17465,N_16672);
nand U18313 (N_18313,N_16230,N_16348);
nand U18314 (N_18314,N_17426,N_16646);
or U18315 (N_18315,N_17994,N_16569);
xnor U18316 (N_18316,N_16087,N_16219);
nor U18317 (N_18317,N_16357,N_17801);
xnor U18318 (N_18318,N_16590,N_16727);
xor U18319 (N_18319,N_17131,N_17942);
and U18320 (N_18320,N_17273,N_17666);
nand U18321 (N_18321,N_17963,N_17953);
nand U18322 (N_18322,N_16116,N_16010);
or U18323 (N_18323,N_17077,N_17172);
and U18324 (N_18324,N_16706,N_17897);
and U18325 (N_18325,N_17816,N_17899);
nand U18326 (N_18326,N_17706,N_17307);
nor U18327 (N_18327,N_16667,N_17127);
xor U18328 (N_18328,N_17877,N_17841);
or U18329 (N_18329,N_17692,N_17391);
nor U18330 (N_18330,N_16282,N_16222);
or U18331 (N_18331,N_16699,N_16458);
nor U18332 (N_18332,N_17249,N_17797);
or U18333 (N_18333,N_16208,N_17084);
nand U18334 (N_18334,N_16254,N_17552);
nor U18335 (N_18335,N_16757,N_17813);
xnor U18336 (N_18336,N_17190,N_17441);
or U18337 (N_18337,N_17069,N_17662);
nor U18338 (N_18338,N_17836,N_17403);
and U18339 (N_18339,N_16181,N_17689);
xnor U18340 (N_18340,N_16938,N_16582);
or U18341 (N_18341,N_17305,N_17900);
xnor U18342 (N_18342,N_17437,N_17609);
or U18343 (N_18343,N_17556,N_16859);
and U18344 (N_18344,N_17907,N_17814);
nor U18345 (N_18345,N_16481,N_16135);
xor U18346 (N_18346,N_17100,N_16000);
nand U18347 (N_18347,N_16515,N_16066);
or U18348 (N_18348,N_16224,N_17796);
or U18349 (N_18349,N_16721,N_17258);
xor U18350 (N_18350,N_17468,N_16077);
nor U18351 (N_18351,N_17914,N_17601);
nand U18352 (N_18352,N_16558,N_17968);
xor U18353 (N_18353,N_17673,N_16793);
or U18354 (N_18354,N_17225,N_17622);
nor U18355 (N_18355,N_16832,N_16568);
or U18356 (N_18356,N_16867,N_17824);
nor U18357 (N_18357,N_16138,N_16888);
nor U18358 (N_18358,N_17159,N_17453);
xor U18359 (N_18359,N_16924,N_16749);
xor U18360 (N_18360,N_16505,N_16654);
and U18361 (N_18361,N_16593,N_16153);
and U18362 (N_18362,N_16445,N_16406);
nand U18363 (N_18363,N_17726,N_17295);
xor U18364 (N_18364,N_16723,N_16776);
xor U18365 (N_18365,N_17382,N_16436);
nand U18366 (N_18366,N_17957,N_16098);
or U18367 (N_18367,N_17531,N_17990);
xor U18368 (N_18368,N_16314,N_17487);
and U18369 (N_18369,N_16308,N_16574);
xor U18370 (N_18370,N_16187,N_17707);
nand U18371 (N_18371,N_17592,N_16786);
and U18372 (N_18372,N_16719,N_16128);
or U18373 (N_18373,N_17188,N_17001);
nand U18374 (N_18374,N_16177,N_16217);
xor U18375 (N_18375,N_17515,N_16297);
nor U18376 (N_18376,N_17891,N_17637);
or U18377 (N_18377,N_17040,N_16176);
xor U18378 (N_18378,N_17030,N_17277);
and U18379 (N_18379,N_16773,N_16309);
xnor U18380 (N_18380,N_17356,N_16196);
or U18381 (N_18381,N_16890,N_16948);
nor U18382 (N_18382,N_17636,N_17966);
and U18383 (N_18383,N_17507,N_17559);
and U18384 (N_18384,N_17757,N_16870);
nand U18385 (N_18385,N_17913,N_16244);
xnor U18386 (N_18386,N_17572,N_16895);
nand U18387 (N_18387,N_17498,N_17864);
nand U18388 (N_18388,N_17862,N_17800);
or U18389 (N_18389,N_17290,N_17641);
nor U18390 (N_18390,N_17650,N_17544);
xnor U18391 (N_18391,N_16279,N_16403);
and U18392 (N_18392,N_17324,N_17013);
xor U18393 (N_18393,N_16266,N_17831);
nand U18394 (N_18394,N_16931,N_17695);
and U18395 (N_18395,N_16579,N_17063);
xor U18396 (N_18396,N_17099,N_17386);
nand U18397 (N_18397,N_16972,N_17364);
or U18398 (N_18398,N_16816,N_17264);
and U18399 (N_18399,N_17893,N_17259);
and U18400 (N_18400,N_16520,N_17353);
xnor U18401 (N_18401,N_17837,N_17102);
nor U18402 (N_18402,N_17613,N_17284);
and U18403 (N_18403,N_16122,N_16923);
nand U18404 (N_18404,N_17377,N_17410);
nand U18405 (N_18405,N_17687,N_16553);
xnor U18406 (N_18406,N_16896,N_17764);
xnor U18407 (N_18407,N_17418,N_16649);
xnor U18408 (N_18408,N_17780,N_16998);
xor U18409 (N_18409,N_17619,N_16425);
nand U18410 (N_18410,N_17896,N_16788);
and U18411 (N_18411,N_16124,N_17889);
nor U18412 (N_18412,N_16696,N_16810);
nor U18413 (N_18413,N_16079,N_16774);
or U18414 (N_18414,N_16578,N_17248);
and U18415 (N_18415,N_16207,N_16738);
and U18416 (N_18416,N_17009,N_16955);
nor U18417 (N_18417,N_17194,N_16985);
nand U18418 (N_18418,N_16025,N_16915);
xor U18419 (N_18419,N_17434,N_17329);
and U18420 (N_18420,N_17162,N_16855);
xnor U18421 (N_18421,N_17485,N_16944);
nand U18422 (N_18422,N_16512,N_17642);
or U18423 (N_18423,N_16694,N_16639);
xor U18424 (N_18424,N_17303,N_16860);
nor U18425 (N_18425,N_17499,N_16146);
nand U18426 (N_18426,N_17772,N_17697);
or U18427 (N_18427,N_16885,N_17588);
or U18428 (N_18428,N_16287,N_16019);
and U18429 (N_18429,N_16471,N_17773);
xor U18430 (N_18430,N_17360,N_16523);
and U18431 (N_18431,N_16642,N_16397);
xor U18432 (N_18432,N_17723,N_17334);
nand U18433 (N_18433,N_16623,N_17644);
nor U18434 (N_18434,N_17076,N_17580);
or U18435 (N_18435,N_17616,N_16063);
or U18436 (N_18436,N_17944,N_16302);
xor U18437 (N_18437,N_16333,N_17492);
xor U18438 (N_18438,N_17369,N_17072);
xnor U18439 (N_18439,N_16950,N_17830);
nor U18440 (N_18440,N_16157,N_16029);
nand U18441 (N_18441,N_17037,N_17984);
and U18442 (N_18442,N_17928,N_16123);
or U18443 (N_18443,N_17003,N_17843);
nor U18444 (N_18444,N_16315,N_16328);
xnor U18445 (N_18445,N_16249,N_17694);
and U18446 (N_18446,N_17501,N_17497);
and U18447 (N_18447,N_16072,N_17678);
nor U18448 (N_18448,N_16708,N_17256);
xnor U18449 (N_18449,N_17443,N_17912);
nor U18450 (N_18450,N_16235,N_16772);
and U18451 (N_18451,N_17378,N_16534);
and U18452 (N_18452,N_16421,N_17911);
nor U18453 (N_18453,N_16958,N_17456);
xnor U18454 (N_18454,N_16703,N_16784);
nor U18455 (N_18455,N_16543,N_16478);
xor U18456 (N_18456,N_16084,N_16180);
xnor U18457 (N_18457,N_17195,N_16882);
and U18458 (N_18458,N_16306,N_17550);
nor U18459 (N_18459,N_16440,N_16830);
and U18460 (N_18460,N_17385,N_16093);
nor U18461 (N_18461,N_17809,N_17146);
xor U18462 (N_18462,N_17051,N_16922);
xor U18463 (N_18463,N_16294,N_16521);
or U18464 (N_18464,N_17972,N_17275);
xnor U18465 (N_18465,N_17537,N_16245);
and U18466 (N_18466,N_16336,N_17338);
xor U18467 (N_18467,N_16737,N_17587);
and U18468 (N_18468,N_16973,N_16178);
nor U18469 (N_18469,N_17812,N_16889);
nand U18470 (N_18470,N_17089,N_16597);
xnor U18471 (N_18471,N_16452,N_16159);
and U18472 (N_18472,N_17308,N_17574);
and U18473 (N_18473,N_16285,N_16483);
xnor U18474 (N_18474,N_16678,N_17345);
or U18475 (N_18475,N_17733,N_16036);
xnor U18476 (N_18476,N_16911,N_17591);
nand U18477 (N_18477,N_17148,N_16559);
or U18478 (N_18478,N_16067,N_16834);
nand U18479 (N_18479,N_16550,N_16307);
xor U18480 (N_18480,N_17321,N_17397);
or U18481 (N_18481,N_16851,N_17664);
xnor U18482 (N_18482,N_17296,N_17064);
nand U18483 (N_18483,N_17472,N_17549);
or U18484 (N_18484,N_16444,N_16229);
or U18485 (N_18485,N_17969,N_17746);
nor U18486 (N_18486,N_16136,N_16030);
nor U18487 (N_18487,N_17445,N_16778);
nand U18488 (N_18488,N_16928,N_16137);
nor U18489 (N_18489,N_17921,N_16736);
xor U18490 (N_18490,N_16959,N_17805);
or U18491 (N_18491,N_16535,N_16783);
and U18492 (N_18492,N_16823,N_17596);
or U18493 (N_18493,N_17590,N_17082);
nor U18494 (N_18494,N_17180,N_16387);
nor U18495 (N_18495,N_17438,N_16105);
nor U18496 (N_18496,N_17028,N_16371);
nand U18497 (N_18497,N_17350,N_17774);
or U18498 (N_18498,N_17551,N_17732);
and U18499 (N_18499,N_16937,N_17705);
nor U18500 (N_18500,N_16525,N_17070);
nand U18501 (N_18501,N_17850,N_16871);
nand U18502 (N_18502,N_16284,N_17847);
nand U18503 (N_18503,N_17822,N_17128);
nand U18504 (N_18504,N_17423,N_17049);
or U18505 (N_18505,N_16760,N_17866);
or U18506 (N_18506,N_17846,N_17411);
nor U18507 (N_18507,N_16800,N_17208);
nand U18508 (N_18508,N_17872,N_16734);
and U18509 (N_18509,N_17436,N_17861);
xor U18510 (N_18510,N_16332,N_16863);
nand U18511 (N_18511,N_17917,N_16142);
xor U18512 (N_18512,N_16894,N_16864);
or U18513 (N_18513,N_16743,N_16023);
and U18514 (N_18514,N_16932,N_16277);
xor U18515 (N_18515,N_16556,N_16771);
or U18516 (N_18516,N_16195,N_16369);
nor U18517 (N_18517,N_16286,N_16154);
nor U18518 (N_18518,N_17239,N_16691);
nor U18519 (N_18519,N_16960,N_16296);
nor U18520 (N_18520,N_17853,N_17352);
nand U18521 (N_18521,N_17611,N_17491);
or U18522 (N_18522,N_17967,N_17735);
nor U18523 (N_18523,N_16172,N_17025);
nor U18524 (N_18524,N_17088,N_17024);
or U18525 (N_18525,N_17688,N_17223);
and U18526 (N_18526,N_17623,N_16747);
nor U18527 (N_18527,N_17280,N_17607);
nor U18528 (N_18528,N_17621,N_17269);
xor U18529 (N_18529,N_16375,N_16384);
nand U18530 (N_18530,N_17298,N_16239);
xor U18531 (N_18531,N_17754,N_17825);
nand U18532 (N_18532,N_17476,N_16780);
nand U18533 (N_18533,N_16542,N_16679);
and U18534 (N_18534,N_17533,N_17659);
or U18535 (N_18535,N_16715,N_16183);
nor U18536 (N_18536,N_16401,N_16050);
xnor U18537 (N_18537,N_16562,N_16530);
nor U18538 (N_18538,N_16378,N_16488);
and U18539 (N_18539,N_16274,N_17811);
nor U18540 (N_18540,N_17540,N_17715);
xnor U18541 (N_18541,N_17770,N_16739);
and U18542 (N_18542,N_16223,N_16607);
and U18543 (N_18543,N_16434,N_16638);
xor U18544 (N_18544,N_16033,N_16477);
or U18545 (N_18545,N_16388,N_17670);
nand U18546 (N_18546,N_17543,N_16081);
and U18547 (N_18547,N_16689,N_16400);
nor U18548 (N_18548,N_16954,N_16547);
nand U18549 (N_18549,N_16549,N_16334);
nand U18550 (N_18550,N_16576,N_17518);
nand U18551 (N_18551,N_17451,N_16161);
nor U18552 (N_18552,N_17478,N_16226);
and U18553 (N_18553,N_17421,N_16514);
nand U18554 (N_18554,N_16104,N_17325);
nand U18555 (N_18555,N_17894,N_16606);
nand U18556 (N_18556,N_17207,N_17165);
nand U18557 (N_18557,N_16978,N_17844);
or U18558 (N_18558,N_17677,N_17660);
nand U18559 (N_18559,N_16170,N_16876);
and U18560 (N_18560,N_16267,N_16656);
xnor U18561 (N_18561,N_17153,N_17752);
and U18562 (N_18562,N_17920,N_16601);
xnor U18563 (N_18563,N_16856,N_16189);
and U18564 (N_18564,N_17971,N_16843);
and U18565 (N_18565,N_16979,N_17854);
xor U18566 (N_18566,N_17257,N_16345);
nor U18567 (N_18567,N_16366,N_17720);
and U18568 (N_18568,N_16395,N_17584);
nor U18569 (N_18569,N_17224,N_17606);
xor U18570 (N_18570,N_16539,N_17977);
xnor U18571 (N_18571,N_17068,N_16532);
or U18572 (N_18572,N_17384,N_16705);
or U18573 (N_18573,N_17712,N_17835);
nor U18574 (N_18574,N_17934,N_17373);
and U18575 (N_18575,N_16311,N_16248);
xor U18576 (N_18576,N_17272,N_17263);
and U18577 (N_18577,N_17276,N_16168);
xor U18578 (N_18578,N_17612,N_17419);
or U18579 (N_18579,N_17133,N_16179);
and U18580 (N_18580,N_16554,N_16099);
nor U18581 (N_18581,N_16303,N_16748);
nor U18582 (N_18582,N_17045,N_17804);
and U18583 (N_18583,N_17675,N_16289);
xor U18584 (N_18584,N_16039,N_16724);
xnor U18585 (N_18585,N_16448,N_16107);
nor U18586 (N_18586,N_17261,N_17122);
xnor U18587 (N_18587,N_17632,N_16686);
or U18588 (N_18588,N_16389,N_16908);
nor U18589 (N_18589,N_16981,N_16255);
or U18590 (N_18590,N_17375,N_17615);
xnor U18591 (N_18591,N_17645,N_17245);
nand U18592 (N_18592,N_16115,N_16927);
nor U18593 (N_18593,N_16265,N_17570);
nand U18594 (N_18594,N_17191,N_16133);
xnor U18595 (N_18595,N_17372,N_17924);
nand U18596 (N_18596,N_17287,N_16561);
nand U18597 (N_18597,N_16365,N_16396);
nor U18598 (N_18598,N_17203,N_17460);
and U18599 (N_18599,N_16383,N_16325);
and U18600 (N_18600,N_17125,N_17021);
nand U18601 (N_18601,N_17892,N_17226);
or U18602 (N_18602,N_16794,N_16982);
xor U18603 (N_18603,N_16531,N_17078);
nor U18604 (N_18604,N_16874,N_16394);
or U18605 (N_18605,N_17199,N_16273);
nor U18606 (N_18606,N_16720,N_17293);
or U18607 (N_18607,N_17568,N_16347);
or U18608 (N_18608,N_17488,N_16393);
nand U18609 (N_18609,N_17608,N_17792);
or U18610 (N_18610,N_17936,N_17469);
and U18611 (N_18611,N_16171,N_16148);
xor U18612 (N_18612,N_16608,N_16907);
and U18613 (N_18613,N_17918,N_16791);
nand U18614 (N_18614,N_17605,N_17827);
nand U18615 (N_18615,N_16151,N_16075);
nor U18616 (N_18616,N_16526,N_16833);
and U18617 (N_18617,N_17173,N_17503);
nand U18618 (N_18618,N_16701,N_16941);
and U18619 (N_18619,N_16809,N_17749);
nand U18620 (N_18620,N_17141,N_16141);
and U18621 (N_18621,N_16493,N_16682);
or U18622 (N_18622,N_17563,N_16237);
xnor U18623 (N_18623,N_16451,N_17374);
xnor U18624 (N_18624,N_16035,N_17450);
and U18625 (N_18625,N_16119,N_17581);
xor U18626 (N_18626,N_16292,N_17166);
nor U18627 (N_18627,N_16898,N_16102);
or U18628 (N_18628,N_16565,N_17665);
and U18629 (N_18629,N_16647,N_17289);
xnor U18630 (N_18630,N_17602,N_16233);
xor U18631 (N_18631,N_17684,N_16474);
xor U18632 (N_18632,N_17031,N_17493);
nand U18633 (N_18633,N_17250,N_17393);
and U18634 (N_18634,N_17222,N_16731);
nor U18635 (N_18635,N_17989,N_16096);
or U18636 (N_18636,N_17789,N_16741);
nor U18637 (N_18637,N_16538,N_17002);
and U18638 (N_18638,N_16169,N_17576);
or U18639 (N_18639,N_17658,N_16439);
nand U18640 (N_18640,N_16746,N_17508);
nand U18641 (N_18641,N_17415,N_17923);
nor U18642 (N_18642,N_16975,N_17786);
xor U18643 (N_18643,N_16442,N_16926);
and U18644 (N_18644,N_17005,N_17661);
xnor U18645 (N_18645,N_17777,N_17904);
nor U18646 (N_18646,N_16796,N_16962);
or U18647 (N_18647,N_16270,N_17220);
and U18648 (N_18648,N_17820,N_16438);
or U18649 (N_18649,N_17054,N_16754);
and U18650 (N_18650,N_16420,N_16174);
xnor U18651 (N_18651,N_17767,N_17007);
and U18652 (N_18652,N_16967,N_17828);
nor U18653 (N_18653,N_17599,N_17237);
or U18654 (N_18654,N_16801,N_16455);
and U18655 (N_18655,N_16589,N_16186);
nand U18656 (N_18656,N_17516,N_16893);
nor U18657 (N_18657,N_16690,N_17903);
nor U18658 (N_18658,N_17679,N_17152);
xor U18659 (N_18659,N_17255,N_16988);
and U18660 (N_18660,N_16787,N_17951);
or U18661 (N_18661,N_17528,N_16283);
nor U18662 (N_18662,N_16062,N_17314);
or U18663 (N_18663,N_17376,N_17011);
or U18664 (N_18664,N_16402,N_16825);
or U18665 (N_18665,N_17511,N_16524);
and U18666 (N_18666,N_16942,N_17803);
and U18667 (N_18667,N_17818,N_17205);
nor U18668 (N_18668,N_16007,N_16323);
or U18669 (N_18669,N_16469,N_16470);
or U18670 (N_18670,N_16450,N_16519);
and U18671 (N_18671,N_16619,N_16454);
or U18672 (N_18672,N_16761,N_17231);
nand U18673 (N_18673,N_17993,N_16566);
xor U18674 (N_18674,N_17440,N_17530);
xor U18675 (N_18675,N_16702,N_17589);
nand U18676 (N_18676,N_17071,N_16996);
nor U18677 (N_18677,N_17554,N_17113);
xor U18678 (N_18678,N_17806,N_16410);
or U18679 (N_18679,N_16300,N_16709);
or U18680 (N_18680,N_17330,N_16074);
nand U18681 (N_18681,N_17626,N_17525);
or U18682 (N_18682,N_17874,N_16957);
and U18683 (N_18683,N_16044,N_16193);
nor U18684 (N_18684,N_16126,N_17594);
nand U18685 (N_18685,N_16166,N_17868);
and U18686 (N_18686,N_16584,N_17246);
nand U18687 (N_18687,N_17212,N_17446);
nand U18688 (N_18688,N_17420,N_17760);
xor U18689 (N_18689,N_16602,N_16160);
xor U18690 (N_18690,N_17545,N_16103);
nor U18691 (N_18691,N_16693,N_17171);
nor U18692 (N_18692,N_16510,N_16211);
and U18693 (N_18693,N_16428,N_17839);
nand U18694 (N_18694,N_16498,N_16006);
and U18695 (N_18695,N_17560,N_16363);
nor U18696 (N_18696,N_16884,N_17915);
or U18697 (N_18697,N_17392,N_17730);
nor U18698 (N_18698,N_16379,N_16637);
nand U18699 (N_18699,N_16615,N_16089);
xor U18700 (N_18700,N_16758,N_16416);
and U18701 (N_18701,N_17428,N_16533);
or U18702 (N_18702,N_16086,N_16022);
xor U18703 (N_18703,N_17898,N_17541);
nand U18704 (N_18704,N_16165,N_16818);
nor U18705 (N_18705,N_16095,N_16604);
or U18706 (N_18706,N_17447,N_16056);
xor U18707 (N_18707,N_16215,N_16069);
and U18708 (N_18708,N_17974,N_17782);
nor U18709 (N_18709,N_17026,N_16966);
and U18710 (N_18710,N_16862,N_17138);
xnor U18711 (N_18711,N_16346,N_16432);
and U18712 (N_18712,N_17406,N_17521);
nand U18713 (N_18713,N_17111,N_16795);
or U18714 (N_18714,N_16609,N_16194);
xnor U18715 (N_18715,N_17279,N_16120);
or U18716 (N_18716,N_17676,N_17046);
nor U18717 (N_18717,N_16935,N_17700);
nand U18718 (N_18718,N_16873,N_16485);
nor U18719 (N_18719,N_17121,N_16290);
nand U18720 (N_18720,N_17922,N_16078);
and U18721 (N_18721,N_16370,N_16560);
nand U18722 (N_18722,N_17235,N_16732);
or U18723 (N_18723,N_17890,N_17674);
xnor U18724 (N_18724,N_16055,N_17201);
nand U18725 (N_18725,N_16583,N_17750);
xor U18726 (N_18726,N_16127,N_17265);
xnor U18727 (N_18727,N_17787,N_17320);
nor U18728 (N_18728,N_17736,N_17630);
or U18729 (N_18729,N_17108,N_16198);
nor U18730 (N_18730,N_16276,N_16620);
and U18731 (N_18731,N_16341,N_16299);
xor U18732 (N_18732,N_16879,N_16088);
or U18733 (N_18733,N_16496,N_17008);
nor U18734 (N_18734,N_16032,N_16351);
xor U18735 (N_18735,N_17988,N_17424);
or U18736 (N_18736,N_17396,N_17629);
and U18737 (N_18737,N_16231,N_17253);
nand U18738 (N_18738,N_17039,N_17719);
and U18739 (N_18739,N_17193,N_17425);
or U18740 (N_18740,N_16511,N_17821);
nand U18741 (N_18741,N_16861,N_16372);
xor U18742 (N_18742,N_17432,N_16014);
or U18743 (N_18743,N_17702,N_16759);
or U18744 (N_18744,N_17949,N_16016);
nand U18745 (N_18745,N_17838,N_17158);
or U18746 (N_18746,N_17370,N_16404);
and U18747 (N_18747,N_17669,N_16149);
and U18748 (N_18748,N_17115,N_17768);
xor U18749 (N_18749,N_17134,N_16866);
and U18750 (N_18750,N_16664,N_16280);
or U18751 (N_18751,N_17883,N_17407);
and U18752 (N_18752,N_17211,N_17389);
nand U18753 (N_18753,N_16900,N_16965);
nand U18754 (N_18754,N_16918,N_16331);
nand U18755 (N_18755,N_17094,N_16422);
nand U18756 (N_18756,N_16205,N_17368);
xnor U18757 (N_18757,N_17761,N_17504);
and U18758 (N_18758,N_16668,N_16536);
and U18759 (N_18759,N_17336,N_17169);
nor U18760 (N_18760,N_17845,N_16768);
and U18761 (N_18761,N_17136,N_17634);
or U18762 (N_18762,N_16356,N_16594);
nor U18763 (N_18763,N_16555,N_17681);
and U18764 (N_18764,N_16462,N_17755);
and U18765 (N_18765,N_16322,N_17505);
nand U18766 (N_18766,N_16484,N_16802);
and U18767 (N_18767,N_17243,N_16658);
or U18768 (N_18768,N_17569,N_17643);
and U18769 (N_18769,N_17577,N_16491);
and U18770 (N_18770,N_17562,N_17080);
xor U18771 (N_18771,N_16272,N_16012);
xor U18772 (N_18772,N_16045,N_17473);
nor U18773 (N_18773,N_17241,N_17232);
or U18774 (N_18774,N_16377,N_16805);
and U18775 (N_18775,N_17387,N_16473);
xor U18776 (N_18776,N_16635,N_16046);
xor U18777 (N_18777,N_17267,N_17510);
or U18778 (N_18778,N_17522,N_16831);
or U18779 (N_18779,N_16676,N_17319);
nand U18780 (N_18780,N_16904,N_17354);
nand U18781 (N_18781,N_17181,N_17933);
xnor U18782 (N_18782,N_17693,N_17405);
nor U18783 (N_18783,N_16835,N_17137);
xor U18784 (N_18784,N_16500,N_16817);
and U18785 (N_18785,N_16080,N_17229);
or U18786 (N_18786,N_17143,N_16977);
or U18787 (N_18787,N_16259,N_16147);
and U18788 (N_18788,N_16185,N_17980);
xor U18789 (N_18789,N_16844,N_16588);
nand U18790 (N_18790,N_17361,N_16826);
xor U18791 (N_18791,N_16509,N_17573);
nor U18792 (N_18792,N_17214,N_17598);
nand U18793 (N_18793,N_17383,N_16423);
and U18794 (N_18794,N_16182,N_17328);
nand U18795 (N_18795,N_17187,N_16313);
xnor U18796 (N_18796,N_16660,N_16162);
nor U18797 (N_18797,N_16745,N_17958);
and U18798 (N_18798,N_17067,N_16782);
or U18799 (N_18799,N_16013,N_17686);
and U18800 (N_18800,N_16204,N_16435);
xor U18801 (N_18801,N_16097,N_16430);
and U18802 (N_18802,N_16291,N_17526);
xor U18803 (N_18803,N_16824,N_16163);
or U18804 (N_18804,N_17781,N_17909);
xor U18805 (N_18805,N_16919,N_16199);
xor U18806 (N_18806,N_17288,N_16009);
nand U18807 (N_18807,N_17351,N_16437);
and U18808 (N_18808,N_17018,N_17744);
nand U18809 (N_18809,N_16627,N_17875);
and U18810 (N_18810,N_17347,N_17902);
or U18811 (N_18811,N_16200,N_17778);
nor U18812 (N_18812,N_16005,N_17262);
or U18813 (N_18813,N_17023,N_16131);
nand U18814 (N_18814,N_16201,N_17177);
nor U18815 (N_18815,N_16071,N_16076);
or U18816 (N_18816,N_16622,N_17093);
xnor U18817 (N_18817,N_17737,N_16242);
or U18818 (N_18818,N_17414,N_17869);
and U18819 (N_18819,N_17461,N_16092);
or U18820 (N_18820,N_16797,N_17044);
nor U18821 (N_18821,N_17863,N_17292);
nand U18822 (N_18822,N_16125,N_16499);
nor U18823 (N_18823,N_17848,N_17919);
xor U18824 (N_18824,N_17946,N_17101);
nor U18825 (N_18825,N_17765,N_16433);
or U18826 (N_18826,N_17682,N_16418);
xnor U18827 (N_18827,N_17657,N_16465);
nand U18828 (N_18828,N_16228,N_16669);
and U18829 (N_18829,N_17341,N_16712);
xnor U18830 (N_18830,N_16529,N_16101);
or U18831 (N_18831,N_16920,N_16361);
xor U18832 (N_18832,N_16976,N_16570);
nor U18833 (N_18833,N_16350,N_16426);
nand U18834 (N_18834,N_17458,N_16711);
or U18835 (N_18835,N_16744,N_17471);
xnor U18836 (N_18836,N_17033,N_17228);
or U18837 (N_18837,N_16933,N_17059);
or U18838 (N_18838,N_17092,N_16917);
xnor U18839 (N_18839,N_16807,N_16502);
nor U18840 (N_18840,N_16804,N_17975);
xnor U18841 (N_18841,N_17322,N_17362);
or U18842 (N_18842,N_17667,N_17097);
and U18843 (N_18843,N_16997,N_16548);
xnor U18844 (N_18844,N_17495,N_17791);
or U18845 (N_18845,N_17390,N_16763);
nand U18846 (N_18846,N_16234,N_16043);
or U18847 (N_18847,N_17753,N_17189);
nand U18848 (N_18848,N_17260,N_16250);
xor U18849 (N_18849,N_16192,N_16618);
or U18850 (N_18850,N_16999,N_16275);
and U18851 (N_18851,N_17006,N_17139);
or U18852 (N_18852,N_17160,N_16653);
or U18853 (N_18853,N_17105,N_17401);
nand U18854 (N_18854,N_16443,N_17857);
nor U18855 (N_18855,N_16770,N_17534);
nand U18856 (N_18856,N_16339,N_16494);
nor U18857 (N_18857,N_16329,N_17930);
nand U18858 (N_18858,N_16507,N_17155);
nand U18859 (N_18859,N_16042,N_17714);
nor U18860 (N_18860,N_17161,N_17935);
or U18861 (N_18861,N_16828,N_16490);
nand U18862 (N_18862,N_16324,N_16633);
and U18863 (N_18863,N_16140,N_17524);
xnor U18864 (N_18864,N_16399,N_17566);
nor U18865 (N_18865,N_16930,N_16468);
nand U18866 (N_18866,N_16190,N_16118);
and U18867 (N_18867,N_16839,N_16909);
xnor U18868 (N_18868,N_16545,N_16964);
or U18869 (N_18869,N_17565,N_16936);
xor U18870 (N_18870,N_16212,N_17710);
or U18871 (N_18871,N_17202,N_17144);
xnor U18872 (N_18872,N_17817,N_16054);
and U18873 (N_18873,N_17490,N_16854);
xnor U18874 (N_18874,N_17481,N_17547);
xnor U18875 (N_18875,N_16777,N_17887);
and U18876 (N_18876,N_16951,N_16728);
or U18877 (N_18877,N_16335,N_17690);
or U18878 (N_18878,N_16475,N_17343);
nand U18879 (N_18879,N_17527,N_16612);
and U18880 (N_18880,N_16392,N_16047);
or U18881 (N_18881,N_16381,N_17363);
xnor U18882 (N_18882,N_16352,N_16278);
xnor U18883 (N_18883,N_16755,N_16903);
nand U18884 (N_18884,N_16052,N_17651);
nor U18885 (N_18885,N_16613,N_17167);
xnor U18886 (N_18886,N_17878,N_17618);
xnor U18887 (N_18887,N_17888,N_17268);
and U18888 (N_18888,N_17344,N_16412);
nor U18889 (N_18889,N_17333,N_16368);
nand U18890 (N_18890,N_16596,N_16320);
nand U18891 (N_18891,N_16288,N_16853);
or U18892 (N_18892,N_16021,N_17057);
nand U18893 (N_18893,N_17119,N_16811);
and U18894 (N_18894,N_17271,N_16405);
and U18895 (N_18895,N_16673,N_17509);
or U18896 (N_18896,N_17776,N_17413);
nand U18897 (N_18897,N_17929,N_17880);
nor U18898 (N_18898,N_17019,N_17123);
and U18899 (N_18899,N_16764,N_17981);
xnor U18900 (N_18900,N_17316,N_16218);
xor U18901 (N_18901,N_16236,N_16497);
and U18902 (N_18902,N_17470,N_16799);
and U18903 (N_18903,N_16947,N_17743);
nand U18904 (N_18904,N_16663,N_16108);
and U18905 (N_18905,N_16031,N_17871);
and U18906 (N_18906,N_16358,N_16616);
nor U18907 (N_18907,N_17992,N_17979);
xnor U18908 (N_18908,N_16197,N_17925);
xor U18909 (N_18909,N_17852,N_17794);
xor U18910 (N_18910,N_16002,N_17683);
xnor U18911 (N_18911,N_17654,N_16710);
nand U18912 (N_18912,N_16726,N_16144);
nand U18913 (N_18913,N_17788,N_16886);
xor U18914 (N_18914,N_17060,N_17931);
nand U18915 (N_18915,N_17983,N_17335);
nand U18916 (N_18916,N_16665,N_16675);
or U18917 (N_18917,N_16139,N_17489);
xnor U18918 (N_18918,N_17130,N_16585);
nor U18919 (N_18919,N_17579,N_17062);
nand U18920 (N_18920,N_16883,N_16956);
nand U18921 (N_18921,N_17986,N_17252);
or U18922 (N_18922,N_17691,N_16362);
xor U18923 (N_18923,N_16892,N_16848);
or U18924 (N_18924,N_16685,N_17242);
xor U18925 (N_18925,N_16969,N_17829);
or U18926 (N_18926,N_16264,N_17459);
xnor U18927 (N_18927,N_16806,N_16714);
or U18928 (N_18928,N_17404,N_17834);
and U18929 (N_18929,N_16360,N_16221);
nand U18930 (N_18930,N_16980,N_17617);
and U18931 (N_18931,N_16008,N_16213);
xor U18932 (N_18932,N_16114,N_17500);
nor U18933 (N_18933,N_17318,N_16018);
xnor U18934 (N_18934,N_17140,N_17184);
nand U18935 (N_18935,N_17079,N_16453);
and U18936 (N_18936,N_16026,N_17120);
and U18937 (N_18937,N_17795,N_16989);
xnor U18938 (N_18938,N_17474,N_16408);
nand U18939 (N_18939,N_17758,N_16963);
and U18940 (N_18940,N_16326,N_17192);
or U18941 (N_18941,N_17183,N_16943);
or U18942 (N_18942,N_17422,N_16599);
nor U18943 (N_18943,N_16038,N_17671);
nor U18944 (N_18944,N_17520,N_17475);
nor U18945 (N_18945,N_16722,N_16210);
xor U18946 (N_18946,N_16766,N_17327);
or U18947 (N_18947,N_16581,N_17098);
or U18948 (N_18948,N_16090,N_16572);
nor U18949 (N_18949,N_17306,N_17939);
nor U18950 (N_18950,N_16842,N_16713);
nor U18951 (N_18951,N_16648,N_16840);
and U18952 (N_18952,N_17010,N_17799);
nand U18953 (N_18953,N_17741,N_16459);
nor U18954 (N_18954,N_17196,N_16385);
nand U18955 (N_18955,N_17197,N_17698);
or U18956 (N_18956,N_17218,N_16058);
and U18957 (N_18957,N_17614,N_16167);
xnor U18958 (N_18958,N_16921,N_16527);
or U18959 (N_18959,N_16518,N_17442);
xnor U18960 (N_18960,N_16150,N_16003);
or U18961 (N_18961,N_16659,N_17604);
and U18962 (N_18962,N_17323,N_17371);
nand U18963 (N_18963,N_16905,N_16256);
and U18964 (N_18964,N_16847,N_17309);
nand U18965 (N_18965,N_16592,N_16697);
nand U18966 (N_18966,N_16716,N_16586);
nor U18967 (N_18967,N_16110,N_17216);
nor U18968 (N_18968,N_16792,N_17870);
and U18969 (N_18969,N_16901,N_16552);
or U18970 (N_18970,N_17536,N_17164);
and U18971 (N_18971,N_17178,N_17721);
and U18972 (N_18972,N_16037,N_17427);
and U18973 (N_18973,N_17635,N_17982);
or U18974 (N_18974,N_16803,N_16064);
and U18975 (N_18975,N_16253,N_16735);
nor U18976 (N_18976,N_16877,N_16145);
nand U18977 (N_18977,N_16733,N_17785);
or U18978 (N_18978,N_17179,N_17230);
or U18979 (N_18979,N_17204,N_17129);
and U18980 (N_18980,N_17337,N_16865);
xnor U18981 (N_18981,N_17876,N_17236);
nand U18982 (N_18982,N_17964,N_17751);
nor U18983 (N_18983,N_17798,N_17477);
xnor U18984 (N_18984,N_16247,N_17412);
xnor U18985 (N_18985,N_16751,N_16260);
nor U18986 (N_18986,N_16813,N_16516);
xor U18987 (N_18987,N_17126,N_17209);
or U18988 (N_18988,N_16725,N_16567);
nor U18989 (N_18989,N_16857,N_16707);
or U18990 (N_18990,N_17135,N_17855);
and U18991 (N_18991,N_16414,N_17210);
xnor U18992 (N_18992,N_17567,N_17342);
and U18993 (N_18993,N_17699,N_16431);
xor U18994 (N_18994,N_16990,N_16338);
nor U18995 (N_18995,N_17639,N_16374);
nand U18996 (N_18996,N_16605,N_16662);
or U18997 (N_18997,N_17066,N_17718);
or U18998 (N_18998,N_16730,N_16912);
xor U18999 (N_18999,N_16617,N_17978);
nand U19000 (N_19000,N_17278,N_16650);
nand U19001 (N_19001,N_17381,N_16252);
nand U19002 (N_19002,N_17259,N_16074);
and U19003 (N_19003,N_16554,N_17289);
nor U19004 (N_19004,N_17443,N_17849);
xnor U19005 (N_19005,N_17853,N_17384);
or U19006 (N_19006,N_17428,N_16510);
xnor U19007 (N_19007,N_17678,N_16183);
or U19008 (N_19008,N_16421,N_16487);
nand U19009 (N_19009,N_17454,N_17255);
nand U19010 (N_19010,N_17922,N_16640);
xor U19011 (N_19011,N_17968,N_17394);
and U19012 (N_19012,N_16509,N_16093);
nand U19013 (N_19013,N_17822,N_17224);
nor U19014 (N_19014,N_17363,N_16443);
and U19015 (N_19015,N_16874,N_17072);
and U19016 (N_19016,N_16813,N_16691);
and U19017 (N_19017,N_16756,N_16674);
xnor U19018 (N_19018,N_17358,N_17089);
xnor U19019 (N_19019,N_16744,N_17625);
and U19020 (N_19020,N_16760,N_17367);
and U19021 (N_19021,N_16938,N_16458);
nand U19022 (N_19022,N_16290,N_16753);
or U19023 (N_19023,N_16573,N_16906);
nor U19024 (N_19024,N_16945,N_16355);
or U19025 (N_19025,N_17041,N_17302);
and U19026 (N_19026,N_17136,N_16865);
and U19027 (N_19027,N_16217,N_17760);
nor U19028 (N_19028,N_17157,N_16562);
nand U19029 (N_19029,N_16068,N_17457);
xnor U19030 (N_19030,N_17511,N_16824);
nand U19031 (N_19031,N_16036,N_16810);
xnor U19032 (N_19032,N_16966,N_16325);
xor U19033 (N_19033,N_16719,N_17235);
nand U19034 (N_19034,N_16364,N_16155);
or U19035 (N_19035,N_16380,N_17923);
or U19036 (N_19036,N_17095,N_17332);
nor U19037 (N_19037,N_17514,N_17071);
xnor U19038 (N_19038,N_16094,N_17171);
xnor U19039 (N_19039,N_16626,N_16618);
or U19040 (N_19040,N_17509,N_16995);
nor U19041 (N_19041,N_17403,N_16642);
nand U19042 (N_19042,N_16454,N_17531);
nor U19043 (N_19043,N_17889,N_16861);
xnor U19044 (N_19044,N_17106,N_16745);
nand U19045 (N_19045,N_17747,N_17152);
and U19046 (N_19046,N_16393,N_17255);
and U19047 (N_19047,N_17544,N_17453);
nor U19048 (N_19048,N_16996,N_17654);
and U19049 (N_19049,N_16642,N_16080);
xnor U19050 (N_19050,N_16761,N_17950);
xnor U19051 (N_19051,N_16889,N_17774);
or U19052 (N_19052,N_17980,N_16741);
xnor U19053 (N_19053,N_17927,N_16557);
nand U19054 (N_19054,N_17189,N_16164);
xnor U19055 (N_19055,N_16592,N_16863);
xor U19056 (N_19056,N_16940,N_17044);
or U19057 (N_19057,N_16556,N_17300);
nor U19058 (N_19058,N_16887,N_17342);
nand U19059 (N_19059,N_16788,N_16604);
xor U19060 (N_19060,N_16475,N_16024);
nor U19061 (N_19061,N_16732,N_16804);
and U19062 (N_19062,N_17094,N_16583);
nor U19063 (N_19063,N_16868,N_16225);
and U19064 (N_19064,N_17358,N_16215);
or U19065 (N_19065,N_16594,N_16912);
or U19066 (N_19066,N_17694,N_17786);
or U19067 (N_19067,N_16033,N_16757);
and U19068 (N_19068,N_16788,N_16423);
nand U19069 (N_19069,N_17744,N_17926);
or U19070 (N_19070,N_16035,N_16588);
nand U19071 (N_19071,N_16073,N_16752);
xor U19072 (N_19072,N_17721,N_16802);
and U19073 (N_19073,N_17368,N_16319);
and U19074 (N_19074,N_16360,N_17030);
nand U19075 (N_19075,N_17728,N_17807);
or U19076 (N_19076,N_16701,N_17965);
nand U19077 (N_19077,N_16770,N_17770);
nor U19078 (N_19078,N_16898,N_17594);
and U19079 (N_19079,N_16111,N_16711);
nand U19080 (N_19080,N_16028,N_16625);
nand U19081 (N_19081,N_17869,N_17911);
or U19082 (N_19082,N_17124,N_16703);
and U19083 (N_19083,N_16358,N_16197);
or U19084 (N_19084,N_16472,N_16727);
nand U19085 (N_19085,N_16723,N_17301);
and U19086 (N_19086,N_17390,N_17506);
nor U19087 (N_19087,N_17750,N_16674);
nand U19088 (N_19088,N_16495,N_17909);
or U19089 (N_19089,N_16088,N_16316);
or U19090 (N_19090,N_16555,N_16338);
nor U19091 (N_19091,N_16724,N_16626);
xnor U19092 (N_19092,N_17815,N_17443);
xor U19093 (N_19093,N_16787,N_16929);
xnor U19094 (N_19094,N_16383,N_16801);
nand U19095 (N_19095,N_16360,N_16046);
nor U19096 (N_19096,N_16659,N_16557);
nor U19097 (N_19097,N_17161,N_16963);
and U19098 (N_19098,N_17940,N_17132);
nand U19099 (N_19099,N_16437,N_17593);
and U19100 (N_19100,N_16042,N_16764);
nor U19101 (N_19101,N_16116,N_16742);
nor U19102 (N_19102,N_17634,N_16425);
and U19103 (N_19103,N_17479,N_17977);
xor U19104 (N_19104,N_17806,N_17890);
nor U19105 (N_19105,N_16300,N_16261);
or U19106 (N_19106,N_16260,N_16428);
and U19107 (N_19107,N_17684,N_16556);
nand U19108 (N_19108,N_16236,N_17928);
or U19109 (N_19109,N_16165,N_16170);
nor U19110 (N_19110,N_17438,N_17596);
nor U19111 (N_19111,N_16611,N_16052);
and U19112 (N_19112,N_17900,N_16165);
nand U19113 (N_19113,N_16652,N_16482);
nand U19114 (N_19114,N_17862,N_16618);
nand U19115 (N_19115,N_17103,N_17224);
nor U19116 (N_19116,N_16424,N_17534);
xor U19117 (N_19117,N_16712,N_17835);
and U19118 (N_19118,N_16724,N_16716);
nand U19119 (N_19119,N_17111,N_16672);
nor U19120 (N_19120,N_16532,N_17438);
xnor U19121 (N_19121,N_17938,N_16180);
or U19122 (N_19122,N_17241,N_17692);
nor U19123 (N_19123,N_17787,N_16565);
or U19124 (N_19124,N_17503,N_17079);
or U19125 (N_19125,N_16700,N_17751);
nand U19126 (N_19126,N_17637,N_17178);
xnor U19127 (N_19127,N_16079,N_16173);
nand U19128 (N_19128,N_17023,N_16308);
and U19129 (N_19129,N_17166,N_17292);
or U19130 (N_19130,N_16989,N_16511);
and U19131 (N_19131,N_16473,N_17667);
nand U19132 (N_19132,N_16272,N_17594);
and U19133 (N_19133,N_17599,N_17721);
and U19134 (N_19134,N_16001,N_17493);
nand U19135 (N_19135,N_16313,N_17864);
nor U19136 (N_19136,N_17020,N_16113);
or U19137 (N_19137,N_16475,N_16091);
nor U19138 (N_19138,N_16944,N_17544);
xor U19139 (N_19139,N_16267,N_16498);
and U19140 (N_19140,N_17436,N_17251);
nand U19141 (N_19141,N_17328,N_16283);
nand U19142 (N_19142,N_16558,N_17647);
nor U19143 (N_19143,N_17977,N_17492);
and U19144 (N_19144,N_17422,N_17667);
xnor U19145 (N_19145,N_17286,N_17988);
and U19146 (N_19146,N_16898,N_16721);
or U19147 (N_19147,N_16450,N_16222);
nor U19148 (N_19148,N_16471,N_16334);
xor U19149 (N_19149,N_16501,N_17231);
nor U19150 (N_19150,N_16728,N_16771);
nor U19151 (N_19151,N_16127,N_16028);
xor U19152 (N_19152,N_17223,N_17552);
nand U19153 (N_19153,N_16349,N_16482);
xor U19154 (N_19154,N_16747,N_17936);
nor U19155 (N_19155,N_16656,N_16222);
and U19156 (N_19156,N_16933,N_16040);
and U19157 (N_19157,N_17701,N_17604);
nand U19158 (N_19158,N_16099,N_17278);
xnor U19159 (N_19159,N_17074,N_16488);
and U19160 (N_19160,N_16673,N_17372);
or U19161 (N_19161,N_17439,N_17374);
nor U19162 (N_19162,N_16491,N_17458);
or U19163 (N_19163,N_17905,N_16117);
or U19164 (N_19164,N_17984,N_16893);
nor U19165 (N_19165,N_16789,N_17801);
nor U19166 (N_19166,N_16936,N_17954);
xnor U19167 (N_19167,N_16780,N_16954);
nand U19168 (N_19168,N_16958,N_16322);
nand U19169 (N_19169,N_16348,N_17028);
or U19170 (N_19170,N_17730,N_16626);
nand U19171 (N_19171,N_17394,N_16420);
or U19172 (N_19172,N_17954,N_16697);
xnor U19173 (N_19173,N_16081,N_16623);
nand U19174 (N_19174,N_17283,N_16444);
and U19175 (N_19175,N_17552,N_17141);
and U19176 (N_19176,N_16696,N_17328);
nor U19177 (N_19177,N_16373,N_16624);
or U19178 (N_19178,N_16310,N_17477);
nand U19179 (N_19179,N_17175,N_17272);
xor U19180 (N_19180,N_16445,N_16666);
nand U19181 (N_19181,N_16960,N_17751);
nand U19182 (N_19182,N_16428,N_17345);
nor U19183 (N_19183,N_17663,N_17323);
or U19184 (N_19184,N_17741,N_16153);
nor U19185 (N_19185,N_16559,N_17194);
nand U19186 (N_19186,N_16124,N_17003);
and U19187 (N_19187,N_16820,N_17104);
and U19188 (N_19188,N_17821,N_16485);
xor U19189 (N_19189,N_17694,N_17900);
nor U19190 (N_19190,N_16564,N_17299);
xnor U19191 (N_19191,N_17200,N_17015);
and U19192 (N_19192,N_16694,N_16068);
nor U19193 (N_19193,N_16526,N_16143);
or U19194 (N_19194,N_17075,N_16288);
and U19195 (N_19195,N_17483,N_17415);
nor U19196 (N_19196,N_17413,N_17318);
xnor U19197 (N_19197,N_16789,N_17635);
and U19198 (N_19198,N_17605,N_16686);
nor U19199 (N_19199,N_17320,N_17646);
nor U19200 (N_19200,N_17654,N_16258);
and U19201 (N_19201,N_17790,N_17939);
nand U19202 (N_19202,N_16740,N_16308);
nand U19203 (N_19203,N_16950,N_17254);
nor U19204 (N_19204,N_16579,N_16604);
and U19205 (N_19205,N_16267,N_16306);
or U19206 (N_19206,N_17487,N_17183);
nand U19207 (N_19207,N_16869,N_17143);
or U19208 (N_19208,N_17016,N_16440);
or U19209 (N_19209,N_16970,N_16978);
or U19210 (N_19210,N_16834,N_17102);
nor U19211 (N_19211,N_16450,N_17618);
nand U19212 (N_19212,N_16980,N_16259);
and U19213 (N_19213,N_16763,N_16579);
nor U19214 (N_19214,N_17854,N_17646);
nand U19215 (N_19215,N_17058,N_16825);
nand U19216 (N_19216,N_17408,N_17117);
xor U19217 (N_19217,N_16195,N_17838);
or U19218 (N_19218,N_16530,N_16299);
nand U19219 (N_19219,N_17881,N_16760);
nand U19220 (N_19220,N_17151,N_16807);
and U19221 (N_19221,N_16724,N_17208);
or U19222 (N_19222,N_16619,N_17579);
nor U19223 (N_19223,N_16473,N_17401);
or U19224 (N_19224,N_16072,N_16753);
and U19225 (N_19225,N_16019,N_17441);
nor U19226 (N_19226,N_17947,N_16704);
or U19227 (N_19227,N_17110,N_16672);
nor U19228 (N_19228,N_17583,N_17755);
xnor U19229 (N_19229,N_16939,N_16756);
or U19230 (N_19230,N_17863,N_17550);
and U19231 (N_19231,N_16947,N_16028);
or U19232 (N_19232,N_16835,N_17528);
nand U19233 (N_19233,N_17054,N_16373);
and U19234 (N_19234,N_17213,N_16582);
or U19235 (N_19235,N_17265,N_16216);
xor U19236 (N_19236,N_17208,N_17201);
nor U19237 (N_19237,N_16281,N_16427);
nor U19238 (N_19238,N_16175,N_16749);
or U19239 (N_19239,N_17480,N_16743);
or U19240 (N_19240,N_16536,N_16165);
and U19241 (N_19241,N_16996,N_17054);
and U19242 (N_19242,N_16815,N_17603);
and U19243 (N_19243,N_17852,N_17413);
xor U19244 (N_19244,N_16284,N_16921);
nand U19245 (N_19245,N_17631,N_16890);
nand U19246 (N_19246,N_16102,N_16333);
xor U19247 (N_19247,N_16734,N_16982);
or U19248 (N_19248,N_17471,N_17381);
and U19249 (N_19249,N_17926,N_17510);
and U19250 (N_19250,N_17668,N_17446);
nand U19251 (N_19251,N_16396,N_16338);
xnor U19252 (N_19252,N_16717,N_17903);
xor U19253 (N_19253,N_16692,N_17626);
xnor U19254 (N_19254,N_16711,N_16871);
nor U19255 (N_19255,N_16021,N_16384);
nor U19256 (N_19256,N_16126,N_17043);
xnor U19257 (N_19257,N_17227,N_16790);
nand U19258 (N_19258,N_17283,N_16498);
nor U19259 (N_19259,N_17165,N_16648);
nand U19260 (N_19260,N_17459,N_16107);
and U19261 (N_19261,N_17485,N_16262);
and U19262 (N_19262,N_16537,N_16610);
or U19263 (N_19263,N_16634,N_17801);
and U19264 (N_19264,N_16956,N_17165);
and U19265 (N_19265,N_16467,N_16916);
nand U19266 (N_19266,N_17917,N_17308);
nor U19267 (N_19267,N_16352,N_16491);
nand U19268 (N_19268,N_16052,N_16885);
nand U19269 (N_19269,N_17597,N_16586);
and U19270 (N_19270,N_17464,N_16923);
xor U19271 (N_19271,N_16495,N_16961);
nor U19272 (N_19272,N_16785,N_16057);
xor U19273 (N_19273,N_17342,N_16954);
xor U19274 (N_19274,N_16231,N_17506);
nor U19275 (N_19275,N_17909,N_17215);
xor U19276 (N_19276,N_17926,N_17713);
xor U19277 (N_19277,N_16696,N_16332);
or U19278 (N_19278,N_17070,N_17685);
and U19279 (N_19279,N_16643,N_17364);
and U19280 (N_19280,N_16504,N_16534);
nand U19281 (N_19281,N_16700,N_16490);
and U19282 (N_19282,N_17268,N_16139);
and U19283 (N_19283,N_16197,N_17010);
or U19284 (N_19284,N_17020,N_17572);
xor U19285 (N_19285,N_16646,N_17315);
xor U19286 (N_19286,N_17134,N_17100);
or U19287 (N_19287,N_16038,N_16579);
nor U19288 (N_19288,N_16913,N_17070);
and U19289 (N_19289,N_16743,N_16364);
xor U19290 (N_19290,N_16387,N_17911);
nand U19291 (N_19291,N_17101,N_16548);
and U19292 (N_19292,N_16213,N_17732);
or U19293 (N_19293,N_17888,N_17708);
nand U19294 (N_19294,N_17067,N_17123);
nor U19295 (N_19295,N_17372,N_16311);
xor U19296 (N_19296,N_16980,N_17729);
xor U19297 (N_19297,N_17773,N_17356);
or U19298 (N_19298,N_17072,N_16549);
nor U19299 (N_19299,N_16005,N_16701);
or U19300 (N_19300,N_17254,N_16206);
nor U19301 (N_19301,N_16367,N_16900);
or U19302 (N_19302,N_17578,N_16800);
nor U19303 (N_19303,N_16488,N_16042);
or U19304 (N_19304,N_16414,N_17220);
and U19305 (N_19305,N_17914,N_17577);
nor U19306 (N_19306,N_16151,N_17620);
nand U19307 (N_19307,N_16538,N_16790);
xor U19308 (N_19308,N_16316,N_16754);
xor U19309 (N_19309,N_17535,N_17035);
or U19310 (N_19310,N_17522,N_17188);
and U19311 (N_19311,N_17612,N_16023);
xnor U19312 (N_19312,N_17480,N_16456);
xor U19313 (N_19313,N_16697,N_16210);
xnor U19314 (N_19314,N_16625,N_16148);
xnor U19315 (N_19315,N_16748,N_16685);
nand U19316 (N_19316,N_16156,N_17808);
nor U19317 (N_19317,N_17048,N_16752);
nand U19318 (N_19318,N_17409,N_16028);
and U19319 (N_19319,N_16893,N_17421);
or U19320 (N_19320,N_17061,N_17683);
and U19321 (N_19321,N_16097,N_16882);
and U19322 (N_19322,N_16382,N_17377);
nand U19323 (N_19323,N_16192,N_17064);
nor U19324 (N_19324,N_17578,N_16019);
and U19325 (N_19325,N_17030,N_17201);
and U19326 (N_19326,N_17411,N_17417);
xnor U19327 (N_19327,N_17837,N_17977);
and U19328 (N_19328,N_16277,N_17096);
nor U19329 (N_19329,N_17936,N_16695);
and U19330 (N_19330,N_17804,N_16741);
or U19331 (N_19331,N_17112,N_16088);
and U19332 (N_19332,N_17637,N_16649);
nand U19333 (N_19333,N_16530,N_16692);
or U19334 (N_19334,N_17861,N_16759);
or U19335 (N_19335,N_16599,N_16181);
or U19336 (N_19336,N_16534,N_16012);
and U19337 (N_19337,N_17665,N_16611);
nor U19338 (N_19338,N_17682,N_16922);
or U19339 (N_19339,N_17356,N_17953);
and U19340 (N_19340,N_16935,N_16766);
nand U19341 (N_19341,N_17696,N_17436);
or U19342 (N_19342,N_17252,N_17363);
and U19343 (N_19343,N_17597,N_17725);
xor U19344 (N_19344,N_17209,N_16668);
and U19345 (N_19345,N_16520,N_17627);
xnor U19346 (N_19346,N_16956,N_16125);
or U19347 (N_19347,N_16784,N_16250);
nor U19348 (N_19348,N_16412,N_16775);
or U19349 (N_19349,N_16305,N_17717);
nor U19350 (N_19350,N_17224,N_17042);
xnor U19351 (N_19351,N_16712,N_16834);
nand U19352 (N_19352,N_16990,N_17070);
xnor U19353 (N_19353,N_17871,N_17345);
or U19354 (N_19354,N_16670,N_16546);
xnor U19355 (N_19355,N_16430,N_16977);
xor U19356 (N_19356,N_17955,N_16516);
and U19357 (N_19357,N_17499,N_16637);
xnor U19358 (N_19358,N_17150,N_16412);
or U19359 (N_19359,N_17372,N_16774);
and U19360 (N_19360,N_17769,N_16461);
nor U19361 (N_19361,N_17082,N_17755);
xor U19362 (N_19362,N_17232,N_16403);
nor U19363 (N_19363,N_16294,N_16169);
nor U19364 (N_19364,N_17436,N_17673);
nand U19365 (N_19365,N_17789,N_16780);
xor U19366 (N_19366,N_16117,N_17749);
xnor U19367 (N_19367,N_16542,N_16192);
xnor U19368 (N_19368,N_17798,N_17890);
or U19369 (N_19369,N_17455,N_17925);
or U19370 (N_19370,N_16305,N_16543);
xor U19371 (N_19371,N_16236,N_17373);
xnor U19372 (N_19372,N_17138,N_16765);
nor U19373 (N_19373,N_17472,N_16828);
nand U19374 (N_19374,N_17369,N_17872);
nor U19375 (N_19375,N_17175,N_16513);
nor U19376 (N_19376,N_17056,N_17186);
nor U19377 (N_19377,N_16187,N_16084);
xor U19378 (N_19378,N_16256,N_16472);
nand U19379 (N_19379,N_16021,N_16639);
nor U19380 (N_19380,N_17215,N_16265);
nand U19381 (N_19381,N_16431,N_16519);
and U19382 (N_19382,N_16422,N_16393);
nor U19383 (N_19383,N_16709,N_16494);
nor U19384 (N_19384,N_16477,N_17354);
nand U19385 (N_19385,N_16512,N_17774);
and U19386 (N_19386,N_17515,N_17814);
xnor U19387 (N_19387,N_16284,N_17295);
nor U19388 (N_19388,N_16672,N_16801);
nand U19389 (N_19389,N_17560,N_17909);
nor U19390 (N_19390,N_16814,N_17266);
and U19391 (N_19391,N_16527,N_17546);
xnor U19392 (N_19392,N_16904,N_16465);
nand U19393 (N_19393,N_16771,N_17820);
nor U19394 (N_19394,N_16133,N_16934);
and U19395 (N_19395,N_16002,N_17436);
and U19396 (N_19396,N_16235,N_16953);
or U19397 (N_19397,N_16340,N_17364);
and U19398 (N_19398,N_16920,N_17984);
nand U19399 (N_19399,N_17911,N_16800);
xnor U19400 (N_19400,N_17677,N_16370);
nor U19401 (N_19401,N_16480,N_16623);
nor U19402 (N_19402,N_16405,N_16493);
nand U19403 (N_19403,N_17296,N_17315);
xor U19404 (N_19404,N_17382,N_16089);
nor U19405 (N_19405,N_16535,N_17443);
nor U19406 (N_19406,N_17825,N_16727);
xor U19407 (N_19407,N_16181,N_16909);
nand U19408 (N_19408,N_17466,N_17101);
or U19409 (N_19409,N_16672,N_16135);
or U19410 (N_19410,N_16531,N_17550);
nand U19411 (N_19411,N_16156,N_17287);
nor U19412 (N_19412,N_17947,N_17550);
nand U19413 (N_19413,N_16457,N_16495);
and U19414 (N_19414,N_17004,N_17231);
or U19415 (N_19415,N_16408,N_16218);
nand U19416 (N_19416,N_16101,N_17944);
nor U19417 (N_19417,N_16596,N_17714);
or U19418 (N_19418,N_17367,N_16558);
nor U19419 (N_19419,N_16096,N_17220);
or U19420 (N_19420,N_16705,N_16555);
xor U19421 (N_19421,N_17585,N_16810);
and U19422 (N_19422,N_16994,N_17089);
nor U19423 (N_19423,N_16093,N_17510);
nand U19424 (N_19424,N_17984,N_17327);
or U19425 (N_19425,N_16358,N_17115);
nor U19426 (N_19426,N_17939,N_16021);
xor U19427 (N_19427,N_17133,N_16235);
xnor U19428 (N_19428,N_17735,N_17098);
nor U19429 (N_19429,N_16295,N_16496);
nand U19430 (N_19430,N_17033,N_16744);
nand U19431 (N_19431,N_16253,N_16397);
and U19432 (N_19432,N_17808,N_16616);
or U19433 (N_19433,N_17752,N_16419);
nor U19434 (N_19434,N_16646,N_17764);
nor U19435 (N_19435,N_16646,N_16667);
nor U19436 (N_19436,N_17278,N_16453);
xor U19437 (N_19437,N_16560,N_16196);
and U19438 (N_19438,N_17310,N_16542);
or U19439 (N_19439,N_17493,N_17728);
or U19440 (N_19440,N_16760,N_17905);
nand U19441 (N_19441,N_17277,N_17387);
and U19442 (N_19442,N_17016,N_16695);
and U19443 (N_19443,N_17289,N_17436);
nand U19444 (N_19444,N_16872,N_17205);
or U19445 (N_19445,N_17783,N_16394);
xnor U19446 (N_19446,N_16768,N_17700);
nor U19447 (N_19447,N_17762,N_16331);
nor U19448 (N_19448,N_16682,N_16615);
xor U19449 (N_19449,N_17949,N_17832);
nand U19450 (N_19450,N_16440,N_17349);
xnor U19451 (N_19451,N_17590,N_17720);
nor U19452 (N_19452,N_16836,N_17185);
nor U19453 (N_19453,N_16039,N_17218);
nor U19454 (N_19454,N_17110,N_17943);
nand U19455 (N_19455,N_17799,N_16535);
xnor U19456 (N_19456,N_16578,N_17193);
and U19457 (N_19457,N_16797,N_16108);
nand U19458 (N_19458,N_17784,N_16364);
nand U19459 (N_19459,N_16431,N_16956);
nor U19460 (N_19460,N_17389,N_16937);
and U19461 (N_19461,N_16242,N_16489);
and U19462 (N_19462,N_16185,N_17303);
nand U19463 (N_19463,N_16691,N_17154);
nand U19464 (N_19464,N_17574,N_16446);
nor U19465 (N_19465,N_17200,N_17803);
xor U19466 (N_19466,N_17582,N_16765);
or U19467 (N_19467,N_16370,N_17278);
or U19468 (N_19468,N_17556,N_16247);
xnor U19469 (N_19469,N_16395,N_17394);
or U19470 (N_19470,N_17049,N_17328);
xnor U19471 (N_19471,N_17932,N_16602);
xor U19472 (N_19472,N_16559,N_17261);
nor U19473 (N_19473,N_16193,N_17449);
nor U19474 (N_19474,N_17310,N_17946);
or U19475 (N_19475,N_16268,N_16963);
and U19476 (N_19476,N_17953,N_16651);
nand U19477 (N_19477,N_17758,N_17648);
nand U19478 (N_19478,N_16626,N_16138);
or U19479 (N_19479,N_17053,N_16667);
nor U19480 (N_19480,N_17173,N_17978);
nor U19481 (N_19481,N_17780,N_16508);
nand U19482 (N_19482,N_16931,N_16991);
nand U19483 (N_19483,N_16593,N_17364);
or U19484 (N_19484,N_16258,N_16836);
nand U19485 (N_19485,N_17268,N_17919);
or U19486 (N_19486,N_17457,N_16296);
nand U19487 (N_19487,N_17272,N_17711);
xor U19488 (N_19488,N_16235,N_17135);
xor U19489 (N_19489,N_17252,N_16493);
and U19490 (N_19490,N_17492,N_17457);
or U19491 (N_19491,N_17467,N_17396);
nor U19492 (N_19492,N_16516,N_16840);
and U19493 (N_19493,N_17035,N_16260);
xnor U19494 (N_19494,N_16530,N_16938);
nand U19495 (N_19495,N_17229,N_16473);
nand U19496 (N_19496,N_17963,N_16815);
xor U19497 (N_19497,N_16511,N_17658);
xor U19498 (N_19498,N_17365,N_17885);
nand U19499 (N_19499,N_16116,N_16092);
xor U19500 (N_19500,N_16540,N_17564);
xor U19501 (N_19501,N_16994,N_16606);
or U19502 (N_19502,N_17980,N_17067);
xnor U19503 (N_19503,N_16839,N_16910);
or U19504 (N_19504,N_16526,N_16259);
nor U19505 (N_19505,N_16024,N_17739);
xor U19506 (N_19506,N_17143,N_17381);
xnor U19507 (N_19507,N_16424,N_16213);
or U19508 (N_19508,N_16237,N_16733);
and U19509 (N_19509,N_16611,N_16833);
or U19510 (N_19510,N_17627,N_16330);
xor U19511 (N_19511,N_17201,N_16191);
nor U19512 (N_19512,N_16818,N_17040);
nor U19513 (N_19513,N_17685,N_16252);
nor U19514 (N_19514,N_17414,N_16888);
or U19515 (N_19515,N_16909,N_17375);
nand U19516 (N_19516,N_17819,N_16861);
or U19517 (N_19517,N_17328,N_17512);
and U19518 (N_19518,N_16758,N_16592);
xor U19519 (N_19519,N_16448,N_16623);
or U19520 (N_19520,N_16539,N_17751);
xor U19521 (N_19521,N_17724,N_17416);
nand U19522 (N_19522,N_17119,N_16985);
nor U19523 (N_19523,N_17015,N_17321);
nand U19524 (N_19524,N_16046,N_17027);
xnor U19525 (N_19525,N_17939,N_17185);
or U19526 (N_19526,N_16500,N_17291);
or U19527 (N_19527,N_17412,N_17842);
xnor U19528 (N_19528,N_17898,N_16267);
nand U19529 (N_19529,N_16897,N_16342);
and U19530 (N_19530,N_16093,N_16260);
nand U19531 (N_19531,N_16633,N_17560);
or U19532 (N_19532,N_17932,N_16594);
or U19533 (N_19533,N_17712,N_16839);
and U19534 (N_19534,N_17244,N_16018);
nand U19535 (N_19535,N_16937,N_16106);
xnor U19536 (N_19536,N_17547,N_16412);
xor U19537 (N_19537,N_17986,N_17842);
nor U19538 (N_19538,N_17583,N_17877);
and U19539 (N_19539,N_16172,N_16005);
and U19540 (N_19540,N_16505,N_17540);
xnor U19541 (N_19541,N_16484,N_16619);
xor U19542 (N_19542,N_16663,N_17959);
and U19543 (N_19543,N_16132,N_16422);
xor U19544 (N_19544,N_16437,N_16660);
nand U19545 (N_19545,N_16502,N_17606);
xnor U19546 (N_19546,N_17668,N_17574);
nand U19547 (N_19547,N_17385,N_16616);
nand U19548 (N_19548,N_16333,N_16348);
nand U19549 (N_19549,N_17233,N_16433);
nor U19550 (N_19550,N_17292,N_17392);
nor U19551 (N_19551,N_17370,N_16675);
nor U19552 (N_19552,N_16769,N_17412);
or U19553 (N_19553,N_16826,N_17910);
or U19554 (N_19554,N_16117,N_17889);
or U19555 (N_19555,N_16129,N_17668);
xor U19556 (N_19556,N_17805,N_16466);
nand U19557 (N_19557,N_17787,N_16320);
or U19558 (N_19558,N_17033,N_17460);
and U19559 (N_19559,N_16158,N_17545);
nand U19560 (N_19560,N_16833,N_17847);
and U19561 (N_19561,N_17575,N_16375);
or U19562 (N_19562,N_16071,N_16446);
or U19563 (N_19563,N_16479,N_17421);
or U19564 (N_19564,N_17526,N_16623);
xor U19565 (N_19565,N_17746,N_17569);
xnor U19566 (N_19566,N_16724,N_16110);
nand U19567 (N_19567,N_16444,N_17496);
nand U19568 (N_19568,N_16494,N_16413);
xor U19569 (N_19569,N_17057,N_17042);
and U19570 (N_19570,N_16091,N_17694);
or U19571 (N_19571,N_17696,N_17412);
xor U19572 (N_19572,N_17788,N_16086);
nand U19573 (N_19573,N_16179,N_16163);
xor U19574 (N_19574,N_17322,N_16284);
and U19575 (N_19575,N_17095,N_16404);
xnor U19576 (N_19576,N_16303,N_17006);
or U19577 (N_19577,N_16895,N_17498);
and U19578 (N_19578,N_16841,N_16610);
and U19579 (N_19579,N_16295,N_17398);
or U19580 (N_19580,N_16218,N_17180);
nor U19581 (N_19581,N_17475,N_16868);
nor U19582 (N_19582,N_16361,N_17189);
nand U19583 (N_19583,N_17652,N_16030);
nor U19584 (N_19584,N_16485,N_17382);
and U19585 (N_19585,N_17799,N_17063);
nor U19586 (N_19586,N_17243,N_17448);
nand U19587 (N_19587,N_17377,N_16728);
or U19588 (N_19588,N_16840,N_17551);
or U19589 (N_19589,N_16474,N_17319);
xor U19590 (N_19590,N_16674,N_17309);
nor U19591 (N_19591,N_16247,N_17882);
or U19592 (N_19592,N_16915,N_17397);
nor U19593 (N_19593,N_17537,N_17907);
xor U19594 (N_19594,N_16604,N_16515);
xor U19595 (N_19595,N_17348,N_17956);
or U19596 (N_19596,N_17561,N_17708);
xor U19597 (N_19597,N_17737,N_16412);
nand U19598 (N_19598,N_16690,N_17720);
nor U19599 (N_19599,N_17372,N_17457);
nor U19600 (N_19600,N_17491,N_16198);
or U19601 (N_19601,N_17618,N_16535);
and U19602 (N_19602,N_17624,N_16501);
nand U19603 (N_19603,N_17159,N_16028);
nand U19604 (N_19604,N_17588,N_16453);
or U19605 (N_19605,N_17739,N_16184);
or U19606 (N_19606,N_16269,N_16262);
nor U19607 (N_19607,N_17492,N_17584);
xor U19608 (N_19608,N_17077,N_17064);
or U19609 (N_19609,N_16078,N_16235);
nand U19610 (N_19610,N_17187,N_16424);
and U19611 (N_19611,N_17471,N_16989);
and U19612 (N_19612,N_17927,N_17203);
and U19613 (N_19613,N_16633,N_16227);
or U19614 (N_19614,N_16060,N_16236);
or U19615 (N_19615,N_17633,N_16799);
xor U19616 (N_19616,N_16723,N_16792);
nor U19617 (N_19617,N_16825,N_17104);
nor U19618 (N_19618,N_16296,N_17909);
or U19619 (N_19619,N_17057,N_16767);
xor U19620 (N_19620,N_16962,N_17317);
nor U19621 (N_19621,N_17588,N_16150);
nor U19622 (N_19622,N_16042,N_17328);
xnor U19623 (N_19623,N_16353,N_16065);
or U19624 (N_19624,N_16409,N_16717);
xor U19625 (N_19625,N_17789,N_17783);
or U19626 (N_19626,N_17965,N_17164);
xor U19627 (N_19627,N_16726,N_17074);
nor U19628 (N_19628,N_17482,N_16391);
or U19629 (N_19629,N_17378,N_16049);
and U19630 (N_19630,N_17460,N_17038);
and U19631 (N_19631,N_17661,N_17688);
nor U19632 (N_19632,N_17263,N_17898);
and U19633 (N_19633,N_16350,N_17670);
and U19634 (N_19634,N_16998,N_16173);
and U19635 (N_19635,N_16983,N_16749);
xnor U19636 (N_19636,N_17288,N_17297);
xnor U19637 (N_19637,N_17565,N_16291);
xnor U19638 (N_19638,N_16192,N_17305);
and U19639 (N_19639,N_16894,N_16221);
nand U19640 (N_19640,N_16573,N_17297);
nand U19641 (N_19641,N_16863,N_16069);
or U19642 (N_19642,N_17247,N_17402);
nand U19643 (N_19643,N_16367,N_16494);
nor U19644 (N_19644,N_16997,N_16854);
nand U19645 (N_19645,N_17226,N_16342);
and U19646 (N_19646,N_16518,N_16844);
nor U19647 (N_19647,N_17454,N_17265);
or U19648 (N_19648,N_17703,N_16463);
nor U19649 (N_19649,N_17295,N_16699);
nor U19650 (N_19650,N_17945,N_17816);
nand U19651 (N_19651,N_16903,N_17766);
or U19652 (N_19652,N_16363,N_17078);
xnor U19653 (N_19653,N_16304,N_17597);
nand U19654 (N_19654,N_17005,N_16869);
xor U19655 (N_19655,N_17052,N_16630);
xnor U19656 (N_19656,N_16024,N_17963);
nand U19657 (N_19657,N_17428,N_17635);
and U19658 (N_19658,N_16904,N_16603);
or U19659 (N_19659,N_17157,N_17241);
nor U19660 (N_19660,N_16759,N_16248);
and U19661 (N_19661,N_17672,N_16991);
or U19662 (N_19662,N_16797,N_17242);
and U19663 (N_19663,N_16575,N_17728);
nor U19664 (N_19664,N_17673,N_16136);
nand U19665 (N_19665,N_17850,N_17743);
nor U19666 (N_19666,N_16357,N_17519);
nand U19667 (N_19667,N_16230,N_16875);
xor U19668 (N_19668,N_17542,N_17339);
or U19669 (N_19669,N_16338,N_16883);
nor U19670 (N_19670,N_17525,N_17372);
and U19671 (N_19671,N_17001,N_16474);
or U19672 (N_19672,N_16354,N_16218);
nand U19673 (N_19673,N_16942,N_17188);
nor U19674 (N_19674,N_16826,N_17521);
nor U19675 (N_19675,N_17204,N_16055);
and U19676 (N_19676,N_17616,N_17348);
or U19677 (N_19677,N_16851,N_17130);
or U19678 (N_19678,N_16588,N_17246);
and U19679 (N_19679,N_16102,N_17515);
or U19680 (N_19680,N_17683,N_17736);
nor U19681 (N_19681,N_17460,N_16520);
xnor U19682 (N_19682,N_17846,N_17589);
nand U19683 (N_19683,N_17395,N_17505);
nor U19684 (N_19684,N_17901,N_16688);
nand U19685 (N_19685,N_16989,N_16244);
xnor U19686 (N_19686,N_17949,N_16098);
nor U19687 (N_19687,N_17884,N_16163);
and U19688 (N_19688,N_16721,N_16929);
nor U19689 (N_19689,N_17505,N_16620);
and U19690 (N_19690,N_17027,N_16728);
and U19691 (N_19691,N_16435,N_16017);
xor U19692 (N_19692,N_16427,N_17064);
or U19693 (N_19693,N_17731,N_16937);
or U19694 (N_19694,N_16487,N_16607);
nand U19695 (N_19695,N_16770,N_16702);
or U19696 (N_19696,N_17804,N_16023);
and U19697 (N_19697,N_17899,N_16395);
nor U19698 (N_19698,N_17142,N_16696);
nor U19699 (N_19699,N_17274,N_16672);
xnor U19700 (N_19700,N_16048,N_17013);
nand U19701 (N_19701,N_17473,N_17582);
and U19702 (N_19702,N_16367,N_16878);
nand U19703 (N_19703,N_16612,N_17131);
nand U19704 (N_19704,N_17480,N_16379);
and U19705 (N_19705,N_16260,N_16686);
or U19706 (N_19706,N_16168,N_16774);
xor U19707 (N_19707,N_16586,N_17666);
xnor U19708 (N_19708,N_16192,N_17462);
xor U19709 (N_19709,N_16622,N_17288);
xor U19710 (N_19710,N_16125,N_17175);
xnor U19711 (N_19711,N_16189,N_16392);
nor U19712 (N_19712,N_16181,N_17222);
nor U19713 (N_19713,N_16385,N_17728);
or U19714 (N_19714,N_16721,N_17802);
xor U19715 (N_19715,N_17302,N_17800);
or U19716 (N_19716,N_17800,N_17891);
and U19717 (N_19717,N_16469,N_17588);
and U19718 (N_19718,N_16362,N_17732);
xor U19719 (N_19719,N_17425,N_16346);
xnor U19720 (N_19720,N_16339,N_17339);
xor U19721 (N_19721,N_17218,N_16708);
nand U19722 (N_19722,N_16693,N_16759);
nor U19723 (N_19723,N_17970,N_16144);
or U19724 (N_19724,N_16995,N_16011);
and U19725 (N_19725,N_17958,N_17465);
or U19726 (N_19726,N_16813,N_16150);
and U19727 (N_19727,N_16488,N_17550);
nor U19728 (N_19728,N_17070,N_17169);
nand U19729 (N_19729,N_17204,N_17693);
and U19730 (N_19730,N_16479,N_17764);
or U19731 (N_19731,N_17418,N_17593);
nor U19732 (N_19732,N_16011,N_17483);
and U19733 (N_19733,N_16832,N_16166);
nand U19734 (N_19734,N_17507,N_17462);
xor U19735 (N_19735,N_17080,N_17674);
xor U19736 (N_19736,N_16371,N_17702);
or U19737 (N_19737,N_17583,N_16806);
nor U19738 (N_19738,N_16131,N_17634);
xnor U19739 (N_19739,N_16324,N_16353);
nor U19740 (N_19740,N_16951,N_17830);
or U19741 (N_19741,N_17645,N_16037);
nor U19742 (N_19742,N_16998,N_17250);
and U19743 (N_19743,N_17762,N_16523);
or U19744 (N_19744,N_17725,N_17310);
or U19745 (N_19745,N_17951,N_16348);
or U19746 (N_19746,N_17237,N_16632);
xor U19747 (N_19747,N_16786,N_16448);
xnor U19748 (N_19748,N_17799,N_16169);
nand U19749 (N_19749,N_16162,N_16226);
xor U19750 (N_19750,N_16253,N_17681);
xor U19751 (N_19751,N_16993,N_17553);
and U19752 (N_19752,N_17536,N_16388);
xnor U19753 (N_19753,N_16705,N_17924);
nand U19754 (N_19754,N_16951,N_16647);
and U19755 (N_19755,N_17370,N_16189);
xnor U19756 (N_19756,N_17827,N_16990);
nand U19757 (N_19757,N_16261,N_17256);
xor U19758 (N_19758,N_17762,N_17953);
and U19759 (N_19759,N_17533,N_16008);
nor U19760 (N_19760,N_17239,N_16856);
or U19761 (N_19761,N_16812,N_16940);
nor U19762 (N_19762,N_16441,N_17100);
nor U19763 (N_19763,N_17626,N_17322);
nand U19764 (N_19764,N_17335,N_16257);
and U19765 (N_19765,N_17063,N_16645);
and U19766 (N_19766,N_16556,N_16808);
nor U19767 (N_19767,N_16757,N_16468);
or U19768 (N_19768,N_16140,N_17351);
or U19769 (N_19769,N_16733,N_16678);
nor U19770 (N_19770,N_17753,N_16311);
or U19771 (N_19771,N_17298,N_16800);
and U19772 (N_19772,N_16200,N_17346);
xnor U19773 (N_19773,N_16982,N_16749);
xor U19774 (N_19774,N_16270,N_17621);
nand U19775 (N_19775,N_16335,N_17298);
and U19776 (N_19776,N_17541,N_17810);
xnor U19777 (N_19777,N_17790,N_17606);
and U19778 (N_19778,N_16905,N_17738);
xor U19779 (N_19779,N_17122,N_16697);
or U19780 (N_19780,N_16831,N_17917);
nor U19781 (N_19781,N_17277,N_17448);
or U19782 (N_19782,N_16665,N_16714);
nand U19783 (N_19783,N_16899,N_17092);
nand U19784 (N_19784,N_17099,N_17128);
and U19785 (N_19785,N_16215,N_16915);
and U19786 (N_19786,N_16987,N_17586);
xnor U19787 (N_19787,N_17569,N_16245);
xnor U19788 (N_19788,N_16449,N_16888);
xnor U19789 (N_19789,N_16468,N_17211);
xor U19790 (N_19790,N_16158,N_17286);
and U19791 (N_19791,N_17146,N_17447);
and U19792 (N_19792,N_16344,N_16316);
nor U19793 (N_19793,N_17288,N_16624);
or U19794 (N_19794,N_16856,N_16650);
nand U19795 (N_19795,N_16415,N_16199);
xor U19796 (N_19796,N_16668,N_17160);
nor U19797 (N_19797,N_16024,N_17924);
nor U19798 (N_19798,N_17844,N_16221);
nor U19799 (N_19799,N_16731,N_17604);
and U19800 (N_19800,N_17672,N_17768);
xor U19801 (N_19801,N_17131,N_17219);
and U19802 (N_19802,N_17270,N_17473);
or U19803 (N_19803,N_16714,N_16132);
or U19804 (N_19804,N_16091,N_17963);
nand U19805 (N_19805,N_17026,N_16113);
nor U19806 (N_19806,N_16257,N_17710);
nor U19807 (N_19807,N_16471,N_16084);
nand U19808 (N_19808,N_16846,N_17453);
or U19809 (N_19809,N_16216,N_16265);
or U19810 (N_19810,N_17495,N_17761);
nor U19811 (N_19811,N_16341,N_17545);
or U19812 (N_19812,N_17817,N_16857);
nand U19813 (N_19813,N_17047,N_16024);
nand U19814 (N_19814,N_17067,N_16247);
or U19815 (N_19815,N_16399,N_17788);
xnor U19816 (N_19816,N_16284,N_17992);
nand U19817 (N_19817,N_16564,N_16245);
nand U19818 (N_19818,N_16710,N_16688);
or U19819 (N_19819,N_16155,N_16583);
or U19820 (N_19820,N_16624,N_17471);
xor U19821 (N_19821,N_17396,N_17501);
nor U19822 (N_19822,N_16398,N_17760);
and U19823 (N_19823,N_16956,N_17671);
xnor U19824 (N_19824,N_17504,N_17052);
and U19825 (N_19825,N_17577,N_17352);
xor U19826 (N_19826,N_17898,N_17628);
nor U19827 (N_19827,N_16765,N_16363);
xnor U19828 (N_19828,N_17731,N_16742);
nor U19829 (N_19829,N_17529,N_17449);
xnor U19830 (N_19830,N_17818,N_17976);
nand U19831 (N_19831,N_16984,N_17940);
or U19832 (N_19832,N_17772,N_17016);
and U19833 (N_19833,N_16502,N_16794);
or U19834 (N_19834,N_16751,N_17885);
xnor U19835 (N_19835,N_17698,N_16616);
nand U19836 (N_19836,N_16252,N_17133);
xor U19837 (N_19837,N_17120,N_17271);
xor U19838 (N_19838,N_16620,N_16550);
nand U19839 (N_19839,N_16721,N_17351);
nor U19840 (N_19840,N_17012,N_17961);
nor U19841 (N_19841,N_17071,N_16497);
nand U19842 (N_19842,N_17189,N_16895);
nand U19843 (N_19843,N_16570,N_16422);
or U19844 (N_19844,N_16364,N_17626);
or U19845 (N_19845,N_17171,N_16190);
nor U19846 (N_19846,N_17156,N_16913);
and U19847 (N_19847,N_16274,N_16732);
or U19848 (N_19848,N_16360,N_16831);
or U19849 (N_19849,N_16170,N_17792);
xor U19850 (N_19850,N_16899,N_16815);
or U19851 (N_19851,N_17312,N_17467);
nor U19852 (N_19852,N_17831,N_16814);
and U19853 (N_19853,N_17444,N_16127);
nand U19854 (N_19854,N_16715,N_16449);
nand U19855 (N_19855,N_17877,N_17733);
nand U19856 (N_19856,N_16337,N_17517);
nand U19857 (N_19857,N_16941,N_16645);
nor U19858 (N_19858,N_17726,N_16353);
nor U19859 (N_19859,N_17384,N_16897);
nor U19860 (N_19860,N_16448,N_17613);
or U19861 (N_19861,N_16799,N_17362);
and U19862 (N_19862,N_16560,N_16543);
or U19863 (N_19863,N_16121,N_16695);
xnor U19864 (N_19864,N_17884,N_17046);
nor U19865 (N_19865,N_16956,N_16984);
nor U19866 (N_19866,N_17334,N_16673);
and U19867 (N_19867,N_16610,N_16903);
xnor U19868 (N_19868,N_16479,N_17424);
nand U19869 (N_19869,N_16367,N_16169);
and U19870 (N_19870,N_16985,N_16943);
or U19871 (N_19871,N_16558,N_17157);
nand U19872 (N_19872,N_17161,N_17583);
and U19873 (N_19873,N_16769,N_17528);
and U19874 (N_19874,N_17000,N_17181);
nor U19875 (N_19875,N_16326,N_17315);
nor U19876 (N_19876,N_16599,N_17132);
and U19877 (N_19877,N_17020,N_16748);
nor U19878 (N_19878,N_17048,N_16723);
and U19879 (N_19879,N_17141,N_17401);
and U19880 (N_19880,N_16670,N_16256);
or U19881 (N_19881,N_16944,N_16001);
or U19882 (N_19882,N_16988,N_16231);
nand U19883 (N_19883,N_17368,N_17003);
or U19884 (N_19884,N_16894,N_16637);
and U19885 (N_19885,N_16837,N_16405);
and U19886 (N_19886,N_16921,N_16794);
nor U19887 (N_19887,N_17148,N_17541);
and U19888 (N_19888,N_16278,N_16530);
and U19889 (N_19889,N_17334,N_16606);
or U19890 (N_19890,N_17619,N_17355);
nand U19891 (N_19891,N_16183,N_17544);
xnor U19892 (N_19892,N_16108,N_17023);
and U19893 (N_19893,N_16267,N_17648);
nand U19894 (N_19894,N_16965,N_17723);
nor U19895 (N_19895,N_17133,N_17507);
or U19896 (N_19896,N_17810,N_16458);
xor U19897 (N_19897,N_16066,N_17011);
or U19898 (N_19898,N_16958,N_16872);
nand U19899 (N_19899,N_17552,N_16300);
nor U19900 (N_19900,N_17817,N_16437);
or U19901 (N_19901,N_17097,N_16429);
nand U19902 (N_19902,N_17754,N_16254);
nand U19903 (N_19903,N_16563,N_17038);
nand U19904 (N_19904,N_17996,N_17487);
and U19905 (N_19905,N_16263,N_16242);
nand U19906 (N_19906,N_17424,N_17001);
xnor U19907 (N_19907,N_16287,N_16930);
and U19908 (N_19908,N_17172,N_17521);
nand U19909 (N_19909,N_16448,N_16721);
and U19910 (N_19910,N_16613,N_17985);
and U19911 (N_19911,N_16995,N_17684);
or U19912 (N_19912,N_16524,N_16452);
xnor U19913 (N_19913,N_16379,N_17628);
nand U19914 (N_19914,N_16868,N_17548);
or U19915 (N_19915,N_16457,N_16797);
xnor U19916 (N_19916,N_16835,N_17610);
nor U19917 (N_19917,N_16427,N_17758);
and U19918 (N_19918,N_17280,N_16659);
nor U19919 (N_19919,N_16569,N_17812);
xor U19920 (N_19920,N_16546,N_16936);
xor U19921 (N_19921,N_16391,N_16265);
xnor U19922 (N_19922,N_17842,N_17166);
or U19923 (N_19923,N_16182,N_16499);
or U19924 (N_19924,N_16491,N_17966);
nand U19925 (N_19925,N_17475,N_17894);
nor U19926 (N_19926,N_17719,N_17846);
and U19927 (N_19927,N_17167,N_17163);
or U19928 (N_19928,N_17467,N_16923);
and U19929 (N_19929,N_17897,N_17991);
nand U19930 (N_19930,N_16258,N_16763);
xor U19931 (N_19931,N_16522,N_16259);
or U19932 (N_19932,N_16069,N_17552);
and U19933 (N_19933,N_17556,N_17039);
nand U19934 (N_19934,N_17159,N_17741);
nand U19935 (N_19935,N_17178,N_17601);
nand U19936 (N_19936,N_16193,N_17787);
xor U19937 (N_19937,N_17251,N_16234);
xnor U19938 (N_19938,N_17979,N_17282);
xor U19939 (N_19939,N_16309,N_17730);
nand U19940 (N_19940,N_16214,N_17557);
xnor U19941 (N_19941,N_16693,N_17341);
and U19942 (N_19942,N_16087,N_16619);
xor U19943 (N_19943,N_16644,N_17004);
or U19944 (N_19944,N_17768,N_17467);
xnor U19945 (N_19945,N_17526,N_16665);
nand U19946 (N_19946,N_16212,N_17893);
nor U19947 (N_19947,N_16273,N_17926);
or U19948 (N_19948,N_16956,N_16447);
nor U19949 (N_19949,N_16517,N_17980);
or U19950 (N_19950,N_17806,N_16916);
and U19951 (N_19951,N_16659,N_16308);
nand U19952 (N_19952,N_16059,N_16684);
xor U19953 (N_19953,N_16451,N_16874);
or U19954 (N_19954,N_17526,N_17905);
and U19955 (N_19955,N_17824,N_17764);
nor U19956 (N_19956,N_16147,N_16879);
xor U19957 (N_19957,N_16645,N_17609);
nor U19958 (N_19958,N_16518,N_17387);
and U19959 (N_19959,N_16655,N_17406);
xor U19960 (N_19960,N_17733,N_16725);
and U19961 (N_19961,N_16169,N_16158);
xnor U19962 (N_19962,N_16532,N_17954);
nor U19963 (N_19963,N_16378,N_16742);
nand U19964 (N_19964,N_16268,N_17431);
nor U19965 (N_19965,N_16769,N_16848);
or U19966 (N_19966,N_17080,N_16181);
and U19967 (N_19967,N_16903,N_17295);
nand U19968 (N_19968,N_17215,N_16554);
and U19969 (N_19969,N_17743,N_17403);
xor U19970 (N_19970,N_16934,N_17244);
or U19971 (N_19971,N_17736,N_16790);
xnor U19972 (N_19972,N_17895,N_17453);
and U19973 (N_19973,N_16991,N_17686);
xnor U19974 (N_19974,N_16479,N_17516);
or U19975 (N_19975,N_16185,N_16400);
or U19976 (N_19976,N_17238,N_17769);
nor U19977 (N_19977,N_16666,N_17459);
and U19978 (N_19978,N_17784,N_17752);
and U19979 (N_19979,N_16468,N_17750);
nand U19980 (N_19980,N_17009,N_17639);
xnor U19981 (N_19981,N_16430,N_17996);
xor U19982 (N_19982,N_16271,N_16413);
xor U19983 (N_19983,N_16104,N_17188);
and U19984 (N_19984,N_16412,N_16534);
nor U19985 (N_19985,N_16756,N_16137);
and U19986 (N_19986,N_16872,N_16816);
nor U19987 (N_19987,N_17533,N_16968);
nand U19988 (N_19988,N_17484,N_17521);
xnor U19989 (N_19989,N_17711,N_16097);
and U19990 (N_19990,N_16918,N_16554);
nand U19991 (N_19991,N_16864,N_17986);
and U19992 (N_19992,N_16476,N_16657);
nor U19993 (N_19993,N_17236,N_17345);
nand U19994 (N_19994,N_17082,N_16187);
and U19995 (N_19995,N_17410,N_17312);
nand U19996 (N_19996,N_16498,N_17614);
xnor U19997 (N_19997,N_16967,N_17687);
nand U19998 (N_19998,N_16373,N_16028);
or U19999 (N_19999,N_17477,N_17962);
xor U20000 (N_20000,N_18509,N_19071);
or U20001 (N_20001,N_18741,N_18133);
nor U20002 (N_20002,N_18989,N_19370);
xnor U20003 (N_20003,N_18297,N_19368);
xor U20004 (N_20004,N_18091,N_19907);
nor U20005 (N_20005,N_19218,N_19652);
nor U20006 (N_20006,N_19022,N_18051);
and U20007 (N_20007,N_18959,N_18074);
nor U20008 (N_20008,N_18916,N_18217);
and U20009 (N_20009,N_19346,N_19797);
and U20010 (N_20010,N_18322,N_18540);
nand U20011 (N_20011,N_19868,N_18777);
nand U20012 (N_20012,N_19972,N_19965);
or U20013 (N_20013,N_18566,N_18276);
nor U20014 (N_20014,N_18819,N_19162);
and U20015 (N_20015,N_18653,N_18801);
nand U20016 (N_20016,N_19026,N_18645);
and U20017 (N_20017,N_18225,N_19188);
xor U20018 (N_20018,N_18579,N_19411);
nor U20019 (N_20019,N_19962,N_18630);
nand U20020 (N_20020,N_19204,N_18414);
and U20021 (N_20021,N_18479,N_19854);
or U20022 (N_20022,N_19436,N_19387);
xnor U20023 (N_20023,N_18665,N_18214);
nor U20024 (N_20024,N_19432,N_19486);
and U20025 (N_20025,N_19722,N_18734);
nand U20026 (N_20026,N_19145,N_18977);
and U20027 (N_20027,N_19817,N_18657);
and U20028 (N_20028,N_19258,N_19135);
and U20029 (N_20029,N_18443,N_19560);
or U20030 (N_20030,N_18692,N_18094);
xor U20031 (N_20031,N_19030,N_18332);
and U20032 (N_20032,N_19597,N_19651);
xnor U20033 (N_20033,N_18289,N_18023);
nor U20034 (N_20034,N_18009,N_18818);
nand U20035 (N_20035,N_18444,N_18054);
and U20036 (N_20036,N_19826,N_18413);
or U20037 (N_20037,N_19142,N_19016);
or U20038 (N_20038,N_19447,N_19985);
or U20039 (N_20039,N_18223,N_18447);
nor U20040 (N_20040,N_18542,N_19910);
nor U20041 (N_20041,N_19841,N_19875);
or U20042 (N_20042,N_18328,N_18427);
nor U20043 (N_20043,N_18713,N_19795);
xnor U20044 (N_20044,N_18753,N_19878);
xor U20045 (N_20045,N_19488,N_19227);
and U20046 (N_20046,N_18655,N_19290);
nand U20047 (N_20047,N_18370,N_18361);
nand U20048 (N_20048,N_18586,N_19784);
and U20049 (N_20049,N_19602,N_19533);
nand U20050 (N_20050,N_18319,N_19889);
xor U20051 (N_20051,N_19173,N_19814);
xor U20052 (N_20052,N_18164,N_19518);
or U20053 (N_20053,N_19916,N_18191);
xor U20054 (N_20054,N_18978,N_19674);
nand U20055 (N_20055,N_18710,N_18382);
nand U20056 (N_20056,N_18696,N_18338);
or U20057 (N_20057,N_19305,N_19561);
and U20058 (N_20058,N_19372,N_18593);
xor U20059 (N_20059,N_18504,N_18458);
or U20060 (N_20060,N_19009,N_19120);
nand U20061 (N_20061,N_19821,N_19452);
nand U20062 (N_20062,N_19014,N_18470);
or U20063 (N_20063,N_18175,N_18534);
nor U20064 (N_20064,N_18851,N_18949);
xnor U20065 (N_20065,N_19017,N_19942);
nor U20066 (N_20066,N_18431,N_18475);
xnor U20067 (N_20067,N_18451,N_19221);
nor U20068 (N_20068,N_18138,N_18092);
nand U20069 (N_20069,N_18111,N_19871);
and U20070 (N_20070,N_19225,N_19152);
or U20071 (N_20071,N_19957,N_19610);
xor U20072 (N_20072,N_18262,N_19523);
nand U20073 (N_20073,N_19006,N_18986);
xnor U20074 (N_20074,N_19742,N_18086);
and U20075 (N_20075,N_18488,N_18997);
nand U20076 (N_20076,N_19124,N_18416);
nor U20077 (N_20077,N_19935,N_18880);
nor U20078 (N_20078,N_18898,N_18562);
nor U20079 (N_20079,N_18599,N_19930);
xnor U20080 (N_20080,N_18151,N_19384);
or U20081 (N_20081,N_19966,N_18429);
or U20082 (N_20082,N_18668,N_19770);
and U20083 (N_20083,N_18169,N_18037);
nand U20084 (N_20084,N_18614,N_19214);
or U20085 (N_20085,N_19856,N_19147);
and U20086 (N_20086,N_19960,N_19051);
or U20087 (N_20087,N_18919,N_18013);
or U20088 (N_20088,N_18893,N_18102);
nand U20089 (N_20089,N_19267,N_18574);
nand U20090 (N_20090,N_18596,N_18926);
nor U20091 (N_20091,N_19213,N_18400);
and U20092 (N_20092,N_18670,N_18639);
nand U20093 (N_20093,N_18021,N_19616);
nor U20094 (N_20094,N_19023,N_19681);
and U20095 (N_20095,N_18501,N_18686);
nor U20096 (N_20096,N_19105,N_19077);
or U20097 (N_20097,N_19280,N_19724);
nand U20098 (N_20098,N_19877,N_18077);
nand U20099 (N_20099,N_18290,N_18136);
or U20100 (N_20100,N_18106,N_19229);
nand U20101 (N_20101,N_19947,N_18031);
or U20102 (N_20102,N_19441,N_19684);
nand U20103 (N_20103,N_18915,N_18292);
and U20104 (N_20104,N_18465,N_19076);
nand U20105 (N_20105,N_19888,N_19198);
or U20106 (N_20106,N_18702,N_19607);
or U20107 (N_20107,N_18863,N_19352);
xnor U20108 (N_20108,N_18493,N_19235);
or U20109 (N_20109,N_18269,N_18385);
or U20110 (N_20110,N_18983,N_18036);
or U20111 (N_20111,N_19970,N_18409);
nand U20112 (N_20112,N_19139,N_19442);
or U20113 (N_20113,N_18640,N_19785);
xor U20114 (N_20114,N_19024,N_19578);
or U20115 (N_20115,N_19589,N_19163);
nand U20116 (N_20116,N_18003,N_19477);
xnor U20117 (N_20117,N_19825,N_19294);
nor U20118 (N_20118,N_19662,N_18236);
and U20119 (N_20119,N_19603,N_18934);
and U20120 (N_20120,N_18399,N_19861);
or U20121 (N_20121,N_19033,N_19881);
and U20122 (N_20122,N_19648,N_18503);
xor U20123 (N_20123,N_18817,N_18519);
or U20124 (N_20124,N_18162,N_18277);
and U20125 (N_20125,N_19391,N_19453);
xnor U20126 (N_20126,N_19563,N_19404);
or U20127 (N_20127,N_18707,N_19159);
and U20128 (N_20128,N_19657,N_19838);
and U20129 (N_20129,N_18766,N_18837);
and U20130 (N_20130,N_19559,N_18324);
and U20131 (N_20131,N_18412,N_18500);
nand U20132 (N_20132,N_18394,N_18224);
xor U20133 (N_20133,N_18812,N_18852);
and U20134 (N_20134,N_19997,N_19679);
nand U20135 (N_20135,N_19572,N_19382);
nand U20136 (N_20136,N_18129,N_19176);
xnor U20137 (N_20137,N_18721,N_18404);
nand U20138 (N_20138,N_18762,N_18219);
or U20139 (N_20139,N_19010,N_19349);
nand U20140 (N_20140,N_19958,N_19999);
or U20141 (N_20141,N_18316,N_19031);
xor U20142 (N_20142,N_18815,N_18284);
and U20143 (N_20143,N_18580,N_19775);
or U20144 (N_20144,N_19101,N_19641);
xor U20145 (N_20145,N_19226,N_18325);
or U20146 (N_20146,N_18103,N_18520);
nand U20147 (N_20147,N_19160,N_18252);
nor U20148 (N_20148,N_18093,N_19203);
or U20149 (N_20149,N_19569,N_19329);
nor U20150 (N_20150,N_19104,N_19579);
or U20151 (N_20151,N_18623,N_18747);
nor U20152 (N_20152,N_19245,N_18468);
xor U20153 (N_20153,N_19738,N_18226);
nand U20154 (N_20154,N_18049,N_19703);
and U20155 (N_20155,N_19315,N_18903);
nor U20156 (N_20156,N_19116,N_19624);
and U20157 (N_20157,N_18795,N_18797);
nand U20158 (N_20158,N_18785,N_19417);
and U20159 (N_20159,N_19704,N_19983);
and U20160 (N_20160,N_18672,N_18492);
or U20161 (N_20161,N_18963,N_18275);
or U20162 (N_20162,N_19260,N_19587);
and U20163 (N_20163,N_19081,N_18460);
or U20164 (N_20164,N_18778,N_18463);
nor U20165 (N_20165,N_18570,N_19098);
nor U20166 (N_20166,N_18867,N_18188);
xor U20167 (N_20167,N_18552,N_19761);
xor U20168 (N_20168,N_19951,N_18397);
nand U20169 (N_20169,N_19783,N_18714);
nand U20170 (N_20170,N_19476,N_18548);
and U20171 (N_20171,N_18078,N_19858);
and U20172 (N_20172,N_19740,N_19397);
nor U20173 (N_20173,N_19255,N_19117);
and U20174 (N_20174,N_18112,N_19677);
nand U20175 (N_20175,N_19181,N_19451);
xor U20176 (N_20176,N_18660,N_18740);
xor U20177 (N_20177,N_19802,N_18245);
and U20178 (N_20178,N_19836,N_19425);
nor U20179 (N_20179,N_19507,N_18287);
xnor U20180 (N_20180,N_19330,N_18845);
xor U20181 (N_20181,N_19720,N_18098);
nor U20182 (N_20182,N_18180,N_19036);
and U20183 (N_20183,N_18947,N_19243);
xnor U20184 (N_20184,N_19727,N_18896);
nor U20185 (N_20185,N_18335,N_18770);
xor U20186 (N_20186,N_19887,N_18241);
xnor U20187 (N_20187,N_18117,N_18899);
nand U20188 (N_20188,N_19992,N_19543);
nor U20189 (N_20189,N_18067,N_19073);
nor U20190 (N_20190,N_19739,N_19583);
nor U20191 (N_20191,N_19465,N_18490);
and U20192 (N_20192,N_18563,N_18514);
nand U20193 (N_20193,N_19601,N_18889);
and U20194 (N_20194,N_19694,N_19427);
or U20195 (N_20195,N_18742,N_19574);
or U20196 (N_20196,N_19599,N_18511);
xnor U20197 (N_20197,N_19787,N_19593);
or U20198 (N_20198,N_18773,N_18123);
nor U20199 (N_20199,N_18113,N_18878);
nand U20200 (N_20200,N_19184,N_18270);
xnor U20201 (N_20201,N_19319,N_18759);
and U20202 (N_20202,N_18288,N_18722);
and U20203 (N_20203,N_19057,N_19710);
nand U20204 (N_20204,N_18296,N_18181);
and U20205 (N_20205,N_19406,N_19899);
xor U20206 (N_20206,N_19067,N_18980);
nand U20207 (N_20207,N_18744,N_19345);
nor U20208 (N_20208,N_18199,N_18318);
and U20209 (N_20209,N_18684,N_19020);
nor U20210 (N_20210,N_19087,N_19242);
or U20211 (N_20211,N_19316,N_18551);
nor U20212 (N_20212,N_18954,N_19037);
and U20213 (N_20213,N_18669,N_18267);
or U20214 (N_20214,N_19860,N_18379);
nor U20215 (N_20215,N_19917,N_18624);
nor U20216 (N_20216,N_19307,N_19004);
nand U20217 (N_20217,N_19180,N_19046);
or U20218 (N_20218,N_19600,N_18302);
nand U20219 (N_20219,N_18046,N_19760);
nand U20220 (N_20220,N_19851,N_19471);
or U20221 (N_20221,N_18621,N_19498);
nor U20222 (N_20222,N_19015,N_18656);
and U20223 (N_20223,N_18786,N_19818);
nor U20224 (N_20224,N_19054,N_18170);
or U20225 (N_20225,N_19019,N_18186);
nand U20226 (N_20226,N_19025,N_18515);
nor U20227 (N_20227,N_18205,N_19482);
nor U20228 (N_20228,N_19671,N_18127);
nand U20229 (N_20229,N_18083,N_18299);
nor U20230 (N_20230,N_19281,N_18626);
nor U20231 (N_20231,N_18158,N_18234);
nor U20232 (N_20232,N_19150,N_19473);
and U20233 (N_20233,N_18587,N_19301);
or U20234 (N_20234,N_19220,N_18301);
nand U20235 (N_20235,N_19847,N_18560);
and U20236 (N_20236,N_19480,N_18888);
nor U20237 (N_20237,N_18754,N_19632);
nor U20238 (N_20238,N_19007,N_18943);
xnor U20239 (N_20239,N_19806,N_18860);
nand U20240 (N_20240,N_18421,N_18765);
nand U20241 (N_20241,N_18368,N_19940);
xnor U20242 (N_20242,N_18798,N_18854);
or U20243 (N_20243,N_19050,N_19536);
nand U20244 (N_20244,N_18891,N_18263);
nand U20245 (N_20245,N_19133,N_19805);
xor U20246 (N_20246,N_19497,N_19164);
nor U20247 (N_20247,N_19200,N_19643);
and U20248 (N_20248,N_19793,N_18163);
nand U20249 (N_20249,N_19604,N_18362);
or U20250 (N_20250,N_19843,N_19396);
nand U20251 (N_20251,N_19222,N_19931);
and U20252 (N_20252,N_19644,N_19709);
or U20253 (N_20253,N_19895,N_19853);
nor U20254 (N_20254,N_18242,N_18244);
and U20255 (N_20255,N_18917,N_18005);
or U20256 (N_20256,N_18209,N_19609);
nand U20257 (N_20257,N_19796,N_19827);
xor U20258 (N_20258,N_19420,N_18255);
or U20259 (N_20259,N_18295,N_18970);
nor U20260 (N_20260,N_19989,N_19371);
nor U20261 (N_20261,N_19144,N_18528);
and U20262 (N_20262,N_18274,N_19364);
or U20263 (N_20263,N_18737,N_19929);
and U20264 (N_20264,N_19238,N_18256);
nor U20265 (N_20265,N_19249,N_19504);
nor U20266 (N_20266,N_19979,N_19637);
nor U20267 (N_20267,N_19663,N_19789);
nand U20268 (N_20268,N_19898,N_19492);
xnor U20269 (N_20269,N_18651,N_19424);
nor U20270 (N_20270,N_19085,N_18197);
xnor U20271 (N_20271,N_19660,N_19062);
or U20272 (N_20272,N_19434,N_18032);
nor U20273 (N_20273,N_19039,N_18182);
and U20274 (N_20274,N_19556,N_19438);
xnor U20275 (N_20275,N_18369,N_19933);
or U20276 (N_20276,N_19283,N_18842);
xor U20277 (N_20277,N_19837,N_18636);
and U20278 (N_20278,N_19575,N_19864);
xnor U20279 (N_20279,N_18512,N_18513);
and U20280 (N_20280,N_19733,N_18827);
or U20281 (N_20281,N_18114,N_19157);
nor U20282 (N_20282,N_18315,N_19303);
nand U20283 (N_20283,N_18559,N_19194);
nor U20284 (N_20284,N_18457,N_19590);
and U20285 (N_20285,N_19361,N_19437);
and U20286 (N_20286,N_18779,N_18706);
xnor U20287 (N_20287,N_19693,N_18533);
nand U20288 (N_20288,N_18131,N_19676);
nor U20289 (N_20289,N_18532,N_19859);
nand U20290 (N_20290,N_18304,N_18972);
and U20291 (N_20291,N_18895,N_19735);
nand U20292 (N_20292,N_18974,N_18990);
or U20293 (N_20293,N_18771,N_19680);
nor U20294 (N_20294,N_18026,N_19585);
xnor U20295 (N_20295,N_19928,N_18576);
or U20296 (N_20296,N_19415,N_18709);
and U20297 (N_20297,N_18703,N_19872);
nor U20298 (N_20298,N_18053,N_19082);
nand U20299 (N_20299,N_18237,N_18671);
xnor U20300 (N_20300,N_19113,N_19755);
nand U20301 (N_20301,N_19513,N_18193);
or U20302 (N_20302,N_18912,N_19586);
nand U20303 (N_20303,N_18584,N_19125);
xor U20304 (N_20304,N_18585,N_19552);
and U20305 (N_20305,N_19926,N_19230);
nor U20306 (N_20306,N_18687,N_19791);
nor U20307 (N_20307,N_19948,N_18134);
nand U20308 (N_20308,N_19698,N_19731);
nor U20309 (N_20309,N_18942,N_19289);
xor U20310 (N_20310,N_18406,N_19469);
nand U20311 (N_20311,N_18824,N_18235);
xor U20312 (N_20312,N_18428,N_18142);
or U20313 (N_20313,N_19723,N_18538);
xor U20314 (N_20314,N_19232,N_18994);
and U20315 (N_20315,N_19654,N_18333);
and U20316 (N_20316,N_18166,N_19626);
nor U20317 (N_20317,N_18122,N_18171);
nand U20318 (N_20318,N_18968,N_18844);
nor U20319 (N_20319,N_18820,N_18178);
nand U20320 (N_20320,N_18985,N_18543);
xor U20321 (N_20321,N_19151,N_18996);
nor U20322 (N_20322,N_18349,N_19196);
xor U20323 (N_20323,N_19711,N_18988);
nand U20324 (N_20324,N_19811,N_19769);
nand U20325 (N_20325,N_19126,N_19865);
or U20326 (N_20326,N_19093,N_18057);
xnor U20327 (N_20327,N_19285,N_19348);
nor U20328 (N_20328,N_18861,N_19029);
nor U20329 (N_20329,N_18008,N_18958);
xnor U20330 (N_20330,N_18139,N_19474);
xor U20331 (N_20331,N_18366,N_19535);
or U20332 (N_20332,N_18089,N_18604);
xor U20333 (N_20333,N_18568,N_19496);
or U20334 (N_20334,N_18575,N_18577);
nand U20335 (N_20335,N_19627,N_19106);
nor U20336 (N_20336,N_19237,N_18869);
or U20337 (N_20337,N_18012,N_18518);
and U20338 (N_20338,N_19166,N_18419);
nor U20339 (N_20339,N_18680,N_19565);
xnor U20340 (N_20340,N_19068,N_18293);
nor U20341 (N_20341,N_19901,N_19870);
nor U20342 (N_20342,N_18910,N_18386);
nand U20343 (N_20343,N_19422,N_19185);
nand U20344 (N_20344,N_18298,N_19075);
nand U20345 (N_20345,N_19692,N_18572);
and U20346 (N_20346,N_19897,N_19146);
or U20347 (N_20347,N_18810,N_19642);
xor U20348 (N_20348,N_19193,N_18351);
and U20349 (N_20349,N_18945,N_19109);
and U20350 (N_20350,N_18323,N_19191);
or U20351 (N_20351,N_19296,N_18115);
nand U20352 (N_20352,N_18251,N_19987);
and U20353 (N_20353,N_19656,N_18360);
and U20354 (N_20354,N_18763,N_19786);
and U20355 (N_20355,N_19538,N_18717);
and U20356 (N_20356,N_19580,N_18477);
xnor U20357 (N_20357,N_19170,N_18220);
nor U20358 (N_20358,N_18811,N_18445);
or U20359 (N_20359,N_18258,N_18177);
nor U20360 (N_20360,N_19276,N_18120);
xor U20361 (N_20361,N_18885,N_18690);
and U20362 (N_20362,N_19129,N_18662);
or U20363 (N_20363,N_19975,N_19325);
nor U20364 (N_20364,N_19508,N_19697);
and U20365 (N_20365,N_18726,N_18682);
and U20366 (N_20366,N_19631,N_18007);
or U20367 (N_20367,N_19069,N_19401);
xnor U20368 (N_20368,N_18618,N_19573);
or U20369 (N_20369,N_18075,N_19089);
or U20370 (N_20370,N_19336,N_18794);
nand U20371 (N_20371,N_18705,N_18000);
and U20372 (N_20372,N_19963,N_19780);
nand U20373 (N_20373,N_19824,N_19219);
and U20374 (N_20374,N_18452,N_19812);
nand U20375 (N_20375,N_19691,N_19835);
nor U20376 (N_20376,N_19460,N_18002);
nand U20377 (N_20377,N_18056,N_18865);
nand U20378 (N_20378,N_19331,N_18321);
or U20379 (N_20379,N_18024,N_19629);
or U20380 (N_20380,N_19155,N_18107);
nor U20381 (N_20381,N_18347,N_19302);
xnor U20382 (N_20382,N_19169,N_18156);
or U20383 (N_20383,N_18087,N_19433);
nand U20384 (N_20384,N_19112,N_18344);
nor U20385 (N_20385,N_18268,N_18495);
or U20386 (N_20386,N_19138,N_18890);
or U20387 (N_20387,N_18161,N_19708);
or U20388 (N_20388,N_19909,N_19628);
or U20389 (N_20389,N_19470,N_18725);
nand U20390 (N_20390,N_19412,N_19746);
xor U20391 (N_20391,N_18948,N_18781);
nor U20392 (N_20392,N_18524,N_18433);
nand U20393 (N_20393,N_19000,N_19056);
and U20394 (N_20394,N_19053,N_18035);
and U20395 (N_20395,N_19322,N_19273);
or U20396 (N_20396,N_19688,N_19202);
and U20397 (N_20397,N_18090,N_19044);
nand U20398 (N_20398,N_19502,N_18357);
nor U20399 (N_20399,N_19955,N_19058);
nor U20400 (N_20400,N_19619,N_19758);
nor U20401 (N_20401,N_18739,N_18531);
or U20402 (N_20402,N_18649,N_18327);
or U20403 (N_20403,N_19675,N_18923);
nor U20404 (N_20404,N_18176,N_18544);
xnor U20405 (N_20405,N_19922,N_19744);
xor U20406 (N_20406,N_19313,N_19996);
nand U20407 (N_20407,N_18654,N_19333);
nand U20408 (N_20408,N_19179,N_18201);
xor U20409 (N_20409,N_18487,N_19696);
xor U20410 (N_20410,N_18044,N_19968);
and U20411 (N_20411,N_18908,N_19403);
nand U20412 (N_20412,N_18783,N_18042);
xor U20413 (N_20413,N_18196,N_19274);
nand U20414 (N_20414,N_18561,N_18461);
and U20415 (N_20415,N_18033,N_18020);
and U20416 (N_20416,N_18588,N_18373);
or U20417 (N_20417,N_19423,N_19409);
nor U20418 (N_20418,N_18305,N_18069);
nor U20419 (N_20419,N_19459,N_19108);
or U20420 (N_20420,N_19500,N_19799);
nand U20421 (N_20421,N_19461,N_19558);
xor U20422 (N_20422,N_19547,N_19653);
nand U20423 (N_20423,N_18486,N_18378);
xor U20424 (N_20424,N_18932,N_18821);
and U20425 (N_20425,N_18745,N_18802);
or U20426 (N_20426,N_19177,N_19041);
and U20427 (N_20427,N_19435,N_18834);
xor U20428 (N_20428,N_18025,N_19367);
or U20429 (N_20429,N_18192,N_19519);
or U20430 (N_20430,N_18935,N_18482);
nor U20431 (N_20431,N_18372,N_18363);
nor U20432 (N_20432,N_18813,N_19750);
or U20433 (N_20433,N_18825,N_18396);
and U20434 (N_20434,N_18689,N_18975);
or U20435 (N_20435,N_19706,N_18125);
nand U20436 (N_20436,N_18901,N_18805);
nor U20437 (N_20437,N_19612,N_19749);
xor U20438 (N_20438,N_18925,N_19205);
xor U20439 (N_20439,N_19291,N_18855);
xor U20440 (N_20440,N_19712,N_18835);
nand U20441 (N_20441,N_19732,N_19820);
or U20442 (N_20442,N_18485,N_18555);
nor U20443 (N_20443,N_18874,N_19130);
nand U20444 (N_20444,N_19974,N_18052);
nand U20445 (N_20445,N_19338,N_19822);
and U20446 (N_20446,N_19293,N_19634);
and U20447 (N_20447,N_19472,N_19766);
nor U20448 (N_20448,N_18006,N_18469);
or U20449 (N_20449,N_19576,N_18157);
and U20450 (N_20450,N_18876,N_18449);
and U20451 (N_20451,N_19702,N_19043);
and U20452 (N_20452,N_19893,N_19534);
nand U20453 (N_20453,N_18198,N_19509);
or U20454 (N_20454,N_19008,N_19807);
or U20455 (N_20455,N_18207,N_18535);
and U20456 (N_20456,N_19879,N_19374);
and U20457 (N_20457,N_18308,N_19553);
and U20458 (N_20458,N_19201,N_19505);
and U20459 (N_20459,N_19114,N_18309);
or U20460 (N_20460,N_18583,N_19834);
or U20461 (N_20461,N_19347,N_19515);
xor U20462 (N_20462,N_18329,N_19055);
and U20463 (N_20463,N_19458,N_18546);
and U20464 (N_20464,N_18539,N_18135);
and U20465 (N_20465,N_18731,N_19862);
or U20466 (N_20466,N_19248,N_18010);
nand U20467 (N_20467,N_19097,N_19686);
or U20468 (N_20468,N_18306,N_18879);
and U20469 (N_20469,N_19259,N_19421);
nor U20470 (N_20470,N_19956,N_19639);
or U20471 (N_20471,N_18909,N_18982);
and U20472 (N_20472,N_19959,N_18119);
and U20473 (N_20473,N_19141,N_18212);
xnor U20474 (N_20474,N_19550,N_19823);
nand U20475 (N_20475,N_19803,N_19532);
nor U20476 (N_20476,N_19771,N_18553);
and U20477 (N_20477,N_19375,N_19905);
nor U20478 (N_20478,N_18516,N_18635);
or U20479 (N_20479,N_19399,N_18679);
nor U20480 (N_20480,N_18247,N_18222);
nor U20481 (N_20481,N_18565,N_19171);
or U20482 (N_20482,N_19183,N_18830);
nand U20483 (N_20483,N_18143,N_18494);
xnor U20484 (N_20484,N_19685,N_19306);
and U20485 (N_20485,N_18420,N_19326);
or U20486 (N_20486,N_18858,N_19236);
xnor U20487 (N_20487,N_18831,N_19650);
xor U20488 (N_20488,N_19883,N_18022);
nand U20489 (N_20489,N_18517,N_18601);
nor U20490 (N_20490,N_19450,N_19045);
xnor U20491 (N_20491,N_19721,N_19393);
and U20492 (N_20492,N_18598,N_19337);
nor U20493 (N_20493,N_19418,N_18856);
nor U20494 (N_20494,N_18132,N_18733);
nor U20495 (N_20495,N_19630,N_19608);
and U20496 (N_20496,N_18497,N_19833);
xor U20497 (N_20497,N_19873,N_18808);
and U20498 (N_20498,N_18659,N_18392);
or U20499 (N_20499,N_18337,N_18791);
xor U20500 (N_20500,N_18594,N_18838);
or U20501 (N_20501,N_19520,N_19491);
nor U20502 (N_20502,N_18937,N_19373);
or U20503 (N_20503,N_19327,N_18833);
nand U20504 (N_20504,N_18278,N_19379);
nand U20505 (N_20505,N_19914,N_18229);
xor U20506 (N_20506,N_19405,N_18780);
or U20507 (N_20507,N_19617,N_19241);
nand U20508 (N_20508,N_18836,N_19388);
xor U20509 (N_20509,N_19455,N_18072);
nor U20510 (N_20510,N_19939,N_19954);
nand U20511 (N_20511,N_19410,N_19064);
or U20512 (N_20512,N_19571,N_18422);
xnor U20513 (N_20513,N_19953,N_18960);
and U20514 (N_20514,N_18806,N_19625);
and U20515 (N_20515,N_18340,N_18853);
or U20516 (N_20516,N_19195,N_18611);
and U20517 (N_20517,N_19778,N_19269);
nand U20518 (N_20518,N_18617,N_19635);
nand U20519 (N_20519,N_18466,N_18582);
nor U20520 (N_20520,N_18050,N_19175);
and U20521 (N_20521,N_18950,N_19620);
nor U20522 (N_20522,N_18969,N_19924);
and U20523 (N_20523,N_18124,N_19121);
nand U20524 (N_20524,N_18695,N_18736);
nand U20525 (N_20525,N_19976,N_19324);
and U20526 (N_20526,N_19557,N_19920);
xor U20527 (N_20527,N_18381,N_19980);
nand U20528 (N_20528,N_19042,N_19264);
or U20529 (N_20529,N_18882,N_18723);
nor U20530 (N_20530,N_19741,N_19541);
xor U20531 (N_20531,N_18663,N_19781);
or U20532 (N_20532,N_19060,N_18254);
nor U20533 (N_20533,N_18259,N_18167);
and U20534 (N_20534,N_18478,N_19658);
nand U20535 (N_20535,N_18631,N_19904);
nand U20536 (N_20536,N_18448,N_19312);
nand U20537 (N_20537,N_18014,N_19209);
xor U20538 (N_20538,N_19079,N_18442);
xor U20539 (N_20539,N_19448,N_18738);
xor U20540 (N_20540,N_18377,N_18265);
nor U20541 (N_20541,N_19757,N_19266);
or U20542 (N_20542,N_18231,N_19478);
nand U20543 (N_20543,N_18992,N_18732);
xor U20544 (N_20544,N_19123,N_19751);
nor U20545 (N_20545,N_19869,N_19849);
and U20546 (N_20546,N_19664,N_19577);
nor U20547 (N_20547,N_19318,N_18375);
nor U20548 (N_20548,N_19288,N_19092);
nor U20549 (N_20549,N_18160,N_18708);
nor U20550 (N_20550,N_19669,N_19896);
and U20551 (N_20551,N_19119,N_18221);
or U20552 (N_20552,N_19483,N_19906);
or U20553 (N_20553,N_18374,N_18210);
nand U20554 (N_20554,N_18841,N_18307);
and U20555 (N_20555,N_19969,N_18048);
xnor U20556 (N_20556,N_19178,N_18294);
nor U20557 (N_20557,N_19408,N_18525);
nor U20558 (N_20558,N_18873,N_18355);
nor U20559 (N_20559,N_19611,N_19485);
or U20560 (N_20560,N_18184,N_19759);
xor U20561 (N_20561,N_18564,N_18547);
and U20562 (N_20562,N_18211,N_19083);
nand U20563 (N_20563,N_19001,N_18676);
nor U20564 (N_20564,N_18571,N_18877);
or U20565 (N_20565,N_18146,N_19982);
xnor U20566 (N_20566,N_19564,N_19103);
xor U20567 (N_20567,N_19528,N_18911);
and U20568 (N_20568,N_19900,N_19429);
or U20569 (N_20569,N_19231,N_18864);
and U20570 (N_20570,N_18589,N_18149);
nand U20571 (N_20571,N_18317,N_18927);
or U20572 (N_20572,N_19463,N_19095);
and U20573 (N_20573,N_19884,N_19311);
nand U20574 (N_20574,N_18350,N_18758);
xnor U20575 (N_20575,N_18467,N_18862);
or U20576 (N_20576,N_18346,N_19386);
or U20577 (N_20577,N_19439,N_19070);
or U20578 (N_20578,N_19810,N_19501);
xnor U20579 (N_20579,N_18929,N_19670);
or U20580 (N_20580,N_19584,N_18541);
or U20581 (N_20581,N_18951,N_19464);
or U20582 (N_20582,N_19490,N_19187);
nor U20583 (N_20583,N_18264,N_18578);
or U20584 (N_20584,N_19445,N_18920);
nor U20585 (N_20585,N_19544,N_18353);
nand U20586 (N_20586,N_19809,N_18314);
and U20587 (N_20587,N_19365,N_18957);
nand U20588 (N_20588,N_18787,N_19678);
nand U20589 (N_20589,N_18913,N_18130);
nor U20590 (N_20590,N_18216,N_18154);
nand U20591 (N_20591,N_18956,N_18790);
nand U20592 (N_20592,N_18061,N_18697);
or U20593 (N_20593,N_19304,N_19765);
nand U20594 (N_20594,N_18857,N_19263);
nor U20595 (N_20595,N_19099,N_19131);
or U20596 (N_20596,N_19494,N_19800);
and U20597 (N_20597,N_18622,N_18886);
and U20598 (N_20598,N_18194,N_19866);
or U20599 (N_20599,N_19546,N_19867);
xor U20600 (N_20600,N_18832,N_18088);
or U20601 (N_20601,N_19134,N_18595);
and U20602 (N_20602,N_18987,N_19936);
xnor U20603 (N_20603,N_18253,N_19287);
nor U20604 (N_20604,N_18489,N_19912);
and U20605 (N_20605,N_18693,N_19852);
xor U20606 (N_20606,N_18148,N_19944);
nor U20607 (N_20607,N_18976,N_18055);
nor U20608 (N_20608,N_18718,N_18724);
nor U20609 (N_20609,N_19923,N_19407);
nand U20610 (N_20610,N_19623,N_18459);
nand U20611 (N_20611,N_18789,N_18675);
nor U20612 (N_20612,N_19199,N_18973);
nand U20613 (N_20613,N_19495,N_18715);
or U20614 (N_20614,N_18408,N_19764);
or U20615 (N_20615,N_18884,N_19941);
and U20616 (N_20616,N_18933,N_18286);
and U20617 (N_20617,N_19212,N_19074);
xor U20618 (N_20618,N_19310,N_18750);
nand U20619 (N_20619,N_18017,N_19950);
nand U20620 (N_20620,N_19137,N_19829);
xnor U20621 (N_20621,N_19548,N_18215);
nand U20622 (N_20622,N_18279,N_19111);
and U20623 (N_20623,N_18632,N_18756);
nand U20624 (N_20624,N_18907,N_19512);
or U20625 (N_20625,N_19385,N_19034);
xnor U20626 (N_20626,N_18735,N_19804);
xor U20627 (N_20627,N_19946,N_18871);
nor U20628 (N_20628,N_18454,N_18613);
nand U20629 (N_20629,N_18894,N_18761);
nand U20630 (N_20630,N_19261,N_18423);
xor U20631 (N_20631,N_18610,N_18848);
nor U20632 (N_20632,N_18557,N_18376);
or U20633 (N_20633,N_19286,N_19581);
or U20634 (N_20634,N_19088,N_19844);
nand U20635 (N_20635,N_18971,N_19275);
nand U20636 (N_20636,N_18185,N_18230);
nor U20637 (N_20637,N_18607,N_18365);
or U20638 (N_20638,N_18764,N_19321);
xor U20639 (N_20639,N_18030,N_19462);
nand U20640 (N_20640,N_18438,N_18788);
or U20641 (N_20641,N_19911,N_18814);
xnor U20642 (N_20642,N_18646,N_18141);
and U20643 (N_20643,N_18108,N_18085);
nor U20644 (N_20644,N_18608,N_19239);
or U20645 (N_20645,N_19748,N_18508);
and U20646 (N_20646,N_18261,N_18628);
nand U20647 (N_20647,N_18402,N_18126);
xnor U20648 (N_20648,N_19446,N_19831);
nor U20649 (N_20649,N_19591,N_18615);
and U20650 (N_20650,N_18206,N_18491);
and U20651 (N_20651,N_19279,N_19908);
xor U20652 (N_20652,N_19211,N_19389);
and U20653 (N_20653,N_19271,N_18850);
and U20654 (N_20654,N_18979,N_18291);
or U20655 (N_20655,N_19078,N_19588);
and U20656 (N_20656,N_19986,N_19467);
xnor U20657 (N_20657,N_19431,N_19390);
or U20658 (N_20658,N_19567,N_19842);
xor U20659 (N_20659,N_18248,N_18768);
xnor U20660 (N_20660,N_18924,N_18415);
nand U20661 (N_20661,N_19278,N_18606);
nor U20662 (N_20662,N_19003,N_18104);
nand U20663 (N_20663,N_19489,N_18473);
nand U20664 (N_20664,N_19270,N_19244);
and U20665 (N_20665,N_18602,N_18743);
xnor U20666 (N_20666,N_19493,N_18354);
or U20667 (N_20667,N_18481,N_18666);
or U20668 (N_20668,N_19207,N_18311);
nor U20669 (N_20669,N_18128,N_18875);
or U20670 (N_20670,N_19882,N_19309);
and U20671 (N_20671,N_19100,N_18434);
nand U20672 (N_20672,N_19094,N_19299);
nor U20673 (N_20673,N_19186,N_18699);
xnor U20674 (N_20674,N_18418,N_19672);
nor U20675 (N_20675,N_18946,N_19376);
nor U20676 (N_20676,N_18064,N_19995);
xnor U20677 (N_20677,N_18001,N_19256);
xnor U20678 (N_20678,N_18059,N_19063);
xnor U20679 (N_20679,N_19782,N_19526);
nand U20680 (N_20680,N_18472,N_19443);
nor U20681 (N_20681,N_19719,N_18550);
nor U20682 (N_20682,N_18905,N_18118);
and U20683 (N_20683,N_19845,N_19894);
xnor U20684 (N_20684,N_19943,N_19091);
nor U20685 (N_20685,N_18147,N_18371);
xnor U20686 (N_20686,N_19254,N_18634);
xnor U20687 (N_20687,N_19216,N_18179);
or U20688 (N_20688,N_19369,N_19340);
and U20689 (N_20689,N_18784,N_18018);
and U20690 (N_20690,N_18661,N_18529);
nor U20691 (N_20691,N_19682,N_18991);
and U20692 (N_20692,N_19210,N_18441);
nand U20693 (N_20693,N_18410,N_18039);
and U20694 (N_20694,N_18549,N_19700);
and U20695 (N_20695,N_18506,N_18208);
nor U20696 (N_20696,N_18407,N_19233);
or U20697 (N_20697,N_18782,N_18100);
and U20698 (N_20698,N_19880,N_18271);
nand U20699 (N_20699,N_19622,N_19456);
nor U20700 (N_20700,N_18080,N_19167);
xor U20701 (N_20701,N_19018,N_18439);
or U20702 (N_20702,N_19351,N_19952);
nor U20703 (N_20703,N_19525,N_19891);
xnor U20704 (N_20704,N_19918,N_19618);
and U20705 (N_20705,N_19876,N_18592);
and U20706 (N_20706,N_19487,N_18073);
xor U20707 (N_20707,N_18799,N_19774);
xnor U20708 (N_20708,N_18719,N_18456);
nor U20709 (N_20709,N_19913,N_19048);
nand U20710 (N_20710,N_19284,N_18900);
and U20711 (N_20711,N_19915,N_19032);
or U20712 (N_20712,N_18720,N_19846);
xor U20713 (N_20713,N_18047,N_19615);
xnor U20714 (N_20714,N_18312,N_18846);
xor U20715 (N_20715,N_19038,N_19208);
or U20716 (N_20716,N_18150,N_18272);
and U20717 (N_20717,N_19265,N_19542);
xnor U20718 (N_20718,N_18966,N_19713);
nand U20719 (N_20719,N_19215,N_18011);
or U20720 (N_20720,N_19839,N_19395);
nor U20721 (N_20721,N_19192,N_19734);
nor U20722 (N_20722,N_19540,N_18172);
or U20723 (N_20723,N_19792,N_18633);
and U20724 (N_20724,N_18266,N_18961);
or U20725 (N_20725,N_19661,N_19440);
xor U20726 (N_20726,N_18203,N_18803);
nand U20727 (N_20727,N_18455,N_18310);
nand U20728 (N_20728,N_19790,N_19383);
nand U20729 (N_20729,N_19503,N_19736);
nand U20730 (N_20730,N_18609,N_19850);
nor U20731 (N_20731,N_19428,N_18521);
or U20732 (N_20732,N_18746,N_19984);
nor U20733 (N_20733,N_18152,N_18173);
and U20734 (N_20734,N_19223,N_19925);
xnor U20735 (N_20735,N_19659,N_19747);
nor U20736 (N_20736,N_19086,N_18183);
or U20737 (N_20737,N_18389,N_19128);
and U20738 (N_20738,N_18605,N_19084);
xnor U20739 (N_20739,N_18367,N_18189);
xnor U20740 (N_20740,N_18105,N_19551);
xnor U20741 (N_20741,N_18897,N_18498);
or U20742 (N_20742,N_19394,N_18313);
nor U20743 (N_20743,N_18462,N_18944);
nand U20744 (N_20744,N_19517,N_19649);
nor U20745 (N_20745,N_19647,N_19339);
or U20746 (N_20746,N_18616,N_19189);
nand U20747 (N_20747,N_19808,N_19705);
or U20748 (N_20748,N_18527,N_18474);
nor U20749 (N_20749,N_19161,N_18597);
nor U20750 (N_20750,N_18393,N_18591);
xnor U20751 (N_20751,N_18336,N_19381);
xnor U20752 (N_20752,N_19168,N_18095);
xnor U20753 (N_20753,N_19689,N_18881);
nand U20754 (N_20754,N_19182,N_18870);
nand U20755 (N_20755,N_19257,N_18545);
or U20756 (N_20756,N_19756,N_19342);
nor U20757 (N_20757,N_19240,N_19272);
or U20758 (N_20758,N_19252,N_18435);
or U20759 (N_20759,N_18070,N_18767);
nor U20760 (N_20760,N_19300,N_18165);
and U20761 (N_20761,N_18330,N_19638);
xnor U20762 (N_20762,N_19971,N_18769);
and U20763 (N_20763,N_19874,N_19118);
or U20764 (N_20764,N_18348,N_19991);
xnor U20765 (N_20765,N_19776,N_19059);
xnor U20766 (N_20766,N_19005,N_19683);
xnor U20767 (N_20767,N_18405,N_18027);
or U20768 (N_20768,N_18711,N_19794);
nand U20769 (N_20769,N_18859,N_19554);
and U20770 (N_20770,N_18849,N_18076);
nand U20771 (N_20771,N_19143,N_18496);
nor U20772 (N_20772,N_19726,N_19320);
xnor U20773 (N_20773,N_18190,N_18619);
nor U20774 (N_20774,N_19707,N_19566);
and U20775 (N_20775,N_19416,N_18984);
xnor U20776 (N_20776,N_18038,N_18260);
xor U20777 (N_20777,N_18751,N_18526);
or U20778 (N_20778,N_19136,N_19754);
nor U20779 (N_20779,N_19919,N_19614);
nor U20780 (N_20780,N_19973,N_19172);
and U20781 (N_20781,N_18345,N_18282);
or U20782 (N_20782,N_18573,N_19398);
nor U20783 (N_20783,N_19021,N_19012);
xnor U20784 (N_20784,N_18417,N_18476);
nand U20785 (N_20785,N_18685,N_19466);
nand U20786 (N_20786,N_18303,N_18648);
nand U20787 (N_20787,N_19268,N_18065);
nand U20788 (N_20788,N_18110,N_19767);
nor U20789 (N_20789,N_18425,N_18536);
nor U20790 (N_20790,N_19414,N_19716);
xor U20791 (N_20791,N_18537,N_18437);
nand U20792 (N_20792,N_18387,N_18729);
xor U20793 (N_20793,N_18383,N_19730);
nor U20794 (N_20794,N_18638,N_19798);
or U20795 (N_20795,N_18257,N_19317);
and U20796 (N_20796,N_18426,N_18530);
and U20797 (N_20797,N_19013,N_19444);
and U20798 (N_20798,N_18644,N_19165);
or U20799 (N_20799,N_19949,N_18941);
or U20800 (N_20800,N_18227,N_18556);
or U20801 (N_20801,N_19562,N_18914);
xor U20802 (N_20802,N_19522,N_19582);
and U20803 (N_20803,N_18712,N_19297);
nor U20804 (N_20804,N_19673,N_19049);
xor U20805 (N_20805,N_18403,N_18678);
and U20806 (N_20806,N_18938,N_19499);
xor U20807 (N_20807,N_18331,N_19636);
nand U20808 (N_20808,N_19568,N_18775);
and U20809 (N_20809,N_18716,N_19938);
xnor U20810 (N_20810,N_18015,N_19655);
and U20811 (N_20811,N_19115,N_19830);
and U20812 (N_20812,N_18174,N_19217);
nand U20813 (N_20813,N_18342,N_19819);
nand U20814 (N_20814,N_19813,N_19282);
or U20815 (N_20815,N_18620,N_19392);
and U20816 (N_20816,N_19606,N_18411);
or U20817 (N_20817,N_18019,N_18213);
xor U20818 (N_20818,N_19080,N_19768);
and U20819 (N_20819,N_19855,N_18364);
and U20820 (N_20820,N_19945,N_19961);
or U20821 (N_20821,N_18872,N_18168);
or U20822 (N_20822,N_18757,N_18847);
nor U20823 (N_20823,N_19350,N_18140);
and U20824 (N_20824,N_19903,N_19621);
and U20825 (N_20825,N_18698,N_18320);
and U20826 (N_20826,N_18034,N_19323);
nor U20827 (N_20827,N_18774,N_18936);
nand U20828 (N_20828,N_19964,N_19530);
xor U20829 (N_20829,N_18424,N_18962);
or U20830 (N_20830,N_18062,N_19902);
nor U20831 (N_20831,N_18683,N_19978);
nor U20832 (N_20832,N_18839,N_19028);
nor U20833 (N_20833,N_18464,N_18674);
xnor U20834 (N_20834,N_18153,N_19449);
and U20835 (N_20835,N_19158,N_18384);
or U20836 (N_20836,N_19539,N_18285);
xnor U20837 (N_20837,N_19356,N_18677);
nand U20838 (N_20838,N_19990,N_18204);
xnor U20839 (N_20839,N_18356,N_19468);
xor U20840 (N_20840,N_18792,N_18999);
nor U20841 (N_20841,N_19545,N_19334);
nor U20842 (N_20842,N_18280,N_19251);
or U20843 (N_20843,N_19481,N_19640);
and U20844 (N_20844,N_19788,N_18101);
nor U20845 (N_20845,N_19344,N_18281);
nor U20846 (N_20846,N_19665,N_19932);
and U20847 (N_20847,N_19246,N_18084);
or U20848 (N_20848,N_18567,N_18641);
xnor U20849 (N_20849,N_18748,N_18430);
nand U20850 (N_20850,N_19419,N_19595);
or U20851 (N_20851,N_19292,N_19832);
xnor U20852 (N_20852,N_18694,N_18471);
or U20853 (N_20853,N_19314,N_18590);
and U20854 (N_20854,N_18600,N_18099);
and U20855 (N_20855,N_19816,N_18728);
or U20856 (N_20856,N_18967,N_19892);
xnor U20857 (N_20857,N_18068,N_18358);
xnor U20858 (N_20858,N_18691,N_18045);
nor U20859 (N_20859,N_19815,N_19362);
xor U20860 (N_20860,N_18800,N_18390);
and U20861 (N_20861,N_18931,N_19475);
xor U20862 (N_20862,N_18200,N_19937);
nand U20863 (N_20863,N_18273,N_19605);
nor U20864 (N_20864,N_18137,N_18028);
xnor U20865 (N_20865,N_18652,N_19457);
nor U20866 (N_20866,N_19594,N_19772);
xor U20867 (N_20867,N_19052,N_19718);
or U20868 (N_20868,N_18388,N_18840);
and U20869 (N_20869,N_18159,N_19378);
nor U20870 (N_20870,N_18843,N_19354);
and U20871 (N_20871,N_19206,N_19529);
nand U20872 (N_20872,N_18510,N_18233);
xnor U20873 (N_20873,N_18238,N_19002);
and U20874 (N_20874,N_19335,N_18569);
xnor U20875 (N_20875,N_18892,N_18612);
nor U20876 (N_20876,N_18866,N_19570);
xor U20877 (N_20877,N_19934,N_18902);
or U20878 (N_20878,N_19531,N_18965);
nor U20879 (N_20879,N_19725,N_19555);
and U20880 (N_20880,N_19174,N_18218);
xnor U20881 (N_20881,N_18642,N_19890);
nand U20882 (N_20882,N_18240,N_18499);
nor U20883 (N_20883,N_18155,N_19359);
or U20884 (N_20884,N_18752,N_19360);
or U20885 (N_20885,N_19592,N_18507);
and U20886 (N_20886,N_18436,N_19977);
and U20887 (N_20887,N_19695,N_18401);
and U20888 (N_20888,N_19549,N_18554);
and U20889 (N_20889,N_18826,N_18776);
or U20890 (N_20890,N_18483,N_19479);
nand U20891 (N_20891,N_18041,N_19096);
xnor U20892 (N_20892,N_19380,N_19763);
nor U20893 (N_20893,N_18300,N_19224);
or U20894 (N_20894,N_19753,N_18829);
xnor U20895 (N_20895,N_18647,N_18955);
nand U20896 (N_20896,N_19484,N_18772);
nor U20897 (N_20897,N_18187,N_19863);
and U20898 (N_20898,N_19332,N_19743);
xor U20899 (N_20899,N_18043,N_19355);
nand U20900 (N_20900,N_19402,N_18998);
nand U20901 (N_20901,N_18239,N_18637);
nor U20902 (N_20902,N_18727,N_19596);
nand U20903 (N_20903,N_19247,N_19885);
xnor U20904 (N_20904,N_19061,N_18995);
nand U20905 (N_20905,N_19035,N_19667);
or U20906 (N_20906,N_19140,N_18804);
nor U20907 (N_20907,N_18522,N_19714);
nand U20908 (N_20908,N_18505,N_18029);
nand U20909 (N_20909,N_19341,N_19828);
xor U20910 (N_20910,N_19737,N_18681);
nand U20911 (N_20911,N_18749,N_18453);
nand U20912 (N_20912,N_18807,N_19127);
nand U20913 (N_20913,N_18664,N_19228);
xnor U20914 (N_20914,N_18981,N_18523);
nand U20915 (N_20915,N_19262,N_19988);
or U20916 (N_20916,N_19102,N_19777);
xnor U20917 (N_20917,N_18730,N_18450);
nand U20918 (N_20918,N_18922,N_18109);
nand U20919 (N_20919,N_18058,N_19065);
or U20920 (N_20920,N_18793,N_18243);
nor U20921 (N_20921,N_19027,N_19308);
xnor U20922 (N_20922,N_19197,N_18249);
nand U20923 (N_20923,N_18939,N_19927);
nor U20924 (N_20924,N_19857,N_19998);
nor U20925 (N_20925,N_18701,N_19298);
or U20926 (N_20926,N_19521,N_18232);
or U20927 (N_20927,N_19701,N_18650);
or U20928 (N_20928,N_19072,N_19295);
xnor U20929 (N_20929,N_18097,N_19762);
xor U20930 (N_20930,N_18816,N_19506);
and U20931 (N_20931,N_19840,N_18066);
nand U20932 (N_20932,N_18480,N_19527);
or U20933 (N_20933,N_19154,N_19426);
nor U20934 (N_20934,N_18016,N_19277);
or U20935 (N_20935,N_18082,N_19668);
xnor U20936 (N_20936,N_18352,N_18339);
nor U20937 (N_20937,N_19779,N_18603);
and U20938 (N_20938,N_18502,N_18246);
nor U20939 (N_20939,N_18116,N_18930);
and U20940 (N_20940,N_19728,N_19454);
nand U20941 (N_20941,N_18796,N_19516);
nor U20942 (N_20942,N_18625,N_19110);
nand U20943 (N_20943,N_19994,N_18380);
or U20944 (N_20944,N_19430,N_18096);
or U20945 (N_20945,N_18334,N_19149);
and U20946 (N_20946,N_18440,N_18283);
or U20947 (N_20947,N_19514,N_18202);
nor U20948 (N_20948,N_19921,N_19353);
nand U20949 (N_20949,N_18809,N_18906);
nor U20950 (N_20950,N_19132,N_19148);
nand U20951 (N_20951,N_19666,N_19122);
nand U20952 (N_20952,N_18760,N_18952);
and U20953 (N_20953,N_18822,N_18629);
and U20954 (N_20954,N_19510,N_18667);
nor U20955 (N_20955,N_18195,N_18921);
nand U20956 (N_20956,N_18823,N_19234);
xor U20957 (N_20957,N_19715,N_18755);
or U20958 (N_20958,N_18904,N_19699);
nor U20959 (N_20959,N_19981,N_19967);
and U20960 (N_20960,N_18250,N_18004);
nand U20961 (N_20961,N_19537,N_19413);
nand U20962 (N_20962,N_19250,N_18643);
and U20963 (N_20963,N_19090,N_19633);
and U20964 (N_20964,N_19153,N_18558);
or U20965 (N_20965,N_18704,N_18121);
xnor U20966 (N_20966,N_19400,N_19745);
nand U20967 (N_20967,N_19066,N_19598);
and U20968 (N_20968,N_19646,N_18953);
xnor U20969 (N_20969,N_18673,N_18228);
or U20970 (N_20970,N_18144,N_19328);
xnor U20971 (N_20971,N_18658,N_18063);
nand U20972 (N_20972,N_18928,N_19190);
or U20973 (N_20973,N_18868,N_18341);
or U20974 (N_20974,N_19253,N_18079);
or U20975 (N_20975,N_18887,N_19156);
nand U20976 (N_20976,N_18359,N_19613);
and U20977 (N_20977,N_18060,N_19524);
and U20978 (N_20978,N_18326,N_19645);
xor U20979 (N_20979,N_18398,N_18432);
or U20980 (N_20980,N_19107,N_19993);
nand U20981 (N_20981,N_18993,N_19752);
nor U20982 (N_20982,N_18828,N_19690);
xor U20983 (N_20983,N_18395,N_18940);
nand U20984 (N_20984,N_19357,N_19366);
nor U20985 (N_20985,N_19358,N_18581);
xnor U20986 (N_20986,N_18484,N_19511);
and U20987 (N_20987,N_18918,N_19773);
and U20988 (N_20988,N_19040,N_19886);
nor U20989 (N_20989,N_19011,N_18627);
xnor U20990 (N_20990,N_18446,N_18071);
nor U20991 (N_20991,N_19343,N_18700);
and U20992 (N_20992,N_19687,N_19363);
nand U20993 (N_20993,N_18040,N_19729);
or U20994 (N_20994,N_19717,N_19848);
and U20995 (N_20995,N_18343,N_19047);
nor U20996 (N_20996,N_19801,N_19377);
xor U20997 (N_20997,N_18145,N_18391);
and U20998 (N_20998,N_18883,N_18964);
xnor U20999 (N_20999,N_18081,N_18688);
nor U21000 (N_21000,N_19372,N_19896);
xnor U21001 (N_21001,N_18191,N_19057);
and U21002 (N_21002,N_19757,N_18990);
nor U21003 (N_21003,N_19895,N_19716);
xnor U21004 (N_21004,N_18031,N_18788);
nor U21005 (N_21005,N_19471,N_19170);
xnor U21006 (N_21006,N_18847,N_19611);
nand U21007 (N_21007,N_19241,N_19024);
nand U21008 (N_21008,N_19892,N_19218);
or U21009 (N_21009,N_18885,N_19729);
xnor U21010 (N_21010,N_19278,N_19931);
and U21011 (N_21011,N_19846,N_19183);
and U21012 (N_21012,N_19598,N_18654);
xnor U21013 (N_21013,N_19016,N_18525);
nand U21014 (N_21014,N_18036,N_19471);
nand U21015 (N_21015,N_19895,N_19745);
xor U21016 (N_21016,N_18040,N_18086);
nand U21017 (N_21017,N_18866,N_19125);
nor U21018 (N_21018,N_18503,N_19100);
xor U21019 (N_21019,N_18428,N_19825);
and U21020 (N_21020,N_18737,N_19175);
or U21021 (N_21021,N_19879,N_18630);
xor U21022 (N_21022,N_18643,N_19305);
nor U21023 (N_21023,N_18103,N_18713);
xnor U21024 (N_21024,N_18482,N_18051);
nor U21025 (N_21025,N_19254,N_18056);
and U21026 (N_21026,N_19277,N_18671);
and U21027 (N_21027,N_19752,N_18421);
and U21028 (N_21028,N_18458,N_19617);
nand U21029 (N_21029,N_18964,N_18935);
xnor U21030 (N_21030,N_19426,N_19632);
xor U21031 (N_21031,N_18244,N_18093);
nor U21032 (N_21032,N_18187,N_18536);
and U21033 (N_21033,N_19533,N_18945);
xor U21034 (N_21034,N_18998,N_19075);
nor U21035 (N_21035,N_18644,N_19814);
nor U21036 (N_21036,N_19590,N_18326);
nor U21037 (N_21037,N_19706,N_19115);
nand U21038 (N_21038,N_18062,N_18769);
and U21039 (N_21039,N_19080,N_19867);
and U21040 (N_21040,N_18560,N_19876);
or U21041 (N_21041,N_18765,N_18291);
or U21042 (N_21042,N_18195,N_19315);
nand U21043 (N_21043,N_18538,N_19939);
nand U21044 (N_21044,N_19026,N_18056);
nand U21045 (N_21045,N_19780,N_18215);
or U21046 (N_21046,N_19853,N_19130);
nor U21047 (N_21047,N_19677,N_19631);
nor U21048 (N_21048,N_18541,N_18424);
and U21049 (N_21049,N_19114,N_19673);
xor U21050 (N_21050,N_18868,N_18697);
nand U21051 (N_21051,N_18181,N_19399);
and U21052 (N_21052,N_18503,N_19697);
and U21053 (N_21053,N_18334,N_18686);
or U21054 (N_21054,N_19776,N_19655);
or U21055 (N_21055,N_19191,N_18359);
xnor U21056 (N_21056,N_19043,N_18470);
or U21057 (N_21057,N_19621,N_19963);
nor U21058 (N_21058,N_19438,N_18419);
or U21059 (N_21059,N_19865,N_18621);
and U21060 (N_21060,N_19601,N_19828);
nor U21061 (N_21061,N_19229,N_19382);
and U21062 (N_21062,N_18994,N_19341);
nand U21063 (N_21063,N_19728,N_18980);
nand U21064 (N_21064,N_19978,N_19209);
nand U21065 (N_21065,N_19668,N_18869);
nor U21066 (N_21066,N_19748,N_19242);
nor U21067 (N_21067,N_19749,N_18842);
nand U21068 (N_21068,N_19202,N_19850);
nor U21069 (N_21069,N_18749,N_19153);
or U21070 (N_21070,N_19610,N_19188);
xnor U21071 (N_21071,N_19670,N_18875);
nor U21072 (N_21072,N_18304,N_18392);
nand U21073 (N_21073,N_18706,N_18656);
nor U21074 (N_21074,N_19593,N_19748);
nand U21075 (N_21075,N_18375,N_18235);
and U21076 (N_21076,N_18137,N_18835);
nand U21077 (N_21077,N_19116,N_19471);
nor U21078 (N_21078,N_18251,N_18333);
nor U21079 (N_21079,N_19219,N_18272);
or U21080 (N_21080,N_19517,N_18830);
nor U21081 (N_21081,N_19263,N_18206);
and U21082 (N_21082,N_18272,N_18044);
xor U21083 (N_21083,N_18577,N_19845);
xor U21084 (N_21084,N_18025,N_18499);
xor U21085 (N_21085,N_18888,N_19743);
or U21086 (N_21086,N_19238,N_19527);
nor U21087 (N_21087,N_19039,N_19598);
or U21088 (N_21088,N_18239,N_18760);
and U21089 (N_21089,N_18135,N_18691);
or U21090 (N_21090,N_18717,N_18246);
or U21091 (N_21091,N_18692,N_18949);
nor U21092 (N_21092,N_19527,N_18218);
xor U21093 (N_21093,N_19388,N_19494);
and U21094 (N_21094,N_18995,N_18534);
nor U21095 (N_21095,N_18985,N_18142);
nor U21096 (N_21096,N_18666,N_18930);
nand U21097 (N_21097,N_18579,N_19142);
or U21098 (N_21098,N_18294,N_19152);
or U21099 (N_21099,N_19870,N_19005);
and U21100 (N_21100,N_19843,N_18441);
or U21101 (N_21101,N_18963,N_19857);
and U21102 (N_21102,N_18032,N_18128);
nor U21103 (N_21103,N_19906,N_19180);
nand U21104 (N_21104,N_18211,N_18677);
nand U21105 (N_21105,N_18600,N_18387);
or U21106 (N_21106,N_18355,N_18138);
or U21107 (N_21107,N_18142,N_18035);
or U21108 (N_21108,N_18222,N_18482);
nand U21109 (N_21109,N_18298,N_19492);
or U21110 (N_21110,N_19369,N_18080);
and U21111 (N_21111,N_19006,N_18725);
nor U21112 (N_21112,N_19907,N_18065);
or U21113 (N_21113,N_18879,N_18562);
nand U21114 (N_21114,N_19465,N_19254);
nor U21115 (N_21115,N_19841,N_19801);
xnor U21116 (N_21116,N_19384,N_19824);
xor U21117 (N_21117,N_18953,N_19894);
xnor U21118 (N_21118,N_18920,N_18644);
xnor U21119 (N_21119,N_19279,N_18889);
and U21120 (N_21120,N_19387,N_18126);
nor U21121 (N_21121,N_19070,N_18587);
or U21122 (N_21122,N_19348,N_19222);
nor U21123 (N_21123,N_19715,N_18291);
nor U21124 (N_21124,N_19010,N_19272);
nor U21125 (N_21125,N_19748,N_19958);
xnor U21126 (N_21126,N_19592,N_18325);
nor U21127 (N_21127,N_18214,N_18962);
nand U21128 (N_21128,N_19542,N_18338);
nor U21129 (N_21129,N_19883,N_19094);
and U21130 (N_21130,N_19652,N_18143);
nor U21131 (N_21131,N_18181,N_18232);
xnor U21132 (N_21132,N_19281,N_19662);
nand U21133 (N_21133,N_19544,N_18480);
and U21134 (N_21134,N_19886,N_19856);
or U21135 (N_21135,N_18957,N_18440);
xnor U21136 (N_21136,N_18427,N_19846);
xor U21137 (N_21137,N_19930,N_18379);
or U21138 (N_21138,N_18468,N_19276);
or U21139 (N_21139,N_18195,N_18673);
or U21140 (N_21140,N_18600,N_19369);
xnor U21141 (N_21141,N_19037,N_18913);
or U21142 (N_21142,N_18958,N_19655);
and U21143 (N_21143,N_19782,N_18480);
or U21144 (N_21144,N_19193,N_19961);
nand U21145 (N_21145,N_18002,N_19745);
and U21146 (N_21146,N_18950,N_18217);
and U21147 (N_21147,N_18483,N_18850);
and U21148 (N_21148,N_18275,N_18182);
or U21149 (N_21149,N_18439,N_19146);
nor U21150 (N_21150,N_18292,N_19985);
nand U21151 (N_21151,N_18469,N_19681);
and U21152 (N_21152,N_19164,N_19063);
nand U21153 (N_21153,N_19100,N_18782);
nor U21154 (N_21154,N_19816,N_18640);
or U21155 (N_21155,N_18347,N_18908);
xor U21156 (N_21156,N_18773,N_18087);
xor U21157 (N_21157,N_19240,N_18861);
nor U21158 (N_21158,N_19268,N_18578);
nand U21159 (N_21159,N_19877,N_18063);
and U21160 (N_21160,N_18366,N_19702);
xor U21161 (N_21161,N_18391,N_19896);
or U21162 (N_21162,N_19084,N_18961);
or U21163 (N_21163,N_19250,N_19481);
xnor U21164 (N_21164,N_19605,N_18412);
nand U21165 (N_21165,N_18622,N_18497);
nand U21166 (N_21166,N_18766,N_19625);
nor U21167 (N_21167,N_18731,N_19270);
xnor U21168 (N_21168,N_18047,N_18849);
and U21169 (N_21169,N_18403,N_18416);
xor U21170 (N_21170,N_18973,N_19323);
nor U21171 (N_21171,N_18856,N_18483);
xnor U21172 (N_21172,N_18329,N_18096);
nand U21173 (N_21173,N_19905,N_19842);
xnor U21174 (N_21174,N_19216,N_18001);
nor U21175 (N_21175,N_19308,N_19990);
and U21176 (N_21176,N_19964,N_19422);
nor U21177 (N_21177,N_18839,N_19312);
xor U21178 (N_21178,N_19137,N_18647);
nor U21179 (N_21179,N_18272,N_18594);
or U21180 (N_21180,N_18507,N_18201);
nor U21181 (N_21181,N_19432,N_19188);
nor U21182 (N_21182,N_19438,N_19545);
xnor U21183 (N_21183,N_19786,N_19278);
nor U21184 (N_21184,N_18074,N_19667);
and U21185 (N_21185,N_19329,N_19851);
nor U21186 (N_21186,N_19881,N_19276);
and U21187 (N_21187,N_19328,N_18031);
xor U21188 (N_21188,N_19562,N_19458);
xor U21189 (N_21189,N_19315,N_19953);
xor U21190 (N_21190,N_18957,N_19540);
xor U21191 (N_21191,N_19325,N_18657);
and U21192 (N_21192,N_19718,N_18323);
nand U21193 (N_21193,N_18996,N_19576);
nor U21194 (N_21194,N_18884,N_18018);
xor U21195 (N_21195,N_19330,N_19217);
xnor U21196 (N_21196,N_18860,N_19199);
or U21197 (N_21197,N_19295,N_18985);
or U21198 (N_21198,N_18495,N_19717);
nand U21199 (N_21199,N_19005,N_19611);
xor U21200 (N_21200,N_18590,N_18066);
nor U21201 (N_21201,N_19258,N_18789);
nor U21202 (N_21202,N_18343,N_18826);
nor U21203 (N_21203,N_18720,N_19302);
and U21204 (N_21204,N_19688,N_18851);
nor U21205 (N_21205,N_19940,N_19094);
and U21206 (N_21206,N_19739,N_19720);
and U21207 (N_21207,N_18327,N_18210);
or U21208 (N_21208,N_19705,N_19111);
and U21209 (N_21209,N_19787,N_18588);
and U21210 (N_21210,N_19582,N_19698);
xor U21211 (N_21211,N_18791,N_19200);
nand U21212 (N_21212,N_19191,N_18652);
or U21213 (N_21213,N_19366,N_18065);
and U21214 (N_21214,N_19919,N_18909);
nor U21215 (N_21215,N_19162,N_19539);
nand U21216 (N_21216,N_18997,N_19993);
or U21217 (N_21217,N_19016,N_18007);
or U21218 (N_21218,N_18076,N_19497);
xnor U21219 (N_21219,N_19737,N_18069);
nand U21220 (N_21220,N_18369,N_19545);
and U21221 (N_21221,N_19961,N_18728);
nand U21222 (N_21222,N_18937,N_18137);
or U21223 (N_21223,N_18263,N_19651);
and U21224 (N_21224,N_19356,N_18346);
nand U21225 (N_21225,N_18640,N_18933);
nor U21226 (N_21226,N_19153,N_18185);
and U21227 (N_21227,N_18267,N_19346);
and U21228 (N_21228,N_19130,N_18755);
nor U21229 (N_21229,N_19326,N_18784);
and U21230 (N_21230,N_19513,N_19706);
xnor U21231 (N_21231,N_19414,N_18963);
and U21232 (N_21232,N_19719,N_18311);
or U21233 (N_21233,N_19091,N_18018);
xor U21234 (N_21234,N_18778,N_18281);
xnor U21235 (N_21235,N_19224,N_18053);
or U21236 (N_21236,N_18274,N_18881);
nor U21237 (N_21237,N_18415,N_18092);
xor U21238 (N_21238,N_19827,N_19486);
nor U21239 (N_21239,N_18466,N_18736);
nand U21240 (N_21240,N_19270,N_19387);
xor U21241 (N_21241,N_18178,N_19267);
xnor U21242 (N_21242,N_19330,N_18293);
nor U21243 (N_21243,N_18677,N_18711);
or U21244 (N_21244,N_19827,N_19906);
or U21245 (N_21245,N_18081,N_19734);
nor U21246 (N_21246,N_18215,N_19351);
nand U21247 (N_21247,N_19128,N_18520);
and U21248 (N_21248,N_19357,N_19208);
nor U21249 (N_21249,N_18171,N_18249);
or U21250 (N_21250,N_18130,N_18925);
or U21251 (N_21251,N_18740,N_18829);
or U21252 (N_21252,N_18413,N_18602);
and U21253 (N_21253,N_18667,N_18850);
nor U21254 (N_21254,N_18723,N_19808);
nand U21255 (N_21255,N_19465,N_18822);
or U21256 (N_21256,N_18212,N_18579);
xnor U21257 (N_21257,N_18965,N_18337);
or U21258 (N_21258,N_19818,N_18210);
xnor U21259 (N_21259,N_19623,N_19684);
and U21260 (N_21260,N_18200,N_18058);
and U21261 (N_21261,N_18110,N_18253);
xnor U21262 (N_21262,N_19595,N_18576);
or U21263 (N_21263,N_19598,N_19569);
xnor U21264 (N_21264,N_18436,N_18991);
and U21265 (N_21265,N_18736,N_19702);
xor U21266 (N_21266,N_19614,N_18341);
xor U21267 (N_21267,N_19139,N_18190);
nor U21268 (N_21268,N_19586,N_19219);
or U21269 (N_21269,N_19332,N_19721);
nand U21270 (N_21270,N_19340,N_19675);
xor U21271 (N_21271,N_19042,N_18069);
nor U21272 (N_21272,N_18426,N_19469);
and U21273 (N_21273,N_18425,N_18872);
xor U21274 (N_21274,N_19158,N_19653);
or U21275 (N_21275,N_18303,N_19151);
and U21276 (N_21276,N_19738,N_18165);
or U21277 (N_21277,N_18138,N_19360);
and U21278 (N_21278,N_19985,N_19006);
xor U21279 (N_21279,N_19247,N_18462);
nand U21280 (N_21280,N_18770,N_18767);
nand U21281 (N_21281,N_18466,N_18982);
nand U21282 (N_21282,N_18828,N_19251);
xnor U21283 (N_21283,N_18223,N_19309);
and U21284 (N_21284,N_18382,N_19360);
nand U21285 (N_21285,N_19092,N_18074);
nand U21286 (N_21286,N_18815,N_18841);
or U21287 (N_21287,N_18574,N_18166);
xor U21288 (N_21288,N_18209,N_18347);
xor U21289 (N_21289,N_19581,N_18596);
nor U21290 (N_21290,N_19733,N_19674);
nor U21291 (N_21291,N_19368,N_18948);
or U21292 (N_21292,N_18860,N_18883);
nand U21293 (N_21293,N_18412,N_19752);
nor U21294 (N_21294,N_19992,N_18916);
nor U21295 (N_21295,N_19154,N_19939);
and U21296 (N_21296,N_18829,N_18581);
xor U21297 (N_21297,N_19474,N_18873);
and U21298 (N_21298,N_19299,N_19627);
and U21299 (N_21299,N_18604,N_18028);
or U21300 (N_21300,N_18607,N_19960);
and U21301 (N_21301,N_18754,N_19024);
nor U21302 (N_21302,N_19171,N_19490);
nand U21303 (N_21303,N_18609,N_18063);
xnor U21304 (N_21304,N_19535,N_18758);
xnor U21305 (N_21305,N_19714,N_18153);
and U21306 (N_21306,N_19119,N_18148);
nand U21307 (N_21307,N_19516,N_18539);
nor U21308 (N_21308,N_18230,N_18947);
or U21309 (N_21309,N_18189,N_18788);
or U21310 (N_21310,N_18978,N_19828);
and U21311 (N_21311,N_19112,N_19555);
or U21312 (N_21312,N_19020,N_19544);
xor U21313 (N_21313,N_18654,N_19002);
xnor U21314 (N_21314,N_19439,N_19296);
nand U21315 (N_21315,N_19468,N_18658);
or U21316 (N_21316,N_18445,N_18355);
and U21317 (N_21317,N_18155,N_18680);
or U21318 (N_21318,N_18827,N_18738);
nor U21319 (N_21319,N_19906,N_19877);
xor U21320 (N_21320,N_19134,N_18748);
xor U21321 (N_21321,N_19682,N_19311);
and U21322 (N_21322,N_19843,N_19448);
or U21323 (N_21323,N_18218,N_18435);
nor U21324 (N_21324,N_19158,N_18407);
xnor U21325 (N_21325,N_19834,N_19677);
and U21326 (N_21326,N_19312,N_18328);
xnor U21327 (N_21327,N_18385,N_19899);
nand U21328 (N_21328,N_18570,N_19504);
or U21329 (N_21329,N_18108,N_18247);
or U21330 (N_21330,N_19419,N_18796);
xor U21331 (N_21331,N_18278,N_18547);
or U21332 (N_21332,N_19069,N_18833);
nor U21333 (N_21333,N_18254,N_18837);
or U21334 (N_21334,N_18743,N_18311);
nand U21335 (N_21335,N_19224,N_18632);
xnor U21336 (N_21336,N_19814,N_19598);
nor U21337 (N_21337,N_19254,N_18679);
xnor U21338 (N_21338,N_19131,N_18329);
nor U21339 (N_21339,N_18279,N_18549);
nand U21340 (N_21340,N_18175,N_19880);
and U21341 (N_21341,N_19744,N_19183);
nand U21342 (N_21342,N_19113,N_18170);
nand U21343 (N_21343,N_18149,N_19388);
nand U21344 (N_21344,N_18673,N_18029);
nand U21345 (N_21345,N_19229,N_19427);
xor U21346 (N_21346,N_18410,N_18080);
nor U21347 (N_21347,N_18127,N_18858);
or U21348 (N_21348,N_18918,N_19687);
nor U21349 (N_21349,N_18087,N_18521);
nor U21350 (N_21350,N_18296,N_19020);
or U21351 (N_21351,N_18728,N_18830);
or U21352 (N_21352,N_18434,N_19926);
xnor U21353 (N_21353,N_19959,N_18974);
nand U21354 (N_21354,N_19419,N_18668);
nor U21355 (N_21355,N_18322,N_19015);
and U21356 (N_21356,N_18300,N_19915);
and U21357 (N_21357,N_18851,N_18555);
nand U21358 (N_21358,N_19746,N_18683);
xor U21359 (N_21359,N_19660,N_19699);
and U21360 (N_21360,N_19370,N_18083);
xor U21361 (N_21361,N_18612,N_18259);
or U21362 (N_21362,N_19691,N_19232);
xnor U21363 (N_21363,N_18722,N_19152);
xnor U21364 (N_21364,N_18393,N_18844);
or U21365 (N_21365,N_18083,N_18382);
nand U21366 (N_21366,N_19264,N_19288);
nor U21367 (N_21367,N_18328,N_18473);
nand U21368 (N_21368,N_19329,N_18896);
and U21369 (N_21369,N_19971,N_18705);
nor U21370 (N_21370,N_18213,N_19243);
nor U21371 (N_21371,N_19119,N_18584);
or U21372 (N_21372,N_18037,N_19039);
nand U21373 (N_21373,N_18582,N_18088);
or U21374 (N_21374,N_18381,N_18444);
and U21375 (N_21375,N_19483,N_19764);
and U21376 (N_21376,N_19383,N_18768);
nor U21377 (N_21377,N_19034,N_19473);
and U21378 (N_21378,N_18508,N_18970);
and U21379 (N_21379,N_19647,N_18197);
nor U21380 (N_21380,N_19638,N_19854);
nor U21381 (N_21381,N_19880,N_19461);
xnor U21382 (N_21382,N_18192,N_18361);
or U21383 (N_21383,N_18925,N_19396);
or U21384 (N_21384,N_19308,N_19524);
or U21385 (N_21385,N_18317,N_19125);
and U21386 (N_21386,N_19783,N_19664);
or U21387 (N_21387,N_18426,N_18281);
and U21388 (N_21388,N_18251,N_19688);
nor U21389 (N_21389,N_19993,N_18674);
nand U21390 (N_21390,N_19298,N_19019);
nor U21391 (N_21391,N_18228,N_18266);
and U21392 (N_21392,N_18088,N_18510);
nand U21393 (N_21393,N_18972,N_18744);
xnor U21394 (N_21394,N_18531,N_19828);
and U21395 (N_21395,N_18459,N_19283);
nand U21396 (N_21396,N_18353,N_18868);
and U21397 (N_21397,N_19626,N_19410);
nand U21398 (N_21398,N_19448,N_18523);
xor U21399 (N_21399,N_19944,N_19508);
xor U21400 (N_21400,N_18560,N_18361);
nand U21401 (N_21401,N_18252,N_19242);
and U21402 (N_21402,N_19974,N_19833);
and U21403 (N_21403,N_18696,N_19727);
xor U21404 (N_21404,N_19522,N_19153);
xor U21405 (N_21405,N_18860,N_18367);
nand U21406 (N_21406,N_18158,N_19032);
nand U21407 (N_21407,N_19042,N_19080);
and U21408 (N_21408,N_19199,N_18155);
and U21409 (N_21409,N_19627,N_19240);
xor U21410 (N_21410,N_18118,N_19012);
and U21411 (N_21411,N_18133,N_19348);
and U21412 (N_21412,N_18050,N_18686);
nor U21413 (N_21413,N_19012,N_18073);
nor U21414 (N_21414,N_19578,N_19303);
nor U21415 (N_21415,N_18641,N_19098);
or U21416 (N_21416,N_19950,N_18584);
and U21417 (N_21417,N_19597,N_19300);
nor U21418 (N_21418,N_18328,N_18064);
nand U21419 (N_21419,N_19107,N_18596);
nand U21420 (N_21420,N_18193,N_19018);
nand U21421 (N_21421,N_19057,N_18898);
xnor U21422 (N_21422,N_19125,N_19443);
and U21423 (N_21423,N_18840,N_19031);
xor U21424 (N_21424,N_19867,N_18077);
and U21425 (N_21425,N_19174,N_19079);
and U21426 (N_21426,N_18432,N_18668);
and U21427 (N_21427,N_19951,N_19071);
and U21428 (N_21428,N_19722,N_19860);
xnor U21429 (N_21429,N_19410,N_19516);
nand U21430 (N_21430,N_19509,N_19276);
or U21431 (N_21431,N_18132,N_18101);
nand U21432 (N_21432,N_18992,N_18608);
nand U21433 (N_21433,N_18031,N_19713);
nor U21434 (N_21434,N_19868,N_19675);
and U21435 (N_21435,N_19223,N_18375);
nor U21436 (N_21436,N_19414,N_19785);
xor U21437 (N_21437,N_19727,N_18307);
nand U21438 (N_21438,N_18305,N_19292);
xor U21439 (N_21439,N_18213,N_19979);
nand U21440 (N_21440,N_19136,N_19475);
nand U21441 (N_21441,N_19393,N_18177);
or U21442 (N_21442,N_18275,N_19629);
or U21443 (N_21443,N_19208,N_19059);
nor U21444 (N_21444,N_18389,N_19078);
nand U21445 (N_21445,N_19673,N_18218);
and U21446 (N_21446,N_18193,N_18460);
xor U21447 (N_21447,N_19352,N_19100);
nor U21448 (N_21448,N_18436,N_19401);
nor U21449 (N_21449,N_19622,N_18643);
nand U21450 (N_21450,N_19118,N_18099);
xor U21451 (N_21451,N_18440,N_19326);
and U21452 (N_21452,N_18816,N_19459);
and U21453 (N_21453,N_18695,N_18452);
and U21454 (N_21454,N_18575,N_19390);
xnor U21455 (N_21455,N_19428,N_18710);
or U21456 (N_21456,N_19250,N_19582);
and U21457 (N_21457,N_18635,N_19964);
nor U21458 (N_21458,N_19725,N_18246);
nand U21459 (N_21459,N_19532,N_18849);
nand U21460 (N_21460,N_18462,N_18629);
and U21461 (N_21461,N_19953,N_19962);
xor U21462 (N_21462,N_19401,N_19639);
xor U21463 (N_21463,N_19362,N_18199);
nand U21464 (N_21464,N_18304,N_19489);
and U21465 (N_21465,N_18534,N_19089);
nand U21466 (N_21466,N_19029,N_19410);
nor U21467 (N_21467,N_19672,N_18423);
and U21468 (N_21468,N_18499,N_19468);
or U21469 (N_21469,N_18405,N_19198);
and U21470 (N_21470,N_18378,N_18148);
xnor U21471 (N_21471,N_19945,N_18437);
nor U21472 (N_21472,N_18682,N_18991);
or U21473 (N_21473,N_19141,N_18856);
or U21474 (N_21474,N_18658,N_19816);
nand U21475 (N_21475,N_18478,N_19003);
nand U21476 (N_21476,N_18279,N_19862);
nand U21477 (N_21477,N_19366,N_19600);
nor U21478 (N_21478,N_18691,N_18197);
and U21479 (N_21479,N_19502,N_18719);
xor U21480 (N_21480,N_18406,N_19601);
and U21481 (N_21481,N_19163,N_19735);
xor U21482 (N_21482,N_18636,N_18006);
nor U21483 (N_21483,N_18618,N_19054);
and U21484 (N_21484,N_19876,N_19101);
and U21485 (N_21485,N_19381,N_18950);
and U21486 (N_21486,N_19665,N_18559);
xor U21487 (N_21487,N_19848,N_18246);
and U21488 (N_21488,N_18994,N_19505);
nand U21489 (N_21489,N_19486,N_19340);
and U21490 (N_21490,N_18707,N_19578);
or U21491 (N_21491,N_18922,N_19046);
and U21492 (N_21492,N_18169,N_18931);
or U21493 (N_21493,N_19293,N_18644);
nand U21494 (N_21494,N_19576,N_18741);
xnor U21495 (N_21495,N_18905,N_19409);
nand U21496 (N_21496,N_19591,N_18773);
and U21497 (N_21497,N_19926,N_19399);
nand U21498 (N_21498,N_19456,N_18088);
nor U21499 (N_21499,N_18392,N_19790);
nor U21500 (N_21500,N_18985,N_19126);
nand U21501 (N_21501,N_18817,N_19744);
nor U21502 (N_21502,N_18887,N_19122);
nand U21503 (N_21503,N_18361,N_18328);
nand U21504 (N_21504,N_18834,N_19121);
nor U21505 (N_21505,N_19814,N_19272);
or U21506 (N_21506,N_19964,N_19500);
xor U21507 (N_21507,N_18298,N_18063);
nor U21508 (N_21508,N_18544,N_19993);
and U21509 (N_21509,N_19478,N_18705);
nand U21510 (N_21510,N_19132,N_18729);
and U21511 (N_21511,N_19506,N_18319);
or U21512 (N_21512,N_18907,N_19369);
nand U21513 (N_21513,N_19939,N_19024);
nor U21514 (N_21514,N_19011,N_19070);
and U21515 (N_21515,N_19227,N_18758);
nand U21516 (N_21516,N_19347,N_18582);
xor U21517 (N_21517,N_18904,N_18069);
xnor U21518 (N_21518,N_19696,N_18930);
or U21519 (N_21519,N_19966,N_19615);
and U21520 (N_21520,N_19335,N_19344);
or U21521 (N_21521,N_19158,N_19051);
nor U21522 (N_21522,N_19757,N_18732);
or U21523 (N_21523,N_18708,N_19381);
or U21524 (N_21524,N_18558,N_19802);
nand U21525 (N_21525,N_19386,N_18291);
nand U21526 (N_21526,N_18679,N_18563);
nor U21527 (N_21527,N_19570,N_19527);
nor U21528 (N_21528,N_18750,N_19391);
or U21529 (N_21529,N_18654,N_19301);
and U21530 (N_21530,N_18020,N_18632);
or U21531 (N_21531,N_19133,N_19539);
and U21532 (N_21532,N_19876,N_18057);
nand U21533 (N_21533,N_19723,N_18244);
nand U21534 (N_21534,N_18921,N_19516);
or U21535 (N_21535,N_19248,N_18324);
and U21536 (N_21536,N_19088,N_18674);
nand U21537 (N_21537,N_18462,N_18619);
xor U21538 (N_21538,N_18158,N_18462);
nand U21539 (N_21539,N_18302,N_19949);
or U21540 (N_21540,N_18340,N_19937);
or U21541 (N_21541,N_19268,N_18908);
nor U21542 (N_21542,N_19250,N_18744);
nor U21543 (N_21543,N_19437,N_19474);
nor U21544 (N_21544,N_19974,N_19454);
nor U21545 (N_21545,N_19792,N_19534);
nor U21546 (N_21546,N_19301,N_19111);
nand U21547 (N_21547,N_18864,N_18543);
nand U21548 (N_21548,N_19577,N_19392);
or U21549 (N_21549,N_19120,N_18642);
nor U21550 (N_21550,N_19468,N_18697);
xnor U21551 (N_21551,N_18439,N_19661);
or U21552 (N_21552,N_18479,N_19245);
and U21553 (N_21553,N_18119,N_19395);
or U21554 (N_21554,N_19817,N_18422);
nand U21555 (N_21555,N_19029,N_18384);
and U21556 (N_21556,N_18574,N_18646);
nand U21557 (N_21557,N_18619,N_19421);
xor U21558 (N_21558,N_18533,N_19910);
nand U21559 (N_21559,N_18938,N_18159);
xor U21560 (N_21560,N_19818,N_19003);
nor U21561 (N_21561,N_19860,N_18499);
nand U21562 (N_21562,N_19111,N_18177);
nand U21563 (N_21563,N_19590,N_19246);
xor U21564 (N_21564,N_19657,N_19201);
xor U21565 (N_21565,N_18825,N_19242);
xor U21566 (N_21566,N_19242,N_18369);
nor U21567 (N_21567,N_18116,N_19020);
or U21568 (N_21568,N_18241,N_18116);
xnor U21569 (N_21569,N_18325,N_18171);
nand U21570 (N_21570,N_18520,N_19230);
xnor U21571 (N_21571,N_19154,N_19086);
nand U21572 (N_21572,N_19671,N_18854);
xor U21573 (N_21573,N_18165,N_18030);
and U21574 (N_21574,N_18214,N_18996);
xnor U21575 (N_21575,N_18813,N_18107);
nand U21576 (N_21576,N_19945,N_18242);
xnor U21577 (N_21577,N_18537,N_18589);
nand U21578 (N_21578,N_18536,N_19954);
nand U21579 (N_21579,N_19542,N_19917);
and U21580 (N_21580,N_18171,N_18288);
xnor U21581 (N_21581,N_19349,N_19083);
xnor U21582 (N_21582,N_18636,N_19339);
xnor U21583 (N_21583,N_19681,N_19128);
nor U21584 (N_21584,N_19540,N_18014);
xor U21585 (N_21585,N_19155,N_19611);
nor U21586 (N_21586,N_19237,N_19527);
and U21587 (N_21587,N_19712,N_19133);
and U21588 (N_21588,N_18470,N_18413);
nand U21589 (N_21589,N_19829,N_19071);
nand U21590 (N_21590,N_19045,N_18114);
nand U21591 (N_21591,N_18709,N_18043);
and U21592 (N_21592,N_19514,N_19659);
and U21593 (N_21593,N_18322,N_18303);
nand U21594 (N_21594,N_18202,N_18359);
xnor U21595 (N_21595,N_18882,N_18183);
or U21596 (N_21596,N_19839,N_19086);
or U21597 (N_21597,N_18611,N_18684);
xor U21598 (N_21598,N_18026,N_18401);
xnor U21599 (N_21599,N_19306,N_18470);
xor U21600 (N_21600,N_19788,N_18234);
nor U21601 (N_21601,N_19626,N_19785);
nand U21602 (N_21602,N_19586,N_19569);
nand U21603 (N_21603,N_18464,N_18632);
and U21604 (N_21604,N_19466,N_18169);
and U21605 (N_21605,N_18742,N_18501);
nand U21606 (N_21606,N_18342,N_18952);
xnor U21607 (N_21607,N_19513,N_19786);
nand U21608 (N_21608,N_19967,N_18764);
nor U21609 (N_21609,N_18184,N_18435);
xor U21610 (N_21610,N_18274,N_19400);
and U21611 (N_21611,N_18092,N_19632);
xnor U21612 (N_21612,N_19579,N_18157);
xor U21613 (N_21613,N_18733,N_18844);
and U21614 (N_21614,N_18224,N_19906);
and U21615 (N_21615,N_18853,N_18772);
and U21616 (N_21616,N_18297,N_19192);
or U21617 (N_21617,N_18024,N_19617);
or U21618 (N_21618,N_18020,N_18825);
nor U21619 (N_21619,N_18845,N_18369);
xor U21620 (N_21620,N_19091,N_19264);
nor U21621 (N_21621,N_19766,N_19847);
nand U21622 (N_21622,N_19522,N_18756);
and U21623 (N_21623,N_18942,N_19501);
xnor U21624 (N_21624,N_18649,N_18451);
and U21625 (N_21625,N_19651,N_19256);
nor U21626 (N_21626,N_18425,N_18949);
nor U21627 (N_21627,N_18333,N_18632);
or U21628 (N_21628,N_18919,N_18129);
and U21629 (N_21629,N_19330,N_18969);
xnor U21630 (N_21630,N_18630,N_19633);
xnor U21631 (N_21631,N_18276,N_18418);
nand U21632 (N_21632,N_18271,N_19766);
and U21633 (N_21633,N_18262,N_19213);
and U21634 (N_21634,N_18503,N_19015);
nand U21635 (N_21635,N_19459,N_18856);
or U21636 (N_21636,N_18064,N_18160);
xnor U21637 (N_21637,N_18330,N_18853);
or U21638 (N_21638,N_18087,N_19539);
xnor U21639 (N_21639,N_19158,N_18638);
nand U21640 (N_21640,N_18953,N_19959);
nor U21641 (N_21641,N_18324,N_19685);
nand U21642 (N_21642,N_18241,N_18829);
nand U21643 (N_21643,N_18583,N_19421);
nand U21644 (N_21644,N_19576,N_18130);
xnor U21645 (N_21645,N_18974,N_18470);
nand U21646 (N_21646,N_19153,N_19455);
xor U21647 (N_21647,N_19078,N_18039);
and U21648 (N_21648,N_18576,N_19053);
xnor U21649 (N_21649,N_19413,N_18215);
nand U21650 (N_21650,N_19814,N_18042);
nor U21651 (N_21651,N_18642,N_18009);
or U21652 (N_21652,N_19769,N_19553);
nand U21653 (N_21653,N_18061,N_19789);
and U21654 (N_21654,N_18831,N_18433);
nor U21655 (N_21655,N_19207,N_18986);
xnor U21656 (N_21656,N_18343,N_18228);
and U21657 (N_21657,N_18002,N_19501);
nor U21658 (N_21658,N_19345,N_19408);
nor U21659 (N_21659,N_18835,N_18551);
or U21660 (N_21660,N_18714,N_19880);
nand U21661 (N_21661,N_18559,N_18297);
nor U21662 (N_21662,N_18704,N_19011);
or U21663 (N_21663,N_19276,N_18529);
nor U21664 (N_21664,N_19469,N_19603);
or U21665 (N_21665,N_18848,N_18237);
or U21666 (N_21666,N_18228,N_18261);
xor U21667 (N_21667,N_18902,N_18276);
xnor U21668 (N_21668,N_19125,N_18370);
nor U21669 (N_21669,N_19364,N_19503);
or U21670 (N_21670,N_19153,N_19815);
and U21671 (N_21671,N_18062,N_19791);
xnor U21672 (N_21672,N_18084,N_19740);
nand U21673 (N_21673,N_19345,N_19360);
or U21674 (N_21674,N_19193,N_19181);
xnor U21675 (N_21675,N_18332,N_19002);
xor U21676 (N_21676,N_19847,N_19233);
or U21677 (N_21677,N_18053,N_19030);
or U21678 (N_21678,N_18180,N_18266);
nor U21679 (N_21679,N_19594,N_19634);
nor U21680 (N_21680,N_18939,N_19452);
and U21681 (N_21681,N_19221,N_19812);
or U21682 (N_21682,N_19238,N_19734);
or U21683 (N_21683,N_18216,N_19857);
or U21684 (N_21684,N_19281,N_18074);
nand U21685 (N_21685,N_19028,N_18721);
nor U21686 (N_21686,N_19431,N_18880);
nand U21687 (N_21687,N_19047,N_18862);
and U21688 (N_21688,N_18290,N_18115);
nand U21689 (N_21689,N_19385,N_19864);
xor U21690 (N_21690,N_19376,N_19924);
and U21691 (N_21691,N_18599,N_18219);
xnor U21692 (N_21692,N_18933,N_18026);
or U21693 (N_21693,N_18224,N_18388);
nor U21694 (N_21694,N_18623,N_18915);
and U21695 (N_21695,N_18513,N_18412);
nor U21696 (N_21696,N_19440,N_19326);
and U21697 (N_21697,N_19319,N_19138);
nand U21698 (N_21698,N_19081,N_18998);
nor U21699 (N_21699,N_18360,N_19633);
or U21700 (N_21700,N_19505,N_19850);
and U21701 (N_21701,N_18026,N_18523);
and U21702 (N_21702,N_19944,N_18815);
nor U21703 (N_21703,N_18953,N_19069);
nand U21704 (N_21704,N_19452,N_18269);
nor U21705 (N_21705,N_18030,N_18346);
xnor U21706 (N_21706,N_19041,N_18915);
xor U21707 (N_21707,N_19596,N_18517);
nor U21708 (N_21708,N_18746,N_18401);
xnor U21709 (N_21709,N_18735,N_19145);
nand U21710 (N_21710,N_18245,N_18734);
xnor U21711 (N_21711,N_18765,N_18618);
and U21712 (N_21712,N_19275,N_19964);
nand U21713 (N_21713,N_19786,N_18123);
or U21714 (N_21714,N_18631,N_19067);
nand U21715 (N_21715,N_19185,N_18290);
or U21716 (N_21716,N_19934,N_19498);
nor U21717 (N_21717,N_19903,N_19538);
or U21718 (N_21718,N_18900,N_18610);
or U21719 (N_21719,N_19200,N_18351);
nor U21720 (N_21720,N_19833,N_19070);
xnor U21721 (N_21721,N_18383,N_18320);
or U21722 (N_21722,N_18036,N_18769);
xnor U21723 (N_21723,N_19151,N_19581);
and U21724 (N_21724,N_19390,N_19123);
nand U21725 (N_21725,N_19136,N_18188);
or U21726 (N_21726,N_18714,N_19172);
nand U21727 (N_21727,N_19525,N_18772);
and U21728 (N_21728,N_18849,N_19762);
xnor U21729 (N_21729,N_19069,N_19400);
nor U21730 (N_21730,N_19602,N_19856);
nand U21731 (N_21731,N_18900,N_19211);
nor U21732 (N_21732,N_19747,N_18322);
or U21733 (N_21733,N_18445,N_18943);
xnor U21734 (N_21734,N_18794,N_19217);
nand U21735 (N_21735,N_19694,N_19790);
and U21736 (N_21736,N_18957,N_19530);
nand U21737 (N_21737,N_19026,N_19681);
and U21738 (N_21738,N_18545,N_19766);
nand U21739 (N_21739,N_18706,N_19763);
or U21740 (N_21740,N_18707,N_18078);
or U21741 (N_21741,N_19833,N_18823);
nor U21742 (N_21742,N_18000,N_18383);
and U21743 (N_21743,N_18580,N_19500);
xnor U21744 (N_21744,N_18744,N_18209);
nor U21745 (N_21745,N_19623,N_19496);
nor U21746 (N_21746,N_18635,N_19218);
nor U21747 (N_21747,N_19338,N_18031);
xor U21748 (N_21748,N_18595,N_19016);
and U21749 (N_21749,N_18752,N_18057);
nor U21750 (N_21750,N_19574,N_18426);
nor U21751 (N_21751,N_18979,N_19791);
and U21752 (N_21752,N_19155,N_19217);
nor U21753 (N_21753,N_18354,N_18656);
nor U21754 (N_21754,N_18801,N_18880);
and U21755 (N_21755,N_18933,N_18990);
xor U21756 (N_21756,N_18848,N_18785);
and U21757 (N_21757,N_18492,N_19791);
or U21758 (N_21758,N_19291,N_19452);
and U21759 (N_21759,N_18630,N_18854);
nor U21760 (N_21760,N_19241,N_18765);
nor U21761 (N_21761,N_19838,N_19436);
or U21762 (N_21762,N_19242,N_19611);
nor U21763 (N_21763,N_19001,N_19979);
nor U21764 (N_21764,N_18147,N_19169);
xnor U21765 (N_21765,N_19787,N_18284);
or U21766 (N_21766,N_19912,N_19406);
nor U21767 (N_21767,N_19974,N_18302);
or U21768 (N_21768,N_18929,N_19229);
nand U21769 (N_21769,N_18463,N_19361);
or U21770 (N_21770,N_18992,N_18739);
xor U21771 (N_21771,N_18522,N_19454);
or U21772 (N_21772,N_19631,N_19003);
nor U21773 (N_21773,N_19141,N_19818);
nand U21774 (N_21774,N_18902,N_18226);
nand U21775 (N_21775,N_19454,N_18875);
xor U21776 (N_21776,N_19782,N_19800);
or U21777 (N_21777,N_19004,N_18463);
nor U21778 (N_21778,N_18108,N_18270);
nor U21779 (N_21779,N_19215,N_19942);
and U21780 (N_21780,N_18895,N_19474);
nor U21781 (N_21781,N_19360,N_18181);
nand U21782 (N_21782,N_18029,N_18627);
nand U21783 (N_21783,N_19583,N_19845);
and U21784 (N_21784,N_19234,N_19861);
nor U21785 (N_21785,N_18399,N_19808);
nor U21786 (N_21786,N_18360,N_18885);
xor U21787 (N_21787,N_19070,N_19619);
xnor U21788 (N_21788,N_18018,N_19236);
xnor U21789 (N_21789,N_18350,N_19943);
nand U21790 (N_21790,N_19349,N_18610);
and U21791 (N_21791,N_19561,N_18273);
xnor U21792 (N_21792,N_18305,N_19722);
or U21793 (N_21793,N_18774,N_19385);
xnor U21794 (N_21794,N_19637,N_18156);
nand U21795 (N_21795,N_18099,N_19212);
or U21796 (N_21796,N_18808,N_18218);
nor U21797 (N_21797,N_19162,N_19286);
nor U21798 (N_21798,N_19992,N_19014);
or U21799 (N_21799,N_19458,N_19661);
xor U21800 (N_21800,N_18360,N_18437);
nand U21801 (N_21801,N_18903,N_19639);
nor U21802 (N_21802,N_18255,N_19328);
nand U21803 (N_21803,N_18267,N_19897);
or U21804 (N_21804,N_18415,N_18254);
or U21805 (N_21805,N_18507,N_19185);
nor U21806 (N_21806,N_19258,N_18837);
xnor U21807 (N_21807,N_18343,N_18404);
and U21808 (N_21808,N_19612,N_18482);
or U21809 (N_21809,N_18874,N_18007);
or U21810 (N_21810,N_18272,N_19324);
xnor U21811 (N_21811,N_19583,N_19206);
nor U21812 (N_21812,N_19494,N_19393);
xnor U21813 (N_21813,N_19355,N_18578);
nor U21814 (N_21814,N_18548,N_18142);
or U21815 (N_21815,N_18129,N_18047);
or U21816 (N_21816,N_19665,N_18805);
xor U21817 (N_21817,N_19074,N_19889);
and U21818 (N_21818,N_18272,N_18888);
nor U21819 (N_21819,N_18314,N_18252);
nor U21820 (N_21820,N_18868,N_18647);
xor U21821 (N_21821,N_19326,N_19439);
nor U21822 (N_21822,N_19386,N_18179);
and U21823 (N_21823,N_18467,N_19455);
and U21824 (N_21824,N_19722,N_19765);
xnor U21825 (N_21825,N_18941,N_18161);
xnor U21826 (N_21826,N_18116,N_18399);
nor U21827 (N_21827,N_18396,N_18057);
nand U21828 (N_21828,N_19153,N_18812);
and U21829 (N_21829,N_19009,N_19966);
xnor U21830 (N_21830,N_18517,N_19843);
or U21831 (N_21831,N_19309,N_19078);
or U21832 (N_21832,N_19027,N_18532);
and U21833 (N_21833,N_19887,N_19893);
nand U21834 (N_21834,N_19513,N_19373);
nand U21835 (N_21835,N_18577,N_19681);
and U21836 (N_21836,N_19087,N_19134);
nand U21837 (N_21837,N_18567,N_19979);
xor U21838 (N_21838,N_18814,N_18182);
nor U21839 (N_21839,N_18270,N_18655);
or U21840 (N_21840,N_19451,N_19854);
xor U21841 (N_21841,N_18218,N_19050);
nor U21842 (N_21842,N_19911,N_18822);
nor U21843 (N_21843,N_18527,N_19468);
or U21844 (N_21844,N_19524,N_18576);
xnor U21845 (N_21845,N_19910,N_19184);
nand U21846 (N_21846,N_18472,N_18588);
nor U21847 (N_21847,N_18933,N_19876);
and U21848 (N_21848,N_19539,N_18812);
nor U21849 (N_21849,N_19499,N_19468);
nor U21850 (N_21850,N_19636,N_18492);
nor U21851 (N_21851,N_19730,N_18999);
xnor U21852 (N_21852,N_19378,N_18971);
nand U21853 (N_21853,N_18491,N_18605);
nor U21854 (N_21854,N_18281,N_18567);
xor U21855 (N_21855,N_18670,N_18989);
or U21856 (N_21856,N_18313,N_19848);
and U21857 (N_21857,N_19825,N_18864);
nor U21858 (N_21858,N_18410,N_18788);
or U21859 (N_21859,N_18901,N_19233);
or U21860 (N_21860,N_19235,N_19487);
xor U21861 (N_21861,N_18090,N_18307);
nand U21862 (N_21862,N_19103,N_19105);
nor U21863 (N_21863,N_19149,N_18138);
nand U21864 (N_21864,N_19247,N_19125);
nand U21865 (N_21865,N_18390,N_18682);
nor U21866 (N_21866,N_19169,N_19250);
nand U21867 (N_21867,N_19839,N_18158);
or U21868 (N_21868,N_18162,N_18089);
and U21869 (N_21869,N_18473,N_18165);
xor U21870 (N_21870,N_19559,N_19810);
and U21871 (N_21871,N_19469,N_18823);
nand U21872 (N_21872,N_18898,N_18134);
nor U21873 (N_21873,N_18221,N_19809);
or U21874 (N_21874,N_19202,N_19111);
or U21875 (N_21875,N_18882,N_19223);
and U21876 (N_21876,N_18978,N_19044);
and U21877 (N_21877,N_19369,N_19762);
nor U21878 (N_21878,N_18662,N_18319);
nor U21879 (N_21879,N_18562,N_18289);
or U21880 (N_21880,N_19348,N_18246);
nor U21881 (N_21881,N_19902,N_18109);
and U21882 (N_21882,N_18443,N_18620);
nor U21883 (N_21883,N_19148,N_19134);
nor U21884 (N_21884,N_18628,N_18900);
nor U21885 (N_21885,N_18068,N_18426);
nor U21886 (N_21886,N_18169,N_18510);
or U21887 (N_21887,N_19744,N_18700);
nor U21888 (N_21888,N_18367,N_19560);
and U21889 (N_21889,N_19352,N_19193);
or U21890 (N_21890,N_19425,N_18677);
and U21891 (N_21891,N_19692,N_18608);
or U21892 (N_21892,N_19900,N_18747);
nor U21893 (N_21893,N_19856,N_18301);
xnor U21894 (N_21894,N_18677,N_19136);
xor U21895 (N_21895,N_19208,N_19037);
nor U21896 (N_21896,N_18806,N_19925);
nand U21897 (N_21897,N_19478,N_19928);
and U21898 (N_21898,N_19614,N_18961);
nand U21899 (N_21899,N_19088,N_19766);
xnor U21900 (N_21900,N_19853,N_18603);
xor U21901 (N_21901,N_18288,N_18386);
and U21902 (N_21902,N_18857,N_18250);
nand U21903 (N_21903,N_18107,N_19311);
or U21904 (N_21904,N_19820,N_18516);
nor U21905 (N_21905,N_19652,N_18740);
nand U21906 (N_21906,N_19862,N_19607);
xnor U21907 (N_21907,N_18047,N_18416);
and U21908 (N_21908,N_18605,N_18179);
xor U21909 (N_21909,N_19162,N_18849);
nand U21910 (N_21910,N_19763,N_19102);
nand U21911 (N_21911,N_18747,N_18895);
and U21912 (N_21912,N_19499,N_19772);
and U21913 (N_21913,N_19771,N_19211);
nand U21914 (N_21914,N_19622,N_19883);
xor U21915 (N_21915,N_19027,N_18400);
nand U21916 (N_21916,N_19384,N_19231);
xnor U21917 (N_21917,N_18802,N_19597);
and U21918 (N_21918,N_19012,N_18126);
nor U21919 (N_21919,N_19353,N_19314);
nand U21920 (N_21920,N_18457,N_18234);
and U21921 (N_21921,N_18189,N_19155);
nor U21922 (N_21922,N_19279,N_18823);
and U21923 (N_21923,N_19409,N_19232);
and U21924 (N_21924,N_19642,N_19900);
nand U21925 (N_21925,N_18870,N_18956);
nor U21926 (N_21926,N_18199,N_18793);
and U21927 (N_21927,N_19025,N_19587);
xor U21928 (N_21928,N_19736,N_19230);
xnor U21929 (N_21929,N_18760,N_18851);
or U21930 (N_21930,N_19833,N_19167);
nand U21931 (N_21931,N_18820,N_18345);
or U21932 (N_21932,N_18571,N_18460);
nor U21933 (N_21933,N_18454,N_18861);
and U21934 (N_21934,N_19441,N_18783);
nand U21935 (N_21935,N_18874,N_19870);
xor U21936 (N_21936,N_19145,N_18395);
xor U21937 (N_21937,N_19038,N_19897);
nor U21938 (N_21938,N_19810,N_19688);
nand U21939 (N_21939,N_18005,N_18672);
nor U21940 (N_21940,N_18215,N_18517);
nor U21941 (N_21941,N_18525,N_19019);
nor U21942 (N_21942,N_18716,N_18068);
and U21943 (N_21943,N_19565,N_19603);
nand U21944 (N_21944,N_19575,N_19589);
or U21945 (N_21945,N_19153,N_19773);
nand U21946 (N_21946,N_19150,N_18433);
nand U21947 (N_21947,N_19632,N_19440);
nand U21948 (N_21948,N_19970,N_18175);
xor U21949 (N_21949,N_18677,N_18321);
nand U21950 (N_21950,N_18580,N_18164);
xnor U21951 (N_21951,N_19506,N_19732);
nor U21952 (N_21952,N_19001,N_19327);
xnor U21953 (N_21953,N_19292,N_18339);
or U21954 (N_21954,N_19832,N_19533);
xnor U21955 (N_21955,N_19452,N_18958);
nand U21956 (N_21956,N_18750,N_19143);
nand U21957 (N_21957,N_19538,N_18553);
nor U21958 (N_21958,N_18713,N_18892);
or U21959 (N_21959,N_18018,N_18838);
nand U21960 (N_21960,N_19797,N_18642);
nand U21961 (N_21961,N_18547,N_19072);
nor U21962 (N_21962,N_18114,N_18196);
nand U21963 (N_21963,N_19993,N_18587);
and U21964 (N_21964,N_18144,N_19074);
and U21965 (N_21965,N_18388,N_19174);
nand U21966 (N_21966,N_19953,N_19083);
nor U21967 (N_21967,N_18430,N_19391);
nand U21968 (N_21968,N_18250,N_18551);
xnor U21969 (N_21969,N_19790,N_19805);
and U21970 (N_21970,N_18964,N_19705);
and U21971 (N_21971,N_19189,N_18613);
nand U21972 (N_21972,N_19472,N_19356);
nand U21973 (N_21973,N_19281,N_18565);
or U21974 (N_21974,N_18554,N_19969);
nand U21975 (N_21975,N_18920,N_18320);
or U21976 (N_21976,N_19719,N_19802);
nor U21977 (N_21977,N_19605,N_18430);
xor U21978 (N_21978,N_18841,N_18502);
xor U21979 (N_21979,N_19601,N_19178);
nor U21980 (N_21980,N_19735,N_19066);
or U21981 (N_21981,N_18687,N_18670);
and U21982 (N_21982,N_18523,N_18218);
xor U21983 (N_21983,N_18465,N_19036);
and U21984 (N_21984,N_19171,N_18512);
nand U21985 (N_21985,N_18433,N_19727);
and U21986 (N_21986,N_18872,N_19513);
and U21987 (N_21987,N_18707,N_18213);
nand U21988 (N_21988,N_18887,N_18885);
xnor U21989 (N_21989,N_18934,N_19711);
or U21990 (N_21990,N_19874,N_18924);
xnor U21991 (N_21991,N_18970,N_19184);
or U21992 (N_21992,N_18522,N_18478);
nand U21993 (N_21993,N_18520,N_18492);
nor U21994 (N_21994,N_18305,N_18010);
xnor U21995 (N_21995,N_19780,N_18121);
xor U21996 (N_21996,N_18300,N_19435);
xnor U21997 (N_21997,N_19319,N_18814);
or U21998 (N_21998,N_18151,N_19996);
nor U21999 (N_21999,N_18389,N_19823);
nor U22000 (N_22000,N_21091,N_20095);
and U22001 (N_22001,N_21162,N_21139);
nor U22002 (N_22002,N_20288,N_21810);
or U22003 (N_22003,N_21489,N_21927);
nor U22004 (N_22004,N_20558,N_20720);
nand U22005 (N_22005,N_21526,N_20213);
xnor U22006 (N_22006,N_21593,N_21147);
and U22007 (N_22007,N_21754,N_20450);
or U22008 (N_22008,N_20191,N_21532);
and U22009 (N_22009,N_20399,N_20397);
xor U22010 (N_22010,N_20634,N_20292);
or U22011 (N_22011,N_21006,N_21327);
nor U22012 (N_22012,N_21846,N_20052);
nand U22013 (N_22013,N_20918,N_21455);
nor U22014 (N_22014,N_20702,N_20856);
xor U22015 (N_22015,N_20482,N_20198);
and U22016 (N_22016,N_21764,N_21932);
nand U22017 (N_22017,N_21521,N_20618);
nand U22018 (N_22018,N_20346,N_20907);
nand U22019 (N_22019,N_20464,N_20815);
and U22020 (N_22020,N_20951,N_21961);
nand U22021 (N_22021,N_21657,N_20961);
and U22022 (N_22022,N_20525,N_20428);
or U22023 (N_22023,N_21705,N_20523);
or U22024 (N_22024,N_20647,N_21237);
and U22025 (N_22025,N_21769,N_20890);
xnor U22026 (N_22026,N_20559,N_21038);
or U22027 (N_22027,N_21684,N_20949);
xor U22028 (N_22028,N_21266,N_21408);
or U22029 (N_22029,N_21074,N_20034);
nand U22030 (N_22030,N_21797,N_20171);
xnor U22031 (N_22031,N_21454,N_20361);
or U22032 (N_22032,N_20929,N_21438);
nand U22033 (N_22033,N_20646,N_20697);
or U22034 (N_22034,N_20148,N_21807);
or U22035 (N_22035,N_20917,N_20294);
or U22036 (N_22036,N_20841,N_20472);
or U22037 (N_22037,N_20109,N_21387);
and U22038 (N_22038,N_21420,N_20817);
nor U22039 (N_22039,N_20133,N_20421);
nand U22040 (N_22040,N_20099,N_21201);
nand U22041 (N_22041,N_20278,N_21771);
or U22042 (N_22042,N_21403,N_21558);
and U22043 (N_22043,N_21843,N_20729);
nor U22044 (N_22044,N_20826,N_21533);
or U22045 (N_22045,N_21209,N_20533);
xor U22046 (N_22046,N_20067,N_20360);
or U22047 (N_22047,N_21992,N_21860);
nand U22048 (N_22048,N_21660,N_21645);
or U22049 (N_22049,N_21149,N_20995);
and U22050 (N_22050,N_21720,N_20740);
nand U22051 (N_22051,N_21443,N_20583);
nand U22052 (N_22052,N_20468,N_21015);
nor U22053 (N_22053,N_20711,N_20478);
nand U22054 (N_22054,N_21844,N_21545);
nor U22055 (N_22055,N_21990,N_20197);
and U22056 (N_22056,N_21626,N_20262);
xnor U22057 (N_22057,N_21603,N_20978);
nor U22058 (N_22058,N_20074,N_20912);
or U22059 (N_22059,N_21869,N_20718);
nor U22060 (N_22060,N_20490,N_21047);
nor U22061 (N_22061,N_20225,N_21013);
nor U22062 (N_22062,N_21244,N_21780);
xnor U22063 (N_22063,N_20120,N_21417);
xor U22064 (N_22064,N_20517,N_21190);
xor U22065 (N_22065,N_21401,N_21111);
nand U22066 (N_22066,N_21738,N_21409);
nand U22067 (N_22067,N_20692,N_21837);
nand U22068 (N_22068,N_20345,N_20727);
or U22069 (N_22069,N_20050,N_20164);
and U22070 (N_22070,N_21043,N_21040);
nand U22071 (N_22071,N_20130,N_21381);
or U22072 (N_22072,N_20215,N_21759);
or U22073 (N_22073,N_21413,N_21317);
nor U22074 (N_22074,N_20513,N_21647);
or U22075 (N_22075,N_20709,N_20924);
xnor U22076 (N_22076,N_21796,N_21475);
xor U22077 (N_22077,N_21178,N_20884);
nand U22078 (N_22078,N_21812,N_20690);
xor U22079 (N_22079,N_21736,N_21156);
nand U22080 (N_22080,N_21734,N_20144);
nand U22081 (N_22081,N_21582,N_20726);
nand U22082 (N_22082,N_21173,N_21763);
nor U22083 (N_22083,N_20366,N_20605);
and U22084 (N_22084,N_21903,N_21511);
nand U22085 (N_22085,N_20454,N_20339);
nor U22086 (N_22086,N_20277,N_20194);
xor U22087 (N_22087,N_21224,N_20804);
xnor U22088 (N_22088,N_21839,N_21329);
or U22089 (N_22089,N_21082,N_21258);
nand U22090 (N_22090,N_21276,N_21599);
and U22091 (N_22091,N_20295,N_20968);
xor U22092 (N_22092,N_21819,N_21658);
or U22093 (N_22093,N_21942,N_21559);
nor U22094 (N_22094,N_21752,N_20160);
or U22095 (N_22095,N_21982,N_20302);
or U22096 (N_22096,N_21654,N_21530);
nor U22097 (N_22097,N_21899,N_20157);
nand U22098 (N_22098,N_20672,N_20211);
and U22099 (N_22099,N_21434,N_21697);
xnor U22100 (N_22100,N_20753,N_21053);
or U22101 (N_22101,N_20424,N_21447);
nand U22102 (N_22102,N_20864,N_20141);
and U22103 (N_22103,N_20934,N_20638);
nand U22104 (N_22104,N_20476,N_21026);
nor U22105 (N_22105,N_20300,N_21663);
or U22106 (N_22106,N_21744,N_20596);
or U22107 (N_22107,N_21066,N_21639);
nand U22108 (N_22108,N_20465,N_20380);
and U22109 (N_22109,N_20694,N_20683);
xnor U22110 (N_22110,N_21775,N_21680);
or U22111 (N_22111,N_21312,N_20081);
nand U22112 (N_22112,N_20955,N_21633);
and U22113 (N_22113,N_20571,N_20987);
xnor U22114 (N_22114,N_21863,N_21348);
nand U22115 (N_22115,N_21490,N_20041);
nor U22116 (N_22116,N_20407,N_20617);
nand U22117 (N_22117,N_20343,N_20106);
xor U22118 (N_22118,N_21277,N_20855);
and U22119 (N_22119,N_21466,N_21161);
or U22120 (N_22120,N_20415,N_20741);
or U22121 (N_22121,N_21056,N_20206);
nand U22122 (N_22122,N_21071,N_20228);
and U22123 (N_22123,N_20770,N_21890);
and U22124 (N_22124,N_20117,N_21773);
or U22125 (N_22125,N_21913,N_20124);
or U22126 (N_22126,N_20187,N_20058);
and U22127 (N_22127,N_20312,N_20422);
and U22128 (N_22128,N_20565,N_21833);
or U22129 (N_22129,N_21830,N_20592);
or U22130 (N_22130,N_21230,N_21172);
nor U22131 (N_22131,N_21701,N_21536);
and U22132 (N_22132,N_20385,N_20750);
nor U22133 (N_22133,N_21527,N_20561);
nand U22134 (N_22134,N_20636,N_20236);
and U22135 (N_22135,N_20042,N_21174);
nand U22136 (N_22136,N_21784,N_20706);
nor U22137 (N_22137,N_20989,N_20892);
and U22138 (N_22138,N_20336,N_21550);
and U22139 (N_22139,N_20326,N_21070);
or U22140 (N_22140,N_20649,N_21130);
xnor U22141 (N_22141,N_20357,N_21624);
nor U22142 (N_22142,N_20296,N_20745);
xor U22143 (N_22143,N_21587,N_21964);
nor U22144 (N_22144,N_20861,N_21044);
and U22145 (N_22145,N_20178,N_21045);
nor U22146 (N_22146,N_21325,N_20797);
and U22147 (N_22147,N_21506,N_21034);
nand U22148 (N_22148,N_20909,N_20051);
nor U22149 (N_22149,N_21105,N_21733);
nor U22150 (N_22150,N_20128,N_21181);
and U22151 (N_22151,N_21416,N_20434);
or U22152 (N_22152,N_20334,N_20545);
xor U22153 (N_22153,N_21858,N_20168);
or U22154 (N_22154,N_20414,N_21137);
or U22155 (N_22155,N_21923,N_21107);
nand U22156 (N_22156,N_20142,N_21922);
xor U22157 (N_22157,N_20504,N_21180);
nand U22158 (N_22158,N_20229,N_20281);
and U22159 (N_22159,N_20367,N_21275);
or U22160 (N_22160,N_21273,N_21169);
xnor U22161 (N_22161,N_20859,N_20405);
xnor U22162 (N_22162,N_20828,N_20274);
xnor U22163 (N_22163,N_21259,N_21248);
and U22164 (N_22164,N_21254,N_20642);
and U22165 (N_22165,N_20879,N_20309);
or U22166 (N_22166,N_21841,N_20010);
or U22167 (N_22167,N_21503,N_20933);
and U22168 (N_22168,N_20678,N_20096);
and U22169 (N_22169,N_21907,N_20568);
and U22170 (N_22170,N_20237,N_20446);
nor U22171 (N_22171,N_21743,N_20598);
nand U22172 (N_22172,N_21620,N_20553);
and U22173 (N_22173,N_20196,N_21065);
and U22174 (N_22174,N_20289,N_21309);
or U22175 (N_22175,N_20611,N_21742);
or U22176 (N_22176,N_21499,N_21129);
or U22177 (N_22177,N_20314,N_21287);
and U22178 (N_22178,N_20716,N_20410);
nand U22179 (N_22179,N_21679,N_21619);
and U22180 (N_22180,N_21621,N_21996);
and U22181 (N_22181,N_21748,N_20976);
nand U22182 (N_22182,N_21076,N_21184);
nand U22183 (N_22183,N_21338,N_21272);
nand U22184 (N_22184,N_21795,N_21449);
or U22185 (N_22185,N_20865,N_21753);
or U22186 (N_22186,N_20789,N_20285);
or U22187 (N_22187,N_21919,N_21410);
xor U22188 (N_22188,N_21954,N_21634);
xnor U22189 (N_22189,N_21198,N_20021);
or U22190 (N_22190,N_20391,N_20805);
xor U22191 (N_22191,N_21234,N_20084);
nor U22192 (N_22192,N_21048,N_21222);
nor U22193 (N_22193,N_20979,N_20313);
or U22194 (N_22194,N_20764,N_21054);
nand U22195 (N_22195,N_20844,N_21363);
xnor U22196 (N_22196,N_21332,N_20891);
nor U22197 (N_22197,N_21579,N_21193);
and U22198 (N_22198,N_21256,N_20355);
or U22199 (N_22199,N_21947,N_21114);
or U22200 (N_22200,N_20423,N_20751);
or U22201 (N_22201,N_21500,N_21788);
nor U22202 (N_22202,N_20994,N_20601);
nor U22203 (N_22203,N_20674,N_21086);
nand U22204 (N_22204,N_21699,N_21480);
and U22205 (N_22205,N_21087,N_21968);
xor U22206 (N_22206,N_20531,N_20658);
xor U22207 (N_22207,N_21873,N_21516);
or U22208 (N_22208,N_20755,N_21977);
and U22209 (N_22209,N_20484,N_21695);
nand U22210 (N_22210,N_20595,N_21625);
and U22211 (N_22211,N_20666,N_21077);
xor U22212 (N_22212,N_20547,N_21594);
nand U22213 (N_22213,N_21959,N_20869);
nand U22214 (N_22214,N_21762,N_20620);
and U22215 (N_22215,N_20433,N_20623);
xnor U22216 (N_22216,N_21975,N_20267);
or U22217 (N_22217,N_20093,N_20455);
or U22218 (N_22218,N_20969,N_20724);
xnor U22219 (N_22219,N_20831,N_21152);
nor U22220 (N_22220,N_21867,N_21084);
and U22221 (N_22221,N_20846,N_20839);
or U22222 (N_22222,N_21909,N_21316);
nand U22223 (N_22223,N_20812,N_20299);
or U22224 (N_22224,N_21378,N_21931);
nor U22225 (N_22225,N_21285,N_20223);
xor U22226 (N_22226,N_21567,N_20039);
and U22227 (N_22227,N_21676,N_20953);
or U22228 (N_22228,N_21106,N_21019);
xnor U22229 (N_22229,N_21556,N_20556);
or U22230 (N_22230,N_20960,N_21974);
nor U22231 (N_22231,N_21962,N_21607);
nand U22232 (N_22232,N_21037,N_21457);
and U22233 (N_22233,N_20973,N_20038);
or U22234 (N_22234,N_20033,N_20681);
and U22235 (N_22235,N_20192,N_20310);
or U22236 (N_22236,N_20108,N_21758);
nand U22237 (N_22237,N_21573,N_21143);
nand U22238 (N_22238,N_20136,N_20721);
xor U22239 (N_22239,N_20972,N_20354);
nand U22240 (N_22240,N_20659,N_21713);
nor U22241 (N_22241,N_20624,N_20537);
and U22242 (N_22242,N_21572,N_21108);
nand U22243 (N_22243,N_21912,N_20503);
xor U22244 (N_22244,N_20358,N_21425);
nand U22245 (N_22245,N_21472,N_20006);
and U22246 (N_22246,N_21007,N_20169);
xnor U22247 (N_22247,N_21249,N_21659);
and U22248 (N_22248,N_21687,N_21896);
or U22249 (N_22249,N_21618,N_21666);
nor U22250 (N_22250,N_21214,N_20102);
nor U22251 (N_22251,N_21051,N_20280);
and U22252 (N_22252,N_20947,N_21269);
xnor U22253 (N_22253,N_20510,N_21100);
or U22254 (N_22254,N_21395,N_20167);
nand U22255 (N_22255,N_20146,N_21350);
xnor U22256 (N_22256,N_21884,N_21940);
nor U22257 (N_22257,N_21081,N_20383);
nor U22258 (N_22258,N_20325,N_21104);
xnor U22259 (N_22259,N_21392,N_21703);
nor U22260 (N_22260,N_20431,N_21941);
nand U22261 (N_22261,N_21757,N_20137);
nor U22262 (N_22262,N_21589,N_21652);
nand U22263 (N_22263,N_21935,N_21386);
or U22264 (N_22264,N_20458,N_20818);
nor U22265 (N_22265,N_20991,N_21630);
and U22266 (N_22266,N_21123,N_20677);
nand U22267 (N_22267,N_21908,N_20737);
xor U22268 (N_22268,N_20785,N_20303);
nor U22269 (N_22269,N_21283,N_20264);
xor U22270 (N_22270,N_20799,N_20212);
and U22271 (N_22271,N_21300,N_20775);
nor U22272 (N_22272,N_20204,N_21134);
nor U22273 (N_22273,N_20530,N_21781);
nor U22274 (N_22274,N_21829,N_21255);
nand U22275 (N_22275,N_21640,N_21548);
and U22276 (N_22276,N_20066,N_20511);
and U22277 (N_22277,N_20263,N_20809);
and U22278 (N_22278,N_21291,N_21356);
nor U22279 (N_22279,N_21646,N_20272);
nand U22280 (N_22280,N_20372,N_21939);
nand U22281 (N_22281,N_21167,N_20044);
and U22282 (N_22282,N_20068,N_20341);
nor U22283 (N_22283,N_20445,N_20221);
or U22284 (N_22284,N_20214,N_20885);
or U22285 (N_22285,N_20413,N_21999);
nor U22286 (N_22286,N_21677,N_20240);
and U22287 (N_22287,N_21280,N_20579);
and U22288 (N_22288,N_21187,N_21967);
nor U22289 (N_22289,N_21011,N_20962);
and U22290 (N_22290,N_21446,N_21813);
nand U22291 (N_22291,N_21750,N_21253);
and U22292 (N_22292,N_20645,N_20493);
and U22293 (N_22293,N_21557,N_21286);
nand U22294 (N_22294,N_20700,N_20937);
or U22295 (N_22295,N_21186,N_20868);
xor U22296 (N_22296,N_20246,N_21430);
or U22297 (N_22297,N_20790,N_21008);
nor U22298 (N_22298,N_21073,N_21802);
nand U22299 (N_22299,N_21487,N_21808);
xnor U22300 (N_22300,N_20535,N_20860);
nor U22301 (N_22301,N_20047,N_21655);
and U22302 (N_22302,N_20779,N_21554);
nand U22303 (N_22303,N_20733,N_20539);
and U22304 (N_22304,N_20092,N_21611);
and U22305 (N_22305,N_20080,N_21668);
or U22306 (N_22306,N_20279,N_21577);
and U22307 (N_22307,N_20111,N_21811);
or U22308 (N_22308,N_20083,N_21433);
and U22309 (N_22309,N_20725,N_20852);
or U22310 (N_22310,N_20963,N_21661);
nor U22311 (N_22311,N_20350,N_20417);
nor U22312 (N_22312,N_21158,N_20575);
xor U22313 (N_22313,N_21140,N_20640);
nand U22314 (N_22314,N_20331,N_20235);
xor U22315 (N_22315,N_20710,N_20232);
nand U22316 (N_22316,N_20479,N_21689);
or U22317 (N_22317,N_20650,N_21882);
xnor U22318 (N_22318,N_20340,N_20249);
nand U22319 (N_22319,N_21918,N_21848);
nor U22320 (N_22320,N_21876,N_20135);
and U22321 (N_22321,N_20996,N_21617);
and U22322 (N_22322,N_20201,N_21385);
xnor U22323 (N_22323,N_21016,N_20125);
and U22324 (N_22324,N_20425,N_21154);
and U22325 (N_22325,N_20820,N_21023);
nand U22326 (N_22326,N_20882,N_21731);
and U22327 (N_22327,N_21060,N_20481);
xnor U22328 (N_22328,N_20532,N_20941);
and U22329 (N_22329,N_20802,N_20398);
and U22330 (N_22330,N_20505,N_21519);
and U22331 (N_22331,N_21473,N_20474);
nor U22332 (N_22332,N_21649,N_20895);
and U22333 (N_22333,N_20762,N_20628);
nor U22334 (N_22334,N_21980,N_21109);
and U22335 (N_22335,N_20631,N_21431);
or U22336 (N_22336,N_21423,N_20563);
or U22337 (N_22337,N_21928,N_21985);
nand U22338 (N_22338,N_21892,N_21801);
or U22339 (N_22339,N_21235,N_21691);
xor U22340 (N_22340,N_20825,N_20848);
or U22341 (N_22341,N_20217,N_21301);
nor U22342 (N_22342,N_20369,N_20477);
or U22343 (N_22343,N_21814,N_20104);
nand U22344 (N_22344,N_21525,N_20959);
nor U22345 (N_22345,N_21274,N_21710);
and U22346 (N_22346,N_21644,N_21906);
or U22347 (N_22347,N_21384,N_21210);
nor U22348 (N_22348,N_21307,N_21776);
nand U22349 (N_22349,N_20669,N_20986);
and U22350 (N_22350,N_20931,N_20463);
nor U22351 (N_22351,N_21756,N_20002);
or U22352 (N_22352,N_20412,N_20456);
and U22353 (N_22353,N_20705,N_21493);
or U22354 (N_22354,N_21783,N_21354);
nor U22355 (N_22355,N_20387,N_21901);
nor U22356 (N_22356,N_21200,N_21747);
nor U22357 (N_22357,N_21546,N_21604);
nand U22358 (N_22358,N_21001,N_21845);
or U22359 (N_22359,N_20319,N_20119);
and U22360 (N_22360,N_21709,N_21563);
nand U22361 (N_22361,N_20956,N_21289);
nor U22362 (N_22362,N_21509,N_21215);
nand U22363 (N_22363,N_21597,N_20379);
and U22364 (N_22364,N_20794,N_21492);
and U22365 (N_22365,N_20181,N_20625);
or U22366 (N_22366,N_21674,N_21010);
and U22367 (N_22367,N_21886,N_20573);
nor U22368 (N_22368,N_21675,N_20787);
and U22369 (N_22369,N_20682,N_21196);
nor U22370 (N_22370,N_21049,N_20247);
and U22371 (N_22371,N_20430,N_20554);
nand U22372 (N_22372,N_20524,N_21406);
nand U22373 (N_22373,N_20166,N_20305);
or U22374 (N_22374,N_20853,N_21791);
nand U22375 (N_22375,N_21826,N_20712);
xnor U22376 (N_22376,N_20306,N_21712);
xnor U22377 (N_22377,N_20622,N_21435);
xnor U22378 (N_22378,N_20233,N_21110);
nor U22379 (N_22379,N_20329,N_20282);
and U22380 (N_22380,N_20534,N_21238);
xnor U22381 (N_22381,N_20159,N_21221);
or U22382 (N_22382,N_20843,N_21426);
or U22383 (N_22383,N_20905,N_21442);
nand U22384 (N_22384,N_20739,N_20644);
nor U22385 (N_22385,N_21566,N_20662);
and U22386 (N_22386,N_21857,N_21916);
nor U22387 (N_22387,N_20046,N_21292);
nor U22388 (N_22388,N_20632,N_20227);
or U22389 (N_22389,N_21456,N_20087);
nor U22390 (N_22390,N_20992,N_21335);
nor U22391 (N_22391,N_20555,N_21495);
nand U22392 (N_22392,N_20985,N_21068);
or U22393 (N_22393,N_21501,N_21393);
and U22394 (N_22394,N_20113,N_21586);
or U22395 (N_22395,N_20834,N_21765);
or U22396 (N_22396,N_20754,N_20833);
nor U22397 (N_22397,N_20795,N_20664);
or U22398 (N_22398,N_21966,N_21798);
xnor U22399 (N_22399,N_20003,N_20471);
and U22400 (N_22400,N_21685,N_21148);
xor U22401 (N_22401,N_20069,N_21127);
and U22402 (N_22402,N_21721,N_21271);
nor U22403 (N_22403,N_20722,N_20293);
or U22404 (N_22404,N_20287,N_20439);
xnor U22405 (N_22405,N_21018,N_20461);
and U22406 (N_22406,N_21041,N_21766);
xor U22407 (N_22407,N_20701,N_21672);
xor U22408 (N_22408,N_21868,N_20320);
nor U22409 (N_22409,N_21090,N_21671);
nor U22410 (N_22410,N_20988,N_21998);
nor U22411 (N_22411,N_20406,N_21203);
nand U22412 (N_22412,N_21092,N_20470);
xnor U22413 (N_22413,N_21000,N_20308);
and U22414 (N_22414,N_21061,N_21079);
xor U22415 (N_22415,N_21543,N_21310);
nor U22416 (N_22416,N_21290,N_21465);
nor U22417 (N_22417,N_20115,N_20656);
and U22418 (N_22418,N_20297,N_20378);
nor U22419 (N_22419,N_20550,N_21165);
and U22420 (N_22420,N_21028,N_20349);
and U22421 (N_22421,N_21881,N_21164);
nand U22422 (N_22422,N_21263,N_21505);
nor U22423 (N_22423,N_21268,N_20452);
nand U22424 (N_22424,N_20184,N_21328);
and U22425 (N_22425,N_21136,N_20543);
nand U22426 (N_22426,N_20043,N_20715);
nor U22427 (N_22427,N_21002,N_21097);
xor U22428 (N_22428,N_20127,N_21827);
nor U22429 (N_22429,N_20457,N_21714);
or U22430 (N_22430,N_20728,N_21265);
or U22431 (N_22431,N_20390,N_20460);
nor U22432 (N_22432,N_20742,N_21179);
xnor U22433 (N_22433,N_21231,N_20506);
xor U22434 (N_22434,N_20266,N_21339);
nor U22435 (N_22435,N_20091,N_21581);
nand U22436 (N_22436,N_21855,N_20679);
nor U22437 (N_22437,N_20210,N_20518);
nor U22438 (N_22438,N_20149,N_21612);
nand U22439 (N_22439,N_20732,N_20777);
xor U22440 (N_22440,N_21202,N_21851);
and U22441 (N_22441,N_21334,N_21828);
nand U22442 (N_22442,N_20730,N_20708);
and U22443 (N_22443,N_20005,N_21306);
nand U22444 (N_22444,N_20322,N_20451);
or U22445 (N_22445,N_21128,N_21119);
and U22446 (N_22446,N_20850,N_21877);
nor U22447 (N_22447,N_20064,N_21570);
xnor U22448 (N_22448,N_20784,N_20330);
nor U22449 (N_22449,N_21146,N_21243);
and U22450 (N_22450,N_20324,N_20667);
nor U22451 (N_22451,N_21004,N_20001);
xor U22452 (N_22452,N_21029,N_21379);
nand U22453 (N_22453,N_21022,N_20065);
or U22454 (N_22454,N_20347,N_21021);
and U22455 (N_22455,N_21514,N_20560);
xor U22456 (N_22456,N_20362,N_20593);
xor U22457 (N_22457,N_20371,N_21949);
and U22458 (N_22458,N_20665,N_20195);
or U22459 (N_22459,N_21321,N_20781);
xor U22460 (N_22460,N_20940,N_20255);
or U22461 (N_22461,N_21643,N_21264);
or U22462 (N_22462,N_21803,N_20791);
or U22463 (N_22463,N_20218,N_20085);
and U22464 (N_22464,N_21656,N_21590);
or U22465 (N_22465,N_20760,N_21834);
or U22466 (N_22466,N_21904,N_21562);
xnor U22467 (N_22467,N_21117,N_20304);
xnor U22468 (N_22468,N_21217,N_21298);
and U22469 (N_22469,N_21358,N_20494);
or U22470 (N_22470,N_21778,N_20581);
nand U22471 (N_22471,N_21101,N_21411);
or U22472 (N_22472,N_21741,N_20007);
and U22473 (N_22473,N_21664,N_20244);
or U22474 (N_22474,N_21177,N_20473);
nand U22475 (N_22475,N_20749,N_20746);
and U22476 (N_22476,N_21580,N_20231);
or U22477 (N_22477,N_20351,N_21088);
nand U22478 (N_22478,N_21318,N_20586);
or U22479 (N_22479,N_20170,N_20911);
and U22480 (N_22480,N_21591,N_20441);
nand U22481 (N_22481,N_20438,N_20926);
or U22482 (N_22482,N_20714,N_20793);
nor U22483 (N_22483,N_21870,N_21461);
and U22484 (N_22484,N_20022,N_21326);
and U22485 (N_22485,N_20747,N_20333);
nand U22486 (N_22486,N_21723,N_20881);
and U22487 (N_22487,N_21915,N_21498);
nor U22488 (N_22488,N_20134,N_20821);
nor U22489 (N_22489,N_20492,N_21629);
and U22490 (N_22490,N_21478,N_20874);
or U22491 (N_22491,N_21208,N_20459);
nor U22492 (N_22492,N_21199,N_21296);
and U22493 (N_22493,N_20079,N_20888);
or U22494 (N_22494,N_20158,N_21937);
nor U22495 (N_22495,N_20938,N_20501);
xor U22496 (N_22496,N_21653,N_21311);
xnor U22497 (N_22497,N_20687,N_20743);
and U22498 (N_22498,N_20110,N_20014);
or U22499 (N_22499,N_20190,N_21902);
or U22500 (N_22500,N_20939,N_20637);
or U22501 (N_22501,N_21031,N_20582);
nand U22502 (N_22502,N_21544,N_21820);
nor U22503 (N_22503,N_20857,N_21491);
and U22504 (N_22504,N_21799,N_20090);
nor U22505 (N_22505,N_21175,N_21840);
or U22506 (N_22506,N_20562,N_21642);
nand U22507 (N_22507,N_20419,N_20020);
xor U22508 (N_22508,N_21122,N_21614);
xnor U22509 (N_22509,N_20162,N_20382);
or U22510 (N_22510,N_20639,N_20498);
nand U22511 (N_22511,N_21365,N_21227);
nor U22512 (N_22512,N_20188,N_20719);
and U22513 (N_22513,N_20619,N_20612);
xnor U22514 (N_22514,N_21341,N_20958);
and U22515 (N_22515,N_21872,N_20353);
and U22516 (N_22516,N_21821,N_20551);
nor U22517 (N_22517,N_20207,N_20591);
nor U22518 (N_22518,N_20851,N_20948);
and U22519 (N_22519,N_21232,N_21602);
nor U22520 (N_22520,N_20177,N_20557);
xor U22521 (N_22521,N_20328,N_20578);
xnor U22522 (N_22522,N_21189,N_20408);
or U22523 (N_22523,N_20840,N_20954);
and U22524 (N_22524,N_20915,N_20147);
or U22525 (N_22525,N_20736,N_21787);
or U22526 (N_22526,N_21694,N_21706);
and U22527 (N_22527,N_21440,N_20898);
xnor U22528 (N_22528,N_21972,N_21046);
nand U22529 (N_22529,N_21481,N_20870);
or U22530 (N_22530,N_21692,N_21971);
nor U22531 (N_22531,N_20604,N_21063);
nand U22532 (N_22532,N_21252,N_21984);
and U22533 (N_22533,N_20290,N_21850);
nand U22534 (N_22534,N_21349,N_20219);
nor U22535 (N_22535,N_21578,N_20862);
nand U22536 (N_22536,N_20768,N_20587);
or U22537 (N_22537,N_21856,N_20925);
or U22538 (N_22538,N_20913,N_20359);
xor U22539 (N_22539,N_21297,N_20698);
nand U22540 (N_22540,N_21118,N_21838);
nand U22541 (N_22541,N_21774,N_20572);
xnor U22542 (N_22542,N_21183,N_21219);
xnor U22543 (N_22543,N_21973,N_20000);
nand U22544 (N_22544,N_21785,N_20153);
nand U22545 (N_22545,N_20783,N_21623);
nor U22546 (N_22546,N_20981,N_20089);
xnor U22547 (N_22547,N_20935,N_21267);
xor U22548 (N_22548,N_21360,N_21375);
or U22549 (N_22549,N_21294,N_21359);
or U22550 (N_22550,N_20151,N_21569);
nor U22551 (N_22551,N_20696,N_20226);
or U22552 (N_22552,N_21236,N_20030);
nor U22553 (N_22553,N_21583,N_21135);
nand U22554 (N_22554,N_21005,N_20552);
and U22555 (N_22555,N_20176,N_21025);
nand U22556 (N_22556,N_20606,N_21042);
nor U22557 (N_22557,N_21057,N_21800);
xor U22558 (N_22558,N_20140,N_21979);
xnor U22559 (N_22559,N_21943,N_21665);
and U22560 (N_22560,N_20138,N_20752);
or U22561 (N_22561,N_21512,N_20590);
nor U22562 (N_22562,N_21476,N_20024);
nand U22563 (N_22563,N_21989,N_20670);
and U22564 (N_22564,N_21729,N_21997);
xor U22565 (N_22565,N_21313,N_20602);
nor U22566 (N_22566,N_21324,N_20114);
and U22567 (N_22567,N_21831,N_20999);
nor U22568 (N_22568,N_21606,N_21960);
nand U22569 (N_22569,N_21616,N_20165);
and U22570 (N_22570,N_20199,N_20835);
and U22571 (N_22571,N_20105,N_20693);
nor U22572 (N_22572,N_21887,N_21024);
and U22573 (N_22573,N_21058,N_20922);
xor U22574 (N_22574,N_20899,N_20971);
nor U22575 (N_22575,N_20529,N_20254);
nand U22576 (N_22576,N_20808,N_20919);
xor U22577 (N_22577,N_21344,N_21418);
and U22578 (N_22578,N_20483,N_21969);
xor U22579 (N_22579,N_21864,N_20538);
xnor U22580 (N_22580,N_21718,N_20923);
xnor U22581 (N_22581,N_21861,N_21247);
or U22582 (N_22582,N_21779,N_20546);
and U22583 (N_22583,N_21510,N_20118);
or U22584 (N_22584,N_20873,N_20758);
or U22585 (N_22585,N_20403,N_21155);
nand U22586 (N_22586,N_21322,N_21362);
nand U22587 (N_22587,N_21717,N_21207);
and U22588 (N_22588,N_20914,N_20467);
and U22589 (N_22589,N_20773,N_20819);
xor U22590 (N_22590,N_20863,N_21059);
or U22591 (N_22591,N_20965,N_20107);
nand U22592 (N_22592,N_20542,N_20876);
and U22593 (N_22593,N_21412,N_20549);
xor U22594 (N_22594,N_21213,N_21529);
nand U22595 (N_22595,N_20763,N_21163);
xnor U22596 (N_22596,N_21853,N_20866);
nand U22597 (N_22597,N_21030,N_20327);
xor U22598 (N_22598,N_21981,N_21995);
or U22599 (N_22599,N_21551,N_20436);
and U22600 (N_22600,N_21879,N_20998);
and U22601 (N_22601,N_21865,N_20364);
and U22602 (N_22602,N_20209,N_20920);
or U22603 (N_22603,N_21535,N_21205);
or U22604 (N_22604,N_20824,N_21955);
and U22605 (N_22605,N_20286,N_21842);
xnor U22606 (N_22606,N_20661,N_21852);
xor U22607 (N_22607,N_20420,N_21683);
nand U22608 (N_22608,N_20376,N_20769);
xor U22609 (N_22609,N_21216,N_20886);
nor U22610 (N_22610,N_20268,N_20009);
xnor U22611 (N_22611,N_20641,N_20256);
nand U22612 (N_22612,N_21737,N_21120);
nand U22613 (N_22613,N_21926,N_20200);
and U22614 (N_22614,N_20018,N_21726);
nor U22615 (N_22615,N_20577,N_21673);
nor U22616 (N_22616,N_20276,N_21330);
nor U22617 (N_22617,N_20528,N_21033);
xor U22618 (N_22618,N_21315,N_20896);
xnor U22619 (N_22619,N_21415,N_21407);
or U22620 (N_22620,N_21399,N_20186);
nand U22621 (N_22621,N_20772,N_20045);
or U22622 (N_22622,N_20713,N_20004);
nor U22623 (N_22623,N_20273,N_21223);
or U22624 (N_22624,N_20977,N_21761);
nand U22625 (N_22625,N_21702,N_20652);
or U22626 (N_22626,N_21809,N_20123);
nand U22627 (N_22627,N_21270,N_20163);
or U22628 (N_22628,N_21956,N_20813);
nor U22629 (N_22629,N_20224,N_20055);
and U22630 (N_22630,N_20208,N_20780);
nor U22631 (N_22631,N_21976,N_21874);
or U22632 (N_22632,N_21866,N_21728);
or U22633 (N_22633,N_21133,N_20589);
nor U22634 (N_22634,N_21421,N_20475);
xnor U22635 (N_22635,N_21441,N_21835);
nand U22636 (N_22636,N_21383,N_21320);
nand U22637 (N_22637,N_21893,N_20830);
or U22638 (N_22638,N_20704,N_21735);
and U22639 (N_22639,N_20626,N_20967);
nor U22640 (N_22640,N_20175,N_20502);
and U22641 (N_22641,N_20395,N_20527);
and U22642 (N_22642,N_21439,N_21637);
nor U22643 (N_22643,N_21934,N_20827);
or U22644 (N_22644,N_20512,N_21014);
nand U22645 (N_22645,N_20121,N_20849);
nand U22646 (N_22646,N_21055,N_21112);
nand U22647 (N_22647,N_20031,N_20983);
and U22648 (N_22648,N_21983,N_20832);
nor U22649 (N_22649,N_21933,N_20767);
nor U22650 (N_22650,N_20259,N_20782);
xnor U22651 (N_22651,N_21518,N_20759);
xor U22652 (N_22652,N_20615,N_20990);
and U22653 (N_22653,N_20040,N_20056);
or U22654 (N_22654,N_21124,N_21131);
xnor U22655 (N_22655,N_21182,N_20396);
nand U22656 (N_22656,N_21085,N_21367);
or U22657 (N_22657,N_21372,N_21513);
nor U22658 (N_22658,N_21126,N_21751);
nand U22659 (N_22659,N_21398,N_21078);
nand U22660 (N_22660,N_20630,N_20970);
nor U22661 (N_22661,N_20062,N_20078);
nor U22662 (N_22662,N_21732,N_21067);
nand U22663 (N_22663,N_21534,N_20388);
xnor U22664 (N_22664,N_20444,N_21062);
xor U22665 (N_22665,N_21825,N_20389);
xnor U22666 (N_22666,N_21246,N_21805);
nor U22667 (N_22667,N_20766,N_20654);
and U22668 (N_22668,N_20703,N_20216);
nand U22669 (N_22669,N_20500,N_21507);
and U22670 (N_22670,N_20317,N_21790);
nor U22671 (N_22671,N_20903,N_20173);
and U22672 (N_22672,N_21782,N_20771);
and U22673 (N_22673,N_21540,N_20875);
or U22674 (N_22674,N_20633,N_21032);
nor U22675 (N_22675,N_21308,N_20801);
nor U22676 (N_22676,N_21584,N_21818);
and U22677 (N_22677,N_20867,N_20570);
xnor U22678 (N_22678,N_20800,N_21470);
nand U22679 (N_22679,N_21965,N_21693);
nor U22680 (N_22680,N_20668,N_21952);
nor U22681 (N_22681,N_21303,N_21613);
nor U22682 (N_22682,N_20097,N_21789);
xor U22683 (N_22683,N_20883,N_20100);
xnor U22684 (N_22684,N_20318,N_20365);
and U22685 (N_22685,N_21553,N_20129);
and U22686 (N_22686,N_21396,N_20348);
nand U22687 (N_22687,N_21257,N_20480);
xor U22688 (N_22688,N_20872,N_21388);
xor U22689 (N_22689,N_21552,N_20516);
or U22690 (N_22690,N_20161,N_20342);
nor U22691 (N_22691,N_20103,N_20323);
or U22692 (N_22692,N_21871,N_21600);
xor U22693 (N_22693,N_21957,N_21592);
xor U22694 (N_22694,N_20250,N_21488);
nor U22695 (N_22695,N_21373,N_21075);
xnor U22696 (N_22696,N_21400,N_21369);
nand U22697 (N_22697,N_20028,N_20540);
nand U22698 (N_22698,N_20026,N_20648);
nor U22699 (N_22699,N_20368,N_20921);
or U22700 (N_22700,N_21382,N_21323);
nand U22701 (N_22701,N_21444,N_20185);
or U22702 (N_22702,N_20806,N_20495);
nand U22703 (N_22703,N_20116,N_21987);
nor U22704 (N_22704,N_20964,N_21069);
nor U22705 (N_22705,N_21794,N_21116);
and U22706 (N_22706,N_21724,N_21849);
xor U22707 (N_22707,N_21686,N_21970);
and U22708 (N_22708,N_20811,N_20269);
nand U22709 (N_22709,N_20150,N_21098);
and U22710 (N_22710,N_21250,N_21351);
nor U22711 (N_22711,N_21740,N_20569);
or U22712 (N_22712,N_21883,N_21404);
xnor U22713 (N_22713,N_20627,N_20798);
nand U22714 (N_22714,N_20520,N_21160);
nor U22715 (N_22715,N_21027,N_20858);
or U22716 (N_22716,N_20691,N_20786);
nor U22717 (N_22717,N_21451,N_20384);
nand U22718 (N_22718,N_20897,N_21547);
nor U22719 (N_22719,N_21854,N_21772);
or U22720 (N_22720,N_21394,N_21428);
or U22721 (N_22721,N_21538,N_20695);
nor U22722 (N_22722,N_21555,N_21093);
nand U22723 (N_22723,N_20507,N_21453);
nand U22724 (N_22724,N_20496,N_21333);
nor U22725 (N_22725,N_20723,N_20966);
nor U22726 (N_22726,N_20462,N_21508);
nor U22727 (N_22727,N_21945,N_21991);
xnor U22728 (N_22728,N_21862,N_20491);
xor U22729 (N_22729,N_20257,N_20241);
and U22730 (N_22730,N_20499,N_21485);
nor U22731 (N_22731,N_20126,N_20437);
nor U22732 (N_22732,N_21727,N_21191);
xor U22733 (N_22733,N_20449,N_20916);
or U22734 (N_22734,N_21064,N_20567);
and U22735 (N_22735,N_21793,N_21337);
and U22736 (N_22736,N_21176,N_20440);
or U22737 (N_22737,N_21459,N_21094);
and U22738 (N_22738,N_20894,N_20796);
nor U22739 (N_22739,N_20077,N_20344);
and U22740 (N_22740,N_20680,N_21598);
and U22741 (N_22741,N_20699,N_21667);
or U22742 (N_22742,N_20984,N_21424);
nand U22743 (N_22743,N_21806,N_21035);
nand U22744 (N_22744,N_21113,N_20526);
and U22745 (N_22745,N_21483,N_20675);
xor U22746 (N_22746,N_20974,N_20576);
nor U22747 (N_22747,N_20222,N_20816);
xnor U22748 (N_22748,N_21786,N_21458);
nor U22749 (N_22749,N_21427,N_20332);
nand U22750 (N_22750,N_20432,N_21142);
and U22751 (N_22751,N_20657,N_20734);
nand U22752 (N_22752,N_21353,N_20242);
xor U22753 (N_22753,N_20610,N_21549);
nor U22754 (N_22754,N_20301,N_20871);
xor U22755 (N_22755,N_20735,N_21627);
nand U22756 (N_22756,N_20778,N_21610);
xor U22757 (N_22757,N_20183,N_20174);
nand U22758 (N_22758,N_21542,N_20075);
and U22759 (N_22759,N_21824,N_20307);
nand U22760 (N_22760,N_21342,N_21102);
nand U22761 (N_22761,N_21494,N_21847);
nor U22762 (N_22762,N_20541,N_21463);
xor U22763 (N_22763,N_20019,N_20316);
and U22764 (N_22764,N_21293,N_21132);
and U22765 (N_22765,N_20243,N_21020);
and U22766 (N_22766,N_20377,N_21419);
xor U22767 (N_22767,N_20603,N_20635);
or U22768 (N_22768,N_20101,N_20270);
nand U22769 (N_22769,N_21361,N_20838);
nand U22770 (N_22770,N_20370,N_21888);
xor U22771 (N_22771,N_21924,N_20205);
xor U22772 (N_22772,N_21823,N_20487);
and U22773 (N_22773,N_21497,N_20321);
and U22774 (N_22774,N_21588,N_21944);
and U22775 (N_22775,N_20847,N_21910);
nor U22776 (N_22776,N_20822,N_21305);
and U22777 (N_22777,N_21938,N_20676);
nand U22778 (N_22778,N_21402,N_20880);
nand U22779 (N_22779,N_21914,N_20514);
xor U22780 (N_22780,N_21719,N_20902);
xor U22781 (N_22781,N_21920,N_20584);
xnor U22782 (N_22782,N_20271,N_20035);
nand U22783 (N_22783,N_20774,N_21988);
or U22784 (N_22784,N_21917,N_21632);
and U22785 (N_22785,N_20234,N_20993);
xor U22786 (N_22786,N_20122,N_20616);
xnor U22787 (N_22787,N_20180,N_20363);
or U22788 (N_22788,N_21897,N_21096);
nor U22789 (N_22789,N_20469,N_21171);
and U22790 (N_22790,N_21080,N_20489);
or U22791 (N_22791,N_21651,N_21436);
xnor U22792 (N_22792,N_21138,N_21448);
or U22793 (N_22793,N_20792,N_21374);
nor U22794 (N_22794,N_21698,N_20519);
and U22795 (N_22795,N_21815,N_20057);
nor U22796 (N_22796,N_21229,N_21150);
xor U22797 (N_22797,N_21141,N_20094);
and U22798 (N_22798,N_20427,N_21523);
nand U22799 (N_22799,N_20008,N_21745);
nor U22800 (N_22800,N_20193,N_20829);
nand U22801 (N_22801,N_21635,N_21777);
xor U22802 (N_22802,N_21768,N_20744);
nand U22803 (N_22803,N_21958,N_21978);
or U22804 (N_22804,N_20453,N_21345);
and U22805 (N_22805,N_20663,N_21211);
and U22806 (N_22806,N_21445,N_20418);
or U22807 (N_22807,N_20284,N_20944);
xor U22808 (N_22808,N_21524,N_21585);
xor U22809 (N_22809,N_21299,N_21304);
nor U22810 (N_22810,N_21605,N_20564);
nor U22811 (N_22811,N_20386,N_20037);
nand U22812 (N_22812,N_20609,N_20076);
and U22813 (N_22813,N_21539,N_21352);
nor U22814 (N_22814,N_20908,N_21464);
or U22815 (N_22815,N_21467,N_20945);
or U22816 (N_22816,N_20607,N_20435);
xnor U22817 (N_22817,N_21357,N_21397);
or U22818 (N_22818,N_21099,N_21260);
xor U22819 (N_22819,N_20155,N_21245);
or U22820 (N_22820,N_20073,N_20088);
xnor U22821 (N_22821,N_20025,N_21159);
or U22822 (N_22822,N_21930,N_20337);
and U22823 (N_22823,N_20261,N_21380);
nand U22824 (N_22824,N_20877,N_21389);
nor U22825 (N_22825,N_20172,N_21678);
and U22826 (N_22826,N_21681,N_20932);
nor U22827 (N_22827,N_20515,N_20260);
or U22828 (N_22828,N_21739,N_21608);
xnor U22829 (N_22829,N_20071,N_20684);
or U22830 (N_22830,N_21218,N_21331);
xnor U22831 (N_22831,N_21204,N_20810);
or U22832 (N_22832,N_21371,N_21262);
nand U22833 (N_22833,N_21880,N_20023);
nor U22834 (N_22834,N_20900,N_21194);
nand U22835 (N_22835,N_20761,N_20011);
nor U22836 (N_22836,N_21638,N_21905);
nand U22837 (N_22837,N_20957,N_20653);
nor U22838 (N_22838,N_21012,N_20952);
xnor U22839 (N_22839,N_21859,N_20239);
or U22840 (N_22840,N_20060,N_20063);
or U22841 (N_22841,N_20521,N_20803);
nor U22842 (N_22842,N_21145,N_20508);
and U22843 (N_22843,N_21284,N_21596);
nand U22844 (N_22844,N_20283,N_21121);
nor U22845 (N_22845,N_20689,N_21891);
or U22846 (N_22846,N_20673,N_20189);
xnor U22847 (N_22847,N_21036,N_21528);
and U22848 (N_22848,N_21366,N_20887);
nor U22849 (N_22849,N_21560,N_21089);
nand U22850 (N_22850,N_21700,N_21471);
xnor U22851 (N_22851,N_21192,N_21708);
or U22852 (N_22852,N_20671,N_20765);
xnor U22853 (N_22853,N_21622,N_20485);
or U22854 (N_22854,N_20145,N_21072);
or U22855 (N_22855,N_21875,N_20497);
nor U22856 (N_22856,N_21894,N_21166);
nor U22857 (N_22857,N_21770,N_21816);
nand U22858 (N_22858,N_21688,N_21911);
nand U22859 (N_22859,N_21746,N_21239);
and U22860 (N_22860,N_21486,N_20132);
and U22861 (N_22861,N_21504,N_20686);
or U22862 (N_22862,N_20613,N_21095);
nand U22863 (N_22863,N_21355,N_21390);
nand U22864 (N_22864,N_21185,N_20930);
and U22865 (N_22865,N_21188,N_21468);
nand U22866 (N_22866,N_21950,N_20685);
xor U22867 (N_22867,N_20082,N_20220);
nor U22868 (N_22868,N_21474,N_21561);
nand U22869 (N_22869,N_21197,N_20904);
nor U22870 (N_22870,N_20402,N_21725);
nand U22871 (N_22871,N_21368,N_21314);
nand U22872 (N_22872,N_20548,N_20013);
nand U22873 (N_22873,N_20566,N_21575);
nor U22874 (N_22874,N_20448,N_20643);
nand U22875 (N_22875,N_21462,N_20447);
or U22876 (N_22876,N_20942,N_20245);
nor U22877 (N_22877,N_20982,N_21225);
nor U22878 (N_22878,N_21730,N_20717);
nand U22879 (N_22879,N_20248,N_20599);
and U22880 (N_22880,N_21749,N_21206);
xnor U22881 (N_22881,N_20143,N_20156);
nor U22882 (N_22882,N_20597,N_20027);
or U22883 (N_22883,N_20352,N_21288);
and U22884 (N_22884,N_21103,N_20651);
nand U22885 (N_22885,N_21115,N_21279);
xor U22886 (N_22886,N_21502,N_21564);
xor U22887 (N_22887,N_21233,N_20585);
nand U22888 (N_22888,N_20392,N_20906);
or U22889 (N_22889,N_21281,N_20776);
nor U22890 (N_22890,N_21568,N_20252);
and U22891 (N_22891,N_21377,N_21986);
xnor U22892 (N_22892,N_20660,N_20910);
or U22893 (N_22893,N_20017,N_21767);
nor U22894 (N_22894,N_21707,N_20373);
nor U22895 (N_22895,N_20182,N_21601);
nor U22896 (N_22896,N_20015,N_20258);
xor U22897 (N_22897,N_20536,N_21669);
xor U22898 (N_22898,N_21157,N_20315);
xnor U22899 (N_22899,N_20036,N_21565);
or U22900 (N_22900,N_21261,N_20488);
nor U22901 (N_22901,N_21477,N_21641);
and U22902 (N_22902,N_20842,N_21083);
xnor U22903 (N_22903,N_20053,N_21520);
xnor U22904 (N_22904,N_21755,N_20975);
xnor U22905 (N_22905,N_21517,N_21993);
or U22906 (N_22906,N_20409,N_21278);
xnor U22907 (N_22907,N_20429,N_20509);
nor U22908 (N_22908,N_21437,N_20061);
xnor U22909 (N_22909,N_21484,N_20574);
nand U22910 (N_22910,N_21878,N_20997);
and U22911 (N_22911,N_20291,N_20072);
or U22912 (N_22912,N_20139,N_20845);
or U22913 (N_22913,N_20154,N_20251);
xnor U22914 (N_22914,N_21391,N_21628);
nand U22915 (N_22915,N_20893,N_20338);
and U22916 (N_22916,N_21364,N_21370);
and U22917 (N_22917,N_21347,N_20265);
xnor U22918 (N_22918,N_21195,N_20621);
or U22919 (N_22919,N_21574,N_20253);
xor U22920 (N_22920,N_20486,N_21895);
or U22921 (N_22921,N_20731,N_21953);
and U22922 (N_22922,N_21609,N_21760);
and U22923 (N_22923,N_21792,N_21994);
nor U22924 (N_22924,N_21496,N_20335);
or U22925 (N_22925,N_21716,N_21125);
nand U22926 (N_22926,N_21240,N_21836);
and U22927 (N_22927,N_20836,N_20901);
nand U22928 (N_22928,N_21670,N_20152);
nor U22929 (N_22929,N_21282,N_20580);
nor U22930 (N_22930,N_20757,N_21242);
or U22931 (N_22931,N_20814,N_21804);
or U22932 (N_22932,N_21636,N_20614);
xor U22933 (N_22933,N_21144,N_20544);
or U22934 (N_22934,N_20275,N_21615);
nand U22935 (N_22935,N_20393,N_20600);
or U22936 (N_22936,N_20426,N_21422);
nand U22937 (N_22937,N_20936,N_21241);
and U22938 (N_22938,N_20837,N_20356);
or U22939 (N_22939,N_21900,N_21948);
and U22940 (N_22940,N_20707,N_20588);
nand U22941 (N_22941,N_21541,N_21832);
and U22942 (N_22942,N_21226,N_20878);
nor U22943 (N_22943,N_21682,N_20098);
nor U22944 (N_22944,N_21936,N_21631);
and U22945 (N_22945,N_21925,N_21017);
nand U22946 (N_22946,N_21039,N_21009);
xor U22947 (N_22947,N_21531,N_20400);
nor U22948 (N_22948,N_20807,N_21662);
xor U22949 (N_22949,N_20629,N_20311);
or U22950 (N_22950,N_21817,N_21722);
nand U22951 (N_22951,N_20012,N_21302);
nand U22952 (N_22952,N_21376,N_20230);
and U22953 (N_22953,N_21715,N_21346);
nor U22954 (N_22954,N_21212,N_21405);
nand U22955 (N_22955,N_21450,N_21469);
nand U22956 (N_22956,N_21295,N_21704);
xor U22957 (N_22957,N_20823,N_20238);
xor U22958 (N_22958,N_21319,N_21648);
and U22959 (N_22959,N_21696,N_20048);
nand U22960 (N_22960,N_20375,N_20943);
and U22961 (N_22961,N_21220,N_21946);
or U22962 (N_22962,N_21050,N_21595);
or U22963 (N_22963,N_20049,N_21921);
nand U22964 (N_22964,N_21336,N_21340);
or U22965 (N_22965,N_21885,N_20738);
or U22966 (N_22966,N_20381,N_20203);
xnor U22967 (N_22967,N_20443,N_21889);
xor U22968 (N_22968,N_21690,N_20950);
and U22969 (N_22969,N_20401,N_21898);
and U22970 (N_22970,N_21515,N_21460);
nand U22971 (N_22971,N_20854,N_20788);
nand U22972 (N_22972,N_21251,N_20059);
or U22973 (N_22973,N_20608,N_21479);
and U22974 (N_22974,N_20522,N_21537);
or U22975 (N_22975,N_21151,N_20980);
nor U22976 (N_22976,N_20889,N_21522);
nand U22977 (N_22977,N_21822,N_21482);
or U22978 (N_22978,N_21963,N_20054);
and U22979 (N_22979,N_20029,N_21168);
nand U22980 (N_22980,N_20688,N_21003);
nor U22981 (N_22981,N_21571,N_20927);
nand U22982 (N_22982,N_20374,N_20032);
xor U22983 (N_22983,N_20946,N_20416);
or U22984 (N_22984,N_20179,N_20298);
xnor U22985 (N_22985,N_20016,N_20928);
xor U22986 (N_22986,N_21170,N_21343);
xnor U22987 (N_22987,N_20112,N_21153);
nand U22988 (N_22988,N_21432,N_20202);
and U22989 (N_22989,N_20394,N_21576);
or U22990 (N_22990,N_21929,N_20466);
nand U22991 (N_22991,N_21650,N_20442);
xnor U22992 (N_22992,N_20070,N_20086);
xor U22993 (N_22993,N_21052,N_21711);
and U22994 (N_22994,N_21414,N_20131);
nand U22995 (N_22995,N_21452,N_20756);
nor U22996 (N_22996,N_20655,N_21429);
nand U22997 (N_22997,N_21951,N_21228);
and U22998 (N_22998,N_20748,N_20404);
xnor U22999 (N_22999,N_20594,N_20411);
and U23000 (N_23000,N_21751,N_20735);
nand U23001 (N_23001,N_21035,N_21755);
and U23002 (N_23002,N_21529,N_20502);
and U23003 (N_23003,N_20445,N_21171);
nand U23004 (N_23004,N_20842,N_20459);
nor U23005 (N_23005,N_20702,N_21040);
xnor U23006 (N_23006,N_21230,N_20031);
or U23007 (N_23007,N_21973,N_20835);
or U23008 (N_23008,N_21305,N_20984);
or U23009 (N_23009,N_20932,N_21515);
or U23010 (N_23010,N_20709,N_21909);
or U23011 (N_23011,N_20415,N_21603);
and U23012 (N_23012,N_21035,N_20391);
xor U23013 (N_23013,N_21648,N_21753);
or U23014 (N_23014,N_20667,N_20195);
or U23015 (N_23015,N_21309,N_20981);
or U23016 (N_23016,N_21457,N_21638);
nor U23017 (N_23017,N_20826,N_20794);
xnor U23018 (N_23018,N_20515,N_21204);
and U23019 (N_23019,N_21566,N_21149);
nor U23020 (N_23020,N_20567,N_21306);
nor U23021 (N_23021,N_21100,N_20834);
nand U23022 (N_23022,N_20552,N_20661);
and U23023 (N_23023,N_20067,N_20856);
and U23024 (N_23024,N_21552,N_20650);
xnor U23025 (N_23025,N_21616,N_21439);
nand U23026 (N_23026,N_21127,N_21846);
or U23027 (N_23027,N_21210,N_21232);
or U23028 (N_23028,N_21737,N_20100);
xnor U23029 (N_23029,N_20021,N_20814);
or U23030 (N_23030,N_21955,N_21236);
or U23031 (N_23031,N_20239,N_20273);
xnor U23032 (N_23032,N_20207,N_20031);
nor U23033 (N_23033,N_21913,N_20783);
or U23034 (N_23034,N_21616,N_20266);
xor U23035 (N_23035,N_21291,N_20340);
nor U23036 (N_23036,N_21202,N_21302);
and U23037 (N_23037,N_20350,N_20689);
nand U23038 (N_23038,N_20886,N_21065);
and U23039 (N_23039,N_21220,N_20456);
and U23040 (N_23040,N_20835,N_21722);
xnor U23041 (N_23041,N_20909,N_21636);
nand U23042 (N_23042,N_20094,N_20137);
or U23043 (N_23043,N_21029,N_20589);
xor U23044 (N_23044,N_21755,N_20671);
nor U23045 (N_23045,N_21506,N_20390);
nand U23046 (N_23046,N_20011,N_21632);
xnor U23047 (N_23047,N_20372,N_21320);
and U23048 (N_23048,N_21282,N_21836);
and U23049 (N_23049,N_20070,N_21232);
xnor U23050 (N_23050,N_20077,N_21835);
or U23051 (N_23051,N_20580,N_20270);
nor U23052 (N_23052,N_21944,N_21904);
xor U23053 (N_23053,N_20080,N_21523);
or U23054 (N_23054,N_20442,N_20417);
or U23055 (N_23055,N_20379,N_20121);
or U23056 (N_23056,N_20886,N_20082);
xnor U23057 (N_23057,N_20269,N_20153);
nor U23058 (N_23058,N_20279,N_20207);
xnor U23059 (N_23059,N_20082,N_20302);
nor U23060 (N_23060,N_20385,N_20348);
nor U23061 (N_23061,N_20096,N_21935);
xor U23062 (N_23062,N_21795,N_21125);
xor U23063 (N_23063,N_21966,N_21587);
nand U23064 (N_23064,N_20167,N_21680);
nor U23065 (N_23065,N_21875,N_21719);
nor U23066 (N_23066,N_21925,N_21520);
and U23067 (N_23067,N_20133,N_21590);
and U23068 (N_23068,N_21816,N_20972);
and U23069 (N_23069,N_20178,N_20989);
xnor U23070 (N_23070,N_21491,N_21547);
nand U23071 (N_23071,N_20165,N_20602);
nor U23072 (N_23072,N_20908,N_20122);
and U23073 (N_23073,N_20763,N_20823);
nand U23074 (N_23074,N_20706,N_21022);
and U23075 (N_23075,N_20286,N_20942);
xnor U23076 (N_23076,N_21737,N_21169);
or U23077 (N_23077,N_21467,N_21740);
xor U23078 (N_23078,N_21308,N_21436);
nor U23079 (N_23079,N_21284,N_20187);
nor U23080 (N_23080,N_20586,N_21338);
nand U23081 (N_23081,N_21315,N_21625);
xnor U23082 (N_23082,N_20863,N_21728);
nand U23083 (N_23083,N_20224,N_20712);
and U23084 (N_23084,N_20608,N_20917);
or U23085 (N_23085,N_21362,N_20936);
and U23086 (N_23086,N_21811,N_21365);
or U23087 (N_23087,N_20108,N_20859);
or U23088 (N_23088,N_20734,N_20487);
nand U23089 (N_23089,N_20068,N_21256);
xor U23090 (N_23090,N_20261,N_20349);
xnor U23091 (N_23091,N_21446,N_21873);
xnor U23092 (N_23092,N_20046,N_20744);
nand U23093 (N_23093,N_21985,N_20820);
and U23094 (N_23094,N_20400,N_20409);
nor U23095 (N_23095,N_21200,N_20840);
nand U23096 (N_23096,N_21431,N_21014);
nor U23097 (N_23097,N_21472,N_20011);
xnor U23098 (N_23098,N_20316,N_21817);
xnor U23099 (N_23099,N_20487,N_21396);
or U23100 (N_23100,N_20669,N_20422);
xnor U23101 (N_23101,N_21575,N_20472);
nor U23102 (N_23102,N_21851,N_21121);
and U23103 (N_23103,N_20089,N_20910);
or U23104 (N_23104,N_20654,N_21458);
nor U23105 (N_23105,N_20897,N_21062);
and U23106 (N_23106,N_20042,N_20362);
or U23107 (N_23107,N_20542,N_21169);
and U23108 (N_23108,N_20301,N_20061);
nand U23109 (N_23109,N_21103,N_21807);
or U23110 (N_23110,N_20903,N_20715);
nand U23111 (N_23111,N_21801,N_21785);
nand U23112 (N_23112,N_20611,N_20730);
and U23113 (N_23113,N_21593,N_20802);
nor U23114 (N_23114,N_20490,N_20636);
nor U23115 (N_23115,N_21232,N_20477);
or U23116 (N_23116,N_21920,N_20564);
nor U23117 (N_23117,N_20699,N_20299);
or U23118 (N_23118,N_20882,N_20331);
and U23119 (N_23119,N_21886,N_21332);
nand U23120 (N_23120,N_21635,N_20703);
nand U23121 (N_23121,N_21236,N_21529);
nand U23122 (N_23122,N_20126,N_20742);
nand U23123 (N_23123,N_20660,N_21915);
nor U23124 (N_23124,N_21432,N_20317);
xor U23125 (N_23125,N_21955,N_20907);
and U23126 (N_23126,N_21688,N_21627);
nand U23127 (N_23127,N_21419,N_21052);
nand U23128 (N_23128,N_21827,N_21812);
or U23129 (N_23129,N_20352,N_20898);
nand U23130 (N_23130,N_21102,N_21363);
or U23131 (N_23131,N_20608,N_21135);
or U23132 (N_23132,N_21493,N_21692);
nor U23133 (N_23133,N_21715,N_21195);
or U23134 (N_23134,N_21955,N_20776);
nor U23135 (N_23135,N_21843,N_21360);
or U23136 (N_23136,N_20521,N_21078);
and U23137 (N_23137,N_21706,N_20644);
nand U23138 (N_23138,N_21216,N_20123);
nor U23139 (N_23139,N_21269,N_20929);
xor U23140 (N_23140,N_20640,N_20316);
nor U23141 (N_23141,N_20988,N_21178);
and U23142 (N_23142,N_20717,N_21575);
or U23143 (N_23143,N_21236,N_21972);
and U23144 (N_23144,N_21918,N_21711);
and U23145 (N_23145,N_21867,N_21429);
and U23146 (N_23146,N_21613,N_20800);
and U23147 (N_23147,N_21673,N_21715);
nand U23148 (N_23148,N_20593,N_20011);
xnor U23149 (N_23149,N_21093,N_21046);
nand U23150 (N_23150,N_20169,N_20330);
xor U23151 (N_23151,N_21110,N_21262);
xnor U23152 (N_23152,N_21378,N_20102);
and U23153 (N_23153,N_20416,N_21477);
xnor U23154 (N_23154,N_21569,N_20587);
nand U23155 (N_23155,N_21408,N_21510);
nor U23156 (N_23156,N_21929,N_20870);
nor U23157 (N_23157,N_21771,N_20300);
nand U23158 (N_23158,N_21057,N_20051);
nor U23159 (N_23159,N_21777,N_20115);
or U23160 (N_23160,N_20995,N_21858);
nor U23161 (N_23161,N_20425,N_20226);
xnor U23162 (N_23162,N_21507,N_20408);
nand U23163 (N_23163,N_21736,N_20374);
and U23164 (N_23164,N_20161,N_21820);
and U23165 (N_23165,N_21966,N_21215);
or U23166 (N_23166,N_20452,N_21602);
nor U23167 (N_23167,N_20479,N_20050);
nor U23168 (N_23168,N_21467,N_21654);
nor U23169 (N_23169,N_20344,N_20652);
xnor U23170 (N_23170,N_21850,N_20532);
nand U23171 (N_23171,N_20949,N_21060);
nor U23172 (N_23172,N_21530,N_21730);
nand U23173 (N_23173,N_21988,N_21636);
or U23174 (N_23174,N_20149,N_21172);
nand U23175 (N_23175,N_21758,N_21123);
xor U23176 (N_23176,N_20655,N_20638);
nand U23177 (N_23177,N_20837,N_21748);
nor U23178 (N_23178,N_21297,N_21854);
and U23179 (N_23179,N_20908,N_21346);
or U23180 (N_23180,N_21331,N_20436);
nand U23181 (N_23181,N_21325,N_20174);
and U23182 (N_23182,N_21571,N_20298);
and U23183 (N_23183,N_21591,N_20405);
nand U23184 (N_23184,N_20056,N_20668);
and U23185 (N_23185,N_21705,N_21486);
nand U23186 (N_23186,N_20596,N_20469);
and U23187 (N_23187,N_21117,N_21913);
xor U23188 (N_23188,N_21930,N_20308);
or U23189 (N_23189,N_21723,N_21887);
nand U23190 (N_23190,N_21089,N_20226);
or U23191 (N_23191,N_21572,N_21631);
or U23192 (N_23192,N_20746,N_20664);
xnor U23193 (N_23193,N_21495,N_20965);
xnor U23194 (N_23194,N_20175,N_20124);
or U23195 (N_23195,N_21293,N_20533);
and U23196 (N_23196,N_20693,N_20664);
xnor U23197 (N_23197,N_20657,N_20745);
xor U23198 (N_23198,N_21486,N_21907);
or U23199 (N_23199,N_21224,N_21870);
and U23200 (N_23200,N_21321,N_20587);
xor U23201 (N_23201,N_20351,N_20558);
xnor U23202 (N_23202,N_20194,N_20274);
and U23203 (N_23203,N_20362,N_21768);
nor U23204 (N_23204,N_20490,N_20051);
nand U23205 (N_23205,N_20163,N_21808);
or U23206 (N_23206,N_20375,N_21716);
or U23207 (N_23207,N_21073,N_20125);
or U23208 (N_23208,N_21109,N_20343);
xor U23209 (N_23209,N_20427,N_21177);
nand U23210 (N_23210,N_21158,N_21078);
or U23211 (N_23211,N_20873,N_20981);
or U23212 (N_23212,N_21583,N_21345);
xnor U23213 (N_23213,N_21654,N_21587);
xnor U23214 (N_23214,N_21912,N_20334);
nor U23215 (N_23215,N_20373,N_21220);
nand U23216 (N_23216,N_21440,N_20400);
xor U23217 (N_23217,N_21929,N_21175);
nor U23218 (N_23218,N_21818,N_21946);
or U23219 (N_23219,N_21208,N_21472);
nor U23220 (N_23220,N_21954,N_21986);
nor U23221 (N_23221,N_20599,N_20342);
nand U23222 (N_23222,N_20427,N_21529);
xnor U23223 (N_23223,N_21007,N_21463);
or U23224 (N_23224,N_20613,N_20164);
xnor U23225 (N_23225,N_21793,N_21085);
nand U23226 (N_23226,N_21028,N_21769);
nand U23227 (N_23227,N_20806,N_21993);
nor U23228 (N_23228,N_20772,N_21601);
and U23229 (N_23229,N_21238,N_21655);
xor U23230 (N_23230,N_20525,N_21569);
xor U23231 (N_23231,N_20353,N_20559);
nor U23232 (N_23232,N_20031,N_21995);
xor U23233 (N_23233,N_21126,N_20430);
or U23234 (N_23234,N_21174,N_21712);
nand U23235 (N_23235,N_20387,N_20749);
xnor U23236 (N_23236,N_20887,N_21447);
or U23237 (N_23237,N_20539,N_21705);
nand U23238 (N_23238,N_21422,N_20127);
xor U23239 (N_23239,N_21809,N_20124);
and U23240 (N_23240,N_21114,N_21651);
nor U23241 (N_23241,N_20333,N_20101);
and U23242 (N_23242,N_20381,N_21735);
xor U23243 (N_23243,N_21653,N_21556);
and U23244 (N_23244,N_20516,N_21056);
nand U23245 (N_23245,N_20321,N_21667);
nor U23246 (N_23246,N_21596,N_21172);
and U23247 (N_23247,N_21910,N_21658);
and U23248 (N_23248,N_20557,N_21094);
nand U23249 (N_23249,N_21810,N_21622);
or U23250 (N_23250,N_21656,N_20430);
xor U23251 (N_23251,N_21472,N_21343);
nand U23252 (N_23252,N_20330,N_20530);
xor U23253 (N_23253,N_20799,N_21916);
and U23254 (N_23254,N_20989,N_20527);
nor U23255 (N_23255,N_20653,N_21967);
xnor U23256 (N_23256,N_20946,N_20126);
and U23257 (N_23257,N_21803,N_20707);
and U23258 (N_23258,N_20215,N_21756);
nand U23259 (N_23259,N_21354,N_21642);
or U23260 (N_23260,N_20739,N_20697);
or U23261 (N_23261,N_21077,N_20877);
or U23262 (N_23262,N_21549,N_21427);
nand U23263 (N_23263,N_20745,N_21694);
nor U23264 (N_23264,N_20069,N_21715);
or U23265 (N_23265,N_21720,N_20216);
xnor U23266 (N_23266,N_20249,N_21816);
xor U23267 (N_23267,N_21608,N_20314);
or U23268 (N_23268,N_21717,N_20386);
and U23269 (N_23269,N_21949,N_20100);
or U23270 (N_23270,N_20941,N_20455);
nor U23271 (N_23271,N_20080,N_20735);
nor U23272 (N_23272,N_21216,N_21865);
xnor U23273 (N_23273,N_21617,N_21913);
and U23274 (N_23274,N_21854,N_21294);
nand U23275 (N_23275,N_21297,N_20419);
nand U23276 (N_23276,N_20126,N_20148);
or U23277 (N_23277,N_20804,N_21900);
nor U23278 (N_23278,N_20133,N_21062);
nor U23279 (N_23279,N_20634,N_20147);
or U23280 (N_23280,N_20545,N_20521);
nor U23281 (N_23281,N_21016,N_20702);
and U23282 (N_23282,N_20937,N_21231);
xor U23283 (N_23283,N_21822,N_20469);
xnor U23284 (N_23284,N_20464,N_20714);
and U23285 (N_23285,N_20409,N_20827);
or U23286 (N_23286,N_21370,N_21076);
nor U23287 (N_23287,N_21327,N_20023);
nand U23288 (N_23288,N_21804,N_21281);
nor U23289 (N_23289,N_20803,N_21701);
xnor U23290 (N_23290,N_20503,N_20508);
nor U23291 (N_23291,N_20374,N_21212);
nor U23292 (N_23292,N_21222,N_21506);
nor U23293 (N_23293,N_20951,N_20237);
xor U23294 (N_23294,N_21251,N_20155);
xor U23295 (N_23295,N_20155,N_20663);
nand U23296 (N_23296,N_21579,N_21053);
xnor U23297 (N_23297,N_20088,N_20198);
nor U23298 (N_23298,N_20510,N_20577);
and U23299 (N_23299,N_21852,N_21554);
nand U23300 (N_23300,N_21731,N_21725);
nand U23301 (N_23301,N_20752,N_20346);
or U23302 (N_23302,N_21538,N_20543);
nand U23303 (N_23303,N_21681,N_21103);
nand U23304 (N_23304,N_21937,N_21481);
nor U23305 (N_23305,N_21473,N_20907);
nor U23306 (N_23306,N_20961,N_21078);
and U23307 (N_23307,N_21426,N_21372);
xnor U23308 (N_23308,N_21241,N_21762);
nor U23309 (N_23309,N_21245,N_20839);
and U23310 (N_23310,N_21727,N_20978);
nand U23311 (N_23311,N_21488,N_20558);
or U23312 (N_23312,N_21043,N_21866);
xor U23313 (N_23313,N_20015,N_21229);
nor U23314 (N_23314,N_21440,N_20916);
or U23315 (N_23315,N_20739,N_21853);
xnor U23316 (N_23316,N_20383,N_20939);
nand U23317 (N_23317,N_20739,N_20142);
and U23318 (N_23318,N_20604,N_20850);
and U23319 (N_23319,N_20668,N_21520);
xnor U23320 (N_23320,N_21428,N_21443);
xor U23321 (N_23321,N_21117,N_21551);
or U23322 (N_23322,N_21778,N_20882);
nor U23323 (N_23323,N_20017,N_21391);
nand U23324 (N_23324,N_21434,N_21135);
nor U23325 (N_23325,N_20199,N_20954);
nor U23326 (N_23326,N_21844,N_21091);
nand U23327 (N_23327,N_20044,N_21318);
and U23328 (N_23328,N_20097,N_21403);
nand U23329 (N_23329,N_20058,N_20483);
nor U23330 (N_23330,N_20642,N_20461);
xnor U23331 (N_23331,N_20852,N_21265);
nor U23332 (N_23332,N_20495,N_21483);
and U23333 (N_23333,N_20887,N_21419);
and U23334 (N_23334,N_20978,N_20132);
nand U23335 (N_23335,N_21914,N_20370);
and U23336 (N_23336,N_21668,N_20518);
nand U23337 (N_23337,N_21000,N_21978);
or U23338 (N_23338,N_21123,N_20569);
xnor U23339 (N_23339,N_20117,N_20743);
or U23340 (N_23340,N_20186,N_21429);
nand U23341 (N_23341,N_20017,N_21927);
or U23342 (N_23342,N_20105,N_20148);
or U23343 (N_23343,N_21627,N_20757);
or U23344 (N_23344,N_21717,N_21516);
and U23345 (N_23345,N_20703,N_21948);
or U23346 (N_23346,N_20631,N_21693);
nand U23347 (N_23347,N_20761,N_20897);
nor U23348 (N_23348,N_20205,N_20802);
and U23349 (N_23349,N_21841,N_21325);
xor U23350 (N_23350,N_21304,N_21349);
xnor U23351 (N_23351,N_21298,N_20739);
nand U23352 (N_23352,N_21253,N_20333);
nand U23353 (N_23353,N_20131,N_20874);
and U23354 (N_23354,N_21732,N_20180);
or U23355 (N_23355,N_21181,N_20973);
or U23356 (N_23356,N_21099,N_20189);
xor U23357 (N_23357,N_21591,N_21730);
or U23358 (N_23358,N_20722,N_20359);
nand U23359 (N_23359,N_20932,N_20310);
nor U23360 (N_23360,N_21342,N_21588);
nor U23361 (N_23361,N_21920,N_21918);
and U23362 (N_23362,N_20932,N_20846);
or U23363 (N_23363,N_21038,N_20134);
nor U23364 (N_23364,N_21240,N_20602);
and U23365 (N_23365,N_21738,N_21677);
or U23366 (N_23366,N_21814,N_20449);
or U23367 (N_23367,N_20273,N_21713);
nor U23368 (N_23368,N_21449,N_20386);
xor U23369 (N_23369,N_20782,N_20978);
and U23370 (N_23370,N_21746,N_21997);
nor U23371 (N_23371,N_21323,N_21944);
nor U23372 (N_23372,N_20940,N_21989);
or U23373 (N_23373,N_20466,N_21187);
xor U23374 (N_23374,N_20816,N_20327);
xor U23375 (N_23375,N_21926,N_20779);
nand U23376 (N_23376,N_21336,N_20601);
or U23377 (N_23377,N_21842,N_20080);
nand U23378 (N_23378,N_21210,N_20664);
and U23379 (N_23379,N_20031,N_20159);
and U23380 (N_23380,N_21592,N_21971);
xnor U23381 (N_23381,N_20350,N_21067);
nand U23382 (N_23382,N_20909,N_20898);
or U23383 (N_23383,N_20296,N_20227);
nand U23384 (N_23384,N_20638,N_21797);
nand U23385 (N_23385,N_21947,N_21465);
or U23386 (N_23386,N_20235,N_20345);
xnor U23387 (N_23387,N_20657,N_21034);
nor U23388 (N_23388,N_21285,N_21578);
xnor U23389 (N_23389,N_20689,N_21716);
nand U23390 (N_23390,N_20930,N_21251);
xnor U23391 (N_23391,N_21435,N_21002);
nor U23392 (N_23392,N_20352,N_20858);
xnor U23393 (N_23393,N_21784,N_20430);
or U23394 (N_23394,N_21200,N_21371);
or U23395 (N_23395,N_21603,N_21814);
or U23396 (N_23396,N_20307,N_20633);
or U23397 (N_23397,N_20908,N_21498);
or U23398 (N_23398,N_21249,N_21094);
xnor U23399 (N_23399,N_21334,N_20531);
nand U23400 (N_23400,N_21727,N_21311);
and U23401 (N_23401,N_21015,N_21660);
nor U23402 (N_23402,N_20242,N_21092);
nor U23403 (N_23403,N_20136,N_20891);
nor U23404 (N_23404,N_20205,N_20836);
xnor U23405 (N_23405,N_20031,N_21481);
and U23406 (N_23406,N_21175,N_20518);
nand U23407 (N_23407,N_20718,N_21867);
or U23408 (N_23408,N_21830,N_21355);
xor U23409 (N_23409,N_20286,N_20614);
xnor U23410 (N_23410,N_21505,N_20140);
nor U23411 (N_23411,N_21018,N_20583);
and U23412 (N_23412,N_20366,N_20131);
or U23413 (N_23413,N_21484,N_20490);
nor U23414 (N_23414,N_21809,N_20451);
and U23415 (N_23415,N_20645,N_20303);
nor U23416 (N_23416,N_21373,N_21194);
and U23417 (N_23417,N_20155,N_21312);
or U23418 (N_23418,N_20098,N_21476);
or U23419 (N_23419,N_21458,N_20021);
xor U23420 (N_23420,N_21784,N_20629);
xnor U23421 (N_23421,N_20543,N_21373);
xor U23422 (N_23422,N_20447,N_21299);
or U23423 (N_23423,N_21779,N_21471);
nand U23424 (N_23424,N_21708,N_21344);
xnor U23425 (N_23425,N_20132,N_20085);
xnor U23426 (N_23426,N_20342,N_21499);
xor U23427 (N_23427,N_20566,N_20757);
nand U23428 (N_23428,N_21746,N_21196);
nand U23429 (N_23429,N_20312,N_21877);
xor U23430 (N_23430,N_20065,N_21689);
nor U23431 (N_23431,N_21898,N_21607);
and U23432 (N_23432,N_21104,N_21012);
or U23433 (N_23433,N_21475,N_20034);
xor U23434 (N_23434,N_20139,N_21708);
and U23435 (N_23435,N_20908,N_20526);
nand U23436 (N_23436,N_20215,N_21524);
nand U23437 (N_23437,N_21323,N_21678);
and U23438 (N_23438,N_20287,N_20991);
nor U23439 (N_23439,N_21690,N_20257);
xnor U23440 (N_23440,N_21741,N_20216);
nor U23441 (N_23441,N_21139,N_21681);
nor U23442 (N_23442,N_21416,N_20933);
nand U23443 (N_23443,N_20697,N_20257);
nand U23444 (N_23444,N_20008,N_20305);
xnor U23445 (N_23445,N_21131,N_20060);
nand U23446 (N_23446,N_20574,N_21538);
nand U23447 (N_23447,N_21873,N_20595);
and U23448 (N_23448,N_20314,N_21932);
or U23449 (N_23449,N_21072,N_21022);
and U23450 (N_23450,N_21466,N_20208);
nor U23451 (N_23451,N_20423,N_20260);
xor U23452 (N_23452,N_20992,N_21056);
nand U23453 (N_23453,N_21560,N_20212);
and U23454 (N_23454,N_20938,N_20421);
nand U23455 (N_23455,N_20318,N_20584);
and U23456 (N_23456,N_21510,N_21405);
or U23457 (N_23457,N_21194,N_21875);
and U23458 (N_23458,N_20242,N_20402);
nand U23459 (N_23459,N_21396,N_20421);
and U23460 (N_23460,N_21207,N_21376);
nor U23461 (N_23461,N_21811,N_21107);
and U23462 (N_23462,N_20258,N_21553);
or U23463 (N_23463,N_20811,N_20989);
and U23464 (N_23464,N_21905,N_21339);
and U23465 (N_23465,N_20731,N_21667);
or U23466 (N_23466,N_21106,N_21725);
or U23467 (N_23467,N_21645,N_20289);
nor U23468 (N_23468,N_21159,N_21238);
and U23469 (N_23469,N_21099,N_21719);
xnor U23470 (N_23470,N_21843,N_21500);
nand U23471 (N_23471,N_20299,N_21931);
and U23472 (N_23472,N_20984,N_20618);
xor U23473 (N_23473,N_20879,N_20030);
xor U23474 (N_23474,N_20063,N_20560);
or U23475 (N_23475,N_20603,N_20012);
or U23476 (N_23476,N_20731,N_21895);
nand U23477 (N_23477,N_20540,N_21932);
xnor U23478 (N_23478,N_21069,N_20476);
xnor U23479 (N_23479,N_20557,N_21795);
and U23480 (N_23480,N_20031,N_20455);
and U23481 (N_23481,N_20305,N_21496);
nand U23482 (N_23482,N_21151,N_20825);
nand U23483 (N_23483,N_20197,N_20263);
and U23484 (N_23484,N_20249,N_21021);
xor U23485 (N_23485,N_20689,N_20375);
nand U23486 (N_23486,N_20670,N_20291);
and U23487 (N_23487,N_21520,N_21154);
xnor U23488 (N_23488,N_20568,N_21641);
nor U23489 (N_23489,N_20436,N_21563);
or U23490 (N_23490,N_21317,N_20778);
xnor U23491 (N_23491,N_20460,N_20505);
xor U23492 (N_23492,N_21504,N_20388);
nand U23493 (N_23493,N_20131,N_20099);
nor U23494 (N_23494,N_21388,N_20934);
nand U23495 (N_23495,N_20161,N_21744);
nand U23496 (N_23496,N_21561,N_21683);
and U23497 (N_23497,N_21998,N_21061);
or U23498 (N_23498,N_21363,N_20582);
or U23499 (N_23499,N_21376,N_21195);
nor U23500 (N_23500,N_20755,N_20631);
nor U23501 (N_23501,N_20026,N_20827);
nand U23502 (N_23502,N_20913,N_20553);
nand U23503 (N_23503,N_21034,N_20199);
nand U23504 (N_23504,N_20570,N_20023);
nand U23505 (N_23505,N_21835,N_20950);
or U23506 (N_23506,N_21306,N_21073);
nand U23507 (N_23507,N_21462,N_21070);
nor U23508 (N_23508,N_21225,N_20318);
or U23509 (N_23509,N_21170,N_21488);
nand U23510 (N_23510,N_20496,N_21877);
nand U23511 (N_23511,N_21007,N_20941);
and U23512 (N_23512,N_20297,N_20655);
nor U23513 (N_23513,N_20578,N_21119);
xor U23514 (N_23514,N_21277,N_20926);
nand U23515 (N_23515,N_21260,N_20051);
and U23516 (N_23516,N_21930,N_20083);
or U23517 (N_23517,N_20739,N_20565);
nand U23518 (N_23518,N_21784,N_20613);
nand U23519 (N_23519,N_20791,N_20997);
xor U23520 (N_23520,N_20938,N_20944);
xnor U23521 (N_23521,N_20933,N_21128);
or U23522 (N_23522,N_21537,N_21910);
nor U23523 (N_23523,N_21793,N_20701);
xor U23524 (N_23524,N_20847,N_20674);
or U23525 (N_23525,N_21935,N_20859);
or U23526 (N_23526,N_20843,N_20925);
and U23527 (N_23527,N_21446,N_20940);
and U23528 (N_23528,N_21648,N_20733);
or U23529 (N_23529,N_20499,N_21406);
and U23530 (N_23530,N_20429,N_21322);
xnor U23531 (N_23531,N_20138,N_21137);
and U23532 (N_23532,N_21099,N_21385);
nand U23533 (N_23533,N_20388,N_21436);
nand U23534 (N_23534,N_20437,N_21807);
nand U23535 (N_23535,N_21829,N_21197);
and U23536 (N_23536,N_20207,N_20974);
or U23537 (N_23537,N_20394,N_20276);
or U23538 (N_23538,N_21870,N_21094);
nor U23539 (N_23539,N_21862,N_20346);
nor U23540 (N_23540,N_20135,N_21460);
and U23541 (N_23541,N_20920,N_21222);
and U23542 (N_23542,N_20195,N_21800);
nor U23543 (N_23543,N_20137,N_20282);
and U23544 (N_23544,N_21388,N_21807);
nor U23545 (N_23545,N_20927,N_20503);
xnor U23546 (N_23546,N_20031,N_20717);
or U23547 (N_23547,N_21273,N_21013);
or U23548 (N_23548,N_20683,N_21116);
and U23549 (N_23549,N_20763,N_21083);
or U23550 (N_23550,N_21604,N_20276);
and U23551 (N_23551,N_21581,N_21815);
or U23552 (N_23552,N_20768,N_21835);
and U23553 (N_23553,N_20731,N_21775);
or U23554 (N_23554,N_20321,N_21035);
nor U23555 (N_23555,N_21429,N_21576);
or U23556 (N_23556,N_21578,N_20858);
xnor U23557 (N_23557,N_20350,N_21571);
or U23558 (N_23558,N_20247,N_21092);
or U23559 (N_23559,N_21333,N_21783);
and U23560 (N_23560,N_21692,N_20629);
and U23561 (N_23561,N_20713,N_20859);
xnor U23562 (N_23562,N_21710,N_21207);
nand U23563 (N_23563,N_21169,N_21789);
nor U23564 (N_23564,N_21273,N_21460);
and U23565 (N_23565,N_20080,N_20700);
and U23566 (N_23566,N_21128,N_20905);
nor U23567 (N_23567,N_20374,N_21847);
and U23568 (N_23568,N_20886,N_20691);
and U23569 (N_23569,N_21787,N_21934);
nand U23570 (N_23570,N_20487,N_21828);
or U23571 (N_23571,N_21201,N_21915);
xor U23572 (N_23572,N_20502,N_20535);
and U23573 (N_23573,N_21742,N_20422);
xor U23574 (N_23574,N_20339,N_21495);
and U23575 (N_23575,N_20074,N_21406);
and U23576 (N_23576,N_20180,N_20190);
and U23577 (N_23577,N_20436,N_20866);
xor U23578 (N_23578,N_20199,N_20573);
and U23579 (N_23579,N_20613,N_21164);
nand U23580 (N_23580,N_20204,N_20655);
and U23581 (N_23581,N_21586,N_20468);
nand U23582 (N_23582,N_21317,N_21712);
xnor U23583 (N_23583,N_21322,N_21910);
nand U23584 (N_23584,N_20292,N_21149);
and U23585 (N_23585,N_20288,N_20172);
or U23586 (N_23586,N_20612,N_20883);
or U23587 (N_23587,N_21807,N_20774);
xor U23588 (N_23588,N_20856,N_20385);
and U23589 (N_23589,N_20063,N_21496);
or U23590 (N_23590,N_20937,N_20393);
or U23591 (N_23591,N_21653,N_20655);
nand U23592 (N_23592,N_20050,N_20780);
or U23593 (N_23593,N_21943,N_20166);
and U23594 (N_23594,N_21162,N_20784);
xor U23595 (N_23595,N_20287,N_21972);
or U23596 (N_23596,N_21024,N_20661);
and U23597 (N_23597,N_20077,N_21948);
nor U23598 (N_23598,N_20312,N_21761);
xnor U23599 (N_23599,N_21883,N_21482);
xnor U23600 (N_23600,N_21437,N_20811);
xor U23601 (N_23601,N_20152,N_20698);
xor U23602 (N_23602,N_20834,N_21033);
and U23603 (N_23603,N_21863,N_20813);
xor U23604 (N_23604,N_20293,N_20142);
or U23605 (N_23605,N_20618,N_20775);
nor U23606 (N_23606,N_20861,N_21458);
and U23607 (N_23607,N_21255,N_20403);
nor U23608 (N_23608,N_21892,N_20392);
nand U23609 (N_23609,N_20266,N_21866);
and U23610 (N_23610,N_20386,N_21702);
nor U23611 (N_23611,N_20324,N_21119);
xnor U23612 (N_23612,N_21274,N_20783);
and U23613 (N_23613,N_20811,N_21738);
xor U23614 (N_23614,N_20521,N_21145);
and U23615 (N_23615,N_21127,N_20097);
or U23616 (N_23616,N_20311,N_21621);
nor U23617 (N_23617,N_21496,N_21101);
nand U23618 (N_23618,N_21162,N_21831);
nor U23619 (N_23619,N_21790,N_21212);
nor U23620 (N_23620,N_21042,N_21762);
nor U23621 (N_23621,N_21792,N_21111);
xnor U23622 (N_23622,N_21894,N_21434);
and U23623 (N_23623,N_21208,N_20246);
and U23624 (N_23624,N_21078,N_20681);
and U23625 (N_23625,N_20934,N_20131);
nor U23626 (N_23626,N_21748,N_20849);
nor U23627 (N_23627,N_21787,N_20532);
and U23628 (N_23628,N_20079,N_21269);
or U23629 (N_23629,N_20308,N_20771);
and U23630 (N_23630,N_20487,N_20793);
or U23631 (N_23631,N_20279,N_21341);
and U23632 (N_23632,N_21345,N_20408);
or U23633 (N_23633,N_21247,N_21802);
xor U23634 (N_23634,N_20017,N_21456);
and U23635 (N_23635,N_21356,N_21384);
xor U23636 (N_23636,N_21536,N_20586);
xor U23637 (N_23637,N_20911,N_21094);
xor U23638 (N_23638,N_21340,N_21830);
nand U23639 (N_23639,N_21928,N_20198);
and U23640 (N_23640,N_21031,N_20392);
nand U23641 (N_23641,N_20167,N_20408);
nand U23642 (N_23642,N_20985,N_21694);
and U23643 (N_23643,N_20834,N_21691);
or U23644 (N_23644,N_21305,N_20152);
nor U23645 (N_23645,N_21345,N_20587);
nor U23646 (N_23646,N_20717,N_21438);
xor U23647 (N_23647,N_20072,N_21907);
or U23648 (N_23648,N_20821,N_20028);
nor U23649 (N_23649,N_20214,N_21928);
xor U23650 (N_23650,N_21888,N_21638);
or U23651 (N_23651,N_20532,N_20492);
nand U23652 (N_23652,N_21471,N_21437);
and U23653 (N_23653,N_20897,N_21294);
and U23654 (N_23654,N_20037,N_21809);
nand U23655 (N_23655,N_21185,N_20067);
and U23656 (N_23656,N_21031,N_20319);
and U23657 (N_23657,N_21386,N_21563);
nand U23658 (N_23658,N_21749,N_20019);
nor U23659 (N_23659,N_21036,N_20963);
xnor U23660 (N_23660,N_20142,N_21994);
xnor U23661 (N_23661,N_20015,N_20162);
xnor U23662 (N_23662,N_20231,N_20119);
xor U23663 (N_23663,N_21607,N_20941);
xor U23664 (N_23664,N_21809,N_21031);
or U23665 (N_23665,N_20405,N_21167);
nand U23666 (N_23666,N_21556,N_20933);
nor U23667 (N_23667,N_21049,N_21327);
xor U23668 (N_23668,N_21728,N_21644);
nand U23669 (N_23669,N_20296,N_21596);
or U23670 (N_23670,N_20329,N_21139);
nor U23671 (N_23671,N_20042,N_20363);
xor U23672 (N_23672,N_21047,N_20531);
or U23673 (N_23673,N_21847,N_21555);
nor U23674 (N_23674,N_20432,N_20008);
nor U23675 (N_23675,N_20299,N_21330);
nor U23676 (N_23676,N_20882,N_21200);
nand U23677 (N_23677,N_21107,N_21720);
xnor U23678 (N_23678,N_21980,N_21550);
nand U23679 (N_23679,N_20355,N_20205);
and U23680 (N_23680,N_20396,N_20091);
nand U23681 (N_23681,N_21320,N_21995);
or U23682 (N_23682,N_20837,N_21499);
and U23683 (N_23683,N_20000,N_20265);
or U23684 (N_23684,N_20741,N_21186);
nor U23685 (N_23685,N_20886,N_20369);
or U23686 (N_23686,N_21411,N_21607);
and U23687 (N_23687,N_21632,N_20446);
nand U23688 (N_23688,N_21194,N_20078);
and U23689 (N_23689,N_20292,N_21050);
xor U23690 (N_23690,N_20381,N_21513);
xnor U23691 (N_23691,N_21837,N_21002);
or U23692 (N_23692,N_20903,N_21571);
nand U23693 (N_23693,N_21866,N_20906);
nor U23694 (N_23694,N_20542,N_20647);
nand U23695 (N_23695,N_20644,N_21631);
or U23696 (N_23696,N_20683,N_20109);
and U23697 (N_23697,N_21932,N_20794);
nor U23698 (N_23698,N_20284,N_20957);
xor U23699 (N_23699,N_20433,N_20824);
xnor U23700 (N_23700,N_20171,N_21365);
or U23701 (N_23701,N_20359,N_20814);
or U23702 (N_23702,N_21947,N_21076);
nor U23703 (N_23703,N_21513,N_21450);
nand U23704 (N_23704,N_20493,N_20324);
and U23705 (N_23705,N_20220,N_20969);
nand U23706 (N_23706,N_20425,N_20157);
xnor U23707 (N_23707,N_20695,N_21643);
nand U23708 (N_23708,N_21068,N_21871);
nand U23709 (N_23709,N_21448,N_20181);
nand U23710 (N_23710,N_21960,N_20691);
nor U23711 (N_23711,N_21009,N_20087);
nand U23712 (N_23712,N_20023,N_20344);
nor U23713 (N_23713,N_20273,N_20873);
xor U23714 (N_23714,N_20833,N_21569);
nand U23715 (N_23715,N_21457,N_20155);
xnor U23716 (N_23716,N_21443,N_21228);
nor U23717 (N_23717,N_20198,N_21759);
or U23718 (N_23718,N_21816,N_20648);
nor U23719 (N_23719,N_21055,N_21820);
nand U23720 (N_23720,N_21035,N_21778);
xnor U23721 (N_23721,N_21971,N_20052);
nor U23722 (N_23722,N_21465,N_21411);
and U23723 (N_23723,N_20701,N_20587);
nand U23724 (N_23724,N_20778,N_21220);
nor U23725 (N_23725,N_21113,N_20671);
nand U23726 (N_23726,N_20897,N_20752);
and U23727 (N_23727,N_20648,N_20749);
xor U23728 (N_23728,N_20643,N_20758);
xnor U23729 (N_23729,N_21071,N_20895);
or U23730 (N_23730,N_20136,N_20052);
nor U23731 (N_23731,N_20917,N_21447);
nor U23732 (N_23732,N_21063,N_20939);
and U23733 (N_23733,N_20485,N_20223);
nor U23734 (N_23734,N_21867,N_21789);
and U23735 (N_23735,N_20441,N_21797);
xor U23736 (N_23736,N_21739,N_21785);
nor U23737 (N_23737,N_21678,N_20993);
nand U23738 (N_23738,N_21362,N_21073);
nand U23739 (N_23739,N_20333,N_20613);
or U23740 (N_23740,N_20788,N_21494);
and U23741 (N_23741,N_20321,N_21207);
and U23742 (N_23742,N_21050,N_21203);
nor U23743 (N_23743,N_21814,N_20953);
xnor U23744 (N_23744,N_20626,N_20898);
and U23745 (N_23745,N_20832,N_20316);
nor U23746 (N_23746,N_20967,N_20433);
nor U23747 (N_23747,N_21518,N_21938);
and U23748 (N_23748,N_20384,N_20241);
or U23749 (N_23749,N_21045,N_20738);
or U23750 (N_23750,N_20862,N_20584);
nand U23751 (N_23751,N_20338,N_20638);
xor U23752 (N_23752,N_20980,N_21428);
nor U23753 (N_23753,N_20614,N_21828);
and U23754 (N_23754,N_21872,N_20169);
nor U23755 (N_23755,N_21497,N_21578);
and U23756 (N_23756,N_21599,N_20516);
nor U23757 (N_23757,N_20177,N_20224);
xnor U23758 (N_23758,N_20941,N_21281);
xnor U23759 (N_23759,N_20922,N_21124);
or U23760 (N_23760,N_20000,N_21237);
nor U23761 (N_23761,N_20044,N_20266);
and U23762 (N_23762,N_20829,N_20076);
nand U23763 (N_23763,N_20762,N_21493);
and U23764 (N_23764,N_20891,N_20041);
and U23765 (N_23765,N_21801,N_21560);
nor U23766 (N_23766,N_20308,N_21252);
nand U23767 (N_23767,N_20036,N_21745);
and U23768 (N_23768,N_21470,N_21862);
nand U23769 (N_23769,N_21364,N_21094);
and U23770 (N_23770,N_21302,N_21318);
nor U23771 (N_23771,N_20952,N_21442);
xnor U23772 (N_23772,N_20112,N_20104);
nand U23773 (N_23773,N_20336,N_21394);
or U23774 (N_23774,N_20817,N_21730);
nand U23775 (N_23775,N_20171,N_21195);
xor U23776 (N_23776,N_21691,N_21575);
and U23777 (N_23777,N_20804,N_20364);
xor U23778 (N_23778,N_20065,N_20488);
nor U23779 (N_23779,N_20622,N_20235);
nand U23780 (N_23780,N_20763,N_20831);
nand U23781 (N_23781,N_21374,N_20048);
or U23782 (N_23782,N_20122,N_20930);
nand U23783 (N_23783,N_21031,N_20524);
nand U23784 (N_23784,N_20454,N_20260);
nor U23785 (N_23785,N_20469,N_20653);
nor U23786 (N_23786,N_21243,N_20230);
xnor U23787 (N_23787,N_21207,N_20946);
xor U23788 (N_23788,N_20558,N_21290);
and U23789 (N_23789,N_20307,N_21904);
and U23790 (N_23790,N_21628,N_20127);
or U23791 (N_23791,N_21235,N_21370);
and U23792 (N_23792,N_21291,N_21026);
or U23793 (N_23793,N_21495,N_20551);
and U23794 (N_23794,N_20841,N_21845);
nand U23795 (N_23795,N_21466,N_21115);
or U23796 (N_23796,N_21628,N_21313);
nor U23797 (N_23797,N_20241,N_21988);
nor U23798 (N_23798,N_21841,N_21692);
nor U23799 (N_23799,N_20626,N_20372);
nand U23800 (N_23800,N_20742,N_20237);
nor U23801 (N_23801,N_20015,N_20942);
xnor U23802 (N_23802,N_20151,N_20982);
or U23803 (N_23803,N_21233,N_21851);
and U23804 (N_23804,N_21573,N_20623);
xor U23805 (N_23805,N_20175,N_21856);
and U23806 (N_23806,N_21609,N_20691);
or U23807 (N_23807,N_21149,N_21132);
and U23808 (N_23808,N_21278,N_21089);
nor U23809 (N_23809,N_21683,N_20599);
and U23810 (N_23810,N_20152,N_20695);
and U23811 (N_23811,N_21031,N_21542);
xor U23812 (N_23812,N_21374,N_20748);
and U23813 (N_23813,N_21873,N_20168);
and U23814 (N_23814,N_21330,N_20347);
nor U23815 (N_23815,N_20598,N_21127);
nor U23816 (N_23816,N_20230,N_20837);
or U23817 (N_23817,N_20931,N_21639);
xor U23818 (N_23818,N_20029,N_21762);
xor U23819 (N_23819,N_20502,N_20949);
nor U23820 (N_23820,N_21253,N_21738);
nand U23821 (N_23821,N_20103,N_21460);
nor U23822 (N_23822,N_21247,N_20208);
or U23823 (N_23823,N_21048,N_20846);
and U23824 (N_23824,N_20023,N_20408);
nor U23825 (N_23825,N_21992,N_20737);
and U23826 (N_23826,N_21328,N_20831);
xor U23827 (N_23827,N_20101,N_20122);
nor U23828 (N_23828,N_21381,N_21548);
nor U23829 (N_23829,N_21114,N_21396);
nor U23830 (N_23830,N_21736,N_21904);
and U23831 (N_23831,N_21421,N_20640);
or U23832 (N_23832,N_20323,N_20909);
nor U23833 (N_23833,N_21645,N_21178);
nor U23834 (N_23834,N_21411,N_20589);
and U23835 (N_23835,N_21695,N_21313);
and U23836 (N_23836,N_21571,N_21892);
and U23837 (N_23837,N_20567,N_21192);
or U23838 (N_23838,N_21957,N_20051);
xnor U23839 (N_23839,N_20221,N_21338);
nand U23840 (N_23840,N_21418,N_21931);
nand U23841 (N_23841,N_21251,N_21696);
xnor U23842 (N_23842,N_21664,N_21760);
and U23843 (N_23843,N_21830,N_21363);
xnor U23844 (N_23844,N_20760,N_21938);
nor U23845 (N_23845,N_21447,N_20376);
or U23846 (N_23846,N_21260,N_20323);
and U23847 (N_23847,N_20025,N_21567);
nand U23848 (N_23848,N_21563,N_21627);
and U23849 (N_23849,N_20884,N_21411);
and U23850 (N_23850,N_21957,N_20763);
nor U23851 (N_23851,N_21780,N_21826);
nor U23852 (N_23852,N_21353,N_21785);
xnor U23853 (N_23853,N_21139,N_21216);
and U23854 (N_23854,N_21884,N_21860);
xor U23855 (N_23855,N_20726,N_21074);
and U23856 (N_23856,N_20357,N_21438);
and U23857 (N_23857,N_21696,N_21474);
nor U23858 (N_23858,N_21257,N_20692);
xnor U23859 (N_23859,N_20518,N_20713);
nor U23860 (N_23860,N_20584,N_21608);
xnor U23861 (N_23861,N_21016,N_20713);
nand U23862 (N_23862,N_20798,N_20564);
xnor U23863 (N_23863,N_20488,N_21692);
and U23864 (N_23864,N_20764,N_21939);
nor U23865 (N_23865,N_21115,N_20808);
xnor U23866 (N_23866,N_20297,N_20436);
nand U23867 (N_23867,N_20773,N_20990);
xnor U23868 (N_23868,N_21934,N_21856);
and U23869 (N_23869,N_21682,N_20406);
nor U23870 (N_23870,N_20701,N_21783);
or U23871 (N_23871,N_21572,N_21412);
nor U23872 (N_23872,N_20576,N_20152);
xor U23873 (N_23873,N_21778,N_21735);
or U23874 (N_23874,N_21975,N_21361);
nor U23875 (N_23875,N_20688,N_20753);
xnor U23876 (N_23876,N_20517,N_21670);
and U23877 (N_23877,N_21476,N_21682);
or U23878 (N_23878,N_20983,N_21806);
or U23879 (N_23879,N_20840,N_21763);
and U23880 (N_23880,N_20244,N_21153);
or U23881 (N_23881,N_20427,N_21103);
xor U23882 (N_23882,N_21670,N_20772);
nor U23883 (N_23883,N_20187,N_20091);
nor U23884 (N_23884,N_21620,N_21056);
nor U23885 (N_23885,N_20110,N_21058);
xor U23886 (N_23886,N_20848,N_21042);
and U23887 (N_23887,N_20535,N_20708);
nand U23888 (N_23888,N_21445,N_20199);
and U23889 (N_23889,N_21741,N_21546);
nand U23890 (N_23890,N_20730,N_20300);
xor U23891 (N_23891,N_20995,N_20269);
and U23892 (N_23892,N_21427,N_20523);
nor U23893 (N_23893,N_21501,N_21075);
nor U23894 (N_23894,N_20268,N_20424);
xnor U23895 (N_23895,N_21101,N_20143);
and U23896 (N_23896,N_20682,N_20469);
nor U23897 (N_23897,N_20138,N_20511);
xnor U23898 (N_23898,N_20017,N_20182);
nand U23899 (N_23899,N_20303,N_21344);
nor U23900 (N_23900,N_20448,N_21492);
or U23901 (N_23901,N_20905,N_21940);
xnor U23902 (N_23902,N_20208,N_21725);
xnor U23903 (N_23903,N_20959,N_20338);
xnor U23904 (N_23904,N_20612,N_21362);
xnor U23905 (N_23905,N_21054,N_21427);
nand U23906 (N_23906,N_20895,N_20566);
or U23907 (N_23907,N_21530,N_21152);
xnor U23908 (N_23908,N_20212,N_21136);
nor U23909 (N_23909,N_20325,N_21864);
and U23910 (N_23910,N_20905,N_20630);
nand U23911 (N_23911,N_21289,N_20832);
nand U23912 (N_23912,N_20772,N_20662);
xnor U23913 (N_23913,N_21984,N_20521);
nor U23914 (N_23914,N_21602,N_21835);
or U23915 (N_23915,N_21285,N_21784);
and U23916 (N_23916,N_21079,N_21375);
and U23917 (N_23917,N_21124,N_20432);
xnor U23918 (N_23918,N_21769,N_20165);
nor U23919 (N_23919,N_21023,N_21194);
and U23920 (N_23920,N_20793,N_20853);
nor U23921 (N_23921,N_20969,N_21892);
xnor U23922 (N_23922,N_20297,N_21876);
and U23923 (N_23923,N_20975,N_20007);
nand U23924 (N_23924,N_21019,N_20909);
and U23925 (N_23925,N_21225,N_20433);
or U23926 (N_23926,N_20676,N_20709);
nor U23927 (N_23927,N_21275,N_20892);
and U23928 (N_23928,N_20900,N_21590);
nand U23929 (N_23929,N_20785,N_20411);
nand U23930 (N_23930,N_21200,N_21466);
nand U23931 (N_23931,N_20542,N_20421);
nand U23932 (N_23932,N_21850,N_21249);
xor U23933 (N_23933,N_20920,N_21989);
nand U23934 (N_23934,N_21869,N_20149);
nand U23935 (N_23935,N_20511,N_21754);
or U23936 (N_23936,N_21542,N_21786);
or U23937 (N_23937,N_21305,N_21953);
nand U23938 (N_23938,N_20721,N_21845);
or U23939 (N_23939,N_21284,N_20090);
nor U23940 (N_23940,N_21050,N_20710);
and U23941 (N_23941,N_21475,N_21385);
nand U23942 (N_23942,N_20063,N_20936);
or U23943 (N_23943,N_20943,N_20198);
nand U23944 (N_23944,N_20662,N_20682);
or U23945 (N_23945,N_20809,N_20391);
nand U23946 (N_23946,N_21942,N_21993);
and U23947 (N_23947,N_20391,N_21741);
xnor U23948 (N_23948,N_21293,N_20088);
nand U23949 (N_23949,N_20702,N_20246);
nand U23950 (N_23950,N_20816,N_21725);
nand U23951 (N_23951,N_21210,N_20244);
or U23952 (N_23952,N_20112,N_20526);
xor U23953 (N_23953,N_21804,N_21769);
nand U23954 (N_23954,N_20756,N_20128);
xor U23955 (N_23955,N_21537,N_20263);
nand U23956 (N_23956,N_20317,N_20630);
xor U23957 (N_23957,N_20909,N_20606);
and U23958 (N_23958,N_20458,N_20002);
nor U23959 (N_23959,N_21476,N_21010);
xor U23960 (N_23960,N_21857,N_21724);
xor U23961 (N_23961,N_21784,N_20425);
nand U23962 (N_23962,N_20056,N_20579);
nor U23963 (N_23963,N_21710,N_21602);
and U23964 (N_23964,N_21062,N_20315);
and U23965 (N_23965,N_20864,N_20492);
or U23966 (N_23966,N_21961,N_20774);
xor U23967 (N_23967,N_21632,N_20587);
or U23968 (N_23968,N_20888,N_21934);
or U23969 (N_23969,N_21795,N_21288);
or U23970 (N_23970,N_21592,N_21849);
xor U23971 (N_23971,N_20597,N_21844);
and U23972 (N_23972,N_20323,N_21072);
and U23973 (N_23973,N_20514,N_20360);
nor U23974 (N_23974,N_20267,N_20105);
and U23975 (N_23975,N_21402,N_20657);
nand U23976 (N_23976,N_20122,N_20768);
nor U23977 (N_23977,N_21709,N_21042);
xnor U23978 (N_23978,N_20795,N_21789);
nor U23979 (N_23979,N_20932,N_21762);
nand U23980 (N_23980,N_20722,N_21719);
xnor U23981 (N_23981,N_20922,N_20992);
nand U23982 (N_23982,N_20945,N_21556);
and U23983 (N_23983,N_21498,N_20680);
nor U23984 (N_23984,N_21454,N_20492);
xnor U23985 (N_23985,N_21395,N_21214);
nor U23986 (N_23986,N_20514,N_20960);
xnor U23987 (N_23987,N_20820,N_20217);
xnor U23988 (N_23988,N_21532,N_20344);
or U23989 (N_23989,N_21804,N_20519);
and U23990 (N_23990,N_20720,N_21741);
nor U23991 (N_23991,N_21851,N_20836);
nand U23992 (N_23992,N_21159,N_21510);
and U23993 (N_23993,N_21090,N_21393);
and U23994 (N_23994,N_21628,N_21098);
xor U23995 (N_23995,N_21609,N_21314);
nand U23996 (N_23996,N_21856,N_20112);
xor U23997 (N_23997,N_21996,N_20267);
or U23998 (N_23998,N_21417,N_20132);
and U23999 (N_23999,N_20691,N_21950);
nand U24000 (N_24000,N_22112,N_22899);
xor U24001 (N_24001,N_22862,N_23715);
nor U24002 (N_24002,N_22333,N_23344);
nor U24003 (N_24003,N_23847,N_23665);
nand U24004 (N_24004,N_22963,N_22053);
xor U24005 (N_24005,N_23519,N_22662);
nand U24006 (N_24006,N_22213,N_22378);
and U24007 (N_24007,N_22238,N_23582);
and U24008 (N_24008,N_22103,N_23701);
and U24009 (N_24009,N_23013,N_22480);
and U24010 (N_24010,N_22125,N_22806);
and U24011 (N_24011,N_23565,N_22031);
and U24012 (N_24012,N_23779,N_23671);
nor U24013 (N_24013,N_22715,N_23879);
and U24014 (N_24014,N_23462,N_23523);
and U24015 (N_24015,N_22878,N_22924);
xnor U24016 (N_24016,N_22360,N_23777);
nand U24017 (N_24017,N_23303,N_23995);
and U24018 (N_24018,N_23645,N_22381);
or U24019 (N_24019,N_22558,N_22855);
xnor U24020 (N_24020,N_23142,N_23722);
nor U24021 (N_24021,N_23283,N_22597);
nor U24022 (N_24022,N_23255,N_23162);
and U24023 (N_24023,N_23504,N_22292);
nand U24024 (N_24024,N_23257,N_23328);
or U24025 (N_24025,N_23029,N_23123);
nand U24026 (N_24026,N_22580,N_23003);
and U24027 (N_24027,N_23108,N_22714);
nand U24028 (N_24028,N_23648,N_23903);
xnor U24029 (N_24029,N_23992,N_23015);
nand U24030 (N_24030,N_23343,N_23240);
and U24031 (N_24031,N_22481,N_23429);
and U24032 (N_24032,N_22359,N_22854);
or U24033 (N_24033,N_23619,N_23865);
and U24034 (N_24034,N_22844,N_23980);
xor U24035 (N_24035,N_22497,N_23376);
or U24036 (N_24036,N_22107,N_23120);
xnor U24037 (N_24037,N_22118,N_22690);
nor U24038 (N_24038,N_23734,N_23791);
and U24039 (N_24039,N_23944,N_22262);
or U24040 (N_24040,N_23494,N_23401);
nor U24041 (N_24041,N_23489,N_22323);
xor U24042 (N_24042,N_23712,N_23687);
nand U24043 (N_24043,N_22958,N_22484);
nand U24044 (N_24044,N_22172,N_22135);
and U24045 (N_24045,N_22666,N_23087);
or U24046 (N_24046,N_22077,N_22365);
nor U24047 (N_24047,N_22021,N_22098);
and U24048 (N_24048,N_22167,N_22014);
or U24049 (N_24049,N_23972,N_22256);
nor U24050 (N_24050,N_23846,N_22618);
nor U24051 (N_24051,N_23655,N_23964);
or U24052 (N_24052,N_23124,N_23908);
and U24053 (N_24053,N_23402,N_22459);
and U24054 (N_24054,N_23993,N_22850);
nor U24055 (N_24055,N_23857,N_23322);
nand U24056 (N_24056,N_23593,N_23793);
nor U24057 (N_24057,N_22034,N_23078);
and U24058 (N_24058,N_22095,N_22489);
nand U24059 (N_24059,N_22569,N_23056);
and U24060 (N_24060,N_23533,N_22140);
nand U24061 (N_24061,N_23602,N_23911);
nand U24062 (N_24062,N_22069,N_23295);
xnor U24063 (N_24063,N_23484,N_22725);
xnor U24064 (N_24064,N_22450,N_22173);
and U24065 (N_24065,N_22555,N_22830);
or U24066 (N_24066,N_23566,N_23986);
and U24067 (N_24067,N_23555,N_22158);
nand U24068 (N_24068,N_22287,N_23158);
nand U24069 (N_24069,N_22334,N_22275);
xor U24070 (N_24070,N_22430,N_22609);
nand U24071 (N_24071,N_22841,N_22169);
nand U24072 (N_24072,N_22039,N_22265);
nor U24073 (N_24073,N_22982,N_23042);
and U24074 (N_24074,N_22547,N_23785);
and U24075 (N_24075,N_23904,N_23239);
nand U24076 (N_24076,N_22196,N_22394);
xor U24077 (N_24077,N_22419,N_23443);
or U24078 (N_24078,N_22961,N_22584);
nor U24079 (N_24079,N_23890,N_22945);
nand U24080 (N_24080,N_22222,N_22980);
nor U24081 (N_24081,N_22412,N_23318);
xor U24082 (N_24082,N_22691,N_23906);
nor U24083 (N_24083,N_22499,N_22187);
and U24084 (N_24084,N_22444,N_23235);
and U24085 (N_24085,N_23333,N_22303);
nand U24086 (N_24086,N_23020,N_23973);
nor U24087 (N_24087,N_22722,N_23083);
or U24088 (N_24088,N_23098,N_23189);
and U24089 (N_24089,N_22792,N_22373);
nand U24090 (N_24090,N_22244,N_23615);
nor U24091 (N_24091,N_23134,N_23735);
or U24092 (N_24092,N_23392,N_22035);
and U24093 (N_24093,N_22608,N_23348);
nand U24094 (N_24094,N_23515,N_22583);
and U24095 (N_24095,N_23104,N_22403);
xor U24096 (N_24096,N_22563,N_23644);
nor U24097 (N_24097,N_22994,N_22747);
and U24098 (N_24098,N_22768,N_22553);
nor U24099 (N_24099,N_23997,N_22533);
nor U24100 (N_24100,N_22905,N_22425);
nor U24101 (N_24101,N_22174,N_22696);
nor U24102 (N_24102,N_22559,N_23834);
nor U24103 (N_24103,N_22352,N_22078);
nor U24104 (N_24104,N_22847,N_22882);
or U24105 (N_24105,N_23856,N_23096);
or U24106 (N_24106,N_23902,N_22818);
nor U24107 (N_24107,N_22976,N_23048);
and U24108 (N_24108,N_23688,N_22826);
xor U24109 (N_24109,N_23070,N_23814);
and U24110 (N_24110,N_23365,N_22736);
or U24111 (N_24111,N_22354,N_23741);
xnor U24112 (N_24112,N_23739,N_23046);
nor U24113 (N_24113,N_23469,N_23706);
or U24114 (N_24114,N_22417,N_22979);
and U24115 (N_24115,N_23625,N_23636);
nand U24116 (N_24116,N_22508,N_22258);
nand U24117 (N_24117,N_22898,N_23862);
or U24118 (N_24118,N_22442,N_23957);
nand U24119 (N_24119,N_22250,N_22219);
nand U24120 (N_24120,N_23710,N_22236);
nand U24121 (N_24121,N_22543,N_22008);
nor U24122 (N_24122,N_23362,N_23642);
or U24123 (N_24123,N_22253,N_23586);
or U24124 (N_24124,N_23258,N_22900);
or U24125 (N_24125,N_22134,N_22539);
or U24126 (N_24126,N_22097,N_23653);
nand U24127 (N_24127,N_22755,N_23437);
nor U24128 (N_24128,N_22279,N_22805);
nor U24129 (N_24129,N_22019,N_22392);
or U24130 (N_24130,N_22398,N_22990);
xor U24131 (N_24131,N_23787,N_22965);
and U24132 (N_24132,N_22717,N_22205);
or U24133 (N_24133,N_23799,N_22320);
or U24134 (N_24134,N_23552,N_23691);
nand U24135 (N_24135,N_23617,N_22836);
xnor U24136 (N_24136,N_22310,N_22564);
nor U24137 (N_24137,N_23403,N_23026);
nor U24138 (N_24138,N_22797,N_23037);
or U24139 (N_24139,N_22502,N_23019);
or U24140 (N_24140,N_23171,N_23749);
xor U24141 (N_24141,N_23748,N_22374);
and U24142 (N_24142,N_23596,N_23971);
and U24143 (N_24143,N_22124,N_23650);
or U24144 (N_24144,N_22052,N_23010);
nand U24145 (N_24145,N_23448,N_22734);
nand U24146 (N_24146,N_23505,N_23346);
xnor U24147 (N_24147,N_22577,N_23826);
nor U24148 (N_24148,N_23413,N_22094);
or U24149 (N_24149,N_23962,N_23990);
nor U24150 (N_24150,N_22991,N_22541);
or U24151 (N_24151,N_22835,N_23601);
xnor U24152 (N_24152,N_22109,N_23639);
or U24153 (N_24153,N_22535,N_23666);
nor U24154 (N_24154,N_23140,N_23440);
nand U24155 (N_24155,N_23316,N_23921);
xnor U24156 (N_24156,N_22877,N_22627);
xor U24157 (N_24157,N_23304,N_22730);
xor U24158 (N_24158,N_23975,N_22229);
nand U24159 (N_24159,N_23811,N_22908);
nor U24160 (N_24160,N_22698,N_22446);
xnor U24161 (N_24161,N_22099,N_23781);
nand U24162 (N_24162,N_23782,N_22410);
nor U24163 (N_24163,N_23294,N_23631);
xor U24164 (N_24164,N_23521,N_23790);
nand U24165 (N_24165,N_22232,N_22353);
and U24166 (N_24166,N_22170,N_22482);
nand U24167 (N_24167,N_23589,N_22514);
and U24168 (N_24168,N_23251,N_23807);
xor U24169 (N_24169,N_22672,N_23212);
nand U24170 (N_24170,N_22478,N_22308);
xnor U24171 (N_24171,N_23732,N_22267);
nand U24172 (N_24172,N_22567,N_23233);
nor U24173 (N_24173,N_22534,N_22026);
nor U24174 (N_24174,N_22131,N_23125);
and U24175 (N_24175,N_23424,N_22351);
nand U24176 (N_24176,N_23496,N_23770);
and U24177 (N_24177,N_23998,N_23062);
xnor U24178 (N_24178,N_22576,N_23818);
xor U24179 (N_24179,N_22944,N_22494);
nor U24180 (N_24180,N_23486,N_22466);
nand U24181 (N_24181,N_22814,N_22677);
nand U24182 (N_24182,N_22361,N_23977);
nand U24183 (N_24183,N_23340,N_22313);
xor U24184 (N_24184,N_23514,N_23036);
nand U24185 (N_24185,N_22380,N_22336);
or U24186 (N_24186,N_22063,N_22532);
nor U24187 (N_24187,N_23680,N_22753);
xor U24188 (N_24188,N_22309,N_23778);
and U24189 (N_24189,N_22975,N_23752);
nor U24190 (N_24190,N_22550,N_23032);
nor U24191 (N_24191,N_22654,N_23827);
and U24192 (N_24192,N_22537,N_23941);
nand U24193 (N_24193,N_22637,N_22349);
xor U24194 (N_24194,N_23077,N_22810);
xor U24195 (N_24195,N_23358,N_22289);
nor U24196 (N_24196,N_23963,N_22556);
nor U24197 (N_24197,N_22795,N_22757);
or U24198 (N_24198,N_23305,N_22782);
or U24199 (N_24199,N_23634,N_22363);
nor U24200 (N_24200,N_23468,N_23877);
nand U24201 (N_24201,N_23268,N_23564);
or U24202 (N_24202,N_22732,N_22910);
or U24203 (N_24203,N_23766,N_23409);
xor U24204 (N_24204,N_22959,N_23111);
xnor U24205 (N_24205,N_22033,N_22355);
or U24206 (N_24206,N_23720,N_23767);
xnor U24207 (N_24207,N_22195,N_23580);
nor U24208 (N_24208,N_22366,N_22004);
and U24209 (N_24209,N_23823,N_23508);
nor U24210 (N_24210,N_23398,N_23873);
nor U24211 (N_24211,N_22611,N_22827);
and U24212 (N_24212,N_23430,N_22492);
or U24213 (N_24213,N_23090,N_23916);
nand U24214 (N_24214,N_22621,N_22766);
nand U24215 (N_24215,N_23058,N_22137);
nand U24216 (N_24216,N_22857,N_22426);
or U24217 (N_24217,N_22807,N_23133);
or U24218 (N_24218,N_23272,N_23273);
or U24219 (N_24219,N_22325,N_22969);
or U24220 (N_24220,N_22274,N_23422);
nand U24221 (N_24221,N_23837,N_23176);
nor U24222 (N_24222,N_22479,N_23731);
and U24223 (N_24223,N_23236,N_22694);
nand U24224 (N_24224,N_23981,N_23578);
or U24225 (N_24225,N_22752,N_23946);
xnor U24226 (N_24226,N_22938,N_22467);
or U24227 (N_24227,N_22346,N_22064);
and U24228 (N_24228,N_22909,N_23892);
nor U24229 (N_24229,N_22529,N_23547);
and U24230 (N_24230,N_22184,N_22188);
or U24231 (N_24231,N_23756,N_22051);
xnor U24232 (N_24232,N_22096,N_23672);
nor U24233 (N_24233,N_22610,N_22458);
xnor U24234 (N_24234,N_22973,N_22845);
xor U24235 (N_24235,N_23792,N_22895);
nand U24236 (N_24236,N_23520,N_22946);
nor U24237 (N_24237,N_22290,N_23727);
xnor U24238 (N_24238,N_23612,N_23454);
and U24239 (N_24239,N_22922,N_23394);
or U24240 (N_24240,N_23016,N_23541);
nor U24241 (N_24241,N_23385,N_22212);
or U24242 (N_24242,N_22582,N_23896);
nor U24243 (N_24243,N_22340,N_22306);
nor U24244 (N_24244,N_22186,N_23412);
and U24245 (N_24245,N_22524,N_22831);
xnor U24246 (N_24246,N_22798,N_23187);
or U24247 (N_24247,N_23050,N_23869);
nand U24248 (N_24248,N_22781,N_22156);
and U24249 (N_24249,N_22804,N_22935);
or U24250 (N_24250,N_23775,N_23771);
and U24251 (N_24251,N_22822,N_23325);
or U24252 (N_24252,N_23806,N_23186);
xnor U24253 (N_24253,N_23185,N_23053);
nor U24254 (N_24254,N_22257,N_22987);
nand U24255 (N_24255,N_22121,N_23945);
or U24256 (N_24256,N_22964,N_23607);
or U24257 (N_24257,N_23389,N_22180);
or U24258 (N_24258,N_23485,N_22668);
xnor U24259 (N_24259,N_23417,N_22389);
and U24260 (N_24260,N_22950,N_23353);
nand U24261 (N_24261,N_22120,N_23191);
xnor U24262 (N_24262,N_23449,N_23065);
or U24263 (N_24263,N_23571,N_22276);
or U24264 (N_24264,N_23632,N_23658);
or U24265 (N_24265,N_23878,N_22476);
nor U24266 (N_24266,N_23306,N_23947);
and U24267 (N_24267,N_22472,N_23382);
xor U24268 (N_24268,N_22228,N_23097);
nand U24269 (N_24269,N_22387,N_23428);
nor U24270 (N_24270,N_22375,N_22903);
nor U24271 (N_24271,N_22519,N_22345);
nand U24272 (N_24272,N_23319,N_22491);
nor U24273 (N_24273,N_23664,N_23587);
or U24274 (N_24274,N_22316,N_23201);
xor U24275 (N_24275,N_22144,N_23024);
nand U24276 (N_24276,N_22161,N_23479);
and U24277 (N_24277,N_22382,N_23717);
and U24278 (N_24278,N_23418,N_23359);
nor U24279 (N_24279,N_23844,N_23331);
or U24280 (N_24280,N_23788,N_23374);
nand U24281 (N_24281,N_23516,N_22934);
or U24282 (N_24282,N_23491,N_23008);
xor U24283 (N_24283,N_22155,N_22673);
or U24284 (N_24284,N_22220,N_22940);
or U24285 (N_24285,N_23184,N_23935);
nand U24286 (N_24286,N_22803,N_22194);
nand U24287 (N_24287,N_22679,N_23646);
nor U24288 (N_24288,N_23853,N_22277);
or U24289 (N_24289,N_22506,N_23202);
xor U24290 (N_24290,N_22025,N_22202);
or U24291 (N_24291,N_22415,N_23859);
xor U24292 (N_24292,N_23982,N_22544);
and U24293 (N_24293,N_23072,N_22066);
and U24294 (N_24294,N_22695,N_23408);
xor U24295 (N_24295,N_22867,N_22809);
nor U24296 (N_24296,N_22931,N_22246);
nor U24297 (N_24297,N_23746,N_22347);
nand U24298 (N_24298,N_23527,N_22581);
nor U24299 (N_24299,N_23014,N_23622);
and U24300 (N_24300,N_23728,N_23657);
or U24301 (N_24301,N_22764,N_23164);
and U24302 (N_24302,N_22210,N_22858);
and U24303 (N_24303,N_22045,N_22302);
xor U24304 (N_24304,N_22438,N_22061);
or U24305 (N_24305,N_22468,N_23545);
or U24306 (N_24306,N_22620,N_23754);
and U24307 (N_24307,N_22086,N_22676);
or U24308 (N_24308,N_22082,N_22475);
and U24309 (N_24309,N_22861,N_22328);
and U24310 (N_24310,N_23914,N_23931);
nand U24311 (N_24311,N_22384,N_23923);
or U24312 (N_24312,N_23425,N_22074);
nand U24313 (N_24313,N_23828,N_22744);
and U24314 (N_24314,N_22105,N_22528);
nor U24315 (N_24315,N_23030,N_22248);
nor U24316 (N_24316,N_22549,N_23167);
nor U24317 (N_24317,N_23172,N_22998);
nand U24318 (N_24318,N_23699,N_23606);
nand U24319 (N_24319,N_22068,N_22562);
nand U24320 (N_24320,N_22988,N_22159);
xor U24321 (N_24321,N_22911,N_22511);
or U24322 (N_24322,N_23116,N_23351);
xnor U24323 (N_24323,N_22111,N_23106);
xor U24324 (N_24324,N_23915,N_22602);
nand U24325 (N_24325,N_23222,N_23949);
nand U24326 (N_24326,N_22326,N_23802);
xor U24327 (N_24327,N_22299,N_22441);
xor U24328 (N_24328,N_22707,N_22293);
xnor U24329 (N_24329,N_23461,N_22759);
or U24330 (N_24330,N_23027,N_23928);
and U24331 (N_24331,N_22593,N_22925);
xnor U24332 (N_24332,N_22190,N_22727);
nor U24333 (N_24333,N_22552,N_23432);
nand U24334 (N_24334,N_22568,N_23157);
and U24335 (N_24335,N_22490,N_23228);
nor U24336 (N_24336,N_23180,N_22525);
or U24337 (N_24337,N_22162,N_23543);
or U24338 (N_24338,N_23289,N_23808);
and U24339 (N_24339,N_23934,N_22623);
nor U24340 (N_24340,N_23721,N_23663);
and U24341 (N_24341,N_23868,N_22728);
nor U24342 (N_24342,N_22050,N_22960);
or U24343 (N_24343,N_23511,N_23965);
nor U24344 (N_24344,N_22197,N_22907);
xnor U24345 (N_24345,N_22780,N_23246);
or U24346 (N_24346,N_23588,N_22136);
xnor U24347 (N_24347,N_23446,N_22070);
or U24348 (N_24348,N_23161,N_23870);
nand U24349 (N_24349,N_23913,N_22284);
and U24350 (N_24350,N_22619,N_23166);
or U24351 (N_24351,N_22800,N_22047);
nor U24352 (N_24352,N_22974,N_23668);
or U24353 (N_24353,N_22551,N_22590);
xnor U24354 (N_24354,N_22904,N_22166);
nand U24355 (N_24355,N_23307,N_22860);
and U24356 (N_24356,N_22680,N_22642);
or U24357 (N_24357,N_23849,N_22407);
xnor U24358 (N_24358,N_23920,N_23135);
or U24359 (N_24359,N_23917,N_22385);
or U24360 (N_24360,N_23276,N_22084);
nor U24361 (N_24361,N_22784,N_22054);
and U24362 (N_24362,N_23576,N_22294);
nand U24363 (N_24363,N_23023,N_23047);
nand U24364 (N_24364,N_22408,N_23570);
and U24365 (N_24365,N_23832,N_22364);
xor U24366 (N_24366,N_23259,N_22887);
nand U24367 (N_24367,N_23009,N_23378);
or U24368 (N_24368,N_22003,N_22080);
nor U24369 (N_24369,N_23585,N_23410);
xor U24370 (N_24370,N_23705,N_23453);
xnor U24371 (N_24371,N_22874,N_22143);
nor U24372 (N_24372,N_23758,N_22215);
xor U24373 (N_24373,N_23460,N_23279);
or U24374 (N_24374,N_22414,N_23375);
or U24375 (N_24375,N_22996,N_22036);
or U24376 (N_24376,N_23616,N_23614);
xnor U24377 (N_24377,N_23144,N_23885);
nor U24378 (N_24378,N_23620,N_23815);
nor U24379 (N_24379,N_22132,N_23136);
and U24380 (N_24380,N_22587,N_22044);
xnor U24381 (N_24381,N_23208,N_22866);
and U24382 (N_24382,N_23232,N_23886);
or U24383 (N_24383,N_23840,N_23299);
nor U24384 (N_24384,N_22972,N_22647);
nand U24385 (N_24385,N_22139,N_23603);
nor U24386 (N_24386,N_22329,N_22702);
or U24387 (N_24387,N_23127,N_22794);
nand U24388 (N_24388,N_23347,N_23247);
nand U24389 (N_24389,N_23107,N_22104);
nand U24390 (N_24390,N_23060,N_22182);
xnor U24391 (N_24391,N_22496,N_22526);
nor U24392 (N_24392,N_23229,N_22625);
and U24393 (N_24393,N_22343,N_22765);
and U24394 (N_24394,N_23761,N_23293);
nor U24395 (N_24395,N_22779,N_22585);
nand U24396 (N_24396,N_22540,N_22149);
and U24397 (N_24397,N_23649,N_22929);
or U24398 (N_24398,N_22049,N_22208);
xnor U24399 (N_24399,N_23260,N_22330);
and U24400 (N_24400,N_22641,N_22761);
nand U24401 (N_24401,N_22775,N_22503);
and U24402 (N_24402,N_22406,N_22242);
nor U24403 (N_24403,N_23237,N_22571);
or U24404 (N_24404,N_23141,N_22421);
xor U24405 (N_24405,N_22470,N_22684);
xor U24406 (N_24406,N_23948,N_22009);
and U24407 (N_24407,N_23031,N_23457);
and U24408 (N_24408,N_23447,N_23226);
xnor U24409 (N_24409,N_23231,N_23804);
xor U24410 (N_24410,N_23464,N_22500);
and U24411 (N_24411,N_23656,N_23909);
nand U24412 (N_24412,N_23381,N_23891);
or U24413 (N_24413,N_23824,N_23597);
nand U24414 (N_24414,N_23415,N_23128);
nor U24415 (N_24415,N_22423,N_23531);
and U24416 (N_24416,N_23436,N_23338);
nand U24417 (N_24417,N_23502,N_22834);
or U24418 (N_24418,N_22314,N_22870);
nand U24419 (N_24419,N_23548,N_23079);
nand U24420 (N_24420,N_23796,N_22443);
nor U24421 (N_24421,N_22282,N_22092);
xnor U24422 (N_24422,N_23575,N_22591);
and U24423 (N_24423,N_23894,N_23843);
and U24424 (N_24424,N_22088,N_22216);
and U24425 (N_24425,N_23354,N_22073);
or U24426 (N_24426,N_22640,N_23472);
and U24427 (N_24427,N_22918,N_23159);
nor U24428 (N_24428,N_23471,N_23757);
nor U24429 (N_24429,N_22914,N_22016);
nor U24430 (N_24430,N_22772,N_22356);
xor U24431 (N_24431,N_23218,N_22157);
nor U24432 (N_24432,N_23590,N_22886);
xnor U24433 (N_24433,N_23776,N_22337);
nand U24434 (N_24434,N_22894,N_22889);
and U24435 (N_24435,N_23759,N_22655);
xnor U24436 (N_24436,N_23966,N_23433);
xor U24437 (N_24437,N_23339,N_23794);
nand U24438 (N_24438,N_23181,N_22967);
xnor U24439 (N_24439,N_23080,N_23309);
and U24440 (N_24440,N_22667,N_22864);
or U24441 (N_24441,N_22520,N_23985);
and U24442 (N_24442,N_23483,N_22659);
xor U24443 (N_24443,N_22418,N_22891);
nor U24444 (N_24444,N_22607,N_23155);
and U24445 (N_24445,N_23740,N_22350);
nor U24446 (N_24446,N_23284,N_23193);
nand U24447 (N_24447,N_23487,N_23373);
xnor U24448 (N_24448,N_22735,N_22951);
and U24449 (N_24449,N_23943,N_22439);
or U24450 (N_24450,N_22601,N_23326);
and U24451 (N_24451,N_22207,N_22454);
or U24452 (N_24452,N_23320,N_23940);
xnor U24453 (N_24453,N_23395,N_22181);
or U24454 (N_24454,N_23988,N_22840);
or U24455 (N_24455,N_22400,N_22079);
or U24456 (N_24456,N_23989,N_22636);
nor U24457 (N_24457,N_23352,N_23608);
or U24458 (N_24458,N_22941,N_22327);
nor U24459 (N_24459,N_22379,N_23881);
nand U24460 (N_24460,N_22661,N_22332);
nor U24461 (N_24461,N_22037,N_22448);
and U24462 (N_24462,N_22395,N_22175);
nor U24463 (N_24463,N_23022,N_23101);
and U24464 (N_24464,N_23368,N_22335);
nor U24465 (N_24465,N_23300,N_23091);
nor U24466 (N_24466,N_22065,N_22291);
or U24467 (N_24467,N_23216,N_22260);
and U24468 (N_24468,N_22505,N_22370);
nand U24469 (N_24469,N_23188,N_23220);
xnor U24470 (N_24470,N_23558,N_22341);
and U24471 (N_24471,N_23540,N_22815);
or U24472 (N_24472,N_22981,N_22763);
nand U24473 (N_24473,N_23704,N_23298);
nand U24474 (N_24474,N_23420,N_22966);
nand U24475 (N_24475,N_23290,N_23482);
xor U24476 (N_24476,N_23900,N_23387);
nor U24477 (N_24477,N_23635,N_23130);
or U24478 (N_24478,N_23979,N_22820);
nand U24479 (N_24479,N_23855,N_22513);
nor U24480 (N_24480,N_23476,N_22594);
xor U24481 (N_24481,N_23081,N_23377);
nand U24482 (N_24482,N_23768,N_23423);
and U24483 (N_24483,N_23152,N_22193);
and U24484 (N_24484,N_23040,N_22849);
nand U24485 (N_24485,N_22487,N_22778);
or U24486 (N_24486,N_23984,N_23711);
and U24487 (N_24487,N_22040,N_22977);
nor U24488 (N_24488,N_23196,N_22437);
xnor U24489 (N_24489,N_22665,N_23114);
nor U24490 (N_24490,N_22739,N_23059);
nand U24491 (N_24491,N_23169,N_22399);
nor U24492 (N_24492,N_23953,N_23380);
nor U24493 (N_24493,N_23694,N_23207);
and U24494 (N_24494,N_23061,N_23473);
or U24495 (N_24495,N_23490,N_23951);
xnor U24496 (N_24496,N_22252,N_22455);
and U24497 (N_24497,N_23875,N_23675);
nand U24498 (N_24498,N_22776,N_23275);
or U24499 (N_24499,N_22606,N_22671);
nand U24500 (N_24500,N_23506,N_22829);
nand U24501 (N_24501,N_22912,N_23282);
nand U24502 (N_24502,N_22152,N_23366);
xnor U24503 (N_24503,N_22984,N_22055);
and U24504 (N_24504,N_22992,N_22843);
nor U24505 (N_24505,N_23274,N_23341);
xnor U24506 (N_24506,N_23241,N_22595);
nand U24507 (N_24507,N_23638,N_22791);
nor U24508 (N_24508,N_22390,N_22978);
nor U24509 (N_24509,N_22114,N_23498);
nor U24510 (N_24510,N_22575,N_23952);
nor U24511 (N_24511,N_22785,N_22522);
nand U24512 (N_24512,N_22129,N_22832);
or U24513 (N_24513,N_23474,N_23442);
or U24514 (N_24514,N_23765,N_22011);
and U24515 (N_24515,N_22243,N_23544);
xor U24516 (N_24516,N_22937,N_23383);
nand U24517 (N_24517,N_22756,N_23678);
xor U24518 (N_24518,N_22823,N_23534);
and U24519 (N_24519,N_22317,N_23831);
xnor U24520 (N_24520,N_22300,N_23335);
and U24521 (N_24521,N_22871,N_22561);
nor U24522 (N_24522,N_22402,N_22957);
or U24523 (N_24523,N_22865,N_23066);
nor U24524 (N_24524,N_23110,N_22932);
and U24525 (N_24525,N_22177,N_23163);
or U24526 (N_24526,N_22001,N_22644);
nand U24527 (N_24527,N_22160,N_23129);
nand U24528 (N_24528,N_22102,N_23390);
nand U24529 (N_24529,N_23367,N_22718);
nand U24530 (N_24530,N_22163,N_22315);
nor U24531 (N_24531,N_23567,N_22268);
or U24532 (N_24532,N_23866,N_23113);
xnor U24533 (N_24533,N_22464,N_23160);
xor U24534 (N_24534,N_22851,N_23327);
and U24535 (N_24535,N_23197,N_22875);
or U24536 (N_24536,N_22751,N_22923);
nand U24537 (N_24537,N_22201,N_22209);
nand U24538 (N_24538,N_22023,N_22793);
nand U24539 (N_24539,N_22653,N_23266);
or U24540 (N_24540,N_23269,N_22447);
and U24541 (N_24541,N_22106,N_23700);
nor U24542 (N_24542,N_23291,N_22573);
or U24543 (N_24543,N_23407,N_23399);
and U24544 (N_24544,N_22812,N_22622);
nand U24545 (N_24545,N_23323,N_23507);
and U24546 (N_24546,N_22451,N_22218);
xnor U24547 (N_24547,N_23252,N_23497);
or U24548 (N_24548,N_23256,N_22926);
nor U24549 (N_24549,N_22726,N_22928);
nor U24550 (N_24550,N_23994,N_23702);
and U24551 (N_24551,N_22687,N_23261);
xnor U24552 (N_24552,N_23254,N_23005);
and U24553 (N_24553,N_22445,N_22678);
and U24554 (N_24554,N_23100,N_23224);
nor U24555 (N_24555,N_22032,N_23411);
nand U24556 (N_24556,N_23876,N_23899);
and U24557 (N_24557,N_23094,N_23139);
nand U24558 (N_24558,N_23204,N_23182);
xnor U24559 (N_24559,N_23809,N_22645);
nor U24560 (N_24560,N_22954,N_22530);
nor U24561 (N_24561,N_23249,N_23679);
or U24562 (N_24562,N_23719,N_23627);
nand U24563 (N_24563,N_23629,N_23686);
and U24564 (N_24564,N_23301,N_22178);
nor U24565 (N_24565,N_22404,N_22231);
xor U24566 (N_24566,N_23174,N_23961);
and U24567 (N_24567,N_22833,N_23084);
or U24568 (N_24568,N_23271,N_22515);
xnor U24569 (N_24569,N_22743,N_22245);
xor U24570 (N_24570,N_23102,N_22081);
xor U24571 (N_24571,N_22435,N_22516);
nand U24572 (N_24572,N_23388,N_22214);
and U24573 (N_24573,N_23810,N_22962);
and U24574 (N_24574,N_23044,N_22546);
xor U24575 (N_24575,N_22719,N_22872);
nand U24576 (N_24576,N_23848,N_22604);
xor U24577 (N_24577,N_23405,N_22372);
xor U24578 (N_24578,N_23747,N_23537);
nand U24579 (N_24579,N_22971,N_23234);
or U24580 (N_24580,N_23082,N_23591);
nand U24581 (N_24581,N_23086,N_23696);
and U24582 (N_24582,N_23604,N_23898);
nor U24583 (N_24583,N_22856,N_23598);
or U24584 (N_24584,N_22183,N_22113);
nand U24585 (N_24585,N_22255,N_23503);
nand U24586 (N_24586,N_22700,N_23991);
or U24587 (N_24587,N_23170,N_23500);
and U24588 (N_24588,N_22838,N_23277);
xor U24589 (N_24589,N_23025,N_22657);
or U24590 (N_24590,N_23970,N_22921);
nor U24591 (N_24591,N_23018,N_23554);
nor U24592 (N_24592,N_22062,N_23557);
or U24593 (N_24593,N_23526,N_23709);
nand U24594 (N_24594,N_22226,N_23292);
nand U24595 (N_24595,N_22397,N_23315);
and U24596 (N_24596,N_22474,N_23336);
and U24597 (N_24597,N_23628,N_23673);
or U24598 (N_24598,N_22767,N_22362);
nor U24599 (N_24599,N_23238,N_22906);
or U24600 (N_24600,N_22651,N_22773);
or U24601 (N_24601,N_23190,N_22367);
nand U24602 (N_24602,N_22386,N_23708);
xnor U24603 (N_24603,N_23613,N_23363);
nor U24604 (N_24604,N_23192,N_22706);
nor U24605 (N_24605,N_22897,N_22432);
nor U24606 (N_24606,N_23073,N_22902);
or U24607 (N_24607,N_22783,N_23835);
nand U24608 (N_24608,N_22709,N_23623);
nor U24609 (N_24609,N_23535,N_23912);
or U24610 (N_24610,N_22745,N_22884);
or U24611 (N_24611,N_22685,N_23099);
nor U24612 (N_24612,N_23021,N_23033);
nor U24613 (N_24613,N_23842,N_23350);
and U24614 (N_24614,N_22022,N_22796);
nor U24615 (N_24615,N_22204,N_23369);
xor U24616 (N_24616,N_22626,N_22087);
nor U24617 (N_24617,N_23074,N_23681);
and U24618 (N_24618,N_22828,N_23556);
or U24619 (N_24619,N_23830,N_22164);
and U24620 (N_24620,N_22704,N_23213);
nor U24621 (N_24621,N_22453,N_22296);
and U24622 (N_24622,N_22883,N_22123);
nand U24623 (N_24623,N_22574,N_23695);
xnor U24624 (N_24624,N_23764,N_22774);
xnor U24625 (N_24625,N_23974,N_23416);
and U24626 (N_24626,N_22554,N_22968);
xor U24627 (N_24627,N_23467,N_23280);
xnor U24628 (N_24628,N_23723,N_23248);
and U24629 (N_24629,N_23225,N_23332);
nand U24630 (N_24630,N_23007,N_23379);
or U24631 (N_24631,N_22072,N_22824);
xor U24632 (N_24632,N_23227,N_23901);
nor U24633 (N_24633,N_22357,N_23513);
xor U24634 (N_24634,N_23684,N_23250);
or U24635 (N_24635,N_22485,N_23041);
nand U24636 (N_24636,N_23813,N_22429);
nand U24637 (N_24637,N_23499,N_23745);
xor U24638 (N_24638,N_22788,N_23357);
xor U24639 (N_24639,N_22873,N_23147);
nand U24640 (N_24640,N_22281,N_22510);
xnor U24641 (N_24641,N_22682,N_23532);
and U24642 (N_24642,N_22885,N_22015);
nor U24643 (N_24643,N_22683,N_23451);
nand U24644 (N_24644,N_23337,N_23897);
xor U24645 (N_24645,N_22427,N_22119);
xnor U24646 (N_24646,N_22813,N_22712);
or U24647 (N_24647,N_23718,N_22191);
nand U24648 (N_24648,N_23450,N_22369);
xor U24649 (N_24649,N_22259,N_22239);
or U24650 (N_24650,N_22280,N_22638);
or U24651 (N_24651,N_23049,N_23780);
xor U24652 (N_24652,N_22311,N_23384);
nand U24653 (N_24653,N_22527,N_23889);
nor U24654 (N_24654,N_23605,N_22473);
nor U24655 (N_24655,N_22307,N_23528);
and U24656 (N_24656,N_22708,N_23334);
and U24657 (N_24657,N_23599,N_22786);
xnor U24658 (N_24658,N_23495,N_23154);
nor U24659 (N_24659,N_22927,N_23795);
or U24660 (N_24660,N_23643,N_23549);
and U24661 (N_24661,N_23397,N_22947);
xor U24662 (N_24662,N_22697,N_23119);
or U24663 (N_24663,N_23117,N_22126);
nor U24664 (N_24664,N_22041,N_22741);
nand U24665 (N_24665,N_23153,N_23214);
and U24666 (N_24666,N_23075,N_23851);
nor U24667 (N_24667,N_22057,N_22699);
or U24668 (N_24668,N_23199,N_23444);
xnor U24669 (N_24669,N_23054,N_23884);
and U24670 (N_24670,N_23624,N_23637);
nand U24671 (N_24671,N_22116,N_22091);
and U24672 (N_24672,N_22254,N_23478);
or U24673 (N_24673,N_22853,N_23165);
nand U24674 (N_24674,N_22770,N_23858);
and U24675 (N_24675,N_22076,N_23414);
nor U24676 (N_24676,N_22933,N_22319);
xor U24677 (N_24677,N_23441,N_23115);
nand U24678 (N_24678,N_22600,N_23034);
nor U24679 (N_24679,N_22028,N_23936);
nand U24680 (N_24680,N_22692,N_23342);
and U24681 (N_24681,N_23685,N_22542);
xnor U24682 (N_24682,N_23743,N_22876);
nor U24683 (N_24683,N_23051,N_22024);
nand U24684 (N_24684,N_22154,N_22842);
or U24685 (N_24685,N_23463,N_22338);
or U24686 (N_24686,N_22557,N_23751);
xor U24687 (N_24687,N_23286,N_23317);
or U24688 (N_24688,N_22913,N_23067);
xnor U24689 (N_24689,N_23435,N_22295);
and U24690 (N_24690,N_22531,N_23011);
or U24691 (N_24691,N_22322,N_22298);
nor U24692 (N_24692,N_22225,N_22789);
nor U24693 (N_24693,N_23297,N_22461);
nor U24694 (N_24694,N_23922,N_22811);
xor U24695 (N_24695,N_22750,N_23179);
and U24696 (N_24696,N_22486,N_22235);
nor U24697 (N_24697,N_23996,N_22101);
nand U24698 (N_24698,N_22413,N_22592);
nand U24699 (N_24699,N_22997,N_22579);
and U24700 (N_24700,N_23553,N_22919);
xnor U24701 (N_24701,N_22716,N_22043);
nand U24702 (N_24702,N_22198,N_23177);
xnor U24703 (N_24703,N_23195,N_23278);
xor U24704 (N_24704,N_22018,N_23670);
nor U24705 (N_24705,N_22648,N_22471);
xor U24706 (N_24706,N_23360,N_22688);
and U24707 (N_24707,N_23784,N_23546);
nor U24708 (N_24708,N_22297,N_23518);
nand U24709 (N_24709,N_23396,N_23355);
xor U24710 (N_24710,N_22819,N_22433);
nor U24711 (N_24711,N_22650,N_22501);
or U24712 (N_24712,N_23404,N_23867);
xor U24713 (N_24713,N_22711,N_23938);
or U24714 (N_24714,N_23002,N_23783);
or U24715 (N_24715,N_23156,N_22507);
nor U24716 (N_24716,N_22955,N_22816);
and U24717 (N_24717,N_22456,N_22589);
and U24718 (N_24718,N_23492,N_22674);
nand U24719 (N_24719,N_22721,N_22771);
and U24720 (N_24720,N_22588,N_23039);
xnor U24721 (N_24721,N_23244,N_23045);
and U24722 (N_24722,N_22288,N_22278);
xor U24723 (N_24723,N_23797,N_22920);
xor U24724 (N_24724,N_22371,N_23812);
nand U24725 (N_24725,N_23919,N_23698);
xnor U24726 (N_24726,N_22790,N_23676);
xnor U24727 (N_24727,N_22029,N_22117);
xnor U24728 (N_24728,N_23329,N_22896);
nor U24729 (N_24729,N_23215,N_22599);
nor U24730 (N_24730,N_22171,N_23968);
or U24731 (N_24731,N_23263,N_23738);
xnor U24732 (N_24732,N_23880,N_22930);
xor U24733 (N_24733,N_22440,N_23559);
nand U24734 (N_24734,N_22042,N_23219);
and U24735 (N_24735,N_23882,N_22879);
xor U24736 (N_24736,N_22237,N_23976);
nand U24737 (N_24737,N_23864,N_23716);
nor U24738 (N_24738,N_22742,N_23458);
nor U24739 (N_24739,N_23434,N_22693);
nand U24740 (N_24740,N_22391,N_23510);
nand U24741 (N_24741,N_22713,N_23910);
xnor U24742 (N_24742,N_22146,N_22837);
and U24743 (N_24743,N_23122,N_22808);
and U24744 (N_24744,N_23311,N_22148);
and U24745 (N_24745,N_23737,N_23438);
nor U24746 (N_24746,N_23550,N_23313);
nor U24747 (N_24747,N_22777,N_22859);
and U24748 (N_24748,N_22628,N_22007);
xor U24749 (N_24749,N_22318,N_23978);
or U24750 (N_24750,N_22634,N_22048);
xnor U24751 (N_24751,N_23640,N_23356);
xnor U24752 (N_24752,N_23076,N_22153);
and U24753 (N_24753,N_23763,N_22321);
or U24754 (N_24754,N_22936,N_23146);
xor U24755 (N_24755,N_23595,N_23308);
nor U24756 (N_24756,N_23223,N_23871);
nor U24757 (N_24757,N_22110,N_23118);
and U24758 (N_24758,N_23137,N_22383);
or U24759 (N_24759,N_23611,N_22629);
xor U24760 (N_24760,N_22710,N_23661);
nor U24761 (N_24761,N_22869,N_23287);
or U24762 (N_24762,N_23296,N_23618);
nor U24763 (N_24763,N_23178,N_22504);
nor U24764 (N_24764,N_22241,N_23925);
and U24765 (N_24765,N_22234,N_22000);
or U24766 (N_24766,N_22787,N_23230);
or U24767 (N_24767,N_22422,N_22460);
nor U24768 (N_24768,N_22956,N_23445);
or U24769 (N_24769,N_22916,N_23651);
or U24770 (N_24770,N_22760,N_22301);
nand U24771 (N_24771,N_22305,N_23427);
nand U24772 (N_24772,N_23092,N_23924);
nor U24773 (N_24773,N_22100,N_23312);
xnor U24774 (N_24774,N_22917,N_23431);
nor U24775 (N_24775,N_22342,N_22452);
or U24776 (N_24776,N_23724,N_22740);
and U24777 (N_24777,N_22283,N_23243);
and U24778 (N_24778,N_22017,N_22151);
and U24779 (N_24779,N_22943,N_22483);
and U24780 (N_24780,N_23609,N_23967);
nand U24781 (N_24781,N_22247,N_23253);
or U24782 (N_24782,N_22825,N_23692);
or U24783 (N_24783,N_22880,N_22586);
and U24784 (N_24784,N_22802,N_23028);
xor U24785 (N_24785,N_22206,N_22457);
xnor U24786 (N_24786,N_23386,N_22881);
xnor U24787 (N_24787,N_22612,N_22738);
nor U24788 (N_24788,N_22339,N_22664);
or U24789 (N_24789,N_23148,N_23063);
or U24790 (N_24790,N_23845,N_23801);
nand U24791 (N_24791,N_22179,N_22401);
xor U24792 (N_24792,N_22075,N_22059);
nor U24793 (N_24793,N_22060,N_23730);
and U24794 (N_24794,N_22388,N_23370);
nor U24795 (N_24795,N_23493,N_23439);
nor U24796 (N_24796,N_23726,N_22536);
and U24797 (N_24797,N_23874,N_22377);
nor U24798 (N_24798,N_22199,N_22846);
and U24799 (N_24799,N_23112,N_22273);
xor U24800 (N_24800,N_23577,N_23211);
and U24801 (N_24801,N_23364,N_23361);
and U24802 (N_24802,N_22901,N_22565);
nand U24803 (N_24803,N_22469,N_22115);
nor U24804 (N_24804,N_22999,N_23551);
and U24805 (N_24805,N_23939,N_23697);
nand U24806 (N_24806,N_23713,N_23035);
xor U24807 (N_24807,N_22888,N_23052);
and U24808 (N_24808,N_23682,N_22890);
or U24809 (N_24809,N_23677,N_23281);
xor U24810 (N_24810,N_22986,N_22240);
nand U24811 (N_24811,N_23774,N_23126);
and U24812 (N_24812,N_23592,N_22639);
nand U24813 (N_24813,N_23683,N_23983);
or U24814 (N_24814,N_22168,N_22548);
xor U24815 (N_24815,N_23905,N_22603);
or U24816 (N_24816,N_22578,N_23574);
nor U24817 (N_24817,N_23466,N_23017);
nand U24818 (N_24818,N_22731,N_22130);
nor U24819 (N_24819,N_22393,N_23524);
xnor U24820 (N_24820,N_23475,N_22724);
xor U24821 (N_24821,N_22434,N_23055);
xor U24822 (N_24822,N_23264,N_23209);
nand U24823 (N_24823,N_23930,N_22405);
xor U24824 (N_24824,N_23480,N_23733);
nor U24825 (N_24825,N_22652,N_23012);
nand U24826 (N_24826,N_22660,N_22085);
nor U24827 (N_24827,N_23406,N_23630);
nor U24828 (N_24828,N_22705,N_23750);
nor U24829 (N_24829,N_23805,N_22010);
and U24830 (N_24830,N_23452,N_23621);
xor U24831 (N_24831,N_23426,N_22436);
xor U24832 (N_24832,N_23854,N_23459);
and U24833 (N_24833,N_22411,N_23674);
and U24834 (N_24834,N_23573,N_22703);
nand U24835 (N_24835,N_22495,N_23955);
nor U24836 (N_24836,N_23689,N_23933);
and U24837 (N_24837,N_22344,N_22449);
nor U24838 (N_24838,N_23302,N_23138);
and U24839 (N_24839,N_23530,N_22509);
nor U24840 (N_24840,N_23456,N_22261);
or U24841 (N_24841,N_23314,N_22013);
nor U24842 (N_24842,N_23088,N_23071);
and U24843 (N_24843,N_23267,N_23131);
nand U24844 (N_24844,N_23669,N_22993);
nand U24845 (N_24845,N_23400,N_22605);
nor U24846 (N_24846,N_23816,N_23956);
nand U24847 (N_24847,N_23762,N_22221);
or U24848 (N_24848,N_23529,N_22733);
nor U24849 (N_24849,N_23470,N_22027);
or U24850 (N_24850,N_22512,N_23539);
nor U24851 (N_24851,N_23667,N_23772);
nor U24852 (N_24852,N_23600,N_22663);
and U24853 (N_24853,N_23690,N_23481);
nor U24854 (N_24854,N_23786,N_23419);
or U24855 (N_24855,N_23206,N_22264);
or U24856 (N_24856,N_22498,N_23391);
xnor U24857 (N_24857,N_22192,N_23926);
or U24858 (N_24858,N_22133,N_23610);
or U24859 (N_24859,N_23883,N_22331);
nor U24860 (N_24860,N_22286,N_22368);
xnor U24861 (N_24861,N_22893,N_22067);
nand U24862 (N_24862,N_23150,N_23149);
nand U24863 (N_24863,N_22038,N_23512);
xor U24864 (N_24864,N_23839,N_22942);
nand U24865 (N_24865,N_23660,N_23105);
nor U24866 (N_24866,N_23477,N_22142);
nand U24867 (N_24867,N_22821,N_22848);
or U24868 (N_24868,N_22312,N_23345);
or U24869 (N_24869,N_22613,N_22203);
or U24870 (N_24870,N_22758,N_22635);
or U24871 (N_24871,N_23714,N_23038);
and U24872 (N_24872,N_23950,N_23833);
or U24873 (N_24873,N_22518,N_22217);
nand U24874 (N_24874,N_22863,N_23194);
and U24875 (N_24875,N_22646,N_23659);
and U24876 (N_24876,N_22633,N_22748);
or U24877 (N_24877,N_23151,N_23310);
or U24878 (N_24878,N_23821,N_23245);
nand U24879 (N_24879,N_23860,N_23542);
nand U24880 (N_24880,N_23927,N_22420);
and U24881 (N_24881,N_22463,N_22669);
nand U24882 (N_24882,N_23217,N_23421);
or U24883 (N_24883,N_22493,N_23579);
nor U24884 (N_24884,N_22989,N_23089);
nand U24885 (N_24885,N_22970,N_23371);
nand U24886 (N_24886,N_23836,N_23887);
or U24887 (N_24887,N_22892,N_22165);
nor U24888 (N_24888,N_23536,N_23999);
nand U24889 (N_24889,N_22200,N_23321);
nand U24890 (N_24890,N_23349,N_23085);
or U24891 (N_24891,N_23561,N_22624);
or U24892 (N_24892,N_22083,N_22723);
xnor U24893 (N_24893,N_23330,N_22058);
nand U24894 (N_24894,N_23562,N_23372);
and U24895 (N_24895,N_22689,N_23095);
or U24896 (N_24896,N_22376,N_23819);
xnor U24897 (N_24897,N_23093,N_22020);
and U24898 (N_24898,N_23817,N_23001);
xor U24899 (N_24899,N_23829,N_23850);
or U24900 (N_24900,N_22431,N_23838);
nor U24901 (N_24901,N_22983,N_23893);
or U24902 (N_24902,N_22030,N_23725);
xor U24903 (N_24903,N_22233,N_23572);
xnor U24904 (N_24904,N_23455,N_23800);
and U24905 (N_24905,N_23863,N_22614);
or U24906 (N_24906,N_23822,N_23581);
nand U24907 (N_24907,N_23270,N_23744);
and U24908 (N_24908,N_22108,N_22598);
and U24909 (N_24909,N_23736,N_23937);
nand U24910 (N_24910,N_23143,N_23198);
nor U24911 (N_24911,N_22396,N_23798);
and U24912 (N_24912,N_23203,N_22224);
nand U24913 (N_24913,N_22523,N_23958);
or U24914 (N_24914,N_23168,N_22560);
nor U24915 (N_24915,N_23633,N_22304);
and U24916 (N_24916,N_23517,N_22089);
nand U24917 (N_24917,N_23987,N_22348);
nand U24918 (N_24918,N_23773,N_22632);
xnor U24919 (N_24919,N_23262,N_22572);
or U24920 (N_24920,N_23132,N_22005);
xor U24921 (N_24921,N_23488,N_22266);
xnor U24922 (N_24922,N_23121,N_22720);
and U24923 (N_24923,N_23626,N_23183);
or U24924 (N_24924,N_23210,N_22093);
and U24925 (N_24925,N_23703,N_23200);
or U24926 (N_24926,N_22729,N_23769);
nor U24927 (N_24927,N_23242,N_22801);
nor U24928 (N_24928,N_23583,N_23175);
xor U24929 (N_24929,N_22939,N_22630);
nor U24930 (N_24930,N_23959,N_22269);
or U24931 (N_24931,N_22952,N_22545);
or U24932 (N_24932,N_23929,N_22737);
nor U24933 (N_24933,N_23043,N_23861);
or U24934 (N_24934,N_23525,N_23755);
or U24935 (N_24935,N_22596,N_22150);
nor U24936 (N_24936,N_22617,N_23825);
nor U24937 (N_24937,N_22128,N_22324);
nor U24938 (N_24938,N_22817,N_22948);
and U24939 (N_24939,N_23841,N_22566);
and U24940 (N_24940,N_22428,N_23465);
nand U24941 (N_24941,N_22211,N_22799);
or U24942 (N_24942,N_23707,N_23647);
xnor U24943 (N_24943,N_23004,N_23064);
and U24944 (N_24944,N_22230,N_22670);
nor U24945 (N_24945,N_23789,N_23852);
and U24946 (N_24946,N_22263,N_23872);
xor U24947 (N_24947,N_22145,N_22147);
or U24948 (N_24948,N_22012,N_22769);
nor U24949 (N_24949,N_22122,N_22189);
nor U24950 (N_24950,N_22656,N_22409);
or U24951 (N_24951,N_22686,N_23820);
nor U24952 (N_24952,N_22270,N_22953);
nand U24953 (N_24953,N_23662,N_22762);
nor U24954 (N_24954,N_23205,N_23594);
and U24955 (N_24955,N_22570,N_22488);
and U24956 (N_24956,N_23538,N_23000);
nand U24957 (N_24957,N_22272,N_23285);
nor U24958 (N_24958,N_23221,N_23563);
or U24959 (N_24959,N_23960,N_22675);
and U24960 (N_24960,N_22227,N_23006);
and U24961 (N_24961,N_23109,N_22915);
xnor U24962 (N_24962,N_23265,N_22249);
nor U24963 (N_24963,N_23888,N_23068);
nor U24964 (N_24964,N_23742,N_22477);
xor U24965 (N_24965,N_22071,N_23324);
or U24966 (N_24966,N_22754,N_22701);
or U24967 (N_24967,N_22176,N_22424);
and U24968 (N_24968,N_22868,N_22995);
nor U24969 (N_24969,N_22949,N_22521);
and U24970 (N_24970,N_23393,N_22358);
and U24971 (N_24971,N_23288,N_22056);
or U24972 (N_24972,N_23895,N_23918);
xor U24973 (N_24973,N_22141,N_22223);
and U24974 (N_24974,N_22517,N_22416);
or U24975 (N_24975,N_23693,N_22285);
and U24976 (N_24976,N_23969,N_23932);
nand U24977 (N_24977,N_22839,N_23501);
and U24978 (N_24978,N_23057,N_23103);
xor U24979 (N_24979,N_23509,N_23652);
nor U24980 (N_24980,N_22046,N_22090);
nand U24981 (N_24981,N_22658,N_22631);
xor U24982 (N_24982,N_22271,N_23760);
xnor U24983 (N_24983,N_22643,N_23803);
or U24984 (N_24984,N_23560,N_22002);
nand U24985 (N_24985,N_22006,N_22985);
xnor U24986 (N_24986,N_22749,N_22127);
and U24987 (N_24987,N_22462,N_23729);
nor U24988 (N_24988,N_22251,N_23069);
nor U24989 (N_24989,N_23145,N_22615);
nand U24990 (N_24990,N_23569,N_22616);
or U24991 (N_24991,N_22681,N_22138);
and U24992 (N_24992,N_23907,N_23641);
or U24993 (N_24993,N_22185,N_22465);
or U24994 (N_24994,N_22538,N_23173);
nor U24995 (N_24995,N_23942,N_23522);
and U24996 (N_24996,N_23654,N_23584);
or U24997 (N_24997,N_22649,N_22746);
nand U24998 (N_24998,N_23954,N_22852);
nand U24999 (N_24999,N_23753,N_23568);
xnor U25000 (N_25000,N_22843,N_23246);
nand U25001 (N_25001,N_23220,N_22023);
or U25002 (N_25002,N_23487,N_23423);
xnor U25003 (N_25003,N_23790,N_22744);
nand U25004 (N_25004,N_22994,N_22711);
nor U25005 (N_25005,N_22216,N_23113);
nand U25006 (N_25006,N_22163,N_23735);
nand U25007 (N_25007,N_23706,N_22135);
nand U25008 (N_25008,N_23186,N_22577);
nand U25009 (N_25009,N_23455,N_23582);
or U25010 (N_25010,N_22323,N_22841);
xor U25011 (N_25011,N_23712,N_23513);
xnor U25012 (N_25012,N_22790,N_23321);
and U25013 (N_25013,N_23226,N_23308);
nand U25014 (N_25014,N_23446,N_22074);
or U25015 (N_25015,N_22953,N_22302);
or U25016 (N_25016,N_22003,N_22326);
nor U25017 (N_25017,N_23005,N_22408);
xnor U25018 (N_25018,N_23997,N_22530);
nor U25019 (N_25019,N_23141,N_22332);
nor U25020 (N_25020,N_22643,N_23368);
and U25021 (N_25021,N_22096,N_23075);
xor U25022 (N_25022,N_22213,N_23852);
nor U25023 (N_25023,N_22847,N_23529);
xor U25024 (N_25024,N_23417,N_22713);
or U25025 (N_25025,N_23005,N_23597);
xnor U25026 (N_25026,N_23375,N_22933);
and U25027 (N_25027,N_23700,N_22400);
nor U25028 (N_25028,N_22781,N_23594);
xnor U25029 (N_25029,N_22661,N_22081);
and U25030 (N_25030,N_22113,N_23120);
or U25031 (N_25031,N_22872,N_23376);
nor U25032 (N_25032,N_23763,N_22275);
and U25033 (N_25033,N_23171,N_22889);
nand U25034 (N_25034,N_22073,N_22333);
or U25035 (N_25035,N_22900,N_23244);
nor U25036 (N_25036,N_22432,N_22825);
and U25037 (N_25037,N_23764,N_23420);
and U25038 (N_25038,N_23394,N_23005);
xnor U25039 (N_25039,N_23501,N_23592);
nand U25040 (N_25040,N_22201,N_22695);
and U25041 (N_25041,N_22381,N_23464);
xor U25042 (N_25042,N_22801,N_23176);
or U25043 (N_25043,N_23572,N_22220);
and U25044 (N_25044,N_22635,N_22023);
nor U25045 (N_25045,N_22652,N_22783);
nand U25046 (N_25046,N_23165,N_23711);
and U25047 (N_25047,N_23117,N_22689);
xnor U25048 (N_25048,N_23243,N_22885);
and U25049 (N_25049,N_22958,N_23091);
or U25050 (N_25050,N_22563,N_23364);
and U25051 (N_25051,N_22462,N_22723);
nand U25052 (N_25052,N_23757,N_22187);
or U25053 (N_25053,N_22011,N_22813);
nor U25054 (N_25054,N_22522,N_22166);
and U25055 (N_25055,N_22055,N_23143);
nand U25056 (N_25056,N_23597,N_23018);
nand U25057 (N_25057,N_23814,N_23158);
nor U25058 (N_25058,N_22502,N_22142);
nor U25059 (N_25059,N_23806,N_23427);
or U25060 (N_25060,N_22983,N_23005);
xor U25061 (N_25061,N_22468,N_23460);
nand U25062 (N_25062,N_23150,N_22431);
or U25063 (N_25063,N_23392,N_23082);
or U25064 (N_25064,N_22000,N_23701);
nor U25065 (N_25065,N_22562,N_22679);
or U25066 (N_25066,N_22585,N_23534);
xnor U25067 (N_25067,N_22103,N_22887);
or U25068 (N_25068,N_22732,N_23970);
xor U25069 (N_25069,N_23550,N_22826);
nand U25070 (N_25070,N_22093,N_22652);
nor U25071 (N_25071,N_23745,N_22131);
xor U25072 (N_25072,N_22103,N_23723);
or U25073 (N_25073,N_22336,N_22608);
nand U25074 (N_25074,N_23906,N_22055);
xnor U25075 (N_25075,N_23327,N_22433);
nor U25076 (N_25076,N_23408,N_23971);
nor U25077 (N_25077,N_22881,N_23665);
xnor U25078 (N_25078,N_22352,N_22789);
and U25079 (N_25079,N_22110,N_23960);
nand U25080 (N_25080,N_22837,N_23628);
nor U25081 (N_25081,N_23299,N_22972);
nand U25082 (N_25082,N_23155,N_22955);
nand U25083 (N_25083,N_23480,N_22763);
xor U25084 (N_25084,N_23232,N_23581);
and U25085 (N_25085,N_22711,N_23990);
and U25086 (N_25086,N_22666,N_22664);
nor U25087 (N_25087,N_23059,N_22853);
and U25088 (N_25088,N_22089,N_22413);
and U25089 (N_25089,N_23969,N_23933);
and U25090 (N_25090,N_23092,N_22124);
nand U25091 (N_25091,N_23890,N_23204);
nor U25092 (N_25092,N_22582,N_22883);
nor U25093 (N_25093,N_23448,N_22079);
or U25094 (N_25094,N_22779,N_23209);
and U25095 (N_25095,N_22626,N_22981);
nand U25096 (N_25096,N_23621,N_23345);
and U25097 (N_25097,N_22605,N_22820);
xnor U25098 (N_25098,N_22006,N_22777);
or U25099 (N_25099,N_23657,N_23766);
xor U25100 (N_25100,N_22063,N_22583);
xor U25101 (N_25101,N_23594,N_23373);
xnor U25102 (N_25102,N_23966,N_23000);
xnor U25103 (N_25103,N_22389,N_22561);
nand U25104 (N_25104,N_22996,N_22270);
xor U25105 (N_25105,N_23667,N_23735);
and U25106 (N_25106,N_23706,N_23408);
and U25107 (N_25107,N_22215,N_23576);
nand U25108 (N_25108,N_22429,N_23048);
nor U25109 (N_25109,N_23514,N_22404);
nor U25110 (N_25110,N_22514,N_22141);
or U25111 (N_25111,N_23977,N_22707);
nor U25112 (N_25112,N_23832,N_22638);
nand U25113 (N_25113,N_23353,N_22470);
nor U25114 (N_25114,N_23729,N_23142);
nor U25115 (N_25115,N_23741,N_23062);
or U25116 (N_25116,N_23150,N_23203);
xor U25117 (N_25117,N_22851,N_22869);
and U25118 (N_25118,N_23428,N_22246);
nor U25119 (N_25119,N_23238,N_23858);
nor U25120 (N_25120,N_22371,N_23192);
nand U25121 (N_25121,N_23177,N_23400);
or U25122 (N_25122,N_22528,N_22702);
and U25123 (N_25123,N_23876,N_23412);
nand U25124 (N_25124,N_22007,N_23333);
and U25125 (N_25125,N_23323,N_22672);
nand U25126 (N_25126,N_22796,N_22425);
or U25127 (N_25127,N_22965,N_22008);
and U25128 (N_25128,N_23864,N_23048);
or U25129 (N_25129,N_22970,N_22766);
xnor U25130 (N_25130,N_23569,N_22872);
and U25131 (N_25131,N_22970,N_23419);
xnor U25132 (N_25132,N_22114,N_22059);
xnor U25133 (N_25133,N_23546,N_22999);
nand U25134 (N_25134,N_22848,N_23303);
nor U25135 (N_25135,N_23880,N_22545);
nor U25136 (N_25136,N_23616,N_23403);
and U25137 (N_25137,N_22528,N_22774);
and U25138 (N_25138,N_23547,N_23474);
xnor U25139 (N_25139,N_22009,N_23607);
nand U25140 (N_25140,N_23949,N_22602);
or U25141 (N_25141,N_22487,N_23929);
nor U25142 (N_25142,N_22009,N_22154);
xnor U25143 (N_25143,N_23942,N_23247);
nand U25144 (N_25144,N_23851,N_23969);
nand U25145 (N_25145,N_23752,N_23995);
or U25146 (N_25146,N_23467,N_23866);
nor U25147 (N_25147,N_22473,N_22666);
or U25148 (N_25148,N_23693,N_23446);
and U25149 (N_25149,N_22627,N_23214);
nand U25150 (N_25150,N_22954,N_22090);
and U25151 (N_25151,N_22755,N_22279);
and U25152 (N_25152,N_23003,N_22367);
and U25153 (N_25153,N_22446,N_22118);
nand U25154 (N_25154,N_23722,N_22874);
xnor U25155 (N_25155,N_23359,N_23262);
nor U25156 (N_25156,N_23797,N_22286);
or U25157 (N_25157,N_23963,N_23185);
nand U25158 (N_25158,N_23841,N_22726);
and U25159 (N_25159,N_22542,N_22954);
nand U25160 (N_25160,N_23196,N_23125);
xnor U25161 (N_25161,N_23064,N_22885);
nor U25162 (N_25162,N_23501,N_23815);
nor U25163 (N_25163,N_23194,N_23462);
and U25164 (N_25164,N_22052,N_23663);
nor U25165 (N_25165,N_22235,N_23660);
and U25166 (N_25166,N_22620,N_23107);
nor U25167 (N_25167,N_22900,N_23180);
or U25168 (N_25168,N_23207,N_23405);
nor U25169 (N_25169,N_22451,N_22367);
nand U25170 (N_25170,N_22491,N_23604);
and U25171 (N_25171,N_22495,N_22577);
or U25172 (N_25172,N_22305,N_23692);
xnor U25173 (N_25173,N_22507,N_22881);
and U25174 (N_25174,N_22866,N_22176);
or U25175 (N_25175,N_23090,N_22788);
and U25176 (N_25176,N_23545,N_23804);
and U25177 (N_25177,N_23313,N_22682);
nand U25178 (N_25178,N_23463,N_22842);
nand U25179 (N_25179,N_22651,N_23163);
nand U25180 (N_25180,N_23785,N_23736);
and U25181 (N_25181,N_23621,N_22755);
and U25182 (N_25182,N_23990,N_22844);
and U25183 (N_25183,N_22120,N_22214);
nor U25184 (N_25184,N_22273,N_23359);
xor U25185 (N_25185,N_23932,N_22935);
or U25186 (N_25186,N_22484,N_22241);
nor U25187 (N_25187,N_22228,N_23532);
xor U25188 (N_25188,N_22874,N_22638);
xnor U25189 (N_25189,N_22492,N_23510);
or U25190 (N_25190,N_22619,N_23561);
nor U25191 (N_25191,N_22348,N_22105);
nand U25192 (N_25192,N_23206,N_23587);
and U25193 (N_25193,N_22044,N_23192);
nor U25194 (N_25194,N_23158,N_22829);
and U25195 (N_25195,N_22331,N_22378);
nand U25196 (N_25196,N_22797,N_22186);
and U25197 (N_25197,N_22393,N_22711);
xnor U25198 (N_25198,N_23376,N_22987);
xnor U25199 (N_25199,N_23256,N_22636);
nand U25200 (N_25200,N_22054,N_23956);
or U25201 (N_25201,N_22682,N_23410);
and U25202 (N_25202,N_23519,N_23613);
nand U25203 (N_25203,N_23263,N_23699);
nor U25204 (N_25204,N_23357,N_23612);
xor U25205 (N_25205,N_23848,N_23500);
nand U25206 (N_25206,N_23558,N_23514);
or U25207 (N_25207,N_23281,N_22471);
nor U25208 (N_25208,N_23414,N_23759);
nor U25209 (N_25209,N_23713,N_22777);
xnor U25210 (N_25210,N_22892,N_22925);
nand U25211 (N_25211,N_22494,N_22118);
or U25212 (N_25212,N_22021,N_22497);
nor U25213 (N_25213,N_23303,N_23835);
nand U25214 (N_25214,N_22450,N_23063);
or U25215 (N_25215,N_22302,N_22098);
nor U25216 (N_25216,N_22538,N_23040);
and U25217 (N_25217,N_22543,N_23662);
nand U25218 (N_25218,N_22928,N_22157);
or U25219 (N_25219,N_23130,N_23056);
xor U25220 (N_25220,N_23322,N_22694);
xor U25221 (N_25221,N_22708,N_22572);
nor U25222 (N_25222,N_23051,N_22970);
and U25223 (N_25223,N_23958,N_22324);
nand U25224 (N_25224,N_22182,N_23661);
xnor U25225 (N_25225,N_22656,N_23817);
or U25226 (N_25226,N_22993,N_22126);
xor U25227 (N_25227,N_23073,N_22879);
nand U25228 (N_25228,N_23541,N_22375);
nor U25229 (N_25229,N_22121,N_23778);
nand U25230 (N_25230,N_22064,N_22108);
nor U25231 (N_25231,N_22003,N_23158);
or U25232 (N_25232,N_22959,N_23699);
and U25233 (N_25233,N_22811,N_22591);
nand U25234 (N_25234,N_23303,N_22897);
xor U25235 (N_25235,N_22718,N_23454);
xnor U25236 (N_25236,N_22581,N_22981);
xnor U25237 (N_25237,N_23192,N_22306);
and U25238 (N_25238,N_22421,N_22231);
xor U25239 (N_25239,N_22861,N_22077);
nor U25240 (N_25240,N_22799,N_23797);
and U25241 (N_25241,N_23264,N_22428);
or U25242 (N_25242,N_23703,N_23652);
nand U25243 (N_25243,N_22617,N_22602);
or U25244 (N_25244,N_23703,N_23995);
nand U25245 (N_25245,N_23170,N_22085);
nand U25246 (N_25246,N_22575,N_23512);
nor U25247 (N_25247,N_22697,N_23592);
xor U25248 (N_25248,N_23663,N_23875);
nor U25249 (N_25249,N_23489,N_22740);
nand U25250 (N_25250,N_23103,N_22732);
xor U25251 (N_25251,N_23916,N_23199);
or U25252 (N_25252,N_23640,N_22675);
and U25253 (N_25253,N_23929,N_23164);
xor U25254 (N_25254,N_22040,N_23848);
nand U25255 (N_25255,N_22489,N_22769);
xnor U25256 (N_25256,N_22179,N_23242);
xor U25257 (N_25257,N_23918,N_22367);
xnor U25258 (N_25258,N_22642,N_22018);
nor U25259 (N_25259,N_22517,N_23791);
nor U25260 (N_25260,N_22798,N_22717);
nor U25261 (N_25261,N_23407,N_22594);
or U25262 (N_25262,N_23333,N_23789);
xor U25263 (N_25263,N_22776,N_23850);
nor U25264 (N_25264,N_22153,N_23272);
and U25265 (N_25265,N_23705,N_23714);
and U25266 (N_25266,N_22140,N_23393);
nor U25267 (N_25267,N_22050,N_23752);
or U25268 (N_25268,N_22511,N_22603);
nand U25269 (N_25269,N_23821,N_22500);
xnor U25270 (N_25270,N_22686,N_23518);
or U25271 (N_25271,N_23152,N_23715);
xor U25272 (N_25272,N_22397,N_23829);
xnor U25273 (N_25273,N_22773,N_23955);
or U25274 (N_25274,N_22850,N_23725);
xnor U25275 (N_25275,N_22475,N_23023);
or U25276 (N_25276,N_23968,N_23964);
and U25277 (N_25277,N_23094,N_22258);
or U25278 (N_25278,N_23998,N_23586);
xnor U25279 (N_25279,N_23419,N_23791);
nand U25280 (N_25280,N_22878,N_23154);
or U25281 (N_25281,N_22925,N_22960);
xor U25282 (N_25282,N_23955,N_22606);
xor U25283 (N_25283,N_23991,N_22953);
nor U25284 (N_25284,N_22867,N_23267);
nor U25285 (N_25285,N_22687,N_23912);
xor U25286 (N_25286,N_22730,N_22266);
or U25287 (N_25287,N_22290,N_22141);
and U25288 (N_25288,N_22397,N_22470);
nand U25289 (N_25289,N_23318,N_23988);
nand U25290 (N_25290,N_23272,N_23383);
nor U25291 (N_25291,N_22350,N_23181);
and U25292 (N_25292,N_22777,N_23908);
xnor U25293 (N_25293,N_22806,N_22691);
and U25294 (N_25294,N_22800,N_23357);
and U25295 (N_25295,N_23896,N_23431);
xor U25296 (N_25296,N_22944,N_22464);
and U25297 (N_25297,N_23802,N_22677);
nor U25298 (N_25298,N_23545,N_23454);
nor U25299 (N_25299,N_23256,N_22200);
nand U25300 (N_25300,N_22535,N_22906);
xnor U25301 (N_25301,N_23537,N_22935);
nand U25302 (N_25302,N_22312,N_23109);
nand U25303 (N_25303,N_23692,N_22523);
or U25304 (N_25304,N_23753,N_22747);
or U25305 (N_25305,N_22735,N_23235);
nand U25306 (N_25306,N_22398,N_22993);
nand U25307 (N_25307,N_23930,N_22606);
nor U25308 (N_25308,N_22132,N_23667);
xnor U25309 (N_25309,N_23027,N_22663);
xor U25310 (N_25310,N_23635,N_22078);
nor U25311 (N_25311,N_22662,N_23270);
nand U25312 (N_25312,N_22392,N_22515);
xnor U25313 (N_25313,N_23242,N_23207);
nand U25314 (N_25314,N_22474,N_22624);
nor U25315 (N_25315,N_22988,N_22070);
nor U25316 (N_25316,N_23941,N_22669);
or U25317 (N_25317,N_22875,N_23548);
nor U25318 (N_25318,N_23990,N_23004);
and U25319 (N_25319,N_23918,N_22768);
and U25320 (N_25320,N_23941,N_23649);
nor U25321 (N_25321,N_22262,N_22680);
nor U25322 (N_25322,N_23288,N_23748);
and U25323 (N_25323,N_22510,N_22467);
nor U25324 (N_25324,N_23328,N_23718);
xor U25325 (N_25325,N_22071,N_22414);
and U25326 (N_25326,N_22475,N_22125);
nand U25327 (N_25327,N_22920,N_23725);
or U25328 (N_25328,N_22064,N_22637);
or U25329 (N_25329,N_23599,N_22047);
and U25330 (N_25330,N_22132,N_23531);
xor U25331 (N_25331,N_22478,N_23382);
xor U25332 (N_25332,N_22177,N_22086);
xnor U25333 (N_25333,N_23054,N_22147);
nand U25334 (N_25334,N_23166,N_22256);
xor U25335 (N_25335,N_23938,N_23360);
or U25336 (N_25336,N_23865,N_23105);
or U25337 (N_25337,N_22039,N_23543);
and U25338 (N_25338,N_23026,N_22456);
or U25339 (N_25339,N_23296,N_22123);
nor U25340 (N_25340,N_22353,N_22210);
xor U25341 (N_25341,N_23669,N_23583);
xnor U25342 (N_25342,N_22768,N_22879);
nand U25343 (N_25343,N_23350,N_23394);
and U25344 (N_25344,N_23457,N_23851);
and U25345 (N_25345,N_22051,N_22173);
xnor U25346 (N_25346,N_23690,N_22945);
xor U25347 (N_25347,N_23799,N_23783);
nand U25348 (N_25348,N_22532,N_23802);
and U25349 (N_25349,N_23145,N_23753);
and U25350 (N_25350,N_23935,N_23814);
and U25351 (N_25351,N_23719,N_22226);
and U25352 (N_25352,N_22385,N_23267);
nand U25353 (N_25353,N_23638,N_22682);
or U25354 (N_25354,N_22361,N_22463);
xnor U25355 (N_25355,N_22124,N_23702);
xnor U25356 (N_25356,N_22147,N_22587);
or U25357 (N_25357,N_23276,N_22710);
xnor U25358 (N_25358,N_23679,N_23771);
or U25359 (N_25359,N_23683,N_22025);
or U25360 (N_25360,N_22634,N_23278);
nand U25361 (N_25361,N_22116,N_22493);
nor U25362 (N_25362,N_23952,N_23473);
nor U25363 (N_25363,N_22108,N_23956);
and U25364 (N_25364,N_22953,N_23011);
or U25365 (N_25365,N_22422,N_22055);
and U25366 (N_25366,N_22184,N_22687);
nand U25367 (N_25367,N_22914,N_22986);
or U25368 (N_25368,N_23278,N_22811);
xor U25369 (N_25369,N_22649,N_22523);
nand U25370 (N_25370,N_23314,N_22510);
or U25371 (N_25371,N_22793,N_22260);
or U25372 (N_25372,N_23080,N_22320);
nand U25373 (N_25373,N_22077,N_22806);
or U25374 (N_25374,N_22859,N_23094);
nor U25375 (N_25375,N_23922,N_22066);
nor U25376 (N_25376,N_22247,N_22392);
or U25377 (N_25377,N_23022,N_22194);
or U25378 (N_25378,N_23736,N_23149);
nand U25379 (N_25379,N_23788,N_22949);
and U25380 (N_25380,N_23063,N_22801);
or U25381 (N_25381,N_23336,N_23391);
or U25382 (N_25382,N_22004,N_23920);
and U25383 (N_25383,N_23155,N_23447);
or U25384 (N_25384,N_23593,N_23772);
xor U25385 (N_25385,N_22312,N_22406);
and U25386 (N_25386,N_23414,N_22870);
or U25387 (N_25387,N_22061,N_23809);
or U25388 (N_25388,N_22918,N_23731);
or U25389 (N_25389,N_23315,N_23254);
or U25390 (N_25390,N_23883,N_22677);
nand U25391 (N_25391,N_22570,N_22323);
or U25392 (N_25392,N_23048,N_23653);
and U25393 (N_25393,N_22227,N_22465);
or U25394 (N_25394,N_22206,N_23624);
and U25395 (N_25395,N_23715,N_22157);
or U25396 (N_25396,N_22274,N_22470);
and U25397 (N_25397,N_23354,N_22949);
and U25398 (N_25398,N_23754,N_23858);
nand U25399 (N_25399,N_22137,N_22305);
or U25400 (N_25400,N_22567,N_22428);
xor U25401 (N_25401,N_23431,N_23169);
xor U25402 (N_25402,N_23124,N_22182);
nand U25403 (N_25403,N_23062,N_22144);
nand U25404 (N_25404,N_22875,N_23359);
nor U25405 (N_25405,N_23418,N_23284);
and U25406 (N_25406,N_22158,N_22171);
nor U25407 (N_25407,N_22625,N_22410);
and U25408 (N_25408,N_22836,N_23892);
nor U25409 (N_25409,N_23776,N_23594);
nand U25410 (N_25410,N_22035,N_22850);
or U25411 (N_25411,N_22333,N_23306);
xor U25412 (N_25412,N_23895,N_23283);
nand U25413 (N_25413,N_22361,N_22644);
nand U25414 (N_25414,N_22912,N_22692);
and U25415 (N_25415,N_22904,N_22340);
and U25416 (N_25416,N_23773,N_22809);
or U25417 (N_25417,N_22464,N_23184);
and U25418 (N_25418,N_23862,N_22473);
xnor U25419 (N_25419,N_23068,N_22989);
or U25420 (N_25420,N_23060,N_22287);
nand U25421 (N_25421,N_23166,N_23761);
nor U25422 (N_25422,N_22962,N_23382);
xnor U25423 (N_25423,N_22201,N_23239);
xor U25424 (N_25424,N_22976,N_23060);
nor U25425 (N_25425,N_23527,N_23892);
or U25426 (N_25426,N_22505,N_23855);
nor U25427 (N_25427,N_23250,N_22847);
xnor U25428 (N_25428,N_23434,N_23156);
and U25429 (N_25429,N_23797,N_23986);
nand U25430 (N_25430,N_22456,N_22491);
and U25431 (N_25431,N_22640,N_22231);
xnor U25432 (N_25432,N_23977,N_23145);
nor U25433 (N_25433,N_23620,N_22786);
nand U25434 (N_25434,N_23571,N_22601);
nor U25435 (N_25435,N_22349,N_23405);
nand U25436 (N_25436,N_23557,N_23842);
and U25437 (N_25437,N_23618,N_22548);
xor U25438 (N_25438,N_22073,N_23513);
or U25439 (N_25439,N_23549,N_22229);
or U25440 (N_25440,N_23874,N_22893);
nor U25441 (N_25441,N_22917,N_23456);
and U25442 (N_25442,N_23970,N_23528);
nand U25443 (N_25443,N_22209,N_22248);
and U25444 (N_25444,N_22786,N_22353);
nor U25445 (N_25445,N_23915,N_23112);
nor U25446 (N_25446,N_22341,N_23771);
xnor U25447 (N_25447,N_23900,N_23797);
xor U25448 (N_25448,N_23877,N_23968);
xor U25449 (N_25449,N_22219,N_22708);
nor U25450 (N_25450,N_22314,N_23536);
or U25451 (N_25451,N_22014,N_22303);
xor U25452 (N_25452,N_22901,N_23306);
and U25453 (N_25453,N_23135,N_23467);
nand U25454 (N_25454,N_23191,N_22525);
xnor U25455 (N_25455,N_22588,N_23958);
nor U25456 (N_25456,N_23685,N_22396);
nor U25457 (N_25457,N_23160,N_23037);
and U25458 (N_25458,N_22931,N_22160);
xnor U25459 (N_25459,N_23527,N_22543);
nor U25460 (N_25460,N_23337,N_22552);
nor U25461 (N_25461,N_22841,N_22143);
nand U25462 (N_25462,N_23117,N_22299);
nor U25463 (N_25463,N_22791,N_22094);
nand U25464 (N_25464,N_23746,N_22716);
nand U25465 (N_25465,N_23121,N_22787);
or U25466 (N_25466,N_22433,N_22336);
or U25467 (N_25467,N_22673,N_22334);
xnor U25468 (N_25468,N_23520,N_22621);
xnor U25469 (N_25469,N_23140,N_22665);
nor U25470 (N_25470,N_22016,N_23807);
xnor U25471 (N_25471,N_23901,N_22357);
and U25472 (N_25472,N_22238,N_23363);
or U25473 (N_25473,N_22196,N_23445);
or U25474 (N_25474,N_23841,N_23629);
and U25475 (N_25475,N_23969,N_22970);
nor U25476 (N_25476,N_22260,N_23147);
xor U25477 (N_25477,N_23511,N_23954);
xnor U25478 (N_25478,N_22154,N_23767);
nor U25479 (N_25479,N_22188,N_23212);
xor U25480 (N_25480,N_23936,N_22370);
xor U25481 (N_25481,N_23968,N_22671);
nor U25482 (N_25482,N_23394,N_23432);
or U25483 (N_25483,N_23398,N_22379);
or U25484 (N_25484,N_23859,N_22384);
xor U25485 (N_25485,N_22206,N_23735);
and U25486 (N_25486,N_22229,N_22095);
nand U25487 (N_25487,N_22541,N_23800);
nand U25488 (N_25488,N_23104,N_22059);
and U25489 (N_25489,N_22012,N_22270);
nor U25490 (N_25490,N_22452,N_23896);
xor U25491 (N_25491,N_23827,N_23249);
and U25492 (N_25492,N_23613,N_23188);
or U25493 (N_25493,N_22755,N_22250);
nand U25494 (N_25494,N_23340,N_22519);
xnor U25495 (N_25495,N_22027,N_22192);
xnor U25496 (N_25496,N_22303,N_22203);
nand U25497 (N_25497,N_22461,N_23272);
or U25498 (N_25498,N_23494,N_22206);
or U25499 (N_25499,N_22315,N_23865);
nand U25500 (N_25500,N_23197,N_23451);
and U25501 (N_25501,N_23479,N_23775);
and U25502 (N_25502,N_22110,N_23884);
nand U25503 (N_25503,N_22051,N_22202);
or U25504 (N_25504,N_23633,N_22069);
nand U25505 (N_25505,N_23238,N_22629);
nand U25506 (N_25506,N_22799,N_22263);
and U25507 (N_25507,N_23118,N_22883);
xor U25508 (N_25508,N_23599,N_22264);
or U25509 (N_25509,N_22222,N_23940);
nand U25510 (N_25510,N_22994,N_23857);
xnor U25511 (N_25511,N_23257,N_22816);
xor U25512 (N_25512,N_23998,N_22628);
and U25513 (N_25513,N_23393,N_22426);
and U25514 (N_25514,N_22923,N_23356);
or U25515 (N_25515,N_23389,N_23292);
nand U25516 (N_25516,N_22758,N_23894);
or U25517 (N_25517,N_23990,N_23729);
xnor U25518 (N_25518,N_22910,N_23119);
and U25519 (N_25519,N_23866,N_22848);
or U25520 (N_25520,N_23977,N_22197);
and U25521 (N_25521,N_22908,N_22224);
nand U25522 (N_25522,N_23552,N_23931);
nand U25523 (N_25523,N_23680,N_22262);
or U25524 (N_25524,N_23645,N_23827);
or U25525 (N_25525,N_22696,N_23424);
nand U25526 (N_25526,N_22194,N_23806);
or U25527 (N_25527,N_23514,N_22954);
xor U25528 (N_25528,N_23787,N_22491);
or U25529 (N_25529,N_22302,N_23674);
or U25530 (N_25530,N_23323,N_22292);
nor U25531 (N_25531,N_23240,N_22247);
and U25532 (N_25532,N_23827,N_22919);
nand U25533 (N_25533,N_22903,N_23032);
nand U25534 (N_25534,N_23060,N_22794);
xnor U25535 (N_25535,N_23028,N_23784);
or U25536 (N_25536,N_23690,N_23474);
xor U25537 (N_25537,N_22313,N_23547);
nor U25538 (N_25538,N_22510,N_23288);
nor U25539 (N_25539,N_22844,N_22673);
xnor U25540 (N_25540,N_23802,N_22995);
and U25541 (N_25541,N_22458,N_23768);
and U25542 (N_25542,N_22626,N_23499);
or U25543 (N_25543,N_23875,N_23773);
and U25544 (N_25544,N_23010,N_22795);
nor U25545 (N_25545,N_22650,N_23477);
nor U25546 (N_25546,N_23202,N_22403);
nor U25547 (N_25547,N_23016,N_23412);
nand U25548 (N_25548,N_22173,N_22254);
and U25549 (N_25549,N_23562,N_23211);
nor U25550 (N_25550,N_23903,N_23932);
and U25551 (N_25551,N_22820,N_23606);
or U25552 (N_25552,N_22108,N_23981);
nor U25553 (N_25553,N_23673,N_23644);
or U25554 (N_25554,N_23764,N_23179);
and U25555 (N_25555,N_22540,N_22761);
xor U25556 (N_25556,N_23002,N_22279);
or U25557 (N_25557,N_22251,N_23192);
nand U25558 (N_25558,N_23989,N_22292);
or U25559 (N_25559,N_23680,N_23809);
and U25560 (N_25560,N_22357,N_22011);
nand U25561 (N_25561,N_22536,N_23585);
and U25562 (N_25562,N_22893,N_22801);
xor U25563 (N_25563,N_23474,N_23067);
or U25564 (N_25564,N_22075,N_23385);
nand U25565 (N_25565,N_23634,N_23743);
or U25566 (N_25566,N_22451,N_23796);
and U25567 (N_25567,N_23223,N_22909);
and U25568 (N_25568,N_22120,N_22887);
nand U25569 (N_25569,N_22218,N_22188);
xnor U25570 (N_25570,N_22072,N_23013);
nand U25571 (N_25571,N_22086,N_23254);
xor U25572 (N_25572,N_23146,N_23322);
or U25573 (N_25573,N_22827,N_22601);
nor U25574 (N_25574,N_23495,N_23737);
and U25575 (N_25575,N_22071,N_22606);
and U25576 (N_25576,N_23743,N_23749);
nand U25577 (N_25577,N_22502,N_22337);
or U25578 (N_25578,N_22230,N_23305);
nor U25579 (N_25579,N_23101,N_22796);
xnor U25580 (N_25580,N_22834,N_23413);
nor U25581 (N_25581,N_22797,N_23688);
nor U25582 (N_25582,N_22976,N_23173);
xor U25583 (N_25583,N_22531,N_22355);
and U25584 (N_25584,N_22697,N_23653);
or U25585 (N_25585,N_23034,N_23768);
nor U25586 (N_25586,N_22962,N_23754);
xor U25587 (N_25587,N_22209,N_23865);
nor U25588 (N_25588,N_23984,N_23968);
nand U25589 (N_25589,N_23072,N_22555);
and U25590 (N_25590,N_22007,N_23063);
nand U25591 (N_25591,N_23452,N_23494);
or U25592 (N_25592,N_22308,N_23365);
and U25593 (N_25593,N_23460,N_23814);
or U25594 (N_25594,N_23666,N_23762);
nor U25595 (N_25595,N_22947,N_23134);
xor U25596 (N_25596,N_22270,N_23256);
nand U25597 (N_25597,N_23157,N_22417);
or U25598 (N_25598,N_22874,N_22334);
nor U25599 (N_25599,N_23204,N_22170);
and U25600 (N_25600,N_23225,N_22371);
nand U25601 (N_25601,N_22013,N_22528);
xor U25602 (N_25602,N_23833,N_22578);
or U25603 (N_25603,N_23425,N_22077);
nand U25604 (N_25604,N_23038,N_23137);
xor U25605 (N_25605,N_23773,N_22056);
or U25606 (N_25606,N_22081,N_22967);
or U25607 (N_25607,N_23667,N_23479);
xor U25608 (N_25608,N_23157,N_23927);
nor U25609 (N_25609,N_23496,N_22038);
or U25610 (N_25610,N_23523,N_22120);
or U25611 (N_25611,N_22336,N_22298);
xor U25612 (N_25612,N_23922,N_22508);
nor U25613 (N_25613,N_22777,N_22683);
and U25614 (N_25614,N_22475,N_22361);
nor U25615 (N_25615,N_22068,N_23945);
and U25616 (N_25616,N_22937,N_23591);
nand U25617 (N_25617,N_22417,N_22880);
nand U25618 (N_25618,N_23289,N_22935);
xor U25619 (N_25619,N_23161,N_23552);
nand U25620 (N_25620,N_22850,N_22198);
and U25621 (N_25621,N_23030,N_23270);
or U25622 (N_25622,N_22736,N_22694);
and U25623 (N_25623,N_23985,N_23267);
xnor U25624 (N_25624,N_22776,N_23074);
xor U25625 (N_25625,N_22957,N_22846);
xor U25626 (N_25626,N_22217,N_23718);
xnor U25627 (N_25627,N_22647,N_22630);
nor U25628 (N_25628,N_22444,N_22285);
nor U25629 (N_25629,N_22859,N_23795);
xnor U25630 (N_25630,N_22727,N_22128);
nand U25631 (N_25631,N_23883,N_23898);
nand U25632 (N_25632,N_22689,N_23391);
xor U25633 (N_25633,N_23062,N_22864);
and U25634 (N_25634,N_22820,N_22950);
xor U25635 (N_25635,N_22345,N_23098);
xnor U25636 (N_25636,N_22523,N_22121);
nor U25637 (N_25637,N_23986,N_22230);
nand U25638 (N_25638,N_22873,N_22009);
nor U25639 (N_25639,N_23447,N_23144);
nor U25640 (N_25640,N_22455,N_23728);
xnor U25641 (N_25641,N_22247,N_23774);
and U25642 (N_25642,N_22862,N_23945);
nand U25643 (N_25643,N_22949,N_22503);
and U25644 (N_25644,N_23183,N_23382);
or U25645 (N_25645,N_23661,N_22885);
or U25646 (N_25646,N_22705,N_23596);
and U25647 (N_25647,N_23469,N_22031);
or U25648 (N_25648,N_22266,N_22285);
nor U25649 (N_25649,N_23902,N_23203);
nand U25650 (N_25650,N_23807,N_23067);
xnor U25651 (N_25651,N_22951,N_22783);
nor U25652 (N_25652,N_22054,N_22112);
and U25653 (N_25653,N_23035,N_22097);
or U25654 (N_25654,N_23944,N_23769);
and U25655 (N_25655,N_22006,N_23880);
nand U25656 (N_25656,N_22055,N_22342);
nand U25657 (N_25657,N_22899,N_22398);
xnor U25658 (N_25658,N_22804,N_22064);
or U25659 (N_25659,N_22562,N_23915);
or U25660 (N_25660,N_23754,N_22518);
nand U25661 (N_25661,N_22944,N_23375);
and U25662 (N_25662,N_23169,N_23963);
and U25663 (N_25663,N_23631,N_23452);
and U25664 (N_25664,N_23156,N_23132);
xor U25665 (N_25665,N_22065,N_23356);
nor U25666 (N_25666,N_23609,N_23234);
or U25667 (N_25667,N_22160,N_22178);
and U25668 (N_25668,N_23960,N_22738);
and U25669 (N_25669,N_22840,N_23760);
nand U25670 (N_25670,N_23302,N_22225);
or U25671 (N_25671,N_22080,N_22247);
nand U25672 (N_25672,N_22300,N_22260);
and U25673 (N_25673,N_22414,N_22302);
and U25674 (N_25674,N_22259,N_23251);
and U25675 (N_25675,N_23892,N_22678);
and U25676 (N_25676,N_22861,N_23759);
nor U25677 (N_25677,N_22709,N_23388);
nor U25678 (N_25678,N_23906,N_22620);
or U25679 (N_25679,N_22499,N_22018);
nor U25680 (N_25680,N_23119,N_22803);
nand U25681 (N_25681,N_22777,N_23024);
nor U25682 (N_25682,N_23436,N_23156);
nor U25683 (N_25683,N_22011,N_23677);
xnor U25684 (N_25684,N_23040,N_22049);
and U25685 (N_25685,N_23229,N_22150);
nor U25686 (N_25686,N_22782,N_22862);
nand U25687 (N_25687,N_22516,N_22816);
xor U25688 (N_25688,N_23340,N_23783);
or U25689 (N_25689,N_23154,N_22267);
nor U25690 (N_25690,N_22356,N_23930);
or U25691 (N_25691,N_23946,N_22218);
or U25692 (N_25692,N_22175,N_23488);
and U25693 (N_25693,N_23879,N_23751);
or U25694 (N_25694,N_22989,N_22294);
xor U25695 (N_25695,N_22783,N_23849);
nor U25696 (N_25696,N_22046,N_23726);
and U25697 (N_25697,N_22148,N_22759);
nor U25698 (N_25698,N_22895,N_23694);
xnor U25699 (N_25699,N_22774,N_23044);
or U25700 (N_25700,N_22000,N_22066);
and U25701 (N_25701,N_23466,N_22457);
or U25702 (N_25702,N_23553,N_23771);
and U25703 (N_25703,N_23056,N_22444);
or U25704 (N_25704,N_23044,N_23474);
xnor U25705 (N_25705,N_22114,N_23167);
or U25706 (N_25706,N_23514,N_23933);
and U25707 (N_25707,N_23755,N_23553);
nor U25708 (N_25708,N_23343,N_22866);
nor U25709 (N_25709,N_23840,N_22748);
xor U25710 (N_25710,N_23503,N_22217);
xnor U25711 (N_25711,N_23310,N_22082);
and U25712 (N_25712,N_22482,N_22702);
nor U25713 (N_25713,N_23270,N_22585);
or U25714 (N_25714,N_22869,N_23897);
xnor U25715 (N_25715,N_23056,N_22864);
nor U25716 (N_25716,N_22647,N_23007);
nor U25717 (N_25717,N_22049,N_22509);
or U25718 (N_25718,N_22489,N_23772);
and U25719 (N_25719,N_23387,N_22718);
or U25720 (N_25720,N_22344,N_22705);
nor U25721 (N_25721,N_23530,N_22269);
nor U25722 (N_25722,N_23481,N_23639);
nor U25723 (N_25723,N_23578,N_23493);
nor U25724 (N_25724,N_22945,N_22948);
nor U25725 (N_25725,N_23084,N_23903);
or U25726 (N_25726,N_22226,N_23264);
and U25727 (N_25727,N_22016,N_22632);
xor U25728 (N_25728,N_23624,N_23918);
or U25729 (N_25729,N_22649,N_23607);
xnor U25730 (N_25730,N_23067,N_23437);
or U25731 (N_25731,N_23590,N_23340);
nand U25732 (N_25732,N_22850,N_23910);
xnor U25733 (N_25733,N_22628,N_23582);
or U25734 (N_25734,N_23041,N_22910);
xor U25735 (N_25735,N_23664,N_22489);
and U25736 (N_25736,N_23660,N_22518);
and U25737 (N_25737,N_22018,N_22170);
nor U25738 (N_25738,N_22141,N_23166);
nand U25739 (N_25739,N_22885,N_22744);
or U25740 (N_25740,N_22980,N_23298);
and U25741 (N_25741,N_23425,N_23866);
xor U25742 (N_25742,N_22352,N_22619);
or U25743 (N_25743,N_22178,N_22813);
and U25744 (N_25744,N_23072,N_23725);
and U25745 (N_25745,N_23169,N_23349);
nand U25746 (N_25746,N_23769,N_22964);
and U25747 (N_25747,N_23903,N_23133);
or U25748 (N_25748,N_22085,N_23477);
and U25749 (N_25749,N_22311,N_23035);
and U25750 (N_25750,N_22650,N_22152);
or U25751 (N_25751,N_23751,N_23798);
nand U25752 (N_25752,N_22939,N_22231);
xor U25753 (N_25753,N_22615,N_22718);
nand U25754 (N_25754,N_23100,N_22200);
nand U25755 (N_25755,N_22027,N_22168);
xnor U25756 (N_25756,N_23417,N_22408);
and U25757 (N_25757,N_22844,N_22226);
nor U25758 (N_25758,N_22599,N_23120);
and U25759 (N_25759,N_22399,N_22410);
or U25760 (N_25760,N_22387,N_23163);
or U25761 (N_25761,N_23858,N_22869);
or U25762 (N_25762,N_23635,N_22004);
or U25763 (N_25763,N_23752,N_23054);
or U25764 (N_25764,N_22312,N_22354);
and U25765 (N_25765,N_23481,N_23253);
or U25766 (N_25766,N_23478,N_22446);
or U25767 (N_25767,N_23100,N_23071);
or U25768 (N_25768,N_22821,N_22110);
and U25769 (N_25769,N_23384,N_23896);
nand U25770 (N_25770,N_22178,N_22557);
xor U25771 (N_25771,N_23343,N_23750);
or U25772 (N_25772,N_23455,N_22383);
nor U25773 (N_25773,N_23160,N_23217);
nor U25774 (N_25774,N_22507,N_22790);
nand U25775 (N_25775,N_22125,N_23684);
and U25776 (N_25776,N_22844,N_23006);
or U25777 (N_25777,N_23621,N_22228);
and U25778 (N_25778,N_22966,N_23920);
and U25779 (N_25779,N_23712,N_22933);
nand U25780 (N_25780,N_23357,N_22767);
and U25781 (N_25781,N_23160,N_23350);
nor U25782 (N_25782,N_22673,N_23990);
or U25783 (N_25783,N_23213,N_23948);
nor U25784 (N_25784,N_23612,N_22326);
or U25785 (N_25785,N_23455,N_23498);
or U25786 (N_25786,N_22136,N_23870);
nand U25787 (N_25787,N_23912,N_23498);
and U25788 (N_25788,N_22800,N_22714);
or U25789 (N_25789,N_22990,N_22570);
and U25790 (N_25790,N_23454,N_22062);
and U25791 (N_25791,N_23633,N_23936);
nor U25792 (N_25792,N_22053,N_23993);
or U25793 (N_25793,N_22380,N_23576);
nand U25794 (N_25794,N_22775,N_23357);
xor U25795 (N_25795,N_23921,N_23781);
nand U25796 (N_25796,N_22222,N_23707);
and U25797 (N_25797,N_22297,N_22400);
nand U25798 (N_25798,N_23834,N_23068);
nand U25799 (N_25799,N_22879,N_22801);
nand U25800 (N_25800,N_23949,N_22841);
and U25801 (N_25801,N_22066,N_23558);
xor U25802 (N_25802,N_22615,N_22762);
or U25803 (N_25803,N_22439,N_22450);
nand U25804 (N_25804,N_22643,N_23087);
or U25805 (N_25805,N_22116,N_22183);
and U25806 (N_25806,N_22255,N_22251);
or U25807 (N_25807,N_23172,N_22301);
nor U25808 (N_25808,N_22917,N_23864);
xor U25809 (N_25809,N_23050,N_23140);
nor U25810 (N_25810,N_22842,N_23786);
and U25811 (N_25811,N_22572,N_22201);
nand U25812 (N_25812,N_22169,N_22852);
nand U25813 (N_25813,N_23075,N_23384);
nand U25814 (N_25814,N_23907,N_23727);
nor U25815 (N_25815,N_23405,N_22465);
nand U25816 (N_25816,N_23585,N_22017);
nand U25817 (N_25817,N_23622,N_22606);
or U25818 (N_25818,N_22929,N_23516);
and U25819 (N_25819,N_23218,N_23084);
nor U25820 (N_25820,N_22670,N_23384);
xor U25821 (N_25821,N_22623,N_23029);
nor U25822 (N_25822,N_22622,N_22778);
nand U25823 (N_25823,N_22954,N_22046);
nor U25824 (N_25824,N_22959,N_23656);
and U25825 (N_25825,N_22558,N_22372);
nor U25826 (N_25826,N_22210,N_22538);
nand U25827 (N_25827,N_23518,N_23152);
xor U25828 (N_25828,N_22282,N_23200);
nor U25829 (N_25829,N_23029,N_23686);
xor U25830 (N_25830,N_22910,N_23447);
and U25831 (N_25831,N_23770,N_23108);
and U25832 (N_25832,N_22994,N_22901);
xor U25833 (N_25833,N_22778,N_23773);
and U25834 (N_25834,N_23230,N_23099);
nand U25835 (N_25835,N_22982,N_23969);
nand U25836 (N_25836,N_22944,N_23673);
nor U25837 (N_25837,N_23694,N_23668);
and U25838 (N_25838,N_23902,N_22195);
or U25839 (N_25839,N_22398,N_23324);
xnor U25840 (N_25840,N_23560,N_22278);
nor U25841 (N_25841,N_22416,N_22672);
and U25842 (N_25842,N_23890,N_22266);
or U25843 (N_25843,N_23142,N_22581);
nor U25844 (N_25844,N_22708,N_23226);
nand U25845 (N_25845,N_23859,N_23291);
and U25846 (N_25846,N_23875,N_23518);
or U25847 (N_25847,N_22915,N_23096);
or U25848 (N_25848,N_22306,N_22863);
nand U25849 (N_25849,N_22622,N_22722);
xnor U25850 (N_25850,N_22976,N_22165);
and U25851 (N_25851,N_23433,N_23657);
nor U25852 (N_25852,N_22904,N_22058);
or U25853 (N_25853,N_23869,N_23020);
nand U25854 (N_25854,N_23121,N_23639);
nor U25855 (N_25855,N_22714,N_22218);
and U25856 (N_25856,N_23918,N_23106);
nand U25857 (N_25857,N_23673,N_23342);
xor U25858 (N_25858,N_23132,N_22345);
and U25859 (N_25859,N_22376,N_22733);
xnor U25860 (N_25860,N_23425,N_23630);
nand U25861 (N_25861,N_22451,N_22492);
nor U25862 (N_25862,N_23536,N_22041);
or U25863 (N_25863,N_22850,N_23533);
or U25864 (N_25864,N_23342,N_22312);
nor U25865 (N_25865,N_22831,N_23583);
nand U25866 (N_25866,N_23569,N_23591);
and U25867 (N_25867,N_22456,N_23466);
nor U25868 (N_25868,N_22520,N_23033);
nand U25869 (N_25869,N_23189,N_23913);
or U25870 (N_25870,N_22571,N_22572);
and U25871 (N_25871,N_22694,N_22130);
or U25872 (N_25872,N_22497,N_22130);
or U25873 (N_25873,N_23366,N_23237);
xor U25874 (N_25874,N_22131,N_22455);
nor U25875 (N_25875,N_23927,N_22019);
xnor U25876 (N_25876,N_23702,N_22327);
xor U25877 (N_25877,N_22781,N_23677);
xor U25878 (N_25878,N_22373,N_22725);
or U25879 (N_25879,N_23028,N_23752);
or U25880 (N_25880,N_22968,N_22239);
nor U25881 (N_25881,N_23227,N_22100);
or U25882 (N_25882,N_23131,N_22549);
and U25883 (N_25883,N_23250,N_23479);
xor U25884 (N_25884,N_22888,N_23175);
nor U25885 (N_25885,N_23838,N_22937);
and U25886 (N_25886,N_22485,N_23079);
or U25887 (N_25887,N_22330,N_23674);
nand U25888 (N_25888,N_23033,N_22527);
and U25889 (N_25889,N_22260,N_22887);
or U25890 (N_25890,N_23979,N_22792);
nand U25891 (N_25891,N_23763,N_23022);
xor U25892 (N_25892,N_22791,N_22663);
nor U25893 (N_25893,N_23922,N_23269);
or U25894 (N_25894,N_23847,N_22301);
nor U25895 (N_25895,N_22197,N_23968);
nor U25896 (N_25896,N_23433,N_23203);
nor U25897 (N_25897,N_22335,N_23724);
or U25898 (N_25898,N_22528,N_23708);
xor U25899 (N_25899,N_22968,N_22062);
nor U25900 (N_25900,N_23650,N_23837);
xor U25901 (N_25901,N_22312,N_22290);
nor U25902 (N_25902,N_22263,N_23462);
xnor U25903 (N_25903,N_22068,N_23407);
and U25904 (N_25904,N_22619,N_23806);
xnor U25905 (N_25905,N_22279,N_22270);
xnor U25906 (N_25906,N_22752,N_23996);
nand U25907 (N_25907,N_23451,N_23607);
or U25908 (N_25908,N_22114,N_23044);
nor U25909 (N_25909,N_22546,N_22975);
xnor U25910 (N_25910,N_23662,N_23990);
xnor U25911 (N_25911,N_23831,N_22079);
or U25912 (N_25912,N_23643,N_23591);
or U25913 (N_25913,N_22109,N_23662);
xor U25914 (N_25914,N_23196,N_22494);
and U25915 (N_25915,N_22605,N_22521);
or U25916 (N_25916,N_22509,N_22746);
or U25917 (N_25917,N_23062,N_23315);
and U25918 (N_25918,N_23512,N_22665);
nor U25919 (N_25919,N_23564,N_23640);
nor U25920 (N_25920,N_23088,N_22755);
or U25921 (N_25921,N_23094,N_23737);
or U25922 (N_25922,N_23186,N_23442);
and U25923 (N_25923,N_22346,N_22018);
and U25924 (N_25924,N_22886,N_23208);
or U25925 (N_25925,N_22807,N_22943);
nand U25926 (N_25926,N_22747,N_22039);
nor U25927 (N_25927,N_22811,N_23053);
nor U25928 (N_25928,N_22343,N_22149);
nor U25929 (N_25929,N_23593,N_23559);
and U25930 (N_25930,N_23399,N_22157);
xor U25931 (N_25931,N_23082,N_23727);
or U25932 (N_25932,N_22917,N_22182);
nand U25933 (N_25933,N_22229,N_22660);
or U25934 (N_25934,N_23882,N_23778);
or U25935 (N_25935,N_22462,N_23250);
nand U25936 (N_25936,N_23702,N_23575);
and U25937 (N_25937,N_22207,N_23715);
or U25938 (N_25938,N_22625,N_22888);
nor U25939 (N_25939,N_23055,N_22729);
nor U25940 (N_25940,N_22479,N_22759);
nand U25941 (N_25941,N_22751,N_23818);
or U25942 (N_25942,N_22920,N_23946);
xor U25943 (N_25943,N_23448,N_23444);
xnor U25944 (N_25944,N_22410,N_23815);
and U25945 (N_25945,N_23882,N_22028);
or U25946 (N_25946,N_23087,N_22545);
or U25947 (N_25947,N_23494,N_22065);
or U25948 (N_25948,N_23588,N_23937);
and U25949 (N_25949,N_22518,N_22540);
nand U25950 (N_25950,N_22618,N_22111);
xor U25951 (N_25951,N_22255,N_23850);
xor U25952 (N_25952,N_23622,N_22428);
nor U25953 (N_25953,N_23007,N_23714);
nand U25954 (N_25954,N_23462,N_22249);
xnor U25955 (N_25955,N_22976,N_22398);
nand U25956 (N_25956,N_22816,N_22885);
nor U25957 (N_25957,N_23088,N_22662);
nor U25958 (N_25958,N_23129,N_22759);
or U25959 (N_25959,N_23960,N_23021);
xnor U25960 (N_25960,N_23284,N_23319);
and U25961 (N_25961,N_22009,N_23484);
nand U25962 (N_25962,N_23985,N_22754);
xnor U25963 (N_25963,N_23131,N_22642);
or U25964 (N_25964,N_23228,N_22618);
and U25965 (N_25965,N_22879,N_22342);
or U25966 (N_25966,N_23138,N_23896);
and U25967 (N_25967,N_23719,N_22255);
and U25968 (N_25968,N_22648,N_22330);
nand U25969 (N_25969,N_23990,N_23020);
nand U25970 (N_25970,N_22106,N_22369);
nand U25971 (N_25971,N_22287,N_23536);
and U25972 (N_25972,N_22978,N_22931);
nand U25973 (N_25973,N_23235,N_22814);
or U25974 (N_25974,N_22429,N_22541);
nand U25975 (N_25975,N_23800,N_22424);
xnor U25976 (N_25976,N_23068,N_22267);
and U25977 (N_25977,N_22475,N_23159);
xor U25978 (N_25978,N_22841,N_22665);
nor U25979 (N_25979,N_23709,N_22811);
xnor U25980 (N_25980,N_22325,N_23025);
or U25981 (N_25981,N_22463,N_23508);
xor U25982 (N_25982,N_23200,N_23093);
and U25983 (N_25983,N_22475,N_23537);
nor U25984 (N_25984,N_22276,N_23891);
or U25985 (N_25985,N_22173,N_23458);
or U25986 (N_25986,N_23368,N_22664);
xnor U25987 (N_25987,N_23366,N_23229);
nor U25988 (N_25988,N_22736,N_23684);
xor U25989 (N_25989,N_23004,N_23181);
nor U25990 (N_25990,N_22934,N_22407);
nand U25991 (N_25991,N_23746,N_23483);
nand U25992 (N_25992,N_23970,N_22917);
nand U25993 (N_25993,N_22709,N_23930);
nand U25994 (N_25994,N_23919,N_23118);
or U25995 (N_25995,N_23589,N_23143);
nand U25996 (N_25996,N_23343,N_23252);
xnor U25997 (N_25997,N_22580,N_23143);
or U25998 (N_25998,N_23222,N_23982);
or U25999 (N_25999,N_22093,N_23519);
nor U26000 (N_26000,N_24668,N_25327);
nor U26001 (N_26001,N_25965,N_25715);
or U26002 (N_26002,N_24683,N_24270);
nor U26003 (N_26003,N_25098,N_24792);
xor U26004 (N_26004,N_24832,N_24046);
xor U26005 (N_26005,N_24526,N_24685);
nor U26006 (N_26006,N_24403,N_25100);
or U26007 (N_26007,N_24550,N_25358);
xor U26008 (N_26008,N_25042,N_25078);
and U26009 (N_26009,N_24687,N_25671);
and U26010 (N_26010,N_24873,N_25780);
xor U26011 (N_26011,N_24437,N_24260);
and U26012 (N_26012,N_24208,N_24932);
xnor U26013 (N_26013,N_25713,N_25422);
nor U26014 (N_26014,N_24926,N_25204);
or U26015 (N_26015,N_25873,N_25882);
xor U26016 (N_26016,N_25834,N_25524);
and U26017 (N_26017,N_24388,N_25970);
nand U26018 (N_26018,N_24364,N_24765);
or U26019 (N_26019,N_24645,N_25310);
xor U26020 (N_26020,N_24348,N_24265);
xor U26021 (N_26021,N_24065,N_25433);
or U26022 (N_26022,N_24961,N_24551);
nor U26023 (N_26023,N_25244,N_24872);
or U26024 (N_26024,N_24578,N_24693);
nand U26025 (N_26025,N_24168,N_24642);
nor U26026 (N_26026,N_24037,N_25034);
nor U26027 (N_26027,N_25370,N_24071);
nand U26028 (N_26028,N_24831,N_24589);
or U26029 (N_26029,N_25598,N_25961);
nand U26030 (N_26030,N_24453,N_25664);
xnor U26031 (N_26031,N_24710,N_25302);
nor U26032 (N_26032,N_24288,N_24828);
or U26033 (N_26033,N_24843,N_24225);
and U26034 (N_26034,N_24134,N_24660);
or U26035 (N_26035,N_24555,N_24395);
or U26036 (N_26036,N_25460,N_25663);
nor U26037 (N_26037,N_25219,N_24301);
and U26038 (N_26038,N_25083,N_25823);
nor U26039 (N_26039,N_24804,N_25454);
nor U26040 (N_26040,N_25164,N_25643);
nand U26041 (N_26041,N_25946,N_24465);
nand U26042 (N_26042,N_25818,N_24684);
and U26043 (N_26043,N_25580,N_25110);
xor U26044 (N_26044,N_24153,N_25257);
nand U26045 (N_26045,N_24862,N_24101);
xnor U26046 (N_26046,N_24688,N_24974);
or U26047 (N_26047,N_25359,N_25594);
nand U26048 (N_26048,N_25046,N_25876);
nor U26049 (N_26049,N_24682,N_25005);
nand U26050 (N_26050,N_24838,N_25154);
xor U26051 (N_26051,N_24175,N_24519);
and U26052 (N_26052,N_24739,N_25155);
nor U26053 (N_26053,N_25086,N_25716);
nor U26054 (N_26054,N_25077,N_25440);
or U26055 (N_26055,N_24598,N_25957);
xnor U26056 (N_26056,N_25981,N_24888);
xor U26057 (N_26057,N_24864,N_24402);
nand U26058 (N_26058,N_25602,N_25347);
nor U26059 (N_26059,N_24481,N_24671);
and U26060 (N_26060,N_24359,N_25536);
and U26061 (N_26061,N_24060,N_25812);
xor U26062 (N_26062,N_24777,N_24507);
xor U26063 (N_26063,N_25101,N_24331);
or U26064 (N_26064,N_24539,N_25528);
nand U26065 (N_26065,N_25997,N_24059);
nor U26066 (N_26066,N_25316,N_25803);
nor U26067 (N_26067,N_25660,N_25915);
and U26068 (N_26068,N_25557,N_25597);
nand U26069 (N_26069,N_25609,N_24869);
and U26070 (N_26070,N_25608,N_25260);
and U26071 (N_26071,N_24074,N_25396);
nand U26072 (N_26072,N_24149,N_24942);
and U26073 (N_26073,N_24773,N_24618);
and U26074 (N_26074,N_25994,N_25030);
nor U26075 (N_26075,N_24644,N_24929);
and U26076 (N_26076,N_24849,N_24103);
and U26077 (N_26077,N_25831,N_25453);
or U26078 (N_26078,N_24444,N_24963);
nand U26079 (N_26079,N_24615,N_25613);
xor U26080 (N_26080,N_25895,N_24523);
and U26081 (N_26081,N_25242,N_25035);
nor U26082 (N_26082,N_25161,N_24357);
xor U26083 (N_26083,N_25920,N_24323);
or U26084 (N_26084,N_24081,N_24480);
nand U26085 (N_26085,N_25369,N_24006);
nor U26086 (N_26086,N_25027,N_25567);
xor U26087 (N_26087,N_24498,N_24104);
nor U26088 (N_26088,N_25292,N_25427);
nand U26089 (N_26089,N_24553,N_25906);
or U26090 (N_26090,N_25145,N_24649);
and U26091 (N_26091,N_25804,N_25061);
or U26092 (N_26092,N_24844,N_25297);
or U26093 (N_26093,N_25252,N_25748);
nand U26094 (N_26094,N_25320,N_25227);
or U26095 (N_26095,N_24312,N_25833);
xor U26096 (N_26096,N_25733,N_25406);
xor U26097 (N_26097,N_25502,N_25714);
nor U26098 (N_26098,N_25472,N_25019);
or U26099 (N_26099,N_25696,N_25197);
xor U26100 (N_26100,N_24825,N_24646);
and U26101 (N_26101,N_24631,N_24425);
nand U26102 (N_26102,N_24909,N_24390);
nand U26103 (N_26103,N_24440,N_24385);
or U26104 (N_26104,N_24545,N_25091);
or U26105 (N_26105,N_24500,N_25317);
nand U26106 (N_26106,N_25312,N_24442);
xnor U26107 (N_26107,N_25857,N_24012);
or U26108 (N_26108,N_25562,N_25322);
xor U26109 (N_26109,N_25796,N_25973);
xor U26110 (N_26110,N_25827,N_24297);
nor U26111 (N_26111,N_24040,N_25868);
or U26112 (N_26112,N_24987,N_25616);
and U26113 (N_26113,N_25699,N_25097);
or U26114 (N_26114,N_24800,N_25072);
or U26115 (N_26115,N_24592,N_24508);
nand U26116 (N_26116,N_25314,N_24347);
or U26117 (N_26117,N_24470,N_24053);
xor U26118 (N_26118,N_24345,N_24915);
and U26119 (N_26119,N_25159,N_25636);
nand U26120 (N_26120,N_24484,N_24491);
nand U26121 (N_26121,N_25753,N_24572);
nand U26122 (N_26122,N_24077,N_24501);
xnor U26123 (N_26123,N_24712,N_24320);
or U26124 (N_26124,N_25913,N_25122);
and U26125 (N_26125,N_25245,N_25179);
and U26126 (N_26126,N_24585,N_25631);
or U26127 (N_26127,N_24304,N_25281);
nand U26128 (N_26128,N_25196,N_25905);
or U26129 (N_26129,N_25492,N_24925);
nand U26130 (N_26130,N_24628,N_24336);
and U26131 (N_26131,N_24866,N_25866);
nand U26132 (N_26132,N_25986,N_24656);
nor U26133 (N_26133,N_25646,N_24289);
or U26134 (N_26134,N_24456,N_25425);
and U26135 (N_26135,N_24709,N_24976);
xnor U26136 (N_26136,N_25150,N_24881);
nor U26137 (N_26137,N_25191,N_25162);
nor U26138 (N_26138,N_25548,N_24159);
xnor U26139 (N_26139,N_24492,N_24648);
xor U26140 (N_26140,N_25878,N_25661);
nand U26141 (N_26141,N_24830,N_25898);
nor U26142 (N_26142,N_25720,N_25681);
and U26143 (N_26143,N_25654,N_24476);
or U26144 (N_26144,N_25067,N_24185);
nor U26145 (N_26145,N_24079,N_25686);
nor U26146 (N_26146,N_24788,N_24227);
or U26147 (N_26147,N_25416,N_24349);
or U26148 (N_26148,N_24769,N_24180);
nor U26149 (N_26149,N_24970,N_25233);
and U26150 (N_26150,N_24250,N_25424);
nand U26151 (N_26151,N_25647,N_25478);
xor U26152 (N_26152,N_25216,N_24150);
or U26153 (N_26153,N_24894,N_24760);
or U26154 (N_26154,N_24510,N_24051);
xnor U26155 (N_26155,N_25723,N_25773);
or U26156 (N_26156,N_24827,N_24382);
nand U26157 (N_26157,N_24174,N_25797);
nand U26158 (N_26158,N_24766,N_25366);
or U26159 (N_26159,N_25467,N_25530);
nand U26160 (N_26160,N_24055,N_25635);
nand U26161 (N_26161,N_25372,N_24067);
nand U26162 (N_26162,N_25465,N_24198);
or U26163 (N_26163,N_24415,N_25822);
nor U26164 (N_26164,N_24647,N_25344);
and U26165 (N_26165,N_24940,N_24494);
and U26166 (N_26166,N_24334,N_25020);
nand U26167 (N_26167,N_25193,N_25328);
and U26168 (N_26168,N_25793,N_25657);
nand U26169 (N_26169,N_24354,N_24262);
nand U26170 (N_26170,N_24002,N_25195);
nand U26171 (N_26171,N_24719,N_25764);
or U26172 (N_26172,N_24109,N_25397);
xnor U26173 (N_26173,N_25023,N_24749);
nor U26174 (N_26174,N_24590,N_24398);
or U26175 (N_26175,N_25772,N_25350);
or U26176 (N_26176,N_25939,N_25937);
nand U26177 (N_26177,N_24633,N_25186);
nand U26178 (N_26178,N_25121,N_24392);
and U26179 (N_26179,N_25256,N_25504);
xnor U26180 (N_26180,N_24840,N_25177);
nor U26181 (N_26181,N_25304,N_24050);
nand U26182 (N_26182,N_25093,N_24732);
xnor U26183 (N_26183,N_24254,N_24112);
xnor U26184 (N_26184,N_25871,N_24764);
or U26185 (N_26185,N_25948,N_25556);
xor U26186 (N_26186,N_25171,N_25590);
nor U26187 (N_26187,N_25208,N_24249);
and U26188 (N_26188,N_25691,N_25514);
nand U26189 (N_26189,N_25968,N_24271);
xor U26190 (N_26190,N_24898,N_24171);
and U26191 (N_26191,N_25993,N_25750);
nand U26192 (N_26192,N_24007,N_24230);
nand U26193 (N_26193,N_25375,N_24218);
nor U26194 (N_26194,N_25865,N_24815);
xnor U26195 (N_26195,N_24938,N_24913);
and U26196 (N_26196,N_24094,N_24975);
or U26197 (N_26197,N_24459,N_25054);
nand U26198 (N_26198,N_25729,N_24653);
nand U26199 (N_26199,N_24274,N_24667);
xor U26200 (N_26200,N_25363,N_24243);
nor U26201 (N_26201,N_24386,N_24856);
nor U26202 (N_26202,N_24641,N_24161);
xor U26203 (N_26203,N_25578,N_25143);
nand U26204 (N_26204,N_24816,N_24814);
xnor U26205 (N_26205,N_24039,N_25711);
nand U26206 (N_26206,N_24833,N_25830);
xnor U26207 (N_26207,N_25167,N_24286);
and U26208 (N_26208,N_25684,N_25785);
nand U26209 (N_26209,N_24203,N_24214);
and U26210 (N_26210,N_24763,N_25658);
or U26211 (N_26211,N_24114,N_24473);
and U26212 (N_26212,N_25979,N_25769);
nor U26213 (N_26213,N_24160,N_24457);
and U26214 (N_26214,N_24583,N_24436);
nand U26215 (N_26215,N_25169,N_25289);
and U26216 (N_26216,N_25763,N_24307);
and U26217 (N_26217,N_24619,N_24129);
nand U26218 (N_26218,N_25563,N_25574);
nor U26219 (N_26219,N_24266,N_24340);
xor U26220 (N_26220,N_24697,N_25561);
xnor U26221 (N_26221,N_24559,N_24217);
or U26222 (N_26222,N_24098,N_24352);
nor U26223 (N_26223,N_24310,N_25974);
nor U26224 (N_26224,N_25168,N_24655);
nand U26225 (N_26225,N_24933,N_25253);
or U26226 (N_26226,N_24955,N_24524);
nand U26227 (N_26227,N_24229,N_24487);
and U26228 (N_26228,N_25910,N_24704);
and U26229 (N_26229,N_24389,N_25479);
nand U26230 (N_26230,N_25632,N_24499);
or U26231 (N_26231,N_25498,N_24634);
or U26232 (N_26232,N_25303,N_25450);
nor U26233 (N_26233,N_24004,N_25903);
and U26234 (N_26234,N_24504,N_25102);
or U26235 (N_26235,N_24371,N_24045);
nor U26236 (N_26236,N_25047,N_24700);
and U26237 (N_26237,N_24096,N_25825);
and U26238 (N_26238,N_24309,N_24991);
or U26239 (N_26239,N_25886,N_25881);
or U26240 (N_26240,N_24698,N_24367);
xnor U26241 (N_26241,N_25079,N_24597);
and U26242 (N_26242,N_25092,N_25458);
and U26243 (N_26243,N_24968,N_25008);
or U26244 (N_26244,N_25839,N_25860);
nand U26245 (N_26245,N_25551,N_25051);
or U26246 (N_26246,N_25338,N_24242);
and U26247 (N_26247,N_25954,N_24326);
or U26248 (N_26248,N_24089,N_25940);
xor U26249 (N_26249,N_25984,N_24443);
or U26250 (N_26250,N_25953,N_24210);
xnor U26251 (N_26251,N_24192,N_24267);
xnor U26252 (N_26252,N_25325,N_24853);
nor U26253 (N_26253,N_24374,N_24522);
or U26254 (N_26254,N_24735,N_24582);
xor U26255 (N_26255,N_25787,N_24954);
nand U26256 (N_26256,N_24958,N_24867);
xnor U26257 (N_26257,N_25529,N_24496);
nand U26258 (N_26258,N_25355,N_25447);
nand U26259 (N_26259,N_25048,N_25956);
nor U26260 (N_26260,N_25717,N_25904);
nor U26261 (N_26261,N_24011,N_24085);
or U26262 (N_26262,N_24211,N_24541);
and U26263 (N_26263,N_25284,N_24802);
xnor U26264 (N_26264,N_24406,N_25482);
or U26265 (N_26265,N_25651,N_24676);
nor U26266 (N_26266,N_24823,N_24429);
or U26267 (N_26267,N_24497,N_24734);
xnor U26268 (N_26268,N_24027,N_24713);
nor U26269 (N_26269,N_25213,N_24943);
or U26270 (N_26270,N_24745,N_25761);
xor U26271 (N_26271,N_25737,N_24154);
nor U26272 (N_26272,N_25487,N_24770);
xnor U26273 (N_26273,N_24222,N_25864);
and U26274 (N_26274,N_25200,N_25669);
and U26275 (N_26275,N_25921,N_25928);
nor U26276 (N_26276,N_25689,N_24474);
nor U26277 (N_26277,N_24675,N_24635);
and U26278 (N_26278,N_25214,N_24957);
and U26279 (N_26279,N_25765,N_24950);
xor U26280 (N_26280,N_25601,N_24155);
nand U26281 (N_26281,N_25138,N_24624);
nand U26282 (N_26282,N_24977,N_24384);
or U26283 (N_26283,N_24543,N_24612);
and U26284 (N_26284,N_24455,N_24517);
or U26285 (N_26285,N_24706,N_25998);
nand U26286 (N_26286,N_25988,N_24681);
nand U26287 (N_26287,N_25523,N_25241);
or U26288 (N_26288,N_24311,N_24292);
or U26289 (N_26289,N_24461,N_24291);
nor U26290 (N_26290,N_24725,N_24337);
nor U26291 (N_26291,N_25116,N_25118);
nor U26292 (N_26292,N_25489,N_24280);
nor U26293 (N_26293,N_25365,N_24136);
nand U26294 (N_26294,N_25468,N_25648);
nand U26295 (N_26295,N_25298,N_25045);
xnor U26296 (N_26296,N_24490,N_25001);
and U26297 (N_26297,N_24730,N_24695);
nor U26298 (N_26298,N_25688,N_25418);
nor U26299 (N_26299,N_25929,N_25739);
nor U26300 (N_26300,N_25942,N_24141);
xnor U26301 (N_26301,N_25476,N_25080);
and U26302 (N_26302,N_24601,N_25278);
or U26303 (N_26303,N_24871,N_25778);
or U26304 (N_26304,N_24509,N_25128);
or U26305 (N_26305,N_24353,N_25238);
and U26306 (N_26306,N_25388,N_25995);
nor U26307 (N_26307,N_24741,N_25519);
xnor U26308 (N_26308,N_24177,N_24690);
or U26309 (N_26309,N_25883,N_24478);
or U26310 (N_26310,N_24076,N_24215);
nand U26311 (N_26311,N_25901,N_24021);
nand U26312 (N_26312,N_24917,N_24463);
or U26313 (N_26313,N_25287,N_24813);
or U26314 (N_26314,N_24801,N_24547);
or U26315 (N_26315,N_24910,N_25638);
xor U26316 (N_26316,N_24277,N_24819);
and U26317 (N_26317,N_24163,N_25889);
nand U26318 (N_26318,N_24752,N_24632);
nor U26319 (N_26319,N_24886,N_25362);
nand U26320 (N_26320,N_24944,N_25849);
nor U26321 (N_26321,N_24300,N_24783);
and U26322 (N_26322,N_25675,N_24761);
xnor U26323 (N_26323,N_24934,N_24213);
nor U26324 (N_26324,N_25496,N_25277);
nand U26325 (N_26325,N_24179,N_24235);
or U26326 (N_26326,N_25539,N_24654);
nor U26327 (N_26327,N_25540,N_25002);
and U26328 (N_26328,N_24658,N_25622);
nor U26329 (N_26329,N_25917,N_24084);
nand U26330 (N_26330,N_24922,N_25776);
xnor U26331 (N_26331,N_24308,N_25781);
xor U26332 (N_26332,N_25335,N_25826);
nor U26333 (N_26333,N_25326,N_24124);
or U26334 (N_26334,N_24475,N_24187);
nand U26335 (N_26335,N_25612,N_25391);
xnor U26336 (N_26336,N_24471,N_25767);
nor U26337 (N_26337,N_25576,N_24998);
or U26338 (N_26338,N_24596,N_25249);
nor U26339 (N_26339,N_24355,N_24803);
or U26340 (N_26340,N_24912,N_24606);
xor U26341 (N_26341,N_24772,N_25718);
and U26342 (N_26342,N_25291,N_25125);
nand U26343 (N_26343,N_25206,N_25924);
or U26344 (N_26344,N_24863,N_24907);
xnor U26345 (N_26345,N_24806,N_24530);
nor U26346 (N_26346,N_25914,N_25059);
nor U26347 (N_26347,N_25095,N_24184);
xnor U26348 (N_26348,N_24993,N_24248);
xor U26349 (N_26349,N_25301,N_24614);
nor U26350 (N_26350,N_24275,N_24052);
xnor U26351 (N_26351,N_25798,N_25403);
xor U26352 (N_26352,N_24268,N_24762);
nor U26353 (N_26353,N_24042,N_25198);
and U26354 (N_26354,N_25599,N_24350);
xnor U26355 (N_26355,N_24768,N_24736);
or U26356 (N_26356,N_24015,N_24148);
or U26357 (N_26357,N_25076,N_24727);
and U26358 (N_26358,N_25336,N_24452);
or U26359 (N_26359,N_25432,N_25633);
and U26360 (N_26360,N_25999,N_24822);
nor U26361 (N_26361,N_25624,N_25157);
xnor U26362 (N_26362,N_25400,N_25248);
or U26363 (N_26363,N_25486,N_25107);
xor U26364 (N_26364,N_24043,N_25677);
nand U26365 (N_26365,N_24733,N_25853);
xor U26366 (N_26366,N_24379,N_24850);
xnor U26367 (N_26367,N_25908,N_25843);
nand U26368 (N_26368,N_25891,N_24721);
and U26369 (N_26369,N_24902,N_24132);
or U26370 (N_26370,N_24238,N_24256);
xnor U26371 (N_26371,N_25783,N_25415);
nor U26372 (N_26372,N_24505,N_25096);
nand U26373 (N_26373,N_24221,N_25232);
and U26374 (N_26374,N_25503,N_25220);
xnor U26375 (N_26375,N_25892,N_24834);
or U26376 (N_26376,N_25189,N_25659);
xor U26377 (N_26377,N_24102,N_24568);
nand U26378 (N_26378,N_25043,N_24092);
nor U26379 (N_26379,N_24513,N_25559);
nand U26380 (N_26380,N_24754,N_25473);
and U26381 (N_26381,N_24692,N_24707);
nor U26382 (N_26382,N_25832,N_24125);
nand U26383 (N_26383,N_25614,N_24278);
and U26384 (N_26384,N_24897,N_24140);
and U26385 (N_26385,N_24376,N_24186);
nor U26386 (N_26386,N_25377,N_25215);
or U26387 (N_26387,N_25817,N_25258);
nand U26388 (N_26388,N_24924,N_25131);
nor U26389 (N_26389,N_25735,N_25603);
or U26390 (N_26390,N_25705,N_25199);
and U26391 (N_26391,N_25394,N_24514);
and U26392 (N_26392,N_25499,N_25084);
nor U26393 (N_26393,N_24023,N_25174);
or U26394 (N_26394,N_24257,N_24144);
or U26395 (N_26395,N_24423,N_24407);
and U26396 (N_26396,N_24380,N_24691);
and U26397 (N_26397,N_25119,N_25931);
and U26398 (N_26398,N_24314,N_24558);
or U26399 (N_26399,N_25751,N_25068);
and U26400 (N_26400,N_25057,N_25533);
nand U26401 (N_26401,N_24338,N_24771);
nand U26402 (N_26402,N_24370,N_25160);
and U26403 (N_26403,N_24036,N_25240);
xnor U26404 (N_26404,N_24193,N_24296);
nand U26405 (N_26405,N_24665,N_24057);
or U26406 (N_26406,N_24176,N_25149);
nor U26407 (N_26407,N_24346,N_24900);
xnor U26408 (N_26408,N_25952,N_25000);
and U26409 (N_26409,N_25025,N_25202);
xnor U26410 (N_26410,N_24188,N_24896);
nor U26411 (N_26411,N_25069,N_24714);
or U26412 (N_26412,N_25139,N_24329);
and U26413 (N_26413,N_25401,N_25254);
nand U26414 (N_26414,N_24466,N_25829);
nand U26415 (N_26415,N_25156,N_24810);
nand U26416 (N_26416,N_25604,N_25879);
nor U26417 (N_26417,N_24638,N_24784);
and U26418 (N_26418,N_25560,N_24626);
nand U26419 (N_26419,N_24737,N_24797);
xnor U26420 (N_26420,N_25074,N_25457);
nor U26421 (N_26421,N_24506,N_24990);
nand U26422 (N_26422,N_25480,N_24117);
xnor U26423 (N_26423,N_25462,N_24041);
xor U26424 (N_26424,N_24333,N_24273);
and U26425 (N_26425,N_25270,N_24200);
nand U26426 (N_26426,N_25211,N_25987);
xor U26427 (N_26427,N_24010,N_25842);
and U26428 (N_26428,N_25615,N_24495);
xor U26429 (N_26429,N_24876,N_24600);
or U26430 (N_26430,N_25869,N_24972);
and U26431 (N_26431,N_24696,N_25407);
nor U26432 (N_26432,N_25029,N_24946);
and U26433 (N_26433,N_25938,N_25591);
nand U26434 (N_26434,N_25740,N_24244);
nor U26435 (N_26435,N_25858,N_25040);
and U26436 (N_26436,N_24608,N_25926);
xor U26437 (N_26437,N_25332,N_25863);
or U26438 (N_26438,N_25255,N_25743);
xor U26439 (N_26439,N_24135,N_24083);
and U26440 (N_26440,N_24557,N_24616);
nand U26441 (N_26441,N_24162,N_24928);
or U26442 (N_26442,N_24575,N_25176);
or U26443 (N_26443,N_25449,N_25746);
and U26444 (N_26444,N_25438,N_24908);
nand U26445 (N_26445,N_24018,N_24556);
xor U26446 (N_26446,N_24584,N_25280);
xor U26447 (N_26447,N_24841,N_25777);
nand U26448 (N_26448,N_24317,N_24272);
nor U26449 (N_26449,N_24165,N_25813);
nor U26450 (N_26450,N_24378,N_25726);
nand U26451 (N_26451,N_25836,N_25958);
xnor U26452 (N_26452,N_25137,N_25634);
nor U26453 (N_26453,N_25044,N_25203);
nor U26454 (N_26454,N_24428,N_24047);
or U26455 (N_26455,N_24574,N_25847);
xnor U26456 (N_26456,N_24534,N_25538);
or U26457 (N_26457,N_25461,N_25809);
nor U26458 (N_26458,N_24486,N_25855);
xnor U26459 (N_26459,N_25299,N_25337);
and U26460 (N_26460,N_24283,N_24857);
xnor U26461 (N_26461,N_24003,N_25972);
or U26462 (N_26462,N_25759,N_24781);
xnor U26463 (N_26463,N_24791,N_25413);
nor U26464 (N_26464,N_25334,N_25437);
and U26465 (N_26465,N_24138,N_24662);
and U26466 (N_26466,N_25704,N_25201);
and U26467 (N_26467,N_24462,N_25824);
or U26468 (N_26468,N_25525,N_24643);
xor U26469 (N_26469,N_24580,N_25545);
xor U26470 (N_26470,N_25349,N_25862);
or U26471 (N_26471,N_25782,N_24468);
and U26472 (N_26472,N_25587,N_24664);
or U26473 (N_26473,N_25786,N_24879);
and U26474 (N_26474,N_25147,N_24670);
xnor U26475 (N_26475,N_25455,N_25410);
nor U26476 (N_26476,N_25535,N_24396);
and U26477 (N_26477,N_25389,N_24438);
or U26478 (N_26478,N_24118,N_25165);
xor U26479 (N_26479,N_24293,N_25816);
xnor U26480 (N_26480,N_25228,N_24531);
nand U26481 (N_26481,N_24884,N_24535);
xnor U26482 (N_26482,N_24228,N_25070);
nand U26483 (N_26483,N_24269,N_25626);
and U26484 (N_26484,N_24564,N_25268);
nor U26485 (N_26485,N_25123,N_25925);
nand U26486 (N_26486,N_24544,N_25295);
and U26487 (N_26487,N_24279,N_24446);
nand U26488 (N_26488,N_24093,N_24511);
and U26489 (N_26489,N_24073,N_24110);
nand U26490 (N_26490,N_25641,N_25129);
nand U26491 (N_26491,N_24702,N_25532);
nor U26492 (N_26492,N_24233,N_25130);
nor U26493 (N_26493,N_25960,N_25546);
nand U26494 (N_26494,N_24448,N_24005);
or U26495 (N_26495,N_25144,N_24008);
nor U26496 (N_26496,N_24893,N_24637);
and U26497 (N_26497,N_24620,N_24542);
xor U26498 (N_26498,N_24516,N_24191);
xnor U26499 (N_26499,N_25194,N_24303);
nor U26500 (N_26500,N_25050,N_24937);
and U26501 (N_26501,N_25710,N_25927);
nor U26502 (N_26502,N_24636,N_25411);
nor U26503 (N_26503,N_25445,N_25703);
nand U26504 (N_26504,N_25431,N_24373);
nand U26505 (N_26505,N_25582,N_24560);
nor U26506 (N_26506,N_25721,N_25500);
and U26507 (N_26507,N_25709,N_25518);
nand U26508 (N_26508,N_24793,N_24593);
and U26509 (N_26509,N_24755,N_25708);
nand U26510 (N_26510,N_24439,N_25941);
nor U26511 (N_26511,N_24756,N_24119);
nand U26512 (N_26512,N_25807,N_24743);
nor U26513 (N_26513,N_24890,N_25021);
and U26514 (N_26514,N_24049,N_25259);
or U26515 (N_26515,N_24969,N_25596);
nand U26516 (N_26516,N_25969,N_24044);
xnor U26517 (N_26517,N_24750,N_25799);
nor U26518 (N_26518,N_25577,N_24066);
nor U26519 (N_26519,N_25592,N_24237);
or U26520 (N_26520,N_25977,N_25630);
or U26521 (N_26521,N_25032,N_24190);
xor U26522 (N_26522,N_25429,N_24325);
or U26523 (N_26523,N_25267,N_25890);
xor U26524 (N_26524,N_24365,N_24571);
xor U26525 (N_26525,N_24835,N_24952);
nor U26526 (N_26526,N_24953,N_24421);
xor U26527 (N_26527,N_24393,N_24128);
xnor U26528 (N_26528,N_24854,N_25667);
nand U26529 (N_26529,N_25343,N_25568);
xnor U26530 (N_26530,N_25944,N_25224);
nand U26531 (N_26531,N_24397,N_25627);
and U26532 (N_26532,N_25618,N_24306);
nor U26533 (N_26533,N_25018,N_25623);
xnor U26534 (N_26534,N_25307,N_24477);
nor U26535 (N_26535,N_24485,N_25439);
and U26536 (N_26536,N_24817,N_25451);
nor U26537 (N_26537,N_25484,N_24137);
or U26538 (N_26538,N_24982,N_24061);
nor U26539 (N_26539,N_24341,N_25132);
nor U26540 (N_26540,N_24552,N_25112);
or U26541 (N_26541,N_24882,N_25013);
or U26542 (N_26542,N_24567,N_25488);
nor U26543 (N_26543,N_24818,N_25838);
nor U26544 (N_26544,N_24581,N_25063);
and U26545 (N_26545,N_25052,N_25346);
nand U26546 (N_26546,N_24070,N_24860);
nand U26547 (N_26547,N_24458,N_25275);
and U26548 (N_26548,N_25585,N_24472);
nor U26549 (N_26549,N_24796,N_25495);
or U26550 (N_26550,N_25153,N_24613);
nor U26551 (N_26551,N_25395,N_24483);
nor U26552 (N_26552,N_25951,N_25474);
nand U26553 (N_26553,N_25846,N_25507);
nand U26554 (N_26554,N_24194,N_24360);
nor U26555 (N_26555,N_24205,N_25007);
nor U26556 (N_26556,N_24410,N_24868);
xor U26557 (N_26557,N_24420,N_24527);
or U26558 (N_26558,N_25134,N_25012);
or U26559 (N_26559,N_24258,N_25991);
and U26560 (N_26560,N_24518,N_25148);
xnor U26561 (N_26561,N_24339,N_24941);
or U26562 (N_26562,N_24610,N_24034);
or U26563 (N_26563,N_24152,N_24234);
nand U26564 (N_26564,N_24259,N_25038);
nand U26565 (N_26565,N_24985,N_24009);
xnor U26566 (N_26566,N_25902,N_25109);
or U26567 (N_26567,N_25885,N_25625);
xnor U26568 (N_26568,N_24605,N_25852);
and U26569 (N_26569,N_25117,N_25617);
nand U26570 (N_26570,N_25205,N_24824);
nand U26571 (N_26571,N_24679,N_24594);
xor U26572 (N_26572,N_25309,N_25877);
and U26573 (N_26573,N_24151,N_24157);
or U26574 (N_26574,N_25771,N_25329);
nand U26575 (N_26575,N_24960,N_25188);
and U26576 (N_26576,N_25581,N_25650);
nand U26577 (N_26577,N_25967,N_25212);
and U26578 (N_26578,N_25405,N_24845);
xnor U26579 (N_26579,N_24609,N_24026);
and U26580 (N_26580,N_25607,N_25649);
xnor U26581 (N_26581,N_24989,N_24859);
nor U26582 (N_26582,N_24097,N_25542);
nor U26583 (N_26583,N_25874,N_25341);
nor U26584 (N_26584,N_24204,N_25360);
nor U26585 (N_26585,N_24263,N_25423);
or U26586 (N_26586,N_25113,N_25099);
nand U26587 (N_26587,N_25975,N_25265);
nand U26588 (N_26588,N_24130,N_25501);
and U26589 (N_26589,N_25722,N_25003);
xnor U26590 (N_26590,N_24146,N_24906);
or U26591 (N_26591,N_25124,N_25262);
or U26592 (N_26592,N_25491,N_24809);
or U26593 (N_26593,N_24842,N_24920);
nor U26594 (N_26594,N_25727,N_24220);
xnor U26595 (N_26595,N_24659,N_24905);
and U26596 (N_26596,N_24903,N_24680);
nor U26597 (N_26597,N_25665,N_24878);
xor U26598 (N_26598,N_25856,N_25835);
nand U26599 (N_26599,N_25393,N_24847);
nand U26600 (N_26600,N_24016,N_25509);
nand U26601 (N_26601,N_24069,N_25558);
and U26602 (N_26602,N_25082,N_25900);
or U26603 (N_26603,N_25758,N_24464);
nor U26604 (N_26604,N_25419,N_24992);
xor U26605 (N_26605,N_24025,N_25251);
xnor U26606 (N_26606,N_24315,N_25642);
or U26607 (N_26607,N_25033,N_24836);
xnor U26608 (N_26608,N_25520,N_24931);
or U26609 (N_26609,N_24100,N_24028);
or U26610 (N_26610,N_25526,N_25364);
nand U26611 (N_26611,N_24122,N_25606);
nand U26612 (N_26612,N_24231,N_24811);
nor U26613 (N_26613,N_25845,N_25800);
and U26614 (N_26614,N_25652,N_24650);
xor U26615 (N_26615,N_24742,N_24058);
and U26616 (N_26616,N_25071,N_25932);
and U26617 (N_26617,N_25290,N_25884);
xor U26618 (N_26618,N_24246,N_25935);
xnor U26619 (N_26619,N_25695,N_24528);
nor U26620 (N_26620,N_24640,N_24035);
and U26621 (N_26621,N_25680,N_24573);
xor U26622 (N_26622,N_25209,N_25512);
and U26623 (N_26623,N_25106,N_25226);
xnor U26624 (N_26624,N_24445,N_24971);
and U26625 (N_26625,N_25912,N_24918);
nand U26626 (N_26626,N_25387,N_24324);
or U26627 (N_26627,N_25983,N_25724);
nor U26628 (N_26628,N_25916,N_24226);
or U26629 (N_26629,N_25506,N_24651);
xor U26630 (N_26630,N_25810,N_25742);
nand U26631 (N_26631,N_24189,N_24720);
xnor U26632 (N_26632,N_25550,N_24216);
nor U26633 (N_26633,N_25471,N_24276);
or U26634 (N_26634,N_25645,N_24726);
nand U26635 (N_26635,N_24449,N_24327);
nand U26636 (N_26636,N_24366,N_24375);
nand U26637 (N_26637,N_25673,N_24082);
nor U26638 (N_26638,N_24075,N_25566);
nor U26639 (N_26639,N_24966,N_25768);
nand U26640 (N_26640,N_25339,N_25296);
and U26641 (N_26641,N_24786,N_24419);
nor U26642 (N_26642,N_24282,N_24252);
xnor U26643 (N_26643,N_24883,N_25412);
and U26644 (N_26644,N_25685,N_24261);
nor U26645 (N_26645,N_24795,N_24489);
nand U26646 (N_26646,N_24673,N_24652);
and U26647 (N_26647,N_25947,N_25039);
nor U26648 (N_26648,N_25547,N_25644);
and U26649 (N_26649,N_24133,N_24875);
and U26650 (N_26650,N_24170,N_25955);
or U26651 (N_26651,N_24923,N_25702);
and U26652 (N_26652,N_24799,N_24024);
and U26653 (N_26653,N_24965,N_25731);
xor U26654 (N_26654,N_24927,N_25971);
and U26655 (N_26655,N_25185,N_25361);
or U26656 (N_26656,N_25732,N_24995);
nor U26657 (N_26657,N_25376,N_24808);
and U26658 (N_26658,N_24617,N_25166);
nand U26659 (N_26659,N_24131,N_25694);
or U26660 (N_26660,N_24166,N_24088);
nor U26661 (N_26661,N_24729,N_25348);
nand U26662 (N_26662,N_25815,N_25894);
nor U26663 (N_26663,N_24358,N_25683);
and U26664 (N_26664,N_25371,N_25064);
or U26665 (N_26665,N_24503,N_24846);
nor U26666 (N_26666,N_25950,N_24408);
nor U26667 (N_26667,N_25183,N_24705);
nor U26668 (N_26668,N_25163,N_25554);
xor U26669 (N_26669,N_24467,N_25805);
or U26670 (N_26670,N_25288,N_25229);
nand U26671 (N_26671,N_24565,N_25263);
nor U26672 (N_26672,N_25841,N_25757);
or U26673 (N_26673,N_24820,N_25340);
nand U26674 (N_26674,N_25584,N_24381);
xnor U26675 (N_26675,N_24426,N_25922);
or U26676 (N_26676,N_25481,N_24945);
xnor U26677 (N_26677,N_24657,N_25893);
nand U26678 (N_26678,N_24430,N_24887);
and U26679 (N_26679,N_24994,N_25861);
xor U26680 (N_26680,N_25662,N_24724);
nor U26681 (N_26681,N_24561,N_25115);
or U26682 (N_26682,N_25088,N_25470);
or U26683 (N_26683,N_25690,N_25837);
or U26684 (N_26684,N_25094,N_25875);
and U26685 (N_26685,N_24677,N_25595);
nand U26686 (N_26686,N_24335,N_24424);
xnor U26687 (N_26687,N_25516,N_24328);
xnor U26688 (N_26688,N_24586,N_25517);
and U26689 (N_26689,N_24629,N_25637);
and U26690 (N_26690,N_25221,N_25321);
or U26691 (N_26691,N_24623,N_25741);
xor U26692 (N_26692,N_25513,N_25918);
nand U26693 (N_26693,N_24372,N_24183);
or U26694 (N_26694,N_24139,N_24973);
and U26695 (N_26695,N_24219,N_24400);
or U26696 (N_26696,N_24078,N_25452);
nand U26697 (N_26697,N_24405,N_24919);
or U26698 (N_26698,N_25420,N_24255);
nand U26699 (N_26699,N_25062,N_24343);
and U26700 (N_26700,N_24758,N_25555);
or U26701 (N_26701,N_25801,N_24232);
nor U26702 (N_26702,N_24111,N_25848);
or U26703 (N_26703,N_25026,N_25009);
xnor U26704 (N_26704,N_25345,N_25192);
and U26705 (N_26705,N_24316,N_24914);
xor U26706 (N_26706,N_25041,N_25402);
and U26707 (N_26707,N_25014,N_25354);
and U26708 (N_26708,N_25324,N_24607);
nor U26709 (N_26709,N_24447,N_24895);
nor U26710 (N_26710,N_25152,N_24356);
nand U26711 (N_26711,N_25575,N_24411);
and U26712 (N_26712,N_25887,N_25565);
nor U26713 (N_26713,N_25693,N_25408);
nor U26714 (N_26714,N_25719,N_24450);
or U26715 (N_26715,N_24959,N_25549);
nand U26716 (N_26716,N_25381,N_24904);
nand U26717 (N_26717,N_24787,N_25282);
xnor U26718 (N_26718,N_24717,N_25850);
nor U26719 (N_26719,N_25146,N_25706);
xnor U26720 (N_26720,N_24570,N_24661);
and U26721 (N_26721,N_25037,N_24779);
nand U26722 (N_26722,N_25428,N_25666);
nand U26723 (N_26723,N_24416,N_24427);
nor U26724 (N_26724,N_24080,N_25754);
xnor U26725 (N_26725,N_24563,N_24602);
nand U26726 (N_26726,N_25670,N_25619);
or U26727 (N_26727,N_24746,N_25621);
or U26728 (N_26728,N_25235,N_24022);
xnor U26729 (N_26729,N_25934,N_25111);
or U26730 (N_26730,N_24672,N_25611);
nor U26731 (N_26731,N_24751,N_25744);
nand U26732 (N_26732,N_24147,N_25114);
nand U26733 (N_26733,N_24482,N_25459);
nor U26734 (N_26734,N_25791,N_25273);
or U26735 (N_26735,N_25392,N_24332);
and U26736 (N_26736,N_24533,N_24996);
nor U26737 (N_26737,N_24167,N_25544);
xor U26738 (N_26738,N_25534,N_24239);
nor U26739 (N_26739,N_24807,N_24409);
or U26740 (N_26740,N_25261,N_25266);
xnor U26741 (N_26741,N_25120,N_24029);
and U26742 (N_26742,N_24798,N_24521);
xor U26743 (N_26743,N_25923,N_25353);
xnor U26744 (N_26744,N_25087,N_24032);
and U26745 (N_26745,N_24718,N_25090);
and U26746 (N_26746,N_25435,N_24997);
and U26747 (N_26747,N_25444,N_24529);
and U26748 (N_26748,N_25223,N_25897);
nand U26749 (N_26749,N_25989,N_25274);
and U26750 (N_26750,N_25015,N_24892);
nor U26751 (N_26751,N_25293,N_25356);
xor U26752 (N_26752,N_24921,N_24851);
and U26753 (N_26753,N_25628,N_24536);
nor U26754 (N_26754,N_25436,N_25531);
or U26755 (N_26755,N_24880,N_24019);
xor U26756 (N_26756,N_25747,N_24302);
xor U26757 (N_26757,N_24778,N_25792);
xor U26758 (N_26758,N_25493,N_24488);
and U26759 (N_26759,N_24566,N_25985);
nor U26760 (N_26760,N_25173,N_24202);
and U26761 (N_26761,N_24064,N_25379);
and U26762 (N_26762,N_25073,N_25521);
xnor U26763 (N_26763,N_24767,N_24178);
or U26764 (N_26764,N_24062,N_25964);
or U26765 (N_26765,N_25443,N_24115);
xor U26766 (N_26766,N_24031,N_24330);
xor U26767 (N_26767,N_25605,N_24759);
and U26768 (N_26768,N_24715,N_24342);
xnor U26769 (N_26769,N_25178,N_25374);
nor U26770 (N_26770,N_25756,N_24020);
nor U26771 (N_26771,N_24740,N_24978);
nor U26772 (N_26772,N_25485,N_25909);
nor U26773 (N_26773,N_24588,N_24962);
or U26774 (N_26774,N_25463,N_25269);
nor U26775 (N_26775,N_24520,N_25933);
xnor U26776 (N_26776,N_24891,N_24394);
nand U26777 (N_26777,N_25655,N_25701);
nand U26778 (N_26778,N_25276,N_25774);
or U26779 (N_26779,N_25180,N_25949);
and U26780 (N_26780,N_24414,N_24587);
nand U26781 (N_26781,N_24264,N_25151);
or U26782 (N_26782,N_25390,N_24121);
nand U26783 (N_26783,N_24852,N_25755);
nand U26784 (N_26784,N_25250,N_24422);
nand U26785 (N_26785,N_25434,N_25430);
nand U26786 (N_26786,N_24579,N_24936);
nand U26787 (N_26787,N_24753,N_25367);
nand U26788 (N_26788,N_24351,N_25734);
nor U26789 (N_26789,N_25243,N_24983);
nand U26790 (N_26790,N_25980,N_25515);
nand U26791 (N_26791,N_25674,N_24195);
nand U26792 (N_26792,N_25060,N_24744);
nor U26793 (N_26793,N_24627,N_24344);
xnor U26794 (N_26794,N_25357,N_25790);
and U26795 (N_26795,N_25342,N_25730);
and U26796 (N_26796,N_24413,N_24604);
xnor U26797 (N_26797,N_25305,N_24432);
or U26798 (N_26798,N_25065,N_24142);
nor U26799 (N_26799,N_24181,N_25368);
nor U26800 (N_26800,N_24086,N_24548);
and U26801 (N_26801,N_25385,N_24113);
xor U26802 (N_26802,N_24251,N_24980);
nor U26803 (N_26803,N_25522,N_24212);
or U26804 (N_26804,N_25351,N_24669);
nand U26805 (N_26805,N_25811,N_24116);
nand U26806 (N_26806,N_25311,N_24383);
and U26807 (N_26807,N_24434,N_25446);
and U26808 (N_26808,N_25085,N_25760);
or U26809 (N_26809,N_25880,N_25103);
xor U26810 (N_26810,N_25058,N_24986);
and U26811 (N_26811,N_25006,N_24247);
or U26812 (N_26812,N_24577,N_25081);
or U26813 (N_26813,N_24537,N_25579);
and U26814 (N_26814,N_25996,N_25511);
nand U26815 (N_26815,N_24591,N_24939);
nor U26816 (N_26816,N_24780,N_24599);
nand U26817 (N_26817,N_25456,N_25225);
xor U26818 (N_26818,N_25022,N_25728);
or U26819 (N_26819,N_24000,N_24127);
nor U26820 (N_26820,N_25246,N_24525);
nor U26821 (N_26821,N_25136,N_24172);
xor U26822 (N_26822,N_25976,N_24964);
nor U26823 (N_26823,N_24391,N_25181);
or U26824 (N_26824,N_24209,N_25158);
nand U26825 (N_26825,N_25589,N_25333);
or U26826 (N_26826,N_24401,N_24666);
or U26827 (N_26827,N_24569,N_24546);
and U26828 (N_26828,N_25919,N_24284);
and U26829 (N_26829,N_24855,N_25135);
nand U26830 (N_26830,N_24611,N_24877);
xor U26831 (N_26831,N_25004,N_25736);
nand U26832 (N_26832,N_25182,N_24173);
nor U26833 (N_26833,N_24441,N_24663);
nor U26834 (N_26834,N_24674,N_25697);
nor U26835 (N_26835,N_24451,N_25795);
nor U26836 (N_26836,N_24789,N_24708);
xor U26837 (N_26837,N_24431,N_25477);
nor U26838 (N_26838,N_25620,N_24865);
xor U26839 (N_26839,N_25784,N_25844);
nor U26840 (N_26840,N_25175,N_24540);
or U26841 (N_26841,N_24145,N_24889);
xor U26842 (N_26842,N_24090,N_25872);
nor U26843 (N_26843,N_25752,N_25264);
nor U26844 (N_26844,N_25089,N_25036);
and U26845 (N_26845,N_24412,N_25682);
nand U26846 (N_26846,N_25237,N_25055);
or U26847 (N_26847,N_25049,N_24502);
or U26848 (N_26848,N_25963,N_25653);
xor U26849 (N_26849,N_24728,N_25802);
or U26850 (N_26850,N_24253,N_25808);
nand U26851 (N_26851,N_24956,N_25207);
nor U26852 (N_26852,N_25788,N_24164);
xnor U26853 (N_26853,N_24236,N_24321);
nor U26854 (N_26854,N_25141,N_25247);
and U26855 (N_26855,N_25399,N_24126);
xor U26856 (N_26856,N_24106,N_25010);
or U26857 (N_26857,N_25414,N_25490);
and U26858 (N_26858,N_25888,N_25541);
and U26859 (N_26859,N_24967,N_24625);
nor U26860 (N_26860,N_25571,N_25378);
xor U26861 (N_26861,N_24001,N_24723);
xnor U26862 (N_26862,N_24701,N_24241);
xnor U26863 (N_26863,N_25108,N_24158);
nand U26864 (N_26864,N_24156,N_25031);
xnor U26865 (N_26865,N_25404,N_24686);
xnor U26866 (N_26866,N_24298,N_25313);
nor U26867 (N_26867,N_25417,N_25896);
xor U26868 (N_26868,N_25140,N_24689);
or U26869 (N_26869,N_24182,N_24095);
xnor U26870 (N_26870,N_25475,N_25992);
nor U26871 (N_26871,N_24532,N_24404);
nand U26872 (N_26872,N_24829,N_24435);
nand U26873 (N_26873,N_24538,N_24072);
and U26874 (N_26874,N_25738,N_25814);
or U26875 (N_26875,N_25943,N_25859);
xor U26876 (N_26876,N_24790,N_25306);
or U26877 (N_26877,N_24948,N_25678);
nand U26878 (N_26878,N_24469,N_25285);
nor U26879 (N_26879,N_25966,N_24313);
or U26880 (N_26880,N_24299,N_24622);
xor U26881 (N_26881,N_25775,N_25466);
nand U26882 (N_26882,N_24988,N_25105);
nor U26883 (N_26883,N_24515,N_24949);
and U26884 (N_26884,N_24861,N_25990);
nor U26885 (N_26885,N_25294,N_24196);
xnor U26886 (N_26886,N_24694,N_25569);
or U26887 (N_26887,N_24711,N_24979);
nor U26888 (N_26888,N_24603,N_25505);
nor U26889 (N_26889,N_24947,N_24123);
or U26890 (N_26890,N_24826,N_25770);
and U26891 (N_26891,N_24722,N_24630);
and U26892 (N_26892,N_24930,N_24285);
or U26893 (N_26893,N_24318,N_24099);
or U26894 (N_26894,N_25629,N_25421);
xnor U26895 (N_26895,N_24731,N_25725);
nand U26896 (N_26896,N_25854,N_25170);
and U26897 (N_26897,N_25300,N_24999);
nor U26898 (N_26898,N_25527,N_24984);
and U26899 (N_26899,N_25588,N_25712);
nor U26900 (N_26900,N_25127,N_24699);
nor U26901 (N_26901,N_25572,N_25279);
nor U26902 (N_26902,N_25469,N_24014);
and U26903 (N_26903,N_24399,N_25331);
nand U26904 (N_26904,N_24319,N_25762);
nand U26905 (N_26905,N_25142,N_25552);
nor U26906 (N_26906,N_25323,N_25442);
and U26907 (N_26907,N_25187,N_25011);
nand U26908 (N_26908,N_24206,N_25497);
nor U26909 (N_26909,N_25016,N_24433);
xnor U26910 (N_26910,N_24899,N_24935);
nor U26911 (N_26911,N_24703,N_24512);
and U26912 (N_26912,N_24107,N_24368);
nand U26913 (N_26913,N_24870,N_25543);
and U26914 (N_26914,N_25789,N_24554);
xnor U26915 (N_26915,N_24782,N_24774);
xor U26916 (N_26916,N_25583,N_24120);
nor U26917 (N_26917,N_25656,N_25867);
and U26918 (N_26918,N_24549,N_25028);
nand U26919 (N_26919,N_25564,N_24287);
xor U26920 (N_26920,N_24201,N_24169);
and U26921 (N_26921,N_24369,N_25610);
and U26922 (N_26922,N_24911,N_25745);
nand U26923 (N_26923,N_25133,N_25840);
xor U26924 (N_26924,N_24197,N_25553);
xor U26925 (N_26925,N_24108,N_25573);
or U26926 (N_26926,N_25352,N_24951);
xor U26927 (N_26927,N_24639,N_24738);
and U26928 (N_26928,N_25510,N_25676);
nand U26929 (N_26929,N_25286,N_24776);
nand U26930 (N_26930,N_25494,N_24812);
xor U26931 (N_26931,N_25749,N_25448);
and U26932 (N_26932,N_24821,N_25380);
nor U26933 (N_26933,N_24087,N_24207);
and U26934 (N_26934,N_24747,N_25959);
nand U26935 (N_26935,N_24848,N_24387);
xor U26936 (N_26936,N_25384,N_25911);
nand U26937 (N_26937,N_25441,N_24013);
nand U26938 (N_26938,N_24377,N_24757);
nor U26939 (N_26939,N_25234,N_25821);
xor U26940 (N_26940,N_25271,N_24479);
or U26941 (N_26941,N_24595,N_24305);
or U26942 (N_26942,N_24240,N_24199);
or U26943 (N_26943,N_25700,N_25017);
or U26944 (N_26944,N_24091,N_24048);
nand U26945 (N_26945,N_24105,N_25398);
nor U26946 (N_26946,N_24562,N_24033);
nand U26947 (N_26947,N_25184,N_25707);
and U26948 (N_26948,N_25794,N_24295);
xor U26949 (N_26949,N_25593,N_25272);
and U26950 (N_26950,N_24063,N_24281);
nand U26951 (N_26951,N_25687,N_24839);
xor U26952 (N_26952,N_25222,N_24858);
or U26953 (N_26953,N_24785,N_24056);
xor U26954 (N_26954,N_25319,N_24716);
xnor U26955 (N_26955,N_25819,N_24748);
xnor U26956 (N_26956,N_25820,N_25907);
or U26957 (N_26957,N_25698,N_25806);
and U26958 (N_26958,N_24017,N_25570);
nand U26959 (N_26959,N_25668,N_25851);
nand U26960 (N_26960,N_25766,N_25236);
and U26961 (N_26961,N_25386,N_25870);
and U26962 (N_26962,N_25672,N_25053);
nor U26963 (N_26963,N_25483,N_25692);
and U26964 (N_26964,N_25828,N_24874);
and U26965 (N_26965,N_25308,N_25230);
nor U26966 (N_26966,N_25383,N_25172);
xor U26967 (N_26967,N_24775,N_24837);
nor U26968 (N_26968,N_24294,N_24454);
nand U26969 (N_26969,N_25982,N_25409);
nor U26970 (N_26970,N_25218,N_25639);
nand U26971 (N_26971,N_25066,N_25190);
nor U26972 (N_26972,N_25315,N_24362);
nand U26973 (N_26973,N_24245,N_24981);
xnor U26974 (N_26974,N_25056,N_25537);
xor U26975 (N_26975,N_24322,N_25373);
nor U26976 (N_26976,N_24885,N_25945);
or U26977 (N_26977,N_24224,N_24794);
nand U26978 (N_26978,N_25586,N_25930);
nor U26979 (N_26979,N_25464,N_25426);
and U26980 (N_26980,N_24621,N_25640);
xor U26981 (N_26981,N_24290,N_24143);
or U26982 (N_26982,N_25899,N_24223);
xor U26983 (N_26983,N_25962,N_25508);
nor U26984 (N_26984,N_24678,N_24418);
nand U26985 (N_26985,N_24460,N_25104);
xor U26986 (N_26986,N_25126,N_25217);
nor U26987 (N_26987,N_24363,N_25075);
xor U26988 (N_26988,N_24068,N_24030);
xor U26989 (N_26989,N_24916,N_25779);
nand U26990 (N_26990,N_25318,N_25330);
xor U26991 (N_26991,N_25239,N_24901);
nand U26992 (N_26992,N_25024,N_25210);
or U26993 (N_26993,N_24493,N_25679);
nand U26994 (N_26994,N_25382,N_24576);
and U26995 (N_26995,N_24054,N_25936);
xnor U26996 (N_26996,N_25283,N_24805);
xor U26997 (N_26997,N_24361,N_24417);
or U26998 (N_26998,N_25231,N_25978);
and U26999 (N_26999,N_25600,N_24038);
or U27000 (N_27000,N_25163,N_25038);
and U27001 (N_27001,N_25816,N_24415);
xnor U27002 (N_27002,N_25247,N_24732);
nand U27003 (N_27003,N_24265,N_24006);
and U27004 (N_27004,N_24347,N_25653);
and U27005 (N_27005,N_25699,N_24657);
or U27006 (N_27006,N_24169,N_24785);
nand U27007 (N_27007,N_24578,N_25375);
nand U27008 (N_27008,N_24319,N_24920);
nor U27009 (N_27009,N_24940,N_24226);
nand U27010 (N_27010,N_25288,N_25904);
or U27011 (N_27011,N_25342,N_25522);
or U27012 (N_27012,N_24995,N_25565);
or U27013 (N_27013,N_25608,N_25328);
nor U27014 (N_27014,N_25876,N_24697);
or U27015 (N_27015,N_24013,N_24334);
nor U27016 (N_27016,N_25567,N_24055);
and U27017 (N_27017,N_25084,N_25779);
nor U27018 (N_27018,N_24516,N_25488);
and U27019 (N_27019,N_24228,N_24110);
nand U27020 (N_27020,N_25035,N_25021);
nor U27021 (N_27021,N_24653,N_25806);
xor U27022 (N_27022,N_25379,N_24858);
nor U27023 (N_27023,N_25625,N_25069);
nand U27024 (N_27024,N_25389,N_24876);
or U27025 (N_27025,N_25864,N_24702);
xor U27026 (N_27026,N_24974,N_24952);
nor U27027 (N_27027,N_24076,N_25736);
xor U27028 (N_27028,N_24395,N_25648);
and U27029 (N_27029,N_24136,N_24389);
xnor U27030 (N_27030,N_24206,N_25535);
and U27031 (N_27031,N_25575,N_24298);
or U27032 (N_27032,N_24004,N_24988);
nor U27033 (N_27033,N_24842,N_25786);
xnor U27034 (N_27034,N_24013,N_24126);
and U27035 (N_27035,N_24292,N_24159);
nand U27036 (N_27036,N_24823,N_24957);
or U27037 (N_27037,N_25491,N_25333);
nor U27038 (N_27038,N_24846,N_24769);
and U27039 (N_27039,N_24459,N_25935);
nand U27040 (N_27040,N_25304,N_24739);
and U27041 (N_27041,N_25958,N_25423);
nor U27042 (N_27042,N_25160,N_25614);
and U27043 (N_27043,N_24843,N_25095);
xor U27044 (N_27044,N_25197,N_24962);
xor U27045 (N_27045,N_24229,N_24516);
and U27046 (N_27046,N_25131,N_24973);
or U27047 (N_27047,N_24487,N_24134);
and U27048 (N_27048,N_24737,N_24842);
nor U27049 (N_27049,N_25770,N_24927);
and U27050 (N_27050,N_25422,N_25092);
and U27051 (N_27051,N_24191,N_25342);
or U27052 (N_27052,N_25812,N_25008);
xnor U27053 (N_27053,N_25927,N_25445);
nor U27054 (N_27054,N_24734,N_25831);
or U27055 (N_27055,N_24207,N_25565);
and U27056 (N_27056,N_25241,N_25505);
and U27057 (N_27057,N_24793,N_24051);
and U27058 (N_27058,N_25761,N_24837);
nor U27059 (N_27059,N_24543,N_25369);
nand U27060 (N_27060,N_25971,N_25513);
and U27061 (N_27061,N_25968,N_24121);
and U27062 (N_27062,N_25953,N_24351);
nand U27063 (N_27063,N_25544,N_25075);
nand U27064 (N_27064,N_25101,N_24009);
or U27065 (N_27065,N_25178,N_24274);
or U27066 (N_27066,N_24744,N_24539);
nand U27067 (N_27067,N_25010,N_24393);
or U27068 (N_27068,N_25252,N_24469);
xnor U27069 (N_27069,N_25910,N_25501);
and U27070 (N_27070,N_24280,N_24533);
xor U27071 (N_27071,N_25810,N_25303);
and U27072 (N_27072,N_24132,N_24654);
xor U27073 (N_27073,N_25961,N_24520);
or U27074 (N_27074,N_24755,N_24711);
and U27075 (N_27075,N_25581,N_24431);
xor U27076 (N_27076,N_25126,N_25574);
nor U27077 (N_27077,N_25244,N_24355);
and U27078 (N_27078,N_25365,N_25927);
nand U27079 (N_27079,N_25291,N_25145);
nor U27080 (N_27080,N_25192,N_25489);
and U27081 (N_27081,N_25974,N_25464);
xor U27082 (N_27082,N_24707,N_24817);
nand U27083 (N_27083,N_24454,N_25127);
nor U27084 (N_27084,N_24324,N_25550);
and U27085 (N_27085,N_24743,N_25737);
or U27086 (N_27086,N_24177,N_24531);
xor U27087 (N_27087,N_24606,N_25753);
or U27088 (N_27088,N_24476,N_25439);
and U27089 (N_27089,N_25522,N_25338);
nand U27090 (N_27090,N_25763,N_24558);
nand U27091 (N_27091,N_24973,N_24676);
xnor U27092 (N_27092,N_25972,N_24535);
nor U27093 (N_27093,N_25166,N_24598);
or U27094 (N_27094,N_25440,N_25027);
nor U27095 (N_27095,N_25432,N_24531);
xor U27096 (N_27096,N_24242,N_24862);
nor U27097 (N_27097,N_24856,N_25906);
xor U27098 (N_27098,N_25270,N_24424);
and U27099 (N_27099,N_24179,N_24156);
xnor U27100 (N_27100,N_24108,N_25453);
nand U27101 (N_27101,N_25178,N_25791);
or U27102 (N_27102,N_24477,N_25993);
and U27103 (N_27103,N_25323,N_24717);
or U27104 (N_27104,N_25575,N_25043);
nor U27105 (N_27105,N_25799,N_24813);
xnor U27106 (N_27106,N_25509,N_25477);
and U27107 (N_27107,N_24554,N_24915);
and U27108 (N_27108,N_24502,N_25675);
and U27109 (N_27109,N_24712,N_24939);
nand U27110 (N_27110,N_24407,N_24006);
or U27111 (N_27111,N_24447,N_24765);
nand U27112 (N_27112,N_25174,N_24601);
and U27113 (N_27113,N_24774,N_24708);
xor U27114 (N_27114,N_25789,N_25057);
and U27115 (N_27115,N_25259,N_25505);
nand U27116 (N_27116,N_25841,N_25131);
and U27117 (N_27117,N_25031,N_25490);
xnor U27118 (N_27118,N_24492,N_24425);
and U27119 (N_27119,N_25392,N_24598);
and U27120 (N_27120,N_24529,N_24764);
xnor U27121 (N_27121,N_25995,N_24371);
nand U27122 (N_27122,N_24367,N_25214);
nor U27123 (N_27123,N_24596,N_24336);
nand U27124 (N_27124,N_25225,N_25738);
nand U27125 (N_27125,N_25024,N_24526);
nor U27126 (N_27126,N_24050,N_24065);
and U27127 (N_27127,N_25215,N_25344);
and U27128 (N_27128,N_24969,N_25977);
nand U27129 (N_27129,N_24760,N_24790);
xor U27130 (N_27130,N_24861,N_25026);
nor U27131 (N_27131,N_24637,N_25399);
and U27132 (N_27132,N_24847,N_25007);
nor U27133 (N_27133,N_24811,N_24144);
and U27134 (N_27134,N_24325,N_24788);
nand U27135 (N_27135,N_24148,N_24782);
or U27136 (N_27136,N_25498,N_25469);
xor U27137 (N_27137,N_24864,N_25538);
or U27138 (N_27138,N_24913,N_24079);
and U27139 (N_27139,N_24890,N_25896);
nor U27140 (N_27140,N_25147,N_25347);
and U27141 (N_27141,N_24526,N_25502);
nor U27142 (N_27142,N_25907,N_24445);
nor U27143 (N_27143,N_24986,N_25490);
and U27144 (N_27144,N_24282,N_25724);
nor U27145 (N_27145,N_25033,N_25093);
xor U27146 (N_27146,N_24191,N_25015);
xor U27147 (N_27147,N_25880,N_25373);
and U27148 (N_27148,N_24542,N_25002);
xnor U27149 (N_27149,N_25302,N_25468);
or U27150 (N_27150,N_25637,N_24344);
and U27151 (N_27151,N_24150,N_25783);
and U27152 (N_27152,N_25281,N_25868);
xnor U27153 (N_27153,N_24249,N_25420);
nand U27154 (N_27154,N_24533,N_25130);
and U27155 (N_27155,N_24700,N_25502);
or U27156 (N_27156,N_24152,N_25511);
and U27157 (N_27157,N_24412,N_24913);
xor U27158 (N_27158,N_24075,N_25056);
nor U27159 (N_27159,N_25082,N_25619);
and U27160 (N_27160,N_24741,N_24833);
and U27161 (N_27161,N_24532,N_25664);
nand U27162 (N_27162,N_24896,N_24791);
nand U27163 (N_27163,N_24758,N_24107);
nand U27164 (N_27164,N_24086,N_24495);
nand U27165 (N_27165,N_24363,N_24340);
and U27166 (N_27166,N_25276,N_25841);
or U27167 (N_27167,N_25797,N_25167);
nand U27168 (N_27168,N_24556,N_24940);
xnor U27169 (N_27169,N_25516,N_25860);
nor U27170 (N_27170,N_24146,N_25923);
nand U27171 (N_27171,N_25759,N_24425);
and U27172 (N_27172,N_25659,N_25245);
and U27173 (N_27173,N_25065,N_24412);
xnor U27174 (N_27174,N_24820,N_24965);
and U27175 (N_27175,N_24651,N_24832);
or U27176 (N_27176,N_25943,N_25476);
nor U27177 (N_27177,N_25402,N_25892);
nand U27178 (N_27178,N_25882,N_25273);
xnor U27179 (N_27179,N_24529,N_24284);
and U27180 (N_27180,N_24136,N_25662);
and U27181 (N_27181,N_24196,N_24568);
or U27182 (N_27182,N_25175,N_24148);
nand U27183 (N_27183,N_25056,N_25953);
nand U27184 (N_27184,N_25444,N_24484);
nand U27185 (N_27185,N_24306,N_25880);
or U27186 (N_27186,N_24221,N_25728);
nand U27187 (N_27187,N_25811,N_25419);
nand U27188 (N_27188,N_25866,N_24959);
or U27189 (N_27189,N_24792,N_25174);
nor U27190 (N_27190,N_24183,N_25262);
nor U27191 (N_27191,N_25104,N_25321);
and U27192 (N_27192,N_25649,N_24806);
or U27193 (N_27193,N_24436,N_25166);
nand U27194 (N_27194,N_25986,N_25076);
and U27195 (N_27195,N_25044,N_24706);
and U27196 (N_27196,N_25679,N_24000);
or U27197 (N_27197,N_24969,N_24589);
xnor U27198 (N_27198,N_25351,N_25933);
and U27199 (N_27199,N_24692,N_24668);
nor U27200 (N_27200,N_25442,N_24886);
and U27201 (N_27201,N_25718,N_24968);
nor U27202 (N_27202,N_25363,N_25015);
nor U27203 (N_27203,N_25090,N_25780);
nor U27204 (N_27204,N_25890,N_25981);
nand U27205 (N_27205,N_24261,N_24139);
nand U27206 (N_27206,N_25535,N_24608);
or U27207 (N_27207,N_24198,N_25751);
nand U27208 (N_27208,N_24638,N_24303);
or U27209 (N_27209,N_24310,N_25630);
and U27210 (N_27210,N_24197,N_24620);
or U27211 (N_27211,N_25120,N_24055);
and U27212 (N_27212,N_25590,N_25909);
nand U27213 (N_27213,N_24065,N_24668);
or U27214 (N_27214,N_24607,N_25915);
or U27215 (N_27215,N_24348,N_24983);
xnor U27216 (N_27216,N_25710,N_24461);
and U27217 (N_27217,N_25560,N_25612);
xor U27218 (N_27218,N_25822,N_24834);
nor U27219 (N_27219,N_25473,N_24987);
nand U27220 (N_27220,N_25632,N_25968);
nor U27221 (N_27221,N_25057,N_24086);
xnor U27222 (N_27222,N_25548,N_24736);
nand U27223 (N_27223,N_24233,N_24174);
nor U27224 (N_27224,N_24336,N_25811);
nor U27225 (N_27225,N_25587,N_25350);
and U27226 (N_27226,N_25797,N_24883);
nor U27227 (N_27227,N_24586,N_24481);
nand U27228 (N_27228,N_25494,N_24331);
or U27229 (N_27229,N_25747,N_25877);
nor U27230 (N_27230,N_25649,N_25442);
nor U27231 (N_27231,N_24801,N_24677);
or U27232 (N_27232,N_24548,N_25107);
nor U27233 (N_27233,N_24385,N_25854);
or U27234 (N_27234,N_24436,N_24654);
nor U27235 (N_27235,N_25371,N_25803);
nor U27236 (N_27236,N_24996,N_25426);
nand U27237 (N_27237,N_24973,N_25865);
nor U27238 (N_27238,N_25163,N_25120);
xor U27239 (N_27239,N_24021,N_24787);
xor U27240 (N_27240,N_25098,N_25170);
xor U27241 (N_27241,N_25096,N_24653);
xnor U27242 (N_27242,N_25957,N_24070);
or U27243 (N_27243,N_24397,N_24217);
xnor U27244 (N_27244,N_25630,N_24216);
xnor U27245 (N_27245,N_25092,N_24084);
xnor U27246 (N_27246,N_25965,N_25895);
and U27247 (N_27247,N_24607,N_25041);
or U27248 (N_27248,N_25236,N_24764);
nand U27249 (N_27249,N_24220,N_25680);
and U27250 (N_27250,N_24806,N_24022);
nand U27251 (N_27251,N_24544,N_25219);
nor U27252 (N_27252,N_25834,N_25943);
xor U27253 (N_27253,N_24549,N_24000);
and U27254 (N_27254,N_25627,N_24579);
and U27255 (N_27255,N_24918,N_24475);
nand U27256 (N_27256,N_25770,N_24985);
xor U27257 (N_27257,N_25832,N_25480);
nor U27258 (N_27258,N_24550,N_25982);
nand U27259 (N_27259,N_25825,N_25167);
xnor U27260 (N_27260,N_24641,N_24168);
nor U27261 (N_27261,N_25698,N_25026);
or U27262 (N_27262,N_25350,N_24521);
xor U27263 (N_27263,N_25854,N_25781);
or U27264 (N_27264,N_24008,N_24480);
xor U27265 (N_27265,N_24276,N_24715);
xor U27266 (N_27266,N_25231,N_25737);
nand U27267 (N_27267,N_25776,N_24739);
or U27268 (N_27268,N_24083,N_25381);
xnor U27269 (N_27269,N_25863,N_25305);
xnor U27270 (N_27270,N_25833,N_25358);
or U27271 (N_27271,N_25347,N_24740);
nand U27272 (N_27272,N_24774,N_24476);
or U27273 (N_27273,N_25038,N_24244);
nor U27274 (N_27274,N_24902,N_24320);
and U27275 (N_27275,N_24315,N_25837);
xor U27276 (N_27276,N_24426,N_24518);
nor U27277 (N_27277,N_25693,N_24690);
xnor U27278 (N_27278,N_24039,N_25809);
nor U27279 (N_27279,N_24064,N_25983);
xor U27280 (N_27280,N_24629,N_25308);
nand U27281 (N_27281,N_24450,N_25250);
and U27282 (N_27282,N_25370,N_25130);
nand U27283 (N_27283,N_25572,N_24400);
nor U27284 (N_27284,N_25311,N_24773);
or U27285 (N_27285,N_24095,N_24508);
nand U27286 (N_27286,N_24225,N_25824);
or U27287 (N_27287,N_25549,N_25854);
nor U27288 (N_27288,N_24430,N_24917);
or U27289 (N_27289,N_24365,N_24190);
xor U27290 (N_27290,N_24291,N_24622);
and U27291 (N_27291,N_25294,N_24998);
and U27292 (N_27292,N_24483,N_25344);
and U27293 (N_27293,N_24679,N_24472);
xor U27294 (N_27294,N_25787,N_24837);
nor U27295 (N_27295,N_25854,N_24809);
or U27296 (N_27296,N_25161,N_24248);
xor U27297 (N_27297,N_24417,N_24614);
or U27298 (N_27298,N_24523,N_24373);
nand U27299 (N_27299,N_25855,N_24471);
xnor U27300 (N_27300,N_24275,N_25159);
nand U27301 (N_27301,N_25142,N_24664);
nand U27302 (N_27302,N_24745,N_25179);
or U27303 (N_27303,N_24836,N_24745);
nand U27304 (N_27304,N_25725,N_24008);
nor U27305 (N_27305,N_24790,N_24118);
nor U27306 (N_27306,N_25507,N_25467);
nor U27307 (N_27307,N_24642,N_25949);
nor U27308 (N_27308,N_25465,N_24570);
nor U27309 (N_27309,N_25224,N_25393);
or U27310 (N_27310,N_24612,N_24101);
or U27311 (N_27311,N_24885,N_25774);
nor U27312 (N_27312,N_24750,N_24968);
or U27313 (N_27313,N_24518,N_25726);
nor U27314 (N_27314,N_24204,N_25593);
or U27315 (N_27315,N_24976,N_25209);
xnor U27316 (N_27316,N_24596,N_25751);
or U27317 (N_27317,N_25477,N_25233);
nor U27318 (N_27318,N_24933,N_25421);
nand U27319 (N_27319,N_25736,N_24111);
nor U27320 (N_27320,N_24705,N_25645);
nor U27321 (N_27321,N_24512,N_24762);
xor U27322 (N_27322,N_24348,N_25392);
nand U27323 (N_27323,N_24633,N_25522);
xnor U27324 (N_27324,N_25980,N_25689);
nand U27325 (N_27325,N_24356,N_24699);
xnor U27326 (N_27326,N_25948,N_24901);
nand U27327 (N_27327,N_24350,N_24793);
and U27328 (N_27328,N_25673,N_25573);
nand U27329 (N_27329,N_25978,N_24212);
or U27330 (N_27330,N_24476,N_24507);
xnor U27331 (N_27331,N_25332,N_25993);
nor U27332 (N_27332,N_25692,N_25443);
nor U27333 (N_27333,N_25438,N_25406);
xor U27334 (N_27334,N_24764,N_24895);
or U27335 (N_27335,N_24614,N_25863);
or U27336 (N_27336,N_25922,N_25241);
nor U27337 (N_27337,N_24311,N_25874);
or U27338 (N_27338,N_24205,N_24975);
and U27339 (N_27339,N_25958,N_24811);
nand U27340 (N_27340,N_24426,N_25623);
and U27341 (N_27341,N_24414,N_25124);
nand U27342 (N_27342,N_24947,N_24816);
or U27343 (N_27343,N_25314,N_25957);
nand U27344 (N_27344,N_25215,N_25765);
and U27345 (N_27345,N_25839,N_25946);
or U27346 (N_27346,N_24334,N_24789);
nor U27347 (N_27347,N_25353,N_24480);
and U27348 (N_27348,N_24019,N_25472);
nand U27349 (N_27349,N_25898,N_24560);
xnor U27350 (N_27350,N_24035,N_25312);
nor U27351 (N_27351,N_25204,N_25043);
or U27352 (N_27352,N_25442,N_24297);
nor U27353 (N_27353,N_25308,N_25405);
and U27354 (N_27354,N_25785,N_24434);
nand U27355 (N_27355,N_25457,N_25090);
nand U27356 (N_27356,N_25050,N_25604);
xnor U27357 (N_27357,N_24279,N_24173);
and U27358 (N_27358,N_24870,N_25942);
nand U27359 (N_27359,N_24668,N_24665);
or U27360 (N_27360,N_24486,N_24434);
nor U27361 (N_27361,N_25934,N_25307);
nand U27362 (N_27362,N_24378,N_25799);
nor U27363 (N_27363,N_24652,N_24654);
or U27364 (N_27364,N_24368,N_25539);
nand U27365 (N_27365,N_25777,N_24541);
xor U27366 (N_27366,N_24444,N_25861);
and U27367 (N_27367,N_24436,N_24622);
nor U27368 (N_27368,N_24462,N_24995);
xor U27369 (N_27369,N_24112,N_24482);
and U27370 (N_27370,N_24757,N_24182);
nand U27371 (N_27371,N_25231,N_25243);
or U27372 (N_27372,N_25275,N_24877);
nand U27373 (N_27373,N_25795,N_25025);
nor U27374 (N_27374,N_25066,N_24729);
or U27375 (N_27375,N_24382,N_24519);
xor U27376 (N_27376,N_25919,N_25008);
nor U27377 (N_27377,N_25740,N_24675);
xnor U27378 (N_27378,N_25644,N_25515);
nor U27379 (N_27379,N_25751,N_25992);
nand U27380 (N_27380,N_24993,N_24615);
and U27381 (N_27381,N_25240,N_25491);
nor U27382 (N_27382,N_24558,N_25147);
nor U27383 (N_27383,N_25248,N_25016);
nor U27384 (N_27384,N_25610,N_25318);
or U27385 (N_27385,N_24646,N_24594);
xnor U27386 (N_27386,N_24257,N_25208);
and U27387 (N_27387,N_25147,N_25954);
and U27388 (N_27388,N_25544,N_24237);
xnor U27389 (N_27389,N_24933,N_24524);
or U27390 (N_27390,N_25005,N_25936);
nor U27391 (N_27391,N_25775,N_25705);
or U27392 (N_27392,N_24405,N_25797);
nor U27393 (N_27393,N_25782,N_24504);
or U27394 (N_27394,N_24639,N_24650);
or U27395 (N_27395,N_24243,N_24881);
nor U27396 (N_27396,N_24382,N_24354);
and U27397 (N_27397,N_25278,N_24534);
and U27398 (N_27398,N_24258,N_24869);
xor U27399 (N_27399,N_25677,N_25520);
and U27400 (N_27400,N_25180,N_24973);
and U27401 (N_27401,N_24072,N_24759);
nor U27402 (N_27402,N_24676,N_24864);
xor U27403 (N_27403,N_25368,N_24704);
and U27404 (N_27404,N_25858,N_24160);
nand U27405 (N_27405,N_25974,N_24758);
xor U27406 (N_27406,N_25825,N_24204);
and U27407 (N_27407,N_24533,N_25315);
nor U27408 (N_27408,N_24545,N_24014);
nand U27409 (N_27409,N_24223,N_25222);
nor U27410 (N_27410,N_25007,N_24216);
xnor U27411 (N_27411,N_25869,N_24302);
xor U27412 (N_27412,N_24234,N_24368);
or U27413 (N_27413,N_24697,N_24534);
xor U27414 (N_27414,N_25819,N_25551);
and U27415 (N_27415,N_25997,N_24631);
or U27416 (N_27416,N_25097,N_24399);
nand U27417 (N_27417,N_25822,N_24264);
and U27418 (N_27418,N_25386,N_25049);
nor U27419 (N_27419,N_25601,N_24365);
and U27420 (N_27420,N_25005,N_25990);
nand U27421 (N_27421,N_24105,N_25443);
nor U27422 (N_27422,N_25299,N_24452);
or U27423 (N_27423,N_24362,N_24100);
nor U27424 (N_27424,N_25652,N_25634);
and U27425 (N_27425,N_24198,N_25669);
nor U27426 (N_27426,N_24464,N_24635);
nand U27427 (N_27427,N_25658,N_25175);
and U27428 (N_27428,N_25194,N_24893);
nand U27429 (N_27429,N_25900,N_25643);
nor U27430 (N_27430,N_24101,N_25857);
xnor U27431 (N_27431,N_24925,N_24888);
and U27432 (N_27432,N_24177,N_25423);
nor U27433 (N_27433,N_25478,N_24925);
and U27434 (N_27434,N_24576,N_25537);
nand U27435 (N_27435,N_24241,N_25137);
and U27436 (N_27436,N_24920,N_24280);
or U27437 (N_27437,N_25211,N_24757);
or U27438 (N_27438,N_24415,N_25351);
nand U27439 (N_27439,N_24685,N_25108);
xnor U27440 (N_27440,N_24821,N_24237);
nor U27441 (N_27441,N_24183,N_25337);
and U27442 (N_27442,N_24996,N_24208);
or U27443 (N_27443,N_24749,N_24333);
nor U27444 (N_27444,N_24457,N_24055);
or U27445 (N_27445,N_25706,N_24791);
and U27446 (N_27446,N_25602,N_25866);
xnor U27447 (N_27447,N_24924,N_24213);
and U27448 (N_27448,N_24155,N_25881);
xnor U27449 (N_27449,N_25940,N_25397);
nand U27450 (N_27450,N_25861,N_24374);
nand U27451 (N_27451,N_24925,N_24154);
nand U27452 (N_27452,N_24020,N_25575);
and U27453 (N_27453,N_24710,N_24465);
or U27454 (N_27454,N_25957,N_25354);
xnor U27455 (N_27455,N_24207,N_25456);
xor U27456 (N_27456,N_24772,N_24732);
nor U27457 (N_27457,N_25024,N_24352);
nand U27458 (N_27458,N_24749,N_24150);
and U27459 (N_27459,N_25342,N_24764);
or U27460 (N_27460,N_25638,N_25342);
nor U27461 (N_27461,N_24711,N_24435);
xor U27462 (N_27462,N_25253,N_25135);
nor U27463 (N_27463,N_24794,N_24200);
nor U27464 (N_27464,N_24739,N_24588);
nand U27465 (N_27465,N_25546,N_24512);
or U27466 (N_27466,N_24565,N_25437);
xor U27467 (N_27467,N_24117,N_25938);
or U27468 (N_27468,N_25989,N_25058);
nand U27469 (N_27469,N_25528,N_25123);
nor U27470 (N_27470,N_24880,N_25346);
nor U27471 (N_27471,N_25036,N_25674);
or U27472 (N_27472,N_24286,N_25263);
nand U27473 (N_27473,N_25386,N_24406);
xor U27474 (N_27474,N_25681,N_25719);
and U27475 (N_27475,N_25678,N_25791);
nand U27476 (N_27476,N_25998,N_24539);
or U27477 (N_27477,N_24261,N_25390);
xnor U27478 (N_27478,N_25126,N_25497);
and U27479 (N_27479,N_25016,N_24785);
nand U27480 (N_27480,N_25816,N_25241);
and U27481 (N_27481,N_24925,N_24430);
and U27482 (N_27482,N_25001,N_24318);
xnor U27483 (N_27483,N_25869,N_24635);
and U27484 (N_27484,N_24575,N_24105);
and U27485 (N_27485,N_25193,N_25907);
or U27486 (N_27486,N_25218,N_25647);
xnor U27487 (N_27487,N_24531,N_25130);
nor U27488 (N_27488,N_25063,N_24750);
or U27489 (N_27489,N_24661,N_25651);
nand U27490 (N_27490,N_24523,N_25699);
or U27491 (N_27491,N_25134,N_24133);
or U27492 (N_27492,N_25377,N_25777);
xor U27493 (N_27493,N_25852,N_25390);
nor U27494 (N_27494,N_25659,N_24703);
xnor U27495 (N_27495,N_24881,N_24122);
nor U27496 (N_27496,N_25390,N_24579);
xnor U27497 (N_27497,N_24864,N_24095);
nor U27498 (N_27498,N_25837,N_24895);
and U27499 (N_27499,N_24183,N_24493);
xnor U27500 (N_27500,N_25390,N_24724);
xnor U27501 (N_27501,N_25232,N_24562);
nor U27502 (N_27502,N_24815,N_25953);
and U27503 (N_27503,N_24283,N_25986);
nand U27504 (N_27504,N_25549,N_25986);
or U27505 (N_27505,N_25269,N_24300);
nor U27506 (N_27506,N_25381,N_25633);
nand U27507 (N_27507,N_24866,N_24301);
nand U27508 (N_27508,N_25628,N_25523);
or U27509 (N_27509,N_25332,N_24097);
xnor U27510 (N_27510,N_25611,N_24142);
xor U27511 (N_27511,N_25684,N_25281);
nand U27512 (N_27512,N_24114,N_25653);
nand U27513 (N_27513,N_24586,N_24886);
xnor U27514 (N_27514,N_25974,N_24742);
nor U27515 (N_27515,N_24543,N_24413);
nor U27516 (N_27516,N_25977,N_24613);
or U27517 (N_27517,N_25312,N_25929);
and U27518 (N_27518,N_24399,N_25384);
nand U27519 (N_27519,N_25969,N_24258);
nand U27520 (N_27520,N_24354,N_24889);
or U27521 (N_27521,N_25105,N_25051);
nand U27522 (N_27522,N_25577,N_24119);
xor U27523 (N_27523,N_24215,N_24488);
xnor U27524 (N_27524,N_25552,N_25768);
nand U27525 (N_27525,N_24509,N_24385);
xor U27526 (N_27526,N_25645,N_24949);
and U27527 (N_27527,N_25248,N_25699);
or U27528 (N_27528,N_24176,N_25224);
nor U27529 (N_27529,N_25534,N_25098);
or U27530 (N_27530,N_25138,N_25509);
nor U27531 (N_27531,N_25094,N_25943);
nand U27532 (N_27532,N_25467,N_24990);
and U27533 (N_27533,N_24089,N_24834);
xnor U27534 (N_27534,N_24115,N_24385);
nor U27535 (N_27535,N_24789,N_25830);
nor U27536 (N_27536,N_25439,N_25485);
xor U27537 (N_27537,N_25708,N_25403);
nand U27538 (N_27538,N_25865,N_24504);
xor U27539 (N_27539,N_24724,N_24283);
and U27540 (N_27540,N_24160,N_25019);
or U27541 (N_27541,N_25889,N_24860);
xor U27542 (N_27542,N_25910,N_25101);
or U27543 (N_27543,N_25349,N_25013);
xor U27544 (N_27544,N_25076,N_24343);
and U27545 (N_27545,N_24549,N_25129);
nor U27546 (N_27546,N_24539,N_25846);
or U27547 (N_27547,N_25921,N_25743);
xnor U27548 (N_27548,N_24380,N_24854);
nand U27549 (N_27549,N_25557,N_24480);
or U27550 (N_27550,N_25115,N_24619);
nand U27551 (N_27551,N_25608,N_25459);
or U27552 (N_27552,N_25499,N_24453);
xnor U27553 (N_27553,N_25624,N_24927);
nand U27554 (N_27554,N_24385,N_25957);
xor U27555 (N_27555,N_24366,N_25924);
and U27556 (N_27556,N_25719,N_25950);
or U27557 (N_27557,N_25175,N_24932);
and U27558 (N_27558,N_24927,N_24078);
and U27559 (N_27559,N_24958,N_24633);
nor U27560 (N_27560,N_24935,N_24179);
or U27561 (N_27561,N_24228,N_24693);
nand U27562 (N_27562,N_25383,N_24038);
xnor U27563 (N_27563,N_25365,N_24071);
nand U27564 (N_27564,N_24897,N_25613);
or U27565 (N_27565,N_25169,N_25950);
nor U27566 (N_27566,N_25107,N_24882);
xor U27567 (N_27567,N_24643,N_25069);
or U27568 (N_27568,N_24952,N_24754);
nor U27569 (N_27569,N_25721,N_24328);
xnor U27570 (N_27570,N_24042,N_24280);
nor U27571 (N_27571,N_25145,N_25377);
nand U27572 (N_27572,N_24290,N_24161);
nand U27573 (N_27573,N_24988,N_25254);
or U27574 (N_27574,N_25347,N_24268);
nand U27575 (N_27575,N_25612,N_24577);
and U27576 (N_27576,N_25661,N_24589);
and U27577 (N_27577,N_25413,N_24272);
and U27578 (N_27578,N_25008,N_25253);
and U27579 (N_27579,N_24391,N_24982);
or U27580 (N_27580,N_24640,N_25650);
xnor U27581 (N_27581,N_25291,N_24996);
or U27582 (N_27582,N_24767,N_24607);
nand U27583 (N_27583,N_24590,N_25525);
or U27584 (N_27584,N_24585,N_24086);
nor U27585 (N_27585,N_24446,N_25363);
or U27586 (N_27586,N_24476,N_24748);
nand U27587 (N_27587,N_25640,N_24528);
and U27588 (N_27588,N_24709,N_25265);
nor U27589 (N_27589,N_24315,N_24967);
nor U27590 (N_27590,N_24795,N_25072);
nor U27591 (N_27591,N_25646,N_25156);
xnor U27592 (N_27592,N_25764,N_25315);
and U27593 (N_27593,N_24523,N_24839);
nand U27594 (N_27594,N_24797,N_24111);
xor U27595 (N_27595,N_25143,N_24966);
and U27596 (N_27596,N_24740,N_24396);
xnor U27597 (N_27597,N_25919,N_24361);
xor U27598 (N_27598,N_24110,N_25169);
nor U27599 (N_27599,N_25018,N_24190);
nor U27600 (N_27600,N_24256,N_25720);
nand U27601 (N_27601,N_24201,N_24009);
nor U27602 (N_27602,N_25534,N_24574);
or U27603 (N_27603,N_24414,N_24984);
and U27604 (N_27604,N_25660,N_25732);
nor U27605 (N_27605,N_25975,N_24326);
xnor U27606 (N_27606,N_25702,N_25249);
nand U27607 (N_27607,N_24687,N_25056);
or U27608 (N_27608,N_24330,N_25915);
and U27609 (N_27609,N_24540,N_25052);
xnor U27610 (N_27610,N_24223,N_25320);
nand U27611 (N_27611,N_25239,N_25906);
or U27612 (N_27612,N_25396,N_24402);
xnor U27613 (N_27613,N_24708,N_25755);
xnor U27614 (N_27614,N_25539,N_24452);
nand U27615 (N_27615,N_25181,N_25393);
nand U27616 (N_27616,N_24257,N_24574);
and U27617 (N_27617,N_25539,N_24771);
or U27618 (N_27618,N_24118,N_24823);
and U27619 (N_27619,N_25580,N_25726);
or U27620 (N_27620,N_24715,N_24740);
and U27621 (N_27621,N_25063,N_25500);
nor U27622 (N_27622,N_24215,N_24854);
nor U27623 (N_27623,N_25978,N_25769);
nand U27624 (N_27624,N_25509,N_25860);
or U27625 (N_27625,N_25560,N_24107);
and U27626 (N_27626,N_25141,N_24779);
nor U27627 (N_27627,N_25006,N_24779);
or U27628 (N_27628,N_25369,N_24881);
or U27629 (N_27629,N_25680,N_24178);
nand U27630 (N_27630,N_24148,N_25755);
xnor U27631 (N_27631,N_24624,N_25166);
or U27632 (N_27632,N_25843,N_25953);
or U27633 (N_27633,N_24000,N_24049);
nand U27634 (N_27634,N_25871,N_24179);
or U27635 (N_27635,N_24638,N_24389);
nor U27636 (N_27636,N_25811,N_25894);
nand U27637 (N_27637,N_25741,N_25114);
xor U27638 (N_27638,N_24926,N_24651);
nor U27639 (N_27639,N_24156,N_24996);
xnor U27640 (N_27640,N_24563,N_24770);
xnor U27641 (N_27641,N_25783,N_25535);
and U27642 (N_27642,N_24058,N_25518);
and U27643 (N_27643,N_24328,N_25839);
or U27644 (N_27644,N_25987,N_25340);
nand U27645 (N_27645,N_25035,N_25190);
xor U27646 (N_27646,N_24762,N_25923);
or U27647 (N_27647,N_24111,N_25389);
nor U27648 (N_27648,N_24818,N_25572);
nand U27649 (N_27649,N_25947,N_24123);
and U27650 (N_27650,N_24521,N_24723);
nand U27651 (N_27651,N_24993,N_25834);
or U27652 (N_27652,N_24616,N_25076);
nor U27653 (N_27653,N_25025,N_25158);
and U27654 (N_27654,N_25960,N_24951);
xor U27655 (N_27655,N_24361,N_24039);
or U27656 (N_27656,N_24255,N_24286);
and U27657 (N_27657,N_24499,N_24574);
and U27658 (N_27658,N_24351,N_24369);
xor U27659 (N_27659,N_24735,N_25619);
xor U27660 (N_27660,N_25849,N_25470);
nor U27661 (N_27661,N_25230,N_24881);
nor U27662 (N_27662,N_24054,N_25550);
and U27663 (N_27663,N_24447,N_25943);
and U27664 (N_27664,N_24544,N_24684);
and U27665 (N_27665,N_24447,N_25136);
xor U27666 (N_27666,N_25234,N_25370);
nand U27667 (N_27667,N_25084,N_24138);
xnor U27668 (N_27668,N_24207,N_25066);
or U27669 (N_27669,N_25791,N_24035);
nor U27670 (N_27670,N_24626,N_25739);
nor U27671 (N_27671,N_24520,N_25595);
xor U27672 (N_27672,N_24808,N_24659);
and U27673 (N_27673,N_25930,N_24141);
nand U27674 (N_27674,N_25262,N_24510);
xor U27675 (N_27675,N_25896,N_24178);
nor U27676 (N_27676,N_25165,N_24051);
or U27677 (N_27677,N_25704,N_24091);
and U27678 (N_27678,N_25183,N_24218);
xnor U27679 (N_27679,N_25436,N_25663);
nand U27680 (N_27680,N_24402,N_25340);
nor U27681 (N_27681,N_25446,N_25325);
nand U27682 (N_27682,N_25639,N_24674);
xnor U27683 (N_27683,N_24743,N_25057);
and U27684 (N_27684,N_24380,N_24373);
xor U27685 (N_27685,N_24390,N_25891);
nand U27686 (N_27686,N_25294,N_24385);
or U27687 (N_27687,N_24275,N_25039);
nor U27688 (N_27688,N_25751,N_25493);
nor U27689 (N_27689,N_24855,N_24407);
or U27690 (N_27690,N_24903,N_25247);
nand U27691 (N_27691,N_24806,N_25287);
nor U27692 (N_27692,N_24253,N_24596);
or U27693 (N_27693,N_24221,N_25317);
nor U27694 (N_27694,N_24756,N_25662);
and U27695 (N_27695,N_24036,N_24267);
nand U27696 (N_27696,N_24715,N_25884);
or U27697 (N_27697,N_24683,N_25930);
and U27698 (N_27698,N_24152,N_24032);
or U27699 (N_27699,N_24505,N_24519);
nand U27700 (N_27700,N_24260,N_25145);
xnor U27701 (N_27701,N_24886,N_24903);
xnor U27702 (N_27702,N_24341,N_24931);
nor U27703 (N_27703,N_24968,N_25263);
xnor U27704 (N_27704,N_24845,N_24704);
xnor U27705 (N_27705,N_24365,N_24252);
and U27706 (N_27706,N_25661,N_25383);
and U27707 (N_27707,N_24773,N_24526);
or U27708 (N_27708,N_24948,N_24402);
or U27709 (N_27709,N_25907,N_24787);
nand U27710 (N_27710,N_25599,N_24683);
and U27711 (N_27711,N_24092,N_25614);
xor U27712 (N_27712,N_24275,N_25056);
nor U27713 (N_27713,N_25427,N_24227);
xnor U27714 (N_27714,N_25533,N_24438);
or U27715 (N_27715,N_24967,N_24335);
nor U27716 (N_27716,N_24410,N_24393);
or U27717 (N_27717,N_24627,N_25075);
nand U27718 (N_27718,N_25958,N_25793);
nand U27719 (N_27719,N_25943,N_24628);
nor U27720 (N_27720,N_25336,N_25834);
nand U27721 (N_27721,N_25139,N_24369);
nand U27722 (N_27722,N_24061,N_25498);
nor U27723 (N_27723,N_25009,N_25338);
nand U27724 (N_27724,N_24071,N_24671);
nand U27725 (N_27725,N_25519,N_25722);
xnor U27726 (N_27726,N_25265,N_24212);
or U27727 (N_27727,N_24072,N_25980);
or U27728 (N_27728,N_25517,N_25358);
or U27729 (N_27729,N_24136,N_25190);
and U27730 (N_27730,N_25851,N_25577);
nand U27731 (N_27731,N_25025,N_24770);
nand U27732 (N_27732,N_24544,N_25363);
xnor U27733 (N_27733,N_24547,N_24350);
xnor U27734 (N_27734,N_25253,N_25918);
and U27735 (N_27735,N_24077,N_24796);
and U27736 (N_27736,N_25061,N_24816);
nand U27737 (N_27737,N_25905,N_25615);
xor U27738 (N_27738,N_25835,N_25708);
or U27739 (N_27739,N_25704,N_24469);
xnor U27740 (N_27740,N_25431,N_24992);
and U27741 (N_27741,N_25091,N_24124);
xnor U27742 (N_27742,N_24425,N_24042);
or U27743 (N_27743,N_24888,N_24880);
and U27744 (N_27744,N_24779,N_24522);
or U27745 (N_27745,N_25502,N_25996);
nor U27746 (N_27746,N_25464,N_24927);
and U27747 (N_27747,N_24170,N_24855);
or U27748 (N_27748,N_25447,N_25677);
and U27749 (N_27749,N_25406,N_24077);
nor U27750 (N_27750,N_24790,N_25340);
xnor U27751 (N_27751,N_24306,N_25518);
nor U27752 (N_27752,N_24671,N_24361);
or U27753 (N_27753,N_25738,N_24596);
and U27754 (N_27754,N_24931,N_24475);
nor U27755 (N_27755,N_24260,N_25127);
xor U27756 (N_27756,N_25481,N_25807);
nor U27757 (N_27757,N_24497,N_25945);
nand U27758 (N_27758,N_25086,N_25777);
and U27759 (N_27759,N_24761,N_25470);
or U27760 (N_27760,N_24022,N_24126);
and U27761 (N_27761,N_24276,N_25092);
and U27762 (N_27762,N_25192,N_25263);
nand U27763 (N_27763,N_24059,N_25235);
nand U27764 (N_27764,N_25616,N_25363);
and U27765 (N_27765,N_25632,N_25368);
and U27766 (N_27766,N_25946,N_25287);
nand U27767 (N_27767,N_24241,N_25715);
nand U27768 (N_27768,N_25554,N_24671);
nor U27769 (N_27769,N_24178,N_25963);
nand U27770 (N_27770,N_25677,N_25633);
or U27771 (N_27771,N_24070,N_25572);
and U27772 (N_27772,N_25681,N_25649);
nor U27773 (N_27773,N_24103,N_24697);
nor U27774 (N_27774,N_25829,N_25986);
or U27775 (N_27775,N_25468,N_24464);
nand U27776 (N_27776,N_25212,N_24617);
xor U27777 (N_27777,N_25207,N_24790);
nand U27778 (N_27778,N_24524,N_24551);
and U27779 (N_27779,N_24912,N_24844);
and U27780 (N_27780,N_24210,N_24253);
or U27781 (N_27781,N_25384,N_24138);
nor U27782 (N_27782,N_25516,N_25429);
nand U27783 (N_27783,N_24092,N_25723);
and U27784 (N_27784,N_24056,N_24990);
nand U27785 (N_27785,N_24439,N_25712);
nor U27786 (N_27786,N_24001,N_25199);
nand U27787 (N_27787,N_25405,N_25491);
or U27788 (N_27788,N_24313,N_25199);
and U27789 (N_27789,N_25416,N_25529);
nor U27790 (N_27790,N_24498,N_24966);
nor U27791 (N_27791,N_25961,N_24873);
or U27792 (N_27792,N_25767,N_25999);
and U27793 (N_27793,N_25399,N_24062);
and U27794 (N_27794,N_25128,N_25268);
xor U27795 (N_27795,N_24845,N_25221);
and U27796 (N_27796,N_24795,N_25511);
nor U27797 (N_27797,N_25672,N_25042);
nor U27798 (N_27798,N_24736,N_24197);
xnor U27799 (N_27799,N_25507,N_24571);
nor U27800 (N_27800,N_25956,N_24772);
and U27801 (N_27801,N_25413,N_24110);
nor U27802 (N_27802,N_25491,N_24471);
or U27803 (N_27803,N_25499,N_25494);
xor U27804 (N_27804,N_25425,N_25605);
or U27805 (N_27805,N_25846,N_25025);
nand U27806 (N_27806,N_25443,N_25925);
and U27807 (N_27807,N_25521,N_25896);
and U27808 (N_27808,N_25950,N_25604);
nand U27809 (N_27809,N_25725,N_24942);
nor U27810 (N_27810,N_25821,N_24781);
nand U27811 (N_27811,N_24910,N_25130);
xor U27812 (N_27812,N_24797,N_25553);
and U27813 (N_27813,N_24909,N_25402);
xor U27814 (N_27814,N_24811,N_25449);
xor U27815 (N_27815,N_24977,N_24831);
and U27816 (N_27816,N_24824,N_24072);
nor U27817 (N_27817,N_24141,N_24035);
nor U27818 (N_27818,N_25477,N_25066);
or U27819 (N_27819,N_25387,N_24240);
nor U27820 (N_27820,N_24645,N_25042);
or U27821 (N_27821,N_25195,N_24106);
nor U27822 (N_27822,N_24958,N_25120);
nor U27823 (N_27823,N_25696,N_24914);
nand U27824 (N_27824,N_24894,N_24194);
xor U27825 (N_27825,N_25247,N_25872);
and U27826 (N_27826,N_24380,N_24558);
nand U27827 (N_27827,N_24530,N_25434);
xor U27828 (N_27828,N_24481,N_25818);
nor U27829 (N_27829,N_25353,N_24858);
nand U27830 (N_27830,N_24225,N_25352);
and U27831 (N_27831,N_25717,N_25491);
xnor U27832 (N_27832,N_25770,N_24406);
xor U27833 (N_27833,N_24818,N_24478);
nor U27834 (N_27834,N_24465,N_25982);
nand U27835 (N_27835,N_25364,N_25894);
nand U27836 (N_27836,N_24735,N_25210);
or U27837 (N_27837,N_25013,N_25466);
xnor U27838 (N_27838,N_25164,N_24292);
and U27839 (N_27839,N_24640,N_25028);
nand U27840 (N_27840,N_25089,N_24144);
xor U27841 (N_27841,N_25022,N_25651);
and U27842 (N_27842,N_24363,N_24753);
or U27843 (N_27843,N_24014,N_25311);
nand U27844 (N_27844,N_25159,N_24919);
nand U27845 (N_27845,N_25657,N_25015);
xor U27846 (N_27846,N_25650,N_25888);
xor U27847 (N_27847,N_25933,N_25010);
nand U27848 (N_27848,N_24684,N_24750);
nand U27849 (N_27849,N_25234,N_24262);
nand U27850 (N_27850,N_24099,N_24778);
nor U27851 (N_27851,N_24563,N_25274);
and U27852 (N_27852,N_25196,N_24039);
or U27853 (N_27853,N_24756,N_25241);
and U27854 (N_27854,N_25936,N_25149);
nor U27855 (N_27855,N_25381,N_24995);
or U27856 (N_27856,N_25045,N_25030);
nand U27857 (N_27857,N_25085,N_25403);
and U27858 (N_27858,N_25630,N_25804);
nor U27859 (N_27859,N_25199,N_24245);
and U27860 (N_27860,N_25859,N_25616);
xnor U27861 (N_27861,N_24725,N_25707);
xor U27862 (N_27862,N_25272,N_25405);
xor U27863 (N_27863,N_25299,N_24292);
xnor U27864 (N_27864,N_25089,N_24538);
xnor U27865 (N_27865,N_25258,N_24296);
nand U27866 (N_27866,N_24602,N_25198);
and U27867 (N_27867,N_24687,N_25310);
xnor U27868 (N_27868,N_25435,N_24839);
nand U27869 (N_27869,N_24279,N_24185);
xnor U27870 (N_27870,N_24898,N_24754);
xnor U27871 (N_27871,N_25966,N_25689);
nand U27872 (N_27872,N_24311,N_24611);
nand U27873 (N_27873,N_25362,N_24086);
nand U27874 (N_27874,N_25125,N_24816);
and U27875 (N_27875,N_24407,N_25241);
xor U27876 (N_27876,N_25031,N_25695);
xor U27877 (N_27877,N_25792,N_25119);
or U27878 (N_27878,N_25938,N_25465);
xnor U27879 (N_27879,N_24929,N_25918);
nor U27880 (N_27880,N_25800,N_25276);
nor U27881 (N_27881,N_25513,N_24929);
and U27882 (N_27882,N_24534,N_25584);
and U27883 (N_27883,N_24853,N_25889);
or U27884 (N_27884,N_25946,N_25022);
or U27885 (N_27885,N_25947,N_25708);
nand U27886 (N_27886,N_25976,N_24133);
nand U27887 (N_27887,N_25866,N_24865);
and U27888 (N_27888,N_25400,N_24560);
nor U27889 (N_27889,N_24786,N_24921);
xor U27890 (N_27890,N_25343,N_25155);
and U27891 (N_27891,N_25136,N_25628);
or U27892 (N_27892,N_25201,N_25784);
nor U27893 (N_27893,N_24483,N_25179);
nand U27894 (N_27894,N_25808,N_24027);
nor U27895 (N_27895,N_25660,N_25073);
and U27896 (N_27896,N_24137,N_24854);
nor U27897 (N_27897,N_24760,N_24499);
and U27898 (N_27898,N_24621,N_24715);
nor U27899 (N_27899,N_25353,N_24335);
xnor U27900 (N_27900,N_24429,N_24456);
and U27901 (N_27901,N_24018,N_24428);
nand U27902 (N_27902,N_25260,N_24113);
or U27903 (N_27903,N_24515,N_24938);
xnor U27904 (N_27904,N_24041,N_24541);
nand U27905 (N_27905,N_25757,N_24632);
xor U27906 (N_27906,N_25095,N_24392);
nor U27907 (N_27907,N_25640,N_25273);
nand U27908 (N_27908,N_25409,N_24235);
and U27909 (N_27909,N_24728,N_24290);
xor U27910 (N_27910,N_25224,N_25658);
or U27911 (N_27911,N_25716,N_24438);
and U27912 (N_27912,N_24264,N_24299);
or U27913 (N_27913,N_25119,N_24911);
or U27914 (N_27914,N_24741,N_24214);
and U27915 (N_27915,N_25145,N_24951);
nor U27916 (N_27916,N_24599,N_25469);
nor U27917 (N_27917,N_24187,N_24278);
and U27918 (N_27918,N_24796,N_25535);
nand U27919 (N_27919,N_25963,N_24779);
or U27920 (N_27920,N_25004,N_24753);
xnor U27921 (N_27921,N_25727,N_24561);
or U27922 (N_27922,N_25947,N_24884);
and U27923 (N_27923,N_24094,N_25067);
xnor U27924 (N_27924,N_25248,N_24663);
or U27925 (N_27925,N_24255,N_24052);
xor U27926 (N_27926,N_25281,N_25331);
nor U27927 (N_27927,N_24883,N_25140);
and U27928 (N_27928,N_24302,N_25970);
xnor U27929 (N_27929,N_25367,N_25759);
xnor U27930 (N_27930,N_25170,N_24112);
nand U27931 (N_27931,N_25108,N_24098);
and U27932 (N_27932,N_25676,N_25584);
nand U27933 (N_27933,N_24815,N_25389);
or U27934 (N_27934,N_24672,N_25954);
or U27935 (N_27935,N_24439,N_24186);
xnor U27936 (N_27936,N_25590,N_24708);
nor U27937 (N_27937,N_25041,N_24762);
nand U27938 (N_27938,N_25472,N_24806);
and U27939 (N_27939,N_24700,N_24744);
nor U27940 (N_27940,N_24633,N_24781);
and U27941 (N_27941,N_25169,N_24945);
nor U27942 (N_27942,N_24631,N_25729);
or U27943 (N_27943,N_24158,N_24471);
nor U27944 (N_27944,N_24869,N_25938);
nor U27945 (N_27945,N_24732,N_25971);
nand U27946 (N_27946,N_25479,N_24403);
nand U27947 (N_27947,N_25521,N_24461);
and U27948 (N_27948,N_24305,N_24633);
nor U27949 (N_27949,N_24340,N_25967);
or U27950 (N_27950,N_25414,N_25142);
nor U27951 (N_27951,N_25433,N_24207);
and U27952 (N_27952,N_24089,N_25546);
nand U27953 (N_27953,N_24672,N_25931);
xor U27954 (N_27954,N_24948,N_24643);
and U27955 (N_27955,N_25088,N_24821);
or U27956 (N_27956,N_24309,N_25224);
nand U27957 (N_27957,N_24257,N_25745);
nand U27958 (N_27958,N_25443,N_25368);
or U27959 (N_27959,N_25289,N_24318);
and U27960 (N_27960,N_25969,N_24491);
xnor U27961 (N_27961,N_24759,N_25169);
or U27962 (N_27962,N_24154,N_24188);
and U27963 (N_27963,N_24580,N_24918);
nor U27964 (N_27964,N_25124,N_25431);
xnor U27965 (N_27965,N_25597,N_25629);
and U27966 (N_27966,N_25219,N_25344);
and U27967 (N_27967,N_24176,N_24771);
or U27968 (N_27968,N_24932,N_24034);
nand U27969 (N_27969,N_24660,N_24417);
xnor U27970 (N_27970,N_24518,N_25786);
or U27971 (N_27971,N_24402,N_25067);
or U27972 (N_27972,N_24583,N_24851);
and U27973 (N_27973,N_24891,N_24258);
nand U27974 (N_27974,N_24865,N_25217);
xnor U27975 (N_27975,N_25280,N_24575);
nand U27976 (N_27976,N_25842,N_24159);
nand U27977 (N_27977,N_25131,N_24375);
nor U27978 (N_27978,N_25900,N_25798);
nor U27979 (N_27979,N_25738,N_25623);
and U27980 (N_27980,N_24488,N_25688);
xor U27981 (N_27981,N_24638,N_25110);
xnor U27982 (N_27982,N_25655,N_24531);
nand U27983 (N_27983,N_24618,N_24647);
xnor U27984 (N_27984,N_25414,N_24038);
nand U27985 (N_27985,N_24426,N_25148);
or U27986 (N_27986,N_25688,N_24094);
nor U27987 (N_27987,N_25598,N_25282);
nor U27988 (N_27988,N_25087,N_25675);
and U27989 (N_27989,N_25837,N_25143);
or U27990 (N_27990,N_24717,N_25702);
and U27991 (N_27991,N_25572,N_25190);
nor U27992 (N_27992,N_25801,N_25198);
xor U27993 (N_27993,N_25227,N_25292);
nor U27994 (N_27994,N_25236,N_24568);
or U27995 (N_27995,N_24543,N_25436);
nand U27996 (N_27996,N_25106,N_25797);
or U27997 (N_27997,N_25805,N_24269);
or U27998 (N_27998,N_25923,N_24478);
and U27999 (N_27999,N_24326,N_25872);
nand U28000 (N_28000,N_26754,N_27038);
nand U28001 (N_28001,N_26622,N_27909);
and U28002 (N_28002,N_27275,N_27488);
nand U28003 (N_28003,N_26810,N_27298);
nand U28004 (N_28004,N_26154,N_27740);
nand U28005 (N_28005,N_27901,N_26297);
nor U28006 (N_28006,N_26058,N_26296);
and U28007 (N_28007,N_27819,N_27782);
and U28008 (N_28008,N_26837,N_27513);
nand U28009 (N_28009,N_27766,N_26174);
nand U28010 (N_28010,N_27630,N_27375);
xnor U28011 (N_28011,N_26488,N_26924);
xor U28012 (N_28012,N_26213,N_27885);
nand U28013 (N_28013,N_27582,N_26564);
nand U28014 (N_28014,N_27129,N_26280);
nand U28015 (N_28015,N_26368,N_26127);
nand U28016 (N_28016,N_26984,N_26653);
and U28017 (N_28017,N_26846,N_27732);
and U28018 (N_28018,N_26133,N_26437);
nor U28019 (N_28019,N_27199,N_27430);
nor U28020 (N_28020,N_27382,N_27510);
and U28021 (N_28021,N_27378,N_27037);
nor U28022 (N_28022,N_27914,N_27136);
or U28023 (N_28023,N_26983,N_27745);
or U28024 (N_28024,N_27683,N_27486);
or U28025 (N_28025,N_26911,N_26552);
nor U28026 (N_28026,N_26500,N_27429);
and U28027 (N_28027,N_26729,N_27159);
xnor U28028 (N_28028,N_26940,N_27703);
and U28029 (N_28029,N_26389,N_27717);
and U28030 (N_28030,N_26966,N_26934);
nor U28031 (N_28031,N_27137,N_26992);
nand U28032 (N_28032,N_26311,N_27534);
and U28033 (N_28033,N_26864,N_26139);
or U28034 (N_28034,N_27074,N_26304);
xnor U28035 (N_28035,N_27781,N_26972);
or U28036 (N_28036,N_26786,N_26167);
nand U28037 (N_28037,N_27157,N_27844);
nand U28038 (N_28038,N_26755,N_26651);
xnor U28039 (N_28039,N_26021,N_26890);
and U28040 (N_28040,N_26737,N_27072);
and U28041 (N_28041,N_26884,N_27975);
nand U28042 (N_28042,N_26387,N_27104);
nand U28043 (N_28043,N_27301,N_27229);
and U28044 (N_28044,N_27684,N_27905);
nor U28045 (N_28045,N_26852,N_27804);
or U28046 (N_28046,N_27539,N_26602);
xnor U28047 (N_28047,N_26218,N_27706);
and U28048 (N_28048,N_26862,N_27964);
nor U28049 (N_28049,N_27259,N_26733);
nand U28050 (N_28050,N_26738,N_27249);
xnor U28051 (N_28051,N_27609,N_27869);
and U28052 (N_28052,N_27695,N_26750);
or U28053 (N_28053,N_27460,N_26912);
nor U28054 (N_28054,N_27134,N_26608);
and U28055 (N_28055,N_26143,N_26455);
nor U28056 (N_28056,N_26854,N_26111);
or U28057 (N_28057,N_27309,N_26956);
xnor U28058 (N_28058,N_27030,N_26996);
or U28059 (N_28059,N_26877,N_26449);
nor U28060 (N_28060,N_27726,N_26509);
or U28061 (N_28061,N_27791,N_27212);
or U28062 (N_28062,N_27682,N_27640);
and U28063 (N_28063,N_27599,N_27768);
and U28064 (N_28064,N_26614,N_27365);
xor U28065 (N_28065,N_27141,N_26530);
and U28066 (N_28066,N_26421,N_27923);
nor U28067 (N_28067,N_26736,N_26981);
nand U28068 (N_28068,N_27800,N_26438);
or U28069 (N_28069,N_26403,N_26201);
or U28070 (N_28070,N_26517,N_27160);
and U28071 (N_28071,N_27542,N_26192);
nor U28072 (N_28072,N_27152,N_26360);
nand U28073 (N_28073,N_27638,N_27431);
xor U28074 (N_28074,N_27451,N_27763);
and U28075 (N_28075,N_26534,N_27960);
or U28076 (N_28076,N_27324,N_26392);
xor U28077 (N_28077,N_27366,N_27364);
nor U28078 (N_28078,N_27256,N_27242);
xnor U28079 (N_28079,N_26629,N_27057);
and U28080 (N_28080,N_27461,N_27776);
xnor U28081 (N_28081,N_26723,N_26978);
nand U28082 (N_28082,N_27773,N_27385);
xnor U28083 (N_28083,N_26856,N_27564);
xor U28084 (N_28084,N_27633,N_26395);
or U28085 (N_28085,N_26533,N_27308);
nor U28086 (N_28086,N_26585,N_27325);
or U28087 (N_28087,N_27926,N_27743);
xnor U28088 (N_28088,N_26943,N_26319);
or U28089 (N_28089,N_26005,N_26334);
nand U28090 (N_28090,N_26496,N_27871);
or U28091 (N_28091,N_26901,N_26107);
or U28092 (N_28092,N_27827,N_27641);
or U28093 (N_28093,N_27171,N_26510);
nor U28094 (N_28094,N_26646,N_26947);
or U28095 (N_28095,N_27658,N_26898);
xnor U28096 (N_28096,N_27462,N_27532);
xnor U28097 (N_28097,N_26427,N_26049);
and U28098 (N_28098,N_27587,N_27016);
nor U28099 (N_28099,N_26958,N_27333);
xnor U28100 (N_28100,N_27233,N_27811);
nand U28101 (N_28101,N_26609,N_26380);
xor U28102 (N_28102,N_26698,N_27036);
nand U28103 (N_28103,N_27696,N_27814);
or U28104 (N_28104,N_26887,N_26477);
nand U28105 (N_28105,N_26807,N_26161);
nor U28106 (N_28106,N_26374,N_26732);
xor U28107 (N_28107,N_26706,N_27055);
nor U28108 (N_28108,N_27762,N_27224);
and U28109 (N_28109,N_26244,N_27268);
nor U28110 (N_28110,N_26386,N_26229);
xor U28111 (N_28111,N_27497,N_26868);
and U28112 (N_28112,N_27345,N_27786);
nand U28113 (N_28113,N_27705,N_26915);
and U28114 (N_28114,N_26397,N_26048);
nand U28115 (N_28115,N_26265,N_27395);
nand U28116 (N_28116,N_27215,N_26444);
and U28117 (N_28117,N_26556,N_27413);
nand U28118 (N_28118,N_27949,N_27691);
nor U28119 (N_28119,N_27779,N_27133);
nor U28120 (N_28120,N_27986,N_26502);
nand U28121 (N_28121,N_27573,N_27329);
xnor U28122 (N_28122,N_27409,N_27481);
nor U28123 (N_28123,N_27759,N_27288);
and U28124 (N_28124,N_27831,N_26962);
or U28125 (N_28125,N_27687,N_26279);
and U28126 (N_28126,N_27485,N_27033);
xor U28127 (N_28127,N_26839,N_27627);
xor U28128 (N_28128,N_26333,N_27521);
xnor U28129 (N_28129,N_27220,N_27116);
nand U28130 (N_28130,N_26591,N_27003);
nor U28131 (N_28131,N_27115,N_26761);
or U28132 (N_28132,N_27803,N_26518);
nand U28133 (N_28133,N_27892,N_26151);
xnor U28134 (N_28134,N_26486,N_26109);
nand U28135 (N_28135,N_27648,N_26480);
nor U28136 (N_28136,N_27203,N_27320);
nand U28137 (N_28137,N_27188,N_26372);
and U28138 (N_28138,N_26687,N_26573);
nand U28139 (N_28139,N_27492,N_26679);
nand U28140 (N_28140,N_27402,N_26011);
and U28141 (N_28141,N_26595,N_26832);
xnor U28142 (N_28142,N_26655,N_27565);
nor U28143 (N_28143,N_26963,N_27290);
xnor U28144 (N_28144,N_26809,N_27164);
xor U28145 (N_28145,N_27541,N_26867);
nand U28146 (N_28146,N_27351,N_27792);
nor U28147 (N_28147,N_27623,N_26147);
and U28148 (N_28148,N_27068,N_27533);
nor U28149 (N_28149,N_26952,N_27647);
nor U28150 (N_28150,N_27246,N_27285);
or U28151 (N_28151,N_26288,N_27213);
nor U28152 (N_28152,N_26578,N_27227);
or U28153 (N_28153,N_26183,N_26788);
and U28154 (N_28154,N_27128,N_26467);
nand U28155 (N_28155,N_27177,N_26598);
or U28156 (N_28156,N_27962,N_26287);
xor U28157 (N_28157,N_27783,N_26880);
nand U28158 (N_28158,N_26835,N_27670);
nand U28159 (N_28159,N_27379,N_27219);
and U28160 (N_28160,N_27459,N_26052);
nor U28161 (N_28161,N_26321,N_26462);
nor U28162 (N_28162,N_26926,N_26769);
or U28163 (N_28163,N_27080,N_27591);
and U28164 (N_28164,N_26762,N_27973);
nand U28165 (N_28165,N_27954,N_27942);
nand U28166 (N_28166,N_26569,N_26199);
xor U28167 (N_28167,N_27702,N_26085);
nand U28168 (N_28168,N_27678,N_27861);
and U28169 (N_28169,N_27383,N_26930);
nand U28170 (N_28170,N_27850,N_26938);
nor U28171 (N_28171,N_26110,N_26941);
nand U28172 (N_28172,N_26450,N_26285);
nand U28173 (N_28173,N_26672,N_26774);
and U28174 (N_28174,N_27515,N_26936);
or U28175 (N_28175,N_27557,N_27833);
or U28176 (N_28176,N_27748,N_27316);
or U28177 (N_28177,N_26231,N_26882);
nand U28178 (N_28178,N_27606,N_26439);
xor U28179 (N_28179,N_27990,N_26253);
and U28180 (N_28180,N_27908,N_27253);
or U28181 (N_28181,N_26155,N_27569);
or U28182 (N_28182,N_26281,N_27929);
xor U28183 (N_28183,N_27966,N_27289);
nand U28184 (N_28184,N_26035,N_27083);
nor U28185 (N_28185,N_26907,N_27730);
nor U28186 (N_28186,N_27019,N_27341);
nor U28187 (N_28187,N_27340,N_26291);
nand U28188 (N_28188,N_27335,N_26243);
or U28189 (N_28189,N_26259,N_27820);
xnor U28190 (N_28190,N_26416,N_27849);
nor U28191 (N_28191,N_27698,N_26019);
and U28192 (N_28192,N_27151,N_26166);
nor U28193 (N_28193,N_26789,N_27053);
nand U28194 (N_28194,N_26588,N_26827);
and U28195 (N_28195,N_26802,N_27173);
or U28196 (N_28196,N_26512,N_26701);
nand U28197 (N_28197,N_27095,N_26193);
or U28198 (N_28198,N_26568,N_26634);
nor U28199 (N_28199,N_26409,N_26454);
or U28200 (N_28200,N_26604,N_26740);
xor U28201 (N_28201,N_26597,N_26337);
or U28202 (N_28202,N_26338,N_27267);
xnor U28203 (N_28203,N_27489,N_27368);
nand U28204 (N_28204,N_27491,N_27765);
or U28205 (N_28205,N_27060,N_27988);
nor U28206 (N_28206,N_26379,N_27423);
or U28207 (N_28207,N_27434,N_27167);
nand U28208 (N_28208,N_27545,N_27848);
or U28209 (N_28209,N_26886,N_27008);
and U28210 (N_28210,N_26982,N_26301);
xor U28211 (N_28211,N_26744,N_26341);
nor U28212 (N_28212,N_26353,N_27111);
xor U28213 (N_28213,N_26267,N_26808);
nor U28214 (N_28214,N_26413,N_26465);
xor U28215 (N_28215,N_27562,N_27651);
nand U28216 (N_28216,N_27657,N_26587);
and U28217 (N_28217,N_26641,N_27297);
nand U28218 (N_28218,N_27887,N_27311);
nor U28219 (N_28219,N_26643,N_27477);
or U28220 (N_28220,N_26866,N_27728);
nor U28221 (N_28221,N_26260,N_26069);
or U28222 (N_28222,N_26734,N_26241);
or U28223 (N_28223,N_27050,N_27493);
xnor U28224 (N_28224,N_26722,N_27663);
and U28225 (N_28225,N_26063,N_27900);
or U28226 (N_28226,N_26519,N_27420);
and U28227 (N_28227,N_27837,N_27868);
and U28228 (N_28228,N_27656,N_27693);
or U28229 (N_28229,N_26405,N_27452);
nand U28230 (N_28230,N_26221,N_27661);
xnor U28231 (N_28231,N_26921,N_26472);
xor U28232 (N_28232,N_27042,N_26136);
and U28233 (N_28233,N_27216,N_27098);
nor U28234 (N_28234,N_26527,N_27495);
nor U28235 (N_28235,N_26357,N_26275);
and U28236 (N_28236,N_26121,N_26092);
xnor U28237 (N_28237,N_27002,N_27147);
xor U28238 (N_28238,N_27807,N_26899);
xor U28239 (N_28239,N_27735,N_26343);
nor U28240 (N_28240,N_27239,N_26094);
and U28241 (N_28241,N_26727,N_26391);
nand U28242 (N_28242,N_26906,N_26836);
or U28243 (N_28243,N_26182,N_27859);
xor U28244 (N_28244,N_27632,N_27376);
and U28245 (N_28245,N_26566,N_26649);
xnor U28246 (N_28246,N_27218,N_27374);
xor U28247 (N_28247,N_26215,N_26950);
and U28248 (N_28248,N_27478,N_27207);
xnor U28249 (N_28249,N_27930,N_27736);
or U28250 (N_28250,N_27816,N_27471);
nand U28251 (N_28251,N_26217,N_27135);
xnor U28252 (N_28252,N_27070,N_26266);
nand U28253 (N_28253,N_27465,N_27982);
and U28254 (N_28254,N_26764,N_26986);
and U28255 (N_28255,N_26441,N_27314);
xor U28256 (N_28256,N_26659,N_27770);
nand U28257 (N_28257,N_27543,N_27397);
and U28258 (N_28258,N_27339,N_26383);
or U28259 (N_28259,N_27643,N_27563);
or U28260 (N_28260,N_26995,N_27404);
or U28261 (N_28261,N_27014,N_27009);
nor U28262 (N_28262,N_26861,N_27834);
nand U28263 (N_28263,N_27694,N_27408);
nand U28264 (N_28264,N_26440,N_26077);
or U28265 (N_28265,N_26696,N_26889);
or U28266 (N_28266,N_27815,N_26328);
or U28267 (N_28267,N_26445,N_26850);
nand U28268 (N_28268,N_26305,N_27716);
nand U28269 (N_28269,N_26900,N_26765);
or U28270 (N_28270,N_27888,N_26689);
nand U28271 (N_28271,N_27855,N_26473);
nand U28272 (N_28272,N_26425,N_27155);
xnor U28273 (N_28273,N_26637,N_27864);
nor U28274 (N_28274,N_26498,N_27051);
or U28275 (N_28275,N_27507,N_26865);
nor U28276 (N_28276,N_26753,N_26317);
xor U28277 (N_28277,N_27798,N_26306);
and U28278 (N_28278,N_27389,N_26909);
xnor U28279 (N_28279,N_27062,N_27778);
nand U28280 (N_28280,N_26088,N_26247);
nand U28281 (N_28281,N_27660,N_27384);
or U28282 (N_28282,N_26821,N_26492);
nand U28283 (N_28283,N_26414,N_27243);
nand U28284 (N_28284,N_26725,N_26490);
or U28285 (N_28285,N_26752,N_27963);
nand U28286 (N_28286,N_27953,N_26522);
or U28287 (N_28287,N_27830,N_27244);
nand U28288 (N_28288,N_27720,N_27056);
and U28289 (N_28289,N_27307,N_26070);
and U28290 (N_28290,N_27787,N_27993);
xor U28291 (N_28291,N_27299,N_26985);
or U28292 (N_28292,N_26816,N_26842);
or U28293 (N_28293,N_26504,N_27904);
nor U28294 (N_28294,N_27022,N_27598);
nand U28295 (N_28295,N_26030,N_27225);
or U28296 (N_28296,N_27553,N_26776);
and U28297 (N_28297,N_26785,N_27483);
nand U28298 (N_28298,N_27951,N_27235);
nand U28299 (N_28299,N_27432,N_27161);
nand U28300 (N_28300,N_27872,N_26156);
nand U28301 (N_28301,N_27040,N_26558);
xor U28302 (N_28302,N_26359,N_26895);
nor U28303 (N_28303,N_27639,N_26536);
nor U28304 (N_28304,N_26153,N_26954);
nor U28305 (N_28305,N_26819,N_27959);
or U28306 (N_28306,N_27920,N_26716);
xnor U28307 (N_28307,N_26951,N_27466);
nand U28308 (N_28308,N_27637,N_26903);
xor U28309 (N_28309,N_27449,N_26666);
nand U28310 (N_28310,N_27645,N_26363);
nor U28311 (N_28311,N_27529,N_27727);
nor U28312 (N_28312,N_27555,N_27097);
nor U28313 (N_28313,N_27439,N_26411);
nor U28314 (N_28314,N_27419,N_27091);
nor U28315 (N_28315,N_26778,N_26024);
nor U28316 (N_28316,N_27210,N_27749);
and U28317 (N_28317,N_27453,N_26162);
xor U28318 (N_28318,N_26757,N_26426);
nor U28319 (N_28319,N_27758,N_26150);
xor U28320 (N_28320,N_26017,N_27857);
nand U28321 (N_28321,N_26942,N_26977);
or U28322 (N_28322,N_26342,N_26097);
and U28323 (N_28323,N_27416,N_27502);
nand U28324 (N_28324,N_27472,N_27407);
nand U28325 (N_28325,N_26925,N_26042);
and U28326 (N_28326,N_26393,N_27596);
xor U28327 (N_28327,N_26245,N_26002);
xor U28328 (N_28328,N_27174,N_27729);
and U28329 (N_28329,N_26571,N_26014);
nand U28330 (N_28330,N_26929,N_27427);
xnor U28331 (N_28331,N_27337,N_26841);
nand U28332 (N_28332,N_27718,N_26505);
nand U28333 (N_28333,N_26482,N_26652);
or U28334 (N_28334,N_26032,N_27832);
and U28335 (N_28335,N_26550,N_26086);
nand U28336 (N_28336,N_26937,N_27989);
and U28337 (N_28337,N_26935,N_26225);
xor U28338 (N_28338,N_26410,N_26731);
and U28339 (N_28339,N_27520,N_26481);
or U28340 (N_28340,N_26545,N_27406);
nor U28341 (N_28341,N_26195,N_26168);
nand U28342 (N_28342,N_26662,N_27058);
and U28343 (N_28343,N_26686,N_27790);
or U28344 (N_28344,N_27899,N_26442);
nor U28345 (N_28345,N_27474,N_27677);
xor U28346 (N_28346,N_27808,N_27613);
nor U28347 (N_28347,N_26083,N_27952);
or U28348 (N_28348,N_26286,N_26623);
or U28349 (N_28349,N_27991,N_26547);
nand U28350 (N_28350,N_27755,N_27913);
nand U28351 (N_28351,N_26313,N_26016);
or U28352 (N_28352,N_27422,N_27655);
xor U28353 (N_28353,N_27286,N_26999);
nor U28354 (N_28354,N_27721,N_26001);
nor U28355 (N_28355,N_26830,N_26255);
nand U28356 (N_28356,N_26600,N_27858);
nand U28357 (N_28357,N_26575,N_26843);
nand U28358 (N_28358,N_26144,N_26431);
xnor U28359 (N_28359,N_26971,N_27110);
xnor U28360 (N_28360,N_27206,N_27874);
nand U28361 (N_28361,N_26152,N_26361);
nor U28362 (N_28362,N_26429,N_26893);
nand U28363 (N_28363,N_27496,N_26916);
nor U28364 (N_28364,N_27047,N_26565);
xor U28365 (N_28365,N_27873,N_27487);
nor U28366 (N_28366,N_26314,N_27204);
nand U28367 (N_28367,N_26117,N_26648);
nor U28368 (N_28368,N_26586,N_27580);
nor U28369 (N_28369,N_26775,N_27636);
xor U28370 (N_28370,N_27594,N_27245);
nor U28371 (N_28371,N_26207,N_27818);
xnor U28372 (N_28372,N_26428,N_27100);
or U28373 (N_28373,N_26399,N_27604);
or U28374 (N_28374,N_27535,N_27400);
or U28375 (N_28375,N_27331,N_27769);
or U28376 (N_28376,N_27073,N_27391);
xor U28377 (N_28377,N_26457,N_26513);
nand U28378 (N_28378,N_27469,N_26746);
or U28379 (N_28379,N_27722,N_27463);
xnor U28380 (N_28380,N_26922,N_27927);
nor U28381 (N_28381,N_26100,N_26344);
nand U28382 (N_28382,N_27775,N_26406);
and U28383 (N_28383,N_26064,N_26040);
nand U28384 (N_28384,N_26268,N_26621);
xor U28385 (N_28385,N_26814,N_27006);
nand U28386 (N_28386,N_26631,N_26851);
or U28387 (N_28387,N_26271,N_27209);
or U28388 (N_28388,N_26087,N_26186);
and U28389 (N_28389,N_27576,N_26329);
nand U28390 (N_28390,N_27078,N_27667);
xor U28391 (N_28391,N_27912,N_26028);
xor U28392 (N_28392,N_26184,N_27847);
and U28393 (N_28393,N_26787,N_27295);
nand U28394 (N_28394,N_27538,N_26347);
and U28395 (N_28395,N_26181,N_26061);
nand U28396 (N_28396,N_27258,N_26499);
or U28397 (N_28397,N_27032,N_26913);
nor U28398 (N_28398,N_26084,N_27659);
nand U28399 (N_28399,N_27123,N_27313);
nor U28400 (N_28400,N_27424,N_26619);
or U28401 (N_28401,N_26415,N_26180);
or U28402 (N_28402,N_26628,N_26220);
or U28403 (N_28403,N_26148,N_27937);
and U28404 (N_28404,N_27554,N_26176);
nor U28405 (N_28405,N_27955,N_27621);
or U28406 (N_28406,N_26918,N_26320);
or U28407 (N_28407,N_26349,N_27387);
nand U28408 (N_28408,N_26233,N_27023);
xnor U28409 (N_28409,N_26538,N_26620);
nor U28410 (N_28410,N_26066,N_27846);
and U28411 (N_28411,N_27697,N_27264);
nand U28412 (N_28412,N_26039,N_26551);
nand U28413 (N_28413,N_27250,N_26091);
or U28414 (N_28414,N_27113,N_27701);
nand U28415 (N_28415,N_26693,N_27059);
or U28416 (N_28416,N_26118,N_26194);
xnor U28417 (N_28417,N_27103,N_27214);
and U28418 (N_28418,N_26549,N_26855);
nand U28419 (N_28419,N_27148,N_27879);
and U28420 (N_28420,N_26015,N_27118);
nand U28421 (N_28421,N_27629,N_26236);
nor U28422 (N_28422,N_27838,N_27644);
xor U28423 (N_28423,N_26307,N_26712);
nor U28424 (N_28424,N_26404,N_27350);
or U28425 (N_28425,N_27079,N_27394);
and U28426 (N_28426,N_27835,N_27131);
nand U28427 (N_28427,N_27165,N_26770);
and U28428 (N_28428,N_26124,N_26171);
nand U28429 (N_28429,N_27983,N_27263);
and U28430 (N_28430,N_27935,N_26593);
or U28431 (N_28431,N_26370,N_26892);
nand U28432 (N_28432,N_27010,N_27524);
nor U28433 (N_28433,N_26535,N_26461);
nand U28434 (N_28434,N_26080,N_27940);
nand U28435 (N_28435,N_26185,N_27150);
or U28436 (N_28436,N_27772,N_27537);
and U28437 (N_28437,N_27168,N_27980);
and U28438 (N_28438,N_26615,N_27579);
and U28439 (N_28439,N_27294,N_27355);
and U28440 (N_28440,N_27447,N_26483);
xor U28441 (N_28441,N_27907,N_26020);
or U28442 (N_28442,N_27611,N_27744);
xor U28443 (N_28443,N_26089,N_26096);
xor U28444 (N_28444,N_27593,N_27190);
xnor U28445 (N_28445,N_27516,N_27984);
or U28446 (N_28446,N_27646,N_27998);
nand U28447 (N_28447,N_27201,N_27519);
nand U28448 (N_28448,N_27618,N_26420);
and U28449 (N_28449,N_26582,N_26661);
or U28450 (N_28450,N_26453,N_27619);
nand U28451 (N_28451,N_26685,N_26874);
or U28452 (N_28452,N_27895,N_27823);
or U28453 (N_28453,N_27902,N_26975);
and U28454 (N_28454,N_26829,N_27863);
xnor U28455 (N_28455,N_27878,N_27300);
and U28456 (N_28456,N_27603,N_26170);
and U28457 (N_28457,N_26682,N_26448);
and U28458 (N_28458,N_27191,N_26710);
and U28459 (N_28459,N_27464,N_27707);
and U28460 (N_28460,N_26468,N_27027);
or U28461 (N_28461,N_26132,N_27075);
and U28462 (N_28462,N_26138,N_27851);
or U28463 (N_28463,N_26447,N_26800);
nor U28464 (N_28464,N_26250,N_26443);
xor U28465 (N_28465,N_27184,N_27883);
nor U28466 (N_28466,N_26635,N_26326);
xor U28467 (N_28467,N_27124,N_27172);
nor U28468 (N_28468,N_26531,N_26396);
nand U28469 (N_28469,N_26650,N_27025);
and U28470 (N_28470,N_26067,N_27319);
xor U28471 (N_28471,N_27310,N_27401);
or U28472 (N_28472,N_26514,N_26456);
nand U28473 (N_28473,N_26799,N_26299);
or U28474 (N_28474,N_26452,N_27653);
xor U28475 (N_28475,N_27399,N_26339);
nand U28476 (N_28476,N_27839,N_26300);
nand U28477 (N_28477,N_27896,N_27845);
nand U28478 (N_28478,N_26025,N_27041);
or U28479 (N_28479,N_26478,N_27518);
xor U28480 (N_28480,N_27026,N_26057);
nor U28481 (N_28481,N_26206,N_27494);
xor U28482 (N_28482,N_27994,N_26703);
nand U28483 (N_28483,N_27737,N_27344);
xnor U28484 (N_28484,N_26923,N_26257);
nand U28485 (N_28485,N_26145,N_26974);
nand U28486 (N_28486,N_26973,N_26708);
nand U28487 (N_28487,N_26702,N_26432);
or U28488 (N_28488,N_27739,N_26402);
or U28489 (N_28489,N_27592,N_26688);
nor U28490 (N_28490,N_27293,N_26106);
or U28491 (N_28491,N_27742,N_27162);
xor U28492 (N_28492,N_27260,N_26993);
nor U28493 (N_28493,N_27931,N_27789);
xnor U28494 (N_28494,N_26237,N_27805);
and U28495 (N_28495,N_27362,N_27018);
nor U28496 (N_28496,N_26601,N_26713);
nor U28497 (N_28497,N_27649,N_26640);
and U28498 (N_28498,N_26959,N_27560);
or U28499 (N_28499,N_27578,N_26436);
xor U28500 (N_28500,N_27514,N_27836);
xnor U28501 (N_28501,N_26605,N_26794);
and U28502 (N_28502,N_26210,N_26563);
and U28503 (N_28503,N_26667,N_27504);
nor U28504 (N_28504,N_26760,N_27719);
nor U28505 (N_28505,N_26278,N_26976);
or U28506 (N_28506,N_26739,N_27232);
xor U28507 (N_28507,N_27187,N_26991);
nand U28508 (N_28508,N_26459,N_26784);
nand U28509 (N_28509,N_27140,N_26828);
xor U28510 (N_28510,N_26212,N_26511);
and U28511 (N_28511,N_27392,N_27715);
and U28512 (N_28512,N_26579,N_27612);
xnor U28513 (N_28513,N_27997,N_26790);
xor U28514 (N_28514,N_26412,N_26859);
nor U28515 (N_28515,N_26818,N_26115);
and U28516 (N_28516,N_26407,N_27457);
xnor U28517 (N_28517,N_27840,N_26366);
nand U28518 (N_28518,N_26242,N_27179);
or U28519 (N_28519,N_27178,N_26998);
or U28520 (N_28520,N_27470,N_26897);
and U28521 (N_28521,N_26105,N_26699);
nand U28522 (N_28522,N_27044,N_27856);
or U28523 (N_28523,N_27733,N_26356);
nand U28524 (N_28524,N_27552,N_27690);
and U28525 (N_28525,N_27312,N_26469);
nand U28526 (N_28526,N_26927,N_27278);
and U28527 (N_28527,N_26369,N_27441);
or U28528 (N_28528,N_27600,N_26801);
or U28529 (N_28529,N_26523,N_26120);
nand U28530 (N_28530,N_26177,N_26798);
xnor U28531 (N_28531,N_26670,N_26264);
nand U28532 (N_28532,N_27043,N_27317);
and U28533 (N_28533,N_26594,N_27622);
and U28534 (N_28534,N_26577,N_26006);
nand U28535 (N_28535,N_27093,N_26081);
nor U28536 (N_28536,N_26041,N_26606);
xnor U28537 (N_28537,N_27999,N_26665);
nand U28538 (N_28538,N_26484,N_26908);
and U28539 (N_28539,N_27922,N_26905);
nor U28540 (N_28540,N_27398,N_26920);
nand U28541 (N_28541,N_27882,N_26308);
and U28542 (N_28542,N_27081,N_26251);
and U28543 (N_28543,N_27315,N_26691);
nand U28544 (N_28544,N_26256,N_26165);
nand U28545 (N_28545,N_26293,N_27825);
nand U28546 (N_28546,N_27455,N_26163);
or U28547 (N_28547,N_26146,N_26692);
nand U28548 (N_28548,N_27328,N_27979);
nor U28549 (N_28549,N_26173,N_26466);
and U28550 (N_28550,N_27327,N_26642);
nor U28551 (N_28551,N_27774,N_26046);
nor U28552 (N_28552,N_26491,N_26673);
nor U28553 (N_28553,N_27567,N_27654);
and U28554 (N_28554,N_26894,N_26274);
nor U28555 (N_28555,N_26433,N_26062);
xnor U28556 (N_28556,N_26134,N_27674);
nand U28557 (N_28557,N_26223,N_26390);
xnor U28558 (N_28558,N_26408,N_27438);
or U28559 (N_28559,N_26953,N_27142);
nand U28560 (N_28560,N_26381,N_27829);
xnor U28561 (N_28561,N_27094,N_27114);
nand U28562 (N_28562,N_27911,N_27146);
or U28563 (N_28563,N_27348,N_27411);
nand U28564 (N_28564,N_26095,N_26844);
xnor U28565 (N_28565,N_26424,N_27467);
nand U28566 (N_28566,N_27699,N_26896);
nor U28567 (N_28567,N_27506,N_27063);
and U28568 (N_28568,N_26188,N_26204);
nor U28569 (N_28569,N_27456,N_26529);
nand U28570 (N_28570,N_26824,N_26949);
and U28571 (N_28571,N_26327,N_27015);
nor U28572 (N_28572,N_26160,N_26200);
nand U28573 (N_28573,N_26572,N_26240);
and U28574 (N_28574,N_27890,N_27120);
xor U28575 (N_28575,N_27082,N_27617);
or U28576 (N_28576,N_26751,N_26811);
nor U28577 (N_28577,N_26745,N_27247);
xnor U28578 (N_28578,N_27117,N_26398);
nand U28579 (N_28579,N_27087,N_26720);
or U28580 (N_28580,N_26671,N_27950);
or U28581 (N_28581,N_26435,N_27415);
nand U28582 (N_28582,N_27499,N_27092);
or U28583 (N_28583,N_27797,N_27035);
and U28584 (N_28584,N_27978,N_27020);
xor U28585 (N_28585,N_26540,N_26989);
or U28586 (N_28586,N_27065,N_26627);
xor U28587 (N_28587,N_26560,N_27522);
nand U28588 (N_28588,N_27601,N_27046);
nor U28589 (N_28589,N_27843,N_27668);
and U28590 (N_28590,N_26633,N_26766);
or U28591 (N_28591,N_27796,N_27628);
or U28592 (N_28592,N_27680,N_26222);
xnor U28593 (N_28593,N_27577,N_27444);
nor U28594 (N_28594,N_26303,N_27149);
nor U28595 (N_28595,N_26495,N_26636);
nor U28596 (N_28596,N_26282,N_26345);
nor U28597 (N_28597,N_26987,N_26365);
xnor U28598 (N_28598,N_27353,N_26475);
nor U28599 (N_28599,N_27048,N_26322);
and U28600 (N_28600,N_26205,N_27028);
nor U28601 (N_28601,N_26711,N_27377);
and U28602 (N_28602,N_27585,N_27476);
and U28603 (N_28603,N_26584,N_27581);
nand U28604 (N_28604,N_27274,N_26822);
nor U28605 (N_28605,N_26626,N_26580);
and U28606 (N_28606,N_26632,N_26817);
nor U28607 (N_28607,N_27970,N_26676);
xnor U28608 (N_28608,N_26371,N_26400);
nor U28609 (N_28609,N_27915,N_26335);
and U28610 (N_28610,N_27143,N_26994);
xor U28611 (N_28611,N_27272,N_27620);
nand U28612 (N_28612,N_26683,N_26142);
and U28613 (N_28613,N_26208,N_26474);
xor U28614 (N_28614,N_27685,N_26252);
nand U28615 (N_28615,N_27996,N_26018);
nand U28616 (N_28616,N_26384,N_27440);
xnor U28617 (N_28617,N_27241,N_26239);
or U28618 (N_28618,N_27788,N_27380);
xnor U28619 (N_28619,N_27139,N_26857);
or U28620 (N_28620,N_26931,N_27854);
nand U28621 (N_28621,N_26112,N_27198);
nor U28622 (N_28622,N_26793,N_27403);
or U28623 (N_28623,N_27662,N_27500);
xnor U28624 (N_28624,N_26516,N_26302);
or U28625 (N_28625,N_27875,N_27976);
and U28626 (N_28626,N_26555,N_27664);
and U28627 (N_28627,N_27547,N_26023);
or U28628 (N_28628,N_27870,N_26561);
xor U28629 (N_28629,N_26780,N_27479);
nand U28630 (N_28630,N_27287,N_27052);
or U28631 (N_28631,N_27793,N_27566);
xor U28632 (N_28632,N_27523,N_27527);
nor U28633 (N_28633,N_27480,N_27666);
and U28634 (N_28634,N_27505,N_27528);
nand U28635 (N_28635,N_27910,N_27031);
nand U28636 (N_28636,N_27090,N_26590);
and U28637 (N_28637,N_27194,N_26284);
nor U28638 (N_28638,N_26610,N_27069);
and U28639 (N_28639,N_26515,N_26885);
xor U28640 (N_28640,N_26726,N_26820);
or U28641 (N_28641,N_27676,N_26616);
or U28642 (N_28642,N_26055,N_27761);
or U28643 (N_28643,N_27433,N_26863);
and U28644 (N_28644,N_27780,N_27549);
and U28645 (N_28645,N_27708,N_26508);
nor U28646 (N_28646,N_27801,N_26771);
nor U28647 (N_28647,N_27202,N_27302);
nand U28648 (N_28648,N_27673,N_26806);
xnor U28649 (N_28649,N_26714,N_27561);
or U28650 (N_28650,N_26728,N_27995);
xnor U28651 (N_28651,N_27417,N_27595);
nand U28652 (N_28652,N_27867,N_27624);
nor U28653 (N_28653,N_26045,N_26669);
and U28654 (N_28654,N_27255,N_26196);
nor U28655 (N_28655,N_27941,N_27709);
and U28656 (N_28656,N_27583,N_27810);
xnor U28657 (N_28657,N_26323,N_27396);
nor U28658 (N_28658,N_26639,N_26493);
nor U28659 (N_28659,N_27919,N_26741);
xor U28660 (N_28660,N_27675,N_27688);
nor U28661 (N_28661,N_27652,N_27332);
or U28662 (N_28662,N_26507,N_27886);
xor U28663 (N_28663,N_26840,N_27751);
and U28664 (N_28664,N_27054,N_27175);
or U28665 (N_28665,N_26487,N_27490);
nand U28666 (N_28666,N_27119,N_26532);
nand U28667 (N_28667,N_26090,N_26460);
nand U28668 (N_28668,N_27346,N_27121);
and U28669 (N_28669,N_26352,N_27437);
xor U28670 (N_28670,N_26261,N_27753);
nor U28671 (N_28671,N_26093,N_27153);
nor U28672 (N_28672,N_27066,N_26946);
and U28673 (N_28673,N_26654,N_27669);
nor U28674 (N_28674,N_27446,N_27359);
xnor U28675 (N_28675,N_26694,N_27323);
nand U28676 (N_28676,N_27711,N_26747);
nor U28677 (N_28677,N_26748,N_27221);
xnor U28678 (N_28678,N_26164,N_27071);
or U28679 (N_28679,N_26122,N_26888);
nand U28680 (N_28680,N_27390,N_27746);
and U28681 (N_28681,N_26316,N_27686);
nor U28682 (N_28682,N_26759,N_26933);
nand U28683 (N_28683,N_27828,N_27358);
nor U28684 (N_28684,N_26684,N_27418);
and U28685 (N_28685,N_27458,N_26000);
and U28686 (N_28686,N_26235,N_27971);
and U28687 (N_28687,N_26612,N_26543);
nand U28688 (N_28688,N_27795,N_26717);
or U28689 (N_28689,N_26141,N_26007);
nand U28690 (N_28690,N_26332,N_27588);
xor U28691 (N_28691,N_26965,N_27145);
nor U28692 (N_28692,N_27096,N_27360);
nor U28693 (N_28693,N_27866,N_27222);
xor U28694 (N_28694,N_27928,N_27454);
nand U28695 (N_28695,N_27713,N_27968);
nor U28696 (N_28696,N_26724,N_26656);
xor U28697 (N_28697,N_26860,N_27361);
nor U28698 (N_28698,N_27958,N_26910);
and U28699 (N_28699,N_26175,N_26607);
xor U28700 (N_28700,N_27240,N_26812);
nand U28701 (N_28701,N_26065,N_27754);
or U28702 (N_28702,N_26743,N_26663);
xnor U28703 (N_28703,N_26346,N_26853);
xor U28704 (N_28704,N_26108,N_27764);
or U28705 (N_28705,N_27414,N_26735);
xor U28706 (N_28706,N_27343,N_26611);
and U28707 (N_28707,N_27180,N_27897);
nor U28708 (N_28708,N_26833,N_27893);
nand U28709 (N_28709,N_27283,N_27934);
or U28710 (N_28710,N_26043,N_26596);
nor U28711 (N_28711,N_26554,N_26129);
nand U28712 (N_28712,N_26119,N_26876);
and U28713 (N_28713,N_26351,N_27330);
xnor U28714 (N_28714,N_27388,N_26388);
xnor U28715 (N_28715,N_27862,N_26869);
or U28716 (N_28716,N_27185,N_26831);
or U28717 (N_28717,N_27517,N_27616);
nand U28718 (N_28718,N_26795,N_27572);
nand U28719 (N_28719,N_27372,N_26574);
or U28720 (N_28720,N_27442,N_26777);
or U28721 (N_28721,N_27105,N_26434);
nand U28722 (N_28722,N_26902,N_26878);
and U28723 (N_28723,N_26047,N_27880);
and U28724 (N_28724,N_26418,N_27948);
nor U28725 (N_28725,N_26417,N_27570);
or U28726 (N_28726,N_26544,N_26715);
and U28727 (N_28727,N_26718,N_26881);
nand U28728 (N_28728,N_26191,N_27672);
nand U28729 (N_28729,N_26362,N_27626);
xor U28730 (N_28730,N_27176,N_27435);
nor U28731 (N_28731,N_27334,N_26254);
and U28732 (N_28732,N_27473,N_26845);
xnor U28733 (N_28733,N_26539,N_26034);
nand U28734 (N_28734,N_27881,N_26294);
nor U28735 (N_28735,N_27607,N_26099);
or U28736 (N_28736,N_27386,N_26618);
nor U28737 (N_28737,N_26458,N_26525);
or U28738 (N_28738,N_26312,N_27004);
nand U28739 (N_28739,N_26354,N_26945);
and U28740 (N_28740,N_26364,N_26003);
xor U28741 (N_28741,N_27785,N_27689);
or U28742 (N_28742,N_27757,N_27428);
nand U28743 (N_28743,N_26246,N_27947);
xor U28744 (N_28744,N_27985,N_27957);
xor U28745 (N_28745,N_26763,N_27076);
nand U28746 (N_28746,N_26036,N_26506);
xnor U28747 (N_28747,N_27536,N_27193);
and U28748 (N_28748,N_26681,N_27602);
or U28749 (N_28749,N_27200,N_26051);
and U28750 (N_28750,N_27605,N_26378);
nor U28751 (N_28751,N_26053,N_27631);
or U28752 (N_28752,N_27826,N_27370);
or U28753 (N_28753,N_27484,N_27099);
xnor U28754 (N_28754,N_26076,N_27182);
nor U28755 (N_28755,N_26697,N_27894);
nor U28756 (N_28756,N_26419,N_26700);
nand U28757 (N_28757,N_26227,N_27842);
or U28758 (N_28758,N_27712,N_27725);
and U28759 (N_28759,N_27251,N_26630);
xor U28760 (N_28760,N_26318,N_26290);
or U28761 (N_28761,N_26870,N_27034);
nor U28762 (N_28762,N_26130,N_27704);
nand U28763 (N_28763,N_27752,N_27898);
or U28764 (N_28764,N_26749,N_26189);
or U28765 (N_28765,N_27347,N_26113);
and U28766 (N_28766,N_26324,N_26270);
nor U28767 (N_28767,N_26834,N_26541);
and U28768 (N_28768,N_27508,N_27166);
nand U28769 (N_28769,N_27525,N_27822);
and U28770 (N_28770,N_26485,N_27551);
nor U28771 (N_28771,N_26008,N_27425);
and U28772 (N_28772,N_26537,N_26273);
or U28773 (N_28773,N_26234,N_27192);
or U28774 (N_28774,N_26309,N_27794);
or U28775 (N_28775,N_26068,N_26224);
nand U28776 (N_28776,N_27812,N_27738);
xnor U28777 (N_28777,N_26140,N_26197);
xnor U28778 (N_28778,N_26263,N_26979);
or U28779 (N_28779,N_27248,N_26781);
xor U28780 (N_28780,N_27938,N_26553);
nand U28781 (N_28781,N_26102,N_27714);
nand U28782 (N_28782,N_27921,N_27183);
nand U28783 (N_28783,N_26980,N_27945);
nand U28784 (N_28784,N_27969,N_27501);
and U28785 (N_28785,N_27336,N_26657);
nand U28786 (N_28786,N_27936,N_26277);
or U28787 (N_28787,N_26026,N_26599);
nor U28788 (N_28788,N_27084,N_26826);
and U28789 (N_28789,N_27266,N_26758);
nand U28790 (N_28790,N_26919,N_26219);
xnor U28791 (N_28791,N_27393,N_27257);
or U28792 (N_28792,N_27526,N_26446);
nor U28793 (N_28793,N_27112,N_27546);
or U28794 (N_28794,N_27981,N_27338);
nand U28795 (N_28795,N_27261,N_27357);
nor U28796 (N_28796,N_27281,N_26709);
nor U28797 (N_28797,N_26211,N_27156);
or U28798 (N_28798,N_27939,N_26178);
nor U28799 (N_28799,N_27642,N_26848);
or U28800 (N_28800,N_27756,N_27817);
xnor U28801 (N_28801,N_26330,N_26451);
or U28802 (N_28802,N_26187,N_26705);
xor U28803 (N_28803,N_26128,N_27877);
nand U28804 (N_28804,N_27558,N_26103);
xnor U28805 (N_28805,N_27001,N_27865);
nand U28806 (N_28806,N_26904,N_27158);
and U28807 (N_28807,N_27809,N_26803);
nor U28808 (N_28808,N_26202,N_26969);
nor U28809 (N_28809,N_27650,N_27292);
xnor U28810 (N_28810,N_26730,N_26203);
or U28811 (N_28811,N_27436,N_26135);
nor U28812 (N_28812,N_26292,N_26079);
and U28813 (N_28813,N_27169,N_27279);
xnor U28814 (N_28814,N_27943,N_26955);
xnor U28815 (N_28815,N_26583,N_26325);
xor U28816 (N_28816,N_27322,N_27064);
or U28817 (N_28817,N_27280,N_26198);
or U28818 (N_28818,N_26603,N_27269);
and U28819 (N_28819,N_27944,N_26276);
xnor U28820 (N_28820,N_27029,N_27369);
or U28821 (N_28821,N_27530,N_26226);
nand U28822 (N_28822,N_27961,N_26230);
nor U28823 (N_28823,N_27681,N_26367);
and U28824 (N_28824,N_26295,N_26073);
nand U28825 (N_28825,N_26805,N_27584);
nand U28826 (N_28826,N_26131,N_27559);
xnor U28827 (N_28827,N_27234,N_27806);
or U28828 (N_28828,N_27130,N_26125);
and U28829 (N_28829,N_26355,N_27061);
xor U28830 (N_28830,N_26858,N_26050);
or U28831 (N_28831,N_26767,N_27767);
xor U28832 (N_28832,N_27217,N_26879);
nand U28833 (N_28833,N_26377,N_27475);
xnor U28834 (N_28834,N_26742,N_26385);
nor U28835 (N_28835,N_26680,N_26964);
and U28836 (N_28836,N_27326,N_26394);
and U28837 (N_28837,N_27821,N_27126);
and U28838 (N_28838,N_27734,N_27967);
nor U28839 (N_28839,N_26891,N_26249);
nand U28840 (N_28840,N_27448,N_27635);
or U28841 (N_28841,N_26075,N_26078);
or U28842 (N_28842,N_27590,N_26348);
nand U28843 (N_28843,N_26423,N_27005);
xor U28844 (N_28844,N_27445,N_27144);
or U28845 (N_28845,N_27860,N_27102);
xnor U28846 (N_28846,N_26037,N_27906);
and U28847 (N_28847,N_26791,N_27853);
xnor U28848 (N_28848,N_27373,N_26847);
and U28849 (N_28849,N_26526,N_27109);
and U28850 (N_28850,N_27889,N_26013);
nand U28851 (N_28851,N_26939,N_27186);
nor U28852 (N_28852,N_27045,N_26567);
and U28853 (N_28853,N_26114,N_26463);
xnor U28854 (N_28854,N_27548,N_26823);
xor U28855 (N_28855,N_27876,N_26340);
xor U28856 (N_28856,N_26873,N_27589);
nand U28857 (N_28857,N_26228,N_26494);
and U28858 (N_28858,N_26072,N_26997);
xor U28859 (N_28859,N_27924,N_27017);
nor U28860 (N_28860,N_27089,N_26358);
nor U28861 (N_28861,N_26559,N_27760);
nand U28862 (N_28862,N_26719,N_26957);
nand U28863 (N_28863,N_27296,N_26875);
nand U28864 (N_28864,N_27610,N_26248);
xor U28865 (N_28865,N_26104,N_26031);
xnor U28866 (N_28866,N_26782,N_27671);
nor U28867 (N_28867,N_26157,N_27597);
xnor U28868 (N_28868,N_26872,N_27132);
nand U28869 (N_28869,N_27917,N_27412);
and U28870 (N_28870,N_26967,N_27273);
or U28871 (N_28871,N_26825,N_26813);
or U28872 (N_28872,N_27512,N_27039);
or U28873 (N_28873,N_26071,N_26677);
or U28874 (N_28874,N_26674,N_27231);
xor U28875 (N_28875,N_27088,N_27170);
and U28876 (N_28876,N_27270,N_26232);
or U28877 (N_28877,N_27304,N_27271);
and U28878 (N_28878,N_26546,N_26613);
nor U28879 (N_28879,N_26638,N_26479);
xnor U28880 (N_28880,N_27731,N_26617);
xnor U28881 (N_28881,N_27747,N_27724);
xor U28882 (N_28882,N_27813,N_27700);
or U28883 (N_28883,N_26027,N_26238);
or U28884 (N_28884,N_26464,N_27154);
xor U28885 (N_28885,N_27205,N_27405);
xor U28886 (N_28886,N_27852,N_27884);
nand U28887 (N_28887,N_26796,N_27086);
xnor U28888 (N_28888,N_26783,N_27049);
xnor U28889 (N_28889,N_26932,N_27181);
or U28890 (N_28890,N_27318,N_26562);
nand U28891 (N_28891,N_26373,N_27498);
xnor U28892 (N_28892,N_27771,N_26658);
nand U28893 (N_28893,N_27349,N_27101);
nand U28894 (N_28894,N_27974,N_26503);
and U28895 (N_28895,N_27107,N_26382);
or U28896 (N_28896,N_27354,N_26336);
nor U28897 (N_28897,N_27007,N_27011);
nand U28898 (N_28898,N_27189,N_27197);
xor U28899 (N_28899,N_27665,N_26289);
or U28900 (N_28900,N_27932,N_26269);
and U28901 (N_28901,N_26792,N_27531);
xor U28902 (N_28902,N_26624,N_27550);
nand U28903 (N_28903,N_26756,N_26647);
nand U28904 (N_28904,N_26917,N_27371);
nand U28905 (N_28905,N_27410,N_27254);
and U28906 (N_28906,N_27237,N_26581);
and U28907 (N_28907,N_27163,N_27556);
and U28908 (N_28908,N_26660,N_26944);
nand U28909 (N_28909,N_26350,N_26060);
nor U28910 (N_28910,N_27024,N_27824);
or U28911 (N_28911,N_27262,N_26098);
or U28912 (N_28912,N_26524,N_26029);
nand U28913 (N_28913,N_27509,N_26116);
xor U28914 (N_28914,N_26179,N_26592);
xnor U28915 (N_28915,N_26883,N_27195);
nand U28916 (N_28916,N_27916,N_27223);
or U28917 (N_28917,N_27965,N_27284);
nand U28918 (N_28918,N_26489,N_27891);
xnor U28919 (N_28919,N_26272,N_27977);
nand U28920 (N_28920,N_26988,N_26430);
nand U28921 (N_28921,N_27925,N_26283);
nand U28922 (N_28922,N_27228,N_26542);
and U28923 (N_28923,N_27077,N_27750);
nor U28924 (N_28924,N_27367,N_26707);
nor U28925 (N_28925,N_26520,N_26815);
nor U28926 (N_28926,N_26158,N_27291);
or U28927 (N_28927,N_27013,N_27571);
nor U28928 (N_28928,N_27540,N_27306);
and U28929 (N_28929,N_27127,N_26914);
and U28930 (N_28930,N_27236,N_27277);
nor U28931 (N_28931,N_27741,N_26644);
and U28932 (N_28932,N_27356,N_26849);
and U28933 (N_28933,N_27614,N_26838);
nor U28934 (N_28934,N_26401,N_26059);
nor U28935 (N_28935,N_27252,N_26668);
nand U28936 (N_28936,N_27679,N_27946);
and U28937 (N_28937,N_27692,N_26961);
nand U28938 (N_28938,N_27067,N_27918);
or U28939 (N_28939,N_26695,N_27710);
and U28940 (N_28940,N_27615,N_26928);
or U28941 (N_28941,N_27625,N_27085);
nand U28942 (N_28942,N_26149,N_27586);
or U28943 (N_28943,N_26331,N_26033);
nand U28944 (N_28944,N_26262,N_26209);
nand U28945 (N_28945,N_26721,N_27352);
and U28946 (N_28946,N_26773,N_27802);
nand U28947 (N_28947,N_26678,N_27933);
and U28948 (N_28948,N_27903,N_27381);
and U28949 (N_28949,N_26779,N_26126);
nand U28950 (N_28950,N_26038,N_27511);
or U28951 (N_28951,N_26471,N_26044);
xor U28952 (N_28952,N_27305,N_26012);
or U28953 (N_28953,N_27125,N_27992);
nor U28954 (N_28954,N_26137,N_26968);
nand U28955 (N_28955,N_26190,N_26169);
and U28956 (N_28956,N_26768,N_27138);
nor U28957 (N_28957,N_27799,N_27000);
and U28958 (N_28958,N_27196,N_27230);
and U28959 (N_28959,N_27987,N_26009);
nand U28960 (N_28960,N_26123,N_26258);
nor U28961 (N_28961,N_26315,N_26159);
xor U28962 (N_28962,N_27021,N_26521);
or U28963 (N_28963,N_26310,N_26216);
and U28964 (N_28964,N_26960,N_27421);
nand U28965 (N_28965,N_26690,N_27723);
nand U28966 (N_28966,N_27574,N_27303);
xor U28967 (N_28967,N_27282,N_26422);
nand U28968 (N_28968,N_26675,N_26557);
or U28969 (N_28969,N_26375,N_26704);
nand U28970 (N_28970,N_27575,N_26476);
and U28971 (N_28971,N_27972,N_26625);
and U28972 (N_28972,N_27321,N_27226);
nor U28973 (N_28973,N_27122,N_26010);
nor U28974 (N_28974,N_27568,N_26172);
and U28975 (N_28975,N_27784,N_26470);
nor U28976 (N_28976,N_26214,N_26871);
nor U28977 (N_28977,N_26497,N_26056);
nor U28978 (N_28978,N_26376,N_27276);
or U28979 (N_28979,N_26101,N_27777);
or U28980 (N_28980,N_26772,N_26570);
nor U28981 (N_28981,N_26548,N_26990);
xor U28982 (N_28982,N_26082,N_27634);
and U28983 (N_28983,N_27012,N_27363);
nor U28984 (N_28984,N_27608,N_27108);
nor U28985 (N_28985,N_26664,N_27544);
nand U28986 (N_28986,N_27468,N_26298);
nand U28987 (N_28987,N_26022,N_27265);
xnor U28988 (N_28988,N_27238,N_26004);
and U28989 (N_28989,N_27482,N_26970);
xor U28990 (N_28990,N_27208,N_27106);
nand U28991 (N_28991,N_27342,N_27956);
nor U28992 (N_28992,N_26797,N_26576);
xnor U28993 (N_28993,N_27426,N_27841);
nor U28994 (N_28994,N_27450,N_26501);
and U28995 (N_28995,N_26645,N_27211);
nand U28996 (N_28996,N_26804,N_26074);
xnor U28997 (N_28997,N_27503,N_27443);
xor U28998 (N_28998,N_26054,N_26948);
or U28999 (N_28999,N_26528,N_26589);
nand U29000 (N_29000,N_26364,N_26946);
xor U29001 (N_29001,N_27035,N_27196);
or U29002 (N_29002,N_27883,N_27974);
or U29003 (N_29003,N_27323,N_27170);
xor U29004 (N_29004,N_26592,N_26585);
xnor U29005 (N_29005,N_26591,N_27526);
nand U29006 (N_29006,N_26521,N_26250);
or U29007 (N_29007,N_27582,N_26837);
or U29008 (N_29008,N_27152,N_27885);
nor U29009 (N_29009,N_27024,N_26870);
and U29010 (N_29010,N_26399,N_26349);
nand U29011 (N_29011,N_26865,N_26360);
and U29012 (N_29012,N_26192,N_27014);
nand U29013 (N_29013,N_27681,N_26900);
xor U29014 (N_29014,N_27736,N_27582);
or U29015 (N_29015,N_27489,N_26796);
nand U29016 (N_29016,N_26251,N_26439);
or U29017 (N_29017,N_27801,N_26385);
xnor U29018 (N_29018,N_27714,N_27476);
and U29019 (N_29019,N_27636,N_27535);
and U29020 (N_29020,N_26430,N_26249);
and U29021 (N_29021,N_26357,N_26506);
nor U29022 (N_29022,N_26529,N_26442);
nor U29023 (N_29023,N_26995,N_26300);
nand U29024 (N_29024,N_27051,N_27832);
or U29025 (N_29025,N_27987,N_27201);
and U29026 (N_29026,N_26777,N_26450);
and U29027 (N_29027,N_27191,N_26208);
or U29028 (N_29028,N_27179,N_27653);
and U29029 (N_29029,N_27442,N_26865);
or U29030 (N_29030,N_27416,N_27829);
xor U29031 (N_29031,N_26808,N_27087);
nor U29032 (N_29032,N_27874,N_26620);
and U29033 (N_29033,N_26962,N_27426);
nor U29034 (N_29034,N_27133,N_26429);
and U29035 (N_29035,N_26992,N_27357);
nor U29036 (N_29036,N_26462,N_27340);
nor U29037 (N_29037,N_26430,N_27499);
nor U29038 (N_29038,N_27710,N_26185);
xor U29039 (N_29039,N_27968,N_26025);
xnor U29040 (N_29040,N_27994,N_26943);
or U29041 (N_29041,N_27223,N_26665);
xor U29042 (N_29042,N_27703,N_26601);
xnor U29043 (N_29043,N_27730,N_27003);
or U29044 (N_29044,N_27340,N_26603);
and U29045 (N_29045,N_26991,N_27927);
xnor U29046 (N_29046,N_27448,N_26476);
or U29047 (N_29047,N_27734,N_26041);
nand U29048 (N_29048,N_26045,N_27759);
nand U29049 (N_29049,N_26455,N_27931);
nand U29050 (N_29050,N_26046,N_26905);
or U29051 (N_29051,N_27071,N_26064);
and U29052 (N_29052,N_26788,N_26079);
xnor U29053 (N_29053,N_26714,N_27583);
nor U29054 (N_29054,N_27729,N_27255);
or U29055 (N_29055,N_27373,N_26653);
nand U29056 (N_29056,N_27392,N_27564);
xor U29057 (N_29057,N_26125,N_26116);
or U29058 (N_29058,N_26612,N_27524);
or U29059 (N_29059,N_27022,N_26997);
xnor U29060 (N_29060,N_26075,N_26412);
nand U29061 (N_29061,N_26024,N_26673);
xnor U29062 (N_29062,N_27775,N_27561);
nor U29063 (N_29063,N_27234,N_26006);
xor U29064 (N_29064,N_26782,N_26520);
nand U29065 (N_29065,N_27474,N_27868);
nor U29066 (N_29066,N_27914,N_26617);
xnor U29067 (N_29067,N_26837,N_26087);
or U29068 (N_29068,N_27748,N_27781);
nand U29069 (N_29069,N_27791,N_27776);
xnor U29070 (N_29070,N_26822,N_27626);
and U29071 (N_29071,N_26787,N_27466);
nand U29072 (N_29072,N_27385,N_27659);
or U29073 (N_29073,N_26603,N_26588);
or U29074 (N_29074,N_26562,N_27125);
nor U29075 (N_29075,N_26798,N_27142);
or U29076 (N_29076,N_27020,N_27846);
or U29077 (N_29077,N_26822,N_26133);
nor U29078 (N_29078,N_27139,N_27022);
and U29079 (N_29079,N_27400,N_27876);
and U29080 (N_29080,N_26231,N_26271);
or U29081 (N_29081,N_27215,N_26814);
nor U29082 (N_29082,N_26519,N_26683);
and U29083 (N_29083,N_27343,N_26341);
nor U29084 (N_29084,N_27890,N_26792);
nand U29085 (N_29085,N_27490,N_26702);
nor U29086 (N_29086,N_27441,N_27568);
nor U29087 (N_29087,N_27532,N_27226);
and U29088 (N_29088,N_27459,N_26408);
xnor U29089 (N_29089,N_27151,N_26598);
nand U29090 (N_29090,N_27141,N_26832);
or U29091 (N_29091,N_26909,N_27503);
and U29092 (N_29092,N_26299,N_26466);
and U29093 (N_29093,N_26332,N_27129);
xnor U29094 (N_29094,N_27914,N_27748);
nand U29095 (N_29095,N_27382,N_27774);
nand U29096 (N_29096,N_27031,N_27045);
and U29097 (N_29097,N_27926,N_26649);
nand U29098 (N_29098,N_26845,N_27560);
xor U29099 (N_29099,N_27014,N_27881);
nand U29100 (N_29100,N_26902,N_26830);
xnor U29101 (N_29101,N_26757,N_27609);
nand U29102 (N_29102,N_26923,N_27726);
nand U29103 (N_29103,N_27381,N_26445);
and U29104 (N_29104,N_27489,N_26547);
xor U29105 (N_29105,N_27700,N_27763);
and U29106 (N_29106,N_26690,N_27438);
and U29107 (N_29107,N_26451,N_27599);
xnor U29108 (N_29108,N_27952,N_26588);
and U29109 (N_29109,N_27240,N_27541);
and U29110 (N_29110,N_26013,N_27668);
xor U29111 (N_29111,N_26383,N_27189);
nand U29112 (N_29112,N_26561,N_27459);
nand U29113 (N_29113,N_27761,N_26476);
or U29114 (N_29114,N_27154,N_27223);
or U29115 (N_29115,N_27191,N_26175);
nand U29116 (N_29116,N_27119,N_27737);
and U29117 (N_29117,N_26550,N_27622);
nor U29118 (N_29118,N_27061,N_26290);
nand U29119 (N_29119,N_27992,N_26172);
nor U29120 (N_29120,N_26150,N_27974);
or U29121 (N_29121,N_26289,N_27011);
nand U29122 (N_29122,N_27304,N_26521);
nor U29123 (N_29123,N_27947,N_26605);
nand U29124 (N_29124,N_27496,N_27284);
xnor U29125 (N_29125,N_26831,N_27780);
nor U29126 (N_29126,N_26724,N_27437);
or U29127 (N_29127,N_27930,N_27853);
xor U29128 (N_29128,N_27419,N_26550);
nor U29129 (N_29129,N_26744,N_26252);
xor U29130 (N_29130,N_26446,N_26468);
nor U29131 (N_29131,N_26791,N_27812);
nor U29132 (N_29132,N_26828,N_27522);
or U29133 (N_29133,N_27256,N_27234);
or U29134 (N_29134,N_27100,N_26486);
nor U29135 (N_29135,N_27798,N_26670);
or U29136 (N_29136,N_26176,N_27103);
nor U29137 (N_29137,N_26907,N_26397);
nand U29138 (N_29138,N_27854,N_27300);
and U29139 (N_29139,N_27646,N_27664);
or U29140 (N_29140,N_26561,N_26848);
xor U29141 (N_29141,N_26235,N_27302);
and U29142 (N_29142,N_26874,N_26852);
and U29143 (N_29143,N_27690,N_27799);
nand U29144 (N_29144,N_26320,N_27283);
nor U29145 (N_29145,N_27322,N_26630);
nor U29146 (N_29146,N_27623,N_27204);
and U29147 (N_29147,N_27821,N_27595);
nor U29148 (N_29148,N_26052,N_26449);
or U29149 (N_29149,N_27085,N_26669);
nand U29150 (N_29150,N_26474,N_27374);
xor U29151 (N_29151,N_26579,N_27586);
and U29152 (N_29152,N_26137,N_26896);
or U29153 (N_29153,N_26165,N_27904);
nor U29154 (N_29154,N_26285,N_27657);
nor U29155 (N_29155,N_26095,N_26507);
and U29156 (N_29156,N_27169,N_26263);
and U29157 (N_29157,N_26362,N_26188);
nor U29158 (N_29158,N_27279,N_27164);
xnor U29159 (N_29159,N_26644,N_27643);
nand U29160 (N_29160,N_26512,N_27452);
or U29161 (N_29161,N_27090,N_26153);
and U29162 (N_29162,N_26587,N_27099);
xor U29163 (N_29163,N_26890,N_27441);
and U29164 (N_29164,N_26708,N_26942);
or U29165 (N_29165,N_26829,N_26579);
xnor U29166 (N_29166,N_26843,N_26618);
or U29167 (N_29167,N_26576,N_27964);
xor U29168 (N_29168,N_27371,N_27563);
and U29169 (N_29169,N_26895,N_26084);
and U29170 (N_29170,N_27606,N_27161);
or U29171 (N_29171,N_26447,N_27742);
nand U29172 (N_29172,N_26283,N_26982);
nand U29173 (N_29173,N_27031,N_27705);
nor U29174 (N_29174,N_27580,N_27796);
nand U29175 (N_29175,N_27316,N_27475);
or U29176 (N_29176,N_26535,N_27239);
nand U29177 (N_29177,N_27917,N_27772);
nor U29178 (N_29178,N_27625,N_26818);
nor U29179 (N_29179,N_26553,N_27084);
or U29180 (N_29180,N_26285,N_26949);
nor U29181 (N_29181,N_27350,N_26556);
nand U29182 (N_29182,N_27662,N_27499);
nor U29183 (N_29183,N_26365,N_26241);
or U29184 (N_29184,N_27736,N_27301);
nor U29185 (N_29185,N_27372,N_27080);
xnor U29186 (N_29186,N_27977,N_27624);
and U29187 (N_29187,N_26361,N_27888);
nand U29188 (N_29188,N_27018,N_26843);
or U29189 (N_29189,N_27506,N_27314);
and U29190 (N_29190,N_27448,N_26924);
xnor U29191 (N_29191,N_26915,N_26027);
xnor U29192 (N_29192,N_27657,N_26694);
nand U29193 (N_29193,N_26190,N_27088);
nand U29194 (N_29194,N_27304,N_26802);
nand U29195 (N_29195,N_26884,N_27167);
xor U29196 (N_29196,N_27795,N_27662);
and U29197 (N_29197,N_27640,N_26609);
or U29198 (N_29198,N_26490,N_26123);
and U29199 (N_29199,N_26537,N_26637);
and U29200 (N_29200,N_26905,N_27617);
and U29201 (N_29201,N_27257,N_27062);
nor U29202 (N_29202,N_27728,N_27304);
nor U29203 (N_29203,N_26054,N_26428);
nor U29204 (N_29204,N_26699,N_26166);
nand U29205 (N_29205,N_26165,N_26179);
or U29206 (N_29206,N_27992,N_27726);
xor U29207 (N_29207,N_26199,N_27014);
or U29208 (N_29208,N_26614,N_26214);
and U29209 (N_29209,N_26300,N_27461);
and U29210 (N_29210,N_27920,N_26205);
nor U29211 (N_29211,N_26266,N_27123);
and U29212 (N_29212,N_27701,N_27957);
nand U29213 (N_29213,N_26284,N_26792);
and U29214 (N_29214,N_26906,N_27202);
nand U29215 (N_29215,N_26606,N_27655);
nand U29216 (N_29216,N_27043,N_26732);
and U29217 (N_29217,N_26453,N_27402);
nor U29218 (N_29218,N_26268,N_27395);
or U29219 (N_29219,N_26281,N_26705);
nand U29220 (N_29220,N_27025,N_27033);
xor U29221 (N_29221,N_26175,N_26228);
and U29222 (N_29222,N_27271,N_26230);
nor U29223 (N_29223,N_26406,N_27361);
and U29224 (N_29224,N_26077,N_27447);
and U29225 (N_29225,N_27528,N_26032);
nor U29226 (N_29226,N_26726,N_26769);
nor U29227 (N_29227,N_27573,N_27336);
and U29228 (N_29228,N_27381,N_26146);
nand U29229 (N_29229,N_27646,N_26599);
nand U29230 (N_29230,N_27050,N_27125);
xor U29231 (N_29231,N_27524,N_26802);
xor U29232 (N_29232,N_27098,N_26578);
xor U29233 (N_29233,N_27078,N_26264);
and U29234 (N_29234,N_26577,N_27016);
or U29235 (N_29235,N_27220,N_26789);
nor U29236 (N_29236,N_27789,N_26104);
and U29237 (N_29237,N_27887,N_27111);
and U29238 (N_29238,N_26890,N_26121);
nor U29239 (N_29239,N_26416,N_27469);
or U29240 (N_29240,N_26427,N_26890);
xnor U29241 (N_29241,N_27383,N_26399);
xnor U29242 (N_29242,N_27809,N_26952);
and U29243 (N_29243,N_26283,N_27872);
or U29244 (N_29244,N_27554,N_27454);
and U29245 (N_29245,N_26335,N_26234);
or U29246 (N_29246,N_26667,N_26488);
or U29247 (N_29247,N_27564,N_27899);
nand U29248 (N_29248,N_27439,N_27773);
nor U29249 (N_29249,N_26207,N_27023);
xor U29250 (N_29250,N_26919,N_27669);
xor U29251 (N_29251,N_26500,N_26299);
nand U29252 (N_29252,N_27239,N_27262);
nor U29253 (N_29253,N_27089,N_27071);
nor U29254 (N_29254,N_26841,N_26298);
xnor U29255 (N_29255,N_26609,N_27336);
xnor U29256 (N_29256,N_27112,N_26390);
nor U29257 (N_29257,N_26418,N_26110);
xor U29258 (N_29258,N_26892,N_26107);
nand U29259 (N_29259,N_26536,N_27390);
and U29260 (N_29260,N_27742,N_26105);
or U29261 (N_29261,N_27329,N_26029);
nand U29262 (N_29262,N_26852,N_26765);
and U29263 (N_29263,N_26277,N_27996);
nand U29264 (N_29264,N_27834,N_26345);
nor U29265 (N_29265,N_27838,N_26124);
nor U29266 (N_29266,N_26404,N_27059);
or U29267 (N_29267,N_27868,N_27280);
nand U29268 (N_29268,N_26566,N_27945);
xor U29269 (N_29269,N_27156,N_27709);
nand U29270 (N_29270,N_26893,N_26795);
nand U29271 (N_29271,N_26003,N_27128);
and U29272 (N_29272,N_26775,N_26170);
xnor U29273 (N_29273,N_26725,N_27985);
nor U29274 (N_29274,N_27323,N_27689);
nor U29275 (N_29275,N_26922,N_26907);
xor U29276 (N_29276,N_27236,N_26784);
nor U29277 (N_29277,N_27252,N_27169);
and U29278 (N_29278,N_26930,N_27041);
and U29279 (N_29279,N_26639,N_27324);
and U29280 (N_29280,N_27266,N_27121);
xor U29281 (N_29281,N_27686,N_27985);
or U29282 (N_29282,N_26605,N_26021);
and U29283 (N_29283,N_27642,N_26567);
nor U29284 (N_29284,N_26667,N_26568);
or U29285 (N_29285,N_27250,N_26160);
and U29286 (N_29286,N_27929,N_26060);
nand U29287 (N_29287,N_27922,N_27790);
and U29288 (N_29288,N_26505,N_26866);
nor U29289 (N_29289,N_27166,N_26456);
and U29290 (N_29290,N_27226,N_27489);
or U29291 (N_29291,N_27721,N_26141);
nand U29292 (N_29292,N_27111,N_27808);
and U29293 (N_29293,N_27388,N_27326);
xor U29294 (N_29294,N_26903,N_27889);
and U29295 (N_29295,N_26993,N_27033);
or U29296 (N_29296,N_27175,N_27806);
xnor U29297 (N_29297,N_26624,N_26670);
or U29298 (N_29298,N_27661,N_26360);
and U29299 (N_29299,N_26691,N_27215);
or U29300 (N_29300,N_26299,N_27148);
or U29301 (N_29301,N_27283,N_27875);
nor U29302 (N_29302,N_27092,N_27412);
and U29303 (N_29303,N_27155,N_26700);
nand U29304 (N_29304,N_27757,N_27147);
nor U29305 (N_29305,N_27325,N_27554);
xnor U29306 (N_29306,N_26197,N_27193);
xnor U29307 (N_29307,N_26441,N_26981);
nor U29308 (N_29308,N_27408,N_27380);
and U29309 (N_29309,N_26220,N_26586);
or U29310 (N_29310,N_27531,N_27176);
xor U29311 (N_29311,N_27452,N_26430);
xor U29312 (N_29312,N_27143,N_26015);
and U29313 (N_29313,N_26261,N_27036);
xnor U29314 (N_29314,N_26242,N_27737);
or U29315 (N_29315,N_27487,N_26831);
nand U29316 (N_29316,N_26309,N_27523);
or U29317 (N_29317,N_27433,N_26424);
xor U29318 (N_29318,N_26081,N_26693);
and U29319 (N_29319,N_26202,N_27414);
xnor U29320 (N_29320,N_26374,N_26976);
nor U29321 (N_29321,N_27158,N_27070);
xor U29322 (N_29322,N_27566,N_26673);
and U29323 (N_29323,N_27392,N_27622);
nand U29324 (N_29324,N_27965,N_26082);
or U29325 (N_29325,N_27326,N_27527);
or U29326 (N_29326,N_26934,N_26766);
and U29327 (N_29327,N_27420,N_27979);
or U29328 (N_29328,N_26120,N_27635);
nand U29329 (N_29329,N_27635,N_26662);
nand U29330 (N_29330,N_27735,N_26794);
xnor U29331 (N_29331,N_27005,N_27555);
and U29332 (N_29332,N_27328,N_26578);
nand U29333 (N_29333,N_27393,N_27236);
xor U29334 (N_29334,N_27357,N_27486);
and U29335 (N_29335,N_27161,N_26250);
xnor U29336 (N_29336,N_27535,N_26743);
nor U29337 (N_29337,N_26547,N_27183);
xor U29338 (N_29338,N_26532,N_26761);
nor U29339 (N_29339,N_27120,N_26915);
nand U29340 (N_29340,N_26089,N_26110);
nor U29341 (N_29341,N_26505,N_26776);
xnor U29342 (N_29342,N_27490,N_27978);
nand U29343 (N_29343,N_26106,N_27653);
xor U29344 (N_29344,N_26937,N_26664);
xnor U29345 (N_29345,N_27063,N_26346);
nor U29346 (N_29346,N_27505,N_26919);
nor U29347 (N_29347,N_27432,N_27086);
nor U29348 (N_29348,N_26669,N_26133);
xor U29349 (N_29349,N_27135,N_26132);
xor U29350 (N_29350,N_27873,N_26170);
or U29351 (N_29351,N_27400,N_27461);
and U29352 (N_29352,N_27171,N_26453);
nor U29353 (N_29353,N_27726,N_26542);
xnor U29354 (N_29354,N_26229,N_27308);
nor U29355 (N_29355,N_26183,N_26416);
xor U29356 (N_29356,N_27417,N_27751);
nor U29357 (N_29357,N_27840,N_27351);
nor U29358 (N_29358,N_26633,N_27607);
nor U29359 (N_29359,N_26853,N_27185);
nor U29360 (N_29360,N_27381,N_27907);
xnor U29361 (N_29361,N_26807,N_26448);
nand U29362 (N_29362,N_27574,N_27754);
nand U29363 (N_29363,N_26710,N_26034);
nor U29364 (N_29364,N_26565,N_27643);
nand U29365 (N_29365,N_27462,N_27456);
xor U29366 (N_29366,N_26470,N_26805);
nor U29367 (N_29367,N_26630,N_26330);
and U29368 (N_29368,N_27553,N_26245);
xnor U29369 (N_29369,N_26344,N_26189);
nor U29370 (N_29370,N_26171,N_27008);
and U29371 (N_29371,N_26391,N_27039);
nor U29372 (N_29372,N_26069,N_27647);
nor U29373 (N_29373,N_27953,N_26971);
or U29374 (N_29374,N_27453,N_27637);
or U29375 (N_29375,N_27785,N_27221);
xnor U29376 (N_29376,N_27157,N_26054);
or U29377 (N_29377,N_27298,N_26041);
and U29378 (N_29378,N_27059,N_27887);
xor U29379 (N_29379,N_26346,N_26369);
xnor U29380 (N_29380,N_26869,N_27616);
xnor U29381 (N_29381,N_26718,N_26633);
and U29382 (N_29382,N_26040,N_27224);
nand U29383 (N_29383,N_26963,N_26824);
and U29384 (N_29384,N_27792,N_26692);
and U29385 (N_29385,N_27631,N_27499);
or U29386 (N_29386,N_26776,N_26895);
nor U29387 (N_29387,N_27859,N_26076);
or U29388 (N_29388,N_26568,N_26594);
xor U29389 (N_29389,N_27476,N_26683);
nor U29390 (N_29390,N_26514,N_27733);
xnor U29391 (N_29391,N_26340,N_27180);
nor U29392 (N_29392,N_27669,N_27132);
or U29393 (N_29393,N_26401,N_26023);
nor U29394 (N_29394,N_27101,N_26822);
nand U29395 (N_29395,N_26546,N_26944);
or U29396 (N_29396,N_26884,N_27429);
xor U29397 (N_29397,N_26465,N_27093);
and U29398 (N_29398,N_27251,N_27533);
nand U29399 (N_29399,N_27561,N_27226);
xnor U29400 (N_29400,N_27967,N_27572);
nor U29401 (N_29401,N_26294,N_26556);
xor U29402 (N_29402,N_26616,N_26536);
and U29403 (N_29403,N_26953,N_27653);
nor U29404 (N_29404,N_27833,N_26252);
nand U29405 (N_29405,N_27051,N_26203);
or U29406 (N_29406,N_27149,N_26775);
nand U29407 (N_29407,N_27169,N_27915);
nor U29408 (N_29408,N_26649,N_27331);
and U29409 (N_29409,N_27377,N_27619);
nand U29410 (N_29410,N_27962,N_27326);
nand U29411 (N_29411,N_26256,N_27195);
xor U29412 (N_29412,N_27799,N_26738);
and U29413 (N_29413,N_27585,N_26803);
nand U29414 (N_29414,N_27652,N_27569);
or U29415 (N_29415,N_27009,N_26678);
nor U29416 (N_29416,N_26608,N_27187);
nor U29417 (N_29417,N_26695,N_26779);
nand U29418 (N_29418,N_26630,N_27456);
xnor U29419 (N_29419,N_26290,N_26885);
xnor U29420 (N_29420,N_27248,N_27807);
nor U29421 (N_29421,N_27799,N_26469);
nor U29422 (N_29422,N_27558,N_27132);
xor U29423 (N_29423,N_26348,N_26251);
or U29424 (N_29424,N_27922,N_27304);
or U29425 (N_29425,N_26311,N_27172);
or U29426 (N_29426,N_27611,N_27672);
or U29427 (N_29427,N_27708,N_27339);
nand U29428 (N_29428,N_27921,N_26949);
xor U29429 (N_29429,N_26715,N_27432);
nor U29430 (N_29430,N_26481,N_26436);
or U29431 (N_29431,N_26908,N_26200);
nand U29432 (N_29432,N_27804,N_27341);
and U29433 (N_29433,N_27877,N_27235);
nor U29434 (N_29434,N_27567,N_26466);
or U29435 (N_29435,N_26996,N_26388);
or U29436 (N_29436,N_26270,N_27206);
and U29437 (N_29437,N_26894,N_26889);
xor U29438 (N_29438,N_27277,N_26342);
nand U29439 (N_29439,N_26529,N_26084);
or U29440 (N_29440,N_27065,N_27208);
or U29441 (N_29441,N_27140,N_26397);
and U29442 (N_29442,N_27981,N_26158);
and U29443 (N_29443,N_26087,N_27713);
and U29444 (N_29444,N_26461,N_27111);
or U29445 (N_29445,N_27910,N_27926);
nand U29446 (N_29446,N_27458,N_26553);
nor U29447 (N_29447,N_26320,N_26378);
nand U29448 (N_29448,N_26848,N_26259);
nor U29449 (N_29449,N_26096,N_27855);
nor U29450 (N_29450,N_27335,N_27795);
xor U29451 (N_29451,N_27727,N_27531);
or U29452 (N_29452,N_27627,N_26135);
nor U29453 (N_29453,N_26332,N_27791);
xnor U29454 (N_29454,N_27190,N_26742);
and U29455 (N_29455,N_26061,N_27998);
nand U29456 (N_29456,N_26114,N_26031);
and U29457 (N_29457,N_27147,N_27388);
xor U29458 (N_29458,N_27212,N_26144);
nor U29459 (N_29459,N_26386,N_26794);
xor U29460 (N_29460,N_26548,N_27154);
xor U29461 (N_29461,N_26395,N_26961);
xor U29462 (N_29462,N_27900,N_26303);
nor U29463 (N_29463,N_26928,N_27244);
and U29464 (N_29464,N_26427,N_26632);
or U29465 (N_29465,N_27776,N_27398);
xor U29466 (N_29466,N_27819,N_27159);
and U29467 (N_29467,N_26566,N_26567);
xor U29468 (N_29468,N_26609,N_26614);
xor U29469 (N_29469,N_26947,N_26501);
and U29470 (N_29470,N_26430,N_26358);
and U29471 (N_29471,N_27119,N_27286);
and U29472 (N_29472,N_26976,N_27643);
nand U29473 (N_29473,N_26021,N_27476);
or U29474 (N_29474,N_27546,N_26347);
xnor U29475 (N_29475,N_26144,N_27501);
xnor U29476 (N_29476,N_26878,N_27350);
or U29477 (N_29477,N_27149,N_27399);
nand U29478 (N_29478,N_26868,N_27766);
xnor U29479 (N_29479,N_26300,N_26293);
and U29480 (N_29480,N_26005,N_26023);
nor U29481 (N_29481,N_26768,N_26285);
or U29482 (N_29482,N_26862,N_27606);
and U29483 (N_29483,N_26922,N_26940);
and U29484 (N_29484,N_27103,N_26283);
xor U29485 (N_29485,N_27576,N_27138);
or U29486 (N_29486,N_26883,N_27577);
nor U29487 (N_29487,N_26471,N_26122);
nor U29488 (N_29488,N_26413,N_26571);
nor U29489 (N_29489,N_26674,N_26993);
xor U29490 (N_29490,N_26695,N_26748);
xnor U29491 (N_29491,N_26729,N_26801);
nor U29492 (N_29492,N_27572,N_27276);
xor U29493 (N_29493,N_27564,N_26909);
nor U29494 (N_29494,N_27627,N_26727);
and U29495 (N_29495,N_26507,N_27653);
or U29496 (N_29496,N_26495,N_26436);
and U29497 (N_29497,N_26257,N_26511);
nor U29498 (N_29498,N_26287,N_26137);
nand U29499 (N_29499,N_27546,N_27595);
nor U29500 (N_29500,N_27192,N_27930);
and U29501 (N_29501,N_27871,N_26277);
and U29502 (N_29502,N_27949,N_26925);
nor U29503 (N_29503,N_27920,N_26490);
nor U29504 (N_29504,N_27223,N_27729);
nor U29505 (N_29505,N_26118,N_26817);
or U29506 (N_29506,N_26404,N_26702);
xnor U29507 (N_29507,N_26684,N_26995);
xnor U29508 (N_29508,N_27119,N_26507);
or U29509 (N_29509,N_26281,N_27890);
nand U29510 (N_29510,N_27971,N_27141);
xor U29511 (N_29511,N_27524,N_26729);
and U29512 (N_29512,N_26851,N_26586);
xor U29513 (N_29513,N_27587,N_27574);
and U29514 (N_29514,N_27154,N_26392);
nand U29515 (N_29515,N_26339,N_26556);
nor U29516 (N_29516,N_27630,N_26479);
or U29517 (N_29517,N_26752,N_27010);
and U29518 (N_29518,N_27034,N_26382);
nand U29519 (N_29519,N_26968,N_27190);
and U29520 (N_29520,N_26828,N_27201);
nor U29521 (N_29521,N_26322,N_27795);
nor U29522 (N_29522,N_27849,N_27331);
nand U29523 (N_29523,N_27910,N_26113);
nor U29524 (N_29524,N_27138,N_26440);
or U29525 (N_29525,N_26796,N_27790);
xnor U29526 (N_29526,N_27198,N_26413);
and U29527 (N_29527,N_26814,N_26869);
or U29528 (N_29528,N_27066,N_26584);
nor U29529 (N_29529,N_26529,N_26251);
or U29530 (N_29530,N_27948,N_26221);
nor U29531 (N_29531,N_26914,N_26685);
nor U29532 (N_29532,N_26121,N_26772);
nand U29533 (N_29533,N_27091,N_26182);
and U29534 (N_29534,N_27516,N_26670);
or U29535 (N_29535,N_26874,N_26465);
and U29536 (N_29536,N_27888,N_26205);
xnor U29537 (N_29537,N_26575,N_27102);
or U29538 (N_29538,N_27143,N_26129);
and U29539 (N_29539,N_27324,N_26941);
and U29540 (N_29540,N_27014,N_26184);
xnor U29541 (N_29541,N_26480,N_27119);
and U29542 (N_29542,N_27310,N_27380);
nor U29543 (N_29543,N_26469,N_26451);
nor U29544 (N_29544,N_27895,N_27049);
and U29545 (N_29545,N_26383,N_27460);
nor U29546 (N_29546,N_26478,N_27538);
and U29547 (N_29547,N_26285,N_27950);
or U29548 (N_29548,N_27088,N_27295);
nand U29549 (N_29549,N_27324,N_27881);
nor U29550 (N_29550,N_27272,N_27022);
xnor U29551 (N_29551,N_26334,N_27393);
nand U29552 (N_29552,N_26384,N_27258);
and U29553 (N_29553,N_26323,N_27795);
nand U29554 (N_29554,N_27170,N_26182);
and U29555 (N_29555,N_26245,N_26514);
or U29556 (N_29556,N_26745,N_26920);
nor U29557 (N_29557,N_27484,N_27546);
and U29558 (N_29558,N_26869,N_27809);
nor U29559 (N_29559,N_27923,N_27043);
xor U29560 (N_29560,N_27250,N_26339);
and U29561 (N_29561,N_26682,N_27323);
or U29562 (N_29562,N_26201,N_26747);
nand U29563 (N_29563,N_26534,N_27881);
or U29564 (N_29564,N_27784,N_26502);
and U29565 (N_29565,N_26671,N_26531);
xor U29566 (N_29566,N_27374,N_26117);
nand U29567 (N_29567,N_27309,N_26819);
and U29568 (N_29568,N_27432,N_27316);
xnor U29569 (N_29569,N_26578,N_27491);
nor U29570 (N_29570,N_27435,N_26527);
and U29571 (N_29571,N_26223,N_26980);
or U29572 (N_29572,N_27604,N_27012);
nor U29573 (N_29573,N_26402,N_27718);
and U29574 (N_29574,N_27084,N_27132);
or U29575 (N_29575,N_27663,N_27916);
and U29576 (N_29576,N_26365,N_27320);
nor U29577 (N_29577,N_26579,N_26277);
and U29578 (N_29578,N_27441,N_27209);
nor U29579 (N_29579,N_27158,N_27234);
nor U29580 (N_29580,N_26747,N_27184);
or U29581 (N_29581,N_27729,N_27857);
xor U29582 (N_29582,N_27856,N_27469);
and U29583 (N_29583,N_27965,N_27986);
xnor U29584 (N_29584,N_26180,N_27645);
or U29585 (N_29585,N_26264,N_27044);
or U29586 (N_29586,N_26362,N_26174);
or U29587 (N_29587,N_26772,N_26681);
xor U29588 (N_29588,N_27385,N_27974);
nand U29589 (N_29589,N_26700,N_27255);
or U29590 (N_29590,N_26844,N_27594);
xnor U29591 (N_29591,N_27047,N_26132);
nor U29592 (N_29592,N_26585,N_27699);
nand U29593 (N_29593,N_26515,N_26413);
xor U29594 (N_29594,N_26626,N_26566);
nand U29595 (N_29595,N_27351,N_27259);
xnor U29596 (N_29596,N_26654,N_26051);
and U29597 (N_29597,N_26338,N_26116);
or U29598 (N_29598,N_26238,N_26020);
nand U29599 (N_29599,N_27987,N_27134);
or U29600 (N_29600,N_26276,N_27090);
xor U29601 (N_29601,N_27999,N_26055);
or U29602 (N_29602,N_27003,N_27115);
and U29603 (N_29603,N_27940,N_26822);
or U29604 (N_29604,N_27856,N_27490);
xnor U29605 (N_29605,N_26854,N_26054);
or U29606 (N_29606,N_27931,N_27230);
xor U29607 (N_29607,N_26173,N_27012);
and U29608 (N_29608,N_27271,N_26836);
and U29609 (N_29609,N_27677,N_26340);
nand U29610 (N_29610,N_26977,N_27636);
nor U29611 (N_29611,N_26119,N_27433);
and U29612 (N_29612,N_26020,N_27305);
nor U29613 (N_29613,N_26588,N_27613);
xor U29614 (N_29614,N_26049,N_26566);
nor U29615 (N_29615,N_26623,N_26130);
or U29616 (N_29616,N_26301,N_27732);
xnor U29617 (N_29617,N_26382,N_27634);
and U29618 (N_29618,N_26477,N_27198);
or U29619 (N_29619,N_26340,N_27678);
nand U29620 (N_29620,N_27910,N_26477);
nor U29621 (N_29621,N_27027,N_27440);
or U29622 (N_29622,N_26769,N_27872);
or U29623 (N_29623,N_26761,N_27240);
or U29624 (N_29624,N_26484,N_26751);
nor U29625 (N_29625,N_27121,N_26505);
or U29626 (N_29626,N_27452,N_26534);
nand U29627 (N_29627,N_27096,N_26632);
xor U29628 (N_29628,N_26098,N_27402);
nor U29629 (N_29629,N_27943,N_27632);
nor U29630 (N_29630,N_26714,N_27001);
xor U29631 (N_29631,N_27327,N_27361);
nor U29632 (N_29632,N_26273,N_27988);
or U29633 (N_29633,N_26290,N_26617);
nand U29634 (N_29634,N_26476,N_26791);
xnor U29635 (N_29635,N_27041,N_27152);
nand U29636 (N_29636,N_26271,N_26037);
and U29637 (N_29637,N_26782,N_26312);
xnor U29638 (N_29638,N_26536,N_27305);
and U29639 (N_29639,N_26144,N_27012);
nand U29640 (N_29640,N_27843,N_26349);
nand U29641 (N_29641,N_26660,N_26253);
and U29642 (N_29642,N_26358,N_26884);
and U29643 (N_29643,N_26408,N_27406);
nor U29644 (N_29644,N_26779,N_27461);
nor U29645 (N_29645,N_26358,N_27020);
and U29646 (N_29646,N_26957,N_26868);
or U29647 (N_29647,N_27581,N_26220);
xor U29648 (N_29648,N_26721,N_27466);
or U29649 (N_29649,N_26143,N_26633);
nor U29650 (N_29650,N_27835,N_26928);
or U29651 (N_29651,N_26934,N_26708);
or U29652 (N_29652,N_26204,N_27674);
and U29653 (N_29653,N_27748,N_27510);
nand U29654 (N_29654,N_26727,N_26013);
nand U29655 (N_29655,N_26248,N_26857);
and U29656 (N_29656,N_27820,N_27664);
or U29657 (N_29657,N_27905,N_27300);
or U29658 (N_29658,N_26749,N_27713);
or U29659 (N_29659,N_27185,N_26047);
nand U29660 (N_29660,N_27261,N_27342);
or U29661 (N_29661,N_27496,N_26220);
nor U29662 (N_29662,N_27188,N_26436);
nor U29663 (N_29663,N_26240,N_27119);
nor U29664 (N_29664,N_26071,N_26925);
or U29665 (N_29665,N_26639,N_26646);
xnor U29666 (N_29666,N_26299,N_26375);
nor U29667 (N_29667,N_26520,N_27988);
xor U29668 (N_29668,N_27226,N_26253);
xnor U29669 (N_29669,N_26643,N_27489);
and U29670 (N_29670,N_27885,N_27928);
and U29671 (N_29671,N_26056,N_27879);
or U29672 (N_29672,N_27361,N_27056);
xor U29673 (N_29673,N_26074,N_27928);
nand U29674 (N_29674,N_26077,N_27904);
xnor U29675 (N_29675,N_27295,N_27656);
nor U29676 (N_29676,N_27975,N_26961);
nand U29677 (N_29677,N_27118,N_27831);
nand U29678 (N_29678,N_27029,N_27328);
or U29679 (N_29679,N_26054,N_26285);
and U29680 (N_29680,N_27422,N_27769);
and U29681 (N_29681,N_27784,N_27239);
nor U29682 (N_29682,N_27370,N_27858);
nand U29683 (N_29683,N_26681,N_27370);
and U29684 (N_29684,N_27370,N_27032);
or U29685 (N_29685,N_27450,N_27735);
nand U29686 (N_29686,N_27459,N_26749);
nor U29687 (N_29687,N_27857,N_27347);
nor U29688 (N_29688,N_27202,N_26013);
and U29689 (N_29689,N_26293,N_27094);
nor U29690 (N_29690,N_27980,N_27876);
nor U29691 (N_29691,N_27418,N_26989);
nor U29692 (N_29692,N_27263,N_26062);
xor U29693 (N_29693,N_26402,N_26647);
nand U29694 (N_29694,N_27035,N_27018);
nand U29695 (N_29695,N_27510,N_27652);
nor U29696 (N_29696,N_26474,N_26016);
or U29697 (N_29697,N_27464,N_26686);
or U29698 (N_29698,N_26638,N_26616);
or U29699 (N_29699,N_27356,N_27755);
nand U29700 (N_29700,N_26370,N_26245);
xnor U29701 (N_29701,N_27324,N_27438);
xor U29702 (N_29702,N_27611,N_26533);
nand U29703 (N_29703,N_26661,N_27926);
and U29704 (N_29704,N_26160,N_26317);
or U29705 (N_29705,N_26528,N_27693);
or U29706 (N_29706,N_26965,N_27539);
xor U29707 (N_29707,N_27388,N_27532);
and U29708 (N_29708,N_27945,N_26573);
xnor U29709 (N_29709,N_27592,N_26453);
nor U29710 (N_29710,N_27868,N_26833);
nor U29711 (N_29711,N_26760,N_26300);
or U29712 (N_29712,N_27070,N_27121);
and U29713 (N_29713,N_27725,N_27822);
nor U29714 (N_29714,N_26902,N_26345);
nand U29715 (N_29715,N_27732,N_27251);
or U29716 (N_29716,N_27405,N_27424);
or U29717 (N_29717,N_27072,N_26055);
nor U29718 (N_29718,N_26133,N_26936);
and U29719 (N_29719,N_26334,N_27586);
or U29720 (N_29720,N_26880,N_27247);
or U29721 (N_29721,N_26508,N_26891);
and U29722 (N_29722,N_27290,N_27220);
and U29723 (N_29723,N_26431,N_27231);
nor U29724 (N_29724,N_27614,N_26923);
nor U29725 (N_29725,N_27196,N_26300);
nor U29726 (N_29726,N_27580,N_27971);
xnor U29727 (N_29727,N_27218,N_26303);
and U29728 (N_29728,N_26826,N_27996);
and U29729 (N_29729,N_27704,N_27572);
nand U29730 (N_29730,N_26284,N_26844);
and U29731 (N_29731,N_26605,N_27685);
xor U29732 (N_29732,N_26057,N_27398);
nor U29733 (N_29733,N_27780,N_27353);
or U29734 (N_29734,N_26864,N_26705);
nor U29735 (N_29735,N_26271,N_26278);
xor U29736 (N_29736,N_26452,N_26598);
and U29737 (N_29737,N_27887,N_27207);
nor U29738 (N_29738,N_26797,N_26751);
and U29739 (N_29739,N_27139,N_27282);
or U29740 (N_29740,N_26103,N_27871);
and U29741 (N_29741,N_26169,N_26286);
nand U29742 (N_29742,N_27916,N_27022);
nor U29743 (N_29743,N_27149,N_26504);
nand U29744 (N_29744,N_27166,N_26436);
nand U29745 (N_29745,N_26837,N_26770);
nor U29746 (N_29746,N_27932,N_26380);
nand U29747 (N_29747,N_26718,N_26410);
or U29748 (N_29748,N_27129,N_27415);
nor U29749 (N_29749,N_26896,N_26425);
nor U29750 (N_29750,N_27891,N_26256);
nor U29751 (N_29751,N_27309,N_27136);
or U29752 (N_29752,N_27550,N_26473);
xnor U29753 (N_29753,N_26491,N_26775);
xnor U29754 (N_29754,N_27191,N_26519);
and U29755 (N_29755,N_27452,N_26427);
nor U29756 (N_29756,N_27698,N_26299);
xnor U29757 (N_29757,N_27568,N_27669);
nand U29758 (N_29758,N_26147,N_26922);
nor U29759 (N_29759,N_26257,N_26742);
nor U29760 (N_29760,N_27430,N_27911);
nand U29761 (N_29761,N_26974,N_26426);
nand U29762 (N_29762,N_26885,N_26393);
or U29763 (N_29763,N_26571,N_26349);
and U29764 (N_29764,N_27533,N_27588);
nand U29765 (N_29765,N_27470,N_26175);
and U29766 (N_29766,N_26275,N_26337);
or U29767 (N_29767,N_27580,N_27724);
or U29768 (N_29768,N_27566,N_27913);
nand U29769 (N_29769,N_26370,N_26633);
nand U29770 (N_29770,N_26522,N_27658);
xnor U29771 (N_29771,N_26693,N_27634);
and U29772 (N_29772,N_26357,N_26283);
and U29773 (N_29773,N_26986,N_27153);
and U29774 (N_29774,N_27022,N_26347);
or U29775 (N_29775,N_26973,N_26542);
or U29776 (N_29776,N_27089,N_27288);
nand U29777 (N_29777,N_27611,N_26270);
or U29778 (N_29778,N_27886,N_27258);
nor U29779 (N_29779,N_26225,N_26895);
and U29780 (N_29780,N_26542,N_27334);
nor U29781 (N_29781,N_26599,N_27743);
nor U29782 (N_29782,N_27578,N_26752);
and U29783 (N_29783,N_27899,N_26311);
nand U29784 (N_29784,N_27323,N_27164);
nand U29785 (N_29785,N_27018,N_26905);
nor U29786 (N_29786,N_26744,N_27199);
nor U29787 (N_29787,N_26026,N_26663);
xnor U29788 (N_29788,N_27265,N_26417);
nand U29789 (N_29789,N_26314,N_26011);
nand U29790 (N_29790,N_26541,N_27388);
xor U29791 (N_29791,N_26032,N_27597);
nor U29792 (N_29792,N_27194,N_26564);
and U29793 (N_29793,N_27585,N_26472);
xor U29794 (N_29794,N_26706,N_26621);
xor U29795 (N_29795,N_26550,N_27972);
nor U29796 (N_29796,N_27658,N_27767);
nand U29797 (N_29797,N_26885,N_27818);
and U29798 (N_29798,N_27945,N_27888);
xnor U29799 (N_29799,N_26178,N_26047);
nor U29800 (N_29800,N_27161,N_27535);
xor U29801 (N_29801,N_26247,N_27626);
xor U29802 (N_29802,N_26419,N_26541);
or U29803 (N_29803,N_27885,N_27404);
nor U29804 (N_29804,N_26998,N_27342);
nand U29805 (N_29805,N_26576,N_26896);
and U29806 (N_29806,N_26454,N_26221);
nand U29807 (N_29807,N_27125,N_26914);
and U29808 (N_29808,N_26774,N_26405);
xnor U29809 (N_29809,N_26550,N_27962);
xnor U29810 (N_29810,N_26971,N_26432);
nand U29811 (N_29811,N_27263,N_26554);
or U29812 (N_29812,N_26830,N_26331);
or U29813 (N_29813,N_27495,N_26964);
nand U29814 (N_29814,N_27112,N_27159);
nand U29815 (N_29815,N_27837,N_26886);
and U29816 (N_29816,N_26766,N_26923);
nand U29817 (N_29817,N_26450,N_27307);
or U29818 (N_29818,N_27170,N_26009);
and U29819 (N_29819,N_26736,N_27810);
nand U29820 (N_29820,N_27695,N_26700);
nand U29821 (N_29821,N_27101,N_27512);
nand U29822 (N_29822,N_27624,N_26421);
and U29823 (N_29823,N_26684,N_27630);
and U29824 (N_29824,N_27656,N_27414);
or U29825 (N_29825,N_26919,N_27640);
nand U29826 (N_29826,N_27816,N_27892);
or U29827 (N_29827,N_27958,N_27771);
nand U29828 (N_29828,N_27693,N_26610);
xnor U29829 (N_29829,N_27806,N_27479);
nor U29830 (N_29830,N_27980,N_26580);
xor U29831 (N_29831,N_26138,N_26654);
xnor U29832 (N_29832,N_27617,N_26901);
and U29833 (N_29833,N_27088,N_26982);
xnor U29834 (N_29834,N_26842,N_27382);
nand U29835 (N_29835,N_26832,N_26239);
nand U29836 (N_29836,N_26996,N_26931);
nor U29837 (N_29837,N_27802,N_27348);
nand U29838 (N_29838,N_27202,N_27847);
and U29839 (N_29839,N_27996,N_26650);
or U29840 (N_29840,N_26563,N_27729);
xnor U29841 (N_29841,N_27779,N_27452);
or U29842 (N_29842,N_27785,N_27076);
nor U29843 (N_29843,N_26685,N_27454);
xor U29844 (N_29844,N_27378,N_27551);
or U29845 (N_29845,N_27594,N_26059);
xnor U29846 (N_29846,N_27852,N_27519);
nand U29847 (N_29847,N_27605,N_26193);
nor U29848 (N_29848,N_27343,N_27404);
and U29849 (N_29849,N_27970,N_27003);
xor U29850 (N_29850,N_26200,N_26964);
or U29851 (N_29851,N_27508,N_27475);
nand U29852 (N_29852,N_27915,N_26016);
xor U29853 (N_29853,N_26063,N_26591);
nand U29854 (N_29854,N_26547,N_26029);
xnor U29855 (N_29855,N_27790,N_27874);
xnor U29856 (N_29856,N_26083,N_27059);
xnor U29857 (N_29857,N_27499,N_26019);
or U29858 (N_29858,N_27424,N_26860);
nor U29859 (N_29859,N_27674,N_26879);
and U29860 (N_29860,N_27489,N_27374);
nor U29861 (N_29861,N_26032,N_27440);
nor U29862 (N_29862,N_27130,N_26818);
and U29863 (N_29863,N_27019,N_26764);
xor U29864 (N_29864,N_26585,N_27960);
and U29865 (N_29865,N_26480,N_27550);
nor U29866 (N_29866,N_27971,N_26757);
nand U29867 (N_29867,N_27974,N_27279);
or U29868 (N_29868,N_27707,N_27914);
xnor U29869 (N_29869,N_27017,N_26531);
or U29870 (N_29870,N_26827,N_27159);
or U29871 (N_29871,N_27568,N_26688);
and U29872 (N_29872,N_26943,N_27816);
and U29873 (N_29873,N_26095,N_26793);
nand U29874 (N_29874,N_26133,N_26646);
and U29875 (N_29875,N_26701,N_26137);
and U29876 (N_29876,N_27925,N_26593);
xnor U29877 (N_29877,N_26977,N_27730);
or U29878 (N_29878,N_26894,N_26276);
or U29879 (N_29879,N_26870,N_27075);
or U29880 (N_29880,N_26943,N_26416);
nand U29881 (N_29881,N_26830,N_27620);
and U29882 (N_29882,N_26800,N_27875);
or U29883 (N_29883,N_26455,N_27394);
nor U29884 (N_29884,N_26178,N_27300);
or U29885 (N_29885,N_27670,N_27424);
nand U29886 (N_29886,N_27628,N_27945);
and U29887 (N_29887,N_27936,N_27381);
nor U29888 (N_29888,N_26900,N_27927);
and U29889 (N_29889,N_27156,N_26838);
nor U29890 (N_29890,N_27654,N_27208);
or U29891 (N_29891,N_27893,N_27018);
nor U29892 (N_29892,N_27633,N_26514);
xor U29893 (N_29893,N_26915,N_27659);
xnor U29894 (N_29894,N_26093,N_26592);
nand U29895 (N_29895,N_27365,N_26989);
or U29896 (N_29896,N_27705,N_27352);
nand U29897 (N_29897,N_27831,N_27888);
xor U29898 (N_29898,N_27188,N_27659);
and U29899 (N_29899,N_27929,N_27674);
or U29900 (N_29900,N_26156,N_26275);
and U29901 (N_29901,N_26077,N_26716);
nor U29902 (N_29902,N_26445,N_27319);
and U29903 (N_29903,N_27290,N_27034);
xor U29904 (N_29904,N_26718,N_27559);
xor U29905 (N_29905,N_27427,N_26611);
nor U29906 (N_29906,N_26575,N_26425);
nor U29907 (N_29907,N_26091,N_26925);
or U29908 (N_29908,N_26700,N_26911);
and U29909 (N_29909,N_26490,N_26177);
and U29910 (N_29910,N_26937,N_26800);
nor U29911 (N_29911,N_26089,N_27724);
and U29912 (N_29912,N_26960,N_27166);
or U29913 (N_29913,N_27656,N_26087);
nor U29914 (N_29914,N_27772,N_27310);
nand U29915 (N_29915,N_26492,N_26870);
xnor U29916 (N_29916,N_26462,N_27162);
nand U29917 (N_29917,N_27538,N_26057);
or U29918 (N_29918,N_26959,N_27556);
and U29919 (N_29919,N_27599,N_27652);
nand U29920 (N_29920,N_27929,N_26252);
nor U29921 (N_29921,N_26275,N_27305);
xnor U29922 (N_29922,N_27438,N_26850);
xnor U29923 (N_29923,N_27793,N_27304);
xor U29924 (N_29924,N_27667,N_27298);
and U29925 (N_29925,N_27626,N_26571);
nor U29926 (N_29926,N_26912,N_27510);
nand U29927 (N_29927,N_27020,N_27325);
and U29928 (N_29928,N_27034,N_26589);
nand U29929 (N_29929,N_27511,N_26237);
nand U29930 (N_29930,N_26652,N_26942);
nand U29931 (N_29931,N_26131,N_26388);
and U29932 (N_29932,N_26700,N_26439);
xnor U29933 (N_29933,N_27269,N_27618);
and U29934 (N_29934,N_26976,N_27947);
and U29935 (N_29935,N_27090,N_26451);
or U29936 (N_29936,N_27429,N_26605);
nor U29937 (N_29937,N_27940,N_26983);
nand U29938 (N_29938,N_27819,N_26610);
nor U29939 (N_29939,N_27704,N_26700);
or U29940 (N_29940,N_27513,N_26926);
xor U29941 (N_29941,N_27294,N_26451);
nand U29942 (N_29942,N_27389,N_26933);
nor U29943 (N_29943,N_26733,N_27536);
nand U29944 (N_29944,N_26257,N_26639);
xor U29945 (N_29945,N_27325,N_26579);
and U29946 (N_29946,N_26109,N_26664);
or U29947 (N_29947,N_26117,N_27791);
nand U29948 (N_29948,N_27266,N_26657);
nor U29949 (N_29949,N_27560,N_27394);
xnor U29950 (N_29950,N_27657,N_26822);
nand U29951 (N_29951,N_27294,N_27575);
or U29952 (N_29952,N_26825,N_27988);
or U29953 (N_29953,N_27623,N_26502);
and U29954 (N_29954,N_26655,N_27019);
or U29955 (N_29955,N_26359,N_26857);
nand U29956 (N_29956,N_27753,N_27860);
nor U29957 (N_29957,N_27150,N_26120);
and U29958 (N_29958,N_26625,N_26974);
and U29959 (N_29959,N_26200,N_27979);
nand U29960 (N_29960,N_26492,N_27591);
nand U29961 (N_29961,N_27896,N_26647);
nor U29962 (N_29962,N_27627,N_27940);
xnor U29963 (N_29963,N_27359,N_26341);
nor U29964 (N_29964,N_27466,N_27662);
and U29965 (N_29965,N_26865,N_26619);
or U29966 (N_29966,N_26869,N_26821);
nor U29967 (N_29967,N_27093,N_26697);
nand U29968 (N_29968,N_27949,N_26819);
nand U29969 (N_29969,N_26397,N_27695);
nor U29970 (N_29970,N_27344,N_26118);
or U29971 (N_29971,N_27230,N_27553);
or U29972 (N_29972,N_27603,N_27349);
or U29973 (N_29973,N_26797,N_26581);
xnor U29974 (N_29974,N_27427,N_27198);
xnor U29975 (N_29975,N_27282,N_26707);
and U29976 (N_29976,N_26264,N_27691);
xnor U29977 (N_29977,N_26423,N_27425);
xor U29978 (N_29978,N_26236,N_26215);
xor U29979 (N_29979,N_26546,N_26437);
or U29980 (N_29980,N_26775,N_26434);
or U29981 (N_29981,N_26685,N_26597);
nor U29982 (N_29982,N_27833,N_26231);
nand U29983 (N_29983,N_26035,N_27463);
nand U29984 (N_29984,N_27147,N_26151);
xnor U29985 (N_29985,N_26512,N_26138);
nor U29986 (N_29986,N_27399,N_27924);
xor U29987 (N_29987,N_26299,N_26031);
or U29988 (N_29988,N_27785,N_26626);
nand U29989 (N_29989,N_27756,N_27441);
nor U29990 (N_29990,N_26014,N_26385);
and U29991 (N_29991,N_27389,N_27984);
or U29992 (N_29992,N_26713,N_27451);
nand U29993 (N_29993,N_26028,N_26937);
and U29994 (N_29994,N_27849,N_26314);
nor U29995 (N_29995,N_27239,N_27406);
nor U29996 (N_29996,N_26272,N_26788);
nand U29997 (N_29997,N_26766,N_26860);
nand U29998 (N_29998,N_26440,N_26577);
or U29999 (N_29999,N_27327,N_26733);
and U30000 (N_30000,N_28551,N_28837);
nand U30001 (N_30001,N_29210,N_29357);
nand U30002 (N_30002,N_29911,N_28416);
xor U30003 (N_30003,N_28607,N_29092);
nor U30004 (N_30004,N_29400,N_28300);
and U30005 (N_30005,N_29855,N_28650);
or U30006 (N_30006,N_29966,N_28344);
nor U30007 (N_30007,N_28747,N_29053);
nand U30008 (N_30008,N_29059,N_29449);
nor U30009 (N_30009,N_28663,N_28867);
and U30010 (N_30010,N_29422,N_29285);
nand U30011 (N_30011,N_28406,N_28053);
xnor U30012 (N_30012,N_28444,N_29964);
xnor U30013 (N_30013,N_28609,N_29645);
or U30014 (N_30014,N_28021,N_29200);
or U30015 (N_30015,N_29773,N_29659);
and U30016 (N_30016,N_28785,N_29873);
and U30017 (N_30017,N_28065,N_28642);
and U30018 (N_30018,N_28799,N_28546);
xnor U30019 (N_30019,N_29105,N_29170);
and U30020 (N_30020,N_29867,N_29483);
or U30021 (N_30021,N_28713,N_28373);
and U30022 (N_30022,N_28701,N_29507);
or U30023 (N_30023,N_28782,N_29700);
xor U30024 (N_30024,N_28221,N_28153);
nand U30025 (N_30025,N_28910,N_28843);
xnor U30026 (N_30026,N_28521,N_28679);
xnor U30027 (N_30027,N_29187,N_29020);
and U30028 (N_30028,N_28139,N_28795);
nor U30029 (N_30029,N_28717,N_29231);
and U30030 (N_30030,N_28338,N_28948);
or U30031 (N_30031,N_29906,N_29260);
xnor U30032 (N_30032,N_29727,N_28417);
nor U30033 (N_30033,N_29537,N_29661);
nor U30034 (N_30034,N_29251,N_28596);
nand U30035 (N_30035,N_29012,N_29632);
nor U30036 (N_30036,N_29191,N_28236);
and U30037 (N_30037,N_29024,N_28572);
nor U30038 (N_30038,N_29453,N_29533);
or U30039 (N_30039,N_28113,N_28363);
nor U30040 (N_30040,N_29874,N_29624);
nor U30041 (N_30041,N_28073,N_29636);
or U30042 (N_30042,N_29499,N_29578);
nand U30043 (N_30043,N_29701,N_29687);
nand U30044 (N_30044,N_29702,N_28577);
xnor U30045 (N_30045,N_29017,N_29154);
nor U30046 (N_30046,N_29775,N_29954);
or U30047 (N_30047,N_28265,N_28762);
nand U30048 (N_30048,N_28168,N_28295);
or U30049 (N_30049,N_28039,N_29279);
nand U30050 (N_30050,N_28158,N_29468);
nand U30051 (N_30051,N_29013,N_29914);
nand U30052 (N_30052,N_29295,N_29014);
and U30053 (N_30053,N_29192,N_29642);
nand U30054 (N_30054,N_29056,N_28240);
xnor U30055 (N_30055,N_29863,N_28237);
nand U30056 (N_30056,N_28958,N_28990);
xor U30057 (N_30057,N_28057,N_29389);
xor U30058 (N_30058,N_28340,N_28419);
nand U30059 (N_30059,N_28014,N_29073);
and U30060 (N_30060,N_29511,N_29590);
xnor U30061 (N_30061,N_29842,N_29823);
nor U30062 (N_30062,N_28219,N_28704);
nand U30063 (N_30063,N_28125,N_28686);
nand U30064 (N_30064,N_28031,N_28768);
or U30065 (N_30065,N_29447,N_29932);
nor U30066 (N_30066,N_29293,N_29054);
xor U30067 (N_30067,N_28227,N_28766);
or U30068 (N_30068,N_28235,N_28844);
nor U30069 (N_30069,N_28116,N_28915);
xor U30070 (N_30070,N_29488,N_29045);
and U30071 (N_30071,N_29060,N_29321);
xor U30072 (N_30072,N_28145,N_29201);
xor U30073 (N_30073,N_29395,N_29322);
and U30074 (N_30074,N_29387,N_28839);
xnor U30075 (N_30075,N_29319,N_29692);
and U30076 (N_30076,N_28093,N_28180);
xnor U30077 (N_30077,N_29156,N_29588);
or U30078 (N_30078,N_28019,N_29253);
nand U30079 (N_30079,N_29610,N_28926);
xnor U30080 (N_30080,N_28507,N_28941);
nand U30081 (N_30081,N_28722,N_29265);
xnor U30082 (N_30082,N_29124,N_29397);
and U30083 (N_30083,N_28710,N_28280);
and U30084 (N_30084,N_29921,N_28973);
xnor U30085 (N_30085,N_28539,N_29847);
xnor U30086 (N_30086,N_29228,N_28288);
xnor U30087 (N_30087,N_28706,N_28956);
or U30088 (N_30088,N_29757,N_29263);
nor U30089 (N_30089,N_29108,N_28677);
nand U30090 (N_30090,N_29621,N_28264);
xor U30091 (N_30091,N_29739,N_28353);
and U30092 (N_30092,N_28105,N_29149);
and U30093 (N_30093,N_28356,N_28693);
nor U30094 (N_30094,N_29190,N_29408);
xor U30095 (N_30095,N_29900,N_28482);
or U30096 (N_30096,N_28770,N_28370);
xnor U30097 (N_30097,N_29478,N_29209);
nand U30098 (N_30098,N_29951,N_28623);
or U30099 (N_30099,N_29480,N_28745);
or U30100 (N_30100,N_28134,N_28436);
nand U30101 (N_30101,N_28684,N_29923);
nor U30102 (N_30102,N_29067,N_29238);
or U30103 (N_30103,N_28649,N_29779);
nand U30104 (N_30104,N_29744,N_29180);
and U30105 (N_30105,N_28873,N_29202);
xnor U30106 (N_30106,N_29297,N_29917);
xnor U30107 (N_30107,N_29382,N_28740);
xor U30108 (N_30108,N_28325,N_28281);
xor U30109 (N_30109,N_28332,N_29840);
nand U30110 (N_30110,N_28369,N_28512);
xor U30111 (N_30111,N_28803,N_29556);
nor U30112 (N_30112,N_28059,N_28083);
xnor U30113 (N_30113,N_29058,N_29814);
or U30114 (N_30114,N_28152,N_29732);
and U30115 (N_30115,N_28510,N_29025);
xnor U30116 (N_30116,N_29879,N_28729);
and U30117 (N_30117,N_29761,N_28568);
xor U30118 (N_30118,N_29805,N_29501);
and U30119 (N_30119,N_28517,N_28895);
and U30120 (N_30120,N_28617,N_28969);
nor U30121 (N_30121,N_28815,N_29926);
nor U30122 (N_30122,N_28646,N_29243);
xor U30123 (N_30123,N_28493,N_29824);
nand U30124 (N_30124,N_29698,N_29361);
xnor U30125 (N_30125,N_29795,N_29432);
nor U30126 (N_30126,N_29208,N_29563);
nand U30127 (N_30127,N_29300,N_29691);
and U30128 (N_30128,N_29554,N_29796);
nand U30129 (N_30129,N_29862,N_28283);
and U30130 (N_30130,N_29089,N_28792);
or U30131 (N_30131,N_29850,N_29822);
nand U30132 (N_30132,N_28167,N_29919);
nor U30133 (N_30133,N_28487,N_28146);
or U30134 (N_30134,N_29327,N_28273);
and U30135 (N_30135,N_28791,N_28372);
xor U30136 (N_30136,N_28006,N_28978);
xnor U30137 (N_30137,N_29689,N_29424);
or U30138 (N_30138,N_28150,N_29820);
or U30139 (N_30139,N_28499,N_28104);
or U30140 (N_30140,N_28140,N_28801);
or U30141 (N_30141,N_29048,N_28212);
nand U30142 (N_30142,N_28409,N_28099);
xnor U30143 (N_30143,N_29249,N_29032);
xor U30144 (N_30144,N_28435,N_29258);
or U30145 (N_30145,N_28060,N_29861);
xnor U30146 (N_30146,N_29317,N_28502);
or U30147 (N_30147,N_29677,N_28095);
xnor U30148 (N_30148,N_28079,N_29753);
xor U30149 (N_30149,N_29530,N_29950);
xor U30150 (N_30150,N_29475,N_28147);
and U30151 (N_30151,N_28560,N_28931);
or U30152 (N_30152,N_28767,N_29776);
and U30153 (N_30153,N_29598,N_29937);
nand U30154 (N_30154,N_28223,N_28511);
nor U30155 (N_30155,N_28622,N_29188);
nor U30156 (N_30156,N_28206,N_28383);
nand U30157 (N_30157,N_28284,N_28028);
and U30158 (N_30158,N_29521,N_29366);
and U30159 (N_30159,N_28169,N_28814);
or U30160 (N_30160,N_28929,N_28933);
or U30161 (N_30161,N_29808,N_29274);
and U30162 (N_30162,N_28580,N_29977);
and U30163 (N_30163,N_29999,N_29819);
xnor U30164 (N_30164,N_29542,N_28869);
nand U30165 (N_30165,N_29070,N_28208);
nand U30166 (N_30166,N_29639,N_29363);
and U30167 (N_30167,N_28821,N_28655);
xnor U30168 (N_30168,N_28637,N_28529);
or U30169 (N_30169,N_28691,N_28769);
or U30170 (N_30170,N_28806,N_29527);
nand U30171 (N_30171,N_29685,N_29371);
nor U30172 (N_30172,N_29536,N_28970);
nor U30173 (N_30173,N_29040,N_29155);
nor U30174 (N_30174,N_28963,N_28640);
nor U30175 (N_30175,N_28524,N_29081);
and U30176 (N_30176,N_29665,N_29232);
nor U30177 (N_30177,N_28976,N_28925);
and U30178 (N_30178,N_28003,N_29303);
or U30179 (N_30179,N_29252,N_28913);
nand U30180 (N_30180,N_28017,N_29318);
and U30181 (N_30181,N_28666,N_29749);
and U30182 (N_30182,N_28457,N_29577);
or U30183 (N_30183,N_29623,N_28016);
nor U30184 (N_30184,N_29888,N_29570);
nand U30185 (N_30185,N_28228,N_29358);
xor U30186 (N_30186,N_29309,N_28946);
nand U30187 (N_30187,N_29953,N_29462);
nor U30188 (N_30188,N_29965,N_29602);
or U30189 (N_30189,N_29375,N_29455);
nand U30190 (N_30190,N_28522,N_28421);
or U30191 (N_30191,N_28519,N_28112);
or U30192 (N_30192,N_28251,N_29370);
and U30193 (N_30193,N_28426,N_29833);
or U30194 (N_30194,N_28615,N_29066);
or U30195 (N_30195,N_29519,N_28709);
nand U30196 (N_30196,N_28097,N_29981);
or U30197 (N_30197,N_28362,N_28050);
nor U30198 (N_30198,N_29930,N_29581);
xnor U30199 (N_30199,N_29244,N_29829);
or U30200 (N_30200,N_28106,N_29420);
and U30201 (N_30201,N_28696,N_29748);
xor U30202 (N_30202,N_28921,N_28117);
nand U30203 (N_30203,N_29254,N_29713);
xor U30204 (N_30204,N_28398,N_29535);
xor U30205 (N_30205,N_29486,N_29747);
nor U30206 (N_30206,N_29770,N_29655);
or U30207 (N_30207,N_29021,N_29611);
nor U30208 (N_30208,N_29794,N_28047);
xor U30209 (N_30209,N_28906,N_29214);
nand U30210 (N_30210,N_29349,N_28465);
nand U30211 (N_30211,N_28191,N_28304);
nor U30212 (N_30212,N_29955,N_29215);
nand U30213 (N_30213,N_28243,N_28350);
and U30214 (N_30214,N_28605,N_28088);
nor U30215 (N_30215,N_28999,N_29520);
nor U30216 (N_30216,N_28532,N_29072);
and U30217 (N_30217,N_29599,N_29163);
xnor U30218 (N_30218,N_28172,N_28305);
and U30219 (N_30219,N_28822,N_29088);
xnor U30220 (N_30220,N_28773,N_29391);
and U30221 (N_30221,N_29377,N_28538);
or U30222 (N_30222,N_28872,N_29138);
xor U30223 (N_30223,N_29696,N_29392);
or U30224 (N_30224,N_28781,N_29401);
nand U30225 (N_30225,N_28788,N_29492);
or U30226 (N_30226,N_29606,N_29760);
nand U30227 (N_30227,N_29927,N_28239);
nand U30228 (N_30228,N_29440,N_29267);
nor U30229 (N_30229,N_28128,N_29076);
xnor U30230 (N_30230,N_29052,N_28625);
nand U30231 (N_30231,N_29347,N_29311);
or U30232 (N_30232,N_28660,N_29225);
and U30233 (N_30233,N_29531,N_28977);
or U30234 (N_30234,N_28996,N_28038);
nand U30235 (N_30235,N_28109,N_28936);
xnor U30236 (N_30236,N_29102,N_28214);
or U30237 (N_30237,N_29079,N_28892);
xor U30238 (N_30238,N_28636,N_29818);
nand U30239 (N_30239,N_29650,N_28780);
and U30240 (N_30240,N_29134,N_29857);
nand U30241 (N_30241,N_29708,N_29826);
nand U30242 (N_30242,N_29771,N_28797);
and U30243 (N_30243,N_28951,N_29470);
nor U30244 (N_30244,N_28087,N_29435);
xnor U30245 (N_30245,N_29278,N_28222);
and U30246 (N_30246,N_29116,N_29041);
xor U30247 (N_30247,N_28588,N_29175);
xnor U30248 (N_30248,N_29684,N_29464);
nor U30249 (N_30249,N_28796,N_29451);
nor U30250 (N_30250,N_28361,N_28474);
or U30251 (N_30251,N_29157,N_28894);
nor U30252 (N_30252,N_29240,N_29114);
nor U30253 (N_30253,N_29712,N_29150);
xor U30254 (N_30254,N_29667,N_29666);
or U30255 (N_30255,N_28012,N_29304);
nor U30256 (N_30256,N_29473,N_28725);
and U30257 (N_30257,N_28441,N_29644);
nand U30258 (N_30258,N_28755,N_29904);
nor U30259 (N_30259,N_28690,N_28863);
nor U30260 (N_30260,N_28248,N_29026);
or U30261 (N_30261,N_28783,N_28396);
and U30262 (N_30262,N_29411,N_29288);
and U30263 (N_30263,N_28364,N_28328);
nand U30264 (N_30264,N_29601,N_28685);
and U30265 (N_30265,N_29809,N_29669);
or U30266 (N_30266,N_28897,N_29484);
nand U30267 (N_30267,N_29446,N_28753);
nand U30268 (N_30268,N_29176,N_29193);
xor U30269 (N_30269,N_29164,N_29165);
nor U30270 (N_30270,N_29364,N_28439);
or U30271 (N_30271,N_29793,N_28726);
xnor U30272 (N_30272,N_29383,N_28149);
nand U30273 (N_30273,N_29963,N_29500);
nand U30274 (N_30274,N_29063,N_28229);
or U30275 (N_30275,N_28262,N_28874);
nor U30276 (N_30276,N_29830,N_29777);
nand U30277 (N_30277,N_28846,N_28671);
and U30278 (N_30278,N_28834,N_28754);
nor U30279 (N_30279,N_29626,N_28041);
and U30280 (N_30280,N_29028,N_28489);
nor U30281 (N_30281,N_28997,N_29907);
nand U30282 (N_30282,N_28478,N_29973);
and U30283 (N_30283,N_29103,N_29434);
xnor U30284 (N_30284,N_29452,N_29365);
or U30285 (N_30285,N_28496,N_28454);
nand U30286 (N_30286,N_29471,N_28296);
or U30287 (N_30287,N_28673,N_28271);
xnor U30288 (N_30288,N_29697,N_29630);
nand U30289 (N_30289,N_29008,N_29920);
nand U30290 (N_30290,N_29186,N_28579);
xor U30291 (N_30291,N_29518,N_28741);
nor U30292 (N_30292,N_29498,N_28422);
and U30293 (N_30293,N_29331,N_28187);
nand U30294 (N_30294,N_28899,N_28807);
xnor U30295 (N_30295,N_29695,N_29234);
xnor U30296 (N_30296,N_29458,N_28358);
xor U30297 (N_30297,N_29791,N_28413);
xnor U30298 (N_30298,N_29001,N_28573);
or U30299 (N_30299,N_28267,N_29346);
nor U30300 (N_30300,N_28937,N_29915);
and U30301 (N_30301,N_29526,N_28838);
and U30302 (N_30302,N_29936,N_28547);
nand U30303 (N_30303,N_28324,N_29198);
xnor U30304 (N_30304,N_29362,N_29142);
and U30305 (N_30305,N_29837,N_29891);
or U30306 (N_30306,N_28136,N_28712);
and U30307 (N_30307,N_28911,N_29709);
and U30308 (N_30308,N_28485,N_28809);
or U30309 (N_30309,N_29417,N_28042);
nor U30310 (N_30310,N_28463,N_28345);
nor U30311 (N_30311,N_28774,N_29958);
or U30312 (N_30312,N_28001,N_28089);
nor U30313 (N_30313,N_28902,N_28680);
nor U30314 (N_30314,N_28476,N_28699);
nor U30315 (N_30315,N_29495,N_28983);
nand U30316 (N_30316,N_28475,N_29427);
and U30317 (N_30317,N_29047,N_28708);
and U30318 (N_30318,N_28692,N_29169);
nand U30319 (N_30319,N_29250,N_28302);
nand U30320 (N_30320,N_29550,N_28366);
xnor U30321 (N_30321,N_28310,N_28077);
or U30322 (N_30322,N_29015,N_29725);
nor U30323 (N_30323,N_28824,N_29849);
nand U30324 (N_30324,N_28918,N_28805);
nor U30325 (N_30325,N_28055,N_29816);
nand U30326 (N_30326,N_28835,N_29568);
or U30327 (N_30327,N_28392,N_28942);
nand U30328 (N_30328,N_29658,N_29046);
and U30329 (N_30329,N_29784,N_28849);
nor U30330 (N_30330,N_29135,N_29848);
or U30331 (N_30331,N_28562,N_29009);
xor U30332 (N_30332,N_28082,N_28051);
xnor U30333 (N_30333,N_29686,N_28058);
nor U30334 (N_30334,N_29136,N_29972);
nor U30335 (N_30335,N_29711,N_28985);
or U30336 (N_30336,N_29384,N_29171);
or U30337 (N_30337,N_28683,N_29141);
or U30338 (N_30338,N_29680,N_29604);
xor U30339 (N_30339,N_29859,N_28081);
xnor U30340 (N_30340,N_28488,N_28832);
nand U30341 (N_30341,N_29738,N_28893);
and U30342 (N_30342,N_29918,N_28148);
and U30343 (N_30343,N_28495,N_29087);
nand U30344 (N_30344,N_28261,N_29160);
nand U30345 (N_30345,N_29031,N_28154);
nand U30346 (N_30346,N_28098,N_28269);
and U30347 (N_30347,N_29742,N_28279);
nor U30348 (N_30348,N_29552,N_28407);
or U30349 (N_30349,N_28275,N_29469);
and U30350 (N_30350,N_28775,N_29553);
and U30351 (N_30351,N_28828,N_29315);
nor U30352 (N_30352,N_28241,N_29995);
nand U30353 (N_30353,N_29673,N_29109);
xnor U30354 (N_30354,N_28584,N_28371);
nand U30355 (N_30355,N_28244,N_28987);
or U30356 (N_30356,N_28757,N_28861);
nor U30357 (N_30357,N_28979,N_28526);
nand U30358 (N_30358,N_28013,N_28292);
nor U30359 (N_30359,N_28581,N_29838);
and U30360 (N_30360,N_29528,N_29864);
xor U30361 (N_30361,N_28141,N_29266);
or U30362 (N_30362,N_28375,N_29654);
xnor U30363 (N_30363,N_29339,N_28595);
xnor U30364 (N_30364,N_28746,N_29797);
nor U30365 (N_30365,N_28367,N_29335);
or U30366 (N_30366,N_29516,N_28204);
xnor U30367 (N_30367,N_29236,N_29120);
nor U30368 (N_30368,N_29651,N_29126);
xnor U30369 (N_30369,N_29781,N_29034);
or U30370 (N_30370,N_28827,N_28319);
nor U30371 (N_30371,N_28068,N_29078);
nor U30372 (N_30372,N_28575,N_29239);
xnor U30373 (N_30373,N_29074,N_29913);
or U30374 (N_30374,N_28491,N_28388);
nor U30375 (N_30375,N_29688,N_28718);
nand U30376 (N_30376,N_28552,N_28880);
nand U30377 (N_30377,N_29312,N_29584);
xnor U30378 (N_30378,N_28322,N_29286);
nor U30379 (N_30379,N_29284,N_28467);
xor U30380 (N_30380,N_28924,N_29121);
and U30381 (N_30381,N_29714,N_29110);
xnor U30382 (N_30382,N_28311,N_28414);
and U30383 (N_30383,N_29298,N_28850);
xor U30384 (N_30384,N_28779,N_28245);
nand U30385 (N_30385,N_29412,N_28549);
nor U30386 (N_30386,N_29737,N_29082);
nor U30387 (N_30387,N_28170,N_28201);
xnor U30388 (N_30388,N_28005,N_28234);
xnor U30389 (N_30389,N_29127,N_28408);
or U30390 (N_30390,N_28972,N_28694);
and U30391 (N_30391,N_29069,N_29752);
xnor U30392 (N_30392,N_28256,N_28614);
nand U30393 (N_30393,N_28096,N_29968);
nor U30394 (N_30394,N_29416,N_29902);
nand U30395 (N_30395,N_29705,N_29050);
nand U30396 (N_30396,N_28558,N_28207);
or U30397 (N_30397,N_29592,N_28069);
nor U30398 (N_30398,N_29523,N_28403);
nor U30399 (N_30399,N_28619,N_28306);
or U30400 (N_30400,N_29117,N_29889);
or U30401 (N_30401,N_28255,N_28515);
xnor U30402 (N_30402,N_29337,N_28216);
or U30403 (N_30403,N_29287,N_28889);
or U30404 (N_30404,N_28871,N_29990);
nand U30405 (N_30405,N_29723,N_29743);
xor U30406 (N_30406,N_28715,N_28765);
xnor U30407 (N_30407,N_28751,N_28732);
xor U30408 (N_30408,N_29494,N_29373);
or U30409 (N_30409,N_29111,N_29821);
nand U30410 (N_30410,N_29546,N_29355);
xnor U30411 (N_30411,N_28784,N_29942);
and U30412 (N_30412,N_28247,N_28115);
xnor U30413 (N_30413,N_29368,N_28545);
xor U30414 (N_30414,N_29242,N_29077);
nor U30415 (N_30415,N_29502,N_29273);
nor U30416 (N_30416,N_28352,N_29998);
xor U30417 (N_30417,N_28600,N_29567);
or U30418 (N_30418,N_29018,N_29896);
nand U30419 (N_30419,N_29947,N_28820);
and U30420 (N_30420,N_29622,N_28862);
and U30421 (N_30421,N_29569,N_28107);
and U30422 (N_30422,N_29813,N_29179);
nand U30423 (N_30423,N_29454,N_28303);
or U30424 (N_30424,N_29575,N_29901);
nand U30425 (N_30425,N_28866,N_29139);
or U30426 (N_30426,N_29100,N_28520);
nand U30427 (N_30427,N_29856,N_29086);
and U30428 (N_30428,N_28811,N_29159);
xor U30429 (N_30429,N_29385,N_29006);
nor U30430 (N_30430,N_28586,N_28940);
nor U30431 (N_30431,N_29969,N_29675);
and U30432 (N_30432,N_28257,N_29378);
and U30433 (N_30433,N_28582,N_28971);
and U30434 (N_30434,N_29130,N_28067);
xnor U30435 (N_30435,N_28503,N_28459);
or U30436 (N_30436,N_28365,N_29294);
xor U30437 (N_30437,N_29674,N_29299);
nand U30438 (N_30438,N_29997,N_29683);
xor U30439 (N_30439,N_29724,N_28653);
nand U30440 (N_30440,N_29011,N_28711);
xor U30441 (N_30441,N_29768,N_28108);
xor U30442 (N_30442,N_28425,N_29756);
and U30443 (N_30443,N_28142,N_29101);
and U30444 (N_30444,N_29634,N_28200);
xor U30445 (N_30445,N_28018,N_29605);
xnor U30446 (N_30446,N_28347,N_29836);
or U30447 (N_30447,N_28852,N_29869);
xnor U30448 (N_30448,N_28737,N_29113);
nand U30449 (N_30449,N_28825,N_29996);
nor U30450 (N_30450,N_29846,N_28613);
or U30451 (N_30451,N_29415,N_29872);
or U30452 (N_30452,N_28597,N_28950);
and U30453 (N_30453,N_29166,N_28492);
and U30454 (N_30454,N_29143,N_29627);
nor U30455 (N_30455,N_28905,N_29852);
or U30456 (N_30456,N_28094,N_28379);
or U30457 (N_30457,N_29459,N_29068);
nor U30458 (N_30458,N_29184,N_28382);
and U30459 (N_30459,N_28631,N_29798);
xnor U30460 (N_30460,N_28213,N_29505);
or U30461 (N_30461,N_28556,N_29587);
or U30462 (N_30462,N_28070,N_29213);
and U30463 (N_30463,N_28635,N_29007);
nor U30464 (N_30464,N_29728,N_29801);
nor U30465 (N_30465,N_29393,N_29477);
xnor U30466 (N_30466,N_28749,N_28943);
nor U30467 (N_30467,N_29931,N_29221);
and U30468 (N_30468,N_28563,N_28953);
or U30469 (N_30469,N_29759,N_28447);
xnor U30470 (N_30470,N_28205,N_28315);
nor U30471 (N_30471,N_28182,N_28968);
xnor U30472 (N_30472,N_29509,N_28896);
and U30473 (N_30473,N_29887,N_28101);
nand U30474 (N_30474,N_28080,N_29197);
nor U30475 (N_30475,N_28599,N_28736);
nor U30476 (N_30476,N_28225,N_28610);
nand U30477 (N_30477,N_29875,N_28842);
nand U30478 (N_30478,N_28831,N_28554);
xor U30479 (N_30479,N_29693,N_28156);
or U30480 (N_30480,N_28567,N_28543);
xor U30481 (N_30481,N_29992,N_28193);
nor U30482 (N_30482,N_28508,N_29983);
nand U30483 (N_30483,N_29628,N_29740);
and U30484 (N_30484,N_28505,N_29617);
xor U30485 (N_30485,N_29409,N_28587);
xnor U30486 (N_30486,N_29196,N_29097);
or U30487 (N_30487,N_29316,N_28010);
nor U30488 (N_30488,N_29430,N_28078);
nand U30489 (N_30489,N_28758,N_28061);
and U30490 (N_30490,N_28286,N_29572);
nand U30491 (N_30491,N_29168,N_29443);
nand U30492 (N_30492,N_29597,N_29181);
xnor U30493 (N_30493,N_29448,N_29720);
and U30494 (N_30494,N_29183,N_29595);
and U30495 (N_30495,N_29125,N_28135);
xor U30496 (N_30496,N_29591,N_28460);
or U30497 (N_30497,N_28639,N_28395);
nand U30498 (N_30498,N_28026,N_28266);
xor U30499 (N_30499,N_29463,N_29676);
nand U30500 (N_30500,N_28993,N_28728);
nor U30501 (N_30501,N_28589,N_29129);
xnor U30502 (N_30502,N_29016,N_28602);
or U30503 (N_30503,N_28131,N_28308);
and U30504 (N_30504,N_29976,N_28721);
and U30505 (N_30505,N_28415,N_29096);
nand U30506 (N_30506,N_29678,N_29679);
or U30507 (N_30507,N_29301,N_29802);
nand U30508 (N_30508,N_29207,N_29340);
nand U30509 (N_30509,N_29508,N_28103);
nor U30510 (N_30510,N_29525,N_29224);
xnor U30511 (N_30511,N_28287,N_28738);
or U30512 (N_30512,N_29195,N_29313);
nor U30513 (N_30513,N_28052,N_29019);
nand U30514 (N_30514,N_29690,N_29490);
nand U30515 (N_30515,N_29276,N_29539);
xor U30516 (N_30516,N_28988,N_29694);
nand U30517 (N_30517,N_29445,N_29903);
or U30518 (N_30518,N_29638,N_29115);
nor U30519 (N_30519,N_29912,N_28272);
or U30520 (N_30520,N_28764,N_29406);
and U30521 (N_30521,N_28934,N_29993);
or U30522 (N_30522,N_29153,N_29226);
nor U30523 (N_30523,N_29418,N_29560);
nand U30524 (N_30524,N_28360,N_28904);
xnor U30525 (N_30525,N_29562,N_28336);
or U30526 (N_30526,N_28298,N_29868);
xor U30527 (N_30527,N_28752,N_29005);
nor U30528 (N_30528,N_28044,N_28611);
nand U30529 (N_30529,N_29767,N_28965);
nand U30530 (N_30530,N_29423,N_28220);
or U30531 (N_30531,N_29608,N_28714);
and U30532 (N_30532,N_28535,N_28119);
or U30533 (N_30533,N_28944,N_29162);
nand U30534 (N_30534,N_28466,N_29330);
nor U30535 (N_30535,N_29147,N_28157);
xor U30536 (N_30536,N_29841,N_28400);
nand U30537 (N_30537,N_29722,N_28217);
xnor U30538 (N_30538,N_28092,N_28129);
xnor U30539 (N_30539,N_28506,N_28618);
nor U30540 (N_30540,N_29899,N_28724);
nor U30541 (N_30541,N_28434,N_28494);
xor U30542 (N_30542,N_28263,N_29039);
or U30543 (N_30543,N_29629,N_29217);
nand U30544 (N_30544,N_28484,N_29940);
or U30545 (N_30545,N_29241,N_28591);
nand U30546 (N_30546,N_29682,N_28645);
xor U30547 (N_30547,N_29637,N_28667);
nor U30548 (N_30548,N_28593,N_29194);
nor U30549 (N_30549,N_29561,N_29600);
and U30550 (N_30550,N_28437,N_28500);
and U30551 (N_30551,N_28030,N_28155);
or U30552 (N_30552,N_28230,N_28354);
nor U30553 (N_30553,N_28163,N_28578);
xnor U30554 (N_30554,N_29437,N_28594);
nand U30555 (N_30555,N_28174,N_29959);
and U30556 (N_30556,N_29898,N_28540);
nand U30557 (N_30557,N_29769,N_28514);
nand U30558 (N_30558,N_28716,N_29717);
nor U30559 (N_30559,N_29538,N_29729);
or U30560 (N_30560,N_29799,N_29710);
or U30561 (N_30561,N_28819,N_29481);
or U30562 (N_30562,N_28975,N_29515);
or U30563 (N_30563,N_29586,N_29544);
nor U30564 (N_30564,N_28110,N_29582);
or U30565 (N_30565,N_28498,N_29594);
or U30566 (N_30566,N_29946,N_29460);
nor U30567 (N_30567,N_29928,N_28789);
nor U30568 (N_30568,N_28702,N_28935);
xnor U30569 (N_30569,N_29027,N_29641);
and U30570 (N_30570,N_29979,N_28960);
nand U30571 (N_30571,N_29185,N_28962);
nand U30572 (N_30572,N_28211,N_28268);
xnor U30573 (N_30573,N_28994,N_29935);
xnor U30574 (N_30574,N_29754,N_28816);
or U30575 (N_30575,N_28008,N_28525);
nor U30576 (N_30576,N_29943,N_29715);
xnor U30577 (N_30577,N_29534,N_29003);
xor U30578 (N_30578,N_28707,N_29716);
and U30579 (N_30579,N_29144,N_28875);
or U30580 (N_30580,N_28812,N_29425);
xnor U30581 (N_30581,N_29132,N_29895);
nand U30582 (N_30582,N_29354,N_29699);
xor U30583 (N_30583,N_29878,N_28561);
and U30584 (N_30584,N_28912,N_29706);
nand U30585 (N_30585,N_29545,N_29800);
or U30586 (N_30586,N_28853,N_28032);
nor U30587 (N_30587,N_29212,N_29825);
nand U30588 (N_30588,N_29524,N_28470);
nand U30589 (N_30589,N_28598,N_28086);
xor U30590 (N_30590,N_29305,N_29944);
nand U30591 (N_30591,N_28900,N_28443);
and U30592 (N_30592,N_28884,N_28652);
nor U30593 (N_30593,N_29886,N_28719);
nor U30594 (N_30594,N_29308,N_29772);
xnor U30595 (N_30595,N_29994,N_29949);
nand U30596 (N_30596,N_28885,N_28674);
nor U30597 (N_30597,N_28034,N_29291);
nor U30598 (N_30598,N_29204,N_29152);
nand U30599 (N_30599,N_29865,N_28374);
nor U30600 (N_30600,N_29510,N_28833);
xnor U30601 (N_30601,N_28793,N_28238);
xnor U30602 (N_30602,N_28293,N_28397);
nand U30603 (N_30603,N_29388,N_28548);
or U30604 (N_30604,N_29557,N_28002);
or U30605 (N_30605,N_28159,N_29272);
and U30606 (N_30606,N_28164,N_28386);
nand U30607 (N_30607,N_28847,N_28995);
and U30608 (N_30608,N_28858,N_28258);
and U30609 (N_30609,N_28813,N_28882);
xor U30610 (N_30610,N_28254,N_28901);
or U30611 (N_30611,N_28818,N_28464);
and U30612 (N_30612,N_29974,N_29573);
xnor U30613 (N_30613,N_29503,N_28542);
xor U30614 (N_30614,N_28695,N_29203);
nand U30615 (N_30615,N_28472,N_29866);
and U30616 (N_30616,N_29222,N_29513);
and U30617 (N_30617,N_29613,N_29877);
nor U30618 (N_30618,N_29961,N_29882);
or U30619 (N_30619,N_28830,N_28859);
and U30620 (N_30620,N_28787,N_29479);
xnor U30621 (N_30621,N_29541,N_29223);
nor U30622 (N_30622,N_28608,N_29952);
or U30623 (N_30623,N_29532,N_28682);
and U30624 (N_30624,N_28848,N_28132);
nand U30625 (N_30625,N_29707,N_28442);
xnor U30626 (N_30626,N_29199,N_29780);
nand U30627 (N_30627,N_28151,N_28423);
nand U30628 (N_30628,N_29247,N_28569);
and U30629 (N_30629,N_28091,N_28864);
or U30630 (N_30630,N_28555,N_28654);
and U30631 (N_30631,N_28744,N_28194);
nand U30632 (N_30632,N_28881,N_29975);
nor U30633 (N_30633,N_29811,N_28318);
xor U30634 (N_30634,N_29971,N_28665);
or U30635 (N_30635,N_29774,N_28176);
nor U30636 (N_30636,N_28772,N_29485);
nor U30637 (N_30637,N_29098,N_28390);
xnor U30638 (N_30638,N_28616,N_29962);
xor U30639 (N_30639,N_28688,N_29646);
or U30640 (N_30640,N_29786,N_28461);
or U30641 (N_30641,N_28226,N_28733);
and U30642 (N_30642,N_28887,N_28160);
xnor U30643 (N_30643,N_29734,N_28120);
and U30644 (N_30644,N_28346,N_29413);
nor U30645 (N_30645,N_28331,N_29985);
nor U30646 (N_30646,N_28840,N_29730);
or U30647 (N_30647,N_29173,N_28453);
nand U30648 (N_30648,N_29967,N_29897);
nor U30649 (N_30649,N_28590,N_28760);
xnor U30650 (N_30650,N_29428,N_29306);
xnor U30651 (N_30651,N_28886,N_29792);
or U30652 (N_30652,N_28536,N_29580);
nor U30653 (N_30653,N_28865,N_28703);
nor U30654 (N_30654,N_28049,N_28659);
nor U30655 (N_30655,N_29038,N_28632);
or U30656 (N_30656,N_29764,N_29419);
xor U30657 (N_30657,N_29934,N_28177);
nor U30658 (N_30658,N_29439,N_28570);
xor U30659 (N_30659,N_29353,N_29328);
and U30660 (N_30660,N_28473,N_28122);
or U30661 (N_30661,N_29653,N_29051);
and U30662 (N_30662,N_28468,N_28748);
xnor U30663 (N_30663,N_28307,N_28198);
nor U30664 (N_30664,N_28984,N_28687);
or U30665 (N_30665,N_29890,N_28197);
nor U30666 (N_30666,N_29004,N_29379);
xnor U30667 (N_30667,N_29270,N_28381);
or U30668 (N_30668,N_28601,N_28877);
and U30669 (N_30669,N_29085,N_28171);
nor U30670 (N_30670,N_28776,N_29657);
and U30671 (N_30671,N_29522,N_28250);
nor U30672 (N_30672,N_28385,N_28242);
and U30673 (N_30673,N_28698,N_28161);
nand U30674 (N_30674,N_29788,N_28991);
and U30675 (N_30675,N_29547,N_29514);
xor U30676 (N_30676,N_28114,N_28072);
nand U30677 (N_30677,N_29467,N_29945);
nor U30678 (N_30678,N_28648,N_29731);
and U30679 (N_30679,N_28841,N_28981);
nor U30680 (N_30680,N_29036,N_29548);
nor U30681 (N_30681,N_29565,N_28604);
nand U30682 (N_30682,N_28127,N_29281);
or U30683 (N_30683,N_28179,N_29652);
nor U30684 (N_30684,N_29262,N_28329);
nand U30685 (N_30685,N_29566,N_29029);
xor U30686 (N_30686,N_28668,N_29892);
nand U30687 (N_30687,N_28011,N_28851);
or U30688 (N_30688,N_29755,N_28339);
and U30689 (N_30689,N_29647,N_28290);
xor U30690 (N_30690,N_28100,N_28947);
or U30691 (N_30691,N_29061,N_29119);
and U30692 (N_30692,N_28641,N_28518);
and U30693 (N_30693,N_29177,N_29719);
and U30694 (N_30694,N_28914,N_28928);
or U30695 (N_30695,N_29910,N_29320);
nor U30696 (N_30696,N_29128,N_28759);
nand U30697 (N_30697,N_29555,N_28927);
or U30698 (N_30698,N_29091,N_29987);
nand U30699 (N_30699,N_28670,N_29075);
nor U30700 (N_30700,N_28855,N_29982);
nor U30701 (N_30701,N_29668,N_28483);
nor U30702 (N_30702,N_28771,N_29881);
nor U30703 (N_30703,N_28253,N_28316);
nor U30704 (N_30704,N_28523,N_29559);
nand U30705 (N_30705,N_28908,N_29472);
xnor U30706 (N_30706,N_28627,N_29663);
xor U30707 (N_30707,N_29506,N_29341);
or U30708 (N_30708,N_28471,N_29431);
and U30709 (N_30709,N_29055,N_29099);
nand U30710 (N_30710,N_29380,N_29736);
or U30711 (N_30711,N_29783,N_28720);
nand U30712 (N_30712,N_28630,N_29733);
nor U30713 (N_30713,N_29381,N_29854);
nand U30714 (N_30714,N_28986,N_29703);
and U30715 (N_30715,N_28188,N_29131);
and U30716 (N_30716,N_28121,N_29465);
nor U30717 (N_30717,N_28451,N_28043);
and U30718 (N_30718,N_28786,N_28676);
or U30719 (N_30719,N_28233,N_28056);
nand U30720 (N_30720,N_29571,N_29302);
nand U30721 (N_30721,N_28430,N_28162);
or U30722 (N_30722,N_28196,N_28531);
or U30723 (N_30723,N_28939,N_28644);
or U30724 (N_30724,N_28138,N_29429);
nand U30725 (N_30725,N_28246,N_29421);
nand U30726 (N_30726,N_29989,N_29758);
or U30727 (N_30727,N_28195,N_28909);
xnor U30728 (N_30728,N_29133,N_29812);
or U30729 (N_30729,N_28084,N_29894);
xnor U30730 (N_30730,N_28628,N_28823);
xnor U30731 (N_30731,N_28359,N_28378);
nor U30732 (N_30732,N_28550,N_29290);
and U30733 (N_30733,N_28009,N_28402);
or U30734 (N_30734,N_28585,N_28651);
xor U30735 (N_30735,N_29118,N_28462);
nor U30736 (N_30736,N_28957,N_28368);
nor U30737 (N_30737,N_28898,N_28559);
or U30738 (N_30738,N_29307,N_29925);
nand U30739 (N_30739,N_29832,N_28612);
or U30740 (N_30740,N_29106,N_29269);
nand U30741 (N_30741,N_28189,N_28301);
nand U30742 (N_30742,N_29329,N_28490);
and U30743 (N_30743,N_28438,N_29596);
and U30744 (N_30744,N_28165,N_29625);
nor U30745 (N_30745,N_29350,N_28046);
or U30746 (N_30746,N_29880,N_28527);
nand U30747 (N_30747,N_28015,N_28890);
xor U30748 (N_30748,N_28565,N_28384);
nand U30749 (N_30749,N_28215,N_28076);
nand U30750 (N_30750,N_28294,N_28090);
nand U30751 (N_30751,N_29885,N_29107);
nor U30752 (N_30752,N_28798,N_28763);
nor U30753 (N_30753,N_28313,N_28184);
xnor U30754 (N_30754,N_28260,N_29292);
and U30755 (N_30755,N_29593,N_28777);
nor U30756 (N_30756,N_28742,N_29333);
nor U30757 (N_30757,N_28357,N_29043);
nand U30758 (N_30758,N_28126,N_29310);
xnor U30759 (N_30759,N_28130,N_29870);
xor U30760 (N_30760,N_28181,N_29620);
nand U30761 (N_30761,N_29750,N_28856);
and U30762 (N_30762,N_28202,N_29908);
xor U30763 (N_30763,N_29718,N_29681);
nand U30764 (N_30764,N_29414,N_28387);
nand U30765 (N_30765,N_28428,N_28066);
nand U30766 (N_30766,N_28802,N_28285);
nand U30767 (N_30767,N_28023,N_29064);
nor U30768 (N_30768,N_29140,N_28399);
nand U30769 (N_30769,N_29970,N_28405);
xor U30770 (N_30770,N_28173,N_28917);
and U30771 (N_30771,N_29390,N_28185);
and U30772 (N_30772,N_29671,N_28961);
and U30773 (N_30773,N_29271,N_29905);
and U30774 (N_30774,N_28320,N_28537);
nor U30775 (N_30775,N_29137,N_29551);
or U30776 (N_30776,N_29504,N_28282);
nand U30777 (N_30777,N_28731,N_28530);
xor U30778 (N_30778,N_29167,N_29789);
nor U30779 (N_30779,N_28700,N_29037);
and U30780 (N_30780,N_29704,N_29255);
xor U30781 (N_30781,N_29104,N_29721);
nand U30782 (N_30782,N_29348,N_29403);
or U30783 (N_30783,N_28449,N_28143);
xnor U30784 (N_30784,N_28333,N_28992);
or U30785 (N_30785,N_29476,N_28064);
nor U30786 (N_30786,N_29489,N_29564);
or U30787 (N_30787,N_29123,N_29145);
nor U30788 (N_30788,N_28528,N_28952);
nand U30789 (N_30789,N_28633,N_28689);
nand U30790 (N_30790,N_28672,N_28903);
or U30791 (N_30791,N_29635,N_28326);
and U30792 (N_30792,N_29860,N_28727);
xnor U30793 (N_30793,N_28183,N_29206);
xor U30794 (N_30794,N_28317,N_29205);
xor U30795 (N_30795,N_29261,N_29071);
and U30796 (N_30796,N_28486,N_29323);
and U30797 (N_30797,N_29456,N_29326);
nand U30798 (N_30798,N_28377,N_28982);
xor U30799 (N_30799,N_28458,N_28062);
and U30800 (N_30800,N_28277,N_28349);
nor U30801 (N_30801,N_29615,N_28907);
nor U30802 (N_30802,N_28643,N_29342);
xnor U30803 (N_30803,N_28063,N_28085);
or U30804 (N_30804,N_28199,N_28418);
nor U30805 (N_30805,N_29616,N_28024);
or U30806 (N_30806,N_29609,N_29189);
nand U30807 (N_30807,N_28868,N_28420);
nand U30808 (N_30808,N_28998,N_29461);
and U30809 (N_30809,N_28888,N_29410);
xor U30810 (N_30810,N_28620,N_28004);
or U30811 (N_30811,N_29049,N_29876);
or U30812 (N_30812,N_29444,N_29324);
xnor U30813 (N_30813,N_29345,N_29803);
nor U30814 (N_30814,N_28955,N_28040);
nor U30815 (N_30815,N_28036,N_29161);
nand U30816 (N_30816,N_28389,N_29497);
xnor U30817 (N_30817,N_28980,N_28954);
nand U30818 (N_30818,N_28959,N_29762);
or U30819 (N_30819,N_29858,N_29182);
and U30820 (N_30820,N_29090,N_28705);
or U30821 (N_30821,N_29585,N_28876);
and U30822 (N_30822,N_29782,N_28299);
and U30823 (N_30823,N_29540,N_28860);
nor U30824 (N_30824,N_28938,N_28949);
and U30825 (N_30825,N_28576,N_28029);
or U30826 (N_30826,N_28678,N_29220);
xnor U30827 (N_30827,N_28571,N_28452);
or U30828 (N_30828,N_29386,N_29612);
nand U30829 (N_30829,N_29778,N_28124);
nand U30830 (N_30830,N_29394,N_28376);
or U30831 (N_30831,N_28075,N_28629);
xor U30832 (N_30832,N_29643,N_29360);
and U30833 (N_30833,N_28323,N_29277);
or U30834 (N_30834,N_29956,N_29065);
or U30835 (N_30835,N_29583,N_29289);
xnor U30836 (N_30836,N_29831,N_28432);
or U30837 (N_30837,N_28845,N_29763);
nor U30838 (N_30838,N_29426,N_28661);
nand U30839 (N_30839,N_29268,N_29325);
and U30840 (N_30840,N_28544,N_29988);
and U30841 (N_30841,N_28501,N_28259);
and U30842 (N_30842,N_29122,N_28252);
and U30843 (N_30843,N_29084,N_28891);
nor U30844 (N_30844,N_28723,N_29589);
nand U30845 (N_30845,N_28133,N_29356);
nor U30846 (N_30846,N_29010,N_29828);
and U30847 (N_30847,N_29670,N_28794);
and U30848 (N_30848,N_29148,N_28810);
nand U30849 (N_30849,N_29924,N_29344);
and U30850 (N_30850,N_29369,N_28658);
and U30851 (N_30851,N_28870,N_29259);
or U30852 (N_30852,N_29033,N_29398);
or U30853 (N_30853,N_28404,N_28020);
nor U30854 (N_30854,N_29282,N_28448);
nor U30855 (N_30855,N_29817,N_28433);
xnor U30856 (N_30856,N_28513,N_28734);
or U30857 (N_30857,N_28817,N_28144);
xor U30858 (N_30858,N_29844,N_28274);
and U30859 (N_30859,N_29022,N_29633);
and U30860 (N_30860,N_29929,N_29853);
and U30861 (N_30861,N_29211,N_28662);
and U30862 (N_30862,N_28348,N_29441);
or U30863 (N_30863,N_28446,N_29576);
or U30864 (N_30864,N_28564,N_28334);
and U30865 (N_30865,N_29672,N_28054);
xnor U30866 (N_30866,N_29941,N_28102);
or U30867 (N_30867,N_28175,N_29248);
and U30868 (N_30868,N_28410,N_28621);
and U30869 (N_30869,N_29491,N_29402);
and U30870 (N_30870,N_29151,N_29960);
nor U30871 (N_30871,N_29396,N_29172);
nand U30872 (N_30872,N_29614,N_29984);
or U30873 (N_30873,N_29035,N_29002);
nand U30874 (N_30874,N_29174,N_29660);
nor U30875 (N_30875,N_28469,N_29986);
and U30876 (N_30876,N_29884,N_29296);
and U30877 (N_30877,N_29235,N_28355);
xor U30878 (N_30878,N_28118,N_28603);
nor U30879 (N_30879,N_28743,N_29023);
nand U30880 (N_30880,N_29916,N_28966);
nor U30881 (N_30881,N_28022,N_29834);
xor U30882 (N_30882,N_28826,N_28341);
and U30883 (N_30883,N_29618,N_29256);
or U30884 (N_30884,N_29804,N_29374);
or U30885 (N_30885,N_28836,N_28210);
nor U30886 (N_30886,N_29493,N_28186);
or U30887 (N_30887,N_28808,N_28401);
xnor U30888 (N_30888,N_29835,N_28697);
xor U30889 (N_30889,N_28756,N_28394);
nor U30890 (N_30890,N_28027,N_29334);
or U30891 (N_30891,N_29280,N_29656);
xor U30892 (N_30892,N_29806,N_28922);
xnor U30893 (N_30893,N_28583,N_29314);
nand U30894 (N_30894,N_28297,N_29543);
nand U30895 (N_30895,N_28923,N_29433);
nor U30896 (N_30896,N_28335,N_28035);
or U30897 (N_30897,N_29957,N_28553);
nand U30898 (N_30898,N_28829,N_29093);
and U30899 (N_30899,N_28739,N_29726);
or U30900 (N_30900,N_29978,N_29457);
and U30901 (N_30901,N_28380,N_29405);
and U30902 (N_30902,N_28541,N_28178);
nor U30903 (N_30903,N_28337,N_28479);
and U30904 (N_30904,N_29466,N_28916);
and U30905 (N_30905,N_28967,N_28276);
or U30906 (N_30906,N_29218,N_29517);
or U30907 (N_30907,N_28624,N_29219);
xor U30908 (N_30908,N_28878,N_29579);
and U30909 (N_30909,N_28045,N_29237);
or U30910 (N_30910,N_29649,N_28638);
and U30911 (N_30911,N_29042,N_29851);
nand U30912 (N_30912,N_28190,N_28879);
or U30913 (N_30913,N_28431,N_29178);
or U30914 (N_30914,N_29246,N_28289);
and U30915 (N_30915,N_29631,N_28456);
xnor U30916 (N_30916,N_28657,N_29512);
nor U30917 (N_30917,N_28270,N_29845);
nand U30918 (N_30918,N_28750,N_28424);
or U30919 (N_30919,N_29741,N_29080);
or U30920 (N_30920,N_29158,N_29227);
or U30921 (N_30921,N_28224,N_28606);
nor U30922 (N_30922,N_29057,N_28391);
nand U30923 (N_30923,N_29939,N_28675);
or U30924 (N_30924,N_28445,N_28761);
nor U30925 (N_30925,N_29839,N_28504);
and U30926 (N_30926,N_28883,N_28989);
and U30927 (N_30927,N_29735,N_28203);
nor U30928 (N_30928,N_29815,N_29746);
or U30929 (N_30929,N_29351,N_29827);
nor U30930 (N_30930,N_28480,N_29619);
xnor U30931 (N_30931,N_29529,N_29474);
xnor U30932 (N_30932,N_29648,N_29146);
nor U30933 (N_30933,N_28209,N_28533);
nor U30934 (N_30934,N_29980,N_28231);
nand U30935 (N_30935,N_28534,N_29790);
nor U30936 (N_30936,N_29376,N_29275);
xnor U30937 (N_30937,N_29336,N_28411);
and U30938 (N_30938,N_29000,N_29662);
nand U30939 (N_30939,N_29938,N_28634);
xor U30940 (N_30940,N_28071,N_29343);
nand U30941 (N_30941,N_29438,N_28974);
xor U30942 (N_30942,N_28000,N_29442);
or U30943 (N_30943,N_28800,N_28074);
nor U30944 (N_30944,N_28429,N_29487);
nor U30945 (N_30945,N_28919,N_29030);
and U30946 (N_30946,N_29766,N_28312);
nand U30947 (N_30947,N_28192,N_29450);
and U30948 (N_30948,N_28566,N_29283);
and U30949 (N_30949,N_28342,N_28007);
and U30950 (N_30950,N_28932,N_29574);
xor U30951 (N_30951,N_28455,N_29871);
nor U30952 (N_30952,N_28656,N_28930);
nor U30953 (N_30953,N_28920,N_29603);
xor U30954 (N_30954,N_28321,N_28669);
and U30955 (N_30955,N_29807,N_28232);
nand U30956 (N_30956,N_28249,N_28048);
and U30957 (N_30957,N_29883,N_29482);
nand U30958 (N_30958,N_28647,N_29094);
or U30959 (N_30959,N_29245,N_28857);
nand U30960 (N_30960,N_29496,N_28291);
nand U30961 (N_30961,N_29062,N_28123);
xor U30962 (N_30962,N_29399,N_29216);
or U30963 (N_30963,N_29785,N_28330);
and U30964 (N_30964,N_28025,N_29787);
nor U30965 (N_30965,N_28309,N_28278);
nor U30966 (N_30966,N_29407,N_29083);
and U30967 (N_30967,N_29607,N_28427);
or U30968 (N_30968,N_29810,N_29745);
nor U30969 (N_30969,N_28343,N_28477);
and U30970 (N_30970,N_29095,N_29922);
nand U30971 (N_30971,N_28804,N_29909);
nor U30972 (N_30972,N_28327,N_29352);
nand U30973 (N_30973,N_29233,N_28516);
xnor U30974 (N_30974,N_29558,N_29664);
and U30975 (N_30975,N_28681,N_28497);
and U30976 (N_30976,N_29230,N_28218);
and U30977 (N_30977,N_29948,N_29338);
xor U30978 (N_30978,N_29112,N_28481);
nand U30979 (N_30979,N_28790,N_29549);
xor U30980 (N_30980,N_28412,N_29893);
nor U30981 (N_30981,N_28440,N_29436);
or U30982 (N_30982,N_28778,N_29372);
nor U30983 (N_30983,N_29044,N_28393);
nand U30984 (N_30984,N_29332,N_28166);
nor U30985 (N_30985,N_29640,N_28735);
nor U30986 (N_30986,N_28137,N_28854);
or U30987 (N_30987,N_28351,N_29264);
xor U30988 (N_30988,N_29933,N_28450);
and U30989 (N_30989,N_28033,N_28664);
xnor U30990 (N_30990,N_28557,N_29751);
nor U30991 (N_30991,N_28964,N_28592);
and U30992 (N_30992,N_28574,N_28037);
nand U30993 (N_30993,N_29359,N_28730);
or U30994 (N_30994,N_29229,N_29991);
or U30995 (N_30995,N_29367,N_28945);
or U30996 (N_30996,N_28111,N_28509);
nor U30997 (N_30997,N_28626,N_29404);
nand U30998 (N_30998,N_28314,N_29843);
nand U30999 (N_30999,N_29257,N_29765);
nand U31000 (N_31000,N_28602,N_28586);
nand U31001 (N_31001,N_29778,N_28209);
xnor U31002 (N_31002,N_28380,N_28619);
nand U31003 (N_31003,N_28784,N_28322);
and U31004 (N_31004,N_28845,N_29697);
xor U31005 (N_31005,N_29034,N_29811);
and U31006 (N_31006,N_29501,N_29146);
or U31007 (N_31007,N_28808,N_28122);
and U31008 (N_31008,N_28397,N_28269);
and U31009 (N_31009,N_29108,N_28918);
and U31010 (N_31010,N_28365,N_29274);
xnor U31011 (N_31011,N_29411,N_29582);
and U31012 (N_31012,N_28155,N_28831);
xor U31013 (N_31013,N_29615,N_29854);
xor U31014 (N_31014,N_29780,N_28850);
nand U31015 (N_31015,N_28634,N_28258);
xor U31016 (N_31016,N_29923,N_29223);
xnor U31017 (N_31017,N_28323,N_28788);
nor U31018 (N_31018,N_28683,N_28487);
and U31019 (N_31019,N_29092,N_28563);
nand U31020 (N_31020,N_28177,N_28550);
and U31021 (N_31021,N_28528,N_28155);
and U31022 (N_31022,N_29180,N_29416);
nand U31023 (N_31023,N_29863,N_29202);
and U31024 (N_31024,N_28555,N_28190);
or U31025 (N_31025,N_28610,N_29733);
and U31026 (N_31026,N_29991,N_28150);
and U31027 (N_31027,N_28616,N_28934);
xor U31028 (N_31028,N_29613,N_28715);
nor U31029 (N_31029,N_28903,N_28099);
nand U31030 (N_31030,N_29609,N_28112);
nor U31031 (N_31031,N_29846,N_28211);
xor U31032 (N_31032,N_28137,N_28628);
and U31033 (N_31033,N_28062,N_29533);
nand U31034 (N_31034,N_29760,N_28155);
nor U31035 (N_31035,N_29518,N_29303);
xnor U31036 (N_31036,N_29131,N_29950);
nand U31037 (N_31037,N_29233,N_28215);
nand U31038 (N_31038,N_28593,N_29532);
nor U31039 (N_31039,N_29505,N_28790);
and U31040 (N_31040,N_29678,N_28172);
nand U31041 (N_31041,N_28542,N_29588);
or U31042 (N_31042,N_28653,N_29186);
or U31043 (N_31043,N_29765,N_29018);
nand U31044 (N_31044,N_29422,N_29748);
xnor U31045 (N_31045,N_29251,N_29325);
or U31046 (N_31046,N_28480,N_28459);
nand U31047 (N_31047,N_29816,N_29464);
nand U31048 (N_31048,N_28188,N_29639);
xnor U31049 (N_31049,N_28318,N_28467);
nor U31050 (N_31050,N_29431,N_29248);
nand U31051 (N_31051,N_28373,N_29816);
and U31052 (N_31052,N_29841,N_29939);
nor U31053 (N_31053,N_29692,N_29122);
and U31054 (N_31054,N_29042,N_28530);
or U31055 (N_31055,N_29934,N_29127);
nand U31056 (N_31056,N_28477,N_29318);
and U31057 (N_31057,N_29284,N_28348);
nand U31058 (N_31058,N_28641,N_28663);
or U31059 (N_31059,N_29831,N_29775);
nor U31060 (N_31060,N_29020,N_29339);
and U31061 (N_31061,N_29778,N_29694);
nand U31062 (N_31062,N_28719,N_29753);
or U31063 (N_31063,N_29239,N_28170);
nor U31064 (N_31064,N_28398,N_28744);
nand U31065 (N_31065,N_28864,N_28932);
nor U31066 (N_31066,N_29881,N_29516);
nor U31067 (N_31067,N_29448,N_28213);
or U31068 (N_31068,N_28527,N_28412);
nand U31069 (N_31069,N_29401,N_29762);
and U31070 (N_31070,N_29094,N_29290);
nor U31071 (N_31071,N_29564,N_29513);
nor U31072 (N_31072,N_29936,N_29130);
nor U31073 (N_31073,N_29545,N_28652);
nor U31074 (N_31074,N_28938,N_29994);
nand U31075 (N_31075,N_28997,N_29842);
nand U31076 (N_31076,N_28405,N_29312);
xnor U31077 (N_31077,N_29862,N_28080);
and U31078 (N_31078,N_29815,N_28200);
nor U31079 (N_31079,N_29658,N_29522);
or U31080 (N_31080,N_28381,N_28411);
and U31081 (N_31081,N_29528,N_29144);
nor U31082 (N_31082,N_29849,N_28387);
xor U31083 (N_31083,N_29972,N_28218);
nor U31084 (N_31084,N_28051,N_28372);
xor U31085 (N_31085,N_29814,N_28072);
xor U31086 (N_31086,N_28289,N_28849);
and U31087 (N_31087,N_28358,N_29899);
and U31088 (N_31088,N_29461,N_29106);
nor U31089 (N_31089,N_28934,N_28086);
xnor U31090 (N_31090,N_29774,N_29037);
nand U31091 (N_31091,N_28492,N_29790);
xnor U31092 (N_31092,N_28514,N_29665);
nand U31093 (N_31093,N_28148,N_28376);
nand U31094 (N_31094,N_29941,N_28256);
xnor U31095 (N_31095,N_29210,N_29852);
nand U31096 (N_31096,N_29012,N_28448);
and U31097 (N_31097,N_28227,N_28897);
xor U31098 (N_31098,N_29658,N_29488);
nor U31099 (N_31099,N_29628,N_28220);
or U31100 (N_31100,N_29739,N_28210);
nand U31101 (N_31101,N_29392,N_29101);
nor U31102 (N_31102,N_28160,N_29125);
nor U31103 (N_31103,N_28942,N_29307);
or U31104 (N_31104,N_29401,N_29840);
nor U31105 (N_31105,N_28239,N_28321);
and U31106 (N_31106,N_29179,N_28172);
xnor U31107 (N_31107,N_28496,N_28192);
or U31108 (N_31108,N_28250,N_28125);
nor U31109 (N_31109,N_28515,N_29556);
nand U31110 (N_31110,N_28070,N_28817);
or U31111 (N_31111,N_28158,N_28755);
nor U31112 (N_31112,N_29227,N_29656);
or U31113 (N_31113,N_29607,N_29951);
nand U31114 (N_31114,N_28743,N_29981);
xor U31115 (N_31115,N_29406,N_29321);
and U31116 (N_31116,N_29008,N_28071);
nand U31117 (N_31117,N_28112,N_28620);
or U31118 (N_31118,N_28617,N_28684);
nand U31119 (N_31119,N_29586,N_28449);
and U31120 (N_31120,N_28870,N_28352);
or U31121 (N_31121,N_28505,N_28989);
xnor U31122 (N_31122,N_28250,N_28251);
xor U31123 (N_31123,N_28340,N_28540);
xor U31124 (N_31124,N_28307,N_28921);
and U31125 (N_31125,N_28940,N_28216);
nor U31126 (N_31126,N_28324,N_29739);
or U31127 (N_31127,N_29176,N_29070);
or U31128 (N_31128,N_28371,N_28098);
nand U31129 (N_31129,N_28460,N_29865);
nor U31130 (N_31130,N_29544,N_28905);
and U31131 (N_31131,N_28095,N_28667);
nand U31132 (N_31132,N_28632,N_29424);
or U31133 (N_31133,N_29177,N_29410);
nand U31134 (N_31134,N_28123,N_29302);
nand U31135 (N_31135,N_29345,N_29916);
nand U31136 (N_31136,N_29552,N_29011);
xnor U31137 (N_31137,N_29404,N_29163);
and U31138 (N_31138,N_29300,N_28216);
nor U31139 (N_31139,N_29235,N_28074);
nand U31140 (N_31140,N_28373,N_29159);
xor U31141 (N_31141,N_29779,N_29681);
nor U31142 (N_31142,N_29225,N_29861);
nor U31143 (N_31143,N_28572,N_29203);
and U31144 (N_31144,N_28788,N_29375);
nand U31145 (N_31145,N_28740,N_28109);
or U31146 (N_31146,N_28506,N_28902);
xnor U31147 (N_31147,N_29853,N_29794);
nor U31148 (N_31148,N_29425,N_28377);
xor U31149 (N_31149,N_29860,N_28224);
and U31150 (N_31150,N_29986,N_29400);
xor U31151 (N_31151,N_28315,N_28788);
nand U31152 (N_31152,N_29390,N_29762);
nor U31153 (N_31153,N_28062,N_28635);
nor U31154 (N_31154,N_28241,N_28842);
or U31155 (N_31155,N_28469,N_28507);
xor U31156 (N_31156,N_28942,N_28527);
or U31157 (N_31157,N_29726,N_29227);
nand U31158 (N_31158,N_28291,N_29801);
nor U31159 (N_31159,N_29883,N_28857);
and U31160 (N_31160,N_28877,N_29785);
and U31161 (N_31161,N_29295,N_29619);
xor U31162 (N_31162,N_29385,N_29435);
nor U31163 (N_31163,N_29253,N_29832);
nor U31164 (N_31164,N_29394,N_29482);
or U31165 (N_31165,N_28501,N_29529);
nand U31166 (N_31166,N_28134,N_29830);
and U31167 (N_31167,N_29225,N_28480);
nor U31168 (N_31168,N_28024,N_29048);
nand U31169 (N_31169,N_28877,N_28496);
or U31170 (N_31170,N_28023,N_29345);
and U31171 (N_31171,N_29719,N_28202);
xor U31172 (N_31172,N_28556,N_29017);
or U31173 (N_31173,N_28394,N_29187);
or U31174 (N_31174,N_28964,N_28676);
xor U31175 (N_31175,N_29637,N_28039);
and U31176 (N_31176,N_28701,N_29654);
nor U31177 (N_31177,N_29229,N_28577);
xor U31178 (N_31178,N_28634,N_28980);
or U31179 (N_31179,N_28062,N_29431);
or U31180 (N_31180,N_28909,N_28060);
xnor U31181 (N_31181,N_28320,N_28419);
xnor U31182 (N_31182,N_28000,N_29134);
and U31183 (N_31183,N_28733,N_28060);
nand U31184 (N_31184,N_29694,N_28435);
xor U31185 (N_31185,N_28152,N_28082);
nand U31186 (N_31186,N_29063,N_28359);
and U31187 (N_31187,N_28082,N_28785);
nor U31188 (N_31188,N_29585,N_28206);
xnor U31189 (N_31189,N_28027,N_28079);
nand U31190 (N_31190,N_29054,N_28215);
and U31191 (N_31191,N_28513,N_29006);
nand U31192 (N_31192,N_29055,N_28584);
or U31193 (N_31193,N_29722,N_28622);
nor U31194 (N_31194,N_28560,N_29827);
or U31195 (N_31195,N_29792,N_28202);
xnor U31196 (N_31196,N_29726,N_28063);
or U31197 (N_31197,N_29034,N_29792);
or U31198 (N_31198,N_29669,N_29176);
nor U31199 (N_31199,N_28173,N_29514);
and U31200 (N_31200,N_29930,N_28326);
xnor U31201 (N_31201,N_29595,N_29254);
or U31202 (N_31202,N_28154,N_28667);
xor U31203 (N_31203,N_29865,N_29097);
xnor U31204 (N_31204,N_28265,N_28619);
xor U31205 (N_31205,N_28216,N_28948);
and U31206 (N_31206,N_28757,N_28534);
nor U31207 (N_31207,N_28824,N_29943);
nor U31208 (N_31208,N_29107,N_28308);
nand U31209 (N_31209,N_28468,N_28363);
xor U31210 (N_31210,N_29624,N_29656);
or U31211 (N_31211,N_29965,N_28457);
nand U31212 (N_31212,N_29868,N_29788);
nand U31213 (N_31213,N_29214,N_29216);
or U31214 (N_31214,N_29182,N_29647);
and U31215 (N_31215,N_29413,N_28952);
and U31216 (N_31216,N_29776,N_28969);
nand U31217 (N_31217,N_29576,N_29869);
nand U31218 (N_31218,N_28281,N_29748);
nand U31219 (N_31219,N_28380,N_28404);
xnor U31220 (N_31220,N_28959,N_28503);
nand U31221 (N_31221,N_29577,N_29827);
xnor U31222 (N_31222,N_29238,N_28304);
xnor U31223 (N_31223,N_29662,N_29583);
or U31224 (N_31224,N_28823,N_28983);
nor U31225 (N_31225,N_29345,N_29378);
and U31226 (N_31226,N_28737,N_28677);
xor U31227 (N_31227,N_28382,N_29400);
xor U31228 (N_31228,N_28657,N_29833);
nand U31229 (N_31229,N_28727,N_28967);
nand U31230 (N_31230,N_29431,N_28880);
xor U31231 (N_31231,N_28910,N_28118);
nor U31232 (N_31232,N_29894,N_29380);
and U31233 (N_31233,N_29991,N_28316);
nand U31234 (N_31234,N_28745,N_28143);
nand U31235 (N_31235,N_28317,N_29587);
nand U31236 (N_31236,N_29217,N_29109);
nor U31237 (N_31237,N_28200,N_28898);
xor U31238 (N_31238,N_28995,N_28398);
nor U31239 (N_31239,N_28965,N_28201);
or U31240 (N_31240,N_28911,N_29157);
nand U31241 (N_31241,N_28209,N_29396);
or U31242 (N_31242,N_28690,N_29088);
xor U31243 (N_31243,N_28515,N_28035);
xnor U31244 (N_31244,N_28970,N_28336);
nand U31245 (N_31245,N_29668,N_29714);
nand U31246 (N_31246,N_29739,N_28384);
nand U31247 (N_31247,N_28089,N_28805);
or U31248 (N_31248,N_28075,N_28306);
xor U31249 (N_31249,N_29396,N_28775);
and U31250 (N_31250,N_29021,N_28927);
xnor U31251 (N_31251,N_29656,N_29194);
and U31252 (N_31252,N_29724,N_29020);
and U31253 (N_31253,N_28428,N_29410);
nor U31254 (N_31254,N_28663,N_29921);
nor U31255 (N_31255,N_29592,N_28495);
or U31256 (N_31256,N_28206,N_28434);
nand U31257 (N_31257,N_28042,N_28616);
nor U31258 (N_31258,N_28795,N_28144);
and U31259 (N_31259,N_29058,N_28354);
and U31260 (N_31260,N_29831,N_28299);
xor U31261 (N_31261,N_29002,N_28793);
and U31262 (N_31262,N_28963,N_29919);
and U31263 (N_31263,N_29102,N_29311);
or U31264 (N_31264,N_29518,N_28556);
nor U31265 (N_31265,N_28209,N_29325);
or U31266 (N_31266,N_28932,N_29102);
xor U31267 (N_31267,N_29310,N_28621);
nor U31268 (N_31268,N_29002,N_29806);
xor U31269 (N_31269,N_29337,N_29380);
xnor U31270 (N_31270,N_29319,N_29256);
nand U31271 (N_31271,N_29623,N_29073);
and U31272 (N_31272,N_29138,N_29752);
or U31273 (N_31273,N_28335,N_28745);
nand U31274 (N_31274,N_29659,N_28762);
xnor U31275 (N_31275,N_28146,N_28781);
nor U31276 (N_31276,N_28370,N_29701);
nor U31277 (N_31277,N_29948,N_28406);
nor U31278 (N_31278,N_29182,N_29133);
nand U31279 (N_31279,N_28641,N_28153);
nor U31280 (N_31280,N_29897,N_29411);
nand U31281 (N_31281,N_29766,N_28529);
nor U31282 (N_31282,N_29296,N_28951);
and U31283 (N_31283,N_28071,N_29376);
xnor U31284 (N_31284,N_29694,N_29424);
xor U31285 (N_31285,N_29050,N_28183);
nand U31286 (N_31286,N_28843,N_28254);
xor U31287 (N_31287,N_29504,N_29834);
and U31288 (N_31288,N_29899,N_29524);
nor U31289 (N_31289,N_28989,N_29682);
xnor U31290 (N_31290,N_29195,N_28022);
and U31291 (N_31291,N_29537,N_29412);
nand U31292 (N_31292,N_29654,N_29274);
and U31293 (N_31293,N_28266,N_28077);
xnor U31294 (N_31294,N_28238,N_29449);
nand U31295 (N_31295,N_28273,N_29739);
nor U31296 (N_31296,N_28854,N_28882);
or U31297 (N_31297,N_29149,N_29520);
xor U31298 (N_31298,N_29871,N_28955);
or U31299 (N_31299,N_28927,N_28089);
or U31300 (N_31300,N_29884,N_29125);
or U31301 (N_31301,N_28286,N_28152);
or U31302 (N_31302,N_29500,N_28982);
nor U31303 (N_31303,N_29579,N_28593);
xnor U31304 (N_31304,N_29105,N_29682);
or U31305 (N_31305,N_29496,N_29674);
xnor U31306 (N_31306,N_28740,N_29751);
and U31307 (N_31307,N_29797,N_28072);
nor U31308 (N_31308,N_29663,N_29575);
xnor U31309 (N_31309,N_28507,N_28800);
nand U31310 (N_31310,N_28946,N_29678);
nand U31311 (N_31311,N_28369,N_28447);
nand U31312 (N_31312,N_29403,N_28849);
nand U31313 (N_31313,N_28335,N_29456);
xnor U31314 (N_31314,N_29962,N_28114);
or U31315 (N_31315,N_29192,N_28380);
xor U31316 (N_31316,N_28248,N_28090);
xor U31317 (N_31317,N_28224,N_29233);
nand U31318 (N_31318,N_29053,N_29348);
nor U31319 (N_31319,N_29375,N_28527);
nor U31320 (N_31320,N_29234,N_29944);
or U31321 (N_31321,N_28318,N_29210);
or U31322 (N_31322,N_28045,N_28042);
xor U31323 (N_31323,N_28226,N_28220);
xor U31324 (N_31324,N_29798,N_28448);
nand U31325 (N_31325,N_29474,N_28219);
and U31326 (N_31326,N_29287,N_29848);
and U31327 (N_31327,N_29773,N_29238);
or U31328 (N_31328,N_28077,N_29828);
xnor U31329 (N_31329,N_28662,N_29583);
nor U31330 (N_31330,N_29424,N_29935);
xnor U31331 (N_31331,N_28428,N_29374);
and U31332 (N_31332,N_29550,N_28759);
nor U31333 (N_31333,N_29964,N_29015);
nand U31334 (N_31334,N_29854,N_28851);
xor U31335 (N_31335,N_28033,N_28631);
nor U31336 (N_31336,N_28120,N_28619);
nor U31337 (N_31337,N_29201,N_29943);
or U31338 (N_31338,N_28927,N_28162);
nand U31339 (N_31339,N_28076,N_29470);
xnor U31340 (N_31340,N_29177,N_29760);
or U31341 (N_31341,N_28119,N_28313);
nor U31342 (N_31342,N_29262,N_28660);
nand U31343 (N_31343,N_28198,N_28818);
nand U31344 (N_31344,N_29191,N_29438);
and U31345 (N_31345,N_28923,N_29766);
nor U31346 (N_31346,N_28669,N_29783);
or U31347 (N_31347,N_28044,N_29395);
nor U31348 (N_31348,N_28076,N_28722);
nand U31349 (N_31349,N_29088,N_29520);
nand U31350 (N_31350,N_28220,N_28558);
nand U31351 (N_31351,N_29154,N_28799);
and U31352 (N_31352,N_28574,N_28016);
nor U31353 (N_31353,N_28390,N_28330);
nand U31354 (N_31354,N_28849,N_28739);
nand U31355 (N_31355,N_29700,N_28749);
nor U31356 (N_31356,N_28799,N_28432);
and U31357 (N_31357,N_29565,N_28703);
xnor U31358 (N_31358,N_29907,N_29963);
or U31359 (N_31359,N_28745,N_28782);
or U31360 (N_31360,N_29787,N_29258);
nor U31361 (N_31361,N_29202,N_28328);
xor U31362 (N_31362,N_28781,N_28455);
nand U31363 (N_31363,N_28406,N_29422);
and U31364 (N_31364,N_28070,N_29909);
or U31365 (N_31365,N_29172,N_28331);
nand U31366 (N_31366,N_29942,N_28176);
and U31367 (N_31367,N_28538,N_28396);
or U31368 (N_31368,N_29483,N_29512);
nand U31369 (N_31369,N_29859,N_28310);
or U31370 (N_31370,N_28837,N_28876);
nand U31371 (N_31371,N_28282,N_28594);
xor U31372 (N_31372,N_28002,N_29562);
xnor U31373 (N_31373,N_29400,N_28871);
nor U31374 (N_31374,N_28240,N_29501);
and U31375 (N_31375,N_29041,N_28306);
and U31376 (N_31376,N_28956,N_28858);
or U31377 (N_31377,N_28727,N_28928);
and U31378 (N_31378,N_28605,N_28978);
nor U31379 (N_31379,N_29638,N_28983);
nand U31380 (N_31380,N_29375,N_28408);
or U31381 (N_31381,N_29415,N_28000);
xor U31382 (N_31382,N_28955,N_28631);
or U31383 (N_31383,N_28674,N_29419);
xor U31384 (N_31384,N_29413,N_28205);
nand U31385 (N_31385,N_29324,N_29829);
xnor U31386 (N_31386,N_29960,N_29127);
xor U31387 (N_31387,N_28691,N_29264);
or U31388 (N_31388,N_29045,N_28001);
or U31389 (N_31389,N_28807,N_29916);
and U31390 (N_31390,N_28216,N_29767);
nor U31391 (N_31391,N_29947,N_28343);
and U31392 (N_31392,N_28736,N_29615);
or U31393 (N_31393,N_29244,N_29805);
and U31394 (N_31394,N_28592,N_29084);
nand U31395 (N_31395,N_28836,N_28024);
and U31396 (N_31396,N_29429,N_29964);
and U31397 (N_31397,N_29212,N_29467);
xor U31398 (N_31398,N_29847,N_28993);
xnor U31399 (N_31399,N_28001,N_29756);
or U31400 (N_31400,N_29660,N_29261);
xor U31401 (N_31401,N_28226,N_28422);
or U31402 (N_31402,N_28892,N_29407);
and U31403 (N_31403,N_28492,N_29353);
nor U31404 (N_31404,N_28214,N_29984);
or U31405 (N_31405,N_29011,N_28356);
nand U31406 (N_31406,N_28845,N_28220);
nand U31407 (N_31407,N_28948,N_29667);
and U31408 (N_31408,N_29621,N_29435);
nor U31409 (N_31409,N_29281,N_29844);
and U31410 (N_31410,N_28337,N_28802);
nor U31411 (N_31411,N_28861,N_29154);
or U31412 (N_31412,N_29627,N_28357);
xor U31413 (N_31413,N_29630,N_29767);
and U31414 (N_31414,N_28690,N_28916);
and U31415 (N_31415,N_28589,N_28420);
xor U31416 (N_31416,N_28433,N_28179);
or U31417 (N_31417,N_29849,N_28248);
nor U31418 (N_31418,N_29481,N_29340);
or U31419 (N_31419,N_29504,N_29210);
nand U31420 (N_31420,N_28726,N_28450);
nand U31421 (N_31421,N_28280,N_29537);
and U31422 (N_31422,N_28348,N_29733);
or U31423 (N_31423,N_28361,N_29817);
or U31424 (N_31424,N_28039,N_28552);
nor U31425 (N_31425,N_29307,N_29543);
nor U31426 (N_31426,N_28190,N_28379);
nor U31427 (N_31427,N_28007,N_28321);
nand U31428 (N_31428,N_29096,N_29350);
or U31429 (N_31429,N_29394,N_28199);
xor U31430 (N_31430,N_29112,N_29110);
nand U31431 (N_31431,N_29470,N_28349);
nand U31432 (N_31432,N_29461,N_28888);
nand U31433 (N_31433,N_29400,N_28614);
or U31434 (N_31434,N_28838,N_28411);
xnor U31435 (N_31435,N_28566,N_29648);
nor U31436 (N_31436,N_29592,N_28714);
xnor U31437 (N_31437,N_29021,N_29516);
or U31438 (N_31438,N_28405,N_29632);
nand U31439 (N_31439,N_29473,N_29585);
xor U31440 (N_31440,N_28728,N_28686);
nor U31441 (N_31441,N_28931,N_28723);
nand U31442 (N_31442,N_28614,N_28494);
nor U31443 (N_31443,N_28602,N_29009);
nor U31444 (N_31444,N_28812,N_28690);
and U31445 (N_31445,N_29100,N_29899);
xnor U31446 (N_31446,N_28834,N_28639);
or U31447 (N_31447,N_28620,N_29333);
nor U31448 (N_31448,N_29134,N_28585);
and U31449 (N_31449,N_28817,N_28686);
nor U31450 (N_31450,N_28223,N_28562);
and U31451 (N_31451,N_29177,N_29435);
and U31452 (N_31452,N_28545,N_28017);
nor U31453 (N_31453,N_28962,N_29518);
nand U31454 (N_31454,N_29311,N_28843);
nand U31455 (N_31455,N_28847,N_28384);
xnor U31456 (N_31456,N_28900,N_28585);
nor U31457 (N_31457,N_29049,N_28446);
xor U31458 (N_31458,N_28158,N_29111);
nor U31459 (N_31459,N_28598,N_29304);
and U31460 (N_31460,N_29641,N_29239);
nand U31461 (N_31461,N_29400,N_28334);
nand U31462 (N_31462,N_29376,N_28871);
nor U31463 (N_31463,N_28482,N_28645);
and U31464 (N_31464,N_28206,N_29694);
nor U31465 (N_31465,N_28228,N_28263);
and U31466 (N_31466,N_29149,N_29516);
nor U31467 (N_31467,N_28987,N_28863);
nand U31468 (N_31468,N_29773,N_29789);
xor U31469 (N_31469,N_29834,N_29909);
and U31470 (N_31470,N_29871,N_29156);
xor U31471 (N_31471,N_29210,N_28494);
xnor U31472 (N_31472,N_29509,N_28473);
or U31473 (N_31473,N_28317,N_29564);
xnor U31474 (N_31474,N_29441,N_28614);
nor U31475 (N_31475,N_28465,N_29920);
or U31476 (N_31476,N_28422,N_29165);
nand U31477 (N_31477,N_28397,N_28299);
xor U31478 (N_31478,N_28166,N_29610);
xnor U31479 (N_31479,N_28123,N_29970);
nor U31480 (N_31480,N_28724,N_28741);
nand U31481 (N_31481,N_29944,N_29974);
nand U31482 (N_31482,N_28299,N_29459);
and U31483 (N_31483,N_29692,N_29279);
and U31484 (N_31484,N_29322,N_29546);
and U31485 (N_31485,N_29572,N_28925);
or U31486 (N_31486,N_29222,N_29837);
or U31487 (N_31487,N_29942,N_28612);
xnor U31488 (N_31488,N_28812,N_29740);
or U31489 (N_31489,N_28880,N_29577);
or U31490 (N_31490,N_29636,N_28742);
nand U31491 (N_31491,N_29681,N_29997);
or U31492 (N_31492,N_28155,N_28599);
nor U31493 (N_31493,N_29558,N_28246);
and U31494 (N_31494,N_29238,N_29588);
nor U31495 (N_31495,N_29246,N_28843);
nand U31496 (N_31496,N_28915,N_28588);
and U31497 (N_31497,N_28142,N_29633);
nand U31498 (N_31498,N_28776,N_29109);
or U31499 (N_31499,N_29490,N_29885);
nor U31500 (N_31500,N_29641,N_28130);
nor U31501 (N_31501,N_29938,N_28471);
and U31502 (N_31502,N_28618,N_28479);
nor U31503 (N_31503,N_29967,N_29204);
nor U31504 (N_31504,N_29206,N_28225);
and U31505 (N_31505,N_28279,N_28446);
xor U31506 (N_31506,N_28426,N_29079);
and U31507 (N_31507,N_28358,N_28878);
xnor U31508 (N_31508,N_29488,N_29792);
or U31509 (N_31509,N_29861,N_29963);
xor U31510 (N_31510,N_28128,N_29008);
or U31511 (N_31511,N_29082,N_28967);
nor U31512 (N_31512,N_29048,N_28408);
and U31513 (N_31513,N_28207,N_29223);
nor U31514 (N_31514,N_28445,N_29577);
or U31515 (N_31515,N_29865,N_28521);
nand U31516 (N_31516,N_28852,N_28932);
and U31517 (N_31517,N_28860,N_29785);
nand U31518 (N_31518,N_28335,N_28190);
or U31519 (N_31519,N_28961,N_29157);
nand U31520 (N_31520,N_28706,N_28808);
nand U31521 (N_31521,N_28587,N_29766);
or U31522 (N_31522,N_29039,N_29820);
nand U31523 (N_31523,N_28758,N_29842);
or U31524 (N_31524,N_29340,N_28675);
nor U31525 (N_31525,N_29490,N_28883);
or U31526 (N_31526,N_28443,N_28576);
nor U31527 (N_31527,N_29834,N_29722);
nor U31528 (N_31528,N_28824,N_29811);
or U31529 (N_31529,N_29720,N_29795);
nand U31530 (N_31530,N_28770,N_29637);
xor U31531 (N_31531,N_29750,N_29385);
nand U31532 (N_31532,N_29825,N_29416);
xor U31533 (N_31533,N_28063,N_29446);
nand U31534 (N_31534,N_28955,N_28004);
and U31535 (N_31535,N_29783,N_28364);
nand U31536 (N_31536,N_29292,N_29913);
and U31537 (N_31537,N_28635,N_29836);
xor U31538 (N_31538,N_28353,N_29501);
or U31539 (N_31539,N_28185,N_28183);
nand U31540 (N_31540,N_29357,N_29339);
and U31541 (N_31541,N_28174,N_28415);
nand U31542 (N_31542,N_29052,N_28022);
xnor U31543 (N_31543,N_29259,N_29474);
nor U31544 (N_31544,N_29782,N_29034);
and U31545 (N_31545,N_28446,N_29446);
nand U31546 (N_31546,N_29075,N_28780);
xnor U31547 (N_31547,N_28480,N_28923);
nand U31548 (N_31548,N_28472,N_29517);
nand U31549 (N_31549,N_28385,N_29507);
and U31550 (N_31550,N_29279,N_28955);
nand U31551 (N_31551,N_29637,N_29463);
nor U31552 (N_31552,N_29836,N_29955);
nor U31553 (N_31553,N_29658,N_28203);
xnor U31554 (N_31554,N_29932,N_28404);
nor U31555 (N_31555,N_29806,N_29264);
and U31556 (N_31556,N_29022,N_29795);
xor U31557 (N_31557,N_28437,N_28014);
nor U31558 (N_31558,N_29748,N_29650);
or U31559 (N_31559,N_28565,N_28489);
and U31560 (N_31560,N_28729,N_28933);
or U31561 (N_31561,N_29581,N_28452);
and U31562 (N_31562,N_29546,N_29545);
xor U31563 (N_31563,N_29515,N_29440);
xor U31564 (N_31564,N_28195,N_29348);
nand U31565 (N_31565,N_29862,N_28955);
or U31566 (N_31566,N_29372,N_29954);
nand U31567 (N_31567,N_28126,N_29198);
or U31568 (N_31568,N_29398,N_29533);
nor U31569 (N_31569,N_28394,N_28808);
and U31570 (N_31570,N_28793,N_29496);
xor U31571 (N_31571,N_29973,N_28758);
or U31572 (N_31572,N_29666,N_29915);
and U31573 (N_31573,N_28030,N_29045);
nand U31574 (N_31574,N_29965,N_28645);
xor U31575 (N_31575,N_28450,N_28883);
xnor U31576 (N_31576,N_29183,N_29851);
nor U31577 (N_31577,N_29228,N_29331);
nand U31578 (N_31578,N_28666,N_29984);
nor U31579 (N_31579,N_29579,N_29926);
nand U31580 (N_31580,N_29306,N_28098);
nand U31581 (N_31581,N_28515,N_29475);
or U31582 (N_31582,N_29308,N_29172);
and U31583 (N_31583,N_29301,N_28806);
or U31584 (N_31584,N_28500,N_29687);
and U31585 (N_31585,N_28487,N_28058);
nand U31586 (N_31586,N_28150,N_29652);
or U31587 (N_31587,N_28459,N_29051);
or U31588 (N_31588,N_29371,N_28474);
nor U31589 (N_31589,N_29032,N_29784);
nor U31590 (N_31590,N_28987,N_29412);
xor U31591 (N_31591,N_28329,N_28152);
nand U31592 (N_31592,N_28475,N_29343);
and U31593 (N_31593,N_28359,N_28446);
nand U31594 (N_31594,N_28352,N_28862);
nand U31595 (N_31595,N_29733,N_28181);
or U31596 (N_31596,N_28919,N_28481);
or U31597 (N_31597,N_28168,N_29333);
nor U31598 (N_31598,N_29878,N_29545);
nand U31599 (N_31599,N_29227,N_28211);
and U31600 (N_31600,N_28163,N_29947);
xnor U31601 (N_31601,N_29165,N_29557);
or U31602 (N_31602,N_28275,N_29992);
nand U31603 (N_31603,N_28739,N_28923);
xnor U31604 (N_31604,N_28095,N_29457);
or U31605 (N_31605,N_29631,N_29964);
nand U31606 (N_31606,N_28051,N_28360);
or U31607 (N_31607,N_28339,N_28873);
and U31608 (N_31608,N_28255,N_28889);
xor U31609 (N_31609,N_28037,N_29455);
and U31610 (N_31610,N_28932,N_29031);
nand U31611 (N_31611,N_29089,N_29509);
nand U31612 (N_31612,N_28139,N_28959);
nand U31613 (N_31613,N_28431,N_28615);
and U31614 (N_31614,N_28115,N_29212);
nand U31615 (N_31615,N_29557,N_28924);
nand U31616 (N_31616,N_28495,N_29609);
xor U31617 (N_31617,N_29715,N_29360);
nand U31618 (N_31618,N_29527,N_28538);
or U31619 (N_31619,N_29342,N_28022);
xor U31620 (N_31620,N_29663,N_29011);
or U31621 (N_31621,N_29297,N_28748);
or U31622 (N_31622,N_28665,N_29275);
or U31623 (N_31623,N_29580,N_29372);
nand U31624 (N_31624,N_28400,N_29469);
or U31625 (N_31625,N_28998,N_29660);
xnor U31626 (N_31626,N_28593,N_28971);
nor U31627 (N_31627,N_29190,N_28828);
nand U31628 (N_31628,N_29166,N_28367);
nand U31629 (N_31629,N_29372,N_29870);
nor U31630 (N_31630,N_28364,N_29252);
and U31631 (N_31631,N_29838,N_28704);
nor U31632 (N_31632,N_29004,N_29508);
or U31633 (N_31633,N_29406,N_29005);
and U31634 (N_31634,N_28582,N_29920);
and U31635 (N_31635,N_28253,N_28524);
and U31636 (N_31636,N_29435,N_28540);
nand U31637 (N_31637,N_29100,N_28724);
xnor U31638 (N_31638,N_29918,N_28781);
nand U31639 (N_31639,N_28507,N_28296);
nor U31640 (N_31640,N_28408,N_29131);
nor U31641 (N_31641,N_28664,N_29098);
xnor U31642 (N_31642,N_28668,N_28421);
xor U31643 (N_31643,N_29236,N_28424);
and U31644 (N_31644,N_28329,N_29908);
nand U31645 (N_31645,N_29226,N_29572);
nor U31646 (N_31646,N_28013,N_29291);
xnor U31647 (N_31647,N_29344,N_28908);
nor U31648 (N_31648,N_29014,N_28105);
and U31649 (N_31649,N_29049,N_29946);
nand U31650 (N_31650,N_28792,N_29444);
xnor U31651 (N_31651,N_28082,N_29457);
nor U31652 (N_31652,N_29442,N_29237);
nand U31653 (N_31653,N_28496,N_29613);
and U31654 (N_31654,N_28405,N_28299);
nand U31655 (N_31655,N_28262,N_28236);
nor U31656 (N_31656,N_29647,N_28560);
nand U31657 (N_31657,N_29756,N_28566);
xor U31658 (N_31658,N_28045,N_28963);
nor U31659 (N_31659,N_29893,N_29963);
and U31660 (N_31660,N_29134,N_29692);
nor U31661 (N_31661,N_29463,N_28976);
nand U31662 (N_31662,N_28510,N_29313);
nor U31663 (N_31663,N_28570,N_29127);
or U31664 (N_31664,N_29469,N_29229);
or U31665 (N_31665,N_28275,N_29538);
nand U31666 (N_31666,N_28244,N_29592);
xor U31667 (N_31667,N_28043,N_29006);
nand U31668 (N_31668,N_28600,N_29660);
or U31669 (N_31669,N_29761,N_29754);
or U31670 (N_31670,N_28815,N_28014);
or U31671 (N_31671,N_29122,N_29076);
xnor U31672 (N_31672,N_28360,N_29941);
or U31673 (N_31673,N_28002,N_28664);
or U31674 (N_31674,N_29664,N_28745);
nand U31675 (N_31675,N_29116,N_28858);
and U31676 (N_31676,N_28220,N_29453);
nand U31677 (N_31677,N_29968,N_28716);
and U31678 (N_31678,N_29911,N_28957);
nand U31679 (N_31679,N_29850,N_29105);
nand U31680 (N_31680,N_29498,N_28995);
and U31681 (N_31681,N_29858,N_29755);
nand U31682 (N_31682,N_28212,N_28610);
nand U31683 (N_31683,N_28239,N_29278);
nand U31684 (N_31684,N_28816,N_28889);
and U31685 (N_31685,N_28287,N_29385);
or U31686 (N_31686,N_29858,N_28338);
and U31687 (N_31687,N_29356,N_29413);
nor U31688 (N_31688,N_29006,N_29739);
or U31689 (N_31689,N_29052,N_28184);
nor U31690 (N_31690,N_28243,N_29246);
nand U31691 (N_31691,N_28799,N_29455);
or U31692 (N_31692,N_29386,N_29566);
nor U31693 (N_31693,N_28628,N_29139);
or U31694 (N_31694,N_29601,N_28600);
nand U31695 (N_31695,N_29882,N_29817);
nand U31696 (N_31696,N_28161,N_28864);
nand U31697 (N_31697,N_28293,N_28880);
nand U31698 (N_31698,N_28163,N_28619);
xor U31699 (N_31699,N_28186,N_28503);
and U31700 (N_31700,N_28927,N_28246);
or U31701 (N_31701,N_28641,N_29870);
or U31702 (N_31702,N_28562,N_29573);
xnor U31703 (N_31703,N_28881,N_29489);
and U31704 (N_31704,N_29133,N_28491);
xnor U31705 (N_31705,N_28789,N_29152);
nand U31706 (N_31706,N_28680,N_28026);
nand U31707 (N_31707,N_29957,N_28625);
nand U31708 (N_31708,N_28587,N_28114);
nor U31709 (N_31709,N_28355,N_29899);
and U31710 (N_31710,N_28406,N_28132);
xnor U31711 (N_31711,N_29387,N_29036);
nand U31712 (N_31712,N_29424,N_29166);
and U31713 (N_31713,N_29462,N_29864);
nand U31714 (N_31714,N_29600,N_29593);
nand U31715 (N_31715,N_28151,N_28324);
or U31716 (N_31716,N_29417,N_28366);
or U31717 (N_31717,N_28149,N_29415);
nand U31718 (N_31718,N_28678,N_29482);
or U31719 (N_31719,N_29625,N_29742);
or U31720 (N_31720,N_29022,N_29240);
nand U31721 (N_31721,N_28811,N_29900);
and U31722 (N_31722,N_28729,N_29659);
or U31723 (N_31723,N_29635,N_29588);
xor U31724 (N_31724,N_28103,N_29604);
and U31725 (N_31725,N_29959,N_28424);
nor U31726 (N_31726,N_28455,N_28300);
or U31727 (N_31727,N_28861,N_29196);
nand U31728 (N_31728,N_28662,N_29100);
or U31729 (N_31729,N_28840,N_29734);
and U31730 (N_31730,N_28835,N_28565);
and U31731 (N_31731,N_29943,N_29358);
and U31732 (N_31732,N_28139,N_28502);
xor U31733 (N_31733,N_28097,N_28096);
xor U31734 (N_31734,N_29791,N_29184);
or U31735 (N_31735,N_29510,N_28941);
nand U31736 (N_31736,N_28459,N_29344);
nor U31737 (N_31737,N_29011,N_28850);
or U31738 (N_31738,N_29922,N_29097);
or U31739 (N_31739,N_28722,N_29966);
nand U31740 (N_31740,N_28464,N_28187);
and U31741 (N_31741,N_28026,N_28976);
nand U31742 (N_31742,N_28705,N_29518);
nor U31743 (N_31743,N_28307,N_29685);
or U31744 (N_31744,N_29068,N_28356);
xor U31745 (N_31745,N_28535,N_29486);
xor U31746 (N_31746,N_28498,N_28942);
and U31747 (N_31747,N_29672,N_29367);
xnor U31748 (N_31748,N_29061,N_28309);
nand U31749 (N_31749,N_29713,N_28827);
nand U31750 (N_31750,N_28182,N_29764);
nor U31751 (N_31751,N_29342,N_28956);
or U31752 (N_31752,N_28188,N_28714);
xor U31753 (N_31753,N_28768,N_28995);
or U31754 (N_31754,N_28853,N_29575);
and U31755 (N_31755,N_29798,N_28432);
nand U31756 (N_31756,N_28131,N_28558);
nor U31757 (N_31757,N_29126,N_29889);
xor U31758 (N_31758,N_28059,N_28719);
or U31759 (N_31759,N_29877,N_29801);
and U31760 (N_31760,N_29251,N_28217);
nor U31761 (N_31761,N_29616,N_29340);
or U31762 (N_31762,N_28684,N_28672);
or U31763 (N_31763,N_29632,N_29945);
xnor U31764 (N_31764,N_28313,N_28924);
nor U31765 (N_31765,N_29271,N_29817);
nor U31766 (N_31766,N_28923,N_28016);
and U31767 (N_31767,N_28107,N_29131);
xnor U31768 (N_31768,N_28553,N_28937);
and U31769 (N_31769,N_29789,N_28961);
or U31770 (N_31770,N_28092,N_29564);
or U31771 (N_31771,N_28521,N_29046);
and U31772 (N_31772,N_29335,N_28067);
and U31773 (N_31773,N_29810,N_29500);
nor U31774 (N_31774,N_28493,N_29906);
xnor U31775 (N_31775,N_28139,N_29702);
xnor U31776 (N_31776,N_28304,N_28912);
nand U31777 (N_31777,N_29157,N_28031);
xor U31778 (N_31778,N_28949,N_28296);
or U31779 (N_31779,N_29426,N_29369);
and U31780 (N_31780,N_28271,N_28197);
nand U31781 (N_31781,N_29865,N_29034);
nor U31782 (N_31782,N_29783,N_28610);
nor U31783 (N_31783,N_29268,N_28190);
nand U31784 (N_31784,N_28115,N_28065);
and U31785 (N_31785,N_28919,N_28908);
nor U31786 (N_31786,N_28696,N_29980);
nand U31787 (N_31787,N_28204,N_28465);
nand U31788 (N_31788,N_28278,N_28793);
or U31789 (N_31789,N_28236,N_28283);
xor U31790 (N_31790,N_29332,N_28185);
xnor U31791 (N_31791,N_29378,N_29452);
or U31792 (N_31792,N_29828,N_29770);
nor U31793 (N_31793,N_29795,N_28516);
nor U31794 (N_31794,N_29637,N_29544);
xnor U31795 (N_31795,N_28647,N_28390);
or U31796 (N_31796,N_28505,N_29871);
xnor U31797 (N_31797,N_29323,N_28675);
or U31798 (N_31798,N_29121,N_28608);
xnor U31799 (N_31799,N_28645,N_29539);
or U31800 (N_31800,N_29779,N_29575);
and U31801 (N_31801,N_29965,N_28720);
nand U31802 (N_31802,N_29804,N_29781);
xnor U31803 (N_31803,N_29531,N_29940);
and U31804 (N_31804,N_28237,N_29313);
nand U31805 (N_31805,N_29873,N_29076);
and U31806 (N_31806,N_28603,N_29590);
nor U31807 (N_31807,N_29271,N_29640);
nor U31808 (N_31808,N_28148,N_29589);
nand U31809 (N_31809,N_29806,N_29847);
xor U31810 (N_31810,N_28530,N_28124);
xnor U31811 (N_31811,N_29800,N_29094);
and U31812 (N_31812,N_29741,N_28217);
or U31813 (N_31813,N_29060,N_28549);
nand U31814 (N_31814,N_28032,N_29057);
and U31815 (N_31815,N_28802,N_29906);
and U31816 (N_31816,N_28257,N_29632);
nor U31817 (N_31817,N_28938,N_28041);
nand U31818 (N_31818,N_29129,N_28318);
xnor U31819 (N_31819,N_28339,N_28140);
or U31820 (N_31820,N_28188,N_29121);
or U31821 (N_31821,N_29655,N_28126);
xnor U31822 (N_31822,N_29442,N_29695);
or U31823 (N_31823,N_28915,N_29650);
nor U31824 (N_31824,N_29596,N_29738);
xor U31825 (N_31825,N_28771,N_28001);
nand U31826 (N_31826,N_28345,N_29697);
nand U31827 (N_31827,N_28786,N_29752);
or U31828 (N_31828,N_28065,N_28459);
nand U31829 (N_31829,N_29860,N_28122);
and U31830 (N_31830,N_28782,N_28063);
nor U31831 (N_31831,N_28505,N_29499);
or U31832 (N_31832,N_29746,N_29073);
xnor U31833 (N_31833,N_28085,N_29301);
or U31834 (N_31834,N_29697,N_28969);
xnor U31835 (N_31835,N_29771,N_28097);
or U31836 (N_31836,N_28550,N_29739);
or U31837 (N_31837,N_29486,N_29054);
xor U31838 (N_31838,N_29960,N_29055);
and U31839 (N_31839,N_28072,N_29384);
and U31840 (N_31840,N_29841,N_28165);
nor U31841 (N_31841,N_28380,N_28301);
and U31842 (N_31842,N_28433,N_29185);
and U31843 (N_31843,N_29844,N_29862);
and U31844 (N_31844,N_28667,N_28512);
and U31845 (N_31845,N_28691,N_29856);
and U31846 (N_31846,N_28850,N_29622);
nor U31847 (N_31847,N_28843,N_29048);
xnor U31848 (N_31848,N_28696,N_29236);
nand U31849 (N_31849,N_28406,N_28146);
or U31850 (N_31850,N_29691,N_28014);
nor U31851 (N_31851,N_28942,N_28444);
nor U31852 (N_31852,N_28815,N_29947);
xnor U31853 (N_31853,N_29358,N_29065);
or U31854 (N_31854,N_28885,N_28340);
and U31855 (N_31855,N_29161,N_28414);
nor U31856 (N_31856,N_29639,N_29880);
and U31857 (N_31857,N_29618,N_29243);
xnor U31858 (N_31858,N_28096,N_29594);
xor U31859 (N_31859,N_28696,N_28404);
and U31860 (N_31860,N_29918,N_28762);
nand U31861 (N_31861,N_28674,N_29677);
xnor U31862 (N_31862,N_29420,N_29950);
and U31863 (N_31863,N_29833,N_28007);
nor U31864 (N_31864,N_28848,N_28252);
or U31865 (N_31865,N_28399,N_29611);
or U31866 (N_31866,N_28657,N_28010);
nand U31867 (N_31867,N_28394,N_29127);
xor U31868 (N_31868,N_28276,N_28227);
or U31869 (N_31869,N_29584,N_29842);
nor U31870 (N_31870,N_29781,N_29425);
or U31871 (N_31871,N_29010,N_29202);
nor U31872 (N_31872,N_29889,N_28913);
nand U31873 (N_31873,N_28013,N_29038);
and U31874 (N_31874,N_29372,N_29516);
xor U31875 (N_31875,N_29821,N_28435);
nand U31876 (N_31876,N_29113,N_28467);
nor U31877 (N_31877,N_28315,N_29746);
or U31878 (N_31878,N_28415,N_28348);
nand U31879 (N_31879,N_29043,N_29247);
xor U31880 (N_31880,N_29785,N_29853);
xnor U31881 (N_31881,N_28933,N_29243);
and U31882 (N_31882,N_28889,N_29791);
xor U31883 (N_31883,N_29141,N_29358);
nand U31884 (N_31884,N_29745,N_28050);
xnor U31885 (N_31885,N_28786,N_28109);
and U31886 (N_31886,N_28981,N_29022);
xor U31887 (N_31887,N_28824,N_28021);
nor U31888 (N_31888,N_28388,N_28471);
nor U31889 (N_31889,N_29861,N_29471);
or U31890 (N_31890,N_29684,N_29744);
xnor U31891 (N_31891,N_29915,N_29898);
nor U31892 (N_31892,N_28702,N_28169);
and U31893 (N_31893,N_29556,N_28384);
or U31894 (N_31894,N_29008,N_29398);
xor U31895 (N_31895,N_28339,N_29258);
xor U31896 (N_31896,N_28763,N_28726);
nand U31897 (N_31897,N_28061,N_28826);
and U31898 (N_31898,N_29254,N_28143);
xnor U31899 (N_31899,N_29048,N_28401);
xnor U31900 (N_31900,N_28949,N_29854);
nor U31901 (N_31901,N_28080,N_29936);
or U31902 (N_31902,N_29676,N_28743);
nor U31903 (N_31903,N_28210,N_28872);
or U31904 (N_31904,N_29398,N_28448);
nand U31905 (N_31905,N_28847,N_28947);
nand U31906 (N_31906,N_29389,N_29835);
nand U31907 (N_31907,N_29448,N_29323);
or U31908 (N_31908,N_28374,N_29100);
nand U31909 (N_31909,N_28311,N_29494);
xor U31910 (N_31910,N_28966,N_29098);
or U31911 (N_31911,N_29568,N_28955);
nand U31912 (N_31912,N_29914,N_28743);
nor U31913 (N_31913,N_29639,N_29106);
and U31914 (N_31914,N_28939,N_28506);
and U31915 (N_31915,N_29446,N_28681);
and U31916 (N_31916,N_29140,N_28512);
xnor U31917 (N_31917,N_28255,N_29953);
nor U31918 (N_31918,N_29457,N_29148);
nor U31919 (N_31919,N_28199,N_28794);
nor U31920 (N_31920,N_29230,N_28656);
nor U31921 (N_31921,N_29549,N_28174);
or U31922 (N_31922,N_28161,N_29290);
or U31923 (N_31923,N_28127,N_28879);
and U31924 (N_31924,N_29590,N_28348);
and U31925 (N_31925,N_29752,N_29232);
nor U31926 (N_31926,N_29017,N_29783);
nand U31927 (N_31927,N_29956,N_29136);
nand U31928 (N_31928,N_28750,N_29538);
or U31929 (N_31929,N_29467,N_28954);
and U31930 (N_31930,N_29744,N_28951);
and U31931 (N_31931,N_28052,N_29495);
and U31932 (N_31932,N_28045,N_29718);
nor U31933 (N_31933,N_28346,N_28349);
and U31934 (N_31934,N_28846,N_29001);
nand U31935 (N_31935,N_29775,N_29397);
nand U31936 (N_31936,N_29414,N_28438);
xor U31937 (N_31937,N_29547,N_29738);
and U31938 (N_31938,N_29940,N_28400);
nand U31939 (N_31939,N_29311,N_29186);
xnor U31940 (N_31940,N_29861,N_28307);
nand U31941 (N_31941,N_28428,N_29324);
nor U31942 (N_31942,N_28411,N_29933);
or U31943 (N_31943,N_29361,N_28140);
and U31944 (N_31944,N_28227,N_28196);
or U31945 (N_31945,N_28159,N_28518);
or U31946 (N_31946,N_28476,N_29057);
xnor U31947 (N_31947,N_29662,N_29240);
and U31948 (N_31948,N_28748,N_29616);
nor U31949 (N_31949,N_29116,N_29322);
or U31950 (N_31950,N_29502,N_29882);
and U31951 (N_31951,N_28686,N_28754);
xnor U31952 (N_31952,N_29131,N_28385);
and U31953 (N_31953,N_29618,N_29649);
xor U31954 (N_31954,N_29507,N_28641);
xnor U31955 (N_31955,N_29710,N_29860);
nor U31956 (N_31956,N_29504,N_29724);
or U31957 (N_31957,N_28843,N_29552);
or U31958 (N_31958,N_29883,N_28847);
nor U31959 (N_31959,N_28216,N_28337);
nor U31960 (N_31960,N_28823,N_28490);
xor U31961 (N_31961,N_28577,N_29971);
or U31962 (N_31962,N_28860,N_29493);
xor U31963 (N_31963,N_28728,N_28351);
nor U31964 (N_31964,N_29390,N_28046);
and U31965 (N_31965,N_28113,N_28417);
or U31966 (N_31966,N_29887,N_28996);
nand U31967 (N_31967,N_29995,N_28723);
and U31968 (N_31968,N_28395,N_28886);
nor U31969 (N_31969,N_29353,N_28617);
nor U31970 (N_31970,N_28482,N_28024);
nand U31971 (N_31971,N_29533,N_28260);
nor U31972 (N_31972,N_29983,N_28732);
nor U31973 (N_31973,N_29050,N_28815);
and U31974 (N_31974,N_29217,N_29548);
or U31975 (N_31975,N_28586,N_28640);
nor U31976 (N_31976,N_28497,N_29833);
nor U31977 (N_31977,N_29023,N_29234);
xor U31978 (N_31978,N_28753,N_29925);
and U31979 (N_31979,N_29108,N_29963);
nand U31980 (N_31980,N_29830,N_29978);
and U31981 (N_31981,N_29888,N_28073);
nor U31982 (N_31982,N_29591,N_29814);
and U31983 (N_31983,N_29576,N_28325);
nor U31984 (N_31984,N_28256,N_29505);
nor U31985 (N_31985,N_28940,N_28436);
nor U31986 (N_31986,N_29742,N_29687);
and U31987 (N_31987,N_29506,N_28361);
xor U31988 (N_31988,N_28491,N_29069);
nor U31989 (N_31989,N_28218,N_29073);
xnor U31990 (N_31990,N_28508,N_29396);
or U31991 (N_31991,N_29698,N_29713);
or U31992 (N_31992,N_28604,N_28827);
or U31993 (N_31993,N_29708,N_29029);
nand U31994 (N_31994,N_28809,N_29384);
or U31995 (N_31995,N_28743,N_28037);
nand U31996 (N_31996,N_29080,N_29687);
xnor U31997 (N_31997,N_29057,N_28803);
nand U31998 (N_31998,N_29410,N_29387);
xnor U31999 (N_31999,N_29150,N_28215);
xnor U32000 (N_32000,N_30762,N_31113);
or U32001 (N_32001,N_31541,N_31462);
xor U32002 (N_32002,N_31271,N_31539);
nor U32003 (N_32003,N_30434,N_31686);
nor U32004 (N_32004,N_30440,N_30379);
nand U32005 (N_32005,N_31122,N_30668);
nand U32006 (N_32006,N_31579,N_31146);
or U32007 (N_32007,N_31816,N_30036);
or U32008 (N_32008,N_30248,N_30627);
or U32009 (N_32009,N_31612,N_31235);
or U32010 (N_32010,N_31528,N_31529);
xnor U32011 (N_32011,N_31034,N_30702);
nand U32012 (N_32012,N_31542,N_30323);
and U32013 (N_32013,N_30209,N_31414);
nand U32014 (N_32014,N_31388,N_30163);
xnor U32015 (N_32015,N_31015,N_31915);
nor U32016 (N_32016,N_30557,N_31137);
nand U32017 (N_32017,N_30381,N_30609);
and U32018 (N_32018,N_31105,N_31030);
or U32019 (N_32019,N_31057,N_30608);
xnor U32020 (N_32020,N_31565,N_30808);
or U32021 (N_32021,N_31705,N_30833);
xor U32022 (N_32022,N_31951,N_31992);
or U32023 (N_32023,N_31071,N_30563);
and U32024 (N_32024,N_31058,N_30536);
nand U32025 (N_32025,N_31925,N_31805);
or U32026 (N_32026,N_30122,N_30394);
or U32027 (N_32027,N_30449,N_30859);
xor U32028 (N_32028,N_31238,N_30635);
xor U32029 (N_32029,N_31524,N_31593);
xnor U32030 (N_32030,N_31179,N_30652);
nand U32031 (N_32031,N_30111,N_31794);
xnor U32032 (N_32032,N_31732,N_30550);
nand U32033 (N_32033,N_31580,N_30099);
and U32034 (N_32034,N_31830,N_30500);
and U32035 (N_32035,N_31770,N_30614);
or U32036 (N_32036,N_30512,N_30301);
nor U32037 (N_32037,N_30357,N_31525);
nor U32038 (N_32038,N_30213,N_30519);
nand U32039 (N_32039,N_31468,N_30399);
nand U32040 (N_32040,N_31018,N_31671);
nand U32041 (N_32041,N_31980,N_31772);
nor U32042 (N_32042,N_30530,N_31591);
nor U32043 (N_32043,N_30998,N_30840);
nor U32044 (N_32044,N_31265,N_30777);
or U32045 (N_32045,N_31160,N_31002);
nand U32046 (N_32046,N_31777,N_31526);
and U32047 (N_32047,N_30715,N_30282);
nor U32048 (N_32048,N_31647,N_31241);
and U32049 (N_32049,N_30793,N_31014);
and U32050 (N_32050,N_31287,N_30830);
nand U32051 (N_32051,N_30191,N_30130);
nand U32052 (N_32052,N_31262,N_31740);
xnor U32053 (N_32053,N_31130,N_30802);
nand U32054 (N_32054,N_30790,N_30135);
xor U32055 (N_32055,N_30052,N_31635);
and U32056 (N_32056,N_30771,N_30789);
nand U32057 (N_32057,N_30606,N_30258);
nor U32058 (N_32058,N_30095,N_31413);
xor U32059 (N_32059,N_31050,N_31890);
nand U32060 (N_32060,N_30016,N_31838);
xnor U32061 (N_32061,N_30646,N_30181);
or U32062 (N_32062,N_31810,N_30089);
nor U32063 (N_32063,N_31346,N_31126);
nand U32064 (N_32064,N_30716,N_31898);
and U32065 (N_32065,N_31857,N_31702);
nand U32066 (N_32066,N_30815,N_31943);
and U32067 (N_32067,N_30478,N_30272);
xor U32068 (N_32068,N_30516,N_30733);
nor U32069 (N_32069,N_30107,N_30642);
or U32070 (N_32070,N_30082,N_30719);
xnor U32071 (N_32071,N_31494,N_31520);
nand U32072 (N_32072,N_31102,N_30755);
or U32073 (N_32073,N_31266,N_30780);
xnor U32074 (N_32074,N_30205,N_30404);
nand U32075 (N_32075,N_31005,N_31922);
xnor U32076 (N_32076,N_31036,N_31779);
and U32077 (N_32077,N_31535,N_30470);
and U32078 (N_32078,N_31751,N_31895);
and U32079 (N_32079,N_30377,N_30703);
nor U32080 (N_32080,N_31795,N_31444);
or U32081 (N_32081,N_30875,N_30838);
and U32082 (N_32082,N_30065,N_30187);
xor U32083 (N_32083,N_30267,N_30832);
xor U32084 (N_32084,N_30523,N_31854);
or U32085 (N_32085,N_30074,N_30141);
nor U32086 (N_32086,N_30583,N_30904);
nor U32087 (N_32087,N_30931,N_31905);
or U32088 (N_32088,N_30582,N_30821);
or U32089 (N_32089,N_30162,N_30012);
nand U32090 (N_32090,N_31493,N_30649);
and U32091 (N_32091,N_31856,N_30910);
and U32092 (N_32092,N_31203,N_31634);
and U32093 (N_32093,N_30237,N_31744);
nor U32094 (N_32094,N_30189,N_30499);
or U32095 (N_32095,N_31986,N_31885);
nor U32096 (N_32096,N_31433,N_31750);
xnor U32097 (N_32097,N_30343,N_30843);
and U32098 (N_32098,N_31068,N_31588);
nor U32099 (N_32099,N_31787,N_31887);
or U32100 (N_32100,N_31465,N_31572);
and U32101 (N_32101,N_31739,N_31631);
nor U32102 (N_32102,N_30678,N_31923);
and U32103 (N_32103,N_30996,N_31935);
or U32104 (N_32104,N_30353,N_30728);
or U32105 (N_32105,N_30326,N_30988);
nor U32106 (N_32106,N_31073,N_30510);
nand U32107 (N_32107,N_30014,N_31913);
or U32108 (N_32108,N_31008,N_31448);
nor U32109 (N_32109,N_31255,N_30552);
nand U32110 (N_32110,N_31275,N_31282);
nor U32111 (N_32111,N_30225,N_31332);
nand U32112 (N_32112,N_30730,N_31485);
and U32113 (N_32113,N_30167,N_30750);
xor U32114 (N_32114,N_31150,N_31630);
xor U32115 (N_32115,N_30503,N_30332);
or U32116 (N_32116,N_30286,N_31285);
nand U32117 (N_32117,N_30134,N_31278);
or U32118 (N_32118,N_30775,N_30660);
and U32119 (N_32119,N_30787,N_30897);
or U32120 (N_32120,N_30373,N_30081);
nand U32121 (N_32121,N_31755,N_30410);
or U32122 (N_32122,N_31984,N_30615);
and U32123 (N_32123,N_30058,N_30864);
nor U32124 (N_32124,N_31428,N_31180);
nor U32125 (N_32125,N_31411,N_31067);
or U32126 (N_32126,N_31820,N_31140);
nand U32127 (N_32127,N_31501,N_30484);
xor U32128 (N_32128,N_30927,N_30232);
nor U32129 (N_32129,N_31195,N_30817);
nand U32130 (N_32130,N_31649,N_31283);
and U32131 (N_32131,N_30898,N_30492);
and U32132 (N_32132,N_31691,N_30184);
or U32133 (N_32133,N_31403,N_31615);
and U32134 (N_32134,N_30212,N_30648);
xnor U32135 (N_32135,N_31892,N_30480);
nand U32136 (N_32136,N_31682,N_30667);
and U32137 (N_32137,N_30863,N_30024);
nand U32138 (N_32138,N_31679,N_31025);
nand U32139 (N_32139,N_31111,N_30294);
and U32140 (N_32140,N_30241,N_30391);
or U32141 (N_32141,N_31599,N_30401);
and U32142 (N_32142,N_30390,N_30069);
nor U32143 (N_32143,N_30372,N_31741);
nor U32144 (N_32144,N_30238,N_31270);
nor U32145 (N_32145,N_31496,N_30255);
and U32146 (N_32146,N_31851,N_31076);
xnor U32147 (N_32147,N_30318,N_30654);
and U32148 (N_32148,N_31037,N_30361);
nand U32149 (N_32149,N_31582,N_30786);
nand U32150 (N_32150,N_30240,N_31212);
nor U32151 (N_32151,N_31985,N_30302);
or U32152 (N_32152,N_31832,N_31746);
nor U32153 (N_32153,N_30370,N_31688);
nand U32154 (N_32154,N_31417,N_30091);
xor U32155 (N_32155,N_31666,N_31609);
xnor U32156 (N_32156,N_31543,N_31365);
or U32157 (N_32157,N_31446,N_31439);
and U32158 (N_32158,N_30713,N_30375);
nand U32159 (N_32159,N_30042,N_30188);
nor U32160 (N_32160,N_30131,N_30059);
and U32161 (N_32161,N_30978,N_30531);
nor U32162 (N_32162,N_30247,N_30958);
nand U32163 (N_32163,N_30949,N_30482);
or U32164 (N_32164,N_30269,N_31979);
nor U32165 (N_32165,N_31155,N_30414);
xor U32166 (N_32166,N_30108,N_30767);
or U32167 (N_32167,N_30013,N_31564);
nor U32168 (N_32168,N_31627,N_30868);
nand U32169 (N_32169,N_30115,N_31606);
and U32170 (N_32170,N_30026,N_31771);
nor U32171 (N_32171,N_30179,N_30537);
nand U32172 (N_32172,N_30270,N_31198);
xor U32173 (N_32173,N_30335,N_31152);
nor U32174 (N_32174,N_30588,N_30097);
and U32175 (N_32175,N_31689,N_30558);
and U32176 (N_32176,N_30275,N_30201);
and U32177 (N_32177,N_31127,N_31183);
nand U32178 (N_32178,N_31167,N_31614);
or U32179 (N_32179,N_30788,N_30710);
nor U32180 (N_32180,N_31483,N_30756);
nor U32181 (N_32181,N_31380,N_31874);
xnor U32182 (N_32182,N_31466,N_31884);
nand U32183 (N_32183,N_30545,N_30214);
xor U32184 (N_32184,N_31157,N_31960);
and U32185 (N_32185,N_31131,N_31250);
nand U32186 (N_32186,N_30643,N_31983);
nor U32187 (N_32187,N_30930,N_31763);
xnor U32188 (N_32188,N_31205,N_31547);
or U32189 (N_32189,N_31228,N_31027);
nand U32190 (N_32190,N_30529,N_30576);
nor U32191 (N_32191,N_31638,N_30975);
and U32192 (N_32192,N_30109,N_31334);
xor U32193 (N_32193,N_30010,N_30995);
or U32194 (N_32194,N_30842,N_31502);
or U32195 (N_32195,N_31648,N_30705);
xnor U32196 (N_32196,N_30421,N_30436);
xor U32197 (N_32197,N_31882,N_30636);
or U32198 (N_32198,N_31031,N_30057);
xnor U32199 (N_32199,N_30561,N_31029);
nor U32200 (N_32200,N_31385,N_30204);
xor U32201 (N_32201,N_31181,N_31191);
or U32202 (N_32202,N_31350,N_31611);
and U32203 (N_32203,N_31459,N_31928);
and U32204 (N_32204,N_30553,N_30701);
and U32205 (N_32205,N_30444,N_30378);
nor U32206 (N_32206,N_31419,N_31909);
nor U32207 (N_32207,N_31296,N_31507);
nor U32208 (N_32208,N_30025,N_30689);
and U32209 (N_32209,N_31092,N_31693);
or U32210 (N_32210,N_30246,N_30918);
and U32211 (N_32211,N_31303,N_30175);
nor U32212 (N_32212,N_30806,N_31783);
or U32213 (N_32213,N_31032,N_30967);
nor U32214 (N_32214,N_31924,N_30263);
and U32215 (N_32215,N_30491,N_30535);
xnor U32216 (N_32216,N_30943,N_30465);
nor U32217 (N_32217,N_30330,N_31775);
and U32218 (N_32218,N_30945,N_31473);
xor U32219 (N_32219,N_30822,N_31197);
or U32220 (N_32220,N_31328,N_30916);
or U32221 (N_32221,N_31964,N_31982);
nand U32222 (N_32222,N_31490,N_30971);
and U32223 (N_32223,N_30083,N_31355);
and U32224 (N_32224,N_30319,N_31194);
and U32225 (N_32225,N_31840,N_31013);
or U32226 (N_32226,N_31276,N_31721);
and U32227 (N_32227,N_30849,N_31584);
nand U32228 (N_32228,N_31121,N_30461);
and U32229 (N_32229,N_30517,N_31399);
xnor U32230 (N_32230,N_31880,N_30070);
xnor U32231 (N_32231,N_31289,N_30487);
xnor U32232 (N_32232,N_31053,N_31696);
xnor U32233 (N_32233,N_31281,N_30939);
xnor U32234 (N_32234,N_30565,N_31240);
and U32235 (N_32235,N_30656,N_31607);
or U32236 (N_32236,N_30028,N_31597);
and U32237 (N_32237,N_30984,N_31400);
xor U32238 (N_32238,N_31457,N_31463);
nand U32239 (N_32239,N_30422,N_31972);
nand U32240 (N_32240,N_30151,N_31672);
xnor U32241 (N_32241,N_30745,N_31046);
xnor U32242 (N_32242,N_30456,N_31384);
xor U32243 (N_32243,N_31142,N_31807);
xnor U32244 (N_32244,N_30546,N_31681);
and U32245 (N_32245,N_31574,N_31001);
xor U32246 (N_32246,N_31519,N_31186);
xnor U32247 (N_32247,N_31107,N_31100);
xnor U32248 (N_32248,N_31104,N_30218);
nand U32249 (N_32249,N_31453,N_31719);
nor U32250 (N_32250,N_31327,N_31475);
or U32251 (N_32251,N_30603,N_31514);
and U32252 (N_32252,N_30432,N_30305);
nor U32253 (N_32253,N_30281,N_30265);
xor U32254 (N_32254,N_30825,N_30908);
nand U32255 (N_32255,N_31349,N_30352);
xnor U32256 (N_32256,N_31782,N_30185);
and U32257 (N_32257,N_30004,N_30841);
and U32258 (N_32258,N_30653,N_31345);
nand U32259 (N_32259,N_31099,N_30862);
nand U32260 (N_32260,N_31673,N_30279);
nand U32261 (N_32261,N_31080,N_31655);
nand U32262 (N_32262,N_30088,N_31546);
xor U32263 (N_32263,N_30828,N_30591);
nand U32264 (N_32264,N_31028,N_30851);
or U32265 (N_32265,N_31523,N_31781);
nor U32266 (N_32266,N_30169,N_30569);
or U32267 (N_32267,N_31054,N_30340);
and U32268 (N_32268,N_30324,N_30779);
nor U32269 (N_32269,N_30623,N_31353);
and U32270 (N_32270,N_31602,N_30865);
nor U32271 (N_32271,N_30783,N_30625);
or U32272 (N_32272,N_31340,N_31190);
and U32273 (N_32273,N_30298,N_31391);
xor U32274 (N_32274,N_31893,N_30941);
nand U32275 (N_32275,N_31961,N_31530);
and U32276 (N_32276,N_30691,N_30549);
and U32277 (N_32277,N_30566,N_30198);
nor U32278 (N_32278,N_31188,N_30003);
nand U32279 (N_32279,N_31814,N_30222);
and U32280 (N_32280,N_30164,N_31035);
nor U32281 (N_32281,N_31094,N_31675);
xnor U32282 (N_32282,N_31762,N_30249);
nor U32283 (N_32283,N_30527,N_31511);
and U32284 (N_32284,N_30006,N_30944);
or U32285 (N_32285,N_31201,N_30980);
nand U32286 (N_32286,N_31562,N_31154);
xnor U32287 (N_32287,N_30758,N_30230);
and U32288 (N_32288,N_30658,N_30721);
or U32289 (N_32289,N_30155,N_31697);
xnor U32290 (N_32290,N_31695,N_31662);
nor U32291 (N_32291,N_30407,N_31173);
nor U32292 (N_32292,N_30384,N_31959);
or U32293 (N_32293,N_30049,N_31970);
and U32294 (N_32294,N_31026,N_31613);
and U32295 (N_32295,N_31791,N_30231);
nand U32296 (N_32296,N_31168,N_31424);
and U32297 (N_32297,N_31643,N_30873);
xor U32298 (N_32298,N_31226,N_30676);
xnor U32299 (N_32299,N_30413,N_31504);
or U32300 (N_32300,N_30562,N_31451);
or U32301 (N_32301,N_30291,N_31687);
nand U32302 (N_32302,N_30210,N_31333);
and U32303 (N_32303,N_31553,N_30419);
or U32304 (N_32304,N_31246,N_31878);
and U32305 (N_32305,N_30112,N_31088);
and U32306 (N_32306,N_30860,N_31087);
xnor U32307 (N_32307,N_30724,N_30071);
or U32308 (N_32308,N_30754,N_31585);
and U32309 (N_32309,N_31033,N_31949);
xor U32310 (N_32310,N_30680,N_30244);
or U32311 (N_32311,N_30388,N_31753);
nor U32312 (N_32312,N_30963,N_30882);
or U32313 (N_32313,N_30035,N_31728);
nor U32314 (N_32314,N_31939,N_31184);
and U32315 (N_32315,N_31512,N_30075);
and U32316 (N_32316,N_31217,N_31086);
or U32317 (N_32317,N_30472,N_30878);
or U32318 (N_32318,N_31847,N_30337);
nor U32319 (N_32319,N_31230,N_31508);
nand U32320 (N_32320,N_31633,N_30956);
xnor U32321 (N_32321,N_31442,N_30901);
and U32322 (N_32322,N_30690,N_31766);
nor U32323 (N_32323,N_30400,N_31552);
or U32324 (N_32324,N_30640,N_31128);
or U32325 (N_32325,N_31236,N_31189);
nor U32326 (N_32326,N_30855,N_31103);
and U32327 (N_32327,N_31263,N_30193);
and U32328 (N_32328,N_30120,N_30183);
or U32329 (N_32329,N_31734,N_30037);
and U32330 (N_32330,N_31848,N_31491);
nand U32331 (N_32331,N_30645,N_31125);
or U32332 (N_32332,N_30348,N_31284);
and U32333 (N_32333,N_30772,N_30338);
and U32334 (N_32334,N_31116,N_31171);
and U32335 (N_32335,N_30002,N_31849);
nand U32336 (N_32336,N_30818,N_30481);
and U32337 (N_32337,N_30458,N_31846);
nand U32338 (N_32338,N_30599,N_31706);
and U32339 (N_32339,N_31802,N_31932);
nor U32340 (N_32340,N_31354,N_30735);
and U32341 (N_32341,N_31917,N_31062);
nand U32342 (N_32342,N_31752,N_30709);
and U32343 (N_32343,N_31590,N_31224);
nor U32344 (N_32344,N_30339,N_31192);
nor U32345 (N_32345,N_31808,N_31726);
or U32346 (N_32346,N_31019,N_30890);
nor U32347 (N_32347,N_31158,N_31676);
xor U32348 (N_32348,N_30176,N_31825);
nand U32349 (N_32349,N_31024,N_31910);
xor U32350 (N_32350,N_30018,N_31845);
nand U32351 (N_32351,N_31377,N_30961);
or U32352 (N_32352,N_30250,N_30784);
nand U32353 (N_32353,N_30251,N_31784);
xnor U32354 (N_32354,N_31310,N_30826);
nand U32355 (N_32355,N_30871,N_30217);
or U32356 (N_32356,N_30239,N_31118);
xor U32357 (N_32357,N_30759,N_30125);
nor U32358 (N_32358,N_31548,N_30448);
nand U32359 (N_32359,N_30885,N_31948);
and U32360 (N_32360,N_31320,N_31498);
or U32361 (N_32361,N_30942,N_31339);
nand U32362 (N_32362,N_30768,N_30453);
nand U32363 (N_32363,N_31251,N_30128);
xnor U32364 (N_32364,N_31718,N_30438);
xnor U32365 (N_32365,N_30977,N_30664);
or U32366 (N_32366,N_30718,N_31670);
or U32367 (N_32367,N_30322,N_31084);
or U32368 (N_32368,N_31011,N_31383);
and U32369 (N_32369,N_30123,N_30328);
xnor U32370 (N_32370,N_30476,N_30396);
and U32371 (N_32371,N_30744,N_30221);
nor U32372 (N_32372,N_30398,N_30200);
nand U32373 (N_32373,N_30146,N_31622);
and U32374 (N_32374,N_30657,N_31692);
or U32375 (N_32375,N_30234,N_31534);
or U32376 (N_32376,N_30661,N_30541);
or U32377 (N_32377,N_30990,N_30397);
xor U32378 (N_32378,N_30451,N_31376);
and U32379 (N_32379,N_30364,N_31947);
or U32380 (N_32380,N_31800,N_31852);
nand U32381 (N_32381,N_30253,N_31363);
and U32382 (N_32382,N_31968,N_30468);
and U32383 (N_32383,N_31841,N_31061);
or U32384 (N_32384,N_31624,N_31039);
or U32385 (N_32385,N_31307,N_31715);
and U32386 (N_32386,N_31147,N_30350);
xnor U32387 (N_32387,N_30900,N_30605);
nand U32388 (N_32388,N_31916,N_31252);
nor U32389 (N_32389,N_31396,N_30720);
nand U32390 (N_32390,N_31469,N_30950);
nand U32391 (N_32391,N_30962,N_30953);
or U32392 (N_32392,N_31709,N_30486);
and U32393 (N_32393,N_30929,N_31204);
xor U32394 (N_32394,N_30224,N_30086);
nor U32395 (N_32395,N_30380,N_30592);
and U32396 (N_32396,N_31669,N_30979);
nor U32397 (N_32397,N_31455,N_31075);
nand U32398 (N_32398,N_31225,N_31934);
nor U32399 (N_32399,N_31954,N_30679);
or U32400 (N_32400,N_31497,N_30921);
or U32401 (N_32401,N_31811,N_30700);
or U32402 (N_32402,N_31097,N_31864);
or U32403 (N_32403,N_30521,N_30880);
or U32404 (N_32404,N_30490,N_30955);
xor U32405 (N_32405,N_30947,N_31489);
or U32406 (N_32406,N_30644,N_30707);
or U32407 (N_32407,N_30113,N_31370);
nand U32408 (N_32408,N_30836,N_31213);
nor U32409 (N_32409,N_31598,N_30677);
nor U32410 (N_32410,N_31269,N_30389);
nand U32411 (N_32411,N_31720,N_30045);
or U32412 (N_32412,N_31569,N_31038);
nor U32413 (N_32413,N_30920,N_30617);
nand U32414 (N_32414,N_30090,N_31667);
xor U32415 (N_32415,N_31358,N_31617);
or U32416 (N_32416,N_30520,N_30584);
nor U32417 (N_32417,N_30093,N_30466);
xnor U32418 (N_32418,N_30911,N_31044);
xnor U32419 (N_32419,N_30494,N_30917);
and U32420 (N_32420,N_30695,N_31821);
nor U32421 (N_32421,N_31366,N_30411);
nand U32422 (N_32422,N_30392,N_31735);
nand U32423 (N_32423,N_30586,N_30489);
nand U32424 (N_32424,N_31659,N_31440);
nor U32425 (N_32425,N_30409,N_30351);
or U32426 (N_32426,N_30874,N_31117);
nand U32427 (N_32427,N_30297,N_31683);
nand U32428 (N_32428,N_30202,N_30360);
and U32429 (N_32429,N_30796,N_31906);
nor U32430 (N_32430,N_30850,N_30064);
nand U32431 (N_32431,N_31244,N_31326);
nor U32432 (N_32432,N_31724,N_30670);
xnor U32433 (N_32433,N_30066,N_30903);
nor U32434 (N_32434,N_31476,N_31685);
nor U32435 (N_32435,N_31610,N_30273);
nand U32436 (N_32436,N_30445,N_30621);
or U32437 (N_32437,N_31101,N_30997);
nand U32438 (N_32438,N_31596,N_30795);
nand U32439 (N_32439,N_31942,N_30534);
and U32440 (N_32440,N_30526,N_30308);
xor U32441 (N_32441,N_30425,N_31888);
nand U32442 (N_32442,N_31889,N_31247);
nand U32443 (N_32443,N_30612,N_30513);
and U32444 (N_32444,N_30861,N_31431);
xor U32445 (N_32445,N_31646,N_31853);
and U32446 (N_32446,N_30501,N_30926);
nor U32447 (N_32447,N_31464,N_30858);
or U32448 (N_32448,N_30116,N_31668);
or U32449 (N_32449,N_30475,N_30647);
xnor U32450 (N_32450,N_31806,N_31799);
nor U32451 (N_32451,N_30206,N_31774);
xor U32452 (N_32452,N_31796,N_31618);
xnor U32453 (N_32453,N_31085,N_31967);
or U32454 (N_32454,N_31239,N_30133);
and U32455 (N_32455,N_31858,N_30355);
xor U32456 (N_32456,N_30103,N_30403);
and U32457 (N_32457,N_31420,N_30300);
nand U32458 (N_32458,N_31313,N_30463);
nor U32459 (N_32459,N_30177,N_30604);
and U32460 (N_32460,N_30104,N_30447);
or U32461 (N_32461,N_31202,N_31876);
nor U32462 (N_32462,N_31051,N_31143);
xor U32463 (N_32463,N_30505,N_30259);
or U32464 (N_32464,N_31778,N_30105);
and U32465 (N_32465,N_30922,N_30946);
xnor U32466 (N_32466,N_30019,N_31318);
xor U32467 (N_32467,N_30011,N_31357);
xor U32468 (N_32468,N_30047,N_31492);
or U32469 (N_32469,N_30727,N_31258);
or U32470 (N_32470,N_30150,N_31515);
nor U32471 (N_32471,N_31738,N_30991);
or U32472 (N_32472,N_31950,N_30067);
nand U32473 (N_32473,N_30051,N_31445);
nand U32474 (N_32474,N_31461,N_31551);
or U32475 (N_32475,N_30687,N_31835);
and U32476 (N_32476,N_30696,N_30325);
nand U32477 (N_32477,N_30595,N_30132);
xnor U32478 (N_32478,N_30738,N_31449);
xor U32479 (N_32479,N_31875,N_31335);
nor U32480 (N_32480,N_30079,N_31479);
nand U32481 (N_32481,N_30342,N_30023);
and U32482 (N_32482,N_30001,N_31120);
or U32483 (N_32483,N_31410,N_31165);
nor U32484 (N_32484,N_31356,N_31394);
nor U32485 (N_32485,N_30987,N_31078);
xnor U32486 (N_32486,N_31723,N_31568);
nor U32487 (N_32487,N_31966,N_31901);
and U32488 (N_32488,N_31973,N_31872);
and U32489 (N_32489,N_30030,N_30233);
or U32490 (N_32490,N_31727,N_30848);
nand U32491 (N_32491,N_31218,N_30094);
xnor U32492 (N_32492,N_30973,N_30285);
nor U32493 (N_32493,N_31867,N_30662);
nor U32494 (N_32494,N_31871,N_31712);
xnor U32495 (N_32495,N_30506,N_30870);
and U32496 (N_32496,N_30005,N_31865);
and U32497 (N_32497,N_31639,N_31291);
xor U32498 (N_32498,N_30428,N_31919);
xnor U32499 (N_32499,N_31556,N_31254);
or U32500 (N_32500,N_30992,N_31533);
and U32501 (N_32501,N_31273,N_30454);
and U32502 (N_32502,N_31834,N_31257);
nand U32503 (N_32503,N_31918,N_30792);
and U32504 (N_32504,N_30226,N_30847);
and U32505 (N_32505,N_31395,N_31698);
xnor U32506 (N_32506,N_31041,N_30554);
or U32507 (N_32507,N_31447,N_30834);
and U32508 (N_32508,N_31881,N_31958);
and U32509 (N_32509,N_30587,N_31725);
or U32510 (N_32510,N_30136,N_30242);
or U32511 (N_32511,N_30682,N_31427);
and U32512 (N_32512,N_30969,N_31119);
and U32513 (N_32513,N_30511,N_31149);
nand U32514 (N_32514,N_31074,N_30736);
and U32515 (N_32515,N_31470,N_30974);
nand U32516 (N_32516,N_31422,N_31883);
xnor U32517 (N_32517,N_30837,N_31629);
and U32518 (N_32518,N_30114,N_31785);
nand U32519 (N_32519,N_31308,N_31900);
nor U32520 (N_32520,N_30277,N_31487);
xor U32521 (N_32521,N_30835,N_31516);
or U32522 (N_32522,N_30876,N_31063);
or U32523 (N_32523,N_31650,N_30178);
xnor U32524 (N_32524,N_31351,N_31256);
nor U32525 (N_32525,N_31651,N_30611);
nor U32526 (N_32526,N_30320,N_30518);
nand U32527 (N_32527,N_31977,N_30256);
nor U32528 (N_32528,N_31962,N_30306);
or U32529 (N_32529,N_31112,N_30892);
or U32530 (N_32530,N_30442,N_30674);
nor U32531 (N_32531,N_30110,N_30443);
nand U32532 (N_32532,N_31049,N_31295);
xnor U32533 (N_32533,N_31645,N_30354);
nand U32534 (N_32534,N_31789,N_30778);
or U32535 (N_32535,N_30219,N_30126);
or U32536 (N_32536,N_30138,N_30692);
xor U32537 (N_32537,N_30699,N_30393);
nand U32538 (N_32538,N_30009,N_31020);
nor U32539 (N_32539,N_30303,N_30000);
and U32540 (N_32540,N_30333,N_31280);
nand U32541 (N_32541,N_30542,N_30170);
and U32542 (N_32542,N_31937,N_30764);
nor U32543 (N_32543,N_31272,N_31747);
or U32544 (N_32544,N_31083,N_31321);
nand U32545 (N_32545,N_30763,N_31368);
and U32546 (N_32546,N_30704,N_31141);
or U32547 (N_32547,N_31843,N_31953);
or U32548 (N_32548,N_31877,N_30675);
nand U32549 (N_32549,N_31628,N_31912);
and U32550 (N_32550,N_30912,N_31344);
nor U32551 (N_32551,N_31133,N_30190);
nor U32552 (N_32552,N_31378,N_31330);
xor U32553 (N_32553,N_31879,N_31981);
nand U32554 (N_32554,N_31581,N_31930);
and U32555 (N_32555,N_30556,N_31660);
or U32556 (N_32556,N_31621,N_30514);
xor U32557 (N_32557,N_31438,N_30469);
or U32558 (N_32558,N_30455,N_31936);
xor U32559 (N_32559,N_31748,N_30495);
xnor U32560 (N_32560,N_30161,N_31249);
nand U32561 (N_32561,N_31801,N_31710);
nand U32562 (N_32562,N_30063,N_30528);
and U32563 (N_32563,N_30797,N_31176);
xnor U32564 (N_32564,N_31975,N_30760);
or U32565 (N_32565,N_31232,N_30525);
or U32566 (N_32566,N_31472,N_30153);
nand U32567 (N_32567,N_31301,N_30382);
nand U32568 (N_32568,N_30799,N_30498);
xor U32569 (N_32569,N_30203,N_31976);
and U32570 (N_32570,N_31373,N_30311);
nand U32571 (N_32571,N_30976,N_31223);
xnor U32572 (N_32572,N_30039,N_30027);
nand U32573 (N_32573,N_30547,N_30235);
and U32574 (N_32574,N_30723,N_30924);
nand U32575 (N_32575,N_31663,N_31043);
nor U32576 (N_32576,N_30522,N_30369);
or U32577 (N_32577,N_30423,N_31517);
or U32578 (N_32578,N_31850,N_30970);
nor U32579 (N_32579,N_30464,N_30923);
or U32580 (N_32580,N_31704,N_30714);
nand U32581 (N_32581,N_30883,N_31279);
or U32582 (N_32582,N_30747,N_30739);
or U32583 (N_32583,N_30952,N_31070);
nor U32584 (N_32584,N_31425,N_30650);
xnor U32585 (N_32585,N_30054,N_31677);
and U32586 (N_32586,N_30618,N_31106);
xnor U32587 (N_32587,N_30571,N_31138);
and U32588 (N_32588,N_31317,N_31381);
nand U32589 (N_32589,N_31578,N_30807);
and U32590 (N_32590,N_31920,N_31729);
xnor U32591 (N_32591,N_30289,N_30895);
or U32592 (N_32592,N_31006,N_30805);
or U32593 (N_32593,N_31343,N_31868);
nand U32594 (N_32594,N_31974,N_31371);
nor U32595 (N_32595,N_30544,N_30909);
nand U32596 (N_32596,N_30568,N_30743);
nand U32597 (N_32597,N_31570,N_31963);
nand U32598 (N_32598,N_30809,N_31759);
and U32599 (N_32599,N_31012,N_31161);
nor U32600 (N_32600,N_30708,N_30770);
xor U32601 (N_32601,N_30508,N_30046);
nand U32602 (N_32602,N_30467,N_30033);
and U32603 (N_32603,N_31148,N_30935);
xnor U32604 (N_32604,N_31072,N_30734);
nand U32605 (N_32605,N_31573,N_31352);
and U32606 (N_32606,N_30336,N_31510);
or U32607 (N_32607,N_30186,N_31136);
and U32608 (N_32608,N_31364,N_31894);
nand U32609 (N_32609,N_30881,N_30507);
or U32610 (N_32610,N_30693,N_30919);
nor U32611 (N_32611,N_30937,N_31393);
or U32612 (N_32612,N_30158,N_30593);
or U32613 (N_32613,N_30385,N_31341);
or U32614 (N_32614,N_31595,N_30257);
nand U32615 (N_32615,N_30543,N_30993);
or U32616 (N_32616,N_31780,N_30358);
and U32617 (N_32617,N_30056,N_31505);
nand U32618 (N_32618,N_31135,N_30574);
and U32619 (N_32619,N_30688,N_30271);
nor U32620 (N_32620,N_31402,N_30575);
or U32621 (N_32621,N_31700,N_31994);
nand U32622 (N_32622,N_30195,N_30345);
xnor U32623 (N_32623,N_30888,N_31575);
and U32624 (N_32624,N_31156,N_30143);
xor U32625 (N_32625,N_30437,N_30139);
xor U32626 (N_32626,N_30034,N_30954);
xor U32627 (N_32627,N_31499,N_31844);
nand U32628 (N_32628,N_30965,N_31379);
nand U32629 (N_32629,N_31248,N_31267);
nor U32630 (N_32630,N_30761,N_31398);
or U32631 (N_32631,N_31899,N_30117);
nand U32632 (N_32632,N_30769,N_30433);
nor U32633 (N_32633,N_30533,N_31713);
or U32634 (N_32634,N_30266,N_30310);
nor U32635 (N_32635,N_31421,N_31897);
xor U32636 (N_32636,N_31817,N_31486);
or U32637 (N_32637,N_31302,N_31227);
nand U32638 (N_32638,N_30020,N_31902);
nand U32639 (N_32639,N_30884,N_31163);
xnor U32640 (N_32640,N_31229,N_31436);
nor U32641 (N_32641,N_30539,N_31815);
nor U32642 (N_32642,N_31208,N_31955);
xor U32643 (N_32643,N_31619,N_30906);
and U32644 (N_32644,N_31684,N_30683);
nor U32645 (N_32645,N_30307,N_31056);
nand U32646 (N_32646,N_30804,N_31500);
and U32647 (N_32647,N_31286,N_30473);
or U32648 (N_32648,N_30100,N_31221);
nor U32649 (N_32649,N_30752,N_31387);
nor U32650 (N_32650,N_30479,N_31312);
or U32651 (N_32651,N_31730,N_30905);
nand U32652 (N_32652,N_30077,N_30934);
or U32653 (N_32653,N_30283,N_30072);
or U32654 (N_32654,N_30773,N_30572);
or U32655 (N_32655,N_31222,N_30907);
xor U32656 (N_32656,N_31717,N_31790);
and U32657 (N_32657,N_30827,N_30729);
xor U32658 (N_32658,N_30068,N_30160);
nor U32659 (N_32659,N_30634,N_30349);
or U32660 (N_32660,N_31561,N_30041);
xnor U32661 (N_32661,N_30395,N_30182);
and U32662 (N_32662,N_31991,N_31060);
or U32663 (N_32663,N_31298,N_30532);
xor U32664 (N_32664,N_30655,N_31082);
or U32665 (N_32665,N_31931,N_30812);
nand U32666 (N_32666,N_30749,N_30474);
nand U32667 (N_32667,N_30994,N_31545);
xor U32668 (N_32668,N_30666,N_31538);
or U32669 (N_32669,N_30483,N_30619);
nand U32670 (N_32670,N_30268,N_31177);
nor U32671 (N_32671,N_30061,N_30597);
or U32672 (N_32672,N_30316,N_30118);
nor U32673 (N_32673,N_30766,N_30989);
nand U32674 (N_32674,N_31605,N_30630);
nand U32675 (N_32675,N_31536,N_31331);
nand U32676 (N_32676,N_30073,N_31151);
nor U32677 (N_32677,N_31798,N_30960);
nand U32678 (N_32678,N_31123,N_30933);
or U32679 (N_32679,N_30972,N_31337);
and U32680 (N_32680,N_30814,N_30600);
xor U32681 (N_32681,N_31603,N_31329);
or U32682 (N_32682,N_31644,N_30021);
xnor U32683 (N_32683,N_31636,N_31434);
and U32684 (N_32684,N_31360,N_30844);
nor U32685 (N_32685,N_31274,N_30867);
nand U32686 (N_32686,N_31592,N_30029);
nand U32687 (N_32687,N_31711,N_31004);
nor U32688 (N_32688,N_30159,N_31773);
nand U32689 (N_32689,N_30872,N_30223);
nand U32690 (N_32690,N_31359,N_31325);
and U32691 (N_32691,N_30999,N_31322);
or U32692 (N_32692,N_30889,N_31145);
nand U32693 (N_32693,N_30147,N_31064);
and U32694 (N_32694,N_31294,N_31124);
xor U32695 (N_32695,N_30887,N_30596);
or U32696 (N_32696,N_30431,N_31999);
nor U32697 (N_32697,N_30781,N_31450);
and U32698 (N_32698,N_31243,N_31827);
xor U32699 (N_32699,N_30315,N_30964);
or U32700 (N_32700,N_31348,N_30594);
nor U32701 (N_32701,N_30524,N_31009);
xor U32702 (N_32702,N_30098,N_30387);
or U32703 (N_32703,N_31742,N_30886);
and U32704 (N_32704,N_31786,N_30435);
and U32705 (N_32705,N_31214,N_30076);
nor U32706 (N_32706,N_30148,N_31386);
nand U32707 (N_32707,N_31429,N_30085);
nor U32708 (N_32708,N_31052,N_31809);
nand U32709 (N_32709,N_31311,N_31209);
or U32710 (N_32710,N_30877,N_31716);
or U32711 (N_32711,N_30607,N_31768);
and U32712 (N_32712,N_30296,N_31109);
and U32713 (N_32713,N_30172,N_31432);
nor U32714 (N_32714,N_31637,N_31532);
and U32715 (N_32715,N_31803,N_31259);
xor U32716 (N_32716,N_30078,N_30839);
or U32717 (N_32717,N_31406,N_30371);
nor U32718 (N_32718,N_30165,N_31993);
nand U32719 (N_32719,N_31245,N_30346);
nor U32720 (N_32720,N_30914,N_31733);
or U32721 (N_32721,N_30515,N_31869);
nand U32722 (N_32722,N_31765,N_30488);
and U32723 (N_32723,N_30044,N_31736);
and U32724 (N_32724,N_31842,N_31306);
xnor U32725 (N_32725,N_31404,N_30441);
nand U32726 (N_32726,N_31220,N_31108);
nand U32727 (N_32727,N_30819,N_30681);
or U32728 (N_32728,N_31836,N_30578);
xnor U32729 (N_32729,N_30902,N_31828);
xor U32730 (N_32730,N_30359,N_30982);
or U32731 (N_32731,N_31558,N_31144);
nand U32732 (N_32732,N_31293,N_31506);
nor U32733 (N_32733,N_31200,N_31090);
xnor U32734 (N_32734,N_30737,N_30928);
xor U32735 (N_32735,N_30040,N_30753);
xor U32736 (N_32736,N_30174,N_30741);
xor U32737 (N_32737,N_31098,N_30717);
nor U32738 (N_32738,N_31374,N_31549);
or U32739 (N_32739,N_30309,N_30813);
and U32740 (N_32740,N_31664,N_30274);
and U32741 (N_32741,N_30856,N_31206);
xnor U32742 (N_32742,N_30430,N_30457);
xnor U32743 (N_32743,N_30412,N_31441);
nor U32744 (N_32744,N_31678,N_31566);
xnor U32745 (N_32745,N_31956,N_30601);
and U32746 (N_32746,N_31513,N_30317);
nand U32747 (N_32747,N_31708,N_30211);
or U32748 (N_32748,N_30450,N_31642);
nor U32749 (N_32749,N_31342,N_31554);
and U32750 (N_32750,N_31196,N_30570);
xor U32751 (N_32751,N_31989,N_31309);
xnor U32752 (N_32752,N_31048,N_31804);
or U32753 (N_32753,N_30555,N_30671);
nand U32754 (N_32754,N_30312,N_30551);
or U32755 (N_32755,N_30573,N_30938);
xnor U32756 (N_32756,N_31047,N_30062);
or U32757 (N_32757,N_31215,N_30262);
xor U32758 (N_32758,N_30386,N_31819);
or U32759 (N_32759,N_31616,N_31714);
xnor U32760 (N_32760,N_30751,N_30694);
and U32761 (N_32761,N_31069,N_31010);
nor U32762 (N_32762,N_31319,N_30293);
and U32763 (N_32763,N_31658,N_31652);
nor U32764 (N_32764,N_30811,N_30869);
or U32765 (N_32765,N_31537,N_31863);
nand U32766 (N_32766,N_30439,N_31761);
and U32767 (N_32767,N_30087,N_31927);
nand U32768 (N_32768,N_30493,N_30227);
xnor U32769 (N_32769,N_30280,N_31757);
or U32770 (N_32770,N_30966,N_30344);
nand U32771 (N_32771,N_30659,N_30803);
nor U32772 (N_32772,N_30260,N_30229);
or U32773 (N_32773,N_31945,N_31587);
and U32774 (N_32774,N_31929,N_31957);
nand U32775 (N_32775,N_30641,N_31277);
nand U32776 (N_32776,N_31521,N_31776);
nand U32777 (N_32777,N_30845,N_30706);
and U32778 (N_32778,N_30329,N_31091);
and U32779 (N_32779,N_31219,N_31680);
nor U32780 (N_32780,N_31769,N_30686);
nor U32781 (N_32781,N_31997,N_30616);
xor U32782 (N_32782,N_31261,N_31187);
nor U32783 (N_32783,N_30102,N_31389);
and U32784 (N_32784,N_30613,N_31722);
nand U32785 (N_32785,N_31169,N_30896);
nand U32786 (N_32786,N_31347,N_31055);
nor U32787 (N_32787,N_30043,N_30427);
nor U32788 (N_32788,N_31021,N_31837);
nand U32789 (N_32789,N_31990,N_31416);
nor U32790 (N_32790,N_30060,N_30048);
nor U32791 (N_32791,N_30168,N_30732);
xnor U32792 (N_32792,N_30022,N_30620);
nand U32793 (N_32793,N_30149,N_31996);
nor U32794 (N_32794,N_30567,N_30331);
nor U32795 (N_32795,N_31016,N_31481);
and U32796 (N_32796,N_30236,N_31132);
xor U32797 (N_32797,N_31153,N_31488);
nand U32798 (N_32798,N_31456,N_30776);
and U32799 (N_32799,N_30502,N_31042);
and U32800 (N_32800,N_30156,N_30560);
nand U32801 (N_32801,N_31608,N_31423);
nor U32802 (N_32802,N_31822,N_31392);
and U32803 (N_32803,N_30794,N_30801);
nand U32804 (N_32804,N_30629,N_31007);
xnor U32805 (N_32805,N_31408,N_30415);
xor U32806 (N_32806,N_31560,N_30957);
and U32807 (N_32807,N_30140,N_31788);
nand U32808 (N_32808,N_31908,N_31401);
nor U32809 (N_32809,N_30637,N_30292);
nor U32810 (N_32810,N_30276,N_31907);
nor U32811 (N_32811,N_30598,N_30624);
and U32812 (N_32812,N_31760,N_30948);
nor U32813 (N_32813,N_31336,N_30940);
xnor U32814 (N_32814,N_30321,N_30846);
or U32815 (N_32815,N_31362,N_30774);
or U32816 (N_32816,N_31745,N_31115);
nor U32817 (N_32817,N_31460,N_31998);
nand U32818 (N_32818,N_30208,N_31182);
nor U32819 (N_32819,N_30711,N_31866);
and U32820 (N_32820,N_31300,N_30383);
or U32821 (N_32821,N_30137,N_31040);
xor U32822 (N_32822,N_30417,N_30622);
nor U32823 (N_32823,N_30638,N_31412);
or U32824 (N_32824,N_30220,N_31764);
nand U32825 (N_32825,N_31657,N_31139);
nand U32826 (N_32826,N_30207,N_30420);
and U32827 (N_32827,N_30632,N_31654);
nor U32828 (N_32828,N_30304,N_31793);
xor U32829 (N_32829,N_31583,N_30893);
nand U32830 (N_32830,N_30084,N_31703);
or U32831 (N_32831,N_30951,N_31600);
nor U32832 (N_32832,N_31965,N_31129);
and U32833 (N_32833,N_30216,N_31454);
or U32834 (N_32834,N_31952,N_31531);
or U32835 (N_32835,N_31731,N_31690);
nor U32836 (N_32836,N_31812,N_30816);
nand U32837 (N_32837,N_31443,N_31264);
or U32838 (N_32838,N_31234,N_30080);
nand U32839 (N_32839,N_30053,N_31813);
nand U32840 (N_32840,N_31435,N_31405);
xnor U32841 (N_32841,N_30365,N_30171);
nand U32842 (N_32842,N_31826,N_31216);
nand U32843 (N_32843,N_31971,N_30477);
and U32844 (N_32844,N_31316,N_31833);
nor U32845 (N_32845,N_30782,N_30050);
nand U32846 (N_32846,N_30899,N_30368);
nor U32847 (N_32847,N_30590,N_31471);
and U32848 (N_32848,N_31601,N_30985);
xnor U32849 (N_32849,N_31114,N_31242);
xnor U32850 (N_32850,N_30347,N_30852);
and U32851 (N_32851,N_30180,N_31586);
or U32852 (N_32852,N_31522,N_31604);
nand U32853 (N_32853,N_31338,N_31134);
or U32854 (N_32854,N_31260,N_31096);
nor U32855 (N_32855,N_31409,N_31211);
nor U32856 (N_32856,N_30626,N_30017);
or U32857 (N_32857,N_31185,N_31495);
nand U32858 (N_32858,N_31017,N_31253);
nand U32859 (N_32859,N_30824,N_31818);
nor U32860 (N_32860,N_30669,N_31767);
and U32861 (N_32861,N_31896,N_31305);
nand U32862 (N_32862,N_31756,N_30356);
or U32863 (N_32863,N_31193,N_31940);
or U32864 (N_32864,N_31323,N_31314);
nor U32865 (N_32865,N_31369,N_31210);
nor U32866 (N_32866,N_31891,N_31987);
xor U32867 (N_32867,N_31870,N_31297);
or U32868 (N_32868,N_30936,N_31641);
xor U32869 (N_32869,N_31292,N_31859);
nor U32870 (N_32870,N_31415,N_31237);
nor U32871 (N_32871,N_31095,N_30791);
xor U32872 (N_32872,N_30261,N_30577);
and U32873 (N_32873,N_30746,N_30610);
xnor U32874 (N_32874,N_31855,N_30426);
xnor U32875 (N_32875,N_31824,N_30959);
and U32876 (N_32876,N_31699,N_31164);
xnor U32877 (N_32877,N_31474,N_31390);
nor U32878 (N_32878,N_30446,N_30968);
or U32879 (N_32879,N_31375,N_31749);
and U32880 (N_32880,N_30418,N_30579);
nand U32881 (N_32881,N_30166,N_31594);
nand U32882 (N_32882,N_30497,N_31110);
xor U32883 (N_32883,N_31299,N_30341);
xor U32884 (N_32884,N_30278,N_30866);
nand U32885 (N_32885,N_30363,N_30462);
or U32886 (N_32886,N_30548,N_30684);
nor U32887 (N_32887,N_31661,N_31509);
nand U32888 (N_32888,N_30032,N_31914);
nor U32889 (N_32889,N_31797,N_31458);
xnor U32890 (N_32890,N_30559,N_31079);
or U32891 (N_32891,N_30374,N_31527);
xor U32892 (N_32892,N_30631,N_30313);
and U32893 (N_32893,N_30096,N_30406);
nand U32894 (N_32894,N_31656,N_30673);
or U32895 (N_32895,N_31478,N_30726);
nor U32896 (N_32896,N_30106,N_30891);
xnor U32897 (N_32897,N_30327,N_30471);
nand U32898 (N_32898,N_30983,N_30157);
nor U32899 (N_32899,N_31921,N_30405);
or U32900 (N_32900,N_31172,N_31290);
and U32901 (N_32901,N_31978,N_31518);
and U32902 (N_32902,N_30007,N_30725);
or U32903 (N_32903,N_31550,N_30252);
and U32904 (N_32904,N_30228,N_31170);
nor U32905 (N_32905,N_30633,N_31304);
or U32906 (N_32906,N_30173,N_30879);
or U32907 (N_32907,N_31372,N_31938);
nand U32908 (N_32908,N_31397,N_31418);
nor U32909 (N_32909,N_30101,N_30376);
and U32910 (N_32910,N_30031,N_31467);
nor U32911 (N_32911,N_31665,N_30459);
nand U32912 (N_32912,N_31452,N_30496);
or U32913 (N_32913,N_31904,N_30121);
or U32914 (N_32914,N_30402,N_30452);
xnor U32915 (N_32915,N_31946,N_31066);
nand U32916 (N_32916,N_30142,N_31839);
and U32917 (N_32917,N_31059,N_30663);
or U32918 (N_32918,N_30820,N_30740);
or U32919 (N_32919,N_30540,N_30823);
nor U32920 (N_32920,N_30299,N_31382);
nand U32921 (N_32921,N_30831,N_30154);
or U32922 (N_32922,N_31674,N_31701);
or U32923 (N_32923,N_30731,N_30127);
nand U32924 (N_32924,N_30665,N_31367);
xor U32925 (N_32925,N_30748,N_31361);
and U32926 (N_32926,N_31911,N_30092);
xor U32927 (N_32927,N_30145,N_30284);
and U32928 (N_32928,N_31503,N_30785);
xor U32929 (N_32929,N_30408,N_30564);
nand U32930 (N_32930,N_30742,N_31862);
nor U32931 (N_32931,N_31555,N_31969);
nor U32932 (N_32932,N_31933,N_31159);
xor U32933 (N_32933,N_30290,N_30651);
xnor U32934 (N_32934,N_31231,N_30589);
xor U32935 (N_32935,N_30055,N_31178);
nor U32936 (N_32936,N_30685,N_31886);
nand U32937 (N_32937,N_30810,N_31540);
xnor U32938 (N_32938,N_30509,N_31944);
xnor U32939 (N_32939,N_31941,N_30424);
nor U32940 (N_32940,N_31166,N_30857);
nand U32941 (N_32941,N_30800,N_31576);
and U32942 (N_32942,N_31625,N_31640);
nand U32943 (N_32943,N_30366,N_30015);
and U32944 (N_32944,N_31482,N_31557);
nor U32945 (N_32945,N_31045,N_31792);
xor U32946 (N_32946,N_31626,N_30367);
and U32947 (N_32947,N_30460,N_30194);
nor U32948 (N_32948,N_30913,N_31288);
nor U32949 (N_32949,N_30504,N_31860);
and U32950 (N_32950,N_30580,N_30416);
xnor U32951 (N_32951,N_30915,N_30981);
nand U32952 (N_32952,N_31563,N_30853);
nor U32953 (N_32953,N_31093,N_30798);
and U32954 (N_32954,N_30287,N_31873);
or U32955 (N_32955,N_30538,N_31577);
nand U32956 (N_32956,N_30243,N_30215);
or U32957 (N_32957,N_31207,N_31707);
nand U32958 (N_32958,N_30628,N_30829);
xor U32959 (N_32959,N_31737,N_30245);
nand U32960 (N_32960,N_30119,N_30722);
xor U32961 (N_32961,N_31199,N_30314);
nand U32962 (N_32962,N_31000,N_31430);
nand U32963 (N_32963,N_31175,N_30712);
or U32964 (N_32964,N_31632,N_30757);
nor U32965 (N_32965,N_31831,N_30854);
xor U32966 (N_32966,N_30197,N_31233);
or U32967 (N_32967,N_30295,N_30008);
and U32968 (N_32968,N_31926,N_31589);
xnor U32969 (N_32969,N_31694,N_31077);
nor U32970 (N_32970,N_31089,N_31571);
or U32971 (N_32971,N_30698,N_31754);
and U32972 (N_32972,N_30196,N_30038);
xnor U32973 (N_32973,N_31003,N_30254);
and U32974 (N_32974,N_31653,N_30334);
nor U32975 (N_32975,N_30485,N_31162);
xor U32976 (N_32976,N_30144,N_31988);
nand U32977 (N_32977,N_31023,N_31861);
and U32978 (N_32978,N_31829,N_30429);
or U32979 (N_32979,N_30288,N_31559);
nor U32980 (N_32980,N_31324,N_30124);
xnor U32981 (N_32981,N_31022,N_31065);
and U32982 (N_32982,N_31620,N_30932);
nor U32983 (N_32983,N_30362,N_31174);
or U32984 (N_32984,N_30925,N_30672);
xor U32985 (N_32985,N_30264,N_31995);
and U32986 (N_32986,N_30894,N_30199);
xor U32987 (N_32987,N_31544,N_31480);
nand U32988 (N_32988,N_31268,N_31484);
or U32989 (N_32989,N_31567,N_31823);
and U32990 (N_32990,N_30129,N_31743);
nor U32991 (N_32991,N_30152,N_31477);
nand U32992 (N_32992,N_31623,N_30602);
nor U32993 (N_32993,N_30192,N_31426);
and U32994 (N_32994,N_30639,N_30697);
nor U32995 (N_32995,N_31081,N_31758);
or U32996 (N_32996,N_30986,N_31903);
nor U32997 (N_32997,N_30581,N_31315);
xnor U32998 (N_32998,N_31407,N_30765);
or U32999 (N_32999,N_30585,N_31437);
or U33000 (N_33000,N_30751,N_30254);
nor U33001 (N_33001,N_30620,N_30998);
nor U33002 (N_33002,N_30979,N_31954);
or U33003 (N_33003,N_31950,N_30581);
and U33004 (N_33004,N_30850,N_30282);
or U33005 (N_33005,N_30199,N_31628);
and U33006 (N_33006,N_30639,N_31160);
xnor U33007 (N_33007,N_30015,N_31893);
nand U33008 (N_33008,N_30994,N_31126);
and U33009 (N_33009,N_30539,N_31044);
nor U33010 (N_33010,N_30135,N_31902);
or U33011 (N_33011,N_30958,N_31587);
or U33012 (N_33012,N_31560,N_31376);
xor U33013 (N_33013,N_31016,N_30112);
and U33014 (N_33014,N_30791,N_30849);
nand U33015 (N_33015,N_31309,N_31099);
and U33016 (N_33016,N_30806,N_31892);
nor U33017 (N_33017,N_30648,N_30403);
xnor U33018 (N_33018,N_31077,N_30727);
xor U33019 (N_33019,N_30584,N_31475);
xor U33020 (N_33020,N_30352,N_31919);
and U33021 (N_33021,N_30349,N_30103);
nand U33022 (N_33022,N_30678,N_30392);
nor U33023 (N_33023,N_31140,N_31606);
or U33024 (N_33024,N_31913,N_30922);
or U33025 (N_33025,N_31698,N_31359);
nor U33026 (N_33026,N_30477,N_31694);
xnor U33027 (N_33027,N_30106,N_30437);
or U33028 (N_33028,N_30463,N_31837);
nand U33029 (N_33029,N_31646,N_31095);
nor U33030 (N_33030,N_30678,N_31318);
nand U33031 (N_33031,N_30954,N_30895);
nor U33032 (N_33032,N_30700,N_30483);
or U33033 (N_33033,N_31598,N_30230);
and U33034 (N_33034,N_31749,N_31236);
nor U33035 (N_33035,N_30133,N_31216);
or U33036 (N_33036,N_31377,N_31405);
or U33037 (N_33037,N_30152,N_30624);
xor U33038 (N_33038,N_31180,N_31294);
and U33039 (N_33039,N_31174,N_31212);
or U33040 (N_33040,N_30176,N_31394);
and U33041 (N_33041,N_30665,N_31588);
nand U33042 (N_33042,N_31025,N_30155);
nand U33043 (N_33043,N_31563,N_31958);
and U33044 (N_33044,N_30744,N_31339);
and U33045 (N_33045,N_30933,N_31945);
or U33046 (N_33046,N_31118,N_30867);
nor U33047 (N_33047,N_30277,N_30715);
xor U33048 (N_33048,N_31860,N_30068);
and U33049 (N_33049,N_31784,N_31841);
and U33050 (N_33050,N_30828,N_30381);
and U33051 (N_33051,N_30709,N_30701);
or U33052 (N_33052,N_30522,N_31799);
xnor U33053 (N_33053,N_31431,N_31240);
nor U33054 (N_33054,N_31234,N_30230);
and U33055 (N_33055,N_31229,N_31058);
or U33056 (N_33056,N_30138,N_30058);
and U33057 (N_33057,N_30939,N_30256);
nor U33058 (N_33058,N_31555,N_30964);
nor U33059 (N_33059,N_30311,N_31803);
nand U33060 (N_33060,N_31897,N_31776);
or U33061 (N_33061,N_31855,N_31263);
nand U33062 (N_33062,N_31346,N_30121);
and U33063 (N_33063,N_30531,N_31876);
or U33064 (N_33064,N_30560,N_31054);
xnor U33065 (N_33065,N_30999,N_30360);
nor U33066 (N_33066,N_30176,N_31602);
nand U33067 (N_33067,N_30842,N_30088);
nor U33068 (N_33068,N_31486,N_30628);
xnor U33069 (N_33069,N_30369,N_31852);
or U33070 (N_33070,N_30108,N_30788);
or U33071 (N_33071,N_31802,N_30346);
and U33072 (N_33072,N_31775,N_30851);
and U33073 (N_33073,N_30038,N_31145);
nand U33074 (N_33074,N_30104,N_30747);
or U33075 (N_33075,N_30542,N_30831);
xnor U33076 (N_33076,N_31110,N_31634);
or U33077 (N_33077,N_30755,N_30563);
nor U33078 (N_33078,N_31035,N_30151);
and U33079 (N_33079,N_31391,N_31523);
xor U33080 (N_33080,N_30178,N_30473);
nand U33081 (N_33081,N_30033,N_30650);
nand U33082 (N_33082,N_31616,N_30260);
nor U33083 (N_33083,N_31760,N_30745);
nand U33084 (N_33084,N_30889,N_31251);
or U33085 (N_33085,N_30557,N_31766);
xnor U33086 (N_33086,N_31363,N_30594);
nand U33087 (N_33087,N_31028,N_31405);
or U33088 (N_33088,N_30331,N_30850);
or U33089 (N_33089,N_31099,N_31223);
and U33090 (N_33090,N_30320,N_31063);
nor U33091 (N_33091,N_31723,N_31857);
nand U33092 (N_33092,N_31894,N_30357);
or U33093 (N_33093,N_30136,N_30755);
xor U33094 (N_33094,N_30203,N_30036);
nor U33095 (N_33095,N_31667,N_30870);
and U33096 (N_33096,N_31455,N_30731);
xnor U33097 (N_33097,N_30572,N_31681);
and U33098 (N_33098,N_31170,N_31009);
nor U33099 (N_33099,N_30261,N_31186);
or U33100 (N_33100,N_30891,N_31086);
nor U33101 (N_33101,N_31513,N_31566);
xnor U33102 (N_33102,N_31068,N_30349);
xor U33103 (N_33103,N_31812,N_30168);
or U33104 (N_33104,N_31016,N_31316);
nor U33105 (N_33105,N_31071,N_30924);
nand U33106 (N_33106,N_30596,N_30484);
nor U33107 (N_33107,N_31911,N_30244);
nand U33108 (N_33108,N_31739,N_31390);
xor U33109 (N_33109,N_30674,N_30799);
xnor U33110 (N_33110,N_30123,N_30840);
and U33111 (N_33111,N_31699,N_30539);
xnor U33112 (N_33112,N_30351,N_30027);
nand U33113 (N_33113,N_30791,N_30817);
or U33114 (N_33114,N_31098,N_30216);
and U33115 (N_33115,N_31617,N_30156);
or U33116 (N_33116,N_30855,N_31243);
xor U33117 (N_33117,N_30644,N_31964);
nor U33118 (N_33118,N_31747,N_31623);
xor U33119 (N_33119,N_31912,N_31816);
or U33120 (N_33120,N_30630,N_31088);
xnor U33121 (N_33121,N_31556,N_31367);
and U33122 (N_33122,N_31445,N_30983);
xnor U33123 (N_33123,N_30088,N_31414);
or U33124 (N_33124,N_30531,N_31093);
nor U33125 (N_33125,N_30334,N_31499);
and U33126 (N_33126,N_30819,N_31148);
or U33127 (N_33127,N_31554,N_30144);
xnor U33128 (N_33128,N_31121,N_31020);
nand U33129 (N_33129,N_31108,N_31717);
and U33130 (N_33130,N_30514,N_31997);
or U33131 (N_33131,N_31721,N_30259);
and U33132 (N_33132,N_30673,N_31496);
xor U33133 (N_33133,N_31259,N_30743);
or U33134 (N_33134,N_31501,N_30358);
or U33135 (N_33135,N_30931,N_31322);
or U33136 (N_33136,N_31088,N_30199);
and U33137 (N_33137,N_30348,N_30419);
and U33138 (N_33138,N_30890,N_30920);
nor U33139 (N_33139,N_30127,N_31304);
nand U33140 (N_33140,N_31117,N_31096);
nor U33141 (N_33141,N_30606,N_31899);
nand U33142 (N_33142,N_31473,N_30541);
or U33143 (N_33143,N_31264,N_31517);
nand U33144 (N_33144,N_30178,N_31572);
nand U33145 (N_33145,N_30697,N_30412);
and U33146 (N_33146,N_31229,N_31893);
and U33147 (N_33147,N_30721,N_30502);
or U33148 (N_33148,N_31795,N_30578);
or U33149 (N_33149,N_30973,N_30903);
nor U33150 (N_33150,N_30004,N_31047);
nand U33151 (N_33151,N_30863,N_30423);
or U33152 (N_33152,N_30986,N_30401);
nand U33153 (N_33153,N_30638,N_31687);
or U33154 (N_33154,N_30416,N_31600);
nor U33155 (N_33155,N_31043,N_31047);
xor U33156 (N_33156,N_30235,N_30075);
nand U33157 (N_33157,N_30170,N_31355);
nand U33158 (N_33158,N_31319,N_30347);
or U33159 (N_33159,N_31107,N_31274);
nor U33160 (N_33160,N_31788,N_30731);
and U33161 (N_33161,N_30918,N_30093);
nor U33162 (N_33162,N_31978,N_30038);
nand U33163 (N_33163,N_30642,N_30882);
and U33164 (N_33164,N_30102,N_31436);
nor U33165 (N_33165,N_31071,N_31849);
or U33166 (N_33166,N_31685,N_31504);
or U33167 (N_33167,N_31205,N_31065);
and U33168 (N_33168,N_30534,N_31078);
nand U33169 (N_33169,N_30587,N_31247);
nor U33170 (N_33170,N_31921,N_30701);
nor U33171 (N_33171,N_31144,N_30959);
nand U33172 (N_33172,N_31151,N_30683);
xor U33173 (N_33173,N_31325,N_30234);
nand U33174 (N_33174,N_31790,N_30900);
nand U33175 (N_33175,N_30965,N_30409);
nand U33176 (N_33176,N_30065,N_31238);
nand U33177 (N_33177,N_30025,N_30760);
or U33178 (N_33178,N_31217,N_30369);
and U33179 (N_33179,N_31011,N_31504);
xor U33180 (N_33180,N_31877,N_31457);
and U33181 (N_33181,N_31838,N_30024);
nand U33182 (N_33182,N_30869,N_31620);
xnor U33183 (N_33183,N_31348,N_30303);
nor U33184 (N_33184,N_31341,N_31696);
nor U33185 (N_33185,N_31006,N_30936);
xor U33186 (N_33186,N_30022,N_31089);
and U33187 (N_33187,N_31306,N_31190);
nor U33188 (N_33188,N_30674,N_30698);
xnor U33189 (N_33189,N_31498,N_30645);
nor U33190 (N_33190,N_30758,N_30215);
nand U33191 (N_33191,N_31636,N_31396);
xor U33192 (N_33192,N_30083,N_30609);
or U33193 (N_33193,N_30776,N_31333);
nor U33194 (N_33194,N_31900,N_31501);
xor U33195 (N_33195,N_31936,N_31900);
or U33196 (N_33196,N_31637,N_30448);
nand U33197 (N_33197,N_30875,N_31736);
xnor U33198 (N_33198,N_30994,N_30484);
or U33199 (N_33199,N_31136,N_30265);
nand U33200 (N_33200,N_31357,N_30518);
and U33201 (N_33201,N_30517,N_31899);
and U33202 (N_33202,N_31196,N_30982);
and U33203 (N_33203,N_31678,N_31856);
nand U33204 (N_33204,N_30255,N_30456);
or U33205 (N_33205,N_31997,N_30751);
xor U33206 (N_33206,N_31495,N_30731);
or U33207 (N_33207,N_30531,N_31845);
and U33208 (N_33208,N_30914,N_31877);
nand U33209 (N_33209,N_31770,N_31572);
and U33210 (N_33210,N_30980,N_30144);
or U33211 (N_33211,N_30055,N_31860);
xor U33212 (N_33212,N_30170,N_30731);
and U33213 (N_33213,N_30054,N_30871);
nand U33214 (N_33214,N_30609,N_30588);
nor U33215 (N_33215,N_31102,N_31836);
or U33216 (N_33216,N_30148,N_30644);
xnor U33217 (N_33217,N_30917,N_30500);
and U33218 (N_33218,N_30495,N_31244);
nor U33219 (N_33219,N_30832,N_30173);
nand U33220 (N_33220,N_31414,N_31506);
and U33221 (N_33221,N_30073,N_31930);
or U33222 (N_33222,N_31180,N_31740);
nor U33223 (N_33223,N_30133,N_30399);
and U33224 (N_33224,N_30739,N_30308);
or U33225 (N_33225,N_31984,N_30468);
nor U33226 (N_33226,N_30964,N_31738);
and U33227 (N_33227,N_31817,N_30529);
xnor U33228 (N_33228,N_31007,N_30604);
or U33229 (N_33229,N_30568,N_31591);
nor U33230 (N_33230,N_31192,N_30307);
xor U33231 (N_33231,N_31911,N_31767);
nand U33232 (N_33232,N_30766,N_30090);
nand U33233 (N_33233,N_31097,N_30147);
nor U33234 (N_33234,N_31536,N_31620);
nand U33235 (N_33235,N_30366,N_31717);
and U33236 (N_33236,N_31259,N_30070);
nor U33237 (N_33237,N_31869,N_30870);
xnor U33238 (N_33238,N_30730,N_31452);
and U33239 (N_33239,N_30855,N_31720);
xnor U33240 (N_33240,N_30696,N_30867);
or U33241 (N_33241,N_31709,N_30385);
xor U33242 (N_33242,N_30192,N_30508);
xor U33243 (N_33243,N_30847,N_31663);
or U33244 (N_33244,N_30878,N_30572);
or U33245 (N_33245,N_30278,N_30221);
nor U33246 (N_33246,N_31499,N_31476);
xor U33247 (N_33247,N_31377,N_30224);
nor U33248 (N_33248,N_30612,N_30383);
xor U33249 (N_33249,N_30905,N_31833);
or U33250 (N_33250,N_30614,N_31344);
nand U33251 (N_33251,N_31076,N_31366);
and U33252 (N_33252,N_30352,N_30744);
nand U33253 (N_33253,N_31223,N_30619);
or U33254 (N_33254,N_31426,N_31493);
and U33255 (N_33255,N_31909,N_30951);
nand U33256 (N_33256,N_30013,N_30791);
nor U33257 (N_33257,N_31438,N_30651);
nand U33258 (N_33258,N_30941,N_30121);
xnor U33259 (N_33259,N_30018,N_30211);
nand U33260 (N_33260,N_31011,N_30719);
xor U33261 (N_33261,N_31185,N_31065);
and U33262 (N_33262,N_31384,N_31130);
xor U33263 (N_33263,N_31682,N_31051);
and U33264 (N_33264,N_30727,N_30919);
nand U33265 (N_33265,N_31013,N_30140);
xnor U33266 (N_33266,N_31952,N_31382);
nor U33267 (N_33267,N_30794,N_31222);
and U33268 (N_33268,N_31121,N_31687);
and U33269 (N_33269,N_31383,N_30119);
nor U33270 (N_33270,N_31489,N_30681);
and U33271 (N_33271,N_31555,N_30434);
or U33272 (N_33272,N_30716,N_30011);
or U33273 (N_33273,N_31420,N_31011);
nand U33274 (N_33274,N_30089,N_31100);
or U33275 (N_33275,N_31032,N_31547);
and U33276 (N_33276,N_31225,N_30870);
or U33277 (N_33277,N_31278,N_31483);
nand U33278 (N_33278,N_31689,N_31167);
and U33279 (N_33279,N_30173,N_30673);
nor U33280 (N_33280,N_30034,N_31521);
xor U33281 (N_33281,N_31434,N_30369);
or U33282 (N_33282,N_31365,N_31518);
or U33283 (N_33283,N_31300,N_31307);
nor U33284 (N_33284,N_30400,N_30736);
nor U33285 (N_33285,N_30148,N_31068);
nor U33286 (N_33286,N_30596,N_31983);
nand U33287 (N_33287,N_31859,N_30706);
and U33288 (N_33288,N_30470,N_30966);
nor U33289 (N_33289,N_31956,N_31275);
nand U33290 (N_33290,N_31944,N_31395);
nor U33291 (N_33291,N_30347,N_31371);
nand U33292 (N_33292,N_31453,N_30933);
nand U33293 (N_33293,N_30387,N_30647);
nand U33294 (N_33294,N_31525,N_30924);
or U33295 (N_33295,N_31049,N_30828);
nand U33296 (N_33296,N_30382,N_31236);
nor U33297 (N_33297,N_30723,N_31662);
and U33298 (N_33298,N_30514,N_31050);
nand U33299 (N_33299,N_30663,N_30825);
xnor U33300 (N_33300,N_30579,N_30680);
nor U33301 (N_33301,N_30308,N_30409);
nor U33302 (N_33302,N_30474,N_30791);
and U33303 (N_33303,N_30493,N_31432);
nand U33304 (N_33304,N_31925,N_30760);
xor U33305 (N_33305,N_30598,N_31367);
or U33306 (N_33306,N_31191,N_31319);
nor U33307 (N_33307,N_30398,N_31320);
or U33308 (N_33308,N_31228,N_30829);
or U33309 (N_33309,N_30005,N_30881);
nand U33310 (N_33310,N_30644,N_30220);
xor U33311 (N_33311,N_31672,N_31915);
nor U33312 (N_33312,N_31938,N_30975);
and U33313 (N_33313,N_30788,N_31758);
xnor U33314 (N_33314,N_31792,N_30218);
nor U33315 (N_33315,N_30387,N_30814);
nor U33316 (N_33316,N_30963,N_31421);
nor U33317 (N_33317,N_30852,N_30578);
or U33318 (N_33318,N_30268,N_31336);
nor U33319 (N_33319,N_30757,N_30335);
or U33320 (N_33320,N_31827,N_31163);
nand U33321 (N_33321,N_30535,N_31241);
and U33322 (N_33322,N_31787,N_30416);
or U33323 (N_33323,N_30826,N_30169);
or U33324 (N_33324,N_30572,N_30425);
nor U33325 (N_33325,N_31271,N_31127);
nor U33326 (N_33326,N_30272,N_31304);
nand U33327 (N_33327,N_31790,N_31709);
xor U33328 (N_33328,N_31826,N_31032);
or U33329 (N_33329,N_30523,N_30663);
nor U33330 (N_33330,N_30301,N_30250);
xnor U33331 (N_33331,N_30755,N_31731);
nand U33332 (N_33332,N_30959,N_31656);
or U33333 (N_33333,N_30747,N_31334);
nand U33334 (N_33334,N_31088,N_30043);
and U33335 (N_33335,N_31332,N_31830);
nor U33336 (N_33336,N_31414,N_31534);
and U33337 (N_33337,N_31512,N_30194);
nor U33338 (N_33338,N_31509,N_30197);
or U33339 (N_33339,N_31564,N_31749);
or U33340 (N_33340,N_31278,N_30227);
nand U33341 (N_33341,N_31392,N_31914);
or U33342 (N_33342,N_30580,N_30287);
or U33343 (N_33343,N_30466,N_31865);
nor U33344 (N_33344,N_31150,N_30169);
or U33345 (N_33345,N_31200,N_31563);
or U33346 (N_33346,N_30129,N_30607);
or U33347 (N_33347,N_30597,N_31248);
and U33348 (N_33348,N_30604,N_30281);
xor U33349 (N_33349,N_31422,N_30989);
or U33350 (N_33350,N_30950,N_30898);
nor U33351 (N_33351,N_31546,N_30892);
nor U33352 (N_33352,N_30779,N_31455);
or U33353 (N_33353,N_30837,N_31137);
nand U33354 (N_33354,N_31038,N_31171);
xor U33355 (N_33355,N_31790,N_30386);
or U33356 (N_33356,N_31096,N_31969);
nor U33357 (N_33357,N_30502,N_30557);
nor U33358 (N_33358,N_31665,N_30464);
nor U33359 (N_33359,N_31498,N_31381);
nand U33360 (N_33360,N_30491,N_31593);
xor U33361 (N_33361,N_31594,N_30261);
or U33362 (N_33362,N_30577,N_30317);
xor U33363 (N_33363,N_31484,N_31784);
nand U33364 (N_33364,N_31131,N_30293);
and U33365 (N_33365,N_31201,N_30987);
nand U33366 (N_33366,N_31455,N_30915);
and U33367 (N_33367,N_31346,N_30122);
nor U33368 (N_33368,N_31026,N_31495);
and U33369 (N_33369,N_30961,N_31829);
or U33370 (N_33370,N_30195,N_31773);
nand U33371 (N_33371,N_31819,N_30014);
or U33372 (N_33372,N_30593,N_30421);
or U33373 (N_33373,N_31571,N_30717);
and U33374 (N_33374,N_31631,N_30851);
xor U33375 (N_33375,N_31422,N_30408);
xnor U33376 (N_33376,N_31958,N_30745);
or U33377 (N_33377,N_31218,N_30038);
or U33378 (N_33378,N_30268,N_31712);
or U33379 (N_33379,N_31862,N_30896);
or U33380 (N_33380,N_31017,N_31514);
or U33381 (N_33381,N_31469,N_31466);
nor U33382 (N_33382,N_31285,N_31027);
and U33383 (N_33383,N_30759,N_30846);
xor U33384 (N_33384,N_31046,N_30080);
xor U33385 (N_33385,N_31539,N_31529);
and U33386 (N_33386,N_31391,N_30218);
or U33387 (N_33387,N_30448,N_31033);
xor U33388 (N_33388,N_31858,N_30800);
or U33389 (N_33389,N_31987,N_31184);
nand U33390 (N_33390,N_30750,N_31570);
or U33391 (N_33391,N_31980,N_31401);
xor U33392 (N_33392,N_31394,N_30615);
xnor U33393 (N_33393,N_31360,N_31452);
xor U33394 (N_33394,N_30236,N_31063);
nand U33395 (N_33395,N_30943,N_31376);
nand U33396 (N_33396,N_30639,N_30545);
or U33397 (N_33397,N_31325,N_31274);
or U33398 (N_33398,N_30612,N_31477);
nor U33399 (N_33399,N_31995,N_30155);
and U33400 (N_33400,N_30412,N_30377);
nand U33401 (N_33401,N_30517,N_30441);
and U33402 (N_33402,N_31544,N_30069);
or U33403 (N_33403,N_31745,N_31730);
nand U33404 (N_33404,N_30617,N_31410);
and U33405 (N_33405,N_31143,N_30557);
xnor U33406 (N_33406,N_31132,N_30046);
and U33407 (N_33407,N_30256,N_30235);
or U33408 (N_33408,N_30299,N_30101);
nor U33409 (N_33409,N_30573,N_30873);
nand U33410 (N_33410,N_30878,N_31363);
xor U33411 (N_33411,N_31461,N_31023);
and U33412 (N_33412,N_30082,N_31666);
nor U33413 (N_33413,N_30941,N_30069);
and U33414 (N_33414,N_30058,N_30878);
xnor U33415 (N_33415,N_30702,N_30706);
or U33416 (N_33416,N_30049,N_30174);
and U33417 (N_33417,N_30019,N_30664);
or U33418 (N_33418,N_30282,N_31759);
xor U33419 (N_33419,N_31954,N_31426);
or U33420 (N_33420,N_30858,N_31940);
xor U33421 (N_33421,N_31950,N_30397);
or U33422 (N_33422,N_31613,N_31358);
or U33423 (N_33423,N_31529,N_30881);
or U33424 (N_33424,N_30135,N_31216);
xnor U33425 (N_33425,N_31744,N_30822);
nand U33426 (N_33426,N_31602,N_31361);
and U33427 (N_33427,N_30544,N_31049);
nand U33428 (N_33428,N_31311,N_31075);
nor U33429 (N_33429,N_31306,N_30035);
nand U33430 (N_33430,N_30505,N_30676);
xor U33431 (N_33431,N_30921,N_30432);
xor U33432 (N_33432,N_31156,N_30064);
and U33433 (N_33433,N_31772,N_30190);
or U33434 (N_33434,N_30030,N_30762);
nor U33435 (N_33435,N_31219,N_31755);
or U33436 (N_33436,N_30344,N_31094);
nand U33437 (N_33437,N_31015,N_31571);
or U33438 (N_33438,N_30283,N_30429);
nor U33439 (N_33439,N_31399,N_30254);
nand U33440 (N_33440,N_30624,N_31098);
or U33441 (N_33441,N_30352,N_31262);
nand U33442 (N_33442,N_30903,N_30815);
and U33443 (N_33443,N_30303,N_31872);
nand U33444 (N_33444,N_30498,N_30893);
nand U33445 (N_33445,N_30602,N_31134);
nand U33446 (N_33446,N_30491,N_30313);
nand U33447 (N_33447,N_31908,N_31887);
or U33448 (N_33448,N_31476,N_30905);
nor U33449 (N_33449,N_30230,N_31630);
and U33450 (N_33450,N_31160,N_31962);
or U33451 (N_33451,N_30916,N_30032);
nand U33452 (N_33452,N_30721,N_31843);
nor U33453 (N_33453,N_30856,N_31165);
xor U33454 (N_33454,N_31660,N_30090);
nor U33455 (N_33455,N_31707,N_31087);
nand U33456 (N_33456,N_30606,N_31266);
xor U33457 (N_33457,N_30815,N_30897);
nor U33458 (N_33458,N_31806,N_30604);
and U33459 (N_33459,N_30981,N_31829);
nor U33460 (N_33460,N_30483,N_31603);
xor U33461 (N_33461,N_31286,N_30880);
nor U33462 (N_33462,N_31457,N_30315);
and U33463 (N_33463,N_30243,N_30848);
nand U33464 (N_33464,N_31416,N_31392);
nor U33465 (N_33465,N_30923,N_31634);
or U33466 (N_33466,N_30835,N_31892);
xor U33467 (N_33467,N_30933,N_31937);
nor U33468 (N_33468,N_31364,N_30290);
nand U33469 (N_33469,N_30194,N_30760);
nand U33470 (N_33470,N_31145,N_31013);
nor U33471 (N_33471,N_30554,N_30874);
nand U33472 (N_33472,N_31860,N_31968);
nor U33473 (N_33473,N_31165,N_30690);
or U33474 (N_33474,N_30773,N_31602);
nand U33475 (N_33475,N_31266,N_31681);
nor U33476 (N_33476,N_30678,N_30496);
or U33477 (N_33477,N_31589,N_30026);
or U33478 (N_33478,N_30820,N_31984);
nor U33479 (N_33479,N_30258,N_30091);
nand U33480 (N_33480,N_30169,N_31673);
or U33481 (N_33481,N_31200,N_30724);
nand U33482 (N_33482,N_30598,N_31921);
xor U33483 (N_33483,N_30602,N_30385);
nor U33484 (N_33484,N_31043,N_31478);
and U33485 (N_33485,N_30534,N_31516);
xor U33486 (N_33486,N_30779,N_30585);
xor U33487 (N_33487,N_31002,N_30772);
nor U33488 (N_33488,N_30183,N_30820);
xnor U33489 (N_33489,N_30360,N_30162);
nor U33490 (N_33490,N_30004,N_31016);
xor U33491 (N_33491,N_30573,N_30482);
nand U33492 (N_33492,N_30594,N_30577);
nand U33493 (N_33493,N_30546,N_31827);
or U33494 (N_33494,N_31503,N_30218);
nor U33495 (N_33495,N_30201,N_31760);
xor U33496 (N_33496,N_30695,N_30924);
xor U33497 (N_33497,N_31584,N_30486);
nand U33498 (N_33498,N_30511,N_30733);
xor U33499 (N_33499,N_30094,N_31088);
nand U33500 (N_33500,N_31617,N_31952);
xor U33501 (N_33501,N_31169,N_31890);
xor U33502 (N_33502,N_30597,N_30655);
or U33503 (N_33503,N_30410,N_30147);
and U33504 (N_33504,N_30380,N_31235);
or U33505 (N_33505,N_31457,N_31694);
nor U33506 (N_33506,N_31618,N_30473);
nor U33507 (N_33507,N_31629,N_30333);
xnor U33508 (N_33508,N_30176,N_30825);
or U33509 (N_33509,N_30498,N_30980);
xor U33510 (N_33510,N_30065,N_30338);
nor U33511 (N_33511,N_30816,N_30184);
xor U33512 (N_33512,N_31570,N_30399);
or U33513 (N_33513,N_30054,N_30953);
or U33514 (N_33514,N_30836,N_31940);
nand U33515 (N_33515,N_31939,N_31553);
xor U33516 (N_33516,N_31997,N_30607);
nand U33517 (N_33517,N_31569,N_30455);
xor U33518 (N_33518,N_30838,N_31614);
xnor U33519 (N_33519,N_30038,N_30155);
or U33520 (N_33520,N_31311,N_30528);
nor U33521 (N_33521,N_30918,N_30247);
nor U33522 (N_33522,N_30365,N_31203);
and U33523 (N_33523,N_31613,N_30975);
and U33524 (N_33524,N_30600,N_31690);
nor U33525 (N_33525,N_31171,N_31767);
nor U33526 (N_33526,N_30395,N_30757);
xor U33527 (N_33527,N_31125,N_31563);
and U33528 (N_33528,N_31527,N_30882);
xnor U33529 (N_33529,N_30499,N_30187);
and U33530 (N_33530,N_30616,N_30816);
xor U33531 (N_33531,N_31427,N_31000);
xor U33532 (N_33532,N_30126,N_30163);
nor U33533 (N_33533,N_30965,N_30536);
and U33534 (N_33534,N_31922,N_31214);
xor U33535 (N_33535,N_30183,N_31125);
nand U33536 (N_33536,N_31443,N_31793);
or U33537 (N_33537,N_31067,N_30777);
xnor U33538 (N_33538,N_30664,N_30018);
and U33539 (N_33539,N_30547,N_30721);
nand U33540 (N_33540,N_30017,N_31409);
xnor U33541 (N_33541,N_30748,N_31496);
nand U33542 (N_33542,N_30613,N_31831);
nand U33543 (N_33543,N_30920,N_31220);
or U33544 (N_33544,N_31760,N_30130);
nor U33545 (N_33545,N_30969,N_30314);
nor U33546 (N_33546,N_31057,N_30150);
nand U33547 (N_33547,N_30728,N_30767);
or U33548 (N_33548,N_30090,N_30392);
or U33549 (N_33549,N_31007,N_30158);
or U33550 (N_33550,N_30364,N_31551);
nand U33551 (N_33551,N_31820,N_30999);
or U33552 (N_33552,N_30306,N_31084);
and U33553 (N_33553,N_31612,N_31797);
nor U33554 (N_33554,N_31660,N_30182);
xnor U33555 (N_33555,N_31864,N_31193);
nor U33556 (N_33556,N_31726,N_31124);
and U33557 (N_33557,N_31214,N_31403);
nor U33558 (N_33558,N_31640,N_30627);
nor U33559 (N_33559,N_30869,N_31577);
or U33560 (N_33560,N_31401,N_30513);
xnor U33561 (N_33561,N_31935,N_30905);
and U33562 (N_33562,N_31633,N_31555);
nor U33563 (N_33563,N_31796,N_31289);
nor U33564 (N_33564,N_30605,N_31812);
nand U33565 (N_33565,N_31871,N_31960);
or U33566 (N_33566,N_30577,N_31657);
nand U33567 (N_33567,N_31292,N_31402);
nand U33568 (N_33568,N_31071,N_31885);
nor U33569 (N_33569,N_31966,N_31909);
and U33570 (N_33570,N_31018,N_31973);
nand U33571 (N_33571,N_30247,N_30745);
nor U33572 (N_33572,N_30453,N_30906);
nand U33573 (N_33573,N_31772,N_30105);
nand U33574 (N_33574,N_30251,N_30517);
and U33575 (N_33575,N_31961,N_31803);
nand U33576 (N_33576,N_30101,N_31388);
or U33577 (N_33577,N_30665,N_30854);
or U33578 (N_33578,N_30798,N_31963);
nor U33579 (N_33579,N_30477,N_30659);
or U33580 (N_33580,N_30554,N_31833);
and U33581 (N_33581,N_30243,N_31805);
or U33582 (N_33582,N_30067,N_30763);
xor U33583 (N_33583,N_31010,N_31809);
xor U33584 (N_33584,N_31321,N_31840);
nand U33585 (N_33585,N_31691,N_31346);
nor U33586 (N_33586,N_30343,N_31754);
or U33587 (N_33587,N_31695,N_30481);
nand U33588 (N_33588,N_31659,N_30332);
xor U33589 (N_33589,N_31819,N_30577);
nand U33590 (N_33590,N_31356,N_30260);
and U33591 (N_33591,N_30602,N_31581);
or U33592 (N_33592,N_31604,N_31307);
nand U33593 (N_33593,N_31046,N_31121);
nor U33594 (N_33594,N_30357,N_30879);
or U33595 (N_33595,N_31541,N_30762);
and U33596 (N_33596,N_30719,N_30338);
or U33597 (N_33597,N_30408,N_31571);
nand U33598 (N_33598,N_31206,N_30777);
and U33599 (N_33599,N_31741,N_31556);
nand U33600 (N_33600,N_30210,N_31622);
nor U33601 (N_33601,N_31467,N_30200);
xnor U33602 (N_33602,N_31814,N_31007);
and U33603 (N_33603,N_30851,N_30051);
xor U33604 (N_33604,N_30322,N_31991);
and U33605 (N_33605,N_31192,N_31464);
and U33606 (N_33606,N_31795,N_30677);
or U33607 (N_33607,N_31358,N_31435);
and U33608 (N_33608,N_30570,N_30281);
nand U33609 (N_33609,N_30723,N_30868);
or U33610 (N_33610,N_30334,N_31910);
xor U33611 (N_33611,N_30683,N_31345);
nand U33612 (N_33612,N_31572,N_30775);
xor U33613 (N_33613,N_31696,N_31941);
or U33614 (N_33614,N_31593,N_30700);
and U33615 (N_33615,N_30570,N_30416);
nand U33616 (N_33616,N_30568,N_30766);
nand U33617 (N_33617,N_31215,N_30106);
xnor U33618 (N_33618,N_31360,N_31138);
xnor U33619 (N_33619,N_30861,N_31705);
and U33620 (N_33620,N_31985,N_30620);
nor U33621 (N_33621,N_31640,N_31487);
and U33622 (N_33622,N_31832,N_30740);
or U33623 (N_33623,N_30486,N_30420);
and U33624 (N_33624,N_31706,N_31884);
xnor U33625 (N_33625,N_31557,N_31954);
and U33626 (N_33626,N_31158,N_31746);
nor U33627 (N_33627,N_31169,N_31535);
nand U33628 (N_33628,N_30201,N_31883);
nor U33629 (N_33629,N_31700,N_31005);
nand U33630 (N_33630,N_30228,N_30912);
and U33631 (N_33631,N_30492,N_30773);
nor U33632 (N_33632,N_31197,N_30795);
or U33633 (N_33633,N_31655,N_30293);
nand U33634 (N_33634,N_30423,N_30848);
or U33635 (N_33635,N_31409,N_31206);
and U33636 (N_33636,N_31482,N_31147);
or U33637 (N_33637,N_31232,N_31753);
and U33638 (N_33638,N_31747,N_31311);
or U33639 (N_33639,N_31716,N_31936);
and U33640 (N_33640,N_31372,N_31746);
nand U33641 (N_33641,N_31445,N_30036);
and U33642 (N_33642,N_30177,N_31408);
nor U33643 (N_33643,N_30318,N_31981);
nor U33644 (N_33644,N_30926,N_31098);
nand U33645 (N_33645,N_30926,N_31316);
xnor U33646 (N_33646,N_31634,N_31285);
and U33647 (N_33647,N_30408,N_30342);
nor U33648 (N_33648,N_30220,N_31891);
or U33649 (N_33649,N_31926,N_31639);
or U33650 (N_33650,N_31912,N_31895);
xnor U33651 (N_33651,N_30269,N_30276);
xnor U33652 (N_33652,N_31273,N_31655);
xor U33653 (N_33653,N_30712,N_30053);
nor U33654 (N_33654,N_30136,N_30757);
xor U33655 (N_33655,N_31259,N_31566);
xnor U33656 (N_33656,N_30937,N_31367);
and U33657 (N_33657,N_31450,N_30942);
nand U33658 (N_33658,N_30470,N_30282);
and U33659 (N_33659,N_30110,N_31257);
or U33660 (N_33660,N_30056,N_31344);
and U33661 (N_33661,N_30717,N_30425);
xor U33662 (N_33662,N_30987,N_31554);
xor U33663 (N_33663,N_30075,N_30998);
or U33664 (N_33664,N_31344,N_31095);
or U33665 (N_33665,N_31457,N_31508);
nand U33666 (N_33666,N_31983,N_31918);
or U33667 (N_33667,N_30404,N_30737);
and U33668 (N_33668,N_31918,N_30927);
nand U33669 (N_33669,N_31018,N_31488);
nand U33670 (N_33670,N_30196,N_30588);
xnor U33671 (N_33671,N_30277,N_31233);
xnor U33672 (N_33672,N_31202,N_30826);
and U33673 (N_33673,N_31923,N_30502);
and U33674 (N_33674,N_31669,N_31721);
nand U33675 (N_33675,N_31079,N_30899);
nor U33676 (N_33676,N_30399,N_31198);
or U33677 (N_33677,N_31626,N_30018);
nor U33678 (N_33678,N_30131,N_31626);
nor U33679 (N_33679,N_30505,N_31645);
xnor U33680 (N_33680,N_30044,N_31386);
nor U33681 (N_33681,N_30426,N_30080);
nor U33682 (N_33682,N_31554,N_30626);
nand U33683 (N_33683,N_31936,N_30285);
or U33684 (N_33684,N_31870,N_31184);
xnor U33685 (N_33685,N_31457,N_31093);
nand U33686 (N_33686,N_30474,N_31866);
xor U33687 (N_33687,N_30799,N_31586);
and U33688 (N_33688,N_31650,N_31116);
or U33689 (N_33689,N_30274,N_30962);
and U33690 (N_33690,N_30092,N_31371);
nor U33691 (N_33691,N_31272,N_31842);
nor U33692 (N_33692,N_31321,N_30143);
xnor U33693 (N_33693,N_30382,N_31403);
nor U33694 (N_33694,N_31456,N_30934);
nand U33695 (N_33695,N_31019,N_30514);
xor U33696 (N_33696,N_30741,N_31045);
xor U33697 (N_33697,N_31537,N_31858);
xor U33698 (N_33698,N_31791,N_31919);
xnor U33699 (N_33699,N_30676,N_30711);
xnor U33700 (N_33700,N_30987,N_30048);
nand U33701 (N_33701,N_31112,N_31793);
xor U33702 (N_33702,N_31460,N_30185);
or U33703 (N_33703,N_30183,N_30406);
and U33704 (N_33704,N_30147,N_31054);
or U33705 (N_33705,N_30681,N_31652);
and U33706 (N_33706,N_31741,N_30299);
and U33707 (N_33707,N_31542,N_30828);
and U33708 (N_33708,N_31533,N_30641);
or U33709 (N_33709,N_30253,N_30652);
xnor U33710 (N_33710,N_31014,N_31767);
and U33711 (N_33711,N_31488,N_30291);
nor U33712 (N_33712,N_31187,N_30353);
nand U33713 (N_33713,N_31982,N_30434);
xor U33714 (N_33714,N_30751,N_30905);
xor U33715 (N_33715,N_30757,N_30123);
or U33716 (N_33716,N_30546,N_31144);
nand U33717 (N_33717,N_31676,N_30082);
and U33718 (N_33718,N_31893,N_30430);
nand U33719 (N_33719,N_31940,N_31123);
and U33720 (N_33720,N_30820,N_30455);
nand U33721 (N_33721,N_30230,N_31315);
or U33722 (N_33722,N_31340,N_30418);
nor U33723 (N_33723,N_31197,N_30824);
xnor U33724 (N_33724,N_30807,N_30689);
nand U33725 (N_33725,N_30583,N_30542);
nand U33726 (N_33726,N_30889,N_30606);
or U33727 (N_33727,N_31589,N_31674);
or U33728 (N_33728,N_30633,N_30066);
and U33729 (N_33729,N_30375,N_30855);
and U33730 (N_33730,N_31034,N_31705);
xnor U33731 (N_33731,N_31873,N_30504);
xor U33732 (N_33732,N_30363,N_30458);
nand U33733 (N_33733,N_31688,N_31024);
or U33734 (N_33734,N_31974,N_31843);
or U33735 (N_33735,N_31342,N_31501);
xor U33736 (N_33736,N_30227,N_31043);
nand U33737 (N_33737,N_31737,N_31953);
xnor U33738 (N_33738,N_30749,N_31815);
nand U33739 (N_33739,N_31363,N_31472);
nor U33740 (N_33740,N_30283,N_31691);
xor U33741 (N_33741,N_31538,N_30941);
and U33742 (N_33742,N_31569,N_31121);
or U33743 (N_33743,N_30493,N_31584);
nand U33744 (N_33744,N_31562,N_30181);
or U33745 (N_33745,N_31074,N_30467);
xor U33746 (N_33746,N_30923,N_30430);
and U33747 (N_33747,N_30748,N_31567);
and U33748 (N_33748,N_31800,N_31034);
nor U33749 (N_33749,N_30058,N_30039);
xnor U33750 (N_33750,N_31575,N_30794);
nor U33751 (N_33751,N_31241,N_31528);
or U33752 (N_33752,N_31347,N_30446);
and U33753 (N_33753,N_30323,N_30855);
xor U33754 (N_33754,N_31052,N_30646);
xnor U33755 (N_33755,N_30208,N_31330);
nor U33756 (N_33756,N_31419,N_30264);
xnor U33757 (N_33757,N_31511,N_31171);
xor U33758 (N_33758,N_31524,N_30810);
nand U33759 (N_33759,N_30333,N_31673);
or U33760 (N_33760,N_31908,N_31350);
nor U33761 (N_33761,N_31804,N_30380);
or U33762 (N_33762,N_31418,N_30761);
nand U33763 (N_33763,N_30467,N_31103);
and U33764 (N_33764,N_31494,N_30128);
xor U33765 (N_33765,N_30423,N_31101);
xnor U33766 (N_33766,N_31977,N_31998);
xnor U33767 (N_33767,N_30983,N_31298);
xor U33768 (N_33768,N_30439,N_30758);
nor U33769 (N_33769,N_30765,N_30505);
or U33770 (N_33770,N_31845,N_31208);
nor U33771 (N_33771,N_30358,N_30804);
nor U33772 (N_33772,N_30452,N_30039);
xor U33773 (N_33773,N_31968,N_30426);
and U33774 (N_33774,N_30543,N_30830);
nor U33775 (N_33775,N_31779,N_31964);
nor U33776 (N_33776,N_30476,N_31412);
and U33777 (N_33777,N_30434,N_30630);
and U33778 (N_33778,N_30233,N_31525);
or U33779 (N_33779,N_31319,N_31251);
nor U33780 (N_33780,N_31090,N_31420);
nor U33781 (N_33781,N_31221,N_31466);
or U33782 (N_33782,N_30693,N_30229);
nand U33783 (N_33783,N_31496,N_30079);
xnor U33784 (N_33784,N_31233,N_31140);
or U33785 (N_33785,N_30882,N_30865);
xor U33786 (N_33786,N_31660,N_30826);
xor U33787 (N_33787,N_30098,N_30023);
or U33788 (N_33788,N_30360,N_30717);
xnor U33789 (N_33789,N_31818,N_31237);
nand U33790 (N_33790,N_30427,N_31742);
nor U33791 (N_33791,N_31346,N_30191);
nand U33792 (N_33792,N_30942,N_30221);
xor U33793 (N_33793,N_30008,N_31184);
and U33794 (N_33794,N_30489,N_31501);
xor U33795 (N_33795,N_31920,N_31461);
or U33796 (N_33796,N_31978,N_30831);
xnor U33797 (N_33797,N_31559,N_30387);
nor U33798 (N_33798,N_30478,N_30857);
nor U33799 (N_33799,N_30044,N_30550);
or U33800 (N_33800,N_31546,N_30072);
xor U33801 (N_33801,N_30574,N_31644);
and U33802 (N_33802,N_30299,N_30053);
or U33803 (N_33803,N_30793,N_30527);
xnor U33804 (N_33804,N_30155,N_31918);
or U33805 (N_33805,N_30564,N_31802);
or U33806 (N_33806,N_30584,N_30535);
and U33807 (N_33807,N_30153,N_30468);
and U33808 (N_33808,N_30215,N_31034);
and U33809 (N_33809,N_31161,N_30849);
nor U33810 (N_33810,N_30111,N_31098);
nor U33811 (N_33811,N_31863,N_31554);
nand U33812 (N_33812,N_30390,N_31066);
xnor U33813 (N_33813,N_31158,N_31284);
or U33814 (N_33814,N_30274,N_30319);
nand U33815 (N_33815,N_30930,N_30320);
or U33816 (N_33816,N_30506,N_31868);
nand U33817 (N_33817,N_30623,N_30761);
or U33818 (N_33818,N_30010,N_31121);
and U33819 (N_33819,N_31059,N_31728);
and U33820 (N_33820,N_31898,N_30610);
and U33821 (N_33821,N_31593,N_31995);
xnor U33822 (N_33822,N_30887,N_31997);
xor U33823 (N_33823,N_31477,N_30698);
or U33824 (N_33824,N_30756,N_30456);
nor U33825 (N_33825,N_31805,N_31644);
nand U33826 (N_33826,N_31029,N_30919);
nand U33827 (N_33827,N_30463,N_31451);
xnor U33828 (N_33828,N_31464,N_30467);
xor U33829 (N_33829,N_30605,N_31054);
and U33830 (N_33830,N_30494,N_30096);
or U33831 (N_33831,N_31274,N_31864);
xnor U33832 (N_33832,N_30287,N_30943);
nor U33833 (N_33833,N_30573,N_31980);
xor U33834 (N_33834,N_31131,N_30161);
nor U33835 (N_33835,N_30303,N_30469);
nand U33836 (N_33836,N_31154,N_30031);
or U33837 (N_33837,N_31948,N_31774);
or U33838 (N_33838,N_30479,N_31282);
nand U33839 (N_33839,N_31462,N_31455);
or U33840 (N_33840,N_31478,N_30078);
and U33841 (N_33841,N_30417,N_30089);
nor U33842 (N_33842,N_31540,N_30204);
and U33843 (N_33843,N_31440,N_31616);
nand U33844 (N_33844,N_30907,N_30226);
nand U33845 (N_33845,N_31656,N_30099);
nand U33846 (N_33846,N_30236,N_31756);
or U33847 (N_33847,N_31925,N_30387);
nor U33848 (N_33848,N_30458,N_30560);
and U33849 (N_33849,N_31132,N_30275);
nor U33850 (N_33850,N_31805,N_31538);
and U33851 (N_33851,N_30151,N_30855);
or U33852 (N_33852,N_30998,N_31662);
xor U33853 (N_33853,N_30709,N_31199);
xnor U33854 (N_33854,N_31924,N_31164);
xnor U33855 (N_33855,N_31907,N_31159);
and U33856 (N_33856,N_31269,N_31490);
nand U33857 (N_33857,N_31557,N_31689);
nor U33858 (N_33858,N_30846,N_31335);
or U33859 (N_33859,N_30370,N_30921);
xor U33860 (N_33860,N_31240,N_31043);
or U33861 (N_33861,N_30733,N_31401);
or U33862 (N_33862,N_30445,N_31445);
or U33863 (N_33863,N_30971,N_31251);
or U33864 (N_33864,N_30888,N_30165);
nand U33865 (N_33865,N_30232,N_31360);
or U33866 (N_33866,N_31764,N_30407);
or U33867 (N_33867,N_31490,N_30448);
and U33868 (N_33868,N_30785,N_31024);
xnor U33869 (N_33869,N_31693,N_30261);
xor U33870 (N_33870,N_31633,N_31495);
nand U33871 (N_33871,N_30371,N_30189);
or U33872 (N_33872,N_30304,N_30198);
nor U33873 (N_33873,N_30902,N_30586);
and U33874 (N_33874,N_30329,N_30962);
and U33875 (N_33875,N_31810,N_30320);
or U33876 (N_33876,N_30112,N_30017);
or U33877 (N_33877,N_31408,N_30347);
or U33878 (N_33878,N_30762,N_30247);
or U33879 (N_33879,N_31354,N_30659);
nand U33880 (N_33880,N_30641,N_31017);
or U33881 (N_33881,N_31742,N_31760);
or U33882 (N_33882,N_30965,N_30973);
nand U33883 (N_33883,N_30145,N_31571);
xor U33884 (N_33884,N_31159,N_31013);
xnor U33885 (N_33885,N_30697,N_30220);
nand U33886 (N_33886,N_31863,N_31103);
or U33887 (N_33887,N_31548,N_31259);
and U33888 (N_33888,N_30701,N_30960);
and U33889 (N_33889,N_30158,N_30875);
nand U33890 (N_33890,N_31768,N_30561);
nor U33891 (N_33891,N_30817,N_30144);
xnor U33892 (N_33892,N_31449,N_30172);
nand U33893 (N_33893,N_30503,N_31641);
nand U33894 (N_33894,N_31806,N_31813);
xnor U33895 (N_33895,N_30618,N_31309);
or U33896 (N_33896,N_30594,N_30248);
and U33897 (N_33897,N_30570,N_30237);
and U33898 (N_33898,N_31541,N_30910);
nor U33899 (N_33899,N_30683,N_30419);
or U33900 (N_33900,N_31919,N_31594);
and U33901 (N_33901,N_31454,N_30692);
or U33902 (N_33902,N_30571,N_30881);
or U33903 (N_33903,N_31772,N_31752);
or U33904 (N_33904,N_30147,N_30753);
or U33905 (N_33905,N_31184,N_30062);
and U33906 (N_33906,N_31510,N_31378);
or U33907 (N_33907,N_31589,N_30731);
xnor U33908 (N_33908,N_31997,N_31080);
and U33909 (N_33909,N_31645,N_30192);
xor U33910 (N_33910,N_30649,N_30479);
nand U33911 (N_33911,N_31674,N_31614);
or U33912 (N_33912,N_31454,N_30320);
xnor U33913 (N_33913,N_31544,N_31277);
or U33914 (N_33914,N_31203,N_31284);
and U33915 (N_33915,N_30914,N_31850);
or U33916 (N_33916,N_31879,N_30855);
or U33917 (N_33917,N_30093,N_31511);
nor U33918 (N_33918,N_31384,N_30728);
or U33919 (N_33919,N_31481,N_31931);
nor U33920 (N_33920,N_30420,N_30525);
nand U33921 (N_33921,N_31551,N_31174);
and U33922 (N_33922,N_31408,N_30237);
nand U33923 (N_33923,N_30240,N_31068);
or U33924 (N_33924,N_31952,N_31506);
xnor U33925 (N_33925,N_30166,N_31598);
or U33926 (N_33926,N_30124,N_30543);
xnor U33927 (N_33927,N_31713,N_30636);
nand U33928 (N_33928,N_30587,N_31955);
and U33929 (N_33929,N_30033,N_31387);
nor U33930 (N_33930,N_31895,N_31409);
nand U33931 (N_33931,N_31506,N_31437);
nand U33932 (N_33932,N_30071,N_31862);
xor U33933 (N_33933,N_31106,N_30776);
xnor U33934 (N_33934,N_31040,N_30701);
and U33935 (N_33935,N_30150,N_30754);
or U33936 (N_33936,N_31631,N_30162);
nand U33937 (N_33937,N_30437,N_31968);
and U33938 (N_33938,N_30439,N_30959);
or U33939 (N_33939,N_30349,N_31532);
and U33940 (N_33940,N_31565,N_31087);
or U33941 (N_33941,N_30001,N_30712);
nor U33942 (N_33942,N_30791,N_30837);
and U33943 (N_33943,N_31376,N_30228);
nor U33944 (N_33944,N_30061,N_31379);
nand U33945 (N_33945,N_31925,N_30042);
nand U33946 (N_33946,N_30658,N_31434);
xnor U33947 (N_33947,N_30584,N_30572);
nand U33948 (N_33948,N_31983,N_31895);
xor U33949 (N_33949,N_31157,N_30575);
xor U33950 (N_33950,N_31182,N_30115);
and U33951 (N_33951,N_30072,N_31893);
nor U33952 (N_33952,N_30131,N_31012);
nor U33953 (N_33953,N_31173,N_31698);
or U33954 (N_33954,N_31978,N_30434);
or U33955 (N_33955,N_31375,N_30236);
nand U33956 (N_33956,N_31455,N_30931);
nor U33957 (N_33957,N_30700,N_30713);
xnor U33958 (N_33958,N_30934,N_31069);
and U33959 (N_33959,N_30637,N_30025);
xnor U33960 (N_33960,N_30981,N_30768);
xor U33961 (N_33961,N_31118,N_31079);
xor U33962 (N_33962,N_31030,N_30470);
or U33963 (N_33963,N_30323,N_30359);
nor U33964 (N_33964,N_30104,N_30541);
and U33965 (N_33965,N_31453,N_30953);
or U33966 (N_33966,N_31888,N_30210);
nand U33967 (N_33967,N_30166,N_31232);
and U33968 (N_33968,N_30220,N_31327);
or U33969 (N_33969,N_31817,N_31933);
or U33970 (N_33970,N_30934,N_31251);
and U33971 (N_33971,N_31586,N_30469);
and U33972 (N_33972,N_30170,N_31639);
nand U33973 (N_33973,N_30642,N_31282);
or U33974 (N_33974,N_30855,N_31888);
nor U33975 (N_33975,N_30138,N_30085);
nand U33976 (N_33976,N_31987,N_30393);
nand U33977 (N_33977,N_30911,N_31965);
nand U33978 (N_33978,N_31162,N_30582);
or U33979 (N_33979,N_31790,N_30433);
nand U33980 (N_33980,N_31285,N_31085);
or U33981 (N_33981,N_30670,N_31093);
nor U33982 (N_33982,N_31743,N_31822);
or U33983 (N_33983,N_31484,N_30136);
and U33984 (N_33984,N_30470,N_30214);
nand U33985 (N_33985,N_30127,N_30005);
and U33986 (N_33986,N_31443,N_30296);
nor U33987 (N_33987,N_31229,N_30828);
and U33988 (N_33988,N_31220,N_30410);
nand U33989 (N_33989,N_30745,N_30969);
nor U33990 (N_33990,N_30193,N_31595);
nand U33991 (N_33991,N_31833,N_30128);
nor U33992 (N_33992,N_31876,N_30870);
nor U33993 (N_33993,N_31164,N_31536);
and U33994 (N_33994,N_31738,N_31934);
or U33995 (N_33995,N_30631,N_30796);
xor U33996 (N_33996,N_31489,N_31306);
and U33997 (N_33997,N_30603,N_31409);
or U33998 (N_33998,N_31409,N_30651);
xor U33999 (N_33999,N_30695,N_30113);
or U34000 (N_34000,N_33170,N_32063);
or U34001 (N_34001,N_32330,N_33434);
and U34002 (N_34002,N_33481,N_32402);
and U34003 (N_34003,N_33265,N_33973);
nor U34004 (N_34004,N_32831,N_32580);
nand U34005 (N_34005,N_32799,N_32228);
and U34006 (N_34006,N_33310,N_32690);
xnor U34007 (N_34007,N_32396,N_33724);
and U34008 (N_34008,N_32768,N_33544);
xor U34009 (N_34009,N_33242,N_33528);
and U34010 (N_34010,N_32339,N_32382);
xnor U34011 (N_34011,N_33953,N_33708);
nand U34012 (N_34012,N_32238,N_33014);
or U34013 (N_34013,N_33781,N_32490);
or U34014 (N_34014,N_33063,N_33568);
or U34015 (N_34015,N_33155,N_32222);
and U34016 (N_34016,N_32877,N_32306);
or U34017 (N_34017,N_32242,N_33886);
nor U34018 (N_34018,N_33513,N_33093);
nor U34019 (N_34019,N_33248,N_32884);
or U34020 (N_34020,N_32621,N_32018);
nand U34021 (N_34021,N_32077,N_33668);
nand U34022 (N_34022,N_32694,N_33349);
nor U34023 (N_34023,N_33984,N_33543);
nand U34024 (N_34024,N_33429,N_33216);
and U34025 (N_34025,N_33793,N_32638);
xnor U34026 (N_34026,N_32950,N_32533);
nor U34027 (N_34027,N_32375,N_32604);
nor U34028 (N_34028,N_32168,N_33979);
xnor U34029 (N_34029,N_32119,N_33833);
nand U34030 (N_34030,N_33713,N_32451);
nand U34031 (N_34031,N_33849,N_32867);
nor U34032 (N_34032,N_33067,N_32160);
and U34033 (N_34033,N_33675,N_32701);
nand U34034 (N_34034,N_32613,N_33076);
nor U34035 (N_34035,N_33844,N_33601);
xnor U34036 (N_34036,N_32996,N_32344);
nand U34037 (N_34037,N_32422,N_32516);
or U34038 (N_34038,N_32629,N_33256);
nor U34039 (N_34039,N_32166,N_32637);
nand U34040 (N_34040,N_32301,N_32194);
nand U34041 (N_34041,N_33400,N_32219);
and U34042 (N_34042,N_32936,N_33191);
xor U34043 (N_34043,N_32591,N_32894);
nand U34044 (N_34044,N_33355,N_33152);
nor U34045 (N_34045,N_32568,N_33402);
and U34046 (N_34046,N_32800,N_33970);
xnor U34047 (N_34047,N_33121,N_32984);
and U34048 (N_34048,N_32079,N_32805);
or U34049 (N_34049,N_33459,N_33512);
nor U34050 (N_34050,N_32379,N_33928);
or U34051 (N_34051,N_32862,N_32214);
or U34052 (N_34052,N_32248,N_32612);
or U34053 (N_34053,N_33674,N_32145);
nor U34054 (N_34054,N_33077,N_33041);
nand U34055 (N_34055,N_33086,N_32947);
or U34056 (N_34056,N_33068,N_33106);
nor U34057 (N_34057,N_32876,N_32466);
nor U34058 (N_34058,N_33754,N_33599);
nor U34059 (N_34059,N_32907,N_33382);
nand U34060 (N_34060,N_33343,N_33908);
and U34061 (N_34061,N_33390,N_32473);
or U34062 (N_34062,N_32897,N_33328);
nand U34063 (N_34063,N_33315,N_33285);
and U34064 (N_34064,N_32929,N_32861);
xor U34065 (N_34065,N_32399,N_32365);
nor U34066 (N_34066,N_33882,N_33160);
and U34067 (N_34067,N_33201,N_33769);
nand U34068 (N_34068,N_33969,N_32348);
and U34069 (N_34069,N_33171,N_32767);
nor U34070 (N_34070,N_33053,N_32529);
nand U34071 (N_34071,N_33709,N_33138);
and U34072 (N_34072,N_33236,N_32276);
or U34073 (N_34073,N_32314,N_32822);
nor U34074 (N_34074,N_33579,N_33013);
nor U34075 (N_34075,N_33592,N_32112);
or U34076 (N_34076,N_32691,N_32810);
xnor U34077 (N_34077,N_32447,N_32474);
nor U34078 (N_34078,N_32974,N_33021);
nor U34079 (N_34079,N_33146,N_32304);
and U34080 (N_34080,N_32842,N_33116);
and U34081 (N_34081,N_33430,N_33375);
and U34082 (N_34082,N_33370,N_33472);
or U34083 (N_34083,N_33190,N_33837);
nand U34084 (N_34084,N_32573,N_33945);
nor U34085 (N_34085,N_32007,N_32679);
xor U34086 (N_34086,N_33271,N_33624);
xnor U34087 (N_34087,N_33123,N_32744);
and U34088 (N_34088,N_32059,N_33727);
or U34089 (N_34089,N_32284,N_32383);
nor U34090 (N_34090,N_33029,N_33504);
nand U34091 (N_34091,N_32987,N_33110);
and U34092 (N_34092,N_32541,N_33209);
or U34093 (N_34093,N_32468,N_32766);
and U34094 (N_34094,N_32983,N_32860);
or U34095 (N_34095,N_33900,N_32985);
nor U34096 (N_34096,N_32662,N_33738);
nand U34097 (N_34097,N_32994,N_33646);
nand U34098 (N_34098,N_32523,N_32427);
xor U34099 (N_34099,N_32013,N_32785);
nor U34100 (N_34100,N_32885,N_32711);
nand U34101 (N_34101,N_33433,N_33862);
nor U34102 (N_34102,N_32132,N_33613);
and U34103 (N_34103,N_32170,N_32764);
xnor U34104 (N_34104,N_32715,N_32808);
nor U34105 (N_34105,N_32589,N_32497);
and U34106 (N_34106,N_32724,N_33350);
nand U34107 (N_34107,N_32827,N_32685);
xor U34108 (N_34108,N_33774,N_33647);
nand U34109 (N_34109,N_32297,N_33949);
nand U34110 (N_34110,N_33748,N_33700);
nor U34111 (N_34111,N_32491,N_33799);
nand U34112 (N_34112,N_32037,N_33241);
or U34113 (N_34113,N_32866,N_33286);
or U34114 (N_34114,N_32239,N_32444);
nor U34115 (N_34115,N_33427,N_33173);
nor U34116 (N_34116,N_33635,N_33258);
and U34117 (N_34117,N_33377,N_33416);
nor U34118 (N_34118,N_33224,N_32051);
nor U34119 (N_34119,N_32780,N_33746);
and U34120 (N_34120,N_32281,N_32957);
and U34121 (N_34121,N_33588,N_33845);
and U34122 (N_34122,N_32187,N_32110);
nand U34123 (N_34123,N_32883,N_33932);
nand U34124 (N_34124,N_33560,N_33387);
and U34125 (N_34125,N_33864,N_33712);
nor U34126 (N_34126,N_32153,N_33643);
and U34127 (N_34127,N_32118,N_33348);
nor U34128 (N_34128,N_32359,N_33743);
xnor U34129 (N_34129,N_32012,N_33361);
nand U34130 (N_34130,N_32113,N_33278);
nand U34131 (N_34131,N_32185,N_32068);
or U34132 (N_34132,N_32259,N_33523);
nor U34133 (N_34133,N_33752,N_33473);
or U34134 (N_34134,N_33688,N_32991);
xnor U34135 (N_34135,N_32158,N_32682);
or U34136 (N_34136,N_32699,N_32421);
nand U34137 (N_34137,N_33820,N_32963);
or U34138 (N_34138,N_32627,N_32943);
xnor U34139 (N_34139,N_32659,N_32846);
xor U34140 (N_34140,N_32819,N_32146);
and U34141 (N_34141,N_32881,N_33642);
nor U34142 (N_34142,N_33567,N_32139);
xor U34143 (N_34143,N_32631,N_33220);
nand U34144 (N_34144,N_33344,N_32485);
nand U34145 (N_34145,N_32742,N_33060);
or U34146 (N_34146,N_32598,N_32961);
and U34147 (N_34147,N_33788,N_33454);
and U34148 (N_34148,N_33693,N_33254);
nor U34149 (N_34149,N_32520,N_32770);
or U34150 (N_34150,N_32835,N_33796);
xor U34151 (N_34151,N_33482,N_32346);
nor U34152 (N_34152,N_33345,N_32845);
nor U34153 (N_34153,N_33916,N_33866);
and U34154 (N_34154,N_32585,N_33011);
nor U34155 (N_34155,N_33234,N_32420);
xor U34156 (N_34156,N_33035,N_33148);
nor U34157 (N_34157,N_32039,N_32385);
and U34158 (N_34158,N_33246,N_33817);
nor U34159 (N_34159,N_33530,N_32456);
nor U34160 (N_34160,N_32056,N_32925);
nor U34161 (N_34161,N_33692,N_32046);
xnor U34162 (N_34162,N_32439,N_33235);
nand U34163 (N_34163,N_33983,N_32206);
or U34164 (N_34164,N_32188,N_32472);
and U34165 (N_34165,N_33919,N_32315);
nor U34166 (N_34166,N_33050,N_32605);
and U34167 (N_34167,N_32036,N_33540);
nor U34168 (N_34168,N_33571,N_32848);
nand U34169 (N_34169,N_32593,N_32600);
nor U34170 (N_34170,N_32436,N_32488);
or U34171 (N_34171,N_33178,N_32745);
or U34172 (N_34172,N_32620,N_32147);
xor U34173 (N_34173,N_33480,N_32644);
and U34174 (N_34174,N_32102,N_33841);
nor U34175 (N_34175,N_33156,N_33912);
nor U34176 (N_34176,N_33701,N_32140);
xnor U34177 (N_34177,N_33852,N_32412);
xnor U34178 (N_34178,N_32483,N_32226);
nor U34179 (N_34179,N_32732,N_33702);
xor U34180 (N_34180,N_32367,N_33356);
nor U34181 (N_34181,N_32834,N_33442);
nand U34182 (N_34182,N_33295,N_32312);
or U34183 (N_34183,N_33891,N_33197);
nand U34184 (N_34184,N_33678,N_33778);
or U34185 (N_34185,N_33651,N_32939);
and U34186 (N_34186,N_33135,N_32434);
and U34187 (N_34187,N_32806,N_33419);
nand U34188 (N_34188,N_33009,N_33058);
or U34189 (N_34189,N_33941,N_32435);
nor U34190 (N_34190,N_32993,N_32671);
xor U34191 (N_34191,N_33398,N_33325);
nor U34192 (N_34192,N_32262,N_32017);
nand U34193 (N_34193,N_32769,N_32651);
nand U34194 (N_34194,N_33477,N_32578);
nor U34195 (N_34195,N_32730,N_32625);
xnor U34196 (N_34196,N_33252,N_32195);
nor U34197 (N_34197,N_32400,N_33463);
nor U34198 (N_34198,N_32997,N_32986);
nor U34199 (N_34199,N_32229,N_32441);
and U34200 (N_34200,N_32771,N_32044);
nor U34201 (N_34201,N_32184,N_33410);
xor U34202 (N_34202,N_32398,N_32511);
nand U34203 (N_34203,N_33054,N_32611);
nor U34204 (N_34204,N_33184,N_33997);
nand U34205 (N_34205,N_33204,N_32521);
or U34206 (N_34206,N_32514,N_32999);
xor U34207 (N_34207,N_32384,N_32614);
or U34208 (N_34208,N_32675,N_32972);
xor U34209 (N_34209,N_33633,N_32820);
nor U34210 (N_34210,N_32791,N_32731);
or U34211 (N_34211,N_33260,N_32905);
and U34212 (N_34212,N_32308,N_32107);
or U34213 (N_34213,N_32967,N_33194);
xor U34214 (N_34214,N_33189,N_33244);
and U34215 (N_34215,N_32221,N_33441);
xor U34216 (N_34216,N_32864,N_33373);
or U34217 (N_34217,N_33968,N_33437);
nor U34218 (N_34218,N_32129,N_33509);
nor U34219 (N_34219,N_33944,N_32413);
xor U34220 (N_34220,N_33545,N_33362);
nor U34221 (N_34221,N_32250,N_32932);
nand U34222 (N_34222,N_32686,N_32215);
nand U34223 (N_34223,N_33306,N_32544);
and U34224 (N_34224,N_32896,N_32193);
xnor U34225 (N_34225,N_33718,N_33091);
nand U34226 (N_34226,N_33906,N_33008);
xnor U34227 (N_34227,N_32000,N_32163);
and U34228 (N_34228,N_33109,N_33609);
xor U34229 (N_34229,N_32200,N_32761);
nand U34230 (N_34230,N_33296,N_32350);
and U34231 (N_34231,N_33280,N_33959);
and U34232 (N_34232,N_32032,N_33962);
or U34233 (N_34233,N_32002,N_32498);
xor U34234 (N_34234,N_32204,N_32325);
nand U34235 (N_34235,N_32403,N_32287);
xor U34236 (N_34236,N_33961,N_32607);
xor U34237 (N_34237,N_33287,N_32151);
nor U34238 (N_34238,N_32295,N_32269);
or U34239 (N_34239,N_33137,N_32760);
and U34240 (N_34240,N_32091,N_32716);
and U34241 (N_34241,N_33233,N_32759);
nand U34242 (N_34242,N_33605,N_32336);
nand U34243 (N_34243,N_32050,N_32366);
nor U34244 (N_34244,N_33208,N_32826);
xnor U34245 (N_34245,N_32735,N_32504);
xnor U34246 (N_34246,N_32500,N_32554);
nor U34247 (N_34247,N_32020,N_33075);
nand U34248 (N_34248,N_32198,N_32829);
nand U34249 (N_34249,N_32092,N_33681);
nand U34250 (N_34250,N_32508,N_33131);
and U34251 (N_34251,N_32847,N_33823);
xor U34252 (N_34252,N_32137,N_32776);
nor U34253 (N_34253,N_33324,N_32237);
xnor U34254 (N_34254,N_33498,N_33818);
xnor U34255 (N_34255,N_32035,N_32841);
or U34256 (N_34256,N_32225,N_32234);
nand U34257 (N_34257,N_32178,N_33124);
xor U34258 (N_34258,N_33819,N_33810);
and U34259 (N_34259,N_32481,N_32177);
or U34260 (N_34260,N_32510,N_33083);
xnor U34261 (N_34261,N_32362,N_33409);
xor U34262 (N_34262,N_32296,N_33861);
nand U34263 (N_34263,N_33689,N_32960);
xor U34264 (N_34264,N_33948,N_33552);
or U34265 (N_34265,N_33604,N_32927);
nand U34266 (N_34266,N_32934,N_32755);
nor U34267 (N_34267,N_32666,N_33654);
xnor U34268 (N_34268,N_32090,N_33226);
or U34269 (N_34269,N_33003,N_32428);
nor U34270 (N_34270,N_33926,N_33040);
xnor U34271 (N_34271,N_33770,N_33016);
nand U34272 (N_34272,N_32734,N_33842);
or U34273 (N_34273,N_33198,N_33839);
or U34274 (N_34274,N_33073,N_32062);
nor U34275 (N_34275,N_32212,N_33612);
and U34276 (N_34276,N_32689,N_33697);
and U34277 (N_34277,N_33631,N_32721);
and U34278 (N_34278,N_32432,N_33267);
nand U34279 (N_34279,N_32626,N_33895);
and U34280 (N_34280,N_33611,N_33221);
or U34281 (N_34281,N_32705,N_32356);
nand U34282 (N_34282,N_32850,N_33090);
nand U34283 (N_34283,N_33294,N_33078);
xor U34284 (N_34284,N_32373,N_32388);
and U34285 (N_34285,N_32702,N_33537);
nand U34286 (N_34286,N_32155,N_32317);
and U34287 (N_34287,N_33158,N_33637);
and U34288 (N_34288,N_33232,N_33307);
nand U34289 (N_34289,N_32190,N_33925);
nor U34290 (N_34290,N_33538,N_33596);
nor U34291 (N_34291,N_33905,N_32571);
and U34292 (N_34292,N_33034,N_32804);
xnor U34293 (N_34293,N_33411,N_33811);
and U34294 (N_34294,N_33780,N_33314);
nor U34295 (N_34295,N_33255,N_32291);
and U34296 (N_34296,N_32293,N_33993);
nand U34297 (N_34297,N_33565,N_33469);
or U34298 (N_34298,N_33079,N_32220);
nor U34299 (N_34299,N_33268,N_33859);
nand U34300 (N_34300,N_32069,N_33533);
or U34301 (N_34301,N_32969,N_32552);
xor U34302 (N_34302,N_32639,N_33087);
xnor U34303 (N_34303,N_32230,N_32501);
and U34304 (N_34304,N_33955,N_32703);
and U34305 (N_34305,N_33435,N_33321);
and U34306 (N_34306,N_33176,N_33134);
nor U34307 (N_34307,N_33212,N_32796);
or U34308 (N_34308,N_33329,N_32323);
nor U34309 (N_34309,N_32469,N_33351);
nand U34310 (N_34310,N_33496,N_32725);
nor U34311 (N_34311,N_33102,N_32249);
nor U34312 (N_34312,N_32455,N_33207);
xor U34313 (N_34313,N_32461,N_32706);
and U34314 (N_34314,N_32213,N_33726);
nand U34315 (N_34315,N_33193,N_32161);
and U34316 (N_34316,N_32545,N_32966);
or U34317 (N_34317,N_33840,N_32824);
nor U34318 (N_34318,N_33829,N_32729);
nand U34319 (N_34319,N_32749,N_33958);
and U34320 (N_34320,N_33696,N_33239);
or U34321 (N_34321,N_32021,N_33036);
nor U34322 (N_34322,N_33966,N_32101);
nor U34323 (N_34323,N_33992,N_33911);
and U34324 (N_34324,N_33714,N_32543);
nand U34325 (N_34325,N_32556,N_32154);
nor U34326 (N_34326,N_32450,N_32289);
nor U34327 (N_34327,N_33118,N_32429);
xnor U34328 (N_34328,N_32658,N_33786);
and U34329 (N_34329,N_33378,N_32442);
xor U34330 (N_34330,N_33535,N_33639);
nand U34331 (N_34331,N_33517,N_32148);
and U34332 (N_34332,N_33047,N_32318);
or U34333 (N_34333,N_33519,N_32437);
or U34334 (N_34334,N_32418,N_33486);
xnor U34335 (N_34335,N_33835,N_33154);
and U34336 (N_34336,N_32913,N_32643);
or U34337 (N_34337,N_33071,N_33673);
nand U34338 (N_34338,N_32888,N_33333);
and U34339 (N_34339,N_32494,N_33264);
and U34340 (N_34340,N_33455,N_32989);
or U34341 (N_34341,N_33334,N_33991);
or U34342 (N_34342,N_32098,N_33698);
nor U34343 (N_34343,N_33153,N_33924);
nor U34344 (N_34344,N_32663,N_32778);
nand U34345 (N_34345,N_32043,N_32417);
nand U34346 (N_34346,N_33299,N_32294);
or U34347 (N_34347,N_33245,N_33465);
nor U34348 (N_34348,N_33619,N_32199);
nor U34349 (N_34349,N_33057,N_32123);
or U34350 (N_34350,N_32622,N_32893);
or U34351 (N_34351,N_32584,N_33331);
and U34352 (N_34352,N_32232,N_33880);
nand U34353 (N_34353,N_32116,N_32870);
xor U34354 (N_34354,N_33423,N_32825);
or U34355 (N_34355,N_32014,N_33479);
nand U34356 (N_34356,N_33061,N_33575);
nand U34357 (N_34357,N_32836,N_32487);
nand U34358 (N_34358,N_33529,N_33359);
nand U34359 (N_34359,N_32134,N_32332);
xnor U34360 (N_34360,N_32914,N_32048);
or U34361 (N_34361,N_32587,N_32650);
xor U34362 (N_34362,N_33098,N_32546);
nor U34363 (N_34363,N_32136,N_33401);
nor U34364 (N_34364,N_33431,N_33518);
or U34365 (N_34365,N_32668,N_32231);
and U34366 (N_34366,N_33775,N_33272);
and U34367 (N_34367,N_33289,N_32677);
nor U34368 (N_34368,N_32211,N_32272);
nand U34369 (N_34369,N_33615,N_32944);
or U34370 (N_34370,N_33822,N_33963);
and U34371 (N_34371,N_32073,N_33937);
xor U34372 (N_34372,N_32575,N_32673);
xnor U34373 (N_34373,N_33873,N_33863);
and U34374 (N_34374,N_33998,N_33987);
xnor U34375 (N_34375,N_32890,N_33921);
nand U34376 (N_34376,N_32784,N_33732);
and U34377 (N_34377,N_32542,N_33199);
nand U34378 (N_34378,N_32124,N_33850);
xor U34379 (N_34379,N_33846,N_32223);
nor U34380 (N_34380,N_32080,N_33650);
xor U34381 (N_34381,N_33574,N_33466);
nor U34382 (N_34382,N_33450,N_32322);
xnor U34383 (N_34383,N_33843,N_33725);
nand U34384 (N_34384,N_33890,N_33894);
nand U34385 (N_34385,N_32548,N_33447);
nor U34386 (N_34386,N_32258,N_32235);
nor U34387 (N_34387,N_33671,N_33132);
xor U34388 (N_34388,N_32875,N_32712);
nor U34389 (N_34389,N_33326,N_32426);
xor U34390 (N_34390,N_32353,N_32696);
and U34391 (N_34391,N_32754,N_32802);
and U34392 (N_34392,N_32126,N_33293);
xor U34393 (N_34393,N_32465,N_32047);
nand U34394 (N_34394,N_33551,N_32979);
nand U34395 (N_34395,N_33300,N_32904);
xnor U34396 (N_34396,N_33169,N_32528);
or U34397 (N_34397,N_33857,N_32395);
nor U34398 (N_34398,N_32719,N_32391);
xor U34399 (N_34399,N_33603,N_33147);
xnor U34400 (N_34400,N_33557,N_33901);
nor U34401 (N_34401,N_32093,N_33658);
xor U34402 (N_34402,N_33468,N_32096);
nor U34403 (N_34403,N_33855,N_33940);
nor U34404 (N_34404,N_33340,N_33030);
nor U34405 (N_34405,N_32029,N_33046);
and U34406 (N_34406,N_33162,N_32164);
nor U34407 (N_34407,N_33273,N_32457);
xnor U34408 (N_34408,N_32409,N_32560);
and U34409 (N_34409,N_32471,N_33974);
nand U34410 (N_34410,N_32181,N_33261);
and U34411 (N_34411,N_32347,N_33577);
nand U34412 (N_34412,N_32801,N_33206);
nor U34413 (N_34413,N_32975,N_33004);
or U34414 (N_34414,N_33525,N_32111);
nor U34415 (N_34415,N_33589,N_33074);
and U34416 (N_34416,N_32486,N_32410);
xor U34417 (N_34417,N_32202,N_33986);
or U34418 (N_34418,N_32290,N_32540);
nand U34419 (N_34419,N_32302,N_33581);
xor U34420 (N_34420,N_33556,N_32513);
nand U34421 (N_34421,N_32815,N_33622);
xnor U34422 (N_34422,N_33656,N_32071);
and U34423 (N_34423,N_33436,N_32128);
nor U34424 (N_34424,N_32493,N_32814);
nand U34425 (N_34425,N_32567,N_32641);
nor U34426 (N_34426,N_33462,N_33122);
and U34427 (N_34427,N_32646,N_32608);
and U34428 (N_34428,N_32592,N_33186);
xnor U34429 (N_34429,N_33794,N_33710);
xnor U34430 (N_34430,N_33425,N_33165);
nor U34431 (N_34431,N_33231,N_32954);
nand U34432 (N_34432,N_32415,N_32443);
or U34433 (N_34433,N_33735,N_32670);
and U34434 (N_34434,N_33586,N_32479);
or U34435 (N_34435,N_33225,N_33745);
nor U34436 (N_34436,N_32937,N_32619);
or U34437 (N_34437,N_33755,N_33716);
or U34438 (N_34438,N_32135,N_33521);
xor U34439 (N_34439,N_33851,N_32590);
nor U34440 (N_34440,N_33027,N_33301);
and U34441 (N_34441,N_33766,N_33797);
or U34442 (N_34442,N_32535,N_32564);
nand U34443 (N_34443,N_33505,N_33825);
nand U34444 (N_34444,N_32865,N_32928);
nand U34445 (N_34445,N_32241,N_32763);
or U34446 (N_34446,N_33747,N_32956);
nand U34447 (N_34447,N_33302,N_32218);
nor U34448 (N_34448,N_32901,N_33493);
or U34449 (N_34449,N_33039,N_33108);
nand U34450 (N_34450,N_32311,N_33044);
nand U34451 (N_34451,N_33376,N_33470);
and U34452 (N_34452,N_33330,N_33412);
nor U34453 (N_34453,N_32786,N_32015);
or U34454 (N_34454,N_32343,N_32746);
xnor U34455 (N_34455,N_33903,N_33621);
and U34456 (N_34456,N_33291,N_32931);
and U34457 (N_34457,N_33790,N_33305);
or U34458 (N_34458,N_33043,N_32374);
and U34459 (N_34459,N_32109,N_33371);
xnor U34460 (N_34460,N_33303,N_32681);
xnor U34461 (N_34461,N_33520,N_33798);
nor U34462 (N_34462,N_32390,N_32852);
nand U34463 (N_34463,N_33451,N_32811);
or U34464 (N_34464,N_33742,N_33446);
nand U34465 (N_34465,N_32171,N_33597);
or U34466 (N_34466,N_33943,N_32175);
and U34467 (N_34467,N_33750,N_33508);
and U34468 (N_34468,N_33690,N_32714);
xor U34469 (N_34469,N_33610,N_32602);
or U34470 (N_34470,N_32738,N_33089);
or U34471 (N_34471,N_33002,N_32741);
xnor U34472 (N_34472,N_32868,N_32874);
nor U34473 (N_34473,N_33276,N_33816);
nand U34474 (N_34474,N_33934,N_33478);
or U34475 (N_34475,N_32698,N_32895);
xnor U34476 (N_34476,N_33595,N_33792);
nor U34477 (N_34477,N_33534,N_33210);
nor U34478 (N_34478,N_32817,N_33187);
nand U34479 (N_34479,N_32462,N_32261);
xnor U34480 (N_34480,N_33795,N_33380);
nor U34481 (N_34481,N_33237,N_32774);
nor U34482 (N_34482,N_33227,N_33358);
nand U34483 (N_34483,N_33616,N_33335);
or U34484 (N_34484,N_32955,N_32618);
xor U34485 (N_34485,N_32022,N_33458);
nand U34486 (N_34486,N_33149,N_33432);
nand U34487 (N_34487,N_33954,N_33219);
and U34488 (N_34488,N_32270,N_32710);
nor U34489 (N_34489,N_33100,N_33125);
xnor U34490 (N_34490,N_33805,N_32089);
nand U34491 (N_34491,N_33767,N_32998);
nor U34492 (N_34492,N_33942,N_32886);
or U34493 (N_34493,N_32354,N_32106);
nand U34494 (N_34494,N_32201,N_33872);
and U34495 (N_34495,N_32803,N_32532);
and U34496 (N_34496,N_33995,N_33449);
nand U34497 (N_34497,N_32665,N_33563);
xor U34498 (N_34498,N_33316,N_33977);
xor U34499 (N_34499,N_33670,N_33284);
nor U34500 (N_34500,N_33001,N_33452);
and U34501 (N_34501,N_32172,N_33308);
or U34502 (N_34502,N_33809,N_33240);
nor U34503 (N_34503,N_33617,N_32962);
and U34504 (N_34504,N_33005,N_33893);
and U34505 (N_34505,N_32011,N_32891);
or U34506 (N_34506,N_33982,N_33645);
nand U34507 (N_34507,N_33394,N_33706);
and U34508 (N_34508,N_32509,N_33368);
nor U34509 (N_34509,N_33672,N_32773);
nand U34510 (N_34510,N_33573,N_32300);
xor U34511 (N_34511,N_32753,N_32086);
nand U34512 (N_34512,N_33322,N_33570);
and U34513 (N_34513,N_32777,N_32949);
or U34514 (N_34514,N_32207,N_33317);
nor U34515 (N_34515,N_32480,N_32349);
xnor U34516 (N_34516,N_32438,N_33623);
or U34517 (N_34517,N_33386,N_32411);
xnor U34518 (N_34518,N_32031,N_32227);
nand U34519 (N_34519,N_33460,N_33023);
xor U34520 (N_34520,N_33103,N_33020);
nor U34521 (N_34521,N_33728,N_32657);
and U34522 (N_34522,N_32327,N_33277);
or U34523 (N_34523,N_33806,N_33608);
nand U34524 (N_34524,N_32019,N_33065);
xnor U34525 (N_34525,N_32722,N_32143);
or U34526 (N_34526,N_32448,N_33641);
xnor U34527 (N_34527,N_32783,N_32727);
and U34528 (N_34528,N_32667,N_32704);
nor U34529 (N_34529,N_32920,N_33657);
or U34530 (N_34530,N_33881,N_32839);
or U34531 (N_34531,N_32209,N_32912);
and U34532 (N_34532,N_33999,N_32557);
xnor U34533 (N_34533,N_33099,N_33707);
nor U34534 (N_34534,N_32977,N_33161);
xor U34535 (N_34535,N_32251,N_33860);
and U34536 (N_34536,N_32572,N_33105);
and U34537 (N_34537,N_33026,N_33682);
or U34538 (N_34538,N_32357,N_32319);
or U34539 (N_34539,N_33323,N_32566);
or U34540 (N_34540,N_33407,N_33485);
xnor U34541 (N_34541,N_32813,N_33628);
nor U34542 (N_34542,N_32088,N_33055);
nor U34543 (N_34543,N_32601,N_33304);
or U34544 (N_34544,N_33753,N_33813);
nor U34545 (N_34545,N_33787,N_32243);
or U34546 (N_34546,N_33909,N_33676);
or U34547 (N_34547,N_32726,N_33789);
and U34548 (N_34548,N_32594,N_32652);
nand U34549 (N_34549,N_32562,N_32024);
and U34550 (N_34550,N_32338,N_32352);
xnor U34551 (N_34551,N_32360,N_33404);
and U34552 (N_34552,N_32597,N_32458);
nor U34553 (N_34553,N_32603,N_33757);
nor U34554 (N_34554,N_32416,N_33988);
xnor U34555 (N_34555,N_32423,N_33388);
and U34556 (N_34556,N_32463,N_33364);
and U34557 (N_34557,N_33907,N_32515);
and U34558 (N_34558,N_33667,N_32064);
nor U34559 (N_34559,N_32616,N_32397);
nor U34560 (N_34560,N_32253,N_32404);
nor U34561 (N_34561,N_32733,N_32747);
or U34562 (N_34562,N_32299,N_32167);
or U34563 (N_34563,N_33389,N_32368);
or U34564 (N_34564,N_32358,N_33956);
nor U34565 (N_34565,N_32271,N_33729);
nand U34566 (N_34566,N_33526,N_32152);
xnor U34567 (N_34567,N_32240,N_33808);
nand U34568 (N_34568,N_32882,N_32782);
or U34569 (N_34569,N_32736,N_32182);
nand U34570 (N_34570,N_32775,N_32538);
xor U34571 (N_34571,N_33952,N_32723);
nand U34572 (N_34572,N_33269,N_32973);
and U34573 (N_34573,N_33347,N_33028);
xnor U34574 (N_34574,N_33374,N_33522);
or U34575 (N_34575,N_33163,N_33064);
xor U34576 (N_34576,N_32709,N_33445);
nand U34577 (N_34577,N_33045,N_32816);
nand U34578 (N_34578,N_33288,N_33136);
or U34579 (N_34579,N_33126,N_33365);
nor U34580 (N_34580,N_33217,N_32133);
nand U34581 (N_34581,N_32203,N_33414);
nand U34582 (N_34582,N_32157,N_32933);
nand U34583 (N_34583,N_32921,N_32869);
xor U34584 (N_34584,N_32549,N_33180);
xor U34585 (N_34585,N_32918,N_33166);
xor U34586 (N_34586,N_33015,N_32807);
and U34587 (N_34587,N_33889,N_32978);
and U34588 (N_34588,N_33483,N_33768);
nor U34589 (N_34589,N_32863,N_32697);
and U34590 (N_34590,N_33413,N_32654);
or U34591 (N_34591,N_33975,N_33555);
or U34592 (N_34592,N_32205,N_32900);
or U34593 (N_34593,N_32174,N_32303);
or U34594 (N_34594,N_32823,N_33687);
nand U34595 (N_34595,N_32908,N_33150);
nor U34596 (N_34596,N_32341,N_33017);
nand U34597 (N_34597,N_33475,N_33765);
nand U34598 (N_34598,N_33168,N_33867);
nor U34599 (N_34599,N_32292,N_33868);
nand U34600 (N_34600,N_32316,N_32305);
or U34601 (N_34601,N_33853,N_33346);
nand U34602 (N_34602,N_32524,N_32162);
nand U34603 (N_34603,N_33721,N_32406);
nor U34604 (N_34604,N_32286,N_32843);
or U34605 (N_34605,N_33532,N_33120);
or U34606 (N_34606,N_32335,N_33274);
nor U34607 (N_34607,N_32700,N_32452);
or U34608 (N_34608,N_33546,N_33205);
and U34609 (N_34609,N_33715,N_32649);
or U34610 (N_34610,N_33403,N_33476);
nor U34611 (N_34611,N_33717,N_33749);
xnor U34612 (N_34612,N_32653,N_32094);
nor U34613 (N_34613,N_33634,N_32298);
nor U34614 (N_34614,N_33764,N_33602);
xor U34615 (N_34615,N_33583,N_32953);
nand U34616 (N_34616,N_33461,N_32169);
and U34617 (N_34617,N_32337,N_33415);
nand U34618 (N_34618,N_32507,N_32288);
xnor U34619 (N_34619,N_32854,N_33874);
nor U34620 (N_34620,N_33640,N_33369);
or U34621 (N_34621,N_32503,N_32923);
or U34622 (N_34622,N_32165,N_32142);
nor U34623 (N_34623,N_33677,N_33549);
xor U34624 (N_34624,N_32027,N_32108);
and U34625 (N_34625,N_33838,N_32630);
xnor U34626 (N_34626,N_32553,N_33569);
nor U34627 (N_34627,N_32282,N_32467);
xor U34628 (N_34628,N_33824,N_33664);
and U34629 (N_34629,N_33737,N_33910);
nor U34630 (N_34630,N_33980,N_32581);
or U34631 (N_34631,N_33510,N_33554);
xnor U34632 (N_34632,N_33627,N_33930);
xor U34633 (N_34633,N_33929,N_32506);
and U34634 (N_34634,N_32256,N_32926);
or U34635 (N_34635,N_33783,N_33699);
or U34636 (N_34636,N_33489,N_33630);
nor U34637 (N_34637,N_33593,N_33270);
nor U34638 (N_34638,N_32309,N_33947);
xor U34639 (N_34639,N_32260,N_33902);
nand U34640 (N_34640,N_32058,N_32559);
or U34641 (N_34641,N_33585,N_32636);
nor U34642 (N_34642,N_32130,N_33502);
nor U34643 (N_34643,N_33366,N_32935);
xor U34644 (N_34644,N_33553,N_33965);
nand U34645 (N_34645,N_33876,N_32797);
and U34646 (N_34646,N_33694,N_33740);
and U34647 (N_34647,N_33066,N_33426);
nand U34648 (N_34648,N_32672,N_33195);
xnor U34649 (N_34649,N_33095,N_32648);
nor U34650 (N_34650,N_32361,N_33457);
nand U34651 (N_34651,N_32010,N_33084);
nor U34652 (N_34652,N_33695,N_33157);
and U34653 (N_34653,N_33311,N_33177);
and U34654 (N_34654,N_33777,N_33140);
and U34655 (N_34655,N_33019,N_32569);
xor U34656 (N_34656,N_32517,N_33878);
nand U34657 (N_34657,N_33736,N_32534);
nor U34658 (N_34658,N_32057,N_33572);
or U34659 (N_34659,N_32083,N_33000);
xnor U34660 (N_34660,N_32656,N_33620);
or U34661 (N_34661,N_33097,N_32006);
and U34662 (N_34662,N_32851,N_33669);
nor U34663 (N_34663,N_32976,N_32042);
or U34664 (N_34664,N_33587,N_32902);
or U34665 (N_34665,N_33875,N_33663);
and U34666 (N_34666,N_33936,N_32247);
xnor U34667 (N_34667,N_32028,N_33547);
nand U34668 (N_34668,N_32389,N_32245);
xnor U34669 (N_34669,N_33497,N_32433);
or U34670 (N_34670,N_33638,N_32454);
xor U34671 (N_34671,N_32586,N_32192);
or U34672 (N_34672,N_33751,N_33514);
and U34673 (N_34673,N_32351,N_33598);
and U34674 (N_34674,N_32906,N_33847);
and U34675 (N_34675,N_33784,N_32100);
or U34676 (N_34676,N_33379,N_32326);
nor U34677 (N_34677,N_32674,N_33957);
xnor U34678 (N_34678,N_33056,N_33275);
nor U34679 (N_34679,N_32609,N_32489);
and U34680 (N_34680,N_33812,N_33491);
and U34681 (N_34681,N_33499,N_33744);
and U34682 (N_34682,N_32264,N_32790);
xor U34683 (N_34683,N_33381,N_32074);
nor U34684 (N_34684,N_32695,N_33309);
nor U34685 (N_34685,N_32159,N_33211);
or U34686 (N_34686,N_32095,N_33524);
and U34687 (N_34687,N_32707,N_32183);
xor U34688 (N_34688,N_33313,N_32830);
nor U34689 (N_34689,N_33443,N_32930);
nand U34690 (N_34690,N_33006,N_32757);
or U34691 (N_34691,N_32916,N_32878);
or U34692 (N_34692,N_32634,N_32196);
nand U34693 (N_34693,N_32512,N_32246);
xnor U34694 (N_34694,N_33978,N_32547);
or U34695 (N_34695,N_33946,N_33629);
or U34696 (N_34696,N_33420,N_32849);
or U34697 (N_34697,N_32115,N_33214);
nand U34698 (N_34698,N_33127,N_33059);
nand U34699 (N_34699,N_33229,N_32342);
nor U34700 (N_34700,N_33051,N_33367);
xnor U34701 (N_34701,N_33660,N_33115);
nor U34702 (N_34702,N_32789,N_32880);
or U34703 (N_34703,N_33967,N_32104);
or U34704 (N_34704,N_33972,N_33856);
and U34705 (N_34705,N_32717,N_33182);
nand U34706 (N_34706,N_33474,N_32224);
nor U34707 (N_34707,N_33771,N_32419);
nand U34708 (N_34708,N_32477,N_32328);
xnor U34709 (N_34709,N_33342,N_33422);
and U34710 (N_34710,N_32889,N_33200);
nand U34711 (N_34711,N_32838,N_33250);
nor U34712 (N_34712,N_32176,N_32750);
nor U34713 (N_34713,N_33785,N_32401);
nor U34714 (N_34714,N_32693,N_33096);
and U34715 (N_34715,N_32278,N_33655);
and U34716 (N_34716,N_32952,N_32550);
xor U34717 (N_34717,N_33418,N_32004);
xnor U34718 (N_34718,N_33659,N_32052);
nand U34719 (N_34719,N_33607,N_32992);
nor U34720 (N_34720,N_32574,N_33396);
or U34721 (N_34721,N_32345,N_32408);
or U34722 (N_34722,N_33828,N_32743);
nand U34723 (N_34723,N_32821,N_33913);
nor U34724 (N_34724,N_33691,N_32633);
or U34725 (N_34725,N_32060,N_32431);
nor U34726 (N_34726,N_32331,N_32023);
and U34727 (N_34727,N_32795,N_32632);
nor U34728 (N_34728,N_33488,N_32186);
or U34729 (N_34729,N_32363,N_33548);
nor U34730 (N_34730,N_33918,N_33142);
xor U34731 (N_34731,N_32475,N_32909);
xor U34732 (N_34732,N_32527,N_32087);
or U34733 (N_34733,N_32505,N_32372);
and U34734 (N_34734,N_33733,N_33703);
and U34735 (N_34735,N_32530,N_32369);
nor U34736 (N_34736,N_32364,N_33636);
and U34737 (N_34737,N_33888,N_32255);
or U34738 (N_34738,N_33814,N_33129);
nand U34739 (N_34739,N_33562,N_33114);
xor U34740 (N_34740,N_32555,N_32499);
and U34741 (N_34741,N_33372,N_33253);
and U34742 (N_34742,N_33052,N_33408);
or U34743 (N_34743,N_33815,N_32208);
nor U34744 (N_34744,N_33531,N_32283);
and U34745 (N_34745,N_32740,N_32536);
nor U34746 (N_34746,N_33834,N_33711);
nand U34747 (N_34747,N_33222,N_32254);
nor U34748 (N_34748,N_33353,N_33025);
or U34749 (N_34749,N_33484,N_33112);
xnor U34750 (N_34750,N_32522,N_33048);
nand U34751 (N_34751,N_32739,N_32951);
or U34752 (N_34752,N_32980,N_32772);
xor U34753 (N_34753,N_32038,N_33337);
nand U34754 (N_34754,N_32781,N_33938);
xnor U34755 (N_34755,N_32809,N_33922);
or U34756 (N_34756,N_32197,N_32669);
nand U34757 (N_34757,N_32968,N_32687);
xor U34758 (N_34758,N_33360,N_33332);
nor U34759 (N_34759,N_32539,N_32525);
xnor U34760 (N_34760,N_32563,N_32313);
nand U34761 (N_34761,N_33800,N_33010);
or U34762 (N_34762,N_33453,N_32217);
nand U34763 (N_34763,N_32635,N_32076);
nand U34764 (N_34764,N_33879,N_32583);
and U34765 (N_34765,N_32072,N_32565);
nand U34766 (N_34766,N_32798,N_33263);
xnor U34767 (N_34767,N_32958,N_33312);
or U34768 (N_34768,N_33456,N_32922);
xnor U34769 (N_34769,N_33128,N_32680);
nand U34770 (N_34770,N_33085,N_33139);
nand U34771 (N_34771,N_33283,N_32856);
or U34772 (N_34772,N_32971,N_33935);
or U34773 (N_34773,N_33803,N_33007);
or U34774 (N_34774,N_33391,N_32762);
nand U34775 (N_34775,N_33092,N_32329);
nand U34776 (N_34776,N_32558,N_32377);
and U34777 (N_34777,N_33072,N_32005);
nor U34778 (N_34778,N_32236,N_33281);
nor U34779 (N_34779,N_32453,N_32582);
nor U34780 (N_34780,N_33320,N_32445);
and U34781 (N_34781,N_33444,N_32459);
and U34782 (N_34782,N_32179,N_32871);
nor U34783 (N_34783,N_33500,N_32683);
or U34784 (N_34784,N_32030,N_32688);
or U34785 (N_34785,N_33985,N_32279);
and U34786 (N_34786,N_32055,N_32097);
nor U34787 (N_34787,N_33492,N_32948);
or U34788 (N_34788,N_33996,N_33722);
and U34789 (N_34789,N_32405,N_32156);
xnor U34790 (N_34790,N_32099,N_33776);
nand U34791 (N_34791,N_32266,N_33393);
nor U34792 (N_34792,N_32233,N_33101);
nand U34793 (N_34793,N_32940,N_33632);
nand U34794 (N_34794,N_33399,N_32857);
nand U34795 (N_34795,N_33832,N_32828);
xnor U34796 (N_34796,N_33680,N_33503);
nand U34797 (N_34797,N_32370,N_33339);
and U34798 (N_34798,N_32941,N_32120);
or U34799 (N_34799,N_33826,N_32765);
and U34800 (N_34800,N_32252,N_33830);
nand U34801 (N_34801,N_33070,N_33282);
nand U34802 (N_34802,N_32033,N_32924);
xor U34803 (N_34803,N_33363,N_33062);
or U34804 (N_34804,N_32518,N_33327);
and U34805 (N_34805,N_32642,N_32588);
or U34806 (N_34806,N_32676,N_33438);
nor U34807 (N_34807,N_33383,N_32873);
nand U34808 (N_34808,N_33836,N_33887);
or U34809 (N_34809,N_33685,N_32320);
or U34810 (N_34810,N_32066,N_32519);
xnor U34811 (N_34811,N_32832,N_32599);
nand U34812 (N_34812,N_32121,N_32016);
and U34813 (N_34813,N_33661,N_33130);
nor U34814 (N_34814,N_33541,N_33897);
and U34815 (N_34815,N_32990,N_33782);
xnor U34816 (N_34816,N_33338,N_33490);
and U34817 (N_34817,N_33884,N_33618);
xnor U34818 (N_34818,N_33406,N_33594);
xor U34819 (N_34819,N_33734,N_32470);
nand U34820 (N_34820,N_32752,N_32794);
nor U34821 (N_34821,N_33759,N_33259);
nand U34822 (N_34822,N_33564,N_33539);
or U34823 (N_34823,N_33183,N_32917);
and U34824 (N_34824,N_32141,N_33181);
or U34825 (N_34825,N_33582,N_33870);
xnor U34826 (N_34826,N_33357,N_33760);
nor U34827 (N_34827,N_33069,N_33644);
or U34828 (N_34828,N_32394,N_33536);
nand U34829 (N_34829,N_33590,N_33440);
xnor U34830 (N_34830,N_32125,N_32959);
xnor U34831 (N_34831,N_32718,N_32144);
xor U34832 (N_34832,N_33352,N_33088);
and U34833 (N_34833,N_32812,N_32105);
xor U34834 (N_34834,N_33584,N_32595);
or U34835 (N_34835,N_32376,N_32070);
nor U34836 (N_34836,N_32065,N_33501);
or U34837 (N_34837,N_33981,N_33515);
xor U34838 (N_34838,N_33506,N_32915);
nor U34839 (N_34839,N_32495,N_32818);
nor U34840 (N_34840,N_32788,N_33266);
and U34841 (N_34841,N_33542,N_33174);
xor U34842 (N_34842,N_33392,N_32430);
nand U34843 (N_34843,N_32647,N_32117);
nor U34844 (N_34844,N_32274,N_33761);
nor U34845 (N_34845,N_32277,N_33896);
nand U34846 (N_34846,N_33223,N_32180);
nand U34847 (N_34847,N_33964,N_33914);
and U34848 (N_34848,N_33037,N_33933);
and U34849 (N_34849,N_32615,N_32756);
and U34850 (N_34850,N_33927,N_33018);
nand U34851 (N_34851,N_32478,N_32275);
nand U34852 (N_34852,N_33885,N_33448);
nand U34853 (N_34853,N_33899,N_32661);
or U34854 (N_34854,N_33257,N_32720);
xnor U34855 (N_34855,N_33033,N_33031);
nand U34856 (N_34856,N_32484,N_33094);
or U34857 (N_34857,N_33550,N_33827);
and U34858 (N_34858,N_33704,N_33117);
nor U34859 (N_34859,N_32628,N_33318);
nor U34860 (N_34860,N_32859,N_33215);
or U34861 (N_34861,N_33107,N_33580);
and U34862 (N_34862,N_33405,N_33939);
nor U34863 (N_34863,N_33119,N_32061);
or U34864 (N_34864,N_32708,N_33871);
xnor U34865 (N_34865,N_32310,N_33080);
nor U34866 (N_34866,N_32887,N_32265);
nand U34867 (N_34867,N_33831,N_33600);
or U34868 (N_34868,N_33424,N_33319);
or U34869 (N_34869,N_33487,N_33606);
or U34870 (N_34870,N_32840,N_33249);
and U34871 (N_34871,N_32728,N_33022);
nand U34872 (N_34872,N_33801,N_33719);
nand U34873 (N_34873,N_32945,N_33960);
or U34874 (N_34874,N_33196,N_33625);
nand U34875 (N_34875,N_32216,N_33917);
nand U34876 (N_34876,N_32610,N_32425);
nand U34877 (N_34877,N_33558,N_33341);
xor U34878 (N_34878,N_32280,N_33683);
nand U34879 (N_34879,N_33559,N_32640);
nor U34880 (N_34880,N_33730,N_32257);
and U34881 (N_34881,N_33989,N_32737);
nor U34882 (N_34882,N_32476,N_32970);
xor U34883 (N_34883,N_33561,N_33763);
and U34884 (N_34884,N_33858,N_32787);
nand U34885 (N_34885,N_33298,N_33976);
or U34886 (N_34886,N_32551,N_32267);
nor U34887 (N_34887,N_33262,N_32321);
xnor U34888 (N_34888,N_32268,N_33614);
or U34889 (N_34889,N_32114,N_33892);
nand U34890 (N_34890,N_32131,N_32081);
or U34891 (N_34891,N_33848,N_33665);
and U34892 (N_34892,N_33649,N_32645);
xnor U34893 (N_34893,N_32150,N_32624);
and U34894 (N_34894,N_32122,N_32713);
and U34895 (N_34895,N_33791,N_32054);
or U34896 (N_34896,N_32570,N_32041);
nor U34897 (N_34897,N_33251,N_32464);
nand U34898 (N_34898,N_32003,N_33218);
nand U34899 (N_34899,N_33779,N_32837);
or U34900 (N_34900,N_32623,N_33731);
xnor U34901 (N_34901,N_32502,N_32078);
xor U34902 (N_34902,N_33038,N_33705);
nor U34903 (N_34903,N_32910,N_33684);
and U34904 (N_34904,N_32378,N_32034);
nor U34905 (N_34905,N_33898,N_33024);
or U34906 (N_34906,N_33081,N_33049);
or U34907 (N_34907,N_32045,N_32355);
xnor U34908 (N_34908,N_33990,N_32324);
or U34909 (N_34909,N_32009,N_33279);
nand U34910 (N_34910,N_33175,N_33111);
xnor U34911 (N_34911,N_32899,N_33804);
and U34912 (N_34912,N_32085,N_33877);
nand U34913 (N_34913,N_32191,N_33290);
or U34914 (N_34914,N_33821,N_33662);
or U34915 (N_34915,N_33297,N_32964);
or U34916 (N_34916,N_33141,N_33395);
or U34917 (N_34917,N_33151,N_32449);
or U34918 (N_34918,N_32001,N_32049);
or U34919 (N_34919,N_33185,N_32040);
or U34920 (N_34920,N_33213,N_33772);
or U34921 (N_34921,N_33920,N_33188);
xor U34922 (N_34922,N_33762,N_33230);
or U34923 (N_34923,N_33243,N_33032);
xnor U34924 (N_34924,N_33950,N_32678);
nor U34925 (N_34925,N_32008,N_33666);
nand U34926 (N_34926,N_32386,N_33566);
or U34927 (N_34927,N_33807,N_33113);
nand U34928 (N_34928,N_32892,N_32460);
or U34929 (N_34929,N_32938,N_32263);
xnor U34930 (N_34930,N_32872,N_33144);
nor U34931 (N_34931,N_32793,N_33336);
nand U34932 (N_34932,N_33723,N_33145);
and U34933 (N_34933,N_33802,N_32684);
nand U34934 (N_34934,N_33203,N_33773);
nand U34935 (N_34935,N_32333,N_33397);
xnor U34936 (N_34936,N_32853,N_33923);
xor U34937 (N_34937,N_32995,N_32655);
nand U34938 (N_34938,N_33385,N_32492);
or U34939 (N_34939,N_32340,N_32285);
and U34940 (N_34940,N_33758,N_33238);
nor U34941 (N_34941,N_32273,N_33865);
xor U34942 (N_34942,N_32903,N_32334);
nor U34943 (N_34943,N_33143,N_32748);
xor U34944 (N_34944,N_32879,N_33591);
nor U34945 (N_34945,N_33172,N_33648);
and U34946 (N_34946,N_32393,N_32189);
and U34947 (N_34947,N_32075,N_32138);
or U34948 (N_34948,N_33384,N_32380);
and U34949 (N_34949,N_32371,N_32664);
nor U34950 (N_34950,N_32526,N_33931);
or U34951 (N_34951,N_33739,N_32392);
xnor U34952 (N_34952,N_32577,N_33994);
nand U34953 (N_34953,N_32025,N_32942);
nor U34954 (N_34954,N_32988,N_32446);
and U34955 (N_34955,N_32210,N_32579);
nand U34956 (N_34956,N_32561,N_32792);
or U34957 (N_34957,N_33292,N_32103);
or U34958 (N_34958,N_33511,N_32244);
xor U34959 (N_34959,N_33012,N_32531);
nand U34960 (N_34960,N_33164,N_32982);
xor U34961 (N_34961,N_32660,N_32173);
or U34962 (N_34962,N_32855,N_32898);
and U34963 (N_34963,N_33527,N_33626);
xor U34964 (N_34964,N_32067,N_33428);
and U34965 (N_34965,N_32482,N_33167);
or U34966 (N_34966,N_33228,N_32758);
xnor U34967 (N_34967,N_33756,N_33741);
xor U34968 (N_34968,N_32606,N_33854);
xor U34969 (N_34969,N_33133,N_32981);
or U34970 (N_34970,N_33202,N_33516);
nand U34971 (N_34971,N_32307,N_32596);
or U34972 (N_34972,N_32946,N_32844);
or U34973 (N_34973,N_32965,N_32911);
nor U34974 (N_34974,N_32576,N_33421);
xor U34975 (N_34975,N_32053,N_33042);
xor U34976 (N_34976,N_33883,N_33439);
and U34977 (N_34977,N_32424,N_32387);
nand U34978 (N_34978,N_33576,N_32496);
nand U34979 (N_34979,N_33467,N_33971);
nor U34980 (N_34980,N_33494,N_33417);
and U34981 (N_34981,N_33578,N_32084);
and U34982 (N_34982,N_32414,N_32751);
or U34983 (N_34983,N_33686,N_33247);
and U34984 (N_34984,N_33652,N_33104);
and U34985 (N_34985,N_32381,N_32617);
xor U34986 (N_34986,N_33904,N_32537);
and U34987 (N_34987,N_33192,N_32692);
nor U34988 (N_34988,N_32919,N_33082);
nor U34989 (N_34989,N_33495,N_32082);
nor U34990 (N_34990,N_33471,N_32127);
nor U34991 (N_34991,N_32407,N_33179);
or U34992 (N_34992,N_33915,N_32858);
nand U34993 (N_34993,N_33507,N_33951);
xnor U34994 (N_34994,N_32026,N_33159);
or U34995 (N_34995,N_32833,N_33720);
and U34996 (N_34996,N_33679,N_32440);
xnor U34997 (N_34997,N_32149,N_33354);
nand U34998 (N_34998,N_33869,N_33464);
nor U34999 (N_34999,N_32779,N_33653);
xor U35000 (N_35000,N_32093,N_33710);
or U35001 (N_35001,N_33139,N_33728);
and U35002 (N_35002,N_33128,N_32441);
nand U35003 (N_35003,N_32667,N_33958);
nand U35004 (N_35004,N_33047,N_32220);
nor U35005 (N_35005,N_33981,N_33321);
nor U35006 (N_35006,N_33873,N_32004);
and U35007 (N_35007,N_33548,N_32386);
and U35008 (N_35008,N_32593,N_33392);
nor U35009 (N_35009,N_32763,N_32059);
nor U35010 (N_35010,N_32228,N_32662);
nor U35011 (N_35011,N_32451,N_32583);
xnor U35012 (N_35012,N_33334,N_33883);
and U35013 (N_35013,N_32333,N_32642);
xor U35014 (N_35014,N_33306,N_32961);
and U35015 (N_35015,N_32986,N_33540);
nand U35016 (N_35016,N_33667,N_32536);
nor U35017 (N_35017,N_33203,N_32094);
nor U35018 (N_35018,N_32364,N_33278);
xor U35019 (N_35019,N_32252,N_33995);
or U35020 (N_35020,N_32626,N_32288);
or U35021 (N_35021,N_32205,N_32949);
nand U35022 (N_35022,N_33887,N_33743);
nor U35023 (N_35023,N_32890,N_32528);
xor U35024 (N_35024,N_32001,N_32327);
xor U35025 (N_35025,N_33666,N_32042);
nand U35026 (N_35026,N_32693,N_32212);
nand U35027 (N_35027,N_33426,N_32916);
nand U35028 (N_35028,N_32338,N_32884);
nand U35029 (N_35029,N_32864,N_33501);
and U35030 (N_35030,N_32190,N_32050);
nor U35031 (N_35031,N_33687,N_33539);
or U35032 (N_35032,N_32850,N_32307);
xor U35033 (N_35033,N_32570,N_33851);
and U35034 (N_35034,N_33538,N_33913);
or U35035 (N_35035,N_32031,N_33778);
nand U35036 (N_35036,N_32397,N_33789);
nor U35037 (N_35037,N_32070,N_33111);
nor U35038 (N_35038,N_32989,N_32141);
and U35039 (N_35039,N_32245,N_32347);
or U35040 (N_35040,N_33429,N_32650);
nor U35041 (N_35041,N_32356,N_32175);
nand U35042 (N_35042,N_32423,N_33367);
nand U35043 (N_35043,N_32771,N_33623);
or U35044 (N_35044,N_32218,N_33318);
xnor U35045 (N_35045,N_32057,N_32144);
xnor U35046 (N_35046,N_32338,N_33921);
and U35047 (N_35047,N_33990,N_33198);
nand U35048 (N_35048,N_33157,N_32671);
nand U35049 (N_35049,N_32689,N_33316);
nand U35050 (N_35050,N_32622,N_33186);
xor U35051 (N_35051,N_32552,N_32219);
nor U35052 (N_35052,N_33964,N_32334);
or U35053 (N_35053,N_32047,N_33385);
or U35054 (N_35054,N_32836,N_32773);
nand U35055 (N_35055,N_33978,N_32102);
or U35056 (N_35056,N_32711,N_32643);
xnor U35057 (N_35057,N_32052,N_33634);
nand U35058 (N_35058,N_32359,N_32082);
nor U35059 (N_35059,N_32260,N_32685);
or U35060 (N_35060,N_33334,N_32581);
and U35061 (N_35061,N_33393,N_32682);
nor U35062 (N_35062,N_32917,N_33082);
nor U35063 (N_35063,N_32270,N_33647);
nor U35064 (N_35064,N_32243,N_33519);
nand U35065 (N_35065,N_33765,N_33985);
nor U35066 (N_35066,N_32348,N_33950);
or U35067 (N_35067,N_32187,N_32755);
and U35068 (N_35068,N_32502,N_33052);
or U35069 (N_35069,N_32607,N_33966);
nor U35070 (N_35070,N_32066,N_32219);
nor U35071 (N_35071,N_33650,N_33096);
or U35072 (N_35072,N_32905,N_32555);
nand U35073 (N_35073,N_33514,N_33540);
nand U35074 (N_35074,N_33471,N_33027);
nand U35075 (N_35075,N_32064,N_33185);
or U35076 (N_35076,N_33518,N_32296);
xor U35077 (N_35077,N_32951,N_32673);
and U35078 (N_35078,N_33097,N_33675);
nand U35079 (N_35079,N_33094,N_33825);
or U35080 (N_35080,N_32240,N_32245);
or U35081 (N_35081,N_33844,N_33365);
nand U35082 (N_35082,N_33964,N_33468);
nand U35083 (N_35083,N_33997,N_32080);
and U35084 (N_35084,N_32073,N_32566);
nor U35085 (N_35085,N_32814,N_32343);
nor U35086 (N_35086,N_33473,N_32362);
nor U35087 (N_35087,N_32163,N_33703);
nor U35088 (N_35088,N_33493,N_33449);
or U35089 (N_35089,N_32235,N_33815);
and U35090 (N_35090,N_32231,N_33311);
and U35091 (N_35091,N_32371,N_32505);
and U35092 (N_35092,N_32461,N_33514);
nand U35093 (N_35093,N_32097,N_33986);
nor U35094 (N_35094,N_32876,N_33532);
and U35095 (N_35095,N_32414,N_33823);
or U35096 (N_35096,N_32763,N_33307);
and U35097 (N_35097,N_33125,N_33715);
xnor U35098 (N_35098,N_33053,N_33062);
or U35099 (N_35099,N_32339,N_32110);
nand U35100 (N_35100,N_32826,N_33028);
nor U35101 (N_35101,N_32538,N_32366);
xnor U35102 (N_35102,N_33806,N_33419);
or U35103 (N_35103,N_32331,N_33587);
or U35104 (N_35104,N_32758,N_32363);
nor U35105 (N_35105,N_32896,N_32066);
nand U35106 (N_35106,N_32369,N_32171);
nor U35107 (N_35107,N_32434,N_32774);
and U35108 (N_35108,N_33071,N_33567);
and U35109 (N_35109,N_32752,N_32316);
xor U35110 (N_35110,N_33473,N_32918);
nand U35111 (N_35111,N_33429,N_32875);
xor U35112 (N_35112,N_33926,N_32106);
and U35113 (N_35113,N_33057,N_32068);
and U35114 (N_35114,N_33989,N_33229);
nor U35115 (N_35115,N_32113,N_32066);
and U35116 (N_35116,N_33648,N_32330);
and U35117 (N_35117,N_33435,N_33093);
xnor U35118 (N_35118,N_32732,N_33247);
xor U35119 (N_35119,N_32481,N_33252);
or U35120 (N_35120,N_33937,N_33671);
and U35121 (N_35121,N_32690,N_32508);
or U35122 (N_35122,N_32780,N_33616);
xor U35123 (N_35123,N_33541,N_32557);
or U35124 (N_35124,N_33461,N_33265);
and U35125 (N_35125,N_32466,N_33512);
and U35126 (N_35126,N_33764,N_32567);
nand U35127 (N_35127,N_33004,N_32601);
or U35128 (N_35128,N_33960,N_33970);
nand U35129 (N_35129,N_33034,N_32657);
xor U35130 (N_35130,N_33456,N_33458);
and U35131 (N_35131,N_33818,N_32108);
nand U35132 (N_35132,N_32819,N_32604);
or U35133 (N_35133,N_32869,N_33261);
and U35134 (N_35134,N_33583,N_33138);
nor U35135 (N_35135,N_33344,N_33183);
or U35136 (N_35136,N_32444,N_32594);
nor U35137 (N_35137,N_33488,N_32986);
nand U35138 (N_35138,N_32660,N_32298);
and U35139 (N_35139,N_33376,N_32049);
or U35140 (N_35140,N_33406,N_32811);
or U35141 (N_35141,N_33637,N_33704);
or U35142 (N_35142,N_33040,N_33452);
nor U35143 (N_35143,N_32563,N_32845);
or U35144 (N_35144,N_32912,N_32847);
nand U35145 (N_35145,N_32686,N_32647);
xor U35146 (N_35146,N_32525,N_33941);
nor U35147 (N_35147,N_33071,N_33756);
nand U35148 (N_35148,N_32062,N_33002);
nand U35149 (N_35149,N_33399,N_33690);
or U35150 (N_35150,N_32641,N_32377);
nand U35151 (N_35151,N_32113,N_32955);
nand U35152 (N_35152,N_32596,N_32262);
xor U35153 (N_35153,N_33834,N_33329);
xor U35154 (N_35154,N_32916,N_32866);
nand U35155 (N_35155,N_32034,N_32065);
nand U35156 (N_35156,N_33488,N_33318);
nor U35157 (N_35157,N_32186,N_32761);
nor U35158 (N_35158,N_32020,N_33045);
xnor U35159 (N_35159,N_32244,N_33774);
and U35160 (N_35160,N_32189,N_33074);
or U35161 (N_35161,N_32434,N_33552);
nor U35162 (N_35162,N_32183,N_33477);
xor U35163 (N_35163,N_32637,N_32382);
nand U35164 (N_35164,N_33143,N_32762);
nor U35165 (N_35165,N_32983,N_33543);
or U35166 (N_35166,N_33455,N_32239);
xor U35167 (N_35167,N_33895,N_33174);
nor U35168 (N_35168,N_33503,N_33566);
xnor U35169 (N_35169,N_32208,N_32602);
nor U35170 (N_35170,N_33323,N_32928);
or U35171 (N_35171,N_32425,N_33985);
xnor U35172 (N_35172,N_33132,N_32795);
and U35173 (N_35173,N_33689,N_33186);
or U35174 (N_35174,N_32089,N_33688);
nor U35175 (N_35175,N_32265,N_33662);
or U35176 (N_35176,N_33174,N_33282);
nand U35177 (N_35177,N_33013,N_32649);
or U35178 (N_35178,N_33026,N_32294);
xnor U35179 (N_35179,N_32681,N_33272);
or U35180 (N_35180,N_33053,N_33518);
nor U35181 (N_35181,N_33231,N_32742);
and U35182 (N_35182,N_32587,N_33666);
nand U35183 (N_35183,N_32605,N_32436);
or U35184 (N_35184,N_33898,N_33422);
xnor U35185 (N_35185,N_33343,N_32358);
xor U35186 (N_35186,N_32437,N_33595);
and U35187 (N_35187,N_32364,N_32517);
nand U35188 (N_35188,N_33883,N_32776);
and U35189 (N_35189,N_33143,N_33648);
or U35190 (N_35190,N_32648,N_33330);
and U35191 (N_35191,N_33033,N_32750);
xor U35192 (N_35192,N_33728,N_32819);
and U35193 (N_35193,N_32171,N_32860);
and U35194 (N_35194,N_32468,N_32402);
nor U35195 (N_35195,N_32955,N_32286);
nor U35196 (N_35196,N_33686,N_32094);
and U35197 (N_35197,N_33965,N_32151);
xnor U35198 (N_35198,N_33689,N_32940);
xor U35199 (N_35199,N_32905,N_32193);
nand U35200 (N_35200,N_32530,N_33056);
and U35201 (N_35201,N_33868,N_32789);
nand U35202 (N_35202,N_33075,N_33937);
and U35203 (N_35203,N_32074,N_32839);
nand U35204 (N_35204,N_33995,N_33038);
and U35205 (N_35205,N_32490,N_32822);
or U35206 (N_35206,N_32639,N_32090);
nand U35207 (N_35207,N_33432,N_33356);
nor U35208 (N_35208,N_33285,N_32705);
and U35209 (N_35209,N_32716,N_33454);
and U35210 (N_35210,N_32805,N_32070);
xnor U35211 (N_35211,N_33747,N_33283);
and U35212 (N_35212,N_33563,N_33463);
or U35213 (N_35213,N_33812,N_32459);
nand U35214 (N_35214,N_33225,N_33039);
xnor U35215 (N_35215,N_32432,N_32376);
and U35216 (N_35216,N_33516,N_33828);
or U35217 (N_35217,N_33911,N_32817);
nor U35218 (N_35218,N_33884,N_32773);
xnor U35219 (N_35219,N_32287,N_33618);
and U35220 (N_35220,N_32992,N_32802);
nand U35221 (N_35221,N_33914,N_32588);
or U35222 (N_35222,N_32809,N_32683);
or U35223 (N_35223,N_32882,N_33655);
nand U35224 (N_35224,N_32515,N_32817);
nor U35225 (N_35225,N_32465,N_32518);
nor U35226 (N_35226,N_33877,N_33522);
nand U35227 (N_35227,N_32989,N_33213);
or U35228 (N_35228,N_32390,N_33074);
xor U35229 (N_35229,N_32871,N_33477);
and U35230 (N_35230,N_32451,N_32240);
nand U35231 (N_35231,N_33508,N_33886);
and U35232 (N_35232,N_32638,N_32324);
or U35233 (N_35233,N_33669,N_32549);
xor U35234 (N_35234,N_33117,N_32352);
or U35235 (N_35235,N_33940,N_33419);
and U35236 (N_35236,N_33493,N_33163);
xnor U35237 (N_35237,N_32564,N_32021);
and U35238 (N_35238,N_33036,N_33916);
xnor U35239 (N_35239,N_32006,N_32296);
or U35240 (N_35240,N_32481,N_33855);
and U35241 (N_35241,N_32810,N_32530);
nand U35242 (N_35242,N_32718,N_32890);
nand U35243 (N_35243,N_32373,N_32302);
nor U35244 (N_35244,N_32949,N_32345);
nor U35245 (N_35245,N_32852,N_33859);
nor U35246 (N_35246,N_32862,N_33276);
nand U35247 (N_35247,N_32689,N_33769);
and U35248 (N_35248,N_33782,N_32706);
nor U35249 (N_35249,N_33186,N_33708);
nor U35250 (N_35250,N_33788,N_32429);
and U35251 (N_35251,N_32438,N_32598);
nor U35252 (N_35252,N_32258,N_32340);
nand U35253 (N_35253,N_32210,N_32385);
and U35254 (N_35254,N_32829,N_33208);
or U35255 (N_35255,N_32433,N_32695);
nor U35256 (N_35256,N_32622,N_32481);
or U35257 (N_35257,N_33958,N_33323);
and U35258 (N_35258,N_33982,N_32377);
or U35259 (N_35259,N_32321,N_32522);
nand U35260 (N_35260,N_33885,N_33485);
or U35261 (N_35261,N_32592,N_32860);
nor U35262 (N_35262,N_32446,N_33968);
nand U35263 (N_35263,N_33033,N_33769);
nor U35264 (N_35264,N_32417,N_32705);
or U35265 (N_35265,N_33073,N_33262);
nand U35266 (N_35266,N_32106,N_33180);
nand U35267 (N_35267,N_33614,N_33396);
and U35268 (N_35268,N_33079,N_33711);
nor U35269 (N_35269,N_32012,N_33329);
and U35270 (N_35270,N_33912,N_32201);
nor U35271 (N_35271,N_33753,N_32386);
and U35272 (N_35272,N_33853,N_32489);
nor U35273 (N_35273,N_33194,N_32773);
and U35274 (N_35274,N_32316,N_32055);
nor U35275 (N_35275,N_33518,N_32513);
nand U35276 (N_35276,N_32866,N_32037);
and U35277 (N_35277,N_33578,N_32498);
xnor U35278 (N_35278,N_32197,N_32124);
or U35279 (N_35279,N_33894,N_32913);
and U35280 (N_35280,N_33802,N_32571);
nand U35281 (N_35281,N_32118,N_33917);
xor U35282 (N_35282,N_33796,N_33443);
nor U35283 (N_35283,N_33443,N_33738);
or U35284 (N_35284,N_33062,N_32194);
xor U35285 (N_35285,N_32532,N_32838);
nand U35286 (N_35286,N_32000,N_33649);
and U35287 (N_35287,N_32944,N_33992);
or U35288 (N_35288,N_32589,N_32853);
xor U35289 (N_35289,N_32256,N_33428);
and U35290 (N_35290,N_32013,N_33054);
or U35291 (N_35291,N_32024,N_33100);
xnor U35292 (N_35292,N_32198,N_33484);
or U35293 (N_35293,N_33544,N_33926);
or U35294 (N_35294,N_32600,N_32919);
or U35295 (N_35295,N_33165,N_32085);
or U35296 (N_35296,N_33268,N_32153);
or U35297 (N_35297,N_33089,N_32731);
xnor U35298 (N_35298,N_32332,N_32254);
xor U35299 (N_35299,N_32655,N_32014);
nor U35300 (N_35300,N_32162,N_33485);
xnor U35301 (N_35301,N_32980,N_33432);
and U35302 (N_35302,N_33938,N_33882);
nor U35303 (N_35303,N_33760,N_33205);
nand U35304 (N_35304,N_32402,N_32952);
and U35305 (N_35305,N_32490,N_33091);
nor U35306 (N_35306,N_33243,N_33333);
and U35307 (N_35307,N_32660,N_33867);
xor U35308 (N_35308,N_33682,N_33109);
nor U35309 (N_35309,N_32882,N_33476);
nand U35310 (N_35310,N_33175,N_32005);
nor U35311 (N_35311,N_32048,N_33148);
and U35312 (N_35312,N_32190,N_32650);
or U35313 (N_35313,N_33169,N_33381);
or U35314 (N_35314,N_32539,N_33873);
nand U35315 (N_35315,N_33718,N_33213);
nor U35316 (N_35316,N_33131,N_33598);
xor U35317 (N_35317,N_33530,N_33268);
or U35318 (N_35318,N_32144,N_32203);
and U35319 (N_35319,N_32282,N_32872);
and U35320 (N_35320,N_33810,N_33891);
and U35321 (N_35321,N_33250,N_32052);
xnor U35322 (N_35322,N_33617,N_33167);
nor U35323 (N_35323,N_32398,N_32710);
xor U35324 (N_35324,N_32868,N_33255);
nor U35325 (N_35325,N_33087,N_33231);
or U35326 (N_35326,N_33548,N_32876);
nor U35327 (N_35327,N_32957,N_32251);
or U35328 (N_35328,N_32115,N_32067);
nor U35329 (N_35329,N_33156,N_33770);
or U35330 (N_35330,N_32692,N_32495);
and U35331 (N_35331,N_33590,N_33608);
xnor U35332 (N_35332,N_32870,N_32222);
nand U35333 (N_35333,N_32210,N_33168);
nand U35334 (N_35334,N_33936,N_32872);
or U35335 (N_35335,N_33693,N_32105);
nand U35336 (N_35336,N_33818,N_32967);
nor U35337 (N_35337,N_33777,N_32272);
nand U35338 (N_35338,N_33996,N_32652);
or U35339 (N_35339,N_33082,N_33802);
nor U35340 (N_35340,N_33117,N_32636);
nor U35341 (N_35341,N_32773,N_32298);
or U35342 (N_35342,N_32097,N_32929);
xnor U35343 (N_35343,N_33933,N_32865);
xor U35344 (N_35344,N_33211,N_33557);
nand U35345 (N_35345,N_32243,N_32954);
nand U35346 (N_35346,N_32389,N_32290);
xnor U35347 (N_35347,N_33421,N_33489);
or U35348 (N_35348,N_33490,N_32415);
and U35349 (N_35349,N_33253,N_33159);
and U35350 (N_35350,N_32818,N_32825);
nor U35351 (N_35351,N_32669,N_33536);
nand U35352 (N_35352,N_32751,N_33026);
xor U35353 (N_35353,N_32126,N_32394);
or U35354 (N_35354,N_33142,N_32168);
nor U35355 (N_35355,N_33064,N_33412);
or U35356 (N_35356,N_33923,N_33056);
and U35357 (N_35357,N_33770,N_32825);
xnor U35358 (N_35358,N_32521,N_32633);
xnor U35359 (N_35359,N_33491,N_33995);
or U35360 (N_35360,N_33862,N_33129);
xnor U35361 (N_35361,N_32763,N_33899);
and U35362 (N_35362,N_32927,N_32131);
xnor U35363 (N_35363,N_32710,N_32697);
or U35364 (N_35364,N_32911,N_32689);
nor U35365 (N_35365,N_33967,N_33537);
xnor U35366 (N_35366,N_33815,N_32172);
and U35367 (N_35367,N_32226,N_32191);
nor U35368 (N_35368,N_33841,N_32687);
or U35369 (N_35369,N_32693,N_33557);
nor U35370 (N_35370,N_32372,N_33055);
or U35371 (N_35371,N_33508,N_32908);
nor U35372 (N_35372,N_33969,N_33124);
nand U35373 (N_35373,N_32969,N_32810);
nor U35374 (N_35374,N_33575,N_33314);
or U35375 (N_35375,N_32598,N_33010);
or U35376 (N_35376,N_32997,N_32106);
and U35377 (N_35377,N_32860,N_33321);
xnor U35378 (N_35378,N_32783,N_32663);
nand U35379 (N_35379,N_33423,N_32495);
and U35380 (N_35380,N_33862,N_32929);
and U35381 (N_35381,N_32572,N_32542);
xnor U35382 (N_35382,N_32248,N_32364);
and U35383 (N_35383,N_33545,N_33486);
or U35384 (N_35384,N_32941,N_33372);
or U35385 (N_35385,N_33723,N_32343);
xor U35386 (N_35386,N_33609,N_32806);
nor U35387 (N_35387,N_33581,N_33806);
xor U35388 (N_35388,N_32789,N_32451);
or U35389 (N_35389,N_33640,N_32659);
and U35390 (N_35390,N_33892,N_33116);
xnor U35391 (N_35391,N_32364,N_32952);
xnor U35392 (N_35392,N_33306,N_32170);
or U35393 (N_35393,N_32445,N_32132);
nand U35394 (N_35394,N_33841,N_33112);
or U35395 (N_35395,N_33059,N_32253);
and U35396 (N_35396,N_33272,N_33928);
nor U35397 (N_35397,N_32787,N_32251);
xor U35398 (N_35398,N_32275,N_32414);
and U35399 (N_35399,N_32065,N_32599);
nor U35400 (N_35400,N_32509,N_32267);
and U35401 (N_35401,N_32332,N_33797);
or U35402 (N_35402,N_33429,N_32860);
and U35403 (N_35403,N_33885,N_32392);
nand U35404 (N_35404,N_32628,N_32458);
and U35405 (N_35405,N_33713,N_32836);
nand U35406 (N_35406,N_32946,N_32254);
or U35407 (N_35407,N_32416,N_33104);
nand U35408 (N_35408,N_33011,N_33785);
or U35409 (N_35409,N_33019,N_33589);
nand U35410 (N_35410,N_33645,N_32708);
xnor U35411 (N_35411,N_32200,N_32101);
nand U35412 (N_35412,N_33786,N_33618);
nor U35413 (N_35413,N_33894,N_32014);
nor U35414 (N_35414,N_32654,N_32652);
or U35415 (N_35415,N_32589,N_33296);
xor U35416 (N_35416,N_32215,N_33860);
and U35417 (N_35417,N_32741,N_33273);
and U35418 (N_35418,N_33671,N_33429);
nand U35419 (N_35419,N_33180,N_32398);
nand U35420 (N_35420,N_33978,N_32176);
nor U35421 (N_35421,N_32068,N_33229);
nand U35422 (N_35422,N_33291,N_32230);
nor U35423 (N_35423,N_32047,N_32817);
and U35424 (N_35424,N_33868,N_32486);
or U35425 (N_35425,N_33964,N_32736);
nor U35426 (N_35426,N_32877,N_32386);
nor U35427 (N_35427,N_33867,N_33111);
or U35428 (N_35428,N_32114,N_32623);
nor U35429 (N_35429,N_32664,N_32714);
nor U35430 (N_35430,N_32389,N_33460);
nor U35431 (N_35431,N_33737,N_33822);
nor U35432 (N_35432,N_33340,N_33276);
nor U35433 (N_35433,N_33825,N_33863);
or U35434 (N_35434,N_33034,N_33604);
nor U35435 (N_35435,N_33122,N_32446);
nor U35436 (N_35436,N_33631,N_32028);
xor U35437 (N_35437,N_32459,N_33151);
and U35438 (N_35438,N_33597,N_32568);
nand U35439 (N_35439,N_33333,N_32517);
or U35440 (N_35440,N_32734,N_33517);
nor U35441 (N_35441,N_33052,N_32361);
nand U35442 (N_35442,N_32985,N_33703);
nor U35443 (N_35443,N_33715,N_33301);
nor U35444 (N_35444,N_33877,N_33644);
or U35445 (N_35445,N_33805,N_33998);
nor U35446 (N_35446,N_32181,N_32245);
nor U35447 (N_35447,N_33409,N_33388);
and U35448 (N_35448,N_32534,N_33888);
nand U35449 (N_35449,N_33578,N_32523);
and U35450 (N_35450,N_33123,N_32851);
nor U35451 (N_35451,N_32031,N_32024);
or U35452 (N_35452,N_32047,N_33620);
xor U35453 (N_35453,N_33517,N_32684);
and U35454 (N_35454,N_33162,N_32165);
nor U35455 (N_35455,N_33727,N_32389);
nor U35456 (N_35456,N_32884,N_32232);
nor U35457 (N_35457,N_33575,N_32589);
nand U35458 (N_35458,N_32197,N_33758);
nand U35459 (N_35459,N_33816,N_33330);
xnor U35460 (N_35460,N_33873,N_33703);
nor U35461 (N_35461,N_32679,N_33815);
and U35462 (N_35462,N_33174,N_33860);
nand U35463 (N_35463,N_33272,N_33881);
nand U35464 (N_35464,N_33539,N_33020);
and U35465 (N_35465,N_33121,N_32852);
xor U35466 (N_35466,N_32605,N_33551);
or U35467 (N_35467,N_33184,N_33594);
nor U35468 (N_35468,N_32620,N_33549);
xor U35469 (N_35469,N_33474,N_32194);
and U35470 (N_35470,N_32796,N_33966);
nor U35471 (N_35471,N_32269,N_32805);
xnor U35472 (N_35472,N_33042,N_32575);
xnor U35473 (N_35473,N_33633,N_32732);
nand U35474 (N_35474,N_33566,N_32792);
or U35475 (N_35475,N_33406,N_33893);
xnor U35476 (N_35476,N_32941,N_32165);
or U35477 (N_35477,N_32040,N_32831);
or U35478 (N_35478,N_32590,N_32631);
and U35479 (N_35479,N_32334,N_33591);
nor U35480 (N_35480,N_33797,N_32922);
nor U35481 (N_35481,N_32371,N_33998);
and U35482 (N_35482,N_32821,N_32586);
xnor U35483 (N_35483,N_33963,N_33330);
or U35484 (N_35484,N_32790,N_33773);
xor U35485 (N_35485,N_32718,N_33160);
or U35486 (N_35486,N_33430,N_33232);
xor U35487 (N_35487,N_32648,N_32972);
xnor U35488 (N_35488,N_33525,N_33769);
or U35489 (N_35489,N_32893,N_33355);
nor U35490 (N_35490,N_33775,N_33580);
nand U35491 (N_35491,N_33030,N_33446);
or U35492 (N_35492,N_33339,N_32534);
xnor U35493 (N_35493,N_33559,N_32069);
nor U35494 (N_35494,N_32672,N_32431);
nor U35495 (N_35495,N_33560,N_32692);
nand U35496 (N_35496,N_33229,N_32572);
nor U35497 (N_35497,N_32455,N_32231);
nor U35498 (N_35498,N_32908,N_33707);
nor U35499 (N_35499,N_33721,N_32049);
nand U35500 (N_35500,N_33570,N_32452);
xnor U35501 (N_35501,N_32712,N_32750);
nand U35502 (N_35502,N_33644,N_32927);
nand U35503 (N_35503,N_32136,N_32051);
nor U35504 (N_35504,N_32764,N_32156);
and U35505 (N_35505,N_33816,N_32017);
and U35506 (N_35506,N_32225,N_33918);
or U35507 (N_35507,N_32682,N_32199);
and U35508 (N_35508,N_32031,N_32094);
nand U35509 (N_35509,N_33524,N_32878);
nor U35510 (N_35510,N_33902,N_33080);
nand U35511 (N_35511,N_32840,N_32440);
nand U35512 (N_35512,N_32678,N_33687);
xnor U35513 (N_35513,N_33384,N_32523);
and U35514 (N_35514,N_33421,N_32492);
xor U35515 (N_35515,N_32046,N_32893);
and U35516 (N_35516,N_33894,N_32586);
nor U35517 (N_35517,N_33692,N_33814);
nor U35518 (N_35518,N_32739,N_33178);
xor U35519 (N_35519,N_33864,N_33940);
or U35520 (N_35520,N_33387,N_33094);
or U35521 (N_35521,N_32290,N_32908);
and U35522 (N_35522,N_33536,N_32097);
xor U35523 (N_35523,N_33622,N_33449);
and U35524 (N_35524,N_32362,N_32898);
nand U35525 (N_35525,N_32127,N_32697);
xnor U35526 (N_35526,N_32240,N_32904);
nor U35527 (N_35527,N_32058,N_32374);
nand U35528 (N_35528,N_33741,N_32034);
nor U35529 (N_35529,N_32697,N_33801);
nor U35530 (N_35530,N_33531,N_32072);
nor U35531 (N_35531,N_32477,N_33730);
and U35532 (N_35532,N_33569,N_33892);
xor U35533 (N_35533,N_32980,N_32913);
nor U35534 (N_35534,N_33214,N_32453);
nand U35535 (N_35535,N_32869,N_32288);
xor U35536 (N_35536,N_32919,N_32725);
xnor U35537 (N_35537,N_33239,N_32033);
nand U35538 (N_35538,N_32242,N_33680);
or U35539 (N_35539,N_32057,N_33592);
nor U35540 (N_35540,N_32581,N_32293);
or U35541 (N_35541,N_32370,N_33682);
and U35542 (N_35542,N_32346,N_32596);
and U35543 (N_35543,N_32240,N_33807);
or U35544 (N_35544,N_33448,N_32881);
nor U35545 (N_35545,N_33149,N_33936);
and U35546 (N_35546,N_33891,N_32539);
xor U35547 (N_35547,N_33402,N_33783);
and U35548 (N_35548,N_32135,N_32359);
nand U35549 (N_35549,N_32721,N_32415);
nor U35550 (N_35550,N_32706,N_32434);
nor U35551 (N_35551,N_32744,N_33481);
nand U35552 (N_35552,N_32205,N_32959);
or U35553 (N_35553,N_32997,N_33144);
nor U35554 (N_35554,N_32331,N_32851);
or U35555 (N_35555,N_32115,N_33261);
or U35556 (N_35556,N_33345,N_33415);
and U35557 (N_35557,N_33338,N_33656);
nand U35558 (N_35558,N_32490,N_32669);
xnor U35559 (N_35559,N_33023,N_32567);
nand U35560 (N_35560,N_32730,N_33102);
nand U35561 (N_35561,N_33370,N_32846);
nor U35562 (N_35562,N_33120,N_32867);
nor U35563 (N_35563,N_33997,N_32989);
and U35564 (N_35564,N_33898,N_32748);
nor U35565 (N_35565,N_33250,N_32270);
or U35566 (N_35566,N_33072,N_32599);
nor U35567 (N_35567,N_32014,N_32828);
nor U35568 (N_35568,N_33988,N_32946);
nand U35569 (N_35569,N_33856,N_33346);
nand U35570 (N_35570,N_33983,N_33843);
or U35571 (N_35571,N_33257,N_32002);
xnor U35572 (N_35572,N_32462,N_32802);
and U35573 (N_35573,N_32597,N_32937);
xor U35574 (N_35574,N_32147,N_33802);
and U35575 (N_35575,N_32903,N_33689);
nor U35576 (N_35576,N_32052,N_32628);
or U35577 (N_35577,N_33143,N_33821);
nand U35578 (N_35578,N_32573,N_33764);
nand U35579 (N_35579,N_32784,N_32772);
nand U35580 (N_35580,N_32814,N_33480);
and U35581 (N_35581,N_32269,N_33359);
or U35582 (N_35582,N_32917,N_32680);
nand U35583 (N_35583,N_33047,N_32874);
or U35584 (N_35584,N_32618,N_32330);
or U35585 (N_35585,N_33311,N_33489);
or U35586 (N_35586,N_33168,N_33046);
nor U35587 (N_35587,N_32640,N_32094);
nand U35588 (N_35588,N_33023,N_32639);
nand U35589 (N_35589,N_33374,N_32222);
or U35590 (N_35590,N_32312,N_32668);
xnor U35591 (N_35591,N_33587,N_32170);
nor U35592 (N_35592,N_33464,N_33693);
xor U35593 (N_35593,N_32333,N_33812);
or U35594 (N_35594,N_32834,N_33189);
nand U35595 (N_35595,N_32690,N_33631);
xnor U35596 (N_35596,N_32760,N_32025);
and U35597 (N_35597,N_32015,N_32279);
or U35598 (N_35598,N_33932,N_33959);
nand U35599 (N_35599,N_32701,N_33737);
nor U35600 (N_35600,N_32891,N_32859);
nand U35601 (N_35601,N_33057,N_33433);
and U35602 (N_35602,N_32255,N_33995);
nor U35603 (N_35603,N_32559,N_33339);
nand U35604 (N_35604,N_32080,N_33885);
or U35605 (N_35605,N_32274,N_32077);
and U35606 (N_35606,N_32765,N_33186);
nand U35607 (N_35607,N_33831,N_32791);
nor U35608 (N_35608,N_32128,N_32320);
and U35609 (N_35609,N_32539,N_32129);
and U35610 (N_35610,N_33773,N_32315);
xor U35611 (N_35611,N_32597,N_32948);
nor U35612 (N_35612,N_32457,N_32810);
and U35613 (N_35613,N_32367,N_33677);
and U35614 (N_35614,N_32451,N_33372);
and U35615 (N_35615,N_32475,N_32012);
nand U35616 (N_35616,N_33044,N_33483);
xor U35617 (N_35617,N_32524,N_32378);
nand U35618 (N_35618,N_33755,N_32680);
or U35619 (N_35619,N_32371,N_33079);
nor U35620 (N_35620,N_33144,N_33775);
and U35621 (N_35621,N_32124,N_32924);
or U35622 (N_35622,N_33939,N_32908);
or U35623 (N_35623,N_32252,N_32852);
nor U35624 (N_35624,N_32786,N_32904);
nand U35625 (N_35625,N_32771,N_33737);
xor U35626 (N_35626,N_33323,N_32224);
and U35627 (N_35627,N_33735,N_33809);
or U35628 (N_35628,N_33325,N_32364);
nand U35629 (N_35629,N_32856,N_32391);
and U35630 (N_35630,N_32759,N_32882);
xnor U35631 (N_35631,N_32139,N_33819);
or U35632 (N_35632,N_33063,N_32928);
xnor U35633 (N_35633,N_32683,N_33175);
nand U35634 (N_35634,N_32435,N_33416);
xnor U35635 (N_35635,N_32588,N_32424);
nor U35636 (N_35636,N_32671,N_32311);
or U35637 (N_35637,N_32783,N_33294);
and U35638 (N_35638,N_33405,N_33081);
nor U35639 (N_35639,N_32525,N_33768);
nor U35640 (N_35640,N_33419,N_33481);
nand U35641 (N_35641,N_33926,N_32484);
xor U35642 (N_35642,N_33480,N_33594);
or U35643 (N_35643,N_32373,N_32772);
and U35644 (N_35644,N_32518,N_32530);
xor U35645 (N_35645,N_33046,N_33401);
or U35646 (N_35646,N_32621,N_32581);
or U35647 (N_35647,N_33841,N_33715);
or U35648 (N_35648,N_33871,N_32980);
or U35649 (N_35649,N_32673,N_33646);
nand U35650 (N_35650,N_33200,N_33258);
and U35651 (N_35651,N_32337,N_33608);
xor U35652 (N_35652,N_33966,N_32870);
nor U35653 (N_35653,N_33339,N_33513);
nand U35654 (N_35654,N_33916,N_32104);
nor U35655 (N_35655,N_32033,N_32920);
nand U35656 (N_35656,N_32225,N_33497);
nor U35657 (N_35657,N_32872,N_33056);
xnor U35658 (N_35658,N_33638,N_33375);
nand U35659 (N_35659,N_32417,N_32841);
or U35660 (N_35660,N_32288,N_33515);
nand U35661 (N_35661,N_33979,N_32899);
or U35662 (N_35662,N_33128,N_33913);
and U35663 (N_35663,N_33511,N_33540);
or U35664 (N_35664,N_32328,N_33467);
and U35665 (N_35665,N_33418,N_32988);
nand U35666 (N_35666,N_32865,N_32402);
or U35667 (N_35667,N_32435,N_33775);
and U35668 (N_35668,N_32628,N_32686);
xor U35669 (N_35669,N_32127,N_33493);
xnor U35670 (N_35670,N_33356,N_33023);
and U35671 (N_35671,N_32805,N_32144);
xor U35672 (N_35672,N_32704,N_32782);
and U35673 (N_35673,N_32673,N_32239);
and U35674 (N_35674,N_32553,N_33738);
xnor U35675 (N_35675,N_32752,N_32578);
and U35676 (N_35676,N_32963,N_32795);
and U35677 (N_35677,N_33630,N_32635);
nor U35678 (N_35678,N_32161,N_33014);
and U35679 (N_35679,N_33573,N_33678);
and U35680 (N_35680,N_33772,N_32850);
nand U35681 (N_35681,N_32051,N_32633);
nor U35682 (N_35682,N_33819,N_33183);
and U35683 (N_35683,N_32128,N_33376);
xor U35684 (N_35684,N_32871,N_33967);
nor U35685 (N_35685,N_32017,N_32556);
nand U35686 (N_35686,N_33506,N_33736);
and U35687 (N_35687,N_32209,N_32404);
xnor U35688 (N_35688,N_32491,N_32800);
and U35689 (N_35689,N_32634,N_32485);
or U35690 (N_35690,N_33323,N_32569);
or U35691 (N_35691,N_33159,N_33270);
nand U35692 (N_35692,N_32584,N_33413);
and U35693 (N_35693,N_33577,N_32459);
nand U35694 (N_35694,N_33557,N_32202);
nand U35695 (N_35695,N_32064,N_33899);
and U35696 (N_35696,N_33676,N_33215);
nand U35697 (N_35697,N_33552,N_32742);
nor U35698 (N_35698,N_33515,N_32293);
and U35699 (N_35699,N_33111,N_33701);
or U35700 (N_35700,N_33440,N_33909);
xor U35701 (N_35701,N_32009,N_33329);
and U35702 (N_35702,N_33956,N_33659);
and U35703 (N_35703,N_33809,N_32596);
and U35704 (N_35704,N_33164,N_33068);
and U35705 (N_35705,N_33037,N_32464);
nand U35706 (N_35706,N_32157,N_33049);
or U35707 (N_35707,N_33484,N_32328);
nand U35708 (N_35708,N_32198,N_32731);
xnor U35709 (N_35709,N_32023,N_32448);
nand U35710 (N_35710,N_32774,N_32642);
xnor U35711 (N_35711,N_32129,N_33237);
nor U35712 (N_35712,N_32419,N_33234);
and U35713 (N_35713,N_33960,N_32473);
xor U35714 (N_35714,N_33632,N_32809);
nor U35715 (N_35715,N_33130,N_32460);
and U35716 (N_35716,N_33978,N_32990);
nand U35717 (N_35717,N_33497,N_32270);
and U35718 (N_35718,N_32064,N_33441);
nand U35719 (N_35719,N_33370,N_33226);
or U35720 (N_35720,N_32814,N_33905);
and U35721 (N_35721,N_32417,N_33659);
xor U35722 (N_35722,N_32474,N_32399);
or U35723 (N_35723,N_33468,N_33956);
nor U35724 (N_35724,N_33054,N_32776);
or U35725 (N_35725,N_33731,N_33116);
xor U35726 (N_35726,N_33978,N_32262);
nor U35727 (N_35727,N_32254,N_33209);
or U35728 (N_35728,N_33320,N_32192);
xor U35729 (N_35729,N_32032,N_33993);
or U35730 (N_35730,N_33011,N_32463);
or U35731 (N_35731,N_33636,N_32646);
and U35732 (N_35732,N_32722,N_33870);
xor U35733 (N_35733,N_33891,N_32528);
and U35734 (N_35734,N_33563,N_32000);
or U35735 (N_35735,N_33823,N_32421);
xnor U35736 (N_35736,N_33343,N_32991);
and U35737 (N_35737,N_32528,N_32053);
nor U35738 (N_35738,N_33755,N_33810);
and U35739 (N_35739,N_32009,N_32932);
and U35740 (N_35740,N_33842,N_33302);
xor U35741 (N_35741,N_33148,N_32612);
xnor U35742 (N_35742,N_32181,N_32204);
and U35743 (N_35743,N_33903,N_33712);
and U35744 (N_35744,N_32708,N_33112);
or U35745 (N_35745,N_32799,N_33559);
and U35746 (N_35746,N_33415,N_33770);
xor U35747 (N_35747,N_32491,N_32468);
nor U35748 (N_35748,N_33766,N_33338);
and U35749 (N_35749,N_32164,N_33470);
nor U35750 (N_35750,N_33592,N_33280);
nand U35751 (N_35751,N_32389,N_33204);
and U35752 (N_35752,N_33776,N_33274);
and U35753 (N_35753,N_32304,N_33029);
and U35754 (N_35754,N_33705,N_32811);
and U35755 (N_35755,N_32417,N_32582);
nand U35756 (N_35756,N_32841,N_32459);
nand U35757 (N_35757,N_32532,N_33903);
or U35758 (N_35758,N_32656,N_33702);
or U35759 (N_35759,N_33352,N_32747);
nor U35760 (N_35760,N_33226,N_32534);
nand U35761 (N_35761,N_32546,N_32349);
and U35762 (N_35762,N_32020,N_33173);
and U35763 (N_35763,N_33026,N_32985);
nor U35764 (N_35764,N_32812,N_32058);
and U35765 (N_35765,N_33249,N_33044);
or U35766 (N_35766,N_32075,N_33430);
nor U35767 (N_35767,N_32483,N_33093);
nor U35768 (N_35768,N_32440,N_32519);
xor U35769 (N_35769,N_32623,N_33985);
or U35770 (N_35770,N_32190,N_33534);
nand U35771 (N_35771,N_32846,N_33529);
nor U35772 (N_35772,N_33771,N_33322);
and U35773 (N_35773,N_33148,N_33910);
and U35774 (N_35774,N_33941,N_33753);
and U35775 (N_35775,N_32626,N_32153);
or U35776 (N_35776,N_32298,N_33276);
or U35777 (N_35777,N_33922,N_33229);
xnor U35778 (N_35778,N_32592,N_32301);
and U35779 (N_35779,N_33812,N_32348);
or U35780 (N_35780,N_33554,N_32895);
or U35781 (N_35781,N_32020,N_33627);
and U35782 (N_35782,N_33945,N_32071);
nand U35783 (N_35783,N_32812,N_32671);
nor U35784 (N_35784,N_32063,N_33045);
xor U35785 (N_35785,N_33109,N_32252);
nand U35786 (N_35786,N_33090,N_32250);
nand U35787 (N_35787,N_33650,N_33956);
nor U35788 (N_35788,N_32469,N_33309);
or U35789 (N_35789,N_32071,N_33265);
or U35790 (N_35790,N_32350,N_32368);
or U35791 (N_35791,N_32106,N_33655);
nor U35792 (N_35792,N_32424,N_33471);
or U35793 (N_35793,N_32509,N_33212);
nor U35794 (N_35794,N_32215,N_33848);
xor U35795 (N_35795,N_32806,N_33817);
xor U35796 (N_35796,N_32471,N_32042);
or U35797 (N_35797,N_33944,N_32609);
xor U35798 (N_35798,N_32369,N_33484);
xor U35799 (N_35799,N_32782,N_33006);
nand U35800 (N_35800,N_33926,N_33776);
xor U35801 (N_35801,N_33929,N_32822);
or U35802 (N_35802,N_32264,N_32563);
or U35803 (N_35803,N_33133,N_32188);
nand U35804 (N_35804,N_32886,N_32079);
and U35805 (N_35805,N_33623,N_33563);
nor U35806 (N_35806,N_32839,N_32383);
nand U35807 (N_35807,N_32515,N_33713);
and U35808 (N_35808,N_33128,N_32452);
and U35809 (N_35809,N_32295,N_32451);
or U35810 (N_35810,N_32413,N_32792);
or U35811 (N_35811,N_32418,N_32055);
or U35812 (N_35812,N_33478,N_32032);
or U35813 (N_35813,N_32496,N_32998);
and U35814 (N_35814,N_32537,N_32675);
nor U35815 (N_35815,N_32604,N_32107);
and U35816 (N_35816,N_33657,N_33855);
and U35817 (N_35817,N_33385,N_33377);
and U35818 (N_35818,N_32834,N_33045);
and U35819 (N_35819,N_32830,N_33867);
xor U35820 (N_35820,N_33181,N_33030);
or U35821 (N_35821,N_33256,N_33900);
or U35822 (N_35822,N_32807,N_33223);
or U35823 (N_35823,N_32557,N_32141);
nor U35824 (N_35824,N_33850,N_32023);
xnor U35825 (N_35825,N_33344,N_33818);
nand U35826 (N_35826,N_33227,N_32120);
nor U35827 (N_35827,N_32550,N_33515);
or U35828 (N_35828,N_33134,N_33174);
nand U35829 (N_35829,N_32839,N_33708);
xnor U35830 (N_35830,N_32019,N_33168);
or U35831 (N_35831,N_32706,N_33407);
xor U35832 (N_35832,N_32845,N_32191);
or U35833 (N_35833,N_33669,N_33178);
nand U35834 (N_35834,N_33595,N_33312);
xnor U35835 (N_35835,N_33376,N_33307);
nand U35836 (N_35836,N_33464,N_32044);
xnor U35837 (N_35837,N_32293,N_33752);
xor U35838 (N_35838,N_32902,N_32293);
or U35839 (N_35839,N_33850,N_33776);
or U35840 (N_35840,N_33030,N_32378);
nand U35841 (N_35841,N_33120,N_32755);
nand U35842 (N_35842,N_32694,N_32360);
nand U35843 (N_35843,N_33046,N_33841);
xor U35844 (N_35844,N_33597,N_33951);
xnor U35845 (N_35845,N_32718,N_33526);
nor U35846 (N_35846,N_33288,N_32777);
nand U35847 (N_35847,N_32015,N_33122);
and U35848 (N_35848,N_32306,N_32374);
or U35849 (N_35849,N_33954,N_32247);
xnor U35850 (N_35850,N_33035,N_32928);
xnor U35851 (N_35851,N_33365,N_32093);
or U35852 (N_35852,N_32602,N_32681);
nand U35853 (N_35853,N_32759,N_33677);
nand U35854 (N_35854,N_33767,N_33681);
and U35855 (N_35855,N_33917,N_33532);
and U35856 (N_35856,N_33495,N_33958);
nand U35857 (N_35857,N_32640,N_33126);
or U35858 (N_35858,N_33732,N_32617);
xnor U35859 (N_35859,N_32748,N_33041);
xnor U35860 (N_35860,N_32481,N_33269);
nand U35861 (N_35861,N_33219,N_33677);
or U35862 (N_35862,N_32881,N_32315);
nor U35863 (N_35863,N_33439,N_32534);
nand U35864 (N_35864,N_32628,N_33929);
and U35865 (N_35865,N_33160,N_32780);
nand U35866 (N_35866,N_32255,N_32937);
and U35867 (N_35867,N_33265,N_33828);
nor U35868 (N_35868,N_32765,N_32914);
xor U35869 (N_35869,N_33551,N_33789);
or U35870 (N_35870,N_32078,N_32316);
or U35871 (N_35871,N_33125,N_33402);
nor U35872 (N_35872,N_33632,N_33907);
or U35873 (N_35873,N_32654,N_32741);
and U35874 (N_35874,N_33415,N_33842);
or U35875 (N_35875,N_32205,N_33577);
or U35876 (N_35876,N_33296,N_33882);
nand U35877 (N_35877,N_32135,N_33443);
xor U35878 (N_35878,N_33136,N_33903);
or U35879 (N_35879,N_32859,N_33221);
and U35880 (N_35880,N_33094,N_33074);
or U35881 (N_35881,N_32009,N_32948);
or U35882 (N_35882,N_32926,N_33333);
and U35883 (N_35883,N_32301,N_32924);
xnor U35884 (N_35884,N_32376,N_32903);
nand U35885 (N_35885,N_32179,N_32464);
or U35886 (N_35886,N_33186,N_32105);
nor U35887 (N_35887,N_32544,N_32897);
nor U35888 (N_35888,N_32090,N_32935);
xor U35889 (N_35889,N_32725,N_33717);
xnor U35890 (N_35890,N_33245,N_32140);
nor U35891 (N_35891,N_32896,N_32342);
nor U35892 (N_35892,N_32748,N_32677);
nor U35893 (N_35893,N_32937,N_32057);
xor U35894 (N_35894,N_33734,N_33612);
nand U35895 (N_35895,N_32952,N_33274);
or U35896 (N_35896,N_32714,N_33919);
or U35897 (N_35897,N_32699,N_32911);
and U35898 (N_35898,N_32738,N_32711);
nand U35899 (N_35899,N_32414,N_33886);
nor U35900 (N_35900,N_32402,N_33606);
nor U35901 (N_35901,N_32189,N_32372);
nor U35902 (N_35902,N_33595,N_32304);
nand U35903 (N_35903,N_32655,N_32437);
nor U35904 (N_35904,N_32149,N_33507);
and U35905 (N_35905,N_33898,N_32870);
nor U35906 (N_35906,N_33886,N_32394);
nand U35907 (N_35907,N_33997,N_32021);
and U35908 (N_35908,N_33973,N_33344);
xnor U35909 (N_35909,N_33282,N_32750);
nand U35910 (N_35910,N_33573,N_32236);
and U35911 (N_35911,N_32367,N_32478);
nand U35912 (N_35912,N_32253,N_33316);
or U35913 (N_35913,N_32209,N_32939);
and U35914 (N_35914,N_32217,N_33642);
nor U35915 (N_35915,N_32315,N_33103);
nor U35916 (N_35916,N_33109,N_32417);
or U35917 (N_35917,N_32390,N_33067);
nor U35918 (N_35918,N_33549,N_32923);
nand U35919 (N_35919,N_33071,N_32796);
and U35920 (N_35920,N_32845,N_32291);
or U35921 (N_35921,N_33213,N_32836);
xnor U35922 (N_35922,N_33982,N_33659);
or U35923 (N_35923,N_33687,N_32350);
nand U35924 (N_35924,N_33861,N_32027);
nor U35925 (N_35925,N_32277,N_32987);
nor U35926 (N_35926,N_33153,N_32911);
nand U35927 (N_35927,N_32995,N_33383);
xor U35928 (N_35928,N_32371,N_33245);
xnor U35929 (N_35929,N_33763,N_32002);
nand U35930 (N_35930,N_32770,N_32228);
nand U35931 (N_35931,N_32997,N_32203);
nand U35932 (N_35932,N_33852,N_33611);
nor U35933 (N_35933,N_33732,N_32154);
or U35934 (N_35934,N_32025,N_32309);
xnor U35935 (N_35935,N_33082,N_33758);
nand U35936 (N_35936,N_32245,N_33469);
nand U35937 (N_35937,N_32964,N_33289);
and U35938 (N_35938,N_32369,N_33751);
xor U35939 (N_35939,N_32678,N_33413);
and U35940 (N_35940,N_32728,N_32456);
and U35941 (N_35941,N_32373,N_32174);
or U35942 (N_35942,N_32538,N_32334);
and U35943 (N_35943,N_33828,N_32930);
xor U35944 (N_35944,N_32202,N_32658);
or U35945 (N_35945,N_32287,N_32292);
or U35946 (N_35946,N_33912,N_32622);
nand U35947 (N_35947,N_33677,N_32963);
xnor U35948 (N_35948,N_33883,N_32122);
and U35949 (N_35949,N_33427,N_32412);
and U35950 (N_35950,N_33035,N_33987);
xor U35951 (N_35951,N_32329,N_33468);
nand U35952 (N_35952,N_32307,N_33790);
nand U35953 (N_35953,N_33965,N_33116);
and U35954 (N_35954,N_33463,N_33212);
nand U35955 (N_35955,N_32502,N_33004);
nor U35956 (N_35956,N_32474,N_33308);
xnor U35957 (N_35957,N_33251,N_32740);
or U35958 (N_35958,N_32854,N_32196);
and U35959 (N_35959,N_32149,N_32194);
and U35960 (N_35960,N_33980,N_32897);
nand U35961 (N_35961,N_33421,N_33145);
nand U35962 (N_35962,N_32012,N_33599);
or U35963 (N_35963,N_32927,N_33543);
nor U35964 (N_35964,N_32053,N_32469);
or U35965 (N_35965,N_32971,N_32018);
or U35966 (N_35966,N_32944,N_32957);
or U35967 (N_35967,N_32127,N_33095);
and U35968 (N_35968,N_33496,N_33484);
and U35969 (N_35969,N_33730,N_33459);
nor U35970 (N_35970,N_33078,N_32950);
xnor U35971 (N_35971,N_33418,N_33331);
nand U35972 (N_35972,N_32718,N_33987);
nand U35973 (N_35973,N_33629,N_32861);
nand U35974 (N_35974,N_32374,N_32333);
or U35975 (N_35975,N_32853,N_33450);
nor U35976 (N_35976,N_33609,N_33825);
nand U35977 (N_35977,N_32801,N_33583);
nand U35978 (N_35978,N_33221,N_32501);
nand U35979 (N_35979,N_32617,N_33177);
and U35980 (N_35980,N_32555,N_33558);
xnor U35981 (N_35981,N_32034,N_33532);
and U35982 (N_35982,N_32381,N_32469);
or U35983 (N_35983,N_32747,N_33836);
and U35984 (N_35984,N_32633,N_33771);
nor U35985 (N_35985,N_33524,N_32539);
or U35986 (N_35986,N_33836,N_33805);
or U35987 (N_35987,N_33257,N_33231);
nor U35988 (N_35988,N_33927,N_33231);
nor U35989 (N_35989,N_33499,N_33760);
and U35990 (N_35990,N_33799,N_33903);
or U35991 (N_35991,N_33047,N_32586);
nand U35992 (N_35992,N_33070,N_33597);
or U35993 (N_35993,N_33348,N_32559);
and U35994 (N_35994,N_32324,N_32659);
or U35995 (N_35995,N_32281,N_33962);
nor U35996 (N_35996,N_32075,N_33856);
xnor U35997 (N_35997,N_33897,N_33631);
nor U35998 (N_35998,N_32287,N_33274);
and U35999 (N_35999,N_33027,N_32359);
nand U36000 (N_36000,N_34648,N_35400);
or U36001 (N_36001,N_35596,N_34964);
nor U36002 (N_36002,N_34764,N_35185);
nand U36003 (N_36003,N_34567,N_35497);
xnor U36004 (N_36004,N_35052,N_34037);
xor U36005 (N_36005,N_34983,N_35305);
and U36006 (N_36006,N_34313,N_35088);
nor U36007 (N_36007,N_35438,N_35409);
or U36008 (N_36008,N_35462,N_35678);
and U36009 (N_36009,N_34322,N_35294);
and U36010 (N_36010,N_35546,N_34548);
and U36011 (N_36011,N_35973,N_34765);
or U36012 (N_36012,N_34333,N_35529);
nor U36013 (N_36013,N_34463,N_35220);
xor U36014 (N_36014,N_34986,N_35507);
nand U36015 (N_36015,N_35420,N_34763);
or U36016 (N_36016,N_34896,N_34932);
and U36017 (N_36017,N_34453,N_34019);
or U36018 (N_36018,N_35388,N_34677);
or U36019 (N_36019,N_35557,N_35085);
or U36020 (N_36020,N_35058,N_34705);
or U36021 (N_36021,N_34342,N_35740);
or U36022 (N_36022,N_34810,N_34020);
or U36023 (N_36023,N_34717,N_35524);
and U36024 (N_36024,N_34258,N_34743);
nand U36025 (N_36025,N_34572,N_34729);
nand U36026 (N_36026,N_35190,N_34637);
xor U36027 (N_36027,N_34994,N_35592);
xnor U36028 (N_36028,N_35101,N_34674);
or U36029 (N_36029,N_35258,N_35315);
nand U36030 (N_36030,N_35251,N_35750);
xor U36031 (N_36031,N_35960,N_34966);
and U36032 (N_36032,N_34452,N_35635);
and U36033 (N_36033,N_35378,N_35779);
nor U36034 (N_36034,N_35715,N_35205);
and U36035 (N_36035,N_34388,N_35152);
xnor U36036 (N_36036,N_34032,N_34784);
nor U36037 (N_36037,N_34337,N_35633);
or U36038 (N_36038,N_34556,N_34590);
or U36039 (N_36039,N_34828,N_34696);
nand U36040 (N_36040,N_34881,N_35062);
and U36041 (N_36041,N_35769,N_34219);
and U36042 (N_36042,N_34553,N_35381);
or U36043 (N_36043,N_34471,N_35788);
xor U36044 (N_36044,N_35784,N_34106);
or U36045 (N_36045,N_34953,N_35235);
nor U36046 (N_36046,N_34546,N_34175);
or U36047 (N_36047,N_35503,N_34458);
and U36048 (N_36048,N_34312,N_34488);
xor U36049 (N_36049,N_34948,N_34104);
and U36050 (N_36050,N_34554,N_35588);
xnor U36051 (N_36051,N_34397,N_34023);
and U36052 (N_36052,N_35585,N_34703);
and U36053 (N_36053,N_34047,N_35215);
nor U36054 (N_36054,N_35419,N_34326);
and U36055 (N_36055,N_34800,N_34196);
and U36056 (N_36056,N_35299,N_35451);
xor U36057 (N_36057,N_34456,N_34699);
and U36058 (N_36058,N_35214,N_34410);
xnor U36059 (N_36059,N_35760,N_34685);
and U36060 (N_36060,N_35375,N_34787);
nand U36061 (N_36061,N_34592,N_35663);
nand U36062 (N_36062,N_35694,N_35486);
nor U36063 (N_36063,N_34933,N_35125);
xor U36064 (N_36064,N_34922,N_34512);
or U36065 (N_36065,N_35802,N_34670);
or U36066 (N_36066,N_35362,N_34140);
and U36067 (N_36067,N_34498,N_34734);
or U36068 (N_36068,N_35081,N_34441);
and U36069 (N_36069,N_34733,N_34054);
nor U36070 (N_36070,N_34578,N_35852);
nand U36071 (N_36071,N_34520,N_35226);
nor U36072 (N_36072,N_35182,N_34347);
and U36073 (N_36073,N_35035,N_34183);
or U36074 (N_36074,N_34804,N_35680);
xnor U36075 (N_36075,N_35474,N_35997);
and U36076 (N_36076,N_35510,N_35581);
and U36077 (N_36077,N_34508,N_35865);
xor U36078 (N_36078,N_35889,N_35595);
nand U36079 (N_36079,N_34877,N_34164);
and U36080 (N_36080,N_35563,N_35422);
nor U36081 (N_36081,N_34404,N_34930);
nor U36082 (N_36082,N_35897,N_34276);
and U36083 (N_36083,N_35791,N_34036);
nand U36084 (N_36084,N_34976,N_34533);
nand U36085 (N_36085,N_35827,N_35238);
xnor U36086 (N_36086,N_34285,N_34735);
and U36087 (N_36087,N_34888,N_35014);
and U36088 (N_36088,N_35519,N_34781);
nor U36089 (N_36089,N_35533,N_35591);
or U36090 (N_36090,N_35725,N_34786);
xor U36091 (N_36091,N_34096,N_34042);
and U36092 (N_36092,N_35331,N_34942);
nand U36093 (N_36093,N_34331,N_35410);
nor U36094 (N_36094,N_35828,N_35677);
nor U36095 (N_36095,N_34751,N_35751);
and U36096 (N_36096,N_35395,N_34177);
and U36097 (N_36097,N_35180,N_35660);
and U36098 (N_36098,N_34330,N_34667);
nand U36099 (N_36099,N_34737,N_34021);
nor U36100 (N_36100,N_35723,N_34704);
nand U36101 (N_36101,N_35261,N_34460);
nor U36102 (N_36102,N_34367,N_34450);
and U36103 (N_36103,N_34466,N_35326);
or U36104 (N_36104,N_34911,N_35396);
nor U36105 (N_36105,N_34311,N_35033);
and U36106 (N_36106,N_34144,N_34345);
xnor U36107 (N_36107,N_35945,N_35860);
nor U36108 (N_36108,N_35262,N_34358);
and U36109 (N_36109,N_35884,N_34831);
or U36110 (N_36110,N_34133,N_34049);
nand U36111 (N_36111,N_34652,N_34418);
xnor U36112 (N_36112,N_35128,N_35109);
or U36113 (N_36113,N_34755,N_35696);
xor U36114 (N_36114,N_34382,N_35228);
nor U36115 (N_36115,N_35253,N_34341);
and U36116 (N_36116,N_34155,N_35891);
or U36117 (N_36117,N_34295,N_34653);
xor U36118 (N_36118,N_35823,N_35758);
nand U36119 (N_36119,N_35389,N_34635);
nor U36120 (N_36120,N_35864,N_35874);
or U36121 (N_36121,N_35602,N_35808);
xor U36122 (N_36122,N_34875,N_34178);
or U36123 (N_36123,N_34034,N_34259);
nand U36124 (N_36124,N_34139,N_35820);
nor U36125 (N_36125,N_34698,N_34129);
xnor U36126 (N_36126,N_35113,N_35916);
nand U36127 (N_36127,N_35787,N_34009);
and U36128 (N_36128,N_35440,N_35626);
and U36129 (N_36129,N_35755,N_35293);
or U36130 (N_36130,N_34641,N_35314);
nor U36131 (N_36131,N_35263,N_34110);
or U36132 (N_36132,N_34477,N_35645);
nand U36133 (N_36133,N_35684,N_34626);
xnor U36134 (N_36134,N_35862,N_34062);
nor U36135 (N_36135,N_35909,N_34437);
and U36136 (N_36136,N_35877,N_34617);
or U36137 (N_36137,N_34662,N_34281);
and U36138 (N_36138,N_34584,N_34519);
xor U36139 (N_36139,N_34610,N_34203);
and U36140 (N_36140,N_35776,N_34803);
and U36141 (N_36141,N_35708,N_34145);
and U36142 (N_36142,N_35495,N_34072);
or U36143 (N_36143,N_34081,N_35778);
and U36144 (N_36144,N_35225,N_35193);
nor U36145 (N_36145,N_35319,N_35196);
xor U36146 (N_36146,N_34629,N_35350);
nand U36147 (N_36147,N_34883,N_35289);
and U36148 (N_36148,N_35150,N_35277);
xor U36149 (N_36149,N_34604,N_35021);
or U36150 (N_36150,N_35686,N_35295);
xor U36151 (N_36151,N_35579,N_35598);
nand U36152 (N_36152,N_35158,N_34832);
nand U36153 (N_36153,N_34492,N_34304);
nor U36154 (N_36154,N_34736,N_34247);
or U36155 (N_36155,N_34860,N_34642);
nand U36156 (N_36156,N_35670,N_35824);
nand U36157 (N_36157,N_35442,N_34945);
xnor U36158 (N_36158,N_35472,N_34030);
and U36159 (N_36159,N_35298,N_35522);
and U36160 (N_36160,N_35988,N_35011);
and U36161 (N_36161,N_34080,N_35348);
nand U36162 (N_36162,N_34613,N_34811);
and U36163 (N_36163,N_35270,N_35993);
nand U36164 (N_36164,N_35232,N_34473);
xnor U36165 (N_36165,N_35071,N_34306);
or U36166 (N_36166,N_35357,N_35108);
or U36167 (N_36167,N_35646,N_34130);
and U36168 (N_36168,N_35325,N_34856);
or U36169 (N_36169,N_34754,N_35673);
and U36170 (N_36170,N_35681,N_35167);
or U36171 (N_36171,N_34076,N_35873);
or U36172 (N_36172,N_34791,N_35500);
or U36173 (N_36173,N_34507,N_35516);
xnor U36174 (N_36174,N_34099,N_34305);
nor U36175 (N_36175,N_34914,N_34093);
nor U36176 (N_36176,N_34277,N_34224);
nand U36177 (N_36177,N_35590,N_35838);
nor U36178 (N_36178,N_35614,N_34833);
and U36179 (N_36179,N_35955,N_34000);
nor U36180 (N_36180,N_34965,N_35609);
nand U36181 (N_36181,N_35918,N_34152);
or U36182 (N_36182,N_35944,N_34317);
or U36183 (N_36183,N_35363,N_34424);
or U36184 (N_36184,N_35795,N_35335);
and U36185 (N_36185,N_35344,N_34264);
xor U36186 (N_36186,N_34121,N_34708);
and U36187 (N_36187,N_34728,N_34352);
and U36188 (N_36188,N_35432,N_35297);
nor U36189 (N_36189,N_34639,N_35127);
nand U36190 (N_36190,N_35327,N_34402);
nor U36191 (N_36191,N_35735,N_34647);
and U36192 (N_36192,N_34527,N_35364);
and U36193 (N_36193,N_35743,N_35722);
nor U36194 (N_36194,N_34475,N_35094);
and U36195 (N_36195,N_35459,N_35867);
and U36196 (N_36196,N_35179,N_34055);
and U36197 (N_36197,N_35580,N_34461);
nor U36198 (N_36198,N_35761,N_34638);
nor U36199 (N_36199,N_34069,N_34627);
xor U36200 (N_36200,N_35981,N_35953);
nand U36201 (N_36201,N_34753,N_34748);
or U36202 (N_36202,N_35834,N_34620);
nand U36203 (N_36203,N_35488,N_34057);
or U36204 (N_36204,N_34371,N_35360);
xnor U36205 (N_36205,N_35672,N_34017);
xnor U36206 (N_36206,N_35917,N_34960);
nand U36207 (N_36207,N_34661,N_34270);
and U36208 (N_36208,N_34513,N_35817);
nand U36209 (N_36209,N_34222,N_35512);
xor U36210 (N_36210,N_35754,N_35281);
or U36211 (N_36211,N_35106,N_34039);
nor U36212 (N_36212,N_35688,N_35222);
and U36213 (N_36213,N_34510,N_34906);
xnor U36214 (N_36214,N_35339,N_34166);
xor U36215 (N_36215,N_35114,N_34937);
nand U36216 (N_36216,N_35923,N_35699);
or U36217 (N_36217,N_35217,N_35068);
nor U36218 (N_36218,N_35998,N_35501);
xnor U36219 (N_36219,N_34710,N_35324);
nor U36220 (N_36220,N_35009,N_34760);
and U36221 (N_36221,N_34016,N_34444);
nor U36222 (N_36222,N_35799,N_35970);
nor U36223 (N_36223,N_34060,N_34842);
and U36224 (N_36224,N_35629,N_34043);
xor U36225 (N_36225,N_34122,N_34141);
xnor U36226 (N_36226,N_35538,N_35583);
and U36227 (N_36227,N_35139,N_34289);
or U36228 (N_36228,N_34795,N_34793);
and U36229 (N_36229,N_35412,N_34845);
nor U36230 (N_36230,N_34103,N_34749);
or U36231 (N_36231,N_35866,N_34984);
nand U36232 (N_36232,N_34923,N_35078);
or U36233 (N_36233,N_34757,N_34282);
and U36234 (N_36234,N_34562,N_35695);
nand U36235 (N_36235,N_35890,N_35551);
nor U36236 (N_36236,N_35941,N_34014);
or U36237 (N_36237,N_34235,N_35702);
nor U36238 (N_36238,N_35482,N_34600);
nand U36239 (N_36239,N_34242,N_34090);
and U36240 (N_36240,N_35285,N_34445);
nand U36241 (N_36241,N_35968,N_34361);
and U36242 (N_36242,N_34830,N_34809);
nand U36243 (N_36243,N_34100,N_34744);
nor U36244 (N_36244,N_35887,N_34821);
and U36245 (N_36245,N_34303,N_35625);
xor U36246 (N_36246,N_35387,N_35355);
and U36247 (N_36247,N_35804,N_34421);
or U36248 (N_36248,N_35184,N_35816);
xor U36249 (N_36249,N_34192,N_34650);
nand U36250 (N_36250,N_34374,N_35521);
or U36251 (N_36251,N_35570,N_34292);
nand U36252 (N_36252,N_34197,N_34890);
xor U36253 (N_36253,N_35553,N_34563);
or U36254 (N_36254,N_35161,N_35675);
or U36255 (N_36255,N_34329,N_34940);
xnor U36256 (N_36256,N_34115,N_35640);
xnor U36257 (N_36257,N_35697,N_35328);
or U36258 (N_36258,N_34646,N_34633);
nor U36259 (N_36259,N_34084,N_35757);
and U36260 (N_36260,N_34171,N_34243);
nand U36261 (N_36261,N_35736,N_35771);
nand U36262 (N_36262,N_34357,N_35075);
nor U36263 (N_36263,N_35634,N_35064);
nor U36264 (N_36264,N_35532,N_34593);
xnor U36265 (N_36265,N_35465,N_35980);
nor U36266 (N_36266,N_34162,N_34676);
nand U36267 (N_36267,N_34978,N_34262);
xnor U36268 (N_36268,N_34112,N_35407);
xor U36269 (N_36269,N_34683,N_35790);
and U36270 (N_36270,N_35651,N_34871);
nor U36271 (N_36271,N_35434,N_35863);
xnor U36272 (N_36272,N_35067,N_34271);
nand U36273 (N_36273,N_34370,N_34430);
xnor U36274 (N_36274,N_35099,N_34193);
nor U36275 (N_36275,N_34490,N_35045);
and U36276 (N_36276,N_35894,N_34949);
nand U36277 (N_36277,N_35227,N_34070);
nor U36278 (N_36278,N_34143,N_34124);
or U36279 (N_36279,N_35025,N_34383);
nand U36280 (N_36280,N_34480,N_34887);
nand U36281 (N_36281,N_35711,N_35798);
and U36282 (N_36282,N_34428,N_35662);
nor U36283 (N_36283,N_34714,N_35069);
and U36284 (N_36284,N_34256,N_35001);
or U36285 (N_36285,N_34866,N_34476);
and U36286 (N_36286,N_34973,N_35470);
xnor U36287 (N_36287,N_34941,N_35812);
and U36288 (N_36288,N_35514,N_35447);
nor U36289 (N_36289,N_34582,N_34869);
nor U36290 (N_36290,N_35936,N_35077);
nand U36291 (N_36291,N_34335,N_34997);
or U36292 (N_36292,N_34950,N_35922);
and U36293 (N_36293,N_35995,N_35034);
nor U36294 (N_36294,N_35908,N_35053);
xnor U36295 (N_36295,N_34979,N_35931);
nor U36296 (N_36296,N_34411,N_34649);
and U36297 (N_36297,N_35836,N_35130);
xnor U36298 (N_36298,N_34939,N_35212);
nand U36299 (N_36299,N_35174,N_34408);
nor U36300 (N_36300,N_35188,N_35103);
and U36301 (N_36301,N_35240,N_35073);
or U36302 (N_36302,N_34798,N_34643);
nand U36303 (N_36303,N_35347,N_35548);
nor U36304 (N_36304,N_35621,N_35803);
nand U36305 (N_36305,N_34403,N_34449);
nor U36306 (N_36306,N_34568,N_35175);
or U36307 (N_36307,N_34154,N_35173);
or U36308 (N_36308,N_34560,N_34198);
and U36309 (N_36309,N_35368,N_35655);
nand U36310 (N_36310,N_35132,N_34829);
nor U36311 (N_36311,N_34697,N_35429);
nor U36312 (N_36312,N_34241,N_35397);
xnor U36313 (N_36313,N_35008,N_35239);
nand U36314 (N_36314,N_34495,N_34390);
nand U36315 (N_36315,N_34136,N_35272);
nor U36316 (N_36316,N_35421,N_34012);
or U36317 (N_36317,N_34426,N_35230);
nor U36318 (N_36318,N_35578,N_35561);
xor U36319 (N_36319,N_35833,N_35839);
and U36320 (N_36320,N_35845,N_34360);
nor U36321 (N_36321,N_34961,N_35079);
xnor U36322 (N_36322,N_35142,N_35479);
and U36323 (N_36323,N_35138,N_35775);
xnor U36324 (N_36324,N_35136,N_35898);
and U36325 (N_36325,N_35747,N_34489);
or U36326 (N_36326,N_34579,N_35408);
or U36327 (N_36327,N_34559,N_34951);
or U36328 (N_36328,N_34327,N_34204);
or U36329 (N_36329,N_34891,N_34297);
nor U36330 (N_36330,N_34314,N_34954);
and U36331 (N_36331,N_34700,N_35907);
nand U36332 (N_36332,N_34834,N_35030);
nand U36333 (N_36333,N_34501,N_34974);
xnor U36334 (N_36334,N_34551,N_34990);
nor U36335 (N_36335,N_35942,N_35712);
and U36336 (N_36336,N_35171,N_35985);
xnor U36337 (N_36337,N_35206,N_35455);
nor U36338 (N_36338,N_35781,N_35559);
or U36339 (N_36339,N_34485,N_35991);
nand U36340 (N_36340,N_34325,N_34011);
and U36341 (N_36341,N_34213,N_35573);
nor U36342 (N_36342,N_35155,N_35117);
nor U36343 (N_36343,N_35544,N_35216);
nand U36344 (N_36344,N_34414,N_34509);
xnor U36345 (N_36345,N_34415,N_35458);
nand U36346 (N_36346,N_34541,N_35032);
nand U36347 (N_36347,N_35252,N_34656);
nor U36348 (N_36348,N_35246,N_35401);
or U36349 (N_36349,N_34826,N_34472);
and U36350 (N_36350,N_35745,N_35149);
xor U36351 (N_36351,N_35168,N_35906);
and U36352 (N_36352,N_35320,N_35160);
and U36353 (N_36353,N_34599,N_35354);
or U36354 (N_36354,N_34678,N_35192);
xor U36355 (N_36355,N_35371,N_35962);
nand U36356 (N_36356,N_35610,N_34251);
or U36357 (N_36357,N_35657,N_35929);
nand U36358 (N_36358,N_35255,N_35382);
or U36359 (N_36359,N_35237,N_34398);
and U36360 (N_36360,N_34928,N_34724);
nand U36361 (N_36361,N_34234,N_34622);
and U36362 (N_36362,N_34601,N_34220);
xor U36363 (N_36363,N_34240,N_35229);
nand U36364 (N_36364,N_34332,N_34064);
xnor U36365 (N_36365,N_35433,N_34246);
or U36366 (N_36366,N_35316,N_34847);
or U36367 (N_36367,N_35893,N_34199);
and U36368 (N_36368,N_35153,N_34176);
xnor U36369 (N_36369,N_34514,N_35207);
nand U36370 (N_36370,N_34655,N_34716);
nand U36371 (N_36371,N_35676,N_34301);
nand U36372 (N_36372,N_35974,N_35063);
or U36373 (N_36373,N_35949,N_34134);
nor U36374 (N_36374,N_34995,N_34401);
xor U36375 (N_36375,N_34651,N_35770);
and U36376 (N_36376,N_35080,N_35477);
nor U36377 (N_36377,N_34713,N_34058);
and U36378 (N_36378,N_34557,N_35273);
nand U36379 (N_36379,N_34442,N_35183);
nor U36380 (N_36380,N_34063,N_34722);
or U36381 (N_36381,N_34107,N_34521);
nor U36382 (N_36382,N_34693,N_34399);
nand U36383 (N_36383,N_34419,N_34434);
nand U36384 (N_36384,N_34392,N_34201);
xnor U36385 (N_36385,N_35964,N_35526);
or U36386 (N_36386,N_34001,N_34355);
xor U36387 (N_36387,N_35056,N_34102);
or U36388 (N_36388,N_34469,N_34863);
nor U36389 (N_36389,N_34307,N_35313);
nand U36390 (N_36390,N_34543,N_34494);
nor U36391 (N_36391,N_35369,N_35878);
nor U36392 (N_36392,N_34943,N_34912);
nand U36393 (N_36393,N_34252,N_35480);
nand U36394 (N_36394,N_35826,N_34537);
xnor U36395 (N_36395,N_34669,N_34539);
xnor U36396 (N_36396,N_35709,N_34846);
nor U36397 (N_36397,N_34815,N_35248);
and U36398 (N_36398,N_34413,N_35885);
xnor U36399 (N_36399,N_35539,N_35679);
or U36400 (N_36400,N_35612,N_34587);
and U36401 (N_36401,N_35797,N_35210);
xor U36402 (N_36402,N_35569,N_35841);
nand U36403 (N_36403,N_35242,N_34179);
or U36404 (N_36404,N_35652,N_35484);
xor U36405 (N_36405,N_34756,N_34731);
nor U36406 (N_36406,N_34095,N_35938);
xnor U36407 (N_36407,N_35850,N_35200);
and U36408 (N_36408,N_35528,N_34464);
and U36409 (N_36409,N_35530,N_35622);
xor U36410 (N_36410,N_35039,N_35300);
or U36411 (N_36411,N_34812,N_35947);
xnor U36412 (N_36412,N_35649,N_34206);
or U36413 (N_36413,N_34901,N_35698);
nor U36414 (N_36414,N_34935,N_35241);
nor U36415 (N_36415,N_34594,N_35456);
xnor U36416 (N_36416,N_34571,N_34376);
nor U36417 (N_36417,N_35624,N_35431);
or U36418 (N_36418,N_34770,N_35815);
xnor U36419 (N_36419,N_35840,N_34819);
nor U36420 (N_36420,N_35303,N_35233);
or U36421 (N_36421,N_35416,N_35567);
nand U36422 (N_36422,N_34718,N_34873);
nor U36423 (N_36423,N_35613,N_34137);
nor U36424 (N_36424,N_34147,N_35558);
or U36425 (N_36425,N_34169,N_35372);
nand U36426 (N_36426,N_35279,N_35140);
xor U36427 (N_36427,N_35854,N_35247);
xnor U36428 (N_36428,N_35888,N_35107);
xnor U36429 (N_36429,N_34422,N_35449);
or U36430 (N_36430,N_35444,N_34393);
xor U36431 (N_36431,N_35910,N_34186);
nand U36432 (N_36432,N_34522,N_34221);
xor U36433 (N_36433,N_35425,N_35837);
and U36434 (N_36434,N_35017,N_35026);
and U36435 (N_36435,N_34423,N_34237);
or U36436 (N_36436,N_35724,N_35478);
nand U36437 (N_36437,N_34944,N_35793);
nand U36438 (N_36438,N_34853,N_34366);
xor U36439 (N_36439,N_35386,N_34050);
nor U36440 (N_36440,N_34151,N_34644);
and U36441 (N_36441,N_35284,N_35915);
or U36442 (N_36442,N_35911,N_34657);
or U36443 (N_36443,N_34381,N_35648);
nand U36444 (N_36444,N_35163,N_34852);
nand U36445 (N_36445,N_34900,N_34859);
nand U36446 (N_36446,N_34205,N_35700);
xor U36447 (N_36447,N_35730,N_35912);
nand U36448 (N_36448,N_34921,N_35036);
xnor U36449 (N_36449,N_34324,N_35738);
nor U36450 (N_36450,N_35647,N_34172);
nand U36451 (N_36451,N_34672,N_34542);
nand U36452 (N_36452,N_34766,N_34577);
nand U36453 (N_36453,N_35047,N_34597);
nor U36454 (N_36454,N_34052,N_35666);
or U36455 (N_36455,N_34336,N_35346);
xor U36456 (N_36456,N_34958,N_34328);
nor U36457 (N_36457,N_34854,N_34068);
or U36458 (N_36458,N_35871,N_35552);
nor U36459 (N_36459,N_35269,N_35411);
and U36460 (N_36460,N_35091,N_35329);
nand U36461 (N_36461,N_34807,N_35321);
and U36462 (N_36462,N_35302,N_35903);
nor U36463 (N_36463,N_35201,N_34132);
nor U36464 (N_36464,N_34455,N_35020);
nand U36465 (N_36465,N_34632,N_35721);
nand U36466 (N_36466,N_35619,N_35731);
or U36467 (N_36467,N_35244,N_34071);
xor U36468 (N_36468,N_35705,N_34759);
nor U36469 (N_36469,N_34163,N_34822);
and U36470 (N_36470,N_35013,N_35366);
and U36471 (N_36471,N_35291,N_35822);
nand U36472 (N_36472,N_34530,N_35924);
and U36473 (N_36473,N_35979,N_35084);
nor U36474 (N_36474,N_34980,N_34797);
xnor U36475 (N_36475,N_34913,N_35134);
and U36476 (N_36476,N_34138,N_34255);
and U36477 (N_36477,N_34712,N_34602);
xnor U36478 (N_36478,N_34308,N_34167);
xor U36479 (N_36479,N_34216,N_35197);
and U36480 (N_36480,N_34992,N_35115);
xor U36481 (N_36481,N_34780,N_35531);
or U36482 (N_36482,N_35390,N_34775);
nand U36483 (N_36483,N_34681,N_35617);
nor U36484 (N_36484,N_34315,N_34908);
xnor U36485 (N_36485,N_34257,N_34882);
and U36486 (N_36486,N_34515,N_34684);
xnor U36487 (N_36487,N_35496,N_35905);
nor U36488 (N_36488,N_34265,N_35102);
and U36489 (N_36489,N_34695,N_35306);
and U36490 (N_36490,N_34555,N_35453);
and U36491 (N_36491,N_35654,N_34767);
or U36492 (N_36492,N_35266,N_35511);
and U36493 (N_36493,N_34396,N_34185);
or U36494 (N_36494,N_34391,N_34209);
nand U36495 (N_36495,N_34769,N_34805);
xnor U36496 (N_36496,N_35967,N_34349);
nor U36497 (N_36497,N_35351,N_34570);
and U36498 (N_36498,N_34416,N_35166);
nand U36499 (N_36499,N_34073,N_35601);
xor U36500 (N_36500,N_35664,N_34660);
and U36501 (N_36501,N_35151,N_34654);
and U36502 (N_36502,N_34245,N_35370);
nor U36503 (N_36503,N_34719,N_35847);
and U36504 (N_36504,N_35975,N_35643);
or U36505 (N_36505,N_34300,N_35628);
xor U36506 (N_36506,N_35318,N_34474);
and U36507 (N_36507,N_34006,N_35504);
nand U36508 (N_36508,N_34915,N_34931);
and U36509 (N_36509,N_35983,N_35323);
nand U36510 (N_36510,N_34895,N_35880);
nor U36511 (N_36511,N_35394,N_34825);
nor U36512 (N_36512,N_35701,N_35704);
nand U36513 (N_36513,N_35104,N_35857);
and U36514 (N_36514,N_34534,N_34086);
nand U36515 (N_36515,N_35756,N_34702);
nor U36516 (N_36516,N_35037,N_34094);
xnor U36517 (N_36517,N_35861,N_34861);
and U36518 (N_36518,N_34864,N_35719);
and U36519 (N_36519,N_35801,N_34850);
or U36520 (N_36520,N_34056,N_34975);
and U36521 (N_36521,N_35460,N_34123);
or U36522 (N_36522,N_34365,N_35288);
nor U36523 (N_36523,N_35987,N_35982);
nand U36524 (N_36524,N_34293,N_34448);
nand U36525 (N_36525,N_35683,N_34212);
xor U36526 (N_36526,N_34015,N_34666);
xnor U36527 (N_36527,N_34027,N_34529);
and U36528 (N_36528,N_35566,N_35165);
nor U36529 (N_36529,N_35195,N_34738);
or U36530 (N_36530,N_34377,N_34260);
nand U36531 (N_36531,N_34089,N_35956);
nor U36532 (N_36532,N_34814,N_35830);
nor U36533 (N_36533,N_34035,N_34857);
nand U36534 (N_36534,N_35574,N_35727);
xnor U36535 (N_36535,N_35012,N_35004);
nand U36536 (N_36536,N_35920,N_34581);
or U36537 (N_36537,N_34506,N_34528);
xor U36538 (N_36538,N_34188,N_35402);
nand U36539 (N_36539,N_34231,N_35976);
nand U36540 (N_36540,N_35439,N_35869);
or U36541 (N_36541,N_35594,N_34761);
nor U36542 (N_36542,N_35659,N_35336);
or U36543 (N_36543,N_35403,N_35523);
and U36544 (N_36544,N_35349,N_35586);
xnor U36545 (N_36545,N_34002,N_35707);
nand U36546 (N_36546,N_35571,N_34927);
nor U36547 (N_36547,N_34824,N_35028);
nand U36548 (N_36548,N_35135,N_34083);
and U36549 (N_36549,N_35882,N_34715);
nand U36550 (N_36550,N_34364,N_34772);
nand U36551 (N_36551,N_34664,N_35280);
and U36552 (N_36552,N_35786,N_35886);
or U36553 (N_36553,N_34195,N_35413);
nor U36554 (N_36554,N_35219,N_35148);
nor U36555 (N_36555,N_34752,N_34631);
nand U36556 (N_36556,N_34372,N_35513);
nand U36557 (N_36557,N_35714,N_34454);
nor U36558 (N_36558,N_34851,N_34777);
nor U36559 (N_36559,N_34689,N_35667);
and U36560 (N_36560,N_34905,N_34972);
or U36561 (N_36561,N_35599,N_34160);
nor U36562 (N_36562,N_35469,N_35876);
nor U36563 (N_36563,N_34538,N_35630);
and U36564 (N_36564,N_35054,N_35352);
and U36565 (N_36565,N_34827,N_34343);
nand U36566 (N_36566,N_34645,N_35928);
and U36567 (N_36567,N_35050,N_34779);
nand U36568 (N_36568,N_34079,N_34947);
and U36569 (N_36569,N_35418,N_35729);
or U36570 (N_36570,N_35508,N_35007);
nand U36571 (N_36571,N_35549,N_34128);
xnor U36572 (N_36572,N_34701,N_35848);
and U36573 (N_36573,N_34707,N_35129);
or U36574 (N_36574,N_35322,N_35384);
and U36575 (N_36575,N_35070,N_34692);
xor U36576 (N_36576,N_34623,N_35061);
or U36577 (N_36577,N_35204,N_35112);
nor U36578 (N_36578,N_35527,N_35464);
and U36579 (N_36579,N_35773,N_34286);
nand U36580 (N_36580,N_35098,N_34608);
nand U36581 (N_36581,N_34720,N_34573);
and U36582 (N_36582,N_34566,N_34158);
nor U36583 (N_36583,N_35520,N_35023);
nand U36584 (N_36584,N_34742,N_35883);
or U36585 (N_36585,N_34173,N_34118);
and U36586 (N_36586,N_35445,N_34855);
xor U36587 (N_36587,N_35074,N_34886);
and U36588 (N_36588,N_35800,N_34182);
and U36589 (N_36589,N_35691,N_35948);
xnor U36590 (N_36590,N_34161,N_35391);
and U36591 (N_36591,N_34278,N_34959);
and U36592 (N_36592,N_34603,N_35337);
and U36593 (N_36593,N_34621,N_35900);
or U36594 (N_36594,N_34338,N_35046);
or U36595 (N_36595,N_34493,N_35042);
or U36596 (N_36596,N_35608,N_35202);
xnor U36597 (N_36597,N_35308,N_35441);
and U36598 (N_36598,N_35385,N_34727);
nor U36599 (N_36599,N_34740,N_35287);
and U36600 (N_36600,N_34074,N_35491);
or U36601 (N_36601,N_35427,N_34502);
and U36602 (N_36602,N_34516,N_34799);
or U36603 (N_36603,N_35952,N_35674);
nor U36604 (N_36604,N_34082,N_34504);
nand U36605 (N_36605,N_35271,N_34993);
nand U36606 (N_36606,N_34598,N_35868);
xor U36607 (N_36607,N_35537,N_35066);
or U36608 (N_36608,N_34936,N_35164);
nand U36609 (N_36609,N_35243,N_34503);
nor U36610 (N_36610,N_34569,N_35525);
and U36611 (N_36611,N_34202,N_35606);
nand U36612 (N_36612,N_35093,N_34899);
nor U36613 (N_36613,N_35428,N_35343);
nor U36614 (N_36614,N_35072,N_35198);
or U36615 (N_36615,N_34535,N_35254);
or U36616 (N_36616,N_34839,N_35710);
xnor U36617 (N_36617,N_35809,N_34823);
xor U36618 (N_36618,N_34575,N_34375);
nand U36619 (N_36619,N_35296,N_34200);
nand U36620 (N_36620,N_34668,N_35119);
and U36621 (N_36621,N_34524,N_34065);
or U36622 (N_36622,N_35746,N_34321);
nand U36623 (N_36623,N_35003,N_34368);
or U36624 (N_36624,N_35006,N_35417);
or U36625 (N_36625,N_34889,N_34564);
nor U36626 (N_36626,N_34412,N_35641);
nor U36627 (N_36627,N_34619,N_35940);
nor U36628 (N_36628,N_34606,N_34773);
xnor U36629 (N_36629,N_35485,N_34790);
nor U36630 (N_36630,N_35703,N_34232);
and U36631 (N_36631,N_34098,N_35310);
nand U36632 (N_36632,N_35250,N_34117);
or U36633 (N_36633,N_35095,N_34999);
xnor U36634 (N_36634,N_34898,N_35116);
xnor U36635 (N_36635,N_34725,N_35065);
nand U36636 (N_36636,N_34148,N_34214);
and U36637 (N_36637,N_35493,N_35002);
and U36638 (N_36638,N_35489,N_35554);
and U36639 (N_36639,N_35260,N_34005);
nand U36640 (N_36640,N_34496,N_35965);
or U36641 (N_36641,N_35209,N_35176);
nor U36642 (N_36642,N_35919,N_35304);
nor U36643 (N_36643,N_34059,N_35022);
nand U36644 (N_36644,N_34732,N_35257);
xnor U36645 (N_36645,N_35133,N_34561);
nor U36646 (N_36646,N_34762,N_35424);
xor U36647 (N_36647,N_35767,N_35494);
nand U36648 (N_36648,N_34316,N_34776);
nor U36649 (N_36649,N_35560,N_34956);
xor U36650 (N_36650,N_35379,N_34425);
or U36651 (N_36651,N_34909,N_35536);
or U36652 (N_36652,N_34585,N_35187);
nor U36653 (N_36653,N_34675,N_35049);
or U36654 (N_36654,N_35990,N_34595);
or U36655 (N_36655,N_34818,N_34998);
nor U36656 (N_36656,N_34659,N_35000);
and U36657 (N_36657,N_34323,N_35332);
and U36658 (N_36658,N_35550,N_35927);
nor U36659 (N_36659,N_35999,N_35143);
or U36660 (N_36660,N_34309,N_35575);
or U36661 (N_36661,N_35818,N_34291);
nand U36662 (N_36662,N_35476,N_35989);
and U36663 (N_36663,N_35656,N_34184);
nand U36664 (N_36664,N_34663,N_35057);
and U36665 (N_36665,N_35110,N_35665);
nand U36666 (N_36666,N_35961,N_34848);
or U36667 (N_36667,N_34236,N_34640);
nand U36668 (N_36668,N_35275,N_34310);
xnor U36669 (N_36669,N_35946,N_35881);
and U36670 (N_36670,N_35256,N_35914);
xor U36671 (N_36671,N_34946,N_34174);
and U36672 (N_36672,N_35301,N_34405);
nand U36673 (N_36673,N_34706,N_34730);
or U36674 (N_36674,N_34849,N_34468);
nand U36675 (N_36675,N_34843,N_34033);
nand U36676 (N_36676,N_35282,N_35939);
xnor U36677 (N_36677,N_35794,N_34283);
and U36678 (N_36678,N_34723,N_34894);
xor U36679 (N_36679,N_34149,N_34439);
nor U36680 (N_36680,N_35123,N_35203);
xnor U36681 (N_36681,N_35807,N_34934);
nand U36682 (N_36682,N_35515,N_35162);
nor U36683 (N_36683,N_35437,N_35650);
or U36684 (N_36684,N_35899,N_34491);
nand U36685 (N_36685,N_34217,N_35189);
xor U36686 (N_36686,N_34273,N_34320);
nor U36687 (N_36687,N_35076,N_35996);
xnor U36688 (N_36688,N_34925,N_35159);
and U36689 (N_36689,N_34482,N_35145);
nor U36690 (N_36690,N_34609,N_35717);
and U36691 (N_36691,N_34348,N_34872);
nor U36692 (N_36692,N_35457,N_35935);
and U36693 (N_36693,N_35157,N_34540);
nand U36694 (N_36694,N_34478,N_34919);
xor U36695 (N_36695,N_35156,N_35631);
and U36696 (N_36696,N_35759,N_35475);
or U36697 (N_36697,N_34181,N_34920);
or U36698 (N_36698,N_34867,N_34596);
xor U36699 (N_36699,N_35858,N_35926);
xor U36700 (N_36700,N_34885,N_34274);
or U36701 (N_36701,N_34747,N_35785);
xnor U36702 (N_36702,N_34862,N_35446);
nand U36703 (N_36703,N_34591,N_34359);
or U36704 (N_36704,N_34996,N_35124);
xnor U36705 (N_36705,N_34782,N_35131);
or U36706 (N_36706,N_34459,N_35685);
or U36707 (N_36707,N_34230,N_34583);
xnor U36708 (N_36708,N_35097,N_34968);
nand U36709 (N_36709,N_34549,N_34385);
nand U36710 (N_36710,N_34844,N_34296);
nand U36711 (N_36711,N_34580,N_34386);
nor U36712 (N_36712,N_34189,N_34431);
nor U36713 (N_36713,N_34438,N_34505);
nand U36714 (N_36714,N_35615,N_34989);
nand U36715 (N_36715,N_34353,N_34146);
nand U36716 (N_36716,N_34446,N_34373);
nor U36717 (N_36717,N_35603,N_34955);
and U36718 (N_36718,N_34957,N_35744);
and U36719 (N_36719,N_35565,N_34962);
nand U36720 (N_36720,N_35792,N_34768);
xor U36721 (N_36721,N_35490,N_34288);
and U36722 (N_36722,N_35627,N_35658);
xor U36723 (N_36723,N_34275,N_35811);
nor U36724 (N_36724,N_34007,N_35542);
and U36725 (N_36725,N_34938,N_34022);
and U36726 (N_36726,N_34101,N_35376);
nand U36727 (N_36727,N_34003,N_35317);
and U36728 (N_36728,N_35623,N_34194);
xnor U36729 (N_36729,N_35436,N_35963);
and U36730 (N_36730,N_35984,N_34774);
and U36731 (N_36731,N_35728,N_35223);
or U36732 (N_36732,N_35932,N_35086);
nand U36733 (N_36733,N_34026,N_35690);
xor U36734 (N_36734,N_34874,N_35562);
nor U36735 (N_36735,N_35443,N_34806);
xnor U36736 (N_36736,N_34119,N_35518);
xnor U36737 (N_36737,N_34350,N_34207);
xor U36738 (N_36738,N_34097,N_34153);
or U36739 (N_36739,N_35435,N_34346);
nor U36740 (N_36740,N_35245,N_35842);
or U36741 (N_36741,N_34407,N_34298);
nor U36742 (N_36742,N_34789,N_34087);
xnor U36743 (N_36743,N_35994,N_35311);
or U36744 (N_36744,N_34040,N_35576);
nand U36745 (N_36745,N_35100,N_35966);
nor U36746 (N_36746,N_34088,N_34536);
nor U36747 (N_36747,N_34272,N_35517);
nand U36748 (N_36748,N_35774,N_34180);
nor U36749 (N_36749,N_34967,N_34671);
nand U36750 (N_36750,N_35831,N_34208);
nand U36751 (N_36751,N_35765,N_34817);
and U36752 (N_36752,N_34612,N_34636);
xor U36753 (N_36753,N_35572,N_35937);
nand U36754 (N_36754,N_35249,N_34982);
xnor U36755 (N_36755,N_35653,N_35682);
xnor U36756 (N_36756,N_35951,N_35796);
and U36757 (N_36757,N_35358,N_35265);
nand U36758 (N_36758,N_35051,N_34126);
xnor U36759 (N_36759,N_34284,N_35309);
nand U36760 (N_36760,N_35734,N_35399);
nor U36761 (N_36761,N_34279,N_34892);
and U36762 (N_36762,N_35930,N_35060);
xor U36763 (N_36763,N_34228,N_34836);
or U36764 (N_36764,N_35902,N_34302);
or U36765 (N_36765,N_35978,N_34447);
xor U36766 (N_36766,N_34053,N_35718);
xor U36767 (N_36767,N_34907,N_35499);
xnor U36768 (N_36768,N_34427,N_34897);
nand U36769 (N_36769,N_35194,N_35359);
or U36770 (N_36770,N_34985,N_34085);
nor U36771 (N_36771,N_34435,N_34218);
xnor U36772 (N_36772,N_35461,N_35846);
and U36773 (N_36773,N_35383,N_35689);
or U36774 (N_36774,N_34165,N_34694);
and U36775 (N_36775,N_34801,N_34253);
nor U36776 (N_36776,N_35921,N_34387);
or U36777 (N_36777,N_35024,N_34389);
or U36778 (N_36778,N_35638,N_35597);
and U36779 (N_36779,N_34618,N_34840);
and U36780 (N_36780,N_34741,N_34268);
xor U36781 (N_36781,N_34837,N_34061);
or U36782 (N_36782,N_35177,N_35829);
or U36783 (N_36783,N_35954,N_35105);
nor U36784 (N_36784,N_34788,N_35430);
nor U36785 (N_36785,N_34025,N_35693);
and U36786 (N_36786,N_34409,N_34589);
nand U36787 (N_36787,N_34248,N_35426);
nand U36788 (N_36788,N_35005,N_34440);
nand U36789 (N_36789,N_35471,N_35120);
or U36790 (N_36790,N_35752,N_35720);
and U36791 (N_36791,N_34249,N_34545);
xnor U36792 (N_36792,N_35768,N_34018);
nor U36793 (N_36793,N_35642,N_34838);
xor U36794 (N_36794,N_35092,N_34918);
and U36795 (N_36795,N_35018,N_34226);
and U36796 (N_36796,N_34868,N_34926);
nor U36797 (N_36797,N_35259,N_35844);
or U36798 (N_36798,N_34150,N_34917);
and U36799 (N_36799,N_34451,N_35904);
or U36800 (N_36800,N_35029,N_35377);
or U36801 (N_36801,N_35556,N_35661);
or U36802 (N_36802,N_35913,N_35713);
and U36803 (N_36803,N_34114,N_35986);
or U36804 (N_36804,N_34356,N_35584);
xnor U36805 (N_36805,N_35669,N_35814);
and U36806 (N_36806,N_34558,N_35487);
nor U36807 (N_36807,N_35353,N_35636);
xnor U36808 (N_36808,N_35716,N_35466);
nor U36809 (N_36809,N_34963,N_34187);
or U36810 (N_36810,N_35819,N_35901);
or U36811 (N_36811,N_34045,N_35468);
and U36812 (N_36812,N_34394,N_34269);
nor U36813 (N_36813,N_35126,N_34462);
and U36814 (N_36814,N_35213,N_34547);
and U36815 (N_36815,N_35498,N_34227);
xor U36816 (N_36816,N_35810,N_34223);
and U36817 (N_36817,N_35568,N_35896);
xnor U36818 (N_36818,N_35041,N_35593);
nand U36819 (N_36819,N_34531,N_34044);
or U36820 (N_36820,N_34624,N_35972);
and U36821 (N_36821,N_35224,N_34778);
xnor U36822 (N_36822,N_34319,N_35692);
nor U36823 (N_36823,N_34916,N_34142);
or U36824 (N_36824,N_34467,N_35856);
nand U36825 (N_36825,N_35925,N_34745);
xor U36826 (N_36826,N_34511,N_35454);
xor U36827 (N_36827,N_34028,N_35154);
and U36828 (N_36828,N_34078,N_35292);
nor U36829 (N_36829,N_35806,N_35121);
xnor U36830 (N_36830,N_34658,N_35741);
nand U36831 (N_36831,N_34457,N_34340);
nor U36832 (N_36832,N_34038,N_35087);
and U36833 (N_36833,N_35600,N_34499);
nand U36834 (N_36834,N_34484,N_34108);
nand U36835 (N_36835,N_35587,N_34135);
or U36836 (N_36836,N_35082,N_35843);
and U36837 (N_36837,N_35969,N_34902);
xor U36838 (N_36838,N_35178,N_34721);
or U36839 (N_36839,N_34417,N_35221);
nand U36840 (N_36840,N_34013,N_34066);
or U36841 (N_36841,N_35473,N_35892);
or U36842 (N_36842,N_35467,N_34969);
nor U36843 (N_36843,N_35763,N_34233);
and U36844 (N_36844,N_35616,N_35509);
nor U36845 (N_36845,N_35211,N_35307);
nor U36846 (N_36846,N_35492,N_34041);
and U36847 (N_36847,N_34544,N_34125);
or U36848 (N_36848,N_35534,N_35543);
nand U36849 (N_36849,N_34429,N_35958);
xor U36850 (N_36850,N_35450,N_34758);
xor U36851 (N_36851,N_34615,N_35933);
or U36852 (N_36852,N_35739,N_34687);
xnor U36853 (N_36853,N_35611,N_35637);
and U36854 (N_36854,N_35234,N_34157);
and U36855 (N_36855,N_34339,N_34820);
and U36856 (N_36856,N_34010,N_34211);
nor U36857 (N_36857,N_35191,N_35398);
xor U36858 (N_36858,N_34031,N_34239);
nor U36859 (N_36859,N_34395,N_34746);
xor U36860 (N_36860,N_34380,N_35483);
nand U36861 (N_36861,N_35766,N_35393);
or U36862 (N_36862,N_35895,N_35423);
nor U36863 (N_36863,N_35541,N_35044);
nor U36864 (N_36864,N_34576,N_34067);
xnor U36865 (N_36865,N_34952,N_34263);
or U36866 (N_36866,N_34479,N_35137);
nor U36867 (N_36867,N_35016,N_34116);
nor U36868 (N_36868,N_34406,N_34525);
and U36869 (N_36869,N_34523,N_34630);
xnor U36870 (N_36870,N_35286,N_34792);
or U36871 (N_36871,N_34254,N_34802);
xor U36872 (N_36872,N_35753,N_35341);
or U36873 (N_36873,N_34518,N_35742);
or U36874 (N_36874,N_34987,N_34628);
nand U36875 (N_36875,N_35380,N_34004);
xnor U36876 (N_36876,N_34878,N_34929);
nand U36877 (N_36877,N_34794,N_34378);
xnor U36878 (N_36878,N_35090,N_35853);
or U36879 (N_36879,N_35312,N_34865);
xnor U36880 (N_36880,N_34229,N_34565);
nor U36881 (N_36881,N_35737,N_34880);
xnor U36882 (N_36882,N_34481,N_35345);
or U36883 (N_36883,N_35789,N_35782);
xor U36884 (N_36884,N_35334,N_35169);
xor U36885 (N_36885,N_35748,N_35540);
or U36886 (N_36886,N_35555,N_34127);
or U36887 (N_36887,N_34048,N_35851);
nand U36888 (N_36888,N_34841,N_35055);
nand U36889 (N_36889,N_35415,N_35089);
xnor U36890 (N_36890,N_35825,N_34977);
and U36891 (N_36891,N_34109,N_34363);
or U36892 (N_36892,N_35992,N_35122);
nand U36893 (N_36893,N_35463,N_35268);
nor U36894 (N_36894,N_35772,N_35236);
nand U36895 (N_36895,N_35832,N_34686);
nor U36896 (N_36896,N_34673,N_34238);
nor U36897 (N_36897,N_35172,N_34470);
or U36898 (N_36898,N_35040,N_34113);
or U36899 (N_36899,N_35333,N_35726);
nand U36900 (N_36900,N_35957,N_34783);
xor U36901 (N_36901,N_34351,N_34487);
nor U36902 (N_36902,N_34354,N_35620);
xor U36903 (N_36903,N_34500,N_35671);
xor U36904 (N_36904,N_35805,N_35448);
nand U36905 (N_36905,N_34287,N_34280);
xor U36906 (N_36906,N_34318,N_34688);
nand U36907 (N_36907,N_35849,N_35605);
and U36908 (N_36908,N_35732,N_34267);
nand U36909 (N_36909,N_35096,N_34517);
and U36910 (N_36910,N_35577,N_35147);
xor U36911 (N_36911,N_34711,N_35502);
xnor U36912 (N_36912,N_34796,N_34443);
xnor U36913 (N_36913,N_34294,N_34835);
nand U36914 (N_36914,N_35392,N_35048);
and U36915 (N_36915,N_34808,N_34893);
nor U36916 (N_36916,N_34215,N_34682);
and U36917 (N_36917,N_34131,N_34362);
and U36918 (N_36918,N_35338,N_35977);
xor U36919 (N_36919,N_34191,N_34210);
or U36920 (N_36920,N_34497,N_35405);
or U36921 (N_36921,N_35414,N_34665);
and U36922 (N_36922,N_35777,N_35404);
and U36923 (N_36923,N_34092,N_34420);
nand U36924 (N_36924,N_34634,N_34159);
nand U36925 (N_36925,N_35934,N_34614);
nor U36926 (N_36926,N_35872,N_34120);
nor U36927 (N_36927,N_35015,N_34290);
nand U36928 (N_36928,N_35181,N_35367);
or U36929 (N_36929,N_34024,N_34244);
or U36930 (N_36930,N_34008,N_34433);
and U36931 (N_36931,N_34884,N_34552);
nor U36932 (N_36932,N_35218,N_35545);
and U36933 (N_36933,N_34046,N_34726);
nor U36934 (N_36934,N_34574,N_34588);
and U36935 (N_36935,N_35146,N_34091);
nor U36936 (N_36936,N_34879,N_35950);
nand U36937 (N_36937,N_35144,N_34970);
nor U36938 (N_36938,N_34077,N_34465);
or U36939 (N_36939,N_34691,N_34690);
nor U36940 (N_36940,N_35859,N_35330);
or U36941 (N_36941,N_35019,N_34105);
xnor U36942 (N_36942,N_34261,N_34250);
or U36943 (N_36943,N_34432,N_35582);
xnor U36944 (N_36944,N_35374,N_35783);
xnor U36945 (N_36945,N_34225,N_35821);
and U36946 (N_36946,N_35264,N_35733);
and U36947 (N_36947,N_34785,N_34910);
nand U36948 (N_36948,N_35010,N_35118);
and U36949 (N_36949,N_35835,N_35547);
and U36950 (N_36950,N_35875,N_34075);
or U36951 (N_36951,N_34903,N_34981);
xnor U36952 (N_36952,N_34379,N_34436);
nor U36953 (N_36953,N_35855,N_34904);
nor U36954 (N_36954,N_34991,N_34988);
xor U36955 (N_36955,N_34739,N_35361);
or U36956 (N_36956,N_34870,N_34611);
xor U36957 (N_36957,N_35943,N_35632);
and U36958 (N_36958,N_34924,N_35278);
nand U36959 (N_36959,N_35639,N_34625);
xor U36960 (N_36960,N_35186,N_35208);
nor U36961 (N_36961,N_35505,N_35059);
nand U36962 (N_36962,N_34679,N_35356);
or U36963 (N_36963,N_35365,N_34111);
nand U36964 (N_36964,N_34400,N_34680);
or U36965 (N_36965,N_35879,N_35506);
nor U36966 (N_36966,N_35083,N_34750);
nor U36967 (N_36967,N_34384,N_34369);
or U36968 (N_36968,N_34532,N_35644);
and U36969 (N_36969,N_34605,N_35027);
nand U36970 (N_36970,N_35267,N_35043);
nand U36971 (N_36971,N_35589,N_34550);
nor U36972 (N_36972,N_35607,N_35749);
xnor U36973 (N_36973,N_35959,N_34858);
and U36974 (N_36974,N_35111,N_35604);
and U36975 (N_36975,N_35762,N_35406);
nor U36976 (N_36976,N_35031,N_34483);
and U36977 (N_36977,N_34168,N_35340);
nor U36978 (N_36978,N_34616,N_34607);
or U36979 (N_36979,N_34876,N_34190);
nand U36980 (N_36980,N_34526,N_35971);
nor U36981 (N_36981,N_35290,N_35780);
nand U36982 (N_36982,N_35342,N_35535);
nand U36983 (N_36983,N_34816,N_35706);
xnor U36984 (N_36984,N_34971,N_34029);
or U36985 (N_36985,N_34771,N_34334);
or U36986 (N_36986,N_35687,N_34486);
or U36987 (N_36987,N_34051,N_34156);
nand U36988 (N_36988,N_35870,N_35764);
xnor U36989 (N_36989,N_35564,N_35199);
nand U36990 (N_36990,N_35274,N_34813);
and U36991 (N_36991,N_34266,N_34586);
nand U36992 (N_36992,N_35276,N_35373);
and U36993 (N_36993,N_35170,N_34170);
and U36994 (N_36994,N_35618,N_34709);
and U36995 (N_36995,N_35038,N_35668);
and U36996 (N_36996,N_34344,N_35481);
or U36997 (N_36997,N_35141,N_35231);
or U36998 (N_36998,N_35283,N_34299);
xnor U36999 (N_36999,N_35813,N_35452);
and U37000 (N_37000,N_35061,N_34294);
nand U37001 (N_37001,N_35700,N_34033);
or U37002 (N_37002,N_34095,N_34407);
or U37003 (N_37003,N_34026,N_35616);
or U37004 (N_37004,N_34088,N_34645);
nor U37005 (N_37005,N_35255,N_34582);
nand U37006 (N_37006,N_34492,N_35848);
nand U37007 (N_37007,N_34623,N_34913);
nor U37008 (N_37008,N_34335,N_34040);
and U37009 (N_37009,N_35429,N_35739);
xor U37010 (N_37010,N_35964,N_35813);
xor U37011 (N_37011,N_34769,N_35639);
nor U37012 (N_37012,N_34069,N_34870);
nand U37013 (N_37013,N_34710,N_34916);
nand U37014 (N_37014,N_34139,N_34556);
xnor U37015 (N_37015,N_35149,N_35906);
and U37016 (N_37016,N_35511,N_35970);
nand U37017 (N_37017,N_35417,N_34764);
or U37018 (N_37018,N_35501,N_34556);
or U37019 (N_37019,N_34531,N_35501);
xnor U37020 (N_37020,N_34128,N_35108);
nor U37021 (N_37021,N_35423,N_35091);
xnor U37022 (N_37022,N_35003,N_34502);
nand U37023 (N_37023,N_34604,N_35583);
nor U37024 (N_37024,N_34390,N_35637);
xnor U37025 (N_37025,N_34596,N_35105);
or U37026 (N_37026,N_35132,N_34028);
or U37027 (N_37027,N_35205,N_35478);
nor U37028 (N_37028,N_34490,N_35583);
nand U37029 (N_37029,N_34476,N_35491);
nor U37030 (N_37030,N_34399,N_34478);
nand U37031 (N_37031,N_34889,N_34012);
xor U37032 (N_37032,N_34062,N_35865);
or U37033 (N_37033,N_35167,N_35429);
nor U37034 (N_37034,N_34886,N_34404);
and U37035 (N_37035,N_35592,N_35138);
nand U37036 (N_37036,N_35824,N_34126);
nor U37037 (N_37037,N_34893,N_35522);
nor U37038 (N_37038,N_35575,N_34148);
xor U37039 (N_37039,N_35901,N_34174);
nor U37040 (N_37040,N_35090,N_34869);
or U37041 (N_37041,N_35331,N_35418);
or U37042 (N_37042,N_34905,N_35041);
nor U37043 (N_37043,N_34211,N_35259);
nor U37044 (N_37044,N_35931,N_34233);
nand U37045 (N_37045,N_35169,N_34772);
nand U37046 (N_37046,N_34143,N_35946);
and U37047 (N_37047,N_34483,N_35337);
or U37048 (N_37048,N_35752,N_34615);
and U37049 (N_37049,N_34551,N_35989);
nor U37050 (N_37050,N_34721,N_35740);
nor U37051 (N_37051,N_34318,N_35250);
nor U37052 (N_37052,N_35323,N_34702);
nand U37053 (N_37053,N_35962,N_34010);
nand U37054 (N_37054,N_34259,N_35536);
or U37055 (N_37055,N_35953,N_35568);
or U37056 (N_37056,N_35459,N_35851);
and U37057 (N_37057,N_35934,N_34465);
xor U37058 (N_37058,N_34537,N_35222);
xnor U37059 (N_37059,N_34483,N_35705);
or U37060 (N_37060,N_34960,N_35778);
and U37061 (N_37061,N_34300,N_35583);
nand U37062 (N_37062,N_34084,N_35083);
nor U37063 (N_37063,N_35399,N_35154);
or U37064 (N_37064,N_35869,N_34128);
or U37065 (N_37065,N_34872,N_34632);
or U37066 (N_37066,N_35065,N_35616);
nand U37067 (N_37067,N_34913,N_34482);
nor U37068 (N_37068,N_34546,N_34420);
xor U37069 (N_37069,N_34330,N_34402);
xor U37070 (N_37070,N_34514,N_34893);
xnor U37071 (N_37071,N_35824,N_34365);
xnor U37072 (N_37072,N_35518,N_34635);
or U37073 (N_37073,N_35091,N_35684);
nand U37074 (N_37074,N_34665,N_34079);
or U37075 (N_37075,N_34475,N_35119);
or U37076 (N_37076,N_34752,N_35673);
or U37077 (N_37077,N_34464,N_35036);
or U37078 (N_37078,N_34341,N_34233);
nor U37079 (N_37079,N_34705,N_35845);
nor U37080 (N_37080,N_34097,N_34403);
nand U37081 (N_37081,N_34734,N_34324);
and U37082 (N_37082,N_35373,N_34462);
nand U37083 (N_37083,N_34862,N_35273);
nand U37084 (N_37084,N_34561,N_35759);
or U37085 (N_37085,N_34266,N_35928);
nor U37086 (N_37086,N_34252,N_35243);
nand U37087 (N_37087,N_34073,N_34627);
or U37088 (N_37088,N_34169,N_35352);
nand U37089 (N_37089,N_35450,N_35465);
xor U37090 (N_37090,N_34483,N_34660);
and U37091 (N_37091,N_34385,N_35276);
nor U37092 (N_37092,N_34444,N_34614);
or U37093 (N_37093,N_34732,N_34110);
nand U37094 (N_37094,N_35300,N_34274);
nand U37095 (N_37095,N_34371,N_34806);
nand U37096 (N_37096,N_34905,N_35954);
or U37097 (N_37097,N_35376,N_35422);
nand U37098 (N_37098,N_34446,N_34651);
xor U37099 (N_37099,N_34007,N_35631);
or U37100 (N_37100,N_34800,N_34954);
nand U37101 (N_37101,N_34587,N_34108);
and U37102 (N_37102,N_35070,N_35026);
nor U37103 (N_37103,N_34305,N_34210);
nand U37104 (N_37104,N_34751,N_35849);
or U37105 (N_37105,N_34037,N_35188);
nor U37106 (N_37106,N_35399,N_35817);
nor U37107 (N_37107,N_35115,N_34268);
nor U37108 (N_37108,N_35784,N_34322);
nand U37109 (N_37109,N_35702,N_35551);
and U37110 (N_37110,N_34701,N_34485);
xnor U37111 (N_37111,N_34733,N_34265);
xnor U37112 (N_37112,N_35084,N_34168);
xnor U37113 (N_37113,N_35282,N_34828);
nor U37114 (N_37114,N_34337,N_34229);
xor U37115 (N_37115,N_35652,N_34823);
or U37116 (N_37116,N_35431,N_35602);
or U37117 (N_37117,N_35346,N_34401);
xnor U37118 (N_37118,N_35126,N_34804);
nand U37119 (N_37119,N_34105,N_34392);
nor U37120 (N_37120,N_34804,N_34579);
xor U37121 (N_37121,N_34461,N_34510);
or U37122 (N_37122,N_35578,N_35433);
nor U37123 (N_37123,N_34574,N_34085);
xor U37124 (N_37124,N_35002,N_35769);
nand U37125 (N_37125,N_35744,N_35708);
or U37126 (N_37126,N_34234,N_35171);
or U37127 (N_37127,N_35861,N_34903);
nor U37128 (N_37128,N_35719,N_34572);
and U37129 (N_37129,N_35380,N_35198);
and U37130 (N_37130,N_34471,N_35218);
nand U37131 (N_37131,N_35451,N_34603);
nand U37132 (N_37132,N_35876,N_34924);
or U37133 (N_37133,N_35444,N_35182);
or U37134 (N_37134,N_35119,N_35631);
or U37135 (N_37135,N_35368,N_35175);
and U37136 (N_37136,N_35230,N_35318);
xnor U37137 (N_37137,N_34945,N_34865);
or U37138 (N_37138,N_34605,N_34797);
nor U37139 (N_37139,N_35002,N_35189);
nand U37140 (N_37140,N_35831,N_35361);
xor U37141 (N_37141,N_34217,N_34978);
nor U37142 (N_37142,N_35650,N_34340);
or U37143 (N_37143,N_35881,N_35816);
and U37144 (N_37144,N_35904,N_34407);
and U37145 (N_37145,N_35618,N_35935);
nand U37146 (N_37146,N_35049,N_34599);
or U37147 (N_37147,N_35271,N_34210);
and U37148 (N_37148,N_35635,N_34707);
and U37149 (N_37149,N_34869,N_34387);
nand U37150 (N_37150,N_34909,N_35792);
nor U37151 (N_37151,N_34225,N_35885);
nand U37152 (N_37152,N_34351,N_35988);
nand U37153 (N_37153,N_34808,N_35616);
nand U37154 (N_37154,N_35546,N_35060);
nand U37155 (N_37155,N_35106,N_35248);
nor U37156 (N_37156,N_35416,N_35845);
xor U37157 (N_37157,N_34927,N_34296);
or U37158 (N_37158,N_34000,N_35193);
and U37159 (N_37159,N_35780,N_34393);
nand U37160 (N_37160,N_34471,N_35238);
or U37161 (N_37161,N_35061,N_35243);
and U37162 (N_37162,N_34512,N_34173);
nand U37163 (N_37163,N_34940,N_34060);
nor U37164 (N_37164,N_34664,N_35521);
or U37165 (N_37165,N_35049,N_35828);
or U37166 (N_37166,N_34010,N_34901);
nand U37167 (N_37167,N_35312,N_35392);
nand U37168 (N_37168,N_35692,N_34812);
xor U37169 (N_37169,N_34989,N_34841);
and U37170 (N_37170,N_34978,N_35779);
nor U37171 (N_37171,N_34251,N_34766);
and U37172 (N_37172,N_34224,N_34025);
nand U37173 (N_37173,N_34496,N_35044);
xnor U37174 (N_37174,N_35700,N_35555);
or U37175 (N_37175,N_34823,N_35216);
xor U37176 (N_37176,N_35863,N_34453);
or U37177 (N_37177,N_34789,N_35446);
xnor U37178 (N_37178,N_34560,N_34696);
xor U37179 (N_37179,N_34715,N_34129);
or U37180 (N_37180,N_35282,N_34088);
nor U37181 (N_37181,N_34234,N_35391);
nor U37182 (N_37182,N_35451,N_34377);
and U37183 (N_37183,N_35181,N_35273);
nand U37184 (N_37184,N_35963,N_35541);
nor U37185 (N_37185,N_34601,N_34246);
nand U37186 (N_37186,N_35805,N_34528);
nand U37187 (N_37187,N_35992,N_34824);
or U37188 (N_37188,N_34780,N_34408);
xnor U37189 (N_37189,N_34014,N_35822);
and U37190 (N_37190,N_35232,N_34425);
nor U37191 (N_37191,N_35056,N_35439);
and U37192 (N_37192,N_35050,N_35909);
or U37193 (N_37193,N_35766,N_35290);
or U37194 (N_37194,N_34689,N_34182);
xnor U37195 (N_37195,N_35212,N_35662);
and U37196 (N_37196,N_35271,N_35690);
nor U37197 (N_37197,N_35539,N_35978);
nor U37198 (N_37198,N_34522,N_34262);
nand U37199 (N_37199,N_35502,N_35270);
xor U37200 (N_37200,N_35924,N_35759);
nand U37201 (N_37201,N_35817,N_35016);
xor U37202 (N_37202,N_34189,N_35593);
and U37203 (N_37203,N_35854,N_35599);
nand U37204 (N_37204,N_34487,N_35766);
nand U37205 (N_37205,N_34172,N_34279);
nand U37206 (N_37206,N_35647,N_35338);
or U37207 (N_37207,N_34956,N_34024);
xnor U37208 (N_37208,N_35184,N_35904);
nor U37209 (N_37209,N_35091,N_35976);
and U37210 (N_37210,N_35716,N_34788);
and U37211 (N_37211,N_34796,N_35532);
or U37212 (N_37212,N_34706,N_35492);
and U37213 (N_37213,N_35978,N_34835);
nor U37214 (N_37214,N_34726,N_35656);
xnor U37215 (N_37215,N_35891,N_35225);
or U37216 (N_37216,N_34034,N_34625);
and U37217 (N_37217,N_34397,N_34589);
nor U37218 (N_37218,N_34485,N_34285);
or U37219 (N_37219,N_34529,N_34023);
and U37220 (N_37220,N_34722,N_35134);
and U37221 (N_37221,N_34241,N_34818);
xnor U37222 (N_37222,N_34966,N_34144);
nor U37223 (N_37223,N_34569,N_34104);
or U37224 (N_37224,N_35514,N_34775);
xnor U37225 (N_37225,N_35462,N_34939);
and U37226 (N_37226,N_34165,N_34342);
xor U37227 (N_37227,N_34880,N_35857);
nand U37228 (N_37228,N_34632,N_34942);
nand U37229 (N_37229,N_35438,N_35530);
nor U37230 (N_37230,N_34045,N_34740);
nor U37231 (N_37231,N_34949,N_34292);
or U37232 (N_37232,N_35505,N_34823);
nor U37233 (N_37233,N_34073,N_35007);
and U37234 (N_37234,N_34167,N_35107);
nor U37235 (N_37235,N_35271,N_34556);
xor U37236 (N_37236,N_34635,N_34483);
and U37237 (N_37237,N_35338,N_35869);
nand U37238 (N_37238,N_34115,N_34749);
or U37239 (N_37239,N_35913,N_34351);
or U37240 (N_37240,N_35581,N_35961);
and U37241 (N_37241,N_34990,N_35482);
xnor U37242 (N_37242,N_35253,N_34762);
nor U37243 (N_37243,N_34180,N_35609);
nand U37244 (N_37244,N_34428,N_34241);
and U37245 (N_37245,N_34747,N_35197);
xnor U37246 (N_37246,N_35358,N_34219);
nand U37247 (N_37247,N_34435,N_35070);
nand U37248 (N_37248,N_34635,N_35069);
nand U37249 (N_37249,N_35732,N_35832);
nor U37250 (N_37250,N_34754,N_34366);
or U37251 (N_37251,N_34354,N_35019);
nor U37252 (N_37252,N_35081,N_35662);
and U37253 (N_37253,N_35158,N_34410);
nand U37254 (N_37254,N_35042,N_34872);
and U37255 (N_37255,N_34528,N_34026);
and U37256 (N_37256,N_35650,N_35874);
nand U37257 (N_37257,N_35500,N_35810);
and U37258 (N_37258,N_34488,N_35694);
nand U37259 (N_37259,N_34769,N_34279);
nor U37260 (N_37260,N_34924,N_35588);
nor U37261 (N_37261,N_34997,N_34511);
nor U37262 (N_37262,N_35359,N_34786);
nand U37263 (N_37263,N_34633,N_35210);
or U37264 (N_37264,N_35221,N_35576);
nand U37265 (N_37265,N_35613,N_34247);
xor U37266 (N_37266,N_34937,N_35346);
xnor U37267 (N_37267,N_34460,N_34218);
nor U37268 (N_37268,N_35647,N_35929);
xnor U37269 (N_37269,N_34119,N_35326);
or U37270 (N_37270,N_34167,N_34225);
nor U37271 (N_37271,N_35810,N_35673);
and U37272 (N_37272,N_35890,N_35011);
nor U37273 (N_37273,N_34431,N_34526);
nor U37274 (N_37274,N_35913,N_35848);
xor U37275 (N_37275,N_35755,N_34043);
xnor U37276 (N_37276,N_35134,N_34598);
xor U37277 (N_37277,N_35343,N_35507);
or U37278 (N_37278,N_35011,N_35781);
and U37279 (N_37279,N_35213,N_34422);
or U37280 (N_37280,N_35654,N_34279);
nand U37281 (N_37281,N_35835,N_34976);
nor U37282 (N_37282,N_34112,N_34601);
and U37283 (N_37283,N_34070,N_35825);
nor U37284 (N_37284,N_35902,N_34633);
nor U37285 (N_37285,N_34967,N_34617);
nor U37286 (N_37286,N_35924,N_34181);
or U37287 (N_37287,N_35133,N_34687);
or U37288 (N_37288,N_35636,N_35343);
or U37289 (N_37289,N_34553,N_35604);
xnor U37290 (N_37290,N_34281,N_35729);
or U37291 (N_37291,N_34460,N_34097);
and U37292 (N_37292,N_34733,N_34767);
xor U37293 (N_37293,N_35204,N_34359);
xnor U37294 (N_37294,N_34950,N_35486);
nor U37295 (N_37295,N_35132,N_35120);
nand U37296 (N_37296,N_34580,N_35381);
or U37297 (N_37297,N_35855,N_35440);
xnor U37298 (N_37298,N_34761,N_35654);
nand U37299 (N_37299,N_34291,N_35413);
nand U37300 (N_37300,N_34833,N_34734);
nor U37301 (N_37301,N_35291,N_35974);
nor U37302 (N_37302,N_34455,N_34758);
or U37303 (N_37303,N_35247,N_35183);
xor U37304 (N_37304,N_34020,N_35952);
and U37305 (N_37305,N_35075,N_34818);
nand U37306 (N_37306,N_34983,N_35367);
nor U37307 (N_37307,N_35156,N_35838);
nor U37308 (N_37308,N_35051,N_35901);
nor U37309 (N_37309,N_35233,N_35903);
and U37310 (N_37310,N_34117,N_34640);
nor U37311 (N_37311,N_34991,N_35929);
xor U37312 (N_37312,N_35222,N_35369);
or U37313 (N_37313,N_35393,N_35947);
or U37314 (N_37314,N_35620,N_34492);
nand U37315 (N_37315,N_35914,N_34814);
nor U37316 (N_37316,N_35661,N_34398);
nor U37317 (N_37317,N_35846,N_35023);
or U37318 (N_37318,N_35798,N_35530);
and U37319 (N_37319,N_34070,N_35672);
xor U37320 (N_37320,N_34572,N_35273);
nand U37321 (N_37321,N_35197,N_35432);
or U37322 (N_37322,N_34520,N_35400);
xnor U37323 (N_37323,N_35384,N_34382);
and U37324 (N_37324,N_34904,N_35978);
nor U37325 (N_37325,N_35982,N_35384);
nand U37326 (N_37326,N_35109,N_34466);
and U37327 (N_37327,N_35848,N_34941);
and U37328 (N_37328,N_34093,N_34460);
nor U37329 (N_37329,N_34990,N_35084);
nor U37330 (N_37330,N_34838,N_34005);
xor U37331 (N_37331,N_34773,N_34390);
and U37332 (N_37332,N_34397,N_35542);
and U37333 (N_37333,N_34248,N_34094);
and U37334 (N_37334,N_35000,N_34386);
and U37335 (N_37335,N_35347,N_34677);
xnor U37336 (N_37336,N_34778,N_34977);
nand U37337 (N_37337,N_34117,N_34752);
nor U37338 (N_37338,N_35526,N_35321);
xnor U37339 (N_37339,N_35562,N_35173);
or U37340 (N_37340,N_34023,N_34553);
nand U37341 (N_37341,N_35663,N_35157);
and U37342 (N_37342,N_35859,N_35684);
and U37343 (N_37343,N_35052,N_34680);
nor U37344 (N_37344,N_35870,N_35252);
nand U37345 (N_37345,N_34063,N_35603);
nand U37346 (N_37346,N_35536,N_34405);
or U37347 (N_37347,N_35765,N_35726);
xnor U37348 (N_37348,N_34329,N_35410);
xor U37349 (N_37349,N_34173,N_34810);
and U37350 (N_37350,N_34460,N_35491);
nand U37351 (N_37351,N_34587,N_34227);
xor U37352 (N_37352,N_34999,N_35014);
nor U37353 (N_37353,N_35874,N_34083);
or U37354 (N_37354,N_34015,N_34830);
or U37355 (N_37355,N_35755,N_35325);
nand U37356 (N_37356,N_34970,N_34757);
nand U37357 (N_37357,N_35073,N_34086);
or U37358 (N_37358,N_34982,N_34305);
nand U37359 (N_37359,N_35685,N_35625);
or U37360 (N_37360,N_34383,N_34970);
nand U37361 (N_37361,N_34877,N_35724);
or U37362 (N_37362,N_34437,N_35866);
nand U37363 (N_37363,N_35944,N_35046);
and U37364 (N_37364,N_35432,N_35361);
or U37365 (N_37365,N_34129,N_35003);
or U37366 (N_37366,N_34977,N_34235);
nand U37367 (N_37367,N_34370,N_35309);
nand U37368 (N_37368,N_34017,N_34151);
nand U37369 (N_37369,N_34985,N_35220);
xor U37370 (N_37370,N_35704,N_34070);
and U37371 (N_37371,N_34493,N_34105);
and U37372 (N_37372,N_34741,N_35803);
or U37373 (N_37373,N_34219,N_35606);
nor U37374 (N_37374,N_34807,N_34552);
nor U37375 (N_37375,N_35823,N_35508);
nor U37376 (N_37376,N_34215,N_35224);
nand U37377 (N_37377,N_34214,N_35053);
or U37378 (N_37378,N_34096,N_35557);
or U37379 (N_37379,N_34757,N_35063);
and U37380 (N_37380,N_34219,N_35272);
nand U37381 (N_37381,N_35716,N_35123);
nand U37382 (N_37382,N_34490,N_35007);
nor U37383 (N_37383,N_34912,N_35462);
nand U37384 (N_37384,N_34004,N_35274);
xor U37385 (N_37385,N_35867,N_34972);
nor U37386 (N_37386,N_35539,N_35551);
nor U37387 (N_37387,N_34588,N_34916);
xnor U37388 (N_37388,N_35126,N_34215);
or U37389 (N_37389,N_34551,N_34573);
xor U37390 (N_37390,N_35368,N_35221);
xnor U37391 (N_37391,N_35557,N_34459);
nand U37392 (N_37392,N_34789,N_34243);
or U37393 (N_37393,N_34829,N_34725);
xor U37394 (N_37394,N_35654,N_34029);
or U37395 (N_37395,N_34006,N_35658);
nand U37396 (N_37396,N_34320,N_35978);
nand U37397 (N_37397,N_34983,N_35455);
nor U37398 (N_37398,N_35825,N_34922);
or U37399 (N_37399,N_34875,N_35002);
and U37400 (N_37400,N_35730,N_34039);
and U37401 (N_37401,N_34245,N_34350);
or U37402 (N_37402,N_35597,N_35922);
nor U37403 (N_37403,N_34628,N_35828);
nor U37404 (N_37404,N_35253,N_34050);
and U37405 (N_37405,N_34643,N_35386);
nor U37406 (N_37406,N_34003,N_35439);
nand U37407 (N_37407,N_34166,N_34118);
nor U37408 (N_37408,N_34484,N_35089);
and U37409 (N_37409,N_35206,N_35718);
xor U37410 (N_37410,N_34417,N_34122);
xor U37411 (N_37411,N_35924,N_34726);
xor U37412 (N_37412,N_35752,N_34258);
nand U37413 (N_37413,N_35141,N_35685);
xnor U37414 (N_37414,N_35882,N_35744);
nand U37415 (N_37415,N_34499,N_35435);
and U37416 (N_37416,N_35978,N_34486);
nor U37417 (N_37417,N_34978,N_34901);
nand U37418 (N_37418,N_35001,N_35370);
nand U37419 (N_37419,N_35561,N_35304);
and U37420 (N_37420,N_34866,N_34300);
xor U37421 (N_37421,N_34056,N_34536);
and U37422 (N_37422,N_34934,N_35011);
nor U37423 (N_37423,N_34842,N_35125);
nand U37424 (N_37424,N_35462,N_34316);
xnor U37425 (N_37425,N_35673,N_35199);
and U37426 (N_37426,N_34590,N_34575);
xnor U37427 (N_37427,N_34590,N_35098);
nand U37428 (N_37428,N_35643,N_35885);
nand U37429 (N_37429,N_35025,N_34565);
or U37430 (N_37430,N_34057,N_35639);
nand U37431 (N_37431,N_34795,N_35357);
and U37432 (N_37432,N_35920,N_35256);
nor U37433 (N_37433,N_35444,N_35165);
and U37434 (N_37434,N_35337,N_34936);
nand U37435 (N_37435,N_34155,N_35743);
nor U37436 (N_37436,N_35904,N_34425);
nor U37437 (N_37437,N_34343,N_34033);
nand U37438 (N_37438,N_35183,N_35863);
nand U37439 (N_37439,N_35239,N_34513);
nor U37440 (N_37440,N_34108,N_35903);
nor U37441 (N_37441,N_34534,N_35563);
and U37442 (N_37442,N_34781,N_34190);
and U37443 (N_37443,N_35815,N_34632);
xor U37444 (N_37444,N_35325,N_34535);
nand U37445 (N_37445,N_35880,N_34938);
nand U37446 (N_37446,N_35336,N_34214);
nand U37447 (N_37447,N_35777,N_35090);
xnor U37448 (N_37448,N_34979,N_34872);
or U37449 (N_37449,N_35995,N_35585);
and U37450 (N_37450,N_35843,N_34756);
nor U37451 (N_37451,N_35751,N_35928);
nor U37452 (N_37452,N_34258,N_35145);
xnor U37453 (N_37453,N_35570,N_35993);
and U37454 (N_37454,N_35053,N_34711);
nor U37455 (N_37455,N_35085,N_34684);
nand U37456 (N_37456,N_35451,N_34970);
xor U37457 (N_37457,N_35503,N_34322);
and U37458 (N_37458,N_35199,N_35983);
and U37459 (N_37459,N_35889,N_35010);
xor U37460 (N_37460,N_34681,N_35703);
or U37461 (N_37461,N_34147,N_34550);
xor U37462 (N_37462,N_35796,N_35116);
or U37463 (N_37463,N_35807,N_34645);
xor U37464 (N_37464,N_35332,N_34170);
nand U37465 (N_37465,N_34835,N_35355);
nand U37466 (N_37466,N_34239,N_35375);
and U37467 (N_37467,N_35261,N_34215);
xnor U37468 (N_37468,N_34369,N_34897);
nor U37469 (N_37469,N_35093,N_35511);
and U37470 (N_37470,N_35753,N_35070);
or U37471 (N_37471,N_34056,N_34216);
nor U37472 (N_37472,N_35686,N_35538);
nand U37473 (N_37473,N_35444,N_34071);
nor U37474 (N_37474,N_34795,N_35188);
and U37475 (N_37475,N_35605,N_35326);
nand U37476 (N_37476,N_35067,N_34366);
and U37477 (N_37477,N_35845,N_34396);
nand U37478 (N_37478,N_34471,N_35527);
or U37479 (N_37479,N_35515,N_35713);
nor U37480 (N_37480,N_34120,N_34725);
or U37481 (N_37481,N_35288,N_34959);
or U37482 (N_37482,N_34678,N_35675);
or U37483 (N_37483,N_34779,N_35182);
nor U37484 (N_37484,N_35990,N_34713);
and U37485 (N_37485,N_35606,N_34640);
nand U37486 (N_37486,N_35171,N_34301);
nand U37487 (N_37487,N_35764,N_34636);
or U37488 (N_37488,N_34084,N_35143);
xnor U37489 (N_37489,N_34307,N_35947);
nand U37490 (N_37490,N_35656,N_35196);
and U37491 (N_37491,N_35572,N_35086);
nor U37492 (N_37492,N_35984,N_35471);
and U37493 (N_37493,N_34961,N_35031);
and U37494 (N_37494,N_34486,N_34887);
nand U37495 (N_37495,N_34581,N_34716);
or U37496 (N_37496,N_34524,N_35895);
nand U37497 (N_37497,N_34848,N_34826);
or U37498 (N_37498,N_35680,N_34340);
or U37499 (N_37499,N_34175,N_35217);
nor U37500 (N_37500,N_34732,N_35167);
nand U37501 (N_37501,N_35065,N_35186);
and U37502 (N_37502,N_34802,N_35535);
or U37503 (N_37503,N_34508,N_35238);
xor U37504 (N_37504,N_34182,N_34943);
xor U37505 (N_37505,N_34242,N_34687);
xnor U37506 (N_37506,N_34061,N_35689);
or U37507 (N_37507,N_35390,N_35615);
nand U37508 (N_37508,N_35422,N_34253);
or U37509 (N_37509,N_35615,N_34688);
nand U37510 (N_37510,N_35996,N_34695);
and U37511 (N_37511,N_35350,N_34073);
xnor U37512 (N_37512,N_35594,N_35782);
and U37513 (N_37513,N_35460,N_34908);
and U37514 (N_37514,N_35408,N_35153);
or U37515 (N_37515,N_35610,N_34821);
or U37516 (N_37516,N_35083,N_34670);
and U37517 (N_37517,N_35057,N_34841);
and U37518 (N_37518,N_34812,N_35317);
or U37519 (N_37519,N_34195,N_34098);
and U37520 (N_37520,N_35027,N_34432);
and U37521 (N_37521,N_35442,N_34372);
xor U37522 (N_37522,N_35098,N_35442);
nor U37523 (N_37523,N_35107,N_34547);
nand U37524 (N_37524,N_35163,N_34886);
nand U37525 (N_37525,N_34878,N_35523);
xor U37526 (N_37526,N_34136,N_34363);
and U37527 (N_37527,N_35414,N_34731);
or U37528 (N_37528,N_35368,N_34166);
nor U37529 (N_37529,N_35695,N_34365);
and U37530 (N_37530,N_34610,N_34301);
nand U37531 (N_37531,N_35876,N_34210);
and U37532 (N_37532,N_35605,N_35592);
xor U37533 (N_37533,N_35596,N_35175);
and U37534 (N_37534,N_34248,N_35207);
and U37535 (N_37535,N_35033,N_34608);
nor U37536 (N_37536,N_34787,N_34225);
nor U37537 (N_37537,N_34627,N_34938);
or U37538 (N_37538,N_35260,N_34577);
nand U37539 (N_37539,N_35252,N_35393);
nand U37540 (N_37540,N_35285,N_34448);
or U37541 (N_37541,N_34886,N_35077);
nand U37542 (N_37542,N_35541,N_34282);
nand U37543 (N_37543,N_34945,N_34518);
xnor U37544 (N_37544,N_34683,N_34511);
or U37545 (N_37545,N_35283,N_34174);
nor U37546 (N_37546,N_35721,N_34216);
xnor U37547 (N_37547,N_35264,N_35752);
or U37548 (N_37548,N_34331,N_34280);
or U37549 (N_37549,N_34289,N_34137);
nand U37550 (N_37550,N_34751,N_35147);
and U37551 (N_37551,N_34992,N_34599);
nor U37552 (N_37552,N_34063,N_35881);
nand U37553 (N_37553,N_34003,N_34389);
nor U37554 (N_37554,N_34250,N_34303);
and U37555 (N_37555,N_35179,N_34765);
and U37556 (N_37556,N_34001,N_35289);
xor U37557 (N_37557,N_35590,N_34615);
nand U37558 (N_37558,N_34924,N_34571);
nor U37559 (N_37559,N_34185,N_35707);
nand U37560 (N_37560,N_34420,N_35589);
xor U37561 (N_37561,N_34450,N_34853);
or U37562 (N_37562,N_34912,N_35630);
nand U37563 (N_37563,N_34636,N_34880);
nor U37564 (N_37564,N_34764,N_35259);
or U37565 (N_37565,N_35548,N_35011);
xnor U37566 (N_37566,N_35496,N_35442);
or U37567 (N_37567,N_34305,N_35804);
nand U37568 (N_37568,N_35921,N_35252);
or U37569 (N_37569,N_35121,N_34202);
nor U37570 (N_37570,N_34961,N_35335);
or U37571 (N_37571,N_35178,N_35636);
nor U37572 (N_37572,N_35976,N_34009);
nand U37573 (N_37573,N_34223,N_34635);
nand U37574 (N_37574,N_34108,N_35240);
xor U37575 (N_37575,N_34565,N_34520);
xnor U37576 (N_37576,N_35675,N_34279);
and U37577 (N_37577,N_35015,N_35938);
or U37578 (N_37578,N_34950,N_34762);
nor U37579 (N_37579,N_35363,N_34503);
and U37580 (N_37580,N_34949,N_35600);
and U37581 (N_37581,N_34792,N_35709);
nand U37582 (N_37582,N_34865,N_35529);
and U37583 (N_37583,N_34016,N_35721);
xnor U37584 (N_37584,N_35085,N_34824);
xnor U37585 (N_37585,N_35035,N_34492);
or U37586 (N_37586,N_35137,N_35188);
nor U37587 (N_37587,N_35185,N_34368);
nor U37588 (N_37588,N_35936,N_34329);
nor U37589 (N_37589,N_34828,N_35888);
nand U37590 (N_37590,N_34740,N_34579);
nand U37591 (N_37591,N_35488,N_34054);
and U37592 (N_37592,N_34343,N_34238);
xnor U37593 (N_37593,N_35705,N_35378);
and U37594 (N_37594,N_34477,N_35277);
and U37595 (N_37595,N_35381,N_34399);
xnor U37596 (N_37596,N_35904,N_34338);
and U37597 (N_37597,N_34958,N_34699);
or U37598 (N_37598,N_34747,N_35088);
or U37599 (N_37599,N_35586,N_35940);
nor U37600 (N_37600,N_34294,N_35183);
nand U37601 (N_37601,N_34990,N_35693);
nor U37602 (N_37602,N_34348,N_34005);
or U37603 (N_37603,N_34992,N_35853);
and U37604 (N_37604,N_35471,N_34227);
nor U37605 (N_37605,N_34813,N_35388);
or U37606 (N_37606,N_35908,N_34833);
and U37607 (N_37607,N_35491,N_34404);
nor U37608 (N_37608,N_35211,N_34262);
and U37609 (N_37609,N_35858,N_35534);
nand U37610 (N_37610,N_34981,N_34769);
or U37611 (N_37611,N_34541,N_35804);
nor U37612 (N_37612,N_35545,N_35746);
and U37613 (N_37613,N_35553,N_35989);
and U37614 (N_37614,N_35873,N_34535);
nand U37615 (N_37615,N_34492,N_34126);
nand U37616 (N_37616,N_34131,N_35862);
or U37617 (N_37617,N_34994,N_34261);
xnor U37618 (N_37618,N_34640,N_34554);
or U37619 (N_37619,N_34776,N_34609);
nand U37620 (N_37620,N_34006,N_34844);
nand U37621 (N_37621,N_35730,N_34739);
or U37622 (N_37622,N_35360,N_35409);
or U37623 (N_37623,N_35279,N_35019);
nor U37624 (N_37624,N_35096,N_35069);
xnor U37625 (N_37625,N_35637,N_34313);
nor U37626 (N_37626,N_34535,N_34575);
nor U37627 (N_37627,N_35277,N_35828);
xor U37628 (N_37628,N_34285,N_35064);
or U37629 (N_37629,N_35812,N_35130);
nand U37630 (N_37630,N_34654,N_34597);
and U37631 (N_37631,N_34377,N_35204);
or U37632 (N_37632,N_34851,N_34459);
or U37633 (N_37633,N_35733,N_34742);
or U37634 (N_37634,N_35531,N_34349);
or U37635 (N_37635,N_35553,N_35319);
and U37636 (N_37636,N_34624,N_35057);
nor U37637 (N_37637,N_34357,N_34530);
xnor U37638 (N_37638,N_35948,N_34224);
and U37639 (N_37639,N_34871,N_34424);
or U37640 (N_37640,N_34487,N_35247);
nor U37641 (N_37641,N_34388,N_34157);
xnor U37642 (N_37642,N_35150,N_35524);
xnor U37643 (N_37643,N_35998,N_35075);
xor U37644 (N_37644,N_35957,N_35537);
nor U37645 (N_37645,N_34712,N_34236);
or U37646 (N_37646,N_34385,N_34079);
or U37647 (N_37647,N_34031,N_35290);
nand U37648 (N_37648,N_34048,N_35840);
nand U37649 (N_37649,N_35073,N_34833);
xnor U37650 (N_37650,N_34387,N_35828);
or U37651 (N_37651,N_34519,N_35536);
nand U37652 (N_37652,N_35736,N_34041);
or U37653 (N_37653,N_35911,N_34698);
and U37654 (N_37654,N_34033,N_34307);
nor U37655 (N_37655,N_35057,N_35794);
nor U37656 (N_37656,N_35141,N_35198);
or U37657 (N_37657,N_35593,N_34987);
nor U37658 (N_37658,N_35497,N_34573);
nand U37659 (N_37659,N_34578,N_35864);
xnor U37660 (N_37660,N_35351,N_34980);
and U37661 (N_37661,N_34674,N_35642);
or U37662 (N_37662,N_35612,N_34117);
nor U37663 (N_37663,N_34863,N_35899);
nand U37664 (N_37664,N_35944,N_34809);
nand U37665 (N_37665,N_34685,N_34533);
or U37666 (N_37666,N_35591,N_35751);
nand U37667 (N_37667,N_34433,N_34481);
and U37668 (N_37668,N_35143,N_35966);
or U37669 (N_37669,N_35047,N_34259);
nor U37670 (N_37670,N_34883,N_34281);
nand U37671 (N_37671,N_34302,N_35504);
nand U37672 (N_37672,N_34644,N_34684);
nor U37673 (N_37673,N_35312,N_34005);
nand U37674 (N_37674,N_35678,N_34897);
xnor U37675 (N_37675,N_35752,N_34029);
nor U37676 (N_37676,N_35074,N_35675);
nand U37677 (N_37677,N_35867,N_34235);
xnor U37678 (N_37678,N_35818,N_34424);
nor U37679 (N_37679,N_35524,N_35695);
nand U37680 (N_37680,N_35567,N_34138);
nand U37681 (N_37681,N_35218,N_35750);
and U37682 (N_37682,N_34986,N_35761);
xor U37683 (N_37683,N_35352,N_34605);
nand U37684 (N_37684,N_35636,N_34874);
nand U37685 (N_37685,N_35261,N_34665);
nand U37686 (N_37686,N_35457,N_35654);
nor U37687 (N_37687,N_35178,N_35388);
nand U37688 (N_37688,N_35714,N_35039);
and U37689 (N_37689,N_34178,N_34415);
nor U37690 (N_37690,N_35411,N_34505);
nor U37691 (N_37691,N_35577,N_35336);
xor U37692 (N_37692,N_34328,N_35259);
or U37693 (N_37693,N_35712,N_35044);
xor U37694 (N_37694,N_34910,N_35220);
nand U37695 (N_37695,N_35532,N_34317);
and U37696 (N_37696,N_35665,N_35069);
or U37697 (N_37697,N_35595,N_34408);
xnor U37698 (N_37698,N_35657,N_35207);
and U37699 (N_37699,N_35017,N_35752);
nor U37700 (N_37700,N_34195,N_34087);
or U37701 (N_37701,N_34614,N_35834);
nor U37702 (N_37702,N_34002,N_35224);
nand U37703 (N_37703,N_35151,N_35645);
nor U37704 (N_37704,N_35509,N_34769);
xor U37705 (N_37705,N_34446,N_34630);
or U37706 (N_37706,N_34597,N_34695);
and U37707 (N_37707,N_35170,N_34497);
nand U37708 (N_37708,N_35420,N_35520);
nand U37709 (N_37709,N_34052,N_35505);
and U37710 (N_37710,N_35983,N_35961);
and U37711 (N_37711,N_34900,N_35927);
or U37712 (N_37712,N_35948,N_34191);
and U37713 (N_37713,N_34670,N_34403);
xnor U37714 (N_37714,N_35019,N_35793);
xnor U37715 (N_37715,N_35480,N_35468);
xor U37716 (N_37716,N_34387,N_34160);
and U37717 (N_37717,N_34663,N_35611);
and U37718 (N_37718,N_35511,N_35827);
nor U37719 (N_37719,N_34506,N_35172);
and U37720 (N_37720,N_35475,N_34089);
and U37721 (N_37721,N_35497,N_34073);
nand U37722 (N_37722,N_34696,N_35027);
and U37723 (N_37723,N_35325,N_34237);
and U37724 (N_37724,N_35875,N_34617);
nand U37725 (N_37725,N_35531,N_34504);
or U37726 (N_37726,N_35816,N_35156);
xnor U37727 (N_37727,N_35636,N_35821);
and U37728 (N_37728,N_35590,N_35809);
and U37729 (N_37729,N_34890,N_35600);
or U37730 (N_37730,N_34625,N_35964);
nor U37731 (N_37731,N_34989,N_34222);
or U37732 (N_37732,N_35010,N_34492);
and U37733 (N_37733,N_34323,N_34213);
nand U37734 (N_37734,N_35908,N_34165);
nand U37735 (N_37735,N_34089,N_35315);
nand U37736 (N_37736,N_35219,N_35262);
xnor U37737 (N_37737,N_35837,N_35212);
or U37738 (N_37738,N_35843,N_35108);
and U37739 (N_37739,N_34210,N_34244);
and U37740 (N_37740,N_34769,N_35075);
and U37741 (N_37741,N_34456,N_35202);
and U37742 (N_37742,N_34856,N_35015);
xnor U37743 (N_37743,N_35541,N_35000);
or U37744 (N_37744,N_35357,N_35619);
nand U37745 (N_37745,N_35965,N_34389);
nor U37746 (N_37746,N_35022,N_34377);
nand U37747 (N_37747,N_35120,N_35339);
or U37748 (N_37748,N_34437,N_34762);
and U37749 (N_37749,N_34018,N_34853);
and U37750 (N_37750,N_34679,N_34655);
nor U37751 (N_37751,N_34263,N_35112);
nand U37752 (N_37752,N_34990,N_35255);
or U37753 (N_37753,N_34792,N_34211);
xor U37754 (N_37754,N_35274,N_34084);
or U37755 (N_37755,N_34503,N_34010);
xnor U37756 (N_37756,N_35253,N_35667);
nand U37757 (N_37757,N_34631,N_35239);
nand U37758 (N_37758,N_35396,N_34083);
nor U37759 (N_37759,N_34896,N_35149);
or U37760 (N_37760,N_34836,N_35559);
and U37761 (N_37761,N_34314,N_34586);
nand U37762 (N_37762,N_35705,N_34336);
xor U37763 (N_37763,N_34934,N_35874);
nor U37764 (N_37764,N_35171,N_35649);
xnor U37765 (N_37765,N_35199,N_34399);
xor U37766 (N_37766,N_34038,N_34358);
nand U37767 (N_37767,N_34879,N_34988);
nand U37768 (N_37768,N_35065,N_35012);
nand U37769 (N_37769,N_35433,N_34381);
nor U37770 (N_37770,N_34182,N_35575);
nand U37771 (N_37771,N_34597,N_34911);
or U37772 (N_37772,N_34631,N_34682);
xnor U37773 (N_37773,N_35754,N_35709);
or U37774 (N_37774,N_34956,N_34239);
or U37775 (N_37775,N_34260,N_34575);
and U37776 (N_37776,N_34156,N_34333);
or U37777 (N_37777,N_34388,N_34586);
or U37778 (N_37778,N_35065,N_35561);
and U37779 (N_37779,N_34416,N_34172);
xnor U37780 (N_37780,N_35097,N_34483);
or U37781 (N_37781,N_35514,N_34453);
xnor U37782 (N_37782,N_34759,N_35919);
xor U37783 (N_37783,N_35430,N_34242);
xor U37784 (N_37784,N_35054,N_35970);
nor U37785 (N_37785,N_35374,N_34905);
nand U37786 (N_37786,N_34673,N_34312);
or U37787 (N_37787,N_35654,N_34514);
xnor U37788 (N_37788,N_34216,N_34089);
and U37789 (N_37789,N_35276,N_34910);
nand U37790 (N_37790,N_34830,N_34634);
or U37791 (N_37791,N_34847,N_34826);
nor U37792 (N_37792,N_35731,N_35126);
xor U37793 (N_37793,N_35769,N_35682);
nand U37794 (N_37794,N_34650,N_35728);
xor U37795 (N_37795,N_35254,N_34283);
nor U37796 (N_37796,N_34392,N_35820);
xnor U37797 (N_37797,N_35537,N_35666);
xnor U37798 (N_37798,N_34235,N_34119);
and U37799 (N_37799,N_35044,N_35149);
nand U37800 (N_37800,N_34943,N_35990);
and U37801 (N_37801,N_35273,N_35959);
or U37802 (N_37802,N_35886,N_35552);
nand U37803 (N_37803,N_34052,N_34667);
xor U37804 (N_37804,N_34255,N_34995);
nor U37805 (N_37805,N_34518,N_34533);
and U37806 (N_37806,N_35148,N_34007);
nor U37807 (N_37807,N_34713,N_35081);
or U37808 (N_37808,N_34401,N_34466);
nand U37809 (N_37809,N_34827,N_34768);
or U37810 (N_37810,N_34398,N_35431);
and U37811 (N_37811,N_34791,N_34282);
nand U37812 (N_37812,N_34095,N_34633);
or U37813 (N_37813,N_35024,N_34956);
and U37814 (N_37814,N_34968,N_34751);
xnor U37815 (N_37815,N_35160,N_35435);
nor U37816 (N_37816,N_35898,N_34189);
xnor U37817 (N_37817,N_34097,N_34183);
nor U37818 (N_37818,N_34255,N_35128);
nor U37819 (N_37819,N_34812,N_34963);
nand U37820 (N_37820,N_35405,N_35894);
nand U37821 (N_37821,N_34147,N_35092);
or U37822 (N_37822,N_34821,N_35366);
nand U37823 (N_37823,N_35135,N_34998);
or U37824 (N_37824,N_35019,N_35111);
nand U37825 (N_37825,N_34323,N_34144);
and U37826 (N_37826,N_34445,N_35970);
or U37827 (N_37827,N_35543,N_34037);
or U37828 (N_37828,N_34761,N_35151);
nand U37829 (N_37829,N_35627,N_35770);
or U37830 (N_37830,N_34343,N_35945);
xor U37831 (N_37831,N_35547,N_35010);
xor U37832 (N_37832,N_35173,N_34403);
or U37833 (N_37833,N_34161,N_34931);
nand U37834 (N_37834,N_35499,N_35953);
nor U37835 (N_37835,N_34638,N_34077);
xnor U37836 (N_37836,N_35490,N_34657);
and U37837 (N_37837,N_35080,N_34508);
nor U37838 (N_37838,N_34423,N_34163);
or U37839 (N_37839,N_34133,N_34823);
nor U37840 (N_37840,N_34651,N_34584);
xnor U37841 (N_37841,N_35566,N_34475);
and U37842 (N_37842,N_34187,N_34300);
nand U37843 (N_37843,N_34433,N_34343);
and U37844 (N_37844,N_34447,N_35847);
xnor U37845 (N_37845,N_34872,N_35987);
and U37846 (N_37846,N_34785,N_34816);
or U37847 (N_37847,N_34836,N_35790);
nor U37848 (N_37848,N_35890,N_34662);
nand U37849 (N_37849,N_35657,N_35845);
nand U37850 (N_37850,N_35705,N_35265);
nor U37851 (N_37851,N_34671,N_34688);
and U37852 (N_37852,N_35294,N_35178);
nor U37853 (N_37853,N_34114,N_35338);
nand U37854 (N_37854,N_34591,N_35151);
nand U37855 (N_37855,N_35487,N_34314);
or U37856 (N_37856,N_35394,N_34749);
nor U37857 (N_37857,N_34816,N_34497);
nor U37858 (N_37858,N_35919,N_35569);
and U37859 (N_37859,N_35735,N_35654);
or U37860 (N_37860,N_34927,N_34468);
or U37861 (N_37861,N_34515,N_35313);
nand U37862 (N_37862,N_35636,N_34142);
nand U37863 (N_37863,N_35221,N_34607);
and U37864 (N_37864,N_34846,N_35531);
and U37865 (N_37865,N_35734,N_35327);
and U37866 (N_37866,N_34341,N_34002);
nand U37867 (N_37867,N_34449,N_35440);
and U37868 (N_37868,N_35797,N_35506);
or U37869 (N_37869,N_34111,N_35525);
xnor U37870 (N_37870,N_35873,N_34786);
nand U37871 (N_37871,N_35601,N_35824);
nand U37872 (N_37872,N_34917,N_35216);
and U37873 (N_37873,N_35510,N_35822);
or U37874 (N_37874,N_35410,N_34146);
and U37875 (N_37875,N_34471,N_35868);
or U37876 (N_37876,N_35754,N_35155);
nor U37877 (N_37877,N_34299,N_34841);
and U37878 (N_37878,N_35444,N_34080);
and U37879 (N_37879,N_35275,N_34229);
or U37880 (N_37880,N_34082,N_34652);
nor U37881 (N_37881,N_34325,N_34225);
or U37882 (N_37882,N_35968,N_34875);
or U37883 (N_37883,N_35971,N_34261);
and U37884 (N_37884,N_35821,N_35275);
nor U37885 (N_37885,N_34735,N_35433);
or U37886 (N_37886,N_34027,N_35798);
nand U37887 (N_37887,N_34988,N_35110);
xor U37888 (N_37888,N_34827,N_34388);
and U37889 (N_37889,N_35896,N_34833);
xor U37890 (N_37890,N_34215,N_34103);
xnor U37891 (N_37891,N_35744,N_34541);
and U37892 (N_37892,N_34334,N_35724);
nand U37893 (N_37893,N_34524,N_35471);
xor U37894 (N_37894,N_34994,N_34065);
and U37895 (N_37895,N_35530,N_34149);
or U37896 (N_37896,N_34961,N_35041);
or U37897 (N_37897,N_34781,N_35279);
or U37898 (N_37898,N_34114,N_34820);
or U37899 (N_37899,N_35489,N_35089);
nand U37900 (N_37900,N_34371,N_35347);
nor U37901 (N_37901,N_34538,N_35100);
nand U37902 (N_37902,N_35383,N_34963);
nand U37903 (N_37903,N_34538,N_34810);
xnor U37904 (N_37904,N_34561,N_35221);
or U37905 (N_37905,N_35556,N_35184);
nand U37906 (N_37906,N_35565,N_35292);
xnor U37907 (N_37907,N_34325,N_34524);
xor U37908 (N_37908,N_35917,N_34055);
or U37909 (N_37909,N_34857,N_35752);
nor U37910 (N_37910,N_35852,N_34553);
nor U37911 (N_37911,N_35191,N_34585);
xnor U37912 (N_37912,N_35277,N_34857);
or U37913 (N_37913,N_35430,N_35767);
and U37914 (N_37914,N_35646,N_35508);
xor U37915 (N_37915,N_34964,N_35938);
nand U37916 (N_37916,N_35806,N_34161);
or U37917 (N_37917,N_35578,N_35077);
and U37918 (N_37918,N_35726,N_34875);
and U37919 (N_37919,N_34110,N_34654);
xnor U37920 (N_37920,N_35697,N_34883);
or U37921 (N_37921,N_34527,N_35135);
nand U37922 (N_37922,N_34701,N_35737);
and U37923 (N_37923,N_34276,N_34828);
and U37924 (N_37924,N_35880,N_35961);
nand U37925 (N_37925,N_34747,N_34790);
or U37926 (N_37926,N_35313,N_34647);
nand U37927 (N_37927,N_35261,N_35850);
nand U37928 (N_37928,N_35850,N_34159);
and U37929 (N_37929,N_35316,N_35253);
and U37930 (N_37930,N_34823,N_35300);
xnor U37931 (N_37931,N_35828,N_35487);
nand U37932 (N_37932,N_34353,N_35269);
and U37933 (N_37933,N_34637,N_34136);
nor U37934 (N_37934,N_34799,N_34951);
nor U37935 (N_37935,N_34240,N_35456);
and U37936 (N_37936,N_35005,N_34620);
or U37937 (N_37937,N_35860,N_34696);
xor U37938 (N_37938,N_34608,N_34038);
nand U37939 (N_37939,N_35258,N_35964);
nand U37940 (N_37940,N_35745,N_34458);
nand U37941 (N_37941,N_35281,N_35385);
xnor U37942 (N_37942,N_35259,N_34418);
xnor U37943 (N_37943,N_34227,N_34833);
and U37944 (N_37944,N_35490,N_35247);
nor U37945 (N_37945,N_35819,N_34741);
nand U37946 (N_37946,N_35990,N_35181);
nor U37947 (N_37947,N_35010,N_35441);
or U37948 (N_37948,N_35465,N_34551);
nand U37949 (N_37949,N_34731,N_34539);
nand U37950 (N_37950,N_34258,N_35120);
nand U37951 (N_37951,N_35465,N_34189);
xor U37952 (N_37952,N_35961,N_35186);
nand U37953 (N_37953,N_35008,N_35549);
or U37954 (N_37954,N_34341,N_35290);
nor U37955 (N_37955,N_35027,N_35797);
or U37956 (N_37956,N_34140,N_34606);
nor U37957 (N_37957,N_35455,N_34772);
or U37958 (N_37958,N_35161,N_34491);
or U37959 (N_37959,N_34690,N_35535);
nand U37960 (N_37960,N_34725,N_35913);
and U37961 (N_37961,N_35790,N_34651);
nand U37962 (N_37962,N_35226,N_34533);
xnor U37963 (N_37963,N_34070,N_34583);
xor U37964 (N_37964,N_35223,N_34013);
nand U37965 (N_37965,N_35525,N_35667);
xnor U37966 (N_37966,N_34548,N_34002);
xor U37967 (N_37967,N_34802,N_35553);
and U37968 (N_37968,N_35726,N_34043);
and U37969 (N_37969,N_34589,N_34348);
nor U37970 (N_37970,N_35931,N_34063);
and U37971 (N_37971,N_35863,N_34644);
or U37972 (N_37972,N_34555,N_35072);
xor U37973 (N_37973,N_35548,N_35495);
and U37974 (N_37974,N_34709,N_34902);
and U37975 (N_37975,N_34945,N_34092);
or U37976 (N_37976,N_35918,N_35545);
and U37977 (N_37977,N_34670,N_35397);
xor U37978 (N_37978,N_34929,N_35915);
nand U37979 (N_37979,N_34554,N_34645);
nor U37980 (N_37980,N_34327,N_35363);
nand U37981 (N_37981,N_34495,N_35870);
or U37982 (N_37982,N_34903,N_34104);
xnor U37983 (N_37983,N_34852,N_35679);
and U37984 (N_37984,N_34489,N_35736);
and U37985 (N_37985,N_35684,N_35422);
and U37986 (N_37986,N_34796,N_34078);
or U37987 (N_37987,N_34722,N_34650);
and U37988 (N_37988,N_34901,N_34989);
xnor U37989 (N_37989,N_34430,N_34092);
xnor U37990 (N_37990,N_35126,N_34062);
xor U37991 (N_37991,N_35627,N_35765);
and U37992 (N_37992,N_34944,N_34530);
and U37993 (N_37993,N_35828,N_34323);
or U37994 (N_37994,N_34606,N_34186);
and U37995 (N_37995,N_35146,N_35211);
xnor U37996 (N_37996,N_35212,N_34863);
nand U37997 (N_37997,N_35624,N_34897);
nand U37998 (N_37998,N_34471,N_34708);
or U37999 (N_37999,N_35295,N_35258);
nor U38000 (N_38000,N_37363,N_37760);
and U38001 (N_38001,N_36866,N_36654);
xnor U38002 (N_38002,N_37731,N_36664);
and U38003 (N_38003,N_37181,N_36646);
or U38004 (N_38004,N_36071,N_36182);
xor U38005 (N_38005,N_36648,N_36483);
and U38006 (N_38006,N_37640,N_36593);
xnor U38007 (N_38007,N_37820,N_37212);
nor U38008 (N_38008,N_36164,N_36374);
nand U38009 (N_38009,N_36158,N_36303);
nand U38010 (N_38010,N_36460,N_36361);
and U38011 (N_38011,N_37400,N_36327);
nor U38012 (N_38012,N_36898,N_37342);
and U38013 (N_38013,N_37126,N_37420);
nor U38014 (N_38014,N_36555,N_37156);
nor U38015 (N_38015,N_37158,N_36272);
xor U38016 (N_38016,N_36538,N_37571);
xor U38017 (N_38017,N_36780,N_37852);
nand U38018 (N_38018,N_36639,N_36293);
nand U38019 (N_38019,N_36045,N_36682);
or U38020 (N_38020,N_36310,N_36473);
and U38021 (N_38021,N_36261,N_37573);
or U38022 (N_38022,N_36104,N_37246);
nor U38023 (N_38023,N_37679,N_36137);
and U38024 (N_38024,N_36521,N_37377);
or U38025 (N_38025,N_36816,N_36305);
and U38026 (N_38026,N_37105,N_37065);
xor U38027 (N_38027,N_36236,N_37556);
or U38028 (N_38028,N_37801,N_37225);
or U38029 (N_38029,N_37694,N_37869);
xor U38030 (N_38030,N_37681,N_36421);
and U38031 (N_38031,N_37079,N_36124);
or U38032 (N_38032,N_36707,N_37486);
and U38033 (N_38033,N_37103,N_36867);
or U38034 (N_38034,N_36763,N_36641);
nor U38035 (N_38035,N_36729,N_36192);
nand U38036 (N_38036,N_37123,N_36714);
xor U38037 (N_38037,N_37879,N_36776);
nand U38038 (N_38038,N_37429,N_36455);
xnor U38039 (N_38039,N_36083,N_37371);
nand U38040 (N_38040,N_37697,N_36434);
nand U38041 (N_38041,N_36069,N_36477);
or U38042 (N_38042,N_36534,N_36435);
xnor U38043 (N_38043,N_36933,N_37992);
and U38044 (N_38044,N_37952,N_37417);
nand U38045 (N_38045,N_37182,N_37289);
and U38046 (N_38046,N_36977,N_36438);
nor U38047 (N_38047,N_36739,N_37498);
nor U38048 (N_38048,N_37629,N_37749);
nor U38049 (N_38049,N_36352,N_36793);
nor U38050 (N_38050,N_37579,N_36895);
xnor U38051 (N_38051,N_37740,N_36291);
xor U38052 (N_38052,N_36587,N_36458);
nor U38053 (N_38053,N_37927,N_37537);
xor U38054 (N_38054,N_36363,N_37496);
nand U38055 (N_38055,N_36114,N_36098);
or U38056 (N_38056,N_37900,N_37948);
nor U38057 (N_38057,N_36650,N_37755);
xnor U38058 (N_38058,N_37903,N_37373);
xnor U38059 (N_38059,N_36903,N_37099);
or U38060 (N_38060,N_36513,N_37138);
or U38061 (N_38061,N_36242,N_37794);
and U38062 (N_38062,N_37557,N_37443);
and U38063 (N_38063,N_37837,N_37616);
xor U38064 (N_38064,N_36338,N_36580);
and U38065 (N_38065,N_36319,N_37863);
and U38066 (N_38066,N_37322,N_37478);
or U38067 (N_38067,N_36336,N_36723);
nor U38068 (N_38068,N_36886,N_36115);
xnor U38069 (N_38069,N_36789,N_36270);
nand U38070 (N_38070,N_36373,N_37015);
xnor U38071 (N_38071,N_36197,N_37303);
nand U38072 (N_38072,N_37328,N_36812);
or U38073 (N_38073,N_36086,N_36616);
nand U38074 (N_38074,N_37608,N_37506);
and U38075 (N_38075,N_36391,N_36476);
and U38076 (N_38076,N_37418,N_37121);
nand U38077 (N_38077,N_36404,N_36875);
nor U38078 (N_38078,N_36378,N_36204);
or U38079 (N_38079,N_37944,N_37764);
or U38080 (N_38080,N_37603,N_37811);
nand U38081 (N_38081,N_37255,N_37871);
or U38082 (N_38082,N_36079,N_37597);
and U38083 (N_38083,N_37386,N_36200);
xor U38084 (N_38084,N_36941,N_36288);
or U38085 (N_38085,N_37058,N_36949);
nor U38086 (N_38086,N_37711,N_37221);
xnor U38087 (N_38087,N_36478,N_36016);
or U38088 (N_38088,N_37489,N_36413);
xnor U38089 (N_38089,N_37440,N_37765);
or U38090 (N_38090,N_37931,N_37922);
or U38091 (N_38091,N_36173,N_37534);
and U38092 (N_38092,N_37753,N_36148);
or U38093 (N_38093,N_37827,N_36068);
xnor U38094 (N_38094,N_37735,N_37487);
and U38095 (N_38095,N_37204,N_37797);
nand U38096 (N_38096,N_36834,N_36915);
and U38097 (N_38097,N_36752,N_37073);
or U38098 (N_38098,N_36582,N_36792);
xor U38099 (N_38099,N_37460,N_37240);
or U38100 (N_38100,N_36120,N_37905);
xnor U38101 (N_38101,N_36202,N_36459);
nor U38102 (N_38102,N_36259,N_36800);
nor U38103 (N_38103,N_37214,N_37913);
or U38104 (N_38104,N_37151,N_36688);
nor U38105 (N_38105,N_36661,N_36076);
and U38106 (N_38106,N_36094,N_37335);
xor U38107 (N_38107,N_37874,N_37552);
nor U38108 (N_38108,N_37631,N_37149);
nor U38109 (N_38109,N_36656,N_37332);
or U38110 (N_38110,N_36316,N_37928);
nand U38111 (N_38111,N_36936,N_36398);
nand U38112 (N_38112,N_36228,N_37048);
or U38113 (N_38113,N_37844,N_36890);
or U38114 (N_38114,N_37865,N_37933);
nor U38115 (N_38115,N_37914,N_37062);
xnor U38116 (N_38116,N_37353,N_36576);
and U38117 (N_38117,N_36484,N_36999);
and U38118 (N_38118,N_36751,N_36395);
and U38119 (N_38119,N_37494,N_36420);
nor U38120 (N_38120,N_36611,N_36328);
nor U38121 (N_38121,N_37106,N_36559);
xnor U38122 (N_38122,N_36469,N_36782);
nor U38123 (N_38123,N_37578,N_36479);
xnor U38124 (N_38124,N_37877,N_37399);
or U38125 (N_38125,N_37680,N_37309);
xor U38126 (N_38126,N_36838,N_36837);
or U38127 (N_38127,N_37887,N_36566);
xnor U38128 (N_38128,N_36618,N_36480);
nor U38129 (N_38129,N_36399,N_37056);
nor U38130 (N_38130,N_37733,N_36110);
nand U38131 (N_38131,N_37997,N_36529);
xor U38132 (N_38132,N_37770,N_37947);
xnor U38133 (N_38133,N_36368,N_36367);
xnor U38134 (N_38134,N_37834,N_37031);
xor U38135 (N_38135,N_37935,N_36452);
xor U38136 (N_38136,N_37012,N_36612);
nor U38137 (N_38137,N_36108,N_36194);
xnor U38138 (N_38138,N_37059,N_36051);
nor U38139 (N_38139,N_37977,N_37361);
xnor U38140 (N_38140,N_36324,N_36926);
xnor U38141 (N_38141,N_36117,N_36931);
nor U38142 (N_38142,N_37554,N_36871);
xnor U38143 (N_38143,N_37684,N_37621);
or U38144 (N_38144,N_37404,N_37160);
or U38145 (N_38145,N_36064,N_36302);
or U38146 (N_38146,N_37370,N_37722);
xor U38147 (N_38147,N_36377,N_36839);
xnor U38148 (N_38148,N_36741,N_36512);
nand U38149 (N_38149,N_37643,N_36041);
and U38150 (N_38150,N_37517,N_37462);
or U38151 (N_38151,N_36526,N_36916);
or U38152 (N_38152,N_36528,N_37108);
nor U38153 (N_38153,N_37210,N_36863);
nor U38154 (N_38154,N_36351,N_36761);
nand U38155 (N_38155,N_37639,N_37209);
and U38156 (N_38156,N_37604,N_36217);
and U38157 (N_38157,N_37347,N_37199);
nand U38158 (N_38158,N_37800,N_36570);
xnor U38159 (N_38159,N_37349,N_36610);
nand U38160 (N_38160,N_36085,N_37841);
xnor U38161 (N_38161,N_36353,N_36457);
nor U38162 (N_38162,N_36870,N_36998);
nor U38163 (N_38163,N_37019,N_37451);
nand U38164 (N_38164,N_36248,N_37043);
or U38165 (N_38165,N_36665,N_36709);
or U38166 (N_38166,N_37367,N_36187);
nor U38167 (N_38167,N_37778,N_36176);
xor U38168 (N_38168,N_36706,N_37713);
xnor U38169 (N_38169,N_37743,N_37061);
and U38170 (N_38170,N_37939,N_36737);
and U38171 (N_38171,N_37127,N_37252);
and U38172 (N_38172,N_37424,N_37553);
and U38173 (N_38173,N_36364,N_37767);
or U38174 (N_38174,N_37021,N_37144);
nand U38175 (N_38175,N_36055,N_36732);
xnor U38176 (N_38176,N_37995,N_37710);
nor U38177 (N_38177,N_37628,N_37086);
xor U38178 (N_38178,N_36784,N_36686);
xnor U38179 (N_38179,N_37412,N_37134);
or U38180 (N_38180,N_36074,N_37752);
nor U38181 (N_38181,N_37320,N_36599);
nand U38182 (N_38182,N_36928,N_36963);
xor U38183 (N_38183,N_36728,N_36198);
nand U38184 (N_38184,N_37002,N_36062);
xnor U38185 (N_38185,N_37279,N_37634);
nand U38186 (N_38186,N_37272,N_37479);
and U38187 (N_38187,N_36472,N_36600);
and U38188 (N_38188,N_37908,N_37202);
nand U38189 (N_38189,N_37244,N_36702);
or U38190 (N_38190,N_37430,N_37191);
and U38191 (N_38191,N_37786,N_36733);
or U38192 (N_38192,N_37981,N_37512);
nand U38193 (N_38193,N_36354,N_37372);
xor U38194 (N_38194,N_37832,N_37861);
nand U38195 (N_38195,N_37164,N_36394);
xnor U38196 (N_38196,N_37276,N_36273);
nand U38197 (N_38197,N_36713,N_37183);
xnor U38198 (N_38198,N_36872,N_37883);
and U38199 (N_38199,N_37060,N_37102);
and U38200 (N_38200,N_36753,N_37354);
nor U38201 (N_38201,N_37780,N_36226);
nor U38202 (N_38202,N_36285,N_36381);
xor U38203 (N_38203,N_36919,N_37890);
or U38204 (N_38204,N_36581,N_36901);
or U38205 (N_38205,N_36255,N_37333);
nand U38206 (N_38206,N_37613,N_36823);
and U38207 (N_38207,N_36216,N_36342);
and U38208 (N_38208,N_37439,N_37216);
or U38209 (N_38209,N_37539,N_37878);
xor U38210 (N_38210,N_36082,N_37720);
nand U38211 (N_38211,N_37366,N_36296);
and U38212 (N_38212,N_36093,N_36408);
xnor U38213 (N_38213,N_37951,N_36005);
xnor U38214 (N_38214,N_36383,N_37943);
and U38215 (N_38215,N_37311,N_36320);
nor U38216 (N_38216,N_36986,N_36636);
and U38217 (N_38217,N_37416,N_36038);
or U38218 (N_38218,N_37566,N_37954);
and U38219 (N_38219,N_37185,N_37583);
and U38220 (N_38220,N_37170,N_37175);
nand U38221 (N_38221,N_37670,N_37859);
nand U38222 (N_38222,N_37484,N_36149);
nor U38223 (N_38223,N_36097,N_36390);
xor U38224 (N_38224,N_37810,N_36230);
and U38225 (N_38225,N_37978,N_37344);
or U38226 (N_38226,N_36846,N_37482);
nor U38227 (N_38227,N_36254,N_36668);
nand U38228 (N_38228,N_37096,N_37337);
nand U38229 (N_38229,N_36043,N_36499);
or U38230 (N_38230,N_37504,N_37660);
and U38231 (N_38231,N_36208,N_37411);
and U38232 (N_38232,N_36498,N_36238);
or U38233 (N_38233,N_36152,N_36918);
and U38234 (N_38234,N_37845,N_36119);
nand U38235 (N_38235,N_36175,N_37916);
nand U38236 (N_38236,N_37074,N_37812);
nand U38237 (N_38237,N_36830,N_37077);
nor U38238 (N_38238,N_36827,N_36500);
nand U38239 (N_38239,N_37113,N_37438);
nand U38240 (N_38240,N_36249,N_37034);
and U38241 (N_38241,N_36315,N_36658);
nor U38242 (N_38242,N_36970,N_37708);
nand U38243 (N_38243,N_37024,N_37783);
nand U38244 (N_38244,N_36579,N_36878);
or U38245 (N_38245,N_36321,N_37107);
or U38246 (N_38246,N_37858,N_37682);
or U38247 (N_38247,N_36196,N_37232);
nor U38248 (N_38248,N_37548,N_37192);
nor U38249 (N_38249,N_37799,N_37120);
nand U38250 (N_38250,N_37261,N_36609);
xnor U38251 (N_38251,N_37251,N_37282);
or U38252 (N_38252,N_37265,N_37757);
and U38253 (N_38253,N_37409,N_36024);
nor U38254 (N_38254,N_37287,N_37104);
nand U38255 (N_38255,N_37166,N_36670);
or U38256 (N_38256,N_37626,N_36298);
xor U38257 (N_38257,N_37092,N_36134);
nand U38258 (N_38258,N_37567,N_37003);
xnor U38259 (N_38259,N_36740,N_36466);
nand U38260 (N_38260,N_37315,N_37041);
or U38261 (N_38261,N_36525,N_37461);
or U38262 (N_38262,N_36461,N_36357);
or U38263 (N_38263,N_36721,N_37758);
and U38264 (N_38264,N_36130,N_36608);
or U38265 (N_38265,N_36814,N_37744);
or U38266 (N_38266,N_37612,N_36962);
or U38267 (N_38267,N_36366,N_36844);
nor U38268 (N_38268,N_37685,N_37676);
nor U38269 (N_38269,N_36450,N_37860);
xor U38270 (N_38270,N_37445,N_37706);
xnor U38271 (N_38271,N_37044,N_37088);
xor U38272 (N_38272,N_37008,N_37394);
nand U38273 (N_38273,N_36719,N_36932);
and U38274 (N_38274,N_36783,N_36794);
xnor U38275 (N_38275,N_36004,N_36125);
or U38276 (N_38276,N_36507,N_36541);
and U38277 (N_38277,N_37924,N_36758);
xor U38278 (N_38278,N_36874,N_37705);
and U38279 (N_38279,N_37205,N_37538);
nand U38280 (N_38280,N_37020,N_36384);
nor U38281 (N_38281,N_37369,N_36821);
xor U38282 (N_38282,N_37678,N_36433);
nand U38283 (N_38283,N_37875,N_37638);
nor U38284 (N_38284,N_36923,N_36245);
and U38285 (N_38285,N_37917,N_36058);
nand U38286 (N_38286,N_37250,N_36442);
xnor U38287 (N_38287,N_37838,N_36141);
nand U38288 (N_38288,N_37340,N_37173);
nand U38289 (N_38289,N_36899,N_37259);
xnor U38290 (N_38290,N_37958,N_37206);
nand U38291 (N_38291,N_36300,N_36205);
xor U38292 (N_38292,N_37081,N_37395);
or U38293 (N_38293,N_37690,N_37379);
or U38294 (N_38294,N_37502,N_36191);
nand U38295 (N_38295,N_37306,N_37715);
xnor U38296 (N_38296,N_37381,N_36703);
xnor U38297 (N_38297,N_36002,N_37280);
or U38298 (N_38298,N_36030,N_36222);
nand U38299 (N_38299,N_36388,N_36974);
nor U38300 (N_38300,N_36166,N_37700);
xor U38301 (N_38301,N_36632,N_36103);
xnor U38302 (N_38302,N_36920,N_36676);
and U38303 (N_38303,N_37421,N_37897);
nor U38304 (N_38304,N_37000,N_37745);
nand U38305 (N_38305,N_36403,N_36123);
xor U38306 (N_38306,N_37599,N_36008);
nand U38307 (N_38307,N_37356,N_37094);
xor U38308 (N_38308,N_37137,N_37862);
nand U38309 (N_38309,N_37892,N_36880);
nand U38310 (N_38310,N_36537,N_36567);
nand U38311 (N_38311,N_37131,N_36971);
or U38312 (N_38312,N_37348,N_37910);
or U38313 (N_38313,N_36511,N_37918);
nand U38314 (N_38314,N_36893,N_37480);
or U38315 (N_38315,N_36588,N_36666);
nor U38316 (N_38316,N_36778,N_36649);
nor U38317 (N_38317,N_37576,N_36536);
and U38318 (N_38318,N_36809,N_36449);
xor U38319 (N_38319,N_36127,N_37437);
and U38320 (N_38320,N_37324,N_37703);
nor U38321 (N_38321,N_37623,N_36023);
nand U38322 (N_38322,N_37806,N_36340);
and U38323 (N_38323,N_36046,N_37655);
and U38324 (N_38324,N_37382,N_36817);
or U38325 (N_38325,N_37876,N_37991);
xor U38326 (N_38326,N_36683,N_36162);
nand U38327 (N_38327,N_36243,N_37581);
nand U38328 (N_38328,N_37920,N_37521);
nor U38329 (N_38329,N_37477,N_36050);
nor U38330 (N_38330,N_37433,N_37835);
and U38331 (N_38331,N_36430,N_37465);
and U38332 (N_38332,N_36463,N_37231);
nand U38333 (N_38333,N_36225,N_36482);
xnor U38334 (N_38334,N_37912,N_36504);
and U38335 (N_38335,N_37789,N_36414);
or U38336 (N_38336,N_36955,N_37965);
or U38337 (N_38337,N_36358,N_36400);
nor U38338 (N_38338,N_37586,N_36060);
and U38339 (N_38339,N_37618,N_37736);
and U38340 (N_38340,N_37526,N_37001);
xnor U38341 (N_38341,N_36172,N_36239);
nor U38342 (N_38342,N_37622,N_37119);
nand U38343 (N_38343,N_36940,N_37392);
xor U38344 (N_38344,N_37211,N_37600);
xor U38345 (N_38345,N_36927,N_37518);
nand U38346 (N_38346,N_36642,N_36750);
and U38347 (N_38347,N_37213,N_37636);
nand U38348 (N_38348,N_37821,N_36096);
xnor U38349 (N_38349,N_37899,N_37803);
or U38350 (N_38350,N_37915,N_37693);
or U38351 (N_38351,N_37063,N_37304);
or U38352 (N_38352,N_37727,N_37963);
and U38353 (N_38353,N_36308,N_36199);
xnor U38354 (N_38354,N_37569,N_37028);
xnor U38355 (N_38355,N_36615,N_36237);
nor U38356 (N_38356,N_37025,N_36271);
or U38357 (N_38357,N_36048,N_36179);
and U38358 (N_38358,N_36685,N_37281);
and U38359 (N_38359,N_36040,N_37692);
xnor U38360 (N_38360,N_36138,N_37666);
and U38361 (N_38361,N_36859,N_36978);
and U38362 (N_38362,N_37241,N_36849);
or U38363 (N_38363,N_36334,N_36563);
and U38364 (N_38364,N_37606,N_37906);
nand U38365 (N_38365,N_37926,N_37426);
or U38366 (N_38366,N_37042,N_36485);
nand U38367 (N_38367,N_36475,N_36335);
and U38368 (N_38368,N_36836,N_36712);
or U38369 (N_38369,N_37667,N_36551);
xnor U38370 (N_38370,N_36195,N_36907);
or U38371 (N_38371,N_37207,N_37949);
or U38372 (N_38372,N_37046,N_36744);
xnor U38373 (N_38373,N_37341,N_36142);
nand U38374 (N_38374,N_37334,N_37974);
and U38375 (N_38375,N_37983,N_36808);
or U38376 (N_38376,N_36885,N_36339);
or U38377 (N_38377,N_36864,N_36211);
and U38378 (N_38378,N_37243,N_36795);
xnor U38379 (N_38379,N_37560,N_36779);
or U38380 (N_38380,N_37169,N_37432);
or U38381 (N_38381,N_37707,N_36307);
or U38382 (N_38382,N_37718,N_36720);
or U38383 (N_38383,N_36690,N_36036);
nor U38384 (N_38384,N_36956,N_36917);
and U38385 (N_38385,N_37793,N_37148);
and U38386 (N_38386,N_36231,N_36798);
nand U38387 (N_38387,N_36277,N_37784);
nand U38388 (N_38388,N_37157,N_37781);
or U38389 (N_38389,N_36715,N_36930);
or U38390 (N_38390,N_36799,N_37428);
nand U38391 (N_38391,N_37085,N_37047);
and U38392 (N_38392,N_36948,N_36323);
nor U38393 (N_38393,N_37474,N_37452);
and U38394 (N_38394,N_36219,N_36356);
nand U38395 (N_38395,N_36185,N_37714);
nand U38396 (N_38396,N_37542,N_36680);
or U38397 (N_38397,N_37234,N_37220);
or U38398 (N_38398,N_36633,N_37768);
and U38399 (N_38399,N_37946,N_36811);
or U38400 (N_38400,N_36681,N_36897);
xnor U38401 (N_38401,N_36329,N_37719);
xor U38402 (N_38402,N_36787,N_37387);
nor U38403 (N_38403,N_37540,N_36547);
xnor U38404 (N_38404,N_37150,N_37141);
and U38405 (N_38405,N_36644,N_36545);
xor U38406 (N_38406,N_36026,N_37193);
nand U38407 (N_38407,N_37605,N_36423);
nor U38408 (N_38408,N_37070,N_37551);
or U38409 (N_38409,N_36032,N_37435);
nor U38410 (N_38410,N_37891,N_36825);
and U38411 (N_38411,N_37338,N_37263);
nor U38412 (N_38412,N_36453,N_36126);
nor U38413 (N_38413,N_36451,N_36969);
xor U38414 (N_38414,N_36934,N_36966);
nand U38415 (N_38415,N_37975,N_37635);
or U38416 (N_38416,N_36170,N_37804);
nand U38417 (N_38417,N_37167,N_37302);
xnor U38418 (N_38418,N_37033,N_37291);
xnor U38419 (N_38419,N_37093,N_36077);
xnor U38420 (N_38420,N_37468,N_36313);
xnor U38421 (N_38421,N_37580,N_37475);
xor U38422 (N_38422,N_36167,N_36154);
and U38423 (N_38423,N_36637,N_37350);
nor U38424 (N_38424,N_36835,N_37796);
nor U38425 (N_38425,N_36330,N_36535);
or U38426 (N_38426,N_36968,N_37275);
and U38427 (N_38427,N_37130,N_37739);
nor U38428 (N_38428,N_36139,N_37203);
nand U38429 (N_38429,N_36441,N_36078);
and U38430 (N_38430,N_36292,N_37762);
xor U38431 (N_38431,N_37738,N_37601);
or U38432 (N_38432,N_36635,N_37530);
xnor U38433 (N_38433,N_36772,N_37159);
or U38434 (N_38434,N_36868,N_37546);
or U38435 (N_38435,N_37614,N_36253);
and U38436 (N_38436,N_37419,N_37620);
nor U38437 (N_38437,N_36505,N_37989);
or U38438 (N_38438,N_37775,N_36274);
nand U38439 (N_38439,N_37030,N_37967);
nand U38440 (N_38440,N_37630,N_37896);
and U38441 (N_38441,N_36251,N_37114);
nor U38442 (N_38442,N_37162,N_36462);
or U38443 (N_38443,N_37375,N_36630);
nand U38444 (N_38444,N_37091,N_37339);
or U38445 (N_38445,N_37893,N_36989);
nand U38446 (N_38446,N_36552,N_37669);
xor U38447 (N_38447,N_36696,N_36544);
xor U38448 (N_38448,N_36426,N_36369);
or U38449 (N_38449,N_36284,N_36748);
and U38450 (N_38450,N_36663,N_37346);
or U38451 (N_38451,N_37592,N_37568);
xnor U38452 (N_38452,N_36877,N_37870);
nand U38453 (N_38453,N_36424,N_37559);
and U38454 (N_38454,N_36781,N_36973);
nor U38455 (N_38455,N_36089,N_37994);
or U38456 (N_38456,N_36726,N_37146);
nor U38457 (N_38457,N_36386,N_37087);
nand U38458 (N_38458,N_36826,N_37505);
nor U38459 (N_38459,N_36954,N_37766);
nand U38460 (N_38460,N_36586,N_36568);
or U38461 (N_38461,N_37442,N_37378);
and U38462 (N_38462,N_36095,N_37808);
and U38463 (N_38463,N_36266,N_36994);
xor U38464 (N_38464,N_36015,N_36193);
or U38465 (N_38465,N_37756,N_36240);
nor U38466 (N_38466,N_37288,N_37436);
xnor U38467 (N_38467,N_36982,N_36052);
or U38468 (N_38468,N_36887,N_36892);
xor U38469 (N_38469,N_37186,N_36786);
nand U38470 (N_38470,N_37902,N_37527);
xor U38471 (N_38471,N_36229,N_37374);
or U38472 (N_38472,N_36156,N_36157);
nand U38473 (N_38473,N_37319,N_37973);
or U38474 (N_38474,N_37197,N_37075);
nand U38475 (N_38475,N_37066,N_36958);
xnor U38476 (N_38476,N_36771,N_37112);
or U38477 (N_38477,N_36571,N_37208);
nor U38478 (N_38478,N_36694,N_36210);
or U38479 (N_38479,N_36606,N_36287);
nor U38480 (N_38480,N_36843,N_36697);
or U38481 (N_38481,N_36133,N_37270);
xor U38482 (N_38482,N_36332,N_37013);
xor U38483 (N_38483,N_37313,N_36489);
or U38484 (N_38484,N_37380,N_37239);
nand U38485 (N_38485,N_36099,N_37410);
nor U38486 (N_38486,N_36092,N_36054);
nand U38487 (N_38487,N_36624,N_36603);
xor U38488 (N_38488,N_36879,N_37993);
and U38489 (N_38489,N_36824,N_36508);
nor U38490 (N_38490,N_37029,N_37330);
or U38491 (N_38491,N_36234,N_36341);
nor U38492 (N_38492,N_36888,N_36080);
or U38493 (N_38493,N_36003,N_36407);
nor U38494 (N_38494,N_36244,N_37423);
nand U38495 (N_38495,N_36594,N_37472);
xnor U38496 (N_38496,N_36850,N_36350);
or U38497 (N_38497,N_37187,N_37189);
nand U38498 (N_38498,N_36510,N_37950);
nand U38499 (N_38499,N_36218,N_36564);
xor U38500 (N_38500,N_37602,N_36359);
xnor U38501 (N_38501,N_36909,N_37940);
or U38502 (N_38502,N_36181,N_36416);
and U38503 (N_38503,N_37444,N_36214);
or U38504 (N_38504,N_36577,N_36344);
or U38505 (N_38505,N_37194,N_37591);
nand U38506 (N_38506,N_36993,N_37519);
nor U38507 (N_38507,N_36981,N_37717);
or U38508 (N_38508,N_36589,N_37391);
xnor U38509 (N_38509,N_36770,N_36280);
xor U38510 (N_38510,N_37278,N_36629);
or U38511 (N_38511,N_37577,N_37064);
or U38512 (N_38512,N_37833,N_36165);
xor U38513 (N_38513,N_36562,N_37133);
xor U38514 (N_38514,N_37358,N_37434);
or U38515 (N_38515,N_37298,N_36118);
nor U38516 (N_38516,N_37990,N_37300);
xnor U38517 (N_38517,N_37052,N_37286);
xnor U38518 (N_38518,N_36749,N_37236);
and U38519 (N_38519,N_36716,N_36803);
and U38520 (N_38520,N_37493,N_37285);
xor U38521 (N_38521,N_36039,N_37389);
nand U38522 (N_38522,N_37171,N_37515);
xnor U38523 (N_38523,N_36531,N_36186);
and U38524 (N_38524,N_36840,N_37938);
and U38525 (N_38525,N_37582,N_36070);
xor U38526 (N_38526,N_36425,N_36634);
nand U38527 (N_38527,N_37721,N_37501);
nand U38528 (N_38528,N_37218,N_37966);
nor U38529 (N_38529,N_37109,N_37617);
xor U38530 (N_38530,N_36705,N_36619);
nor U38531 (N_38531,N_37176,N_37364);
or U38532 (N_38532,N_37791,N_37326);
nand U38533 (N_38533,N_36263,N_37007);
xor U38534 (N_38534,N_36346,N_36747);
and U38535 (N_38535,N_36943,N_36660);
or U38536 (N_38536,N_36044,N_37649);
or U38537 (N_38537,N_37704,N_37587);
or U38538 (N_38538,N_36042,N_37098);
xor U38539 (N_38539,N_36131,N_37135);
xor U38540 (N_38540,N_37469,N_36791);
and U38541 (N_38541,N_37427,N_36622);
nand U38542 (N_38542,N_36757,N_36860);
nand U38543 (N_38543,N_36105,N_36375);
or U38544 (N_38544,N_36520,N_37425);
and U38545 (N_38545,N_36807,N_37365);
or U38546 (N_38546,N_36597,N_36276);
and U38547 (N_38547,N_37139,N_36075);
nor U38548 (N_38548,N_36805,N_36659);
xnor U38549 (N_38549,N_36617,N_36992);
nand U38550 (N_38550,N_36675,N_36699);
and U38551 (N_38551,N_36470,N_36309);
xor U38552 (N_38552,N_36760,N_37084);
nand U38553 (N_38553,N_37491,N_37688);
xnor U38554 (N_38554,N_36620,N_37217);
nand U38555 (N_38555,N_37823,N_37561);
or U38556 (N_38556,N_37671,N_37633);
xnor U38557 (N_38557,N_37528,N_37509);
or U38558 (N_38558,N_36647,N_36959);
nor U38559 (N_38559,N_37274,N_36657);
nor U38560 (N_38560,N_37772,N_36471);
nor U38561 (N_38561,N_36360,N_36365);
xnor U38562 (N_38562,N_37941,N_37525);
or U38563 (N_38563,N_37408,N_36961);
nand U38564 (N_38564,N_37809,N_36372);
xnor U38565 (N_38565,N_37450,N_36059);
nor U38566 (N_38566,N_36415,N_37415);
or U38567 (N_38567,N_36178,N_36155);
and U38568 (N_38568,N_36667,N_36711);
or U38569 (N_38569,N_36049,N_37401);
nand U38570 (N_38570,N_37894,N_37889);
and U38571 (N_38571,N_37867,N_36802);
xor U38572 (N_38572,N_37463,N_36402);
nand U38573 (N_38573,N_36322,N_37352);
xor U38574 (N_38574,N_37422,N_36088);
xor U38575 (N_38575,N_37122,N_36221);
xnor U38576 (N_38576,N_37619,N_37513);
xnor U38577 (N_38577,N_36698,N_37459);
xor U38578 (N_38578,N_36742,N_36393);
nor U38579 (N_38579,N_37650,N_36876);
or U38580 (N_38580,N_36700,N_36701);
or U38581 (N_38581,N_37492,N_36905);
and U38582 (N_38582,N_37572,N_36819);
nor U38583 (N_38583,N_37689,N_37053);
xnor U38584 (N_38584,N_36829,N_37174);
xnor U38585 (N_38585,N_37283,N_36061);
nand U38586 (N_38586,N_37730,N_36965);
or U38587 (N_38587,N_37564,N_36072);
xnor U38588 (N_38588,N_36012,N_36765);
nand U38589 (N_38589,N_37657,N_37787);
xor U38590 (N_38590,N_37447,N_37027);
nor U38591 (N_38591,N_37257,N_37233);
nor U38592 (N_38592,N_36774,N_36314);
and U38593 (N_38593,N_36540,N_36730);
nand U38594 (N_38594,N_37839,N_36623);
nand U38595 (N_38595,N_37840,N_37520);
or U38596 (N_38596,N_36831,N_37884);
nand U38597 (N_38597,N_36975,N_37881);
xor U38598 (N_38598,N_37842,N_37987);
nor U38599 (N_38599,N_37040,N_36847);
xnor U38600 (N_38600,N_37725,N_37111);
nor U38601 (N_38601,N_36924,N_37153);
and U38602 (N_38602,N_37729,N_37662);
nand U38603 (N_38603,N_36001,N_37035);
and U38604 (N_38604,N_36736,N_37998);
and U38605 (N_38605,N_36613,N_37846);
or U38606 (N_38606,N_36953,N_37069);
or U38607 (N_38607,N_37790,N_37831);
or U38608 (N_38608,N_36517,N_37850);
nand U38609 (N_38609,N_36704,N_36628);
nor U38610 (N_38610,N_37558,N_37481);
nand U38611 (N_38611,N_37290,N_37226);
nand U38612 (N_38612,N_36527,N_37855);
or U38613 (N_38613,N_36188,N_36392);
nand U38614 (N_38614,N_36295,N_37888);
or U38615 (N_38615,N_36267,N_37594);
nor U38616 (N_38616,N_36651,N_36548);
and U38617 (N_38617,N_36145,N_36047);
xor U38618 (N_38618,N_36672,N_37014);
and U38619 (N_38619,N_37868,N_36007);
and U38620 (N_38620,N_37996,N_37807);
nand U38621 (N_38621,N_37663,N_36025);
nand U38622 (N_38622,N_36265,N_37570);
nand U38623 (N_38623,N_36519,N_36768);
nor U38624 (N_38624,N_37665,N_36561);
or U38625 (N_38625,N_37822,N_36448);
xnor U38626 (N_38626,N_37536,N_36769);
xor U38627 (N_38627,N_37609,N_37118);
xnor U38628 (N_38628,N_36873,N_37407);
or U38629 (N_38629,N_37813,N_37644);
xor U38630 (N_38630,N_36283,N_37051);
xor U38631 (N_38631,N_37050,N_37698);
nand U38632 (N_38632,N_37488,N_37872);
and U38633 (N_38633,N_36278,N_37383);
nor U38634 (N_38634,N_36067,N_36911);
nand U38635 (N_38635,N_36788,N_37238);
xnor U38636 (N_38636,N_36935,N_37593);
or U38637 (N_38637,N_37266,N_36967);
xnor U38638 (N_38638,N_36669,N_37351);
xor U38639 (N_38639,N_36852,N_37017);
xor U38640 (N_38640,N_37936,N_36257);
or U38641 (N_38641,N_37545,N_36607);
or U38642 (N_38642,N_37163,N_36147);
xnor U38643 (N_38643,N_36590,N_37155);
or U38644 (N_38644,N_37110,N_37724);
nor U38645 (N_38645,N_36260,N_36979);
nand U38646 (N_38646,N_36550,N_36546);
nand U38647 (N_38647,N_37885,N_37985);
xnor U38648 (N_38648,N_36311,N_36858);
and U38649 (N_38649,N_37988,N_36947);
nor U38650 (N_38650,N_36759,N_36515);
nand U38651 (N_38651,N_36183,N_37925);
nand U38652 (N_38652,N_36174,N_36585);
or U38653 (N_38653,N_36286,N_36756);
nand U38654 (N_38654,N_36964,N_37200);
or U38655 (N_38655,N_37161,N_37843);
nor U38656 (N_38656,N_37544,N_37005);
nor U38657 (N_38657,N_37959,N_37853);
or U38658 (N_38658,N_37907,N_36972);
or U38659 (N_38659,N_37723,N_36207);
nor U38660 (N_38660,N_36764,N_36212);
or U38661 (N_38661,N_37262,N_37750);
xnor U38662 (N_38662,N_36401,N_37495);
nand U38663 (N_38663,N_37984,N_37245);
nor U38664 (N_38664,N_36678,N_37627);
and U38665 (N_38665,N_37271,N_36417);
or U38666 (N_38666,N_37777,N_37934);
or U38667 (N_38667,N_36865,N_37754);
and U38668 (N_38668,N_37590,N_36734);
nor U38669 (N_38669,N_37360,N_37886);
and U38670 (N_38670,N_37343,N_37466);
or U38671 (N_38671,N_36722,N_37699);
nand U38672 (N_38672,N_36299,N_36397);
nor U38673 (N_38673,N_36674,N_37403);
nor U38674 (N_38674,N_37847,N_37969);
nand U38675 (N_38675,N_36312,N_36497);
and U38676 (N_38676,N_37734,N_36396);
and U38677 (N_38677,N_37763,N_37901);
or U38678 (N_38678,N_37816,N_37100);
xor U38679 (N_38679,N_36592,N_37476);
xnor U38680 (N_38680,N_36558,N_36250);
xnor U38681 (N_38681,N_37022,N_37143);
and U38682 (N_38682,N_36379,N_37054);
and U38683 (N_38683,N_37230,N_37406);
nand U38684 (N_38684,N_37072,N_37986);
nor U38685 (N_38685,N_37632,N_37761);
nor U38686 (N_38686,N_37522,N_36922);
nor U38687 (N_38687,N_37611,N_36626);
or U38688 (N_38688,N_37097,N_36810);
nand U38689 (N_38689,N_37728,N_36503);
and U38690 (N_38690,N_36428,N_36833);
nor U38691 (N_38691,N_36921,N_37909);
nand U38692 (N_38692,N_37805,N_36985);
and U38693 (N_38693,N_36988,N_36136);
nand U38694 (N_38694,N_37359,N_37184);
or U38695 (N_38695,N_36213,N_36410);
nand U38696 (N_38696,N_37323,N_37857);
and U38697 (N_38697,N_36894,N_37937);
xnor U38698 (N_38698,N_37325,N_36021);
nor U38699 (N_38699,N_37129,N_37747);
or U38700 (N_38700,N_37771,N_37543);
nand U38701 (N_38701,N_36362,N_37999);
or U38702 (N_38702,N_37152,N_37011);
and U38703 (N_38703,N_37575,N_37248);
nor U38704 (N_38704,N_36530,N_37067);
nor U38705 (N_38705,N_36692,N_36000);
nor U38706 (N_38706,N_36813,N_37535);
nor U38707 (N_38707,N_37227,N_37312);
nor U38708 (N_38708,N_37751,N_37267);
nand U38709 (N_38709,N_37929,N_36144);
and U38710 (N_38710,N_37955,N_36708);
xor U38711 (N_38711,N_37836,N_36355);
nand U38712 (N_38712,N_37895,N_36556);
or U38713 (N_38713,N_37641,N_36853);
nand U38714 (N_38714,N_37136,N_37490);
and U38715 (N_38715,N_36621,N_37555);
xnor U38716 (N_38716,N_37547,N_36412);
and U38717 (N_38717,N_37904,N_36184);
and U38718 (N_38718,N_36575,N_37854);
nand U38719 (N_38719,N_37453,N_36804);
nand U38720 (N_38720,N_36146,N_37132);
nand U38721 (N_38721,N_36960,N_36602);
or U38722 (N_38722,N_37782,N_36671);
xnor U38723 (N_38723,N_36345,N_36891);
nand U38724 (N_38724,N_36081,N_36738);
nand U38725 (N_38725,N_37637,N_37675);
nor U38726 (N_38726,N_36631,N_37701);
nand U38727 (N_38727,N_36106,N_37414);
and U38728 (N_38728,N_36349,N_36939);
or U38729 (N_38729,N_36854,N_37457);
and U38730 (N_38730,N_36533,N_36673);
nand U38731 (N_38731,N_37759,N_37180);
and U38732 (N_38732,N_36495,N_36896);
xor U38733 (N_38733,N_36380,N_37864);
and U38734 (N_38734,N_37652,N_37769);
and U38735 (N_38735,N_37076,N_36437);
xor U38736 (N_38736,N_37260,N_37574);
nor U38737 (N_38737,N_37508,N_37658);
and U38738 (N_38738,N_37686,N_37672);
xnor U38739 (N_38739,N_37829,N_37661);
and U38740 (N_38740,N_36029,N_37045);
xor U38741 (N_38741,N_36444,N_36325);
nand U38742 (N_38742,N_37659,N_36822);
and U38743 (N_38743,N_36492,N_37625);
nand U38744 (N_38744,N_37455,N_36168);
nand U38745 (N_38745,N_36033,N_37957);
and U38746 (N_38746,N_36605,N_36496);
xor U38747 (N_38747,N_36902,N_36851);
nand U38748 (N_38748,N_37932,N_36601);
nand U38749 (N_38749,N_36584,N_37026);
and U38750 (N_38750,N_36481,N_37898);
nand U38751 (N_38751,N_37215,N_37584);
nor U38752 (N_38752,N_36832,N_36035);
or U38753 (N_38753,N_37953,N_37533);
and U38754 (N_38754,N_37329,N_36331);
xnor U38755 (N_38755,N_36129,N_37078);
or U38756 (N_38756,N_36275,N_37009);
and U38757 (N_38757,N_37023,N_36806);
or U38758 (N_38758,N_37516,N_37776);
xor U38759 (N_38759,N_36997,N_37253);
nand U38760 (N_38760,N_36522,N_36405);
nor U38761 (N_38761,N_36991,N_37080);
nand U38762 (N_38762,N_36762,N_37458);
nand U38763 (N_38763,N_37830,N_37038);
or U38764 (N_38764,N_37177,N_36456);
nand U38765 (N_38765,N_37824,N_37273);
nor U38766 (N_38766,N_37980,N_36290);
or U38767 (N_38767,N_36718,N_37773);
or U38768 (N_38768,N_37039,N_37198);
xor U38769 (N_38769,N_37172,N_36486);
nand U38770 (N_38770,N_36856,N_37237);
xnor U38771 (N_38771,N_36957,N_37376);
nand U38772 (N_38772,N_36010,N_37355);
nand U38773 (N_38773,N_36906,N_36506);
xnor U38774 (N_38774,N_36018,N_36848);
nor U38775 (N_38775,N_37413,N_36980);
nor U38776 (N_38776,N_36467,N_37195);
nor U38777 (N_38777,N_36385,N_37645);
or U38778 (N_38778,N_36766,N_36938);
or U38779 (N_38779,N_37677,N_36301);
nor U38780 (N_38780,N_37802,N_37817);
xor U38781 (N_38781,N_37511,N_36925);
nor U38782 (N_38782,N_36189,N_36256);
xor U38783 (N_38783,N_37873,N_36910);
nor U38784 (N_38784,N_36767,N_36343);
xnor U38785 (N_38785,N_37647,N_37882);
or U38786 (N_38786,N_36857,N_37446);
nor U38787 (N_38787,N_37654,N_37396);
nand U38788 (N_38788,N_37589,N_37090);
and U38789 (N_38789,N_37115,N_37398);
or U38790 (N_38790,N_36017,N_37345);
or U38791 (N_38791,N_37235,N_37964);
nand U38792 (N_38792,N_37297,N_36518);
xor U38793 (N_38793,N_36818,N_36090);
xnor U38794 (N_38794,N_37196,N_37128);
and U38795 (N_38795,N_37385,N_36532);
and U38796 (N_38796,N_36710,N_37971);
nand U38797 (N_38797,N_36262,N_37968);
nand U38798 (N_38798,N_37301,N_37036);
xor U38799 (N_38799,N_36717,N_36491);
xor U38800 (N_38800,N_36474,N_37010);
nand U38801 (N_38801,N_37317,N_36439);
and U38802 (N_38802,N_37483,N_37454);
nand U38803 (N_38803,N_36493,N_36501);
nor U38804 (N_38804,N_36727,N_36102);
nand U38805 (N_38805,N_36468,N_36745);
xnor U38806 (N_38806,N_36371,N_37229);
and U38807 (N_38807,N_37792,N_37284);
and U38808 (N_38808,N_36289,N_36464);
nand U38809 (N_38809,N_36057,N_37314);
and U38810 (N_38810,N_37055,N_36112);
xor U38811 (N_38811,N_37610,N_37656);
xnor U38812 (N_38812,N_37254,N_37642);
nand U38813 (N_38813,N_36775,N_36143);
or U38814 (N_38814,N_37397,N_37646);
and U38815 (N_38815,N_36785,N_36169);
nor U38816 (N_38816,N_36264,N_37588);
nor U38817 (N_38817,N_37956,N_37124);
nand U38818 (N_38818,N_36845,N_37307);
or U38819 (N_38819,N_36445,N_37178);
nor U38820 (N_38820,N_37390,N_36904);
nand U38821 (N_38821,N_37624,N_37930);
or U38822 (N_38822,N_36755,N_37222);
nor U38823 (N_38823,N_36912,N_37702);
or U38824 (N_38824,N_36889,N_37321);
or U38825 (N_38825,N_36494,N_36107);
nor U38826 (N_38826,N_36573,N_36908);
and U38827 (N_38827,N_36122,N_37921);
nand U38828 (N_38828,N_36790,N_36422);
xnor U38829 (N_38829,N_36427,N_36801);
nand U38830 (N_38830,N_37532,N_36135);
or U38831 (N_38831,N_36163,N_36797);
or U38832 (N_38832,N_36006,N_36796);
nor U38833 (N_38833,N_37256,N_36294);
and U38834 (N_38834,N_37471,N_37919);
xor U38835 (N_38835,N_36348,N_37695);
xor U38836 (N_38836,N_37006,N_36990);
or U38837 (N_38837,N_36389,N_37531);
nand U38838 (N_38838,N_37467,N_36337);
or U38839 (N_38839,N_36731,N_37741);
or U38840 (N_38840,N_37336,N_37595);
nand U38841 (N_38841,N_37037,N_36553);
or U38842 (N_38842,N_37798,N_37826);
or U38843 (N_38843,N_36031,N_36828);
xnor U38844 (N_38844,N_37393,N_36215);
nand U38845 (N_38845,N_36524,N_36279);
and U38846 (N_38846,N_36454,N_36113);
xor U38847 (N_38847,N_37541,N_37550);
and U38848 (N_38848,N_37125,N_37982);
and U38849 (N_38849,N_36447,N_36574);
nand U38850 (N_38850,N_37598,N_37848);
nand U38851 (N_38851,N_36883,N_37316);
or U38852 (N_38852,N_36028,N_36679);
xor U38853 (N_38853,N_37368,N_37165);
or U38854 (N_38854,N_36869,N_37585);
xnor U38855 (N_38855,N_36735,N_36233);
xor U38856 (N_38856,N_37529,N_36227);
nor U38857 (N_38857,N_36223,N_37089);
xor U38858 (N_38858,N_36662,N_37562);
and U38859 (N_38859,N_37327,N_36132);
and U38860 (N_38860,N_36627,N_36693);
and U38861 (N_38861,N_37737,N_36100);
or U38862 (N_38862,N_37849,N_36151);
and U38863 (N_38863,N_36695,N_37071);
xor U38864 (N_38864,N_36440,N_36101);
and U38865 (N_38865,N_37179,N_37709);
nor U38866 (N_38866,N_36569,N_37224);
xor U38867 (N_38867,N_37305,N_36638);
or U38868 (N_38868,N_36514,N_36190);
nor U38869 (N_38869,N_36900,N_36252);
xor U38870 (N_38870,N_37673,N_36560);
or U38871 (N_38871,N_36037,N_37972);
nor U38872 (N_38872,N_36542,N_37615);
nor U38873 (N_38873,N_37295,N_36241);
nand U38874 (N_38874,N_36543,N_37083);
nand U38875 (N_38875,N_37318,N_36984);
or U38876 (N_38876,N_37648,N_37473);
xor U38877 (N_38877,N_37814,N_36554);
or U38878 (N_38878,N_37292,N_37716);
nor U38879 (N_38879,N_37004,N_36614);
nand U38880 (N_38880,N_37880,N_37268);
or U38881 (N_38881,N_37819,N_36746);
nand U38882 (N_38882,N_36946,N_37497);
and U38883 (N_38883,N_36128,N_37405);
nor U38884 (N_38884,N_36884,N_36652);
nor U38885 (N_38885,N_37507,N_36247);
nor U38886 (N_38886,N_37795,N_36655);
nand U38887 (N_38887,N_37746,N_37960);
or U38888 (N_38888,N_37742,N_37362);
and U38889 (N_38889,N_37095,N_37828);
or U38890 (N_38890,N_36604,N_37524);
or U38891 (N_38891,N_37510,N_37464);
or U38892 (N_38892,N_36625,N_37825);
xor U38893 (N_38893,N_36161,N_37016);
and U38894 (N_38894,N_37596,N_36282);
and U38895 (N_38895,N_36490,N_37549);
nand U38896 (N_38896,N_36258,N_36596);
and U38897 (N_38897,N_36009,N_37142);
and U38898 (N_38898,N_37962,N_36557);
xor U38899 (N_38899,N_37116,N_37563);
or U38900 (N_38900,N_36370,N_36976);
or U38901 (N_38901,N_36937,N_36539);
xor U38902 (N_38902,N_37696,N_37201);
and U38903 (N_38903,N_37082,N_36689);
xnor U38904 (N_38904,N_36171,N_37154);
or U38905 (N_38905,N_36436,N_36591);
nand U38906 (N_38906,N_36983,N_36140);
or U38907 (N_38907,N_37310,N_36022);
or U38908 (N_38908,N_36431,N_36297);
nor U38909 (N_38909,N_36177,N_36502);
or U38910 (N_38910,N_37815,N_36109);
nand U38911 (N_38911,N_36201,N_36995);
nor U38912 (N_38912,N_37294,N_37269);
nor U38913 (N_38913,N_37431,N_36306);
and U38914 (N_38914,N_37140,N_36509);
and U38915 (N_38915,N_36987,N_36326);
nand U38916 (N_38916,N_37945,N_36862);
xor U38917 (N_38917,N_36773,N_37168);
nor U38918 (N_38918,N_36583,N_37691);
nor U38919 (N_38919,N_36053,N_37057);
nand U38920 (N_38920,N_36418,N_37223);
nor U38921 (N_38921,N_36516,N_36160);
xnor U38922 (N_38922,N_36091,N_37961);
nor U38923 (N_38923,N_37503,N_37188);
nor U38924 (N_38924,N_36684,N_37911);
nor U38925 (N_38925,N_36565,N_37296);
or U38926 (N_38926,N_36653,N_36232);
xor U38927 (N_38927,N_36073,N_36150);
xor U38928 (N_38928,N_37032,N_36406);
nand U38929 (N_38929,N_37856,N_37774);
nor U38930 (N_38930,N_36645,N_36206);
and U38931 (N_38931,N_36443,N_36111);
nor U38932 (N_38932,N_36034,N_36376);
nor U38933 (N_38933,N_36013,N_36929);
or U38934 (N_38934,N_37249,N_37147);
and U38935 (N_38935,N_37788,N_37402);
nor U38936 (N_38936,N_36224,N_36153);
nor U38937 (N_38937,N_37441,N_37456);
and U38938 (N_38938,N_37785,N_37117);
or U38939 (N_38939,N_36011,N_36996);
nand U38940 (N_38940,N_36725,N_37748);
nor U38941 (N_38941,N_36387,N_36317);
xor U38942 (N_38942,N_37331,N_37651);
nand U38943 (N_38943,N_37499,N_37258);
xor U38944 (N_38944,N_37190,N_37388);
and U38945 (N_38945,N_36855,N_36572);
xnor U38946 (N_38946,N_36595,N_36121);
nor U38947 (N_38947,N_36268,N_37687);
nor U38948 (N_38948,N_36116,N_36382);
or U38949 (N_38949,N_36056,N_37277);
and U38950 (N_38950,N_37308,N_37145);
and U38951 (N_38951,N_37049,N_37674);
nor U38952 (N_38952,N_36066,N_36842);
nand U38953 (N_38953,N_36446,N_36411);
nand U38954 (N_38954,N_36203,N_36777);
nand U38955 (N_38955,N_36304,N_37668);
xnor U38956 (N_38956,N_36677,N_36318);
nand U38957 (N_38957,N_37979,N_36881);
xor U38958 (N_38958,N_37101,N_37293);
or U38959 (N_38959,N_36269,N_37970);
nor U38960 (N_38960,N_36027,N_36180);
nand U38961 (N_38961,N_36084,N_36640);
or U38962 (N_38962,N_36952,N_36951);
and U38963 (N_38963,N_36087,N_37500);
xor U38964 (N_38964,N_37448,N_36488);
and U38965 (N_38965,N_36419,N_37976);
or U38966 (N_38966,N_36429,N_36014);
and U38967 (N_38967,N_37942,N_36019);
nand U38968 (N_38968,N_37712,N_36942);
nand U38969 (N_38969,N_36063,N_37664);
and U38970 (N_38970,N_36815,N_37514);
nor U38971 (N_38971,N_37247,N_37357);
nor U38972 (N_38972,N_37470,N_36409);
xnor U38973 (N_38973,N_36523,N_36691);
nor U38974 (N_38974,N_36598,N_37068);
or U38975 (N_38975,N_37683,N_37732);
and U38976 (N_38976,N_36914,N_36432);
nand U38977 (N_38977,N_37726,N_36246);
or U38978 (N_38978,N_36743,N_36159);
or U38979 (N_38979,N_36465,N_37523);
or U38980 (N_38980,N_37485,N_36841);
or U38981 (N_38981,N_37449,N_36209);
nand U38982 (N_38982,N_36687,N_36820);
nor U38983 (N_38983,N_37779,N_36944);
xnor U38984 (N_38984,N_36754,N_36333);
or U38985 (N_38985,N_36347,N_36724);
and U38986 (N_38986,N_37299,N_37228);
nor U38987 (N_38987,N_37018,N_36235);
nand U38988 (N_38988,N_37818,N_37866);
nand U38989 (N_38989,N_36578,N_36487);
nor U38990 (N_38990,N_37219,N_37264);
or U38991 (N_38991,N_36950,N_36549);
and U38992 (N_38992,N_36861,N_37242);
and U38993 (N_38993,N_36945,N_37565);
nor U38994 (N_38994,N_37851,N_37384);
or U38995 (N_38995,N_36065,N_36643);
nand U38996 (N_38996,N_36020,N_37923);
and U38997 (N_38997,N_36281,N_36220);
nor U38998 (N_38998,N_36913,N_36882);
nor U38999 (N_38999,N_37653,N_37607);
or U39000 (N_39000,N_36356,N_37894);
nor U39001 (N_39001,N_37518,N_37816);
xor U39002 (N_39002,N_36523,N_36973);
and U39003 (N_39003,N_37780,N_37136);
and U39004 (N_39004,N_37370,N_36754);
nor U39005 (N_39005,N_36804,N_37025);
nor U39006 (N_39006,N_37455,N_36108);
and U39007 (N_39007,N_37669,N_36684);
xnor U39008 (N_39008,N_37214,N_36569);
nand U39009 (N_39009,N_36859,N_36000);
or U39010 (N_39010,N_37908,N_36098);
and U39011 (N_39011,N_37930,N_36770);
or U39012 (N_39012,N_36965,N_37426);
or U39013 (N_39013,N_37232,N_36861);
nor U39014 (N_39014,N_37224,N_36226);
xnor U39015 (N_39015,N_37372,N_36365);
or U39016 (N_39016,N_36704,N_36868);
xor U39017 (N_39017,N_36177,N_37147);
nor U39018 (N_39018,N_36311,N_36851);
nand U39019 (N_39019,N_36158,N_36343);
or U39020 (N_39020,N_36916,N_36504);
xor U39021 (N_39021,N_37312,N_37843);
nand U39022 (N_39022,N_36605,N_36136);
xnor U39023 (N_39023,N_36660,N_36786);
nor U39024 (N_39024,N_36904,N_36039);
xor U39025 (N_39025,N_37777,N_36799);
nor U39026 (N_39026,N_37908,N_37710);
and U39027 (N_39027,N_36807,N_36052);
nor U39028 (N_39028,N_36827,N_36637);
and U39029 (N_39029,N_36279,N_37534);
xor U39030 (N_39030,N_36864,N_36064);
nor U39031 (N_39031,N_37397,N_37106);
nand U39032 (N_39032,N_37630,N_36156);
xor U39033 (N_39033,N_36412,N_37891);
xnor U39034 (N_39034,N_37871,N_36424);
and U39035 (N_39035,N_36173,N_36940);
nor U39036 (N_39036,N_37950,N_36879);
and U39037 (N_39037,N_37597,N_37814);
nand U39038 (N_39038,N_36443,N_37789);
and U39039 (N_39039,N_36711,N_37285);
or U39040 (N_39040,N_36529,N_37868);
xnor U39041 (N_39041,N_36733,N_37188);
and U39042 (N_39042,N_37439,N_37288);
or U39043 (N_39043,N_37493,N_36329);
and U39044 (N_39044,N_36699,N_37992);
and U39045 (N_39045,N_36581,N_37199);
nand U39046 (N_39046,N_37886,N_36149);
xnor U39047 (N_39047,N_36616,N_37812);
nand U39048 (N_39048,N_36960,N_37549);
nand U39049 (N_39049,N_37535,N_37407);
and U39050 (N_39050,N_36864,N_37412);
and U39051 (N_39051,N_36221,N_37424);
nor U39052 (N_39052,N_37443,N_37529);
and U39053 (N_39053,N_37032,N_37298);
or U39054 (N_39054,N_36899,N_37863);
and U39055 (N_39055,N_37673,N_36184);
nor U39056 (N_39056,N_37338,N_36288);
or U39057 (N_39057,N_37717,N_36060);
nand U39058 (N_39058,N_36286,N_37537);
xnor U39059 (N_39059,N_37337,N_36566);
nor U39060 (N_39060,N_37101,N_37879);
nor U39061 (N_39061,N_37223,N_37772);
nor U39062 (N_39062,N_36119,N_36089);
nand U39063 (N_39063,N_36390,N_36725);
xor U39064 (N_39064,N_36003,N_36117);
nor U39065 (N_39065,N_36632,N_37711);
nor U39066 (N_39066,N_37584,N_36162);
nand U39067 (N_39067,N_36490,N_36542);
and U39068 (N_39068,N_36210,N_37832);
or U39069 (N_39069,N_36744,N_37323);
and U39070 (N_39070,N_36807,N_37662);
xor U39071 (N_39071,N_36292,N_37431);
nor U39072 (N_39072,N_37408,N_36584);
or U39073 (N_39073,N_36324,N_36430);
and U39074 (N_39074,N_37516,N_37624);
nor U39075 (N_39075,N_37386,N_36021);
or U39076 (N_39076,N_37491,N_37026);
nor U39077 (N_39077,N_36171,N_36442);
nand U39078 (N_39078,N_37824,N_37213);
and U39079 (N_39079,N_37403,N_37399);
nand U39080 (N_39080,N_37861,N_37055);
or U39081 (N_39081,N_36507,N_36763);
or U39082 (N_39082,N_36594,N_37273);
or U39083 (N_39083,N_37323,N_36111);
and U39084 (N_39084,N_36601,N_36566);
nor U39085 (N_39085,N_36451,N_37971);
or U39086 (N_39086,N_37144,N_37393);
and U39087 (N_39087,N_37959,N_36978);
nand U39088 (N_39088,N_36273,N_36199);
nor U39089 (N_39089,N_36121,N_36572);
and U39090 (N_39090,N_37147,N_36518);
or U39091 (N_39091,N_36439,N_36727);
nor U39092 (N_39092,N_36523,N_36308);
or U39093 (N_39093,N_36679,N_37274);
nand U39094 (N_39094,N_37157,N_37603);
nand U39095 (N_39095,N_37220,N_36977);
and U39096 (N_39096,N_37155,N_37447);
nor U39097 (N_39097,N_36994,N_36741);
xnor U39098 (N_39098,N_37144,N_37655);
or U39099 (N_39099,N_36610,N_37779);
xnor U39100 (N_39100,N_36575,N_36423);
nor U39101 (N_39101,N_37593,N_37090);
xnor U39102 (N_39102,N_37070,N_36558);
nor U39103 (N_39103,N_36134,N_36565);
nand U39104 (N_39104,N_37314,N_37915);
xnor U39105 (N_39105,N_36212,N_37446);
xnor U39106 (N_39106,N_37618,N_36657);
or U39107 (N_39107,N_36388,N_37403);
or U39108 (N_39108,N_37009,N_36478);
nand U39109 (N_39109,N_37728,N_37957);
nand U39110 (N_39110,N_37130,N_36124);
and U39111 (N_39111,N_36453,N_36695);
nand U39112 (N_39112,N_36757,N_37240);
nor U39113 (N_39113,N_36414,N_36059);
and U39114 (N_39114,N_36560,N_36052);
and U39115 (N_39115,N_37958,N_37106);
and U39116 (N_39116,N_37806,N_37230);
nor U39117 (N_39117,N_36686,N_37685);
and U39118 (N_39118,N_37343,N_36989);
nor U39119 (N_39119,N_37439,N_36142);
nor U39120 (N_39120,N_37186,N_36834);
nor U39121 (N_39121,N_37548,N_37972);
xor U39122 (N_39122,N_36123,N_37072);
nor U39123 (N_39123,N_37486,N_36084);
nand U39124 (N_39124,N_37565,N_36304);
or U39125 (N_39125,N_37513,N_37249);
and U39126 (N_39126,N_36408,N_36895);
xnor U39127 (N_39127,N_36961,N_36590);
and U39128 (N_39128,N_36841,N_37388);
xnor U39129 (N_39129,N_37506,N_36939);
and U39130 (N_39130,N_36819,N_36146);
nor U39131 (N_39131,N_36843,N_37111);
nand U39132 (N_39132,N_37029,N_36873);
nand U39133 (N_39133,N_36388,N_36134);
or U39134 (N_39134,N_37791,N_36456);
or U39135 (N_39135,N_36640,N_36167);
and U39136 (N_39136,N_36182,N_37604);
nand U39137 (N_39137,N_36368,N_36937);
nor U39138 (N_39138,N_36551,N_37025);
nand U39139 (N_39139,N_37510,N_36604);
nor U39140 (N_39140,N_36200,N_37839);
or U39141 (N_39141,N_36944,N_36789);
nor U39142 (N_39142,N_36086,N_36040);
and U39143 (N_39143,N_36941,N_36769);
nand U39144 (N_39144,N_36469,N_36145);
or U39145 (N_39145,N_36783,N_37913);
nand U39146 (N_39146,N_37661,N_37719);
xnor U39147 (N_39147,N_37403,N_36235);
and U39148 (N_39148,N_36491,N_36942);
and U39149 (N_39149,N_37101,N_37584);
nand U39150 (N_39150,N_36095,N_37823);
or U39151 (N_39151,N_37066,N_37015);
nand U39152 (N_39152,N_37831,N_36795);
nand U39153 (N_39153,N_37077,N_36499);
nor U39154 (N_39154,N_36296,N_36559);
or U39155 (N_39155,N_37279,N_37547);
xor U39156 (N_39156,N_37195,N_36780);
nand U39157 (N_39157,N_36199,N_36718);
and U39158 (N_39158,N_37000,N_37394);
and U39159 (N_39159,N_37898,N_37384);
and U39160 (N_39160,N_36251,N_36687);
and U39161 (N_39161,N_37469,N_36547);
and U39162 (N_39162,N_36613,N_36096);
and U39163 (N_39163,N_37625,N_37342);
xor U39164 (N_39164,N_36740,N_36778);
xor U39165 (N_39165,N_37743,N_37549);
and U39166 (N_39166,N_36465,N_36544);
nand U39167 (N_39167,N_37474,N_36311);
or U39168 (N_39168,N_36568,N_37507);
or U39169 (N_39169,N_37065,N_37047);
nor U39170 (N_39170,N_36291,N_37800);
xnor U39171 (N_39171,N_36994,N_37994);
or U39172 (N_39172,N_37967,N_36350);
xor U39173 (N_39173,N_36496,N_36238);
and U39174 (N_39174,N_37733,N_37563);
and U39175 (N_39175,N_37300,N_37680);
nor U39176 (N_39176,N_37109,N_37859);
nand U39177 (N_39177,N_36153,N_36374);
and U39178 (N_39178,N_37465,N_36533);
xor U39179 (N_39179,N_36582,N_36091);
and U39180 (N_39180,N_37107,N_36042);
nand U39181 (N_39181,N_37123,N_36276);
and U39182 (N_39182,N_36358,N_37103);
xor U39183 (N_39183,N_36219,N_37823);
nand U39184 (N_39184,N_37947,N_36876);
nand U39185 (N_39185,N_36722,N_37834);
nand U39186 (N_39186,N_37306,N_36993);
xor U39187 (N_39187,N_37826,N_37767);
or U39188 (N_39188,N_36572,N_37936);
nand U39189 (N_39189,N_36937,N_36220);
nand U39190 (N_39190,N_36235,N_37124);
nor U39191 (N_39191,N_37249,N_36294);
and U39192 (N_39192,N_37015,N_37486);
or U39193 (N_39193,N_37565,N_36800);
nand U39194 (N_39194,N_36472,N_36809);
xnor U39195 (N_39195,N_36400,N_37355);
nor U39196 (N_39196,N_37287,N_37226);
or U39197 (N_39197,N_37002,N_37899);
and U39198 (N_39198,N_36687,N_36516);
and U39199 (N_39199,N_37608,N_36856);
nand U39200 (N_39200,N_36150,N_37119);
or U39201 (N_39201,N_36499,N_37099);
and U39202 (N_39202,N_36792,N_36423);
and U39203 (N_39203,N_36621,N_37524);
nor U39204 (N_39204,N_37583,N_36891);
nor U39205 (N_39205,N_36622,N_37490);
xor U39206 (N_39206,N_37271,N_36016);
and U39207 (N_39207,N_37979,N_37174);
and U39208 (N_39208,N_37000,N_37282);
or U39209 (N_39209,N_36013,N_37588);
or U39210 (N_39210,N_37191,N_37822);
nand U39211 (N_39211,N_36502,N_37802);
and U39212 (N_39212,N_36503,N_36390);
nand U39213 (N_39213,N_36494,N_37148);
xor U39214 (N_39214,N_37397,N_37026);
nand U39215 (N_39215,N_36780,N_36662);
xnor U39216 (N_39216,N_37360,N_37718);
nor U39217 (N_39217,N_37395,N_37533);
nor U39218 (N_39218,N_37313,N_37605);
or U39219 (N_39219,N_36134,N_37041);
and U39220 (N_39220,N_36333,N_37471);
xor U39221 (N_39221,N_36176,N_36942);
and U39222 (N_39222,N_37118,N_37142);
or U39223 (N_39223,N_37592,N_36584);
or U39224 (N_39224,N_37135,N_36696);
nand U39225 (N_39225,N_36763,N_36606);
nand U39226 (N_39226,N_37522,N_37138);
and U39227 (N_39227,N_36774,N_36991);
nor U39228 (N_39228,N_37106,N_36356);
and U39229 (N_39229,N_36015,N_37638);
nand U39230 (N_39230,N_36042,N_36998);
nand U39231 (N_39231,N_37155,N_37194);
nor U39232 (N_39232,N_36886,N_37444);
or U39233 (N_39233,N_36831,N_36942);
nor U39234 (N_39234,N_36983,N_37651);
and U39235 (N_39235,N_37957,N_36723);
xnor U39236 (N_39236,N_37966,N_36525);
nand U39237 (N_39237,N_37926,N_36618);
nor U39238 (N_39238,N_36684,N_37282);
and U39239 (N_39239,N_36171,N_37803);
or U39240 (N_39240,N_36543,N_36821);
and U39241 (N_39241,N_36619,N_36239);
and U39242 (N_39242,N_37596,N_36915);
or U39243 (N_39243,N_36238,N_36458);
xor U39244 (N_39244,N_37959,N_37729);
nor U39245 (N_39245,N_37519,N_37355);
nand U39246 (N_39246,N_36799,N_36125);
nand U39247 (N_39247,N_36866,N_37584);
nand U39248 (N_39248,N_36439,N_36403);
or U39249 (N_39249,N_37479,N_37654);
and U39250 (N_39250,N_37191,N_37989);
xor U39251 (N_39251,N_37279,N_36105);
and U39252 (N_39252,N_37629,N_36734);
or U39253 (N_39253,N_36377,N_36093);
nor U39254 (N_39254,N_36424,N_36535);
nand U39255 (N_39255,N_36835,N_36138);
nor U39256 (N_39256,N_36072,N_36992);
nor U39257 (N_39257,N_36924,N_36038);
or U39258 (N_39258,N_36210,N_36941);
or U39259 (N_39259,N_37933,N_36813);
and U39260 (N_39260,N_36988,N_37746);
or U39261 (N_39261,N_37014,N_37930);
and U39262 (N_39262,N_36887,N_36959);
and U39263 (N_39263,N_36324,N_36797);
and U39264 (N_39264,N_36773,N_37654);
and U39265 (N_39265,N_37994,N_36306);
nand U39266 (N_39266,N_37376,N_37210);
nand U39267 (N_39267,N_37575,N_37554);
and U39268 (N_39268,N_36576,N_36794);
nor U39269 (N_39269,N_37447,N_37778);
xor U39270 (N_39270,N_36896,N_36572);
xnor U39271 (N_39271,N_37174,N_36071);
and U39272 (N_39272,N_36114,N_36515);
xnor U39273 (N_39273,N_37029,N_37585);
nand U39274 (N_39274,N_36169,N_36643);
and U39275 (N_39275,N_36071,N_36727);
xor U39276 (N_39276,N_36099,N_37771);
nor U39277 (N_39277,N_36088,N_36413);
and U39278 (N_39278,N_36710,N_36730);
nand U39279 (N_39279,N_37503,N_36680);
xor U39280 (N_39280,N_37444,N_37116);
nand U39281 (N_39281,N_37872,N_37581);
nor U39282 (N_39282,N_36382,N_37497);
or U39283 (N_39283,N_37022,N_37081);
or U39284 (N_39284,N_36913,N_36208);
or U39285 (N_39285,N_37902,N_36398);
xor U39286 (N_39286,N_36996,N_37622);
xor U39287 (N_39287,N_36217,N_36187);
nand U39288 (N_39288,N_37721,N_36866);
xnor U39289 (N_39289,N_36250,N_36182);
nand U39290 (N_39290,N_36862,N_36085);
nor U39291 (N_39291,N_36963,N_37023);
or U39292 (N_39292,N_37376,N_37565);
nor U39293 (N_39293,N_36862,N_36116);
nand U39294 (N_39294,N_37549,N_36042);
xnor U39295 (N_39295,N_37429,N_37926);
nor U39296 (N_39296,N_36720,N_37194);
xor U39297 (N_39297,N_37391,N_37067);
or U39298 (N_39298,N_37065,N_36333);
or U39299 (N_39299,N_36287,N_37541);
or U39300 (N_39300,N_37029,N_36679);
nor U39301 (N_39301,N_36225,N_36432);
xnor U39302 (N_39302,N_36090,N_36156);
and U39303 (N_39303,N_36616,N_36458);
nor U39304 (N_39304,N_37108,N_36778);
and U39305 (N_39305,N_37331,N_36453);
or U39306 (N_39306,N_37797,N_37039);
nand U39307 (N_39307,N_36177,N_37203);
nand U39308 (N_39308,N_36727,N_37125);
xor U39309 (N_39309,N_36309,N_36515);
xnor U39310 (N_39310,N_36183,N_37974);
nand U39311 (N_39311,N_37454,N_37800);
and U39312 (N_39312,N_37646,N_37921);
xnor U39313 (N_39313,N_37602,N_37574);
nand U39314 (N_39314,N_36153,N_37480);
nand U39315 (N_39315,N_36983,N_37094);
nand U39316 (N_39316,N_37766,N_37741);
nor U39317 (N_39317,N_36699,N_36347);
xnor U39318 (N_39318,N_37912,N_36771);
nor U39319 (N_39319,N_37963,N_36809);
nand U39320 (N_39320,N_36512,N_36182);
and U39321 (N_39321,N_37812,N_37843);
nand U39322 (N_39322,N_36673,N_37524);
and U39323 (N_39323,N_37420,N_37160);
xor U39324 (N_39324,N_37696,N_36589);
nand U39325 (N_39325,N_36999,N_36851);
or U39326 (N_39326,N_36812,N_36056);
xor U39327 (N_39327,N_37724,N_36619);
and U39328 (N_39328,N_36776,N_36810);
xnor U39329 (N_39329,N_37532,N_36830);
and U39330 (N_39330,N_37476,N_36199);
and U39331 (N_39331,N_37916,N_36807);
nor U39332 (N_39332,N_37828,N_37418);
or U39333 (N_39333,N_36925,N_37336);
and U39334 (N_39334,N_37891,N_36629);
nor U39335 (N_39335,N_37476,N_37603);
xnor U39336 (N_39336,N_36318,N_36277);
xnor U39337 (N_39337,N_36828,N_37792);
and U39338 (N_39338,N_36350,N_37618);
nand U39339 (N_39339,N_36161,N_36056);
nor U39340 (N_39340,N_36564,N_36253);
and U39341 (N_39341,N_36693,N_36037);
or U39342 (N_39342,N_36463,N_36653);
and U39343 (N_39343,N_36844,N_37836);
or U39344 (N_39344,N_36933,N_36690);
xor U39345 (N_39345,N_36350,N_37806);
nor U39346 (N_39346,N_36116,N_36313);
nand U39347 (N_39347,N_37283,N_36702);
or U39348 (N_39348,N_37197,N_37969);
or U39349 (N_39349,N_37298,N_37517);
nor U39350 (N_39350,N_36503,N_37034);
nor U39351 (N_39351,N_37805,N_37669);
nor U39352 (N_39352,N_36677,N_36843);
nor U39353 (N_39353,N_37786,N_37466);
or U39354 (N_39354,N_36584,N_36489);
nand U39355 (N_39355,N_36086,N_37692);
nor U39356 (N_39356,N_36549,N_37899);
xor U39357 (N_39357,N_37876,N_36922);
or U39358 (N_39358,N_37619,N_36426);
xnor U39359 (N_39359,N_36340,N_37099);
xor U39360 (N_39360,N_36783,N_37490);
and U39361 (N_39361,N_37646,N_36819);
nor U39362 (N_39362,N_37208,N_37418);
nor U39363 (N_39363,N_36419,N_37286);
or U39364 (N_39364,N_37470,N_37787);
nand U39365 (N_39365,N_36958,N_37340);
or U39366 (N_39366,N_37120,N_37391);
or U39367 (N_39367,N_37019,N_37577);
and U39368 (N_39368,N_36714,N_37719);
nor U39369 (N_39369,N_37642,N_37119);
nand U39370 (N_39370,N_36916,N_37880);
xnor U39371 (N_39371,N_36014,N_36543);
nor U39372 (N_39372,N_37722,N_37662);
xor U39373 (N_39373,N_37553,N_37484);
xnor U39374 (N_39374,N_37792,N_37084);
xnor U39375 (N_39375,N_36791,N_37503);
xor U39376 (N_39376,N_37307,N_37243);
xor U39377 (N_39377,N_36029,N_37867);
nor U39378 (N_39378,N_36232,N_36908);
or U39379 (N_39379,N_36389,N_36650);
and U39380 (N_39380,N_37356,N_36768);
nor U39381 (N_39381,N_37763,N_37687);
or U39382 (N_39382,N_36005,N_36447);
nand U39383 (N_39383,N_37775,N_36503);
xor U39384 (N_39384,N_37695,N_36269);
and U39385 (N_39385,N_36025,N_36796);
and U39386 (N_39386,N_37880,N_37024);
nand U39387 (N_39387,N_37070,N_36561);
or U39388 (N_39388,N_36521,N_36032);
nand U39389 (N_39389,N_37391,N_37080);
and U39390 (N_39390,N_37835,N_36720);
xnor U39391 (N_39391,N_36448,N_36589);
and U39392 (N_39392,N_37327,N_37801);
nor U39393 (N_39393,N_37667,N_36514);
nor U39394 (N_39394,N_36854,N_36745);
nor U39395 (N_39395,N_37920,N_36366);
or U39396 (N_39396,N_37919,N_36858);
nor U39397 (N_39397,N_37208,N_36668);
nor U39398 (N_39398,N_37506,N_37124);
or U39399 (N_39399,N_36913,N_37819);
or U39400 (N_39400,N_36200,N_36953);
nand U39401 (N_39401,N_36592,N_37252);
nand U39402 (N_39402,N_36421,N_37721);
nor U39403 (N_39403,N_37440,N_37885);
or U39404 (N_39404,N_36216,N_37906);
xor U39405 (N_39405,N_36846,N_36872);
and U39406 (N_39406,N_36650,N_37652);
or U39407 (N_39407,N_36192,N_36588);
or U39408 (N_39408,N_36894,N_37982);
xor U39409 (N_39409,N_37893,N_36480);
and U39410 (N_39410,N_36011,N_36846);
nand U39411 (N_39411,N_36601,N_36599);
xnor U39412 (N_39412,N_36313,N_37478);
nand U39413 (N_39413,N_37911,N_36883);
and U39414 (N_39414,N_37288,N_37129);
and U39415 (N_39415,N_36022,N_37323);
xor U39416 (N_39416,N_37371,N_37883);
nor U39417 (N_39417,N_36946,N_37825);
nor U39418 (N_39418,N_37998,N_36542);
nand U39419 (N_39419,N_37378,N_37270);
and U39420 (N_39420,N_36322,N_36802);
xnor U39421 (N_39421,N_36411,N_36092);
and U39422 (N_39422,N_37534,N_37111);
xor U39423 (N_39423,N_36486,N_37863);
nand U39424 (N_39424,N_36546,N_37475);
or U39425 (N_39425,N_37916,N_36273);
xnor U39426 (N_39426,N_36208,N_36904);
xor U39427 (N_39427,N_37438,N_37645);
or U39428 (N_39428,N_36680,N_36027);
xnor U39429 (N_39429,N_36831,N_36055);
and U39430 (N_39430,N_36694,N_36953);
nand U39431 (N_39431,N_37990,N_36993);
nor U39432 (N_39432,N_37507,N_37930);
nand U39433 (N_39433,N_37325,N_37955);
or U39434 (N_39434,N_36512,N_36346);
and U39435 (N_39435,N_37114,N_37017);
xor U39436 (N_39436,N_37282,N_37752);
nand U39437 (N_39437,N_36509,N_36475);
xor U39438 (N_39438,N_37537,N_36462);
and U39439 (N_39439,N_36550,N_36673);
nor U39440 (N_39440,N_37603,N_36845);
nand U39441 (N_39441,N_36876,N_36732);
or U39442 (N_39442,N_36763,N_36301);
nor U39443 (N_39443,N_36626,N_36496);
nor U39444 (N_39444,N_36622,N_36570);
nor U39445 (N_39445,N_36660,N_36990);
xor U39446 (N_39446,N_37704,N_36261);
or U39447 (N_39447,N_36292,N_37590);
xnor U39448 (N_39448,N_36883,N_37071);
and U39449 (N_39449,N_36430,N_37092);
or U39450 (N_39450,N_37960,N_37777);
xnor U39451 (N_39451,N_37670,N_37513);
xor U39452 (N_39452,N_37637,N_37243);
xor U39453 (N_39453,N_37929,N_37705);
and U39454 (N_39454,N_36848,N_37739);
xor U39455 (N_39455,N_37678,N_37278);
nand U39456 (N_39456,N_37843,N_37187);
nand U39457 (N_39457,N_37667,N_37567);
nor U39458 (N_39458,N_37084,N_37049);
and U39459 (N_39459,N_37038,N_36431);
and U39460 (N_39460,N_36019,N_37066);
or U39461 (N_39461,N_37197,N_36976);
or U39462 (N_39462,N_37865,N_36113);
nor U39463 (N_39463,N_37461,N_37640);
and U39464 (N_39464,N_36308,N_37047);
xnor U39465 (N_39465,N_36048,N_36416);
xor U39466 (N_39466,N_36762,N_36412);
nand U39467 (N_39467,N_36235,N_37805);
nand U39468 (N_39468,N_36589,N_36175);
nor U39469 (N_39469,N_37631,N_37773);
nand U39470 (N_39470,N_36291,N_37304);
xnor U39471 (N_39471,N_37479,N_37553);
and U39472 (N_39472,N_36116,N_37933);
nand U39473 (N_39473,N_36490,N_37783);
nor U39474 (N_39474,N_36225,N_36395);
nor U39475 (N_39475,N_37816,N_36555);
nor U39476 (N_39476,N_37937,N_36373);
nor U39477 (N_39477,N_36004,N_36098);
and U39478 (N_39478,N_36019,N_37934);
xnor U39479 (N_39479,N_37041,N_36618);
nor U39480 (N_39480,N_36310,N_37074);
xnor U39481 (N_39481,N_37198,N_36572);
xor U39482 (N_39482,N_36108,N_36026);
xor U39483 (N_39483,N_37366,N_37474);
nor U39484 (N_39484,N_36771,N_37716);
or U39485 (N_39485,N_37973,N_37146);
and U39486 (N_39486,N_36179,N_37109);
and U39487 (N_39487,N_37062,N_36947);
or U39488 (N_39488,N_36417,N_36846);
or U39489 (N_39489,N_37385,N_36573);
nor U39490 (N_39490,N_36769,N_36125);
nor U39491 (N_39491,N_36431,N_37218);
and U39492 (N_39492,N_36224,N_36644);
xnor U39493 (N_39493,N_37908,N_36546);
nand U39494 (N_39494,N_37019,N_37723);
or U39495 (N_39495,N_37383,N_37022);
or U39496 (N_39496,N_37151,N_36175);
xor U39497 (N_39497,N_36523,N_37193);
xor U39498 (N_39498,N_37306,N_36293);
nand U39499 (N_39499,N_36158,N_37096);
and U39500 (N_39500,N_37588,N_36103);
and U39501 (N_39501,N_37863,N_36608);
nand U39502 (N_39502,N_37841,N_37568);
or U39503 (N_39503,N_36409,N_37837);
and U39504 (N_39504,N_37376,N_36954);
nand U39505 (N_39505,N_37998,N_36628);
nor U39506 (N_39506,N_37211,N_36561);
xor U39507 (N_39507,N_37348,N_37347);
and U39508 (N_39508,N_37177,N_37244);
nor U39509 (N_39509,N_37991,N_37663);
or U39510 (N_39510,N_37429,N_37515);
and U39511 (N_39511,N_37970,N_36760);
and U39512 (N_39512,N_37136,N_36435);
nor U39513 (N_39513,N_37287,N_36730);
xor U39514 (N_39514,N_37970,N_36829);
nand U39515 (N_39515,N_36473,N_37902);
nor U39516 (N_39516,N_37054,N_37692);
and U39517 (N_39517,N_36756,N_37755);
xor U39518 (N_39518,N_36842,N_36217);
xnor U39519 (N_39519,N_37966,N_37520);
nor U39520 (N_39520,N_36242,N_36251);
nand U39521 (N_39521,N_37340,N_36354);
nor U39522 (N_39522,N_37540,N_37292);
xor U39523 (N_39523,N_36477,N_37199);
or U39524 (N_39524,N_37337,N_37776);
nor U39525 (N_39525,N_36680,N_36505);
nor U39526 (N_39526,N_36835,N_37827);
or U39527 (N_39527,N_37729,N_37409);
and U39528 (N_39528,N_37420,N_36217);
and U39529 (N_39529,N_36068,N_36866);
xor U39530 (N_39530,N_37635,N_37824);
xor U39531 (N_39531,N_37544,N_37866);
nand U39532 (N_39532,N_37643,N_36455);
nand U39533 (N_39533,N_36328,N_36795);
nand U39534 (N_39534,N_37435,N_36814);
nand U39535 (N_39535,N_36535,N_37772);
xnor U39536 (N_39536,N_36012,N_37056);
nand U39537 (N_39537,N_37020,N_36640);
and U39538 (N_39538,N_36805,N_37278);
xnor U39539 (N_39539,N_37229,N_37512);
xnor U39540 (N_39540,N_37877,N_36973);
xnor U39541 (N_39541,N_37779,N_37490);
nand U39542 (N_39542,N_36465,N_36043);
nor U39543 (N_39543,N_36721,N_36665);
nand U39544 (N_39544,N_37404,N_37289);
xnor U39545 (N_39545,N_36705,N_36999);
nor U39546 (N_39546,N_37534,N_36850);
nor U39547 (N_39547,N_37591,N_37939);
xnor U39548 (N_39548,N_36970,N_37584);
xnor U39549 (N_39549,N_36265,N_36060);
nor U39550 (N_39550,N_37054,N_36666);
and U39551 (N_39551,N_37138,N_37919);
nor U39552 (N_39552,N_36970,N_36661);
xor U39553 (N_39553,N_37428,N_37565);
nor U39554 (N_39554,N_37643,N_37853);
and U39555 (N_39555,N_36428,N_36265);
nor U39556 (N_39556,N_36375,N_37143);
or U39557 (N_39557,N_37500,N_36098);
or U39558 (N_39558,N_37716,N_37532);
nand U39559 (N_39559,N_37324,N_36842);
or U39560 (N_39560,N_36377,N_36604);
xnor U39561 (N_39561,N_37137,N_37952);
xnor U39562 (N_39562,N_37062,N_36738);
xnor U39563 (N_39563,N_37979,N_36607);
xnor U39564 (N_39564,N_36153,N_36511);
xnor U39565 (N_39565,N_37297,N_36499);
and U39566 (N_39566,N_37532,N_37198);
nand U39567 (N_39567,N_37288,N_37256);
or U39568 (N_39568,N_37098,N_36307);
nor U39569 (N_39569,N_37790,N_37267);
nor U39570 (N_39570,N_36035,N_37272);
and U39571 (N_39571,N_36767,N_37475);
or U39572 (N_39572,N_37721,N_36768);
nand U39573 (N_39573,N_36992,N_36419);
and U39574 (N_39574,N_36189,N_36117);
or U39575 (N_39575,N_36346,N_36564);
or U39576 (N_39576,N_37310,N_36987);
nand U39577 (N_39577,N_37990,N_37882);
xnor U39578 (N_39578,N_36405,N_36762);
nor U39579 (N_39579,N_37894,N_36630);
and U39580 (N_39580,N_37065,N_37151);
and U39581 (N_39581,N_37532,N_36285);
xor U39582 (N_39582,N_37577,N_36215);
nor U39583 (N_39583,N_36758,N_37130);
and U39584 (N_39584,N_37214,N_37148);
xor U39585 (N_39585,N_36530,N_37282);
xor U39586 (N_39586,N_37564,N_37085);
and U39587 (N_39587,N_36617,N_37013);
or U39588 (N_39588,N_37845,N_37551);
nand U39589 (N_39589,N_37690,N_37046);
xnor U39590 (N_39590,N_37795,N_36932);
and U39591 (N_39591,N_37688,N_37142);
nor U39592 (N_39592,N_37967,N_37787);
xor U39593 (N_39593,N_37327,N_36560);
and U39594 (N_39594,N_36860,N_36626);
nand U39595 (N_39595,N_36291,N_36733);
xor U39596 (N_39596,N_37995,N_37419);
nor U39597 (N_39597,N_37315,N_37691);
xor U39598 (N_39598,N_36595,N_37086);
or U39599 (N_39599,N_36466,N_37591);
nor U39600 (N_39600,N_37494,N_36883);
or U39601 (N_39601,N_36622,N_36634);
or U39602 (N_39602,N_37876,N_37960);
nand U39603 (N_39603,N_37082,N_37321);
or U39604 (N_39604,N_37016,N_37346);
or U39605 (N_39605,N_36417,N_37054);
nor U39606 (N_39606,N_36898,N_37860);
xor U39607 (N_39607,N_37306,N_37422);
or U39608 (N_39608,N_37464,N_36949);
and U39609 (N_39609,N_36196,N_36899);
nand U39610 (N_39610,N_36683,N_36248);
nor U39611 (N_39611,N_37388,N_36951);
or U39612 (N_39612,N_36559,N_36311);
nor U39613 (N_39613,N_37983,N_36899);
xor U39614 (N_39614,N_37210,N_36241);
nand U39615 (N_39615,N_37444,N_36394);
nand U39616 (N_39616,N_36703,N_37321);
nor U39617 (N_39617,N_37666,N_36856);
nand U39618 (N_39618,N_37881,N_36548);
nand U39619 (N_39619,N_37808,N_37916);
and U39620 (N_39620,N_37931,N_37711);
nor U39621 (N_39621,N_36600,N_36407);
xnor U39622 (N_39622,N_36307,N_37152);
and U39623 (N_39623,N_36498,N_37417);
xor U39624 (N_39624,N_36745,N_37474);
and U39625 (N_39625,N_36428,N_36090);
and U39626 (N_39626,N_37215,N_37101);
or U39627 (N_39627,N_37620,N_36312);
and U39628 (N_39628,N_36194,N_36778);
nand U39629 (N_39629,N_36516,N_36197);
xnor U39630 (N_39630,N_36614,N_37042);
nand U39631 (N_39631,N_36830,N_37613);
nand U39632 (N_39632,N_37471,N_37836);
nor U39633 (N_39633,N_37477,N_36379);
nand U39634 (N_39634,N_36470,N_36664);
nor U39635 (N_39635,N_36781,N_37115);
nor U39636 (N_39636,N_37840,N_36577);
nand U39637 (N_39637,N_37288,N_37477);
or U39638 (N_39638,N_36175,N_37022);
nor U39639 (N_39639,N_36242,N_37898);
xor U39640 (N_39640,N_37300,N_36128);
and U39641 (N_39641,N_36607,N_36088);
or U39642 (N_39642,N_36300,N_36655);
xor U39643 (N_39643,N_36284,N_36199);
xnor U39644 (N_39644,N_36830,N_37309);
nor U39645 (N_39645,N_36252,N_37892);
nor U39646 (N_39646,N_37425,N_37104);
xnor U39647 (N_39647,N_36054,N_36042);
and U39648 (N_39648,N_36657,N_36978);
nand U39649 (N_39649,N_37716,N_36824);
and U39650 (N_39650,N_36776,N_36114);
and U39651 (N_39651,N_37025,N_36291);
nand U39652 (N_39652,N_37838,N_36833);
or U39653 (N_39653,N_36483,N_37900);
or U39654 (N_39654,N_36155,N_36546);
or U39655 (N_39655,N_37891,N_36358);
xor U39656 (N_39656,N_37169,N_36018);
xnor U39657 (N_39657,N_36046,N_37254);
or U39658 (N_39658,N_37060,N_36576);
and U39659 (N_39659,N_36583,N_37003);
or U39660 (N_39660,N_36365,N_36095);
or U39661 (N_39661,N_37767,N_37915);
xor U39662 (N_39662,N_37028,N_36453);
or U39663 (N_39663,N_37926,N_36360);
or U39664 (N_39664,N_37256,N_37453);
nand U39665 (N_39665,N_36283,N_36459);
xor U39666 (N_39666,N_36764,N_37936);
or U39667 (N_39667,N_36154,N_37684);
nor U39668 (N_39668,N_36670,N_36493);
nor U39669 (N_39669,N_36623,N_36118);
or U39670 (N_39670,N_36281,N_37857);
nand U39671 (N_39671,N_36448,N_36562);
nand U39672 (N_39672,N_37111,N_36453);
xnor U39673 (N_39673,N_37252,N_36478);
xnor U39674 (N_39674,N_37602,N_36875);
nor U39675 (N_39675,N_36864,N_37417);
nor U39676 (N_39676,N_37581,N_36118);
or U39677 (N_39677,N_37820,N_36566);
nor U39678 (N_39678,N_36359,N_37004);
nand U39679 (N_39679,N_36746,N_36871);
nand U39680 (N_39680,N_37270,N_37843);
nand U39681 (N_39681,N_37466,N_37530);
and U39682 (N_39682,N_37250,N_37596);
or U39683 (N_39683,N_36801,N_37974);
nor U39684 (N_39684,N_36306,N_37725);
nand U39685 (N_39685,N_37982,N_37845);
xor U39686 (N_39686,N_37258,N_36394);
xor U39687 (N_39687,N_36628,N_36698);
nor U39688 (N_39688,N_37227,N_36560);
xnor U39689 (N_39689,N_37364,N_36142);
or U39690 (N_39690,N_37518,N_37402);
or U39691 (N_39691,N_36668,N_37859);
nor U39692 (N_39692,N_37568,N_37609);
xor U39693 (N_39693,N_37094,N_37820);
and U39694 (N_39694,N_37333,N_36244);
and U39695 (N_39695,N_37170,N_37051);
nor U39696 (N_39696,N_36036,N_36724);
xor U39697 (N_39697,N_37566,N_36491);
nor U39698 (N_39698,N_37510,N_37726);
and U39699 (N_39699,N_36166,N_37989);
and U39700 (N_39700,N_37091,N_36802);
xor U39701 (N_39701,N_37092,N_37849);
nor U39702 (N_39702,N_36537,N_36812);
or U39703 (N_39703,N_37137,N_37959);
or U39704 (N_39704,N_36147,N_36376);
xnor U39705 (N_39705,N_37998,N_37170);
xor U39706 (N_39706,N_36016,N_37382);
nor U39707 (N_39707,N_37350,N_37772);
xnor U39708 (N_39708,N_36917,N_37777);
and U39709 (N_39709,N_36885,N_36820);
and U39710 (N_39710,N_36449,N_36684);
nand U39711 (N_39711,N_37245,N_36464);
and U39712 (N_39712,N_36976,N_37811);
nor U39713 (N_39713,N_37072,N_37678);
and U39714 (N_39714,N_36181,N_36168);
and U39715 (N_39715,N_37750,N_36609);
and U39716 (N_39716,N_37721,N_36571);
nand U39717 (N_39717,N_36326,N_37837);
and U39718 (N_39718,N_37257,N_37054);
xnor U39719 (N_39719,N_36214,N_36180);
and U39720 (N_39720,N_36027,N_37698);
xor U39721 (N_39721,N_37126,N_36895);
and U39722 (N_39722,N_36153,N_37120);
or U39723 (N_39723,N_36434,N_37185);
or U39724 (N_39724,N_36571,N_36535);
xor U39725 (N_39725,N_37209,N_36898);
nor U39726 (N_39726,N_37249,N_37221);
nand U39727 (N_39727,N_36189,N_36642);
or U39728 (N_39728,N_37164,N_36320);
nor U39729 (N_39729,N_37667,N_36744);
xnor U39730 (N_39730,N_37090,N_36588);
xnor U39731 (N_39731,N_37965,N_37894);
and U39732 (N_39732,N_37723,N_36018);
nand U39733 (N_39733,N_37631,N_37630);
and U39734 (N_39734,N_37967,N_36466);
or U39735 (N_39735,N_36005,N_36063);
xor U39736 (N_39736,N_36105,N_36469);
nand U39737 (N_39737,N_37289,N_36055);
and U39738 (N_39738,N_36091,N_37311);
nand U39739 (N_39739,N_36107,N_37415);
nand U39740 (N_39740,N_36988,N_37176);
nand U39741 (N_39741,N_37038,N_37513);
or U39742 (N_39742,N_37757,N_37475);
xnor U39743 (N_39743,N_37516,N_36368);
nor U39744 (N_39744,N_37773,N_37449);
nor U39745 (N_39745,N_37957,N_37574);
xor U39746 (N_39746,N_36078,N_36747);
or U39747 (N_39747,N_37240,N_36270);
xnor U39748 (N_39748,N_36903,N_36653);
and U39749 (N_39749,N_37890,N_36579);
and U39750 (N_39750,N_36131,N_36298);
or U39751 (N_39751,N_37039,N_37527);
and U39752 (N_39752,N_37785,N_36501);
nor U39753 (N_39753,N_37928,N_37987);
or U39754 (N_39754,N_36907,N_37079);
or U39755 (N_39755,N_37015,N_37240);
nor U39756 (N_39756,N_36291,N_37532);
and U39757 (N_39757,N_37142,N_36807);
nand U39758 (N_39758,N_36484,N_37471);
nor U39759 (N_39759,N_36894,N_37029);
nor U39760 (N_39760,N_36205,N_37159);
or U39761 (N_39761,N_37023,N_36373);
and U39762 (N_39762,N_37853,N_37532);
nand U39763 (N_39763,N_37966,N_37762);
nor U39764 (N_39764,N_37166,N_37298);
nand U39765 (N_39765,N_37112,N_36475);
or U39766 (N_39766,N_36413,N_37375);
xnor U39767 (N_39767,N_37763,N_36524);
nand U39768 (N_39768,N_36818,N_36242);
xor U39769 (N_39769,N_37261,N_36817);
nor U39770 (N_39770,N_37548,N_37809);
and U39771 (N_39771,N_36799,N_36484);
or U39772 (N_39772,N_36555,N_36978);
nor U39773 (N_39773,N_36542,N_37908);
or U39774 (N_39774,N_37365,N_36418);
xnor U39775 (N_39775,N_37744,N_36718);
xor U39776 (N_39776,N_37866,N_37262);
nand U39777 (N_39777,N_36732,N_37813);
or U39778 (N_39778,N_36737,N_37701);
or U39779 (N_39779,N_37341,N_36466);
and U39780 (N_39780,N_37181,N_36822);
or U39781 (N_39781,N_37078,N_36027);
nor U39782 (N_39782,N_37001,N_37087);
nor U39783 (N_39783,N_36465,N_37771);
xor U39784 (N_39784,N_36110,N_37392);
and U39785 (N_39785,N_36111,N_36296);
xnor U39786 (N_39786,N_36027,N_37154);
or U39787 (N_39787,N_36340,N_36612);
and U39788 (N_39788,N_37269,N_37264);
nand U39789 (N_39789,N_36327,N_36554);
xnor U39790 (N_39790,N_36125,N_36961);
xnor U39791 (N_39791,N_36713,N_36034);
or U39792 (N_39792,N_36255,N_37536);
xnor U39793 (N_39793,N_37765,N_36796);
and U39794 (N_39794,N_36674,N_37863);
xor U39795 (N_39795,N_36909,N_36711);
nor U39796 (N_39796,N_36647,N_36010);
nor U39797 (N_39797,N_37079,N_36645);
or U39798 (N_39798,N_36435,N_36366);
xnor U39799 (N_39799,N_37280,N_36255);
and U39800 (N_39800,N_37686,N_36702);
and U39801 (N_39801,N_36755,N_36399);
xor U39802 (N_39802,N_37517,N_37377);
or U39803 (N_39803,N_36743,N_36329);
or U39804 (N_39804,N_36942,N_36251);
xnor U39805 (N_39805,N_36399,N_36566);
nor U39806 (N_39806,N_36970,N_37164);
nand U39807 (N_39807,N_37149,N_37716);
xor U39808 (N_39808,N_36075,N_37220);
or U39809 (N_39809,N_36583,N_36615);
or U39810 (N_39810,N_37284,N_36743);
nor U39811 (N_39811,N_36304,N_36928);
and U39812 (N_39812,N_37161,N_36768);
xnor U39813 (N_39813,N_37111,N_36354);
and U39814 (N_39814,N_36376,N_37687);
xnor U39815 (N_39815,N_37031,N_37016);
xnor U39816 (N_39816,N_37095,N_36066);
nand U39817 (N_39817,N_36352,N_36387);
and U39818 (N_39818,N_36446,N_36160);
nand U39819 (N_39819,N_37419,N_37591);
or U39820 (N_39820,N_37225,N_37991);
nand U39821 (N_39821,N_36765,N_37154);
nor U39822 (N_39822,N_37620,N_36122);
nor U39823 (N_39823,N_36027,N_36804);
nor U39824 (N_39824,N_37758,N_37429);
and U39825 (N_39825,N_37470,N_36582);
and U39826 (N_39826,N_36866,N_36300);
nand U39827 (N_39827,N_37541,N_37359);
nor U39828 (N_39828,N_37586,N_36728);
and U39829 (N_39829,N_37540,N_36319);
xnor U39830 (N_39830,N_37536,N_37560);
nand U39831 (N_39831,N_37647,N_37222);
or U39832 (N_39832,N_36743,N_36612);
nand U39833 (N_39833,N_36529,N_36289);
nand U39834 (N_39834,N_36086,N_36118);
or U39835 (N_39835,N_36308,N_36801);
nor U39836 (N_39836,N_37608,N_37277);
nand U39837 (N_39837,N_36761,N_36112);
or U39838 (N_39838,N_37840,N_37805);
xor U39839 (N_39839,N_36003,N_36891);
and U39840 (N_39840,N_37475,N_36101);
and U39841 (N_39841,N_36117,N_36830);
nor U39842 (N_39842,N_37029,N_37919);
and U39843 (N_39843,N_37407,N_37717);
nand U39844 (N_39844,N_36628,N_36433);
or U39845 (N_39845,N_37701,N_36339);
nand U39846 (N_39846,N_37306,N_37831);
and U39847 (N_39847,N_36071,N_36533);
nor U39848 (N_39848,N_37980,N_36418);
and U39849 (N_39849,N_37503,N_37698);
or U39850 (N_39850,N_36035,N_37437);
and U39851 (N_39851,N_37790,N_37778);
or U39852 (N_39852,N_36577,N_36858);
and U39853 (N_39853,N_36162,N_36388);
or U39854 (N_39854,N_37265,N_37428);
or U39855 (N_39855,N_36756,N_36736);
or U39856 (N_39856,N_36811,N_37025);
xor U39857 (N_39857,N_36248,N_36729);
xnor U39858 (N_39858,N_36574,N_36697);
nand U39859 (N_39859,N_36584,N_36639);
and U39860 (N_39860,N_36281,N_36611);
nor U39861 (N_39861,N_36736,N_36587);
or U39862 (N_39862,N_37565,N_37586);
nand U39863 (N_39863,N_37194,N_37571);
or U39864 (N_39864,N_36235,N_37346);
or U39865 (N_39865,N_36861,N_37564);
xnor U39866 (N_39866,N_37642,N_37771);
xor U39867 (N_39867,N_36602,N_37689);
nand U39868 (N_39868,N_36670,N_37002);
or U39869 (N_39869,N_36275,N_36925);
nor U39870 (N_39870,N_36534,N_37860);
xor U39871 (N_39871,N_36814,N_37724);
nand U39872 (N_39872,N_37875,N_36827);
and U39873 (N_39873,N_36742,N_36629);
or U39874 (N_39874,N_37210,N_37353);
or U39875 (N_39875,N_37607,N_36029);
nor U39876 (N_39876,N_36691,N_37508);
xor U39877 (N_39877,N_36992,N_36246);
and U39878 (N_39878,N_36510,N_36958);
and U39879 (N_39879,N_36389,N_36475);
nor U39880 (N_39880,N_36204,N_36948);
or U39881 (N_39881,N_36553,N_37898);
or U39882 (N_39882,N_37081,N_36136);
or U39883 (N_39883,N_37753,N_36146);
nand U39884 (N_39884,N_36775,N_37864);
nor U39885 (N_39885,N_37586,N_37133);
and U39886 (N_39886,N_36364,N_37076);
and U39887 (N_39887,N_36687,N_36900);
nor U39888 (N_39888,N_36744,N_36691);
nand U39889 (N_39889,N_37222,N_36124);
and U39890 (N_39890,N_37387,N_36257);
xnor U39891 (N_39891,N_37306,N_37886);
or U39892 (N_39892,N_36903,N_37004);
or U39893 (N_39893,N_36633,N_36101);
nand U39894 (N_39894,N_36064,N_37428);
or U39895 (N_39895,N_36953,N_37599);
xor U39896 (N_39896,N_37857,N_37888);
or U39897 (N_39897,N_37658,N_37434);
and U39898 (N_39898,N_36696,N_36324);
xor U39899 (N_39899,N_37147,N_37488);
and U39900 (N_39900,N_37461,N_36688);
nand U39901 (N_39901,N_37215,N_36754);
nand U39902 (N_39902,N_37190,N_37545);
xnor U39903 (N_39903,N_36277,N_36769);
or U39904 (N_39904,N_36296,N_36999);
xor U39905 (N_39905,N_37493,N_36094);
nor U39906 (N_39906,N_37871,N_37703);
nor U39907 (N_39907,N_36799,N_36329);
or U39908 (N_39908,N_36562,N_37511);
nor U39909 (N_39909,N_37213,N_36821);
nor U39910 (N_39910,N_36081,N_37530);
or U39911 (N_39911,N_36348,N_37283);
xnor U39912 (N_39912,N_37901,N_37254);
or U39913 (N_39913,N_36559,N_37380);
xnor U39914 (N_39914,N_37699,N_37896);
nand U39915 (N_39915,N_36732,N_37774);
or U39916 (N_39916,N_37029,N_37778);
or U39917 (N_39917,N_37416,N_36603);
or U39918 (N_39918,N_37142,N_36762);
nand U39919 (N_39919,N_36965,N_37877);
nor U39920 (N_39920,N_36459,N_36506);
nor U39921 (N_39921,N_37142,N_36144);
or U39922 (N_39922,N_36946,N_36159);
or U39923 (N_39923,N_37188,N_37774);
nand U39924 (N_39924,N_37188,N_37351);
xnor U39925 (N_39925,N_37229,N_36727);
nand U39926 (N_39926,N_37825,N_37134);
or U39927 (N_39927,N_37653,N_37847);
and U39928 (N_39928,N_37183,N_37013);
or U39929 (N_39929,N_37707,N_36633);
or U39930 (N_39930,N_36007,N_37702);
xnor U39931 (N_39931,N_36279,N_36449);
or U39932 (N_39932,N_37813,N_37447);
and U39933 (N_39933,N_36300,N_36096);
nor U39934 (N_39934,N_37941,N_36567);
nor U39935 (N_39935,N_37185,N_36258);
nor U39936 (N_39936,N_37639,N_36616);
nor U39937 (N_39937,N_37544,N_36095);
nor U39938 (N_39938,N_37385,N_36074);
nand U39939 (N_39939,N_37838,N_36425);
nor U39940 (N_39940,N_36170,N_36469);
nor U39941 (N_39941,N_36605,N_37722);
and U39942 (N_39942,N_36875,N_36047);
or U39943 (N_39943,N_36733,N_37762);
and U39944 (N_39944,N_37337,N_36367);
or U39945 (N_39945,N_36688,N_36489);
and U39946 (N_39946,N_36489,N_37745);
nor U39947 (N_39947,N_37526,N_36692);
or U39948 (N_39948,N_36785,N_36289);
xor U39949 (N_39949,N_36949,N_36463);
nand U39950 (N_39950,N_36210,N_36783);
or U39951 (N_39951,N_37235,N_36664);
or U39952 (N_39952,N_37969,N_37485);
and U39953 (N_39953,N_36556,N_37332);
or U39954 (N_39954,N_36476,N_37181);
nor U39955 (N_39955,N_37498,N_37613);
and U39956 (N_39956,N_36533,N_36390);
xor U39957 (N_39957,N_36982,N_37120);
and U39958 (N_39958,N_37178,N_37159);
or U39959 (N_39959,N_36961,N_36499);
xor U39960 (N_39960,N_37144,N_36697);
nor U39961 (N_39961,N_36756,N_36043);
or U39962 (N_39962,N_37659,N_37824);
nor U39963 (N_39963,N_36819,N_36252);
xor U39964 (N_39964,N_37451,N_36700);
xor U39965 (N_39965,N_36520,N_36515);
nand U39966 (N_39966,N_36608,N_36415);
nor U39967 (N_39967,N_36754,N_37702);
xnor U39968 (N_39968,N_36096,N_37659);
and U39969 (N_39969,N_37031,N_36849);
nor U39970 (N_39970,N_37857,N_36915);
nor U39971 (N_39971,N_36780,N_36328);
and U39972 (N_39972,N_37293,N_37459);
and U39973 (N_39973,N_37205,N_37775);
or U39974 (N_39974,N_36495,N_37742);
and U39975 (N_39975,N_37242,N_36778);
nand U39976 (N_39976,N_36833,N_37756);
nand U39977 (N_39977,N_37416,N_37216);
nand U39978 (N_39978,N_36278,N_37760);
nor U39979 (N_39979,N_36385,N_36225);
or U39980 (N_39980,N_37300,N_36901);
nor U39981 (N_39981,N_37176,N_37335);
nor U39982 (N_39982,N_37483,N_36231);
and U39983 (N_39983,N_37631,N_36530);
and U39984 (N_39984,N_36452,N_37843);
xnor U39985 (N_39985,N_36140,N_37736);
or U39986 (N_39986,N_37414,N_36425);
nor U39987 (N_39987,N_37000,N_36294);
or U39988 (N_39988,N_37810,N_37265);
nand U39989 (N_39989,N_36705,N_36116);
or U39990 (N_39990,N_37659,N_36769);
xor U39991 (N_39991,N_36422,N_36832);
nor U39992 (N_39992,N_37308,N_37103);
and U39993 (N_39993,N_37354,N_37348);
and U39994 (N_39994,N_37456,N_36099);
xor U39995 (N_39995,N_36969,N_36402);
nor U39996 (N_39996,N_36358,N_36763);
or U39997 (N_39997,N_37232,N_37973);
nand U39998 (N_39998,N_36984,N_37589);
nand U39999 (N_39999,N_36139,N_36256);
and U40000 (N_40000,N_39340,N_38134);
nor U40001 (N_40001,N_39658,N_39174);
or U40002 (N_40002,N_39436,N_38831);
or U40003 (N_40003,N_39718,N_38342);
nor U40004 (N_40004,N_39118,N_39938);
nand U40005 (N_40005,N_39389,N_39593);
and U40006 (N_40006,N_39988,N_38926);
nor U40007 (N_40007,N_38072,N_39797);
or U40008 (N_40008,N_39401,N_39335);
or U40009 (N_40009,N_39303,N_39461);
and U40010 (N_40010,N_38776,N_38992);
xnor U40011 (N_40011,N_39835,N_39367);
nand U40012 (N_40012,N_38521,N_39199);
nand U40013 (N_40013,N_39032,N_39384);
nor U40014 (N_40014,N_38848,N_38091);
nand U40015 (N_40015,N_39509,N_39779);
or U40016 (N_40016,N_38287,N_38759);
or U40017 (N_40017,N_38253,N_38105);
and U40018 (N_40018,N_39641,N_38034);
or U40019 (N_40019,N_39715,N_38353);
nor U40020 (N_40020,N_38839,N_38191);
nand U40021 (N_40021,N_38911,N_38099);
nor U40022 (N_40022,N_38995,N_39404);
and U40023 (N_40023,N_39852,N_39838);
nor U40024 (N_40024,N_39589,N_38966);
nor U40025 (N_40025,N_39728,N_39172);
nor U40026 (N_40026,N_39189,N_38943);
xnor U40027 (N_40027,N_38504,N_39685);
or U40028 (N_40028,N_38798,N_38586);
and U40029 (N_40029,N_38960,N_38818);
or U40030 (N_40030,N_38567,N_39037);
xor U40031 (N_40031,N_39081,N_39661);
nand U40032 (N_40032,N_38994,N_38860);
and U40033 (N_40033,N_39135,N_38052);
xnor U40034 (N_40034,N_38165,N_39517);
xor U40035 (N_40035,N_39977,N_39616);
nand U40036 (N_40036,N_38632,N_38406);
nand U40037 (N_40037,N_38724,N_39433);
and U40038 (N_40038,N_39333,N_39855);
or U40039 (N_40039,N_38872,N_38178);
xor U40040 (N_40040,N_39448,N_39612);
nor U40041 (N_40041,N_39360,N_39343);
xnor U40042 (N_40042,N_39020,N_38520);
nand U40043 (N_40043,N_39765,N_39870);
nor U40044 (N_40044,N_38955,N_39746);
xnor U40045 (N_40045,N_38298,N_39643);
xnor U40046 (N_40046,N_38918,N_39444);
nand U40047 (N_40047,N_38453,N_39426);
or U40048 (N_40048,N_39435,N_38999);
xor U40049 (N_40049,N_39165,N_38501);
and U40050 (N_40050,N_38833,N_39899);
or U40051 (N_40051,N_39709,N_38998);
nor U40052 (N_40052,N_38325,N_39656);
or U40053 (N_40053,N_38046,N_39609);
nor U40054 (N_40054,N_38115,N_39791);
nand U40055 (N_40055,N_38448,N_38183);
nand U40056 (N_40056,N_39341,N_39566);
xor U40057 (N_40057,N_38132,N_38804);
xor U40058 (N_40058,N_38543,N_38514);
nor U40059 (N_40059,N_38161,N_39066);
xor U40060 (N_40060,N_38479,N_39753);
and U40061 (N_40061,N_38174,N_39901);
nand U40062 (N_40062,N_39153,N_38013);
or U40063 (N_40063,N_38440,N_39088);
and U40064 (N_40064,N_39913,N_39140);
nand U40065 (N_40065,N_38476,N_39083);
or U40066 (N_40066,N_39922,N_38513);
nor U40067 (N_40067,N_39447,N_38620);
or U40068 (N_40068,N_38944,N_39871);
or U40069 (N_40069,N_39608,N_39904);
and U40070 (N_40070,N_39575,N_39001);
or U40071 (N_40071,N_38541,N_39991);
nor U40072 (N_40072,N_38332,N_38748);
xor U40073 (N_40073,N_39339,N_38761);
nand U40074 (N_40074,N_38016,N_39815);
nand U40075 (N_40075,N_39613,N_39460);
nand U40076 (N_40076,N_39758,N_39085);
xnor U40077 (N_40077,N_38750,N_38713);
nand U40078 (N_40078,N_38899,N_39308);
and U40079 (N_40079,N_38626,N_39722);
nand U40080 (N_40080,N_38411,N_39209);
or U40081 (N_40081,N_39620,N_39796);
nor U40082 (N_40082,N_38009,N_38117);
nand U40083 (N_40083,N_39252,N_38442);
xnor U40084 (N_40084,N_39601,N_38840);
nand U40085 (N_40085,N_39158,N_39406);
and U40086 (N_40086,N_39025,N_38335);
nor U40087 (N_40087,N_38649,N_38341);
and U40088 (N_40088,N_38255,N_38515);
or U40089 (N_40089,N_38116,N_39091);
and U40090 (N_40090,N_39498,N_38517);
and U40091 (N_40091,N_39466,N_38392);
nand U40092 (N_40092,N_38668,N_39468);
or U40093 (N_40093,N_38801,N_39271);
nand U40094 (N_40094,N_38763,N_38607);
and U40095 (N_40095,N_39992,N_38712);
xor U40096 (N_40096,N_38153,N_38524);
nor U40097 (N_40097,N_39955,N_38928);
or U40098 (N_40098,N_39840,N_39306);
xor U40099 (N_40099,N_39663,N_38493);
and U40100 (N_40100,N_39314,N_38130);
nor U40101 (N_40101,N_39800,N_39947);
and U40102 (N_40102,N_38989,N_38721);
nand U40103 (N_40103,N_38551,N_39615);
and U40104 (N_40104,N_39634,N_39078);
xnor U40105 (N_40105,N_38273,N_39205);
nand U40106 (N_40106,N_39607,N_38963);
nand U40107 (N_40107,N_38283,N_38006);
and U40108 (N_40108,N_38187,N_38980);
xor U40109 (N_40109,N_39095,N_38876);
nor U40110 (N_40110,N_38741,N_39286);
and U40111 (N_40111,N_38317,N_39524);
or U40112 (N_40112,N_38048,N_39945);
nor U40113 (N_40113,N_39154,N_38002);
nand U40114 (N_40114,N_38791,N_39263);
nor U40115 (N_40115,N_39261,N_39320);
and U40116 (N_40116,N_39833,N_38704);
nor U40117 (N_40117,N_38157,N_38619);
nor U40118 (N_40118,N_39757,N_39281);
and U40119 (N_40119,N_38962,N_39850);
nand U40120 (N_40120,N_39808,N_38398);
nor U40121 (N_40121,N_39238,N_38077);
and U40122 (N_40122,N_39255,N_39481);
and U40123 (N_40123,N_39843,N_38289);
and U40124 (N_40124,N_39486,N_38576);
or U40125 (N_40125,N_38901,N_39542);
and U40126 (N_40126,N_39701,N_39812);
xor U40127 (N_40127,N_39492,N_38202);
or U40128 (N_40128,N_38836,N_39953);
nand U40129 (N_40129,N_38420,N_39573);
or U40130 (N_40130,N_38486,N_39549);
nand U40131 (N_40131,N_38393,N_38527);
nor U40132 (N_40132,N_39457,N_38718);
nand U40133 (N_40133,N_39366,N_38078);
xnor U40134 (N_40134,N_38060,N_38413);
nor U40135 (N_40135,N_39532,N_39914);
and U40136 (N_40136,N_39847,N_39372);
nor U40137 (N_40137,N_39786,N_38868);
xnor U40138 (N_40138,N_38376,N_39398);
xnor U40139 (N_40139,N_38772,N_39592);
and U40140 (N_40140,N_39379,N_39386);
xnor U40141 (N_40141,N_39163,N_39275);
nor U40142 (N_40142,N_39240,N_39645);
and U40143 (N_40143,N_39980,N_39957);
and U40144 (N_40144,N_39694,N_38326);
nor U40145 (N_40145,N_38577,N_39396);
xnor U40146 (N_40146,N_38700,N_38644);
nand U40147 (N_40147,N_38354,N_39302);
nor U40148 (N_40148,N_38595,N_39693);
and U40149 (N_40149,N_38321,N_38940);
and U40150 (N_40150,N_39635,N_39142);
and U40151 (N_40151,N_39007,N_39581);
xnor U40152 (N_40152,N_39124,N_39235);
nand U40153 (N_40153,N_39941,N_38399);
nor U40154 (N_40154,N_38710,N_38604);
nand U40155 (N_40155,N_39846,N_38093);
or U40156 (N_40156,N_38278,N_38234);
or U40157 (N_40157,N_38225,N_39056);
or U40158 (N_40158,N_38871,N_38020);
nor U40159 (N_40159,N_39310,N_39782);
nand U40160 (N_40160,N_39723,N_39221);
nand U40161 (N_40161,N_39096,N_39951);
nor U40162 (N_40162,N_39917,N_38591);
nand U40163 (N_40163,N_39546,N_38931);
xnor U40164 (N_40164,N_39826,N_39767);
and U40165 (N_40165,N_38065,N_38059);
and U40166 (N_40166,N_38461,N_39052);
or U40167 (N_40167,N_39650,N_38687);
nand U40168 (N_40168,N_38869,N_38032);
nor U40169 (N_40169,N_39336,N_39241);
or U40170 (N_40170,N_38482,N_38507);
nor U40171 (N_40171,N_39283,N_39337);
or U40172 (N_40172,N_38137,N_38478);
nor U40173 (N_40173,N_38382,N_38436);
or U40174 (N_40174,N_38435,N_39187);
or U40175 (N_40175,N_38570,N_39582);
xor U40176 (N_40176,N_38374,N_38328);
and U40177 (N_40177,N_39887,N_38303);
xor U40178 (N_40178,N_39895,N_38754);
nand U40179 (N_40179,N_38867,N_39894);
xnor U40180 (N_40180,N_38813,N_38574);
xnor U40181 (N_40181,N_38343,N_38533);
nor U40182 (N_40182,N_38673,N_39692);
nand U40183 (N_40183,N_38601,N_39752);
or U40184 (N_40184,N_38133,N_38734);
or U40185 (N_40185,N_39878,N_38177);
nor U40186 (N_40186,N_38686,N_39113);
or U40187 (N_40187,N_39060,N_38952);
nor U40188 (N_40188,N_39505,N_38490);
nor U40189 (N_40189,N_38864,N_38910);
nand U40190 (N_40190,N_39246,N_39157);
nor U40191 (N_40191,N_39045,N_38347);
or U40192 (N_40192,N_39217,N_39961);
or U40193 (N_40193,N_38351,N_39857);
and U40194 (N_40194,N_38651,N_38349);
and U40195 (N_40195,N_39536,N_38879);
and U40196 (N_40196,N_38689,N_38635);
or U40197 (N_40197,N_38770,N_39934);
and U40198 (N_40198,N_39868,N_39872);
and U40199 (N_40199,N_39256,N_39079);
or U40200 (N_40200,N_38360,N_39130);
and U40201 (N_40201,N_39028,N_39185);
or U40202 (N_40202,N_39167,N_38402);
nand U40203 (N_40203,N_39368,N_38642);
nand U40204 (N_40204,N_39430,N_38881);
and U40205 (N_40205,N_38258,N_38290);
or U40206 (N_40206,N_39743,N_39983);
or U40207 (N_40207,N_39484,N_38694);
nor U40208 (N_40208,N_39465,N_38544);
xnor U40209 (N_40209,N_38025,N_38978);
or U40210 (N_40210,N_38053,N_39734);
xor U40211 (N_40211,N_38859,N_39363);
nand U40212 (N_40212,N_39540,N_39984);
nand U40213 (N_40213,N_39301,N_38502);
or U40214 (N_40214,N_38780,N_38891);
xnor U40215 (N_40215,N_38387,N_38481);
nor U40216 (N_40216,N_39383,N_38222);
nor U40217 (N_40217,N_38268,N_38766);
nor U40218 (N_40218,N_38208,N_39048);
xor U40219 (N_40219,N_39668,N_39086);
xnor U40220 (N_40220,N_38193,N_38449);
or U40221 (N_40221,N_39018,N_38646);
nor U40222 (N_40222,N_39664,N_38975);
xnor U40223 (N_40223,N_38143,N_39968);
xor U40224 (N_40224,N_39770,N_39330);
or U40225 (N_40225,N_39538,N_38716);
nor U40226 (N_40226,N_38030,N_38681);
xor U40227 (N_40227,N_38226,N_38622);
xor U40228 (N_40228,N_39175,N_38429);
xnor U40229 (N_40229,N_39952,N_39541);
or U40230 (N_40230,N_38498,N_38707);
and U40231 (N_40231,N_39925,N_38275);
and U40232 (N_40232,N_38196,N_39138);
xor U40233 (N_40233,N_38739,N_39422);
nand U40234 (N_40234,N_38499,N_39215);
nor U40235 (N_40235,N_38372,N_38516);
or U40236 (N_40236,N_38634,N_38898);
and U40237 (N_40237,N_38631,N_38170);
or U40238 (N_40238,N_39188,N_38896);
or U40239 (N_40239,N_39585,N_39982);
xnor U40240 (N_40240,N_38924,N_38799);
or U40241 (N_40241,N_39376,N_38331);
xor U40242 (N_40242,N_38835,N_39706);
nand U40243 (N_40243,N_38333,N_39662);
or U40244 (N_40244,N_39967,N_38200);
or U40245 (N_40245,N_38519,N_39322);
nor U40246 (N_40246,N_38271,N_39935);
xor U40247 (N_40247,N_38259,N_39229);
nand U40248 (N_40248,N_38982,N_39013);
nand U40249 (N_40249,N_39417,N_39733);
xnor U40250 (N_40250,N_38756,N_39773);
or U40251 (N_40251,N_39489,N_38042);
nand U40252 (N_40252,N_39618,N_39251);
nand U40253 (N_40253,N_38054,N_39137);
and U40254 (N_40254,N_38542,N_38854);
or U40255 (N_40255,N_38862,N_38787);
xnor U40256 (N_40256,N_39795,N_39245);
xor U40257 (N_40257,N_38785,N_39766);
nor U40258 (N_40258,N_38659,N_39463);
xor U40259 (N_40259,N_38929,N_38480);
nand U40260 (N_40260,N_38796,N_39660);
nor U40261 (N_40261,N_39802,N_38579);
nand U40262 (N_40262,N_38532,N_39429);
and U40263 (N_40263,N_38452,N_38865);
xnor U40264 (N_40264,N_39327,N_39555);
nand U40265 (N_40265,N_39006,N_39160);
or U40266 (N_40266,N_39792,N_39544);
xnor U40267 (N_40267,N_38397,N_38883);
xnor U40268 (N_40268,N_38845,N_39563);
or U40269 (N_40269,N_39510,N_38746);
and U40270 (N_40270,N_39731,N_39208);
nand U40271 (N_40271,N_38367,N_38221);
nor U40272 (N_40272,N_39801,N_38385);
nand U40273 (N_40273,N_39464,N_39885);
xor U40274 (N_40274,N_39110,N_39491);
nor U40275 (N_40275,N_38555,N_39749);
nor U40276 (N_40276,N_39506,N_39487);
nand U40277 (N_40277,N_38007,N_39450);
and U40278 (N_40278,N_39195,N_39811);
xor U40279 (N_40279,N_38286,N_38458);
and U40280 (N_40280,N_38008,N_39114);
nor U40281 (N_40281,N_38483,N_38970);
and U40282 (N_40282,N_39845,N_38923);
nor U40283 (N_40283,N_39479,N_39459);
nor U40284 (N_40284,N_39619,N_38892);
nor U40285 (N_40285,N_38122,N_38578);
nand U40286 (N_40286,N_38152,N_38214);
or U40287 (N_40287,N_38597,N_39316);
xnor U40288 (N_40288,N_39649,N_39416);
xor U40289 (N_40289,N_39102,N_39219);
or U40290 (N_40290,N_39184,N_38070);
or U40291 (N_40291,N_39046,N_38968);
or U40292 (N_40292,N_38320,N_38834);
nor U40293 (N_40293,N_38523,N_39453);
xnor U40294 (N_40294,N_39321,N_38653);
or U40295 (N_40295,N_39891,N_39994);
or U40296 (N_40296,N_38997,N_38223);
and U40297 (N_40297,N_39446,N_38582);
nor U40298 (N_40298,N_38991,N_38274);
xnor U40299 (N_40299,N_38920,N_38293);
xnor U40300 (N_40300,N_38670,N_38497);
and U40301 (N_40301,N_38095,N_39213);
and U40302 (N_40302,N_39823,N_39710);
and U40303 (N_40303,N_38186,N_38264);
nor U40304 (N_40304,N_39974,N_38184);
nand U40305 (N_40305,N_39674,N_39061);
nand U40306 (N_40306,N_38658,N_39837);
nand U40307 (N_40307,N_39965,N_38121);
and U40308 (N_40308,N_38907,N_39120);
nor U40309 (N_40309,N_39307,N_38028);
or U40310 (N_40310,N_38055,N_39351);
or U40311 (N_40311,N_38814,N_38365);
nand U40312 (N_40312,N_39586,N_39033);
or U40313 (N_40313,N_38897,N_38003);
nand U40314 (N_40314,N_38702,N_39519);
nand U40315 (N_40315,N_39841,N_38381);
and U40316 (N_40316,N_39182,N_39880);
nand U40317 (N_40317,N_38654,N_39741);
nor U40318 (N_40318,N_38618,N_39525);
and U40319 (N_40319,N_39583,N_39101);
nand U40320 (N_40320,N_38204,N_38949);
xnor U40321 (N_40321,N_39671,N_39739);
nand U40322 (N_40322,N_39365,N_39295);
nand U40323 (N_40323,N_39866,N_39909);
nand U40324 (N_40324,N_39171,N_39625);
nor U40325 (N_40325,N_38890,N_39075);
and U40326 (N_40326,N_39642,N_38842);
nor U40327 (N_40327,N_38518,N_38408);
xnor U40328 (N_40328,N_39599,N_38806);
nor U40329 (N_40329,N_38637,N_38339);
and U40330 (N_40330,N_38786,N_39144);
or U40331 (N_40331,N_38154,N_39572);
nand U40332 (N_40332,N_38050,N_38069);
or U40333 (N_40333,N_38424,N_39640);
xnor U40334 (N_40334,N_38005,N_38605);
and U40335 (N_40335,N_38305,N_39777);
nand U40336 (N_40336,N_39997,N_38781);
nand U40337 (N_40337,N_39636,N_38693);
and U40338 (N_40338,N_38948,N_39035);
xnor U40339 (N_40339,N_38855,N_38951);
xor U40340 (N_40340,N_38248,N_38568);
or U40341 (N_40341,N_39548,N_39959);
nor U40342 (N_40342,N_39702,N_38464);
nor U40343 (N_40343,N_38128,N_39989);
and U40344 (N_40344,N_39305,N_38941);
nand U40345 (N_40345,N_38004,N_38740);
nand U40346 (N_40346,N_38236,N_38086);
nor U40347 (N_40347,N_39017,N_38846);
xor U40348 (N_40348,N_39304,N_38548);
and U40349 (N_40349,N_38987,N_38676);
xnor U40350 (N_40350,N_38388,N_38986);
nor U40351 (N_40351,N_38024,N_38348);
nand U40352 (N_40352,N_39788,N_38830);
and U40353 (N_40353,N_39131,N_38051);
and U40354 (N_40354,N_39454,N_38156);
and U40355 (N_40355,N_38324,N_38088);
nor U40356 (N_40356,N_38001,N_39287);
xnor U40357 (N_40357,N_39162,N_39699);
and U40358 (N_40358,N_39031,N_38616);
nand U40359 (N_40359,N_38337,N_38412);
or U40360 (N_40360,N_38329,N_38663);
nor U40361 (N_40361,N_39345,N_39467);
nor U40362 (N_40362,N_38664,N_39207);
nor U40363 (N_40363,N_39520,N_38703);
nand U40364 (N_40364,N_39041,N_38213);
nand U40365 (N_40365,N_38491,N_39318);
nor U40366 (N_40366,N_39818,N_38485);
nand U40367 (N_40367,N_39423,N_39108);
nor U40368 (N_40368,N_39996,N_38843);
xnor U40369 (N_40369,N_39611,N_38100);
xnor U40370 (N_40370,N_39192,N_39203);
xor U40371 (N_40371,N_39022,N_38742);
xnor U40372 (N_40372,N_39755,N_38506);
xnor U40373 (N_40373,N_39587,N_38185);
or U40374 (N_40374,N_39886,N_39312);
nand U40375 (N_40375,N_39276,N_38147);
nor U40376 (N_40376,N_39648,N_39150);
nor U40377 (N_40377,N_38407,N_38808);
and U40378 (N_40378,N_38035,N_38589);
or U40379 (N_40379,N_39356,N_38768);
or U40380 (N_40380,N_39862,N_39064);
nor U40381 (N_40381,N_38953,N_39839);
or U40382 (N_40382,N_39329,N_38254);
xor U40383 (N_40383,N_39844,N_39300);
or U40384 (N_40384,N_39169,N_39482);
nor U40385 (N_40385,N_39958,N_38379);
nor U40386 (N_40386,N_38231,N_39905);
or U40387 (N_40387,N_38224,N_38063);
xnor U40388 (N_40388,N_38580,N_38179);
or U40389 (N_40389,N_39206,N_39919);
and U40390 (N_40390,N_38957,N_38217);
nor U40391 (N_40391,N_39605,N_39652);
and U40392 (N_40392,N_38295,N_39698);
or U40393 (N_40393,N_39265,N_38014);
or U40394 (N_40394,N_39684,N_39093);
and U40395 (N_40395,N_39474,N_39512);
or U40396 (N_40396,N_39610,N_39347);
or U40397 (N_40397,N_38723,N_38391);
nand U40398 (N_40398,N_38935,N_38358);
nand U40399 (N_40399,N_38389,N_38084);
or U40400 (N_40400,N_38730,N_39145);
and U40401 (N_40401,N_38309,N_39393);
or U40402 (N_40402,N_38075,N_39883);
xor U40403 (N_40403,N_38067,N_39139);
xnor U40404 (N_40404,N_38299,N_38036);
nor U40405 (N_40405,N_39385,N_39125);
and U40406 (N_40406,N_39696,N_38585);
and U40407 (N_40407,N_38056,N_38431);
and U40408 (N_40408,N_38038,N_39803);
nor U40409 (N_40409,N_39440,N_38531);
xnor U40410 (N_40410,N_39279,N_39469);
xnor U40411 (N_40411,N_39787,N_39253);
nor U40412 (N_40412,N_39745,N_39087);
nand U40413 (N_40413,N_38569,N_39570);
nand U40414 (N_40414,N_39239,N_38300);
or U40415 (N_40415,N_39972,N_38743);
xnor U40416 (N_40416,N_39831,N_38500);
nand U40417 (N_40417,N_38540,N_39703);
or U40418 (N_40418,N_39545,N_38522);
and U40419 (N_40419,N_39257,N_38171);
nor U40420 (N_40420,N_38410,N_39721);
and U40421 (N_40421,N_39686,N_39039);
nor U40422 (N_40422,N_38241,N_38247);
nor U40423 (N_40423,N_39621,N_39242);
or U40424 (N_40424,N_38593,N_38624);
nor U40425 (N_40425,N_38755,N_39875);
and U40426 (N_40426,N_39355,N_38908);
or U40427 (N_40427,N_38824,N_39956);
nor U40428 (N_40428,N_39558,N_39727);
nor U40429 (N_40429,N_39359,N_38047);
or U40430 (N_40430,N_38666,N_39748);
nor U40431 (N_40431,N_38158,N_39147);
or U40432 (N_40432,N_38765,N_39771);
nand U40433 (N_40433,N_38334,N_39551);
xnor U40434 (N_40434,N_38262,N_39907);
xnor U40435 (N_40435,N_38136,N_39237);
nand U40436 (N_40436,N_38802,N_39051);
nand U40437 (N_40437,N_38190,N_38964);
nor U40438 (N_40438,N_38795,N_38769);
or U40439 (N_40439,N_38071,N_39906);
and U40440 (N_40440,N_39604,N_39678);
nand U40441 (N_40441,N_39915,N_38076);
or U40442 (N_40442,N_39044,N_39342);
and U40443 (N_40443,N_39471,N_38895);
and U40444 (N_40444,N_39438,N_38124);
and U40445 (N_40445,N_39122,N_38318);
nor U40446 (N_40446,N_39954,N_38400);
nand U40447 (N_40447,N_38445,N_38394);
nor U40448 (N_40448,N_39470,N_38120);
and U40449 (N_40449,N_38371,N_39387);
nand U40450 (N_40450,N_39580,N_38692);
nor U40451 (N_40451,N_39836,N_39704);
or U40452 (N_40452,N_39735,N_39230);
or U40453 (N_40453,N_39233,N_39754);
or U40454 (N_40454,N_39282,N_39234);
and U40455 (N_40455,N_38894,N_39884);
nor U40456 (N_40456,N_38817,N_38396);
and U40457 (N_40457,N_39432,N_38415);
nor U40458 (N_40458,N_39247,N_39560);
xnor U40459 (N_40459,N_38288,N_39810);
and U40460 (N_40460,N_39346,N_38074);
xnor U40461 (N_40461,N_38725,N_38797);
and U40462 (N_40462,N_38705,N_39651);
nor U40463 (N_40463,N_38229,N_38904);
nor U40464 (N_40464,N_38592,N_39311);
nand U40465 (N_40465,N_38749,N_39106);
nand U40466 (N_40466,N_39034,N_38427);
or U40467 (N_40467,N_38494,N_39159);
nand U40468 (N_40468,N_38656,N_39778);
and U40469 (N_40469,N_39588,N_39198);
and U40470 (N_40470,N_38773,N_39976);
nand U40471 (N_40471,N_38108,N_39614);
nand U40472 (N_40472,N_38905,N_38210);
or U40473 (N_40473,N_39394,N_39969);
nor U40474 (N_40474,N_38131,N_39567);
nand U40475 (N_40475,N_39893,N_39419);
nand U40476 (N_40476,N_38990,N_38344);
xnor U40477 (N_40477,N_39561,N_39049);
and U40478 (N_40478,N_39437,N_39116);
or U40479 (N_40479,N_38403,N_38701);
nand U40480 (N_40480,N_39071,N_38123);
nor U40481 (N_40481,N_38432,N_38675);
xnor U40482 (N_40482,N_39100,N_38691);
xor U40483 (N_40483,N_38726,N_38249);
nor U40484 (N_40484,N_39507,N_39082);
or U40485 (N_40485,N_39181,N_39050);
or U40486 (N_40486,N_38419,N_38356);
xnor U40487 (N_40487,N_38425,N_39768);
or U40488 (N_40488,N_38972,N_39737);
nor U40489 (N_40489,N_38097,N_39962);
or U40490 (N_40490,N_39814,N_39534);
xor U40491 (N_40491,N_39485,N_38714);
or U40492 (N_40492,N_38914,N_38564);
nor U40493 (N_40493,N_39497,N_38612);
and U40494 (N_40494,N_38484,N_39655);
xnor U40495 (N_40495,N_38023,N_38826);
xnor U40496 (N_40496,N_39632,N_38877);
nand U40497 (N_40497,N_39092,N_39008);
and U40498 (N_40498,N_39602,N_38764);
or U40499 (N_40499,N_38212,N_38201);
or U40500 (N_40500,N_38731,N_39564);
or U40501 (N_40501,N_39097,N_39284);
nor U40502 (N_40502,N_38832,N_39756);
nand U40503 (N_40503,N_38010,N_39799);
nand U40504 (N_40504,N_38652,N_38438);
xnor U40505 (N_40505,N_38465,N_38118);
or U40506 (N_40506,N_38974,N_39099);
xor U40507 (N_40507,N_39590,N_39848);
or U40508 (N_40508,N_38810,N_38946);
nand U40509 (N_40509,N_38672,N_38709);
and U40510 (N_40510,N_39708,N_39726);
or U40511 (N_40511,N_38129,N_39005);
xnor U40512 (N_40512,N_38757,N_39920);
nand U40513 (N_40513,N_38472,N_39073);
and U40514 (N_40514,N_39231,N_39515);
xor U40515 (N_40515,N_38092,N_39784);
or U40516 (N_40516,N_38279,N_38244);
or U40517 (N_40517,N_39921,N_38019);
and U40518 (N_40518,N_39764,N_38243);
xor U40519 (N_40519,N_39016,N_38357);
or U40520 (N_40520,N_38469,N_38111);
nand U40521 (N_40521,N_38690,N_38550);
or U40522 (N_40522,N_38621,N_38993);
and U40523 (N_40523,N_39720,N_39596);
or U40524 (N_40524,N_39993,N_38058);
nand U40525 (N_40525,N_39760,N_39900);
xor U40526 (N_40526,N_38599,N_39413);
nand U40527 (N_40527,N_38715,N_39015);
or U40528 (N_40528,N_38655,N_38537);
and U40529 (N_40529,N_38738,N_39297);
nor U40530 (N_40530,N_39559,N_38082);
and U40531 (N_40531,N_39547,N_38525);
or U40532 (N_40532,N_39488,N_38777);
nand U40533 (N_40533,N_39112,N_38146);
nand U40534 (N_40534,N_39828,N_38641);
nor U40535 (N_40535,N_38811,N_38127);
and U40536 (N_40536,N_39888,N_39995);
nor U40537 (N_40537,N_38784,N_39123);
xor U40538 (N_40538,N_39508,N_38083);
or U40539 (N_40539,N_39821,N_38857);
and U40540 (N_40540,N_39290,N_39697);
xnor U40541 (N_40541,N_39793,N_38984);
nor U40542 (N_40542,N_39289,N_39908);
or U40543 (N_40543,N_38109,N_39115);
nor U40544 (N_40544,N_39970,N_39223);
nand U40545 (N_40545,N_39830,N_38409);
xor U40546 (N_40546,N_38346,N_39388);
xnor U40547 (N_40547,N_38487,N_38677);
xnor U40548 (N_40548,N_39724,N_39527);
and U40549 (N_40549,N_38792,N_38245);
nor U40550 (N_40550,N_39148,N_38218);
xnor U40551 (N_40551,N_38821,N_39228);
nor U40552 (N_40552,N_38080,N_39877);
xor U40553 (N_40553,N_39254,N_39042);
or U40554 (N_40554,N_38355,N_38031);
nand U40555 (N_40555,N_39317,N_39332);
nor U40556 (N_40556,N_38386,N_38026);
and U40557 (N_40557,N_39725,N_38638);
nand U40558 (N_40558,N_38660,N_39695);
or U40559 (N_40559,N_38837,N_39903);
nor U40560 (N_40560,N_39058,N_39111);
nor U40561 (N_40561,N_38603,N_39445);
nand U40562 (N_40562,N_39334,N_39455);
or U40563 (N_40563,N_39981,N_39842);
xnor U40564 (N_40564,N_39260,N_38774);
and U40565 (N_40565,N_38874,N_39392);
and U40566 (N_40566,N_38625,N_38720);
xor U40567 (N_40567,N_39529,N_38467);
and U40568 (N_40568,N_38119,N_39535);
and U40569 (N_40569,N_38140,N_39029);
nand U40570 (N_40570,N_39288,N_39565);
or U40571 (N_40571,N_39522,N_39076);
or U40572 (N_40572,N_38462,N_38535);
and U40573 (N_40573,N_38292,N_38062);
xnor U40574 (N_40574,N_39227,N_39713);
xnor U40575 (N_40575,N_38882,N_39026);
and U40576 (N_40576,N_39405,N_38858);
or U40577 (N_40577,N_39141,N_38437);
nor U40578 (N_40578,N_39552,N_38340);
and U40579 (N_40579,N_39068,N_38611);
xor U40580 (N_40580,N_38889,N_38615);
nand U40581 (N_40581,N_38979,N_38022);
nor U40582 (N_40582,N_39923,N_39249);
xnor U40583 (N_40583,N_39262,N_39644);
xor U40584 (N_40584,N_38238,N_39133);
or U40585 (N_40585,N_39313,N_39918);
or U40586 (N_40586,N_39070,N_39439);
nand U40587 (N_40587,N_39390,N_39420);
xnor U40588 (N_40588,N_38044,N_39860);
or U40589 (N_40589,N_38678,N_38144);
or U40590 (N_40590,N_39666,N_39940);
nor U40591 (N_40591,N_39785,N_38565);
and U40592 (N_40592,N_39688,N_38285);
nand U40593 (N_40593,N_39654,N_39428);
and U40594 (N_40594,N_38639,N_39309);
and U40595 (N_40595,N_38913,N_39578);
or U40596 (N_40596,N_38197,N_39942);
nor U40597 (N_40597,N_38073,N_39441);
xor U40598 (N_40598,N_38150,N_38719);
xnor U40599 (N_40599,N_39117,N_38581);
xnor U40600 (N_40600,N_39371,N_39858);
and U40601 (N_40601,N_38316,N_39819);
or U40602 (N_40602,N_39944,N_38861);
nand U40603 (N_40603,N_39873,N_38457);
nand U40604 (N_40604,N_38096,N_39569);
or U40605 (N_40605,N_39218,N_38182);
or U40606 (N_40606,N_38079,N_38260);
or U40607 (N_40607,N_39344,N_39002);
nor U40608 (N_40608,N_38369,N_39730);
nand U40609 (N_40609,N_39946,N_38870);
xor U40610 (N_40610,N_39010,N_38732);
and U40611 (N_40611,N_39280,N_38647);
and U40612 (N_40612,N_38922,N_39809);
or U40613 (N_40613,N_39272,N_38230);
xor U40614 (N_40614,N_38168,N_39259);
nor U40615 (N_40615,N_39084,N_38319);
nand U40616 (N_40616,N_38027,N_38819);
or U40617 (N_40617,N_39667,N_38426);
xor U40618 (N_40618,N_39691,N_39794);
nand U40619 (N_40619,N_38711,N_39062);
or U40620 (N_40620,N_39606,N_38312);
nor U40621 (N_40621,N_39817,N_39630);
nand U40622 (N_40622,N_38825,N_39986);
and U40623 (N_40623,N_38294,N_38444);
and U40624 (N_40624,N_38206,N_39869);
nor U40625 (N_40625,N_39751,N_39562);
nand U40626 (N_40626,N_39483,N_38104);
or U40627 (N_40627,N_39867,N_38471);
or U40628 (N_40628,N_38509,N_39038);
xnor U40629 (N_40629,N_38976,N_38788);
and U40630 (N_40630,N_39633,N_39623);
or U40631 (N_40631,N_39292,N_38545);
nor U40632 (N_40632,N_38417,N_38822);
or U40633 (N_40633,N_39960,N_39072);
or U40634 (N_40634,N_38688,N_39659);
and U40635 (N_40635,N_38181,N_38101);
xnor U40636 (N_40636,N_38893,N_38477);
and U40637 (N_40637,N_38511,N_38528);
nor U40638 (N_40638,N_38744,N_38866);
nor U40639 (N_40639,N_39502,N_38682);
xor U40640 (N_40640,N_38735,N_39975);
xnor U40641 (N_40641,N_39700,N_39763);
xnor U40642 (N_40642,N_38627,N_39762);
xnor U40643 (N_40643,N_39665,N_39397);
or U40644 (N_40644,N_38841,N_38640);
or U40645 (N_40645,N_39626,N_38113);
and U40646 (N_40646,N_38915,N_38175);
and U40647 (N_40647,N_39186,N_38958);
or U40648 (N_40648,N_39790,N_38561);
and U40649 (N_40649,N_38362,N_39200);
and U40650 (N_40650,N_39680,N_39403);
nand U40651 (N_40651,N_38267,N_38233);
and U40652 (N_40652,N_39494,N_39622);
xor U40653 (N_40653,N_39518,N_39411);
xnor U40654 (N_40654,N_39637,N_38404);
and U40655 (N_40655,N_38207,N_38423);
and U40656 (N_40656,N_39493,N_39772);
nand U40657 (N_40657,N_38148,N_38138);
xor U40658 (N_40658,N_39243,N_38421);
nand U40659 (N_40659,N_38803,N_38336);
nor U40660 (N_40660,N_39834,N_38198);
nor U40661 (N_40661,N_38695,N_38930);
nor U40662 (N_40662,N_38401,N_38040);
or U40663 (N_40663,N_39382,N_39151);
and U40664 (N_40664,N_38173,N_38800);
xor U40665 (N_40665,N_39822,N_38375);
or U40666 (N_40666,N_39224,N_39407);
nor U40667 (N_40667,N_39155,N_39014);
nand U40668 (N_40668,N_38160,N_39456);
nor U40669 (N_40669,N_39750,N_38727);
xnor U40670 (N_40670,N_39496,N_39375);
or U40671 (N_40671,N_38380,N_38219);
nor U40672 (N_40672,N_39876,N_39963);
or U40673 (N_40673,N_39504,N_39040);
or U40674 (N_40674,N_39011,N_39672);
and U40675 (N_40675,N_38239,N_39180);
nor U40676 (N_40676,N_38888,N_39916);
and U40677 (N_40677,N_39629,N_38282);
xnor U40678 (N_40678,N_39377,N_38588);
xor U40679 (N_40679,N_38849,N_39516);
or U40680 (N_40680,N_39879,N_39299);
xor U40681 (N_40681,N_39554,N_39973);
or U40682 (N_40682,N_38526,N_39030);
or U40683 (N_40683,N_38240,N_39820);
nor U40684 (N_40684,N_39882,N_38546);
and U40685 (N_40685,N_39191,N_38037);
nand U40686 (N_40686,N_38917,N_39473);
nand U40687 (N_40687,N_38405,N_38838);
and U40688 (N_40688,N_39043,N_39268);
nor U40689 (N_40689,N_38662,N_39220);
xnor U40690 (N_40690,N_38696,N_39897);
nor U40691 (N_40691,N_39478,N_38189);
or U40692 (N_40692,N_38139,N_38395);
or U40693 (N_40693,N_38228,N_38508);
nor U40694 (N_40694,N_39712,N_38880);
nor U40695 (N_40695,N_38195,N_38163);
or U40696 (N_40696,N_39451,N_39326);
or U40697 (N_40697,N_39270,N_38456);
nand U40698 (N_40698,N_38623,N_39789);
or U40699 (N_40699,N_38203,N_39232);
or U40700 (N_40700,N_39222,N_38011);
nor U40701 (N_40701,N_38311,N_39971);
or U40702 (N_40702,N_38628,N_38556);
or U40703 (N_40703,N_39269,N_38752);
or U40704 (N_40704,N_39550,N_39285);
and U40705 (N_40705,N_39059,N_38614);
nand U40706 (N_40706,N_39019,N_38815);
or U40707 (N_40707,N_39274,N_38359);
xor U40708 (N_40708,N_38112,N_38505);
nor U40709 (N_40709,N_38503,N_38909);
and U40710 (N_40710,N_39267,N_38211);
and U40711 (N_40711,N_38064,N_39472);
and U40712 (N_40712,N_39399,N_39670);
xor U40713 (N_40713,N_38296,N_38906);
and U40714 (N_40714,N_39832,N_38793);
nand U40715 (N_40715,N_39168,N_38617);
xor U40716 (N_40716,N_38280,N_39930);
nand U40717 (N_40717,N_39553,N_38600);
or U40718 (N_40718,N_38377,N_38878);
nor U40719 (N_40719,N_39744,N_39804);
nor U40720 (N_40720,N_39475,N_38145);
xnor U40721 (N_40721,N_39107,N_39631);
or U40722 (N_40722,N_39036,N_38159);
and U40723 (N_40723,N_39805,N_39024);
or U40724 (N_40724,N_39719,N_39501);
nor U40725 (N_40725,N_38256,N_39859);
and U40726 (N_40726,N_38114,N_38081);
or U40727 (N_40727,N_39943,N_38571);
nand U40728 (N_40728,N_39236,N_39617);
xnor U40729 (N_40729,N_39003,N_38149);
nor U40730 (N_40730,N_38033,N_39597);
and U40731 (N_40731,N_38916,N_38277);
nor U40732 (N_40732,N_39369,N_38900);
nor U40733 (N_40733,N_38717,N_39856);
and U40734 (N_40734,N_38657,N_38553);
xnor U40735 (N_40735,N_39226,N_38169);
nor U40736 (N_40736,N_39931,N_38085);
nand U40737 (N_40737,N_39273,N_38057);
or U40738 (N_40738,N_38135,N_38679);
or U40739 (N_40739,N_38554,N_38066);
and U40740 (N_40740,N_38330,N_38852);
or U40741 (N_40741,N_38039,N_38665);
xor U40742 (N_40742,N_38306,N_39452);
and U40743 (N_40743,N_39216,N_39362);
nor U40744 (N_40744,N_38783,N_39783);
nand U40745 (N_40745,N_39530,N_39121);
nor U40746 (N_40746,N_39646,N_38434);
nand U40747 (N_40747,N_38251,N_39932);
or U40748 (N_40748,N_39600,N_38270);
or U40749 (N_40749,N_39149,N_38630);
and U40750 (N_40750,N_38301,N_39250);
and U40751 (N_40751,N_39531,N_38068);
nor U40752 (N_40752,N_38087,N_39080);
xor U40753 (N_40753,N_39395,N_39427);
xor U40754 (N_40754,N_38674,N_38643);
nand U40755 (N_40755,N_39928,N_38463);
and U40756 (N_40756,N_38954,N_39598);
or U40757 (N_40757,N_39769,N_38566);
nor U40758 (N_40758,N_39194,N_39047);
or U40759 (N_40759,N_38323,N_39556);
or U40760 (N_40760,N_38350,N_39687);
nand U40761 (N_40761,N_39924,N_38661);
and U40762 (N_40762,N_38390,N_39296);
nor U40763 (N_40763,N_38094,N_38728);
nand U40764 (N_40764,N_39964,N_39381);
nor U40765 (N_40765,N_39103,N_39829);
nand U40766 (N_40766,N_39409,N_39244);
or U40767 (N_40767,N_39816,N_38558);
or U40768 (N_40768,N_38043,N_38921);
or U40769 (N_40769,N_38368,N_39863);
and U40770 (N_40770,N_38552,N_39864);
xor U40771 (N_40771,N_38733,N_38667);
nand U40772 (N_40772,N_39780,N_38789);
nor U40773 (N_40773,N_38090,N_38000);
nand U40774 (N_40774,N_38758,N_38606);
xnor U40775 (N_40775,N_39513,N_39813);
nor U40776 (N_40776,N_39874,N_39676);
nor U40777 (N_40777,N_39069,N_39476);
nand U40778 (N_40778,N_38856,N_39480);
xor U40779 (N_40779,N_38162,N_38823);
nand U40780 (N_40780,N_39063,N_39258);
and U40781 (N_40781,N_39679,N_38942);
nor U40782 (N_40782,N_38041,N_38447);
nand U40783 (N_40783,N_38753,N_39523);
nand U40784 (N_40784,N_39357,N_39806);
or U40785 (N_40785,N_38345,N_38562);
and U40786 (N_40786,N_39098,N_38771);
xor U40787 (N_40787,N_39421,N_38816);
nand U40788 (N_40788,N_38422,N_39057);
nand U40789 (N_40789,N_38778,N_39136);
nand U40790 (N_40790,N_38863,N_38314);
nor U40791 (N_40791,N_39176,N_39759);
nor U40792 (N_40792,N_38613,N_39543);
or U40793 (N_40793,N_38110,N_39023);
nand U40794 (N_40794,N_39639,N_38947);
xnor U40795 (N_40795,N_38061,N_38973);
or U40796 (N_40796,N_39910,N_38281);
nor U40797 (N_40797,N_39425,N_38936);
and U40798 (N_40798,N_39911,N_39865);
or U40799 (N_40799,N_39374,N_39214);
nor U40800 (N_40800,N_38807,N_38308);
or U40801 (N_40801,N_39774,N_39156);
xor U40802 (N_40802,N_38965,N_39349);
nor U40803 (N_40803,N_38475,N_39415);
xor U40804 (N_40804,N_38560,N_39657);
nand U40805 (N_40805,N_38530,N_39851);
nor U40806 (N_40806,N_38790,N_38107);
xor U40807 (N_40807,N_38549,N_39638);
and U40808 (N_40808,N_38373,N_38102);
or U40809 (N_40809,N_38933,N_38598);
or U40810 (N_40810,N_38805,N_39539);
or U40811 (N_40811,N_39164,N_38363);
nand U40812 (N_40812,N_38383,N_38474);
or U40813 (N_40813,N_39177,N_39576);
and U40814 (N_40814,N_38302,N_39449);
nand U40815 (N_40815,N_38945,N_39190);
xnor U40816 (N_40816,N_38782,N_38470);
and U40817 (N_40817,N_38384,N_38310);
nor U40818 (N_40818,N_38468,N_38985);
and U40819 (N_40819,N_39711,N_39591);
nand U40820 (N_40820,N_38547,N_38850);
nand U40821 (N_40821,N_38583,N_39825);
nor U40822 (N_40822,N_39537,N_38125);
or U40823 (N_40823,N_39211,N_38209);
or U40824 (N_40824,N_38820,N_38418);
or U40825 (N_40825,N_38433,N_39210);
and U40826 (N_40826,N_39294,N_38017);
nand U40827 (N_40827,N_38884,N_39690);
xor U40828 (N_40828,N_39736,N_38454);
or U40829 (N_40829,N_38141,N_39849);
xor U40830 (N_40830,N_39315,N_39526);
xor U40831 (N_40831,N_38736,N_38012);
nor U40832 (N_40832,N_39054,N_39978);
and U40833 (N_40833,N_39328,N_39798);
nor U40834 (N_40834,N_38563,N_39714);
xor U40835 (N_40835,N_38594,N_39400);
or U40836 (N_40836,N_39414,N_38250);
nand U40837 (N_40837,N_38459,N_38779);
and U40838 (N_40838,N_38492,N_39161);
xnor U40839 (N_40839,N_38443,N_39775);
xor U40840 (N_40840,N_39264,N_38015);
nand U40841 (N_40841,N_38648,N_39854);
nor U40842 (N_40842,N_39682,N_39890);
and U40843 (N_40843,N_38446,N_39248);
and U40844 (N_40844,N_38451,N_38671);
and U40845 (N_40845,N_39109,N_39183);
xnor U40846 (N_40846,N_38737,N_39179);
xor U40847 (N_40847,N_39926,N_38559);
or U40848 (N_40848,N_38847,N_39933);
nand U40849 (N_40849,N_38257,N_38235);
xnor U40850 (N_40850,N_38473,N_38366);
and U40851 (N_40851,N_39533,N_39134);
and U40852 (N_40852,N_39594,N_39021);
nor U40853 (N_40853,N_38370,N_38747);
xnor U40854 (N_40854,N_38529,N_38266);
nor U40855 (N_40855,N_38988,N_38155);
and U40856 (N_40856,N_38199,N_39225);
and U40857 (N_40857,N_39577,N_39999);
nand U40858 (N_40858,N_38416,N_38751);
xnor U40859 (N_40859,N_39380,N_39027);
nand U40860 (N_40860,N_39579,N_39937);
xnor U40861 (N_40861,N_38575,N_38636);
and U40862 (N_40862,N_39126,N_38961);
nand U40863 (N_40863,N_38633,N_38885);
and U40864 (N_40864,N_38338,N_39584);
or U40865 (N_40865,N_38441,N_38996);
nor U40866 (N_40866,N_39074,N_38886);
nand U40867 (N_40867,N_39511,N_39827);
xor U40868 (N_40868,N_39090,N_38698);
and U40869 (N_40869,N_38969,N_38722);
xnor U40870 (N_40870,N_39500,N_39776);
and U40871 (N_40871,N_38937,N_38510);
nand U40872 (N_40872,N_38246,N_38304);
and U40873 (N_40873,N_38538,N_39603);
nor U40874 (N_40874,N_39681,N_39129);
xor U40875 (N_40875,N_38950,N_39065);
and U40876 (N_40876,N_38194,N_39683);
nand U40877 (N_40877,N_39132,N_39325);
or U40878 (N_40878,N_38488,N_38103);
nand U40879 (N_40879,N_39170,N_38142);
or U40880 (N_40880,N_39009,N_38284);
nor U40881 (N_40881,N_39673,N_38450);
or U40882 (N_40882,N_39717,N_38045);
nor U40883 (N_40883,N_39528,N_39353);
xnor U40884 (N_40884,N_38853,N_38602);
and U40885 (N_40885,N_38959,N_38166);
nor U40886 (N_40886,N_38767,N_38466);
xor U40887 (N_40887,N_39738,N_39761);
and U40888 (N_40888,N_39094,N_39178);
nor U40889 (N_40889,N_39378,N_38242);
nor U40890 (N_40890,N_39571,N_39293);
and U40891 (N_40891,N_39927,N_39807);
nor U40892 (N_40892,N_38925,N_38939);
xor U40893 (N_40893,N_38699,N_38828);
and U40894 (N_40894,N_38361,N_38938);
or U40895 (N_40895,N_39053,N_39373);
nand U40896 (N_40896,N_39521,N_39939);
nand U40897 (N_40897,N_39324,N_38460);
nand U40898 (N_40898,N_38430,N_38192);
nor U40899 (N_40899,N_38512,N_39689);
nand U40900 (N_40900,N_38645,N_39338);
or U40901 (N_40901,N_39004,N_38495);
or U40902 (N_40902,N_39193,N_38934);
xor U40903 (N_40903,N_38584,N_38291);
and U40904 (N_40904,N_38352,N_38098);
nor U40905 (N_40905,N_39628,N_38534);
and U40906 (N_40906,N_39998,N_38812);
and U40907 (N_40907,N_38227,N_39412);
xor U40908 (N_40908,N_39458,N_38851);
and U40909 (N_40909,N_38414,N_38983);
nand U40910 (N_40910,N_38089,N_39732);
nand U40911 (N_40911,N_39442,N_39152);
and U40912 (N_40912,N_39361,N_38215);
xnor U40913 (N_40913,N_38029,N_38903);
xor U40914 (N_40914,N_38729,N_38313);
nand U40915 (N_40915,N_38697,N_39499);
nor U40916 (N_40916,N_39012,N_39350);
xnor U40917 (N_40917,N_38685,N_39298);
or U40918 (N_40918,N_38276,N_39747);
xnor U40919 (N_40919,N_38573,N_39881);
nand U40920 (N_40920,N_38018,N_38809);
and U40921 (N_40921,N_38745,N_38232);
xnor U40922 (N_40922,N_38557,N_39077);
nor U40923 (N_40923,N_38428,N_39443);
nand U40924 (N_40924,N_39431,N_38496);
or U40925 (N_40925,N_39568,N_38590);
and U40926 (N_40926,N_38151,N_39966);
or U40927 (N_40927,N_39204,N_38261);
nand U40928 (N_40928,N_38269,N_39669);
and U40929 (N_40929,N_38364,N_39902);
xnor U40930 (N_40930,N_39781,N_39647);
and U40931 (N_40931,N_38049,N_39370);
nor U40932 (N_40932,N_38760,N_38180);
or U40933 (N_40933,N_38971,N_38873);
or U40934 (N_40934,N_38684,N_39627);
xnor U40935 (N_40935,N_39402,N_39462);
nor U40936 (N_40936,N_39089,N_39212);
xor U40937 (N_40937,N_38827,N_39896);
xnor U40938 (N_40938,N_39127,N_39119);
or U40939 (N_40939,N_39861,N_39348);
xor U40940 (N_40940,N_39323,N_38216);
or U40941 (N_40941,N_38977,N_38188);
nand U40942 (N_40942,N_39824,N_39912);
and U40943 (N_40943,N_38126,N_39000);
xnor U40944 (N_40944,N_39892,N_39477);
nor U40945 (N_40945,N_39705,N_39557);
nand U40946 (N_40946,N_39990,N_38164);
and U40947 (N_40947,N_38967,N_38680);
nand U40948 (N_40948,N_39277,N_39503);
nor U40949 (N_40949,N_38237,N_39201);
nor U40950 (N_40950,N_38172,N_39364);
nand U40951 (N_40951,N_39889,N_39202);
xor U40952 (N_40952,N_38297,N_39434);
nor U40953 (N_40953,N_38794,N_39319);
and U40954 (N_40954,N_39418,N_38265);
xnor U40955 (N_40955,N_38021,N_38252);
nand U40956 (N_40956,N_39067,N_38912);
nor U40957 (N_40957,N_39987,N_39675);
and U40958 (N_40958,N_38539,N_38263);
nor U40959 (N_40959,N_39291,N_38315);
and U40960 (N_40960,N_39985,N_39595);
nor U40961 (N_40961,N_38378,N_39166);
nor U40962 (N_40962,N_38706,N_38439);
xnor U40963 (N_40963,N_38932,N_39853);
nor U40964 (N_40964,N_39742,N_38956);
or U40965 (N_40965,N_38844,N_38536);
or U40966 (N_40966,N_39936,N_39624);
nand U40967 (N_40967,N_39495,N_38608);
or U40968 (N_40968,N_39173,N_38919);
nand U40969 (N_40969,N_39408,N_39352);
nand U40970 (N_40970,N_39358,N_38762);
xnor U40971 (N_40971,N_39716,N_38489);
and U40972 (N_40972,N_38887,N_39146);
nor U40973 (N_40973,N_39740,N_38205);
nor U40974 (N_40974,N_38902,N_39574);
xor U40975 (N_40975,N_38650,N_39331);
xnor U40976 (N_40976,N_39898,N_39949);
and U40977 (N_40977,N_39055,N_38572);
or U40978 (N_40978,N_38775,N_38708);
nand U40979 (N_40979,N_38596,N_39979);
nor U40980 (N_40980,N_39104,N_39929);
or U40981 (N_40981,N_39707,N_38220);
or U40982 (N_40982,N_39677,N_38587);
and U40983 (N_40983,N_39950,N_38610);
or U40984 (N_40984,N_39653,N_39105);
or U40985 (N_40985,N_39490,N_38927);
nor U40986 (N_40986,N_39424,N_38829);
nor U40987 (N_40987,N_39948,N_38609);
nor U40988 (N_40988,N_39143,N_39196);
or U40989 (N_40989,N_38106,N_38683);
or U40990 (N_40990,N_38272,N_38176);
xnor U40991 (N_40991,N_38981,N_39266);
and U40992 (N_40992,N_38307,N_39354);
and U40993 (N_40993,N_38875,N_38669);
nor U40994 (N_40994,N_39391,N_39729);
or U40995 (N_40995,N_39278,N_39128);
nor U40996 (N_40996,N_39197,N_38629);
and U40997 (N_40997,N_38167,N_39410);
nand U40998 (N_40998,N_38327,N_38322);
nand U40999 (N_40999,N_38455,N_39514);
xnor U41000 (N_41000,N_38189,N_39293);
or U41001 (N_41001,N_38166,N_39787);
nand U41002 (N_41002,N_38727,N_39637);
nand U41003 (N_41003,N_38391,N_38418);
nor U41004 (N_41004,N_39871,N_38167);
and U41005 (N_41005,N_38756,N_39785);
and U41006 (N_41006,N_38797,N_38025);
or U41007 (N_41007,N_39469,N_38138);
nand U41008 (N_41008,N_38870,N_38036);
and U41009 (N_41009,N_38532,N_39846);
xnor U41010 (N_41010,N_38145,N_39015);
nor U41011 (N_41011,N_39889,N_38825);
or U41012 (N_41012,N_38288,N_39371);
nand U41013 (N_41013,N_38684,N_39655);
xnor U41014 (N_41014,N_38553,N_39316);
xnor U41015 (N_41015,N_39747,N_38727);
nor U41016 (N_41016,N_39984,N_39821);
or U41017 (N_41017,N_38199,N_39142);
or U41018 (N_41018,N_38612,N_38753);
nor U41019 (N_41019,N_38109,N_38191);
or U41020 (N_41020,N_39317,N_39870);
or U41021 (N_41021,N_39283,N_39047);
and U41022 (N_41022,N_39037,N_39945);
and U41023 (N_41023,N_38602,N_39436);
and U41024 (N_41024,N_38955,N_38306);
xor U41025 (N_41025,N_39266,N_38159);
nor U41026 (N_41026,N_39394,N_39366);
and U41027 (N_41027,N_39387,N_39164);
and U41028 (N_41028,N_38049,N_39756);
and U41029 (N_41029,N_38810,N_38692);
nand U41030 (N_41030,N_38080,N_38918);
nor U41031 (N_41031,N_39779,N_39215);
or U41032 (N_41032,N_38393,N_38593);
nand U41033 (N_41033,N_39180,N_38426);
nand U41034 (N_41034,N_38118,N_39406);
xnor U41035 (N_41035,N_39499,N_39015);
nand U41036 (N_41036,N_39498,N_38314);
nand U41037 (N_41037,N_39969,N_38723);
or U41038 (N_41038,N_38030,N_39034);
and U41039 (N_41039,N_38114,N_38774);
xor U41040 (N_41040,N_38696,N_38312);
or U41041 (N_41041,N_39050,N_38187);
xor U41042 (N_41042,N_39854,N_38518);
or U41043 (N_41043,N_39873,N_38312);
and U41044 (N_41044,N_38341,N_38688);
nand U41045 (N_41045,N_38308,N_38036);
nor U41046 (N_41046,N_39804,N_38824);
or U41047 (N_41047,N_39202,N_38397);
nor U41048 (N_41048,N_39110,N_38809);
and U41049 (N_41049,N_39163,N_39950);
or U41050 (N_41050,N_38811,N_38216);
nand U41051 (N_41051,N_38328,N_39693);
or U41052 (N_41052,N_39427,N_39544);
nand U41053 (N_41053,N_39567,N_38479);
nor U41054 (N_41054,N_38595,N_38893);
nor U41055 (N_41055,N_38081,N_39845);
nor U41056 (N_41056,N_39508,N_39198);
and U41057 (N_41057,N_38209,N_39452);
nand U41058 (N_41058,N_39133,N_39472);
xor U41059 (N_41059,N_39653,N_38997);
nor U41060 (N_41060,N_38762,N_39771);
nand U41061 (N_41061,N_38486,N_38195);
nor U41062 (N_41062,N_38010,N_39270);
nor U41063 (N_41063,N_38425,N_38740);
xnor U41064 (N_41064,N_38099,N_39605);
and U41065 (N_41065,N_38740,N_38260);
nand U41066 (N_41066,N_39160,N_38349);
or U41067 (N_41067,N_38208,N_38617);
nor U41068 (N_41068,N_38572,N_39504);
or U41069 (N_41069,N_39265,N_39699);
nand U41070 (N_41070,N_39328,N_38356);
nand U41071 (N_41071,N_38139,N_39217);
nand U41072 (N_41072,N_38413,N_38038);
or U41073 (N_41073,N_38339,N_38263);
nor U41074 (N_41074,N_38239,N_38893);
or U41075 (N_41075,N_39678,N_38781);
and U41076 (N_41076,N_39999,N_39142);
nor U41077 (N_41077,N_39205,N_38382);
or U41078 (N_41078,N_39272,N_39222);
xnor U41079 (N_41079,N_39747,N_38716);
or U41080 (N_41080,N_38568,N_38377);
xnor U41081 (N_41081,N_39578,N_39613);
nor U41082 (N_41082,N_39948,N_38343);
nand U41083 (N_41083,N_38571,N_39988);
nand U41084 (N_41084,N_39097,N_39517);
or U41085 (N_41085,N_38393,N_39588);
xor U41086 (N_41086,N_38263,N_39339);
nand U41087 (N_41087,N_39544,N_39961);
or U41088 (N_41088,N_38186,N_39442);
xor U41089 (N_41089,N_39065,N_38743);
or U41090 (N_41090,N_39573,N_38619);
or U41091 (N_41091,N_39558,N_38614);
xnor U41092 (N_41092,N_38325,N_39367);
nor U41093 (N_41093,N_38573,N_39274);
or U41094 (N_41094,N_38310,N_38814);
and U41095 (N_41095,N_39385,N_39667);
nor U41096 (N_41096,N_39193,N_38020);
nand U41097 (N_41097,N_39014,N_39030);
and U41098 (N_41098,N_38825,N_38915);
nand U41099 (N_41099,N_38451,N_39780);
or U41100 (N_41100,N_38351,N_38135);
nor U41101 (N_41101,N_38086,N_39247);
or U41102 (N_41102,N_38151,N_39361);
nor U41103 (N_41103,N_39215,N_38506);
nor U41104 (N_41104,N_39981,N_38226);
and U41105 (N_41105,N_39432,N_38171);
or U41106 (N_41106,N_39914,N_38816);
nand U41107 (N_41107,N_38897,N_38962);
and U41108 (N_41108,N_38004,N_39528);
nand U41109 (N_41109,N_38191,N_38133);
xor U41110 (N_41110,N_39712,N_39452);
xor U41111 (N_41111,N_39918,N_39259);
or U41112 (N_41112,N_39872,N_38306);
and U41113 (N_41113,N_39610,N_39164);
nor U41114 (N_41114,N_39191,N_39443);
or U41115 (N_41115,N_38299,N_39398);
and U41116 (N_41116,N_39695,N_39067);
xnor U41117 (N_41117,N_38448,N_38793);
and U41118 (N_41118,N_38303,N_38573);
nor U41119 (N_41119,N_39509,N_39329);
xor U41120 (N_41120,N_38373,N_38152);
xnor U41121 (N_41121,N_39497,N_39592);
nand U41122 (N_41122,N_39383,N_39620);
and U41123 (N_41123,N_39281,N_38980);
and U41124 (N_41124,N_39407,N_39578);
and U41125 (N_41125,N_39271,N_38187);
and U41126 (N_41126,N_38726,N_38993);
xnor U41127 (N_41127,N_38724,N_38736);
nand U41128 (N_41128,N_39375,N_38178);
and U41129 (N_41129,N_39783,N_39889);
nor U41130 (N_41130,N_38785,N_39515);
and U41131 (N_41131,N_38939,N_39773);
xnor U41132 (N_41132,N_39866,N_38982);
xor U41133 (N_41133,N_38518,N_39886);
nand U41134 (N_41134,N_38275,N_38891);
nor U41135 (N_41135,N_39831,N_39920);
nand U41136 (N_41136,N_39022,N_38788);
and U41137 (N_41137,N_38913,N_38694);
or U41138 (N_41138,N_39549,N_38425);
nor U41139 (N_41139,N_39153,N_39584);
or U41140 (N_41140,N_39670,N_39635);
xnor U41141 (N_41141,N_38963,N_39609);
or U41142 (N_41142,N_38047,N_39452);
xor U41143 (N_41143,N_38430,N_38321);
or U41144 (N_41144,N_38188,N_39123);
nor U41145 (N_41145,N_38006,N_39096);
and U41146 (N_41146,N_38649,N_38238);
or U41147 (N_41147,N_38495,N_38299);
and U41148 (N_41148,N_38433,N_39840);
nand U41149 (N_41149,N_38287,N_38792);
nand U41150 (N_41150,N_38583,N_39121);
and U41151 (N_41151,N_38974,N_38045);
nand U41152 (N_41152,N_39610,N_39846);
or U41153 (N_41153,N_38143,N_38997);
nand U41154 (N_41154,N_38971,N_38758);
nand U41155 (N_41155,N_38167,N_39506);
and U41156 (N_41156,N_39764,N_39171);
nor U41157 (N_41157,N_38796,N_39057);
xor U41158 (N_41158,N_38394,N_38218);
nor U41159 (N_41159,N_38805,N_38637);
nor U41160 (N_41160,N_39541,N_39282);
xnor U41161 (N_41161,N_39886,N_39985);
or U41162 (N_41162,N_39620,N_39608);
and U41163 (N_41163,N_38525,N_39780);
and U41164 (N_41164,N_38280,N_38580);
xor U41165 (N_41165,N_38284,N_39885);
xnor U41166 (N_41166,N_38153,N_39502);
nor U41167 (N_41167,N_39813,N_38709);
and U41168 (N_41168,N_39302,N_39713);
or U41169 (N_41169,N_38097,N_39345);
nand U41170 (N_41170,N_38853,N_38774);
or U41171 (N_41171,N_39984,N_39497);
nor U41172 (N_41172,N_39112,N_38902);
or U41173 (N_41173,N_39090,N_39138);
or U41174 (N_41174,N_38064,N_39790);
and U41175 (N_41175,N_38375,N_39910);
nor U41176 (N_41176,N_39988,N_39706);
or U41177 (N_41177,N_38295,N_39137);
xnor U41178 (N_41178,N_38943,N_39810);
xor U41179 (N_41179,N_39266,N_39945);
and U41180 (N_41180,N_39283,N_38299);
xnor U41181 (N_41181,N_38490,N_38413);
nor U41182 (N_41182,N_38459,N_39058);
nand U41183 (N_41183,N_39704,N_39583);
nor U41184 (N_41184,N_39789,N_39513);
nor U41185 (N_41185,N_39477,N_38448);
or U41186 (N_41186,N_38470,N_38602);
xnor U41187 (N_41187,N_39805,N_38238);
nor U41188 (N_41188,N_39201,N_39338);
nand U41189 (N_41189,N_39183,N_38019);
and U41190 (N_41190,N_38052,N_39381);
and U41191 (N_41191,N_38871,N_39976);
nand U41192 (N_41192,N_38702,N_38739);
nand U41193 (N_41193,N_39596,N_39265);
nand U41194 (N_41194,N_38859,N_39706);
xor U41195 (N_41195,N_38104,N_38887);
xnor U41196 (N_41196,N_39330,N_39454);
or U41197 (N_41197,N_38434,N_38529);
nand U41198 (N_41198,N_39933,N_38624);
or U41199 (N_41199,N_39921,N_39420);
and U41200 (N_41200,N_39840,N_38831);
xnor U41201 (N_41201,N_39539,N_38276);
nor U41202 (N_41202,N_38029,N_38202);
and U41203 (N_41203,N_38502,N_39417);
nor U41204 (N_41204,N_38558,N_38883);
and U41205 (N_41205,N_38175,N_38264);
nor U41206 (N_41206,N_38506,N_38712);
nor U41207 (N_41207,N_38415,N_38589);
xnor U41208 (N_41208,N_39883,N_38772);
xnor U41209 (N_41209,N_39806,N_38504);
or U41210 (N_41210,N_38239,N_39761);
nand U41211 (N_41211,N_38313,N_39630);
or U41212 (N_41212,N_38516,N_38674);
nor U41213 (N_41213,N_38590,N_38517);
xnor U41214 (N_41214,N_39727,N_39257);
and U41215 (N_41215,N_39505,N_38418);
nor U41216 (N_41216,N_38667,N_39932);
and U41217 (N_41217,N_39735,N_38306);
xnor U41218 (N_41218,N_39654,N_38387);
nand U41219 (N_41219,N_39678,N_38391);
xor U41220 (N_41220,N_38861,N_39279);
or U41221 (N_41221,N_39734,N_39564);
nor U41222 (N_41222,N_38793,N_38814);
nor U41223 (N_41223,N_38948,N_38666);
and U41224 (N_41224,N_38573,N_39983);
nor U41225 (N_41225,N_38762,N_38702);
nand U41226 (N_41226,N_39028,N_39786);
xor U41227 (N_41227,N_38558,N_38900);
or U41228 (N_41228,N_38386,N_39198);
xor U41229 (N_41229,N_39435,N_39950);
nand U41230 (N_41230,N_39067,N_39923);
xnor U41231 (N_41231,N_39028,N_39409);
xor U41232 (N_41232,N_39641,N_38169);
and U41233 (N_41233,N_39615,N_39271);
and U41234 (N_41234,N_39042,N_38983);
and U41235 (N_41235,N_38139,N_38960);
nor U41236 (N_41236,N_39263,N_39251);
nor U41237 (N_41237,N_39710,N_39422);
or U41238 (N_41238,N_39219,N_39800);
or U41239 (N_41239,N_39687,N_39551);
xnor U41240 (N_41240,N_38015,N_39124);
or U41241 (N_41241,N_39454,N_39612);
nand U41242 (N_41242,N_38852,N_38034);
or U41243 (N_41243,N_39526,N_38353);
xnor U41244 (N_41244,N_39893,N_39722);
and U41245 (N_41245,N_38833,N_39333);
or U41246 (N_41246,N_38942,N_39612);
xor U41247 (N_41247,N_38860,N_38068);
nand U41248 (N_41248,N_39139,N_38848);
and U41249 (N_41249,N_38352,N_39814);
or U41250 (N_41250,N_38785,N_38281);
and U41251 (N_41251,N_38513,N_39664);
and U41252 (N_41252,N_39970,N_38887);
xor U41253 (N_41253,N_38995,N_38230);
xnor U41254 (N_41254,N_39909,N_39646);
and U41255 (N_41255,N_39310,N_39982);
nand U41256 (N_41256,N_38431,N_39790);
nor U41257 (N_41257,N_38189,N_39020);
nand U41258 (N_41258,N_38194,N_39754);
nor U41259 (N_41259,N_39128,N_39665);
xor U41260 (N_41260,N_38824,N_39502);
nor U41261 (N_41261,N_38110,N_38064);
and U41262 (N_41262,N_39608,N_38414);
and U41263 (N_41263,N_38265,N_38920);
and U41264 (N_41264,N_39489,N_39298);
and U41265 (N_41265,N_38176,N_38980);
xor U41266 (N_41266,N_39625,N_38771);
nand U41267 (N_41267,N_39579,N_39111);
and U41268 (N_41268,N_38668,N_38014);
nor U41269 (N_41269,N_39737,N_39391);
xnor U41270 (N_41270,N_39772,N_38851);
xnor U41271 (N_41271,N_39308,N_39814);
and U41272 (N_41272,N_39793,N_38668);
xnor U41273 (N_41273,N_39175,N_38021);
xnor U41274 (N_41274,N_39535,N_39476);
or U41275 (N_41275,N_38403,N_38757);
and U41276 (N_41276,N_38806,N_39722);
xor U41277 (N_41277,N_39291,N_39068);
or U41278 (N_41278,N_38615,N_38501);
xor U41279 (N_41279,N_39807,N_38399);
xor U41280 (N_41280,N_38657,N_39687);
xor U41281 (N_41281,N_39188,N_38782);
nand U41282 (N_41282,N_38613,N_38982);
or U41283 (N_41283,N_39218,N_38541);
xor U41284 (N_41284,N_38058,N_39526);
or U41285 (N_41285,N_39597,N_38173);
and U41286 (N_41286,N_39931,N_39355);
or U41287 (N_41287,N_39739,N_39388);
nand U41288 (N_41288,N_38012,N_39775);
and U41289 (N_41289,N_38818,N_39352);
nor U41290 (N_41290,N_39163,N_39486);
or U41291 (N_41291,N_39922,N_38273);
nand U41292 (N_41292,N_39394,N_39142);
nor U41293 (N_41293,N_39667,N_38664);
nor U41294 (N_41294,N_39544,N_38967);
xnor U41295 (N_41295,N_38808,N_38246);
and U41296 (N_41296,N_39066,N_39651);
and U41297 (N_41297,N_39346,N_39307);
nor U41298 (N_41298,N_39936,N_38550);
nor U41299 (N_41299,N_39895,N_39986);
and U41300 (N_41300,N_38793,N_38821);
or U41301 (N_41301,N_38688,N_38837);
and U41302 (N_41302,N_39034,N_38250);
nor U41303 (N_41303,N_39769,N_39523);
and U41304 (N_41304,N_38098,N_39814);
nor U41305 (N_41305,N_38185,N_39158);
and U41306 (N_41306,N_39646,N_38723);
nand U41307 (N_41307,N_38762,N_38593);
and U41308 (N_41308,N_39824,N_39984);
nand U41309 (N_41309,N_39148,N_39077);
or U41310 (N_41310,N_39140,N_39496);
xnor U41311 (N_41311,N_39987,N_39641);
or U41312 (N_41312,N_38269,N_38498);
nand U41313 (N_41313,N_38017,N_38392);
or U41314 (N_41314,N_38581,N_38712);
xor U41315 (N_41315,N_38960,N_39458);
nand U41316 (N_41316,N_38643,N_38711);
and U41317 (N_41317,N_39732,N_38807);
and U41318 (N_41318,N_39364,N_38296);
and U41319 (N_41319,N_38264,N_39073);
xor U41320 (N_41320,N_39410,N_39177);
xor U41321 (N_41321,N_39611,N_38683);
nor U41322 (N_41322,N_39077,N_39034);
xnor U41323 (N_41323,N_38273,N_39670);
xnor U41324 (N_41324,N_39917,N_38467);
nor U41325 (N_41325,N_38157,N_38590);
nand U41326 (N_41326,N_39729,N_38149);
nand U41327 (N_41327,N_38946,N_39943);
and U41328 (N_41328,N_38503,N_38647);
nor U41329 (N_41329,N_39772,N_38515);
or U41330 (N_41330,N_39484,N_39510);
or U41331 (N_41331,N_39259,N_39409);
and U41332 (N_41332,N_39476,N_39895);
nand U41333 (N_41333,N_39269,N_39729);
or U41334 (N_41334,N_38926,N_39531);
nand U41335 (N_41335,N_39346,N_39266);
nand U41336 (N_41336,N_38779,N_39624);
and U41337 (N_41337,N_39817,N_38045);
and U41338 (N_41338,N_39352,N_39293);
and U41339 (N_41339,N_39498,N_39784);
or U41340 (N_41340,N_38223,N_39837);
nand U41341 (N_41341,N_38921,N_39036);
xor U41342 (N_41342,N_39637,N_39024);
and U41343 (N_41343,N_39846,N_39529);
xnor U41344 (N_41344,N_38118,N_39887);
xor U41345 (N_41345,N_38676,N_38369);
xnor U41346 (N_41346,N_39838,N_39881);
nand U41347 (N_41347,N_38421,N_39418);
nand U41348 (N_41348,N_38129,N_38820);
nand U41349 (N_41349,N_39726,N_39741);
nor U41350 (N_41350,N_39059,N_38720);
nand U41351 (N_41351,N_39309,N_38957);
nor U41352 (N_41352,N_39809,N_39635);
nor U41353 (N_41353,N_38569,N_38181);
nor U41354 (N_41354,N_38033,N_38332);
or U41355 (N_41355,N_38313,N_39295);
nor U41356 (N_41356,N_38048,N_38308);
xnor U41357 (N_41357,N_39373,N_39930);
nor U41358 (N_41358,N_38880,N_39409);
xor U41359 (N_41359,N_38278,N_38740);
and U41360 (N_41360,N_39853,N_39434);
nand U41361 (N_41361,N_39464,N_38176);
nor U41362 (N_41362,N_38261,N_39435);
and U41363 (N_41363,N_38917,N_39890);
and U41364 (N_41364,N_39601,N_39874);
xnor U41365 (N_41365,N_38533,N_39267);
nor U41366 (N_41366,N_38291,N_39371);
nor U41367 (N_41367,N_39127,N_39299);
and U41368 (N_41368,N_39300,N_39024);
and U41369 (N_41369,N_39590,N_38353);
or U41370 (N_41370,N_39848,N_39378);
and U41371 (N_41371,N_39398,N_38435);
nand U41372 (N_41372,N_38904,N_38185);
or U41373 (N_41373,N_39462,N_39617);
or U41374 (N_41374,N_39424,N_39482);
nor U41375 (N_41375,N_38295,N_38836);
or U41376 (N_41376,N_39812,N_39685);
and U41377 (N_41377,N_38110,N_39045);
and U41378 (N_41378,N_39659,N_39300);
and U41379 (N_41379,N_39421,N_38089);
xnor U41380 (N_41380,N_39195,N_38387);
nor U41381 (N_41381,N_39725,N_38043);
xor U41382 (N_41382,N_38886,N_38406);
and U41383 (N_41383,N_38852,N_38880);
or U41384 (N_41384,N_38200,N_39208);
or U41385 (N_41385,N_38988,N_38875);
nor U41386 (N_41386,N_38196,N_39478);
xnor U41387 (N_41387,N_39263,N_39840);
nor U41388 (N_41388,N_38743,N_39488);
and U41389 (N_41389,N_38366,N_39068);
and U41390 (N_41390,N_38572,N_39163);
nor U41391 (N_41391,N_39404,N_39381);
or U41392 (N_41392,N_39380,N_39245);
xnor U41393 (N_41393,N_39481,N_38609);
and U41394 (N_41394,N_38807,N_39434);
xor U41395 (N_41395,N_38274,N_38500);
xor U41396 (N_41396,N_38851,N_39560);
and U41397 (N_41397,N_39342,N_38611);
nand U41398 (N_41398,N_39632,N_38746);
xnor U41399 (N_41399,N_39041,N_38329);
xor U41400 (N_41400,N_38334,N_38957);
or U41401 (N_41401,N_39106,N_39458);
or U41402 (N_41402,N_38639,N_39571);
or U41403 (N_41403,N_39429,N_38392);
xor U41404 (N_41404,N_39537,N_38243);
nor U41405 (N_41405,N_39747,N_39396);
nor U41406 (N_41406,N_38098,N_38151);
nor U41407 (N_41407,N_39850,N_39831);
and U41408 (N_41408,N_38378,N_39164);
nand U41409 (N_41409,N_39518,N_38343);
and U41410 (N_41410,N_38205,N_38183);
nand U41411 (N_41411,N_39940,N_39906);
nand U41412 (N_41412,N_39501,N_38944);
or U41413 (N_41413,N_38602,N_38801);
and U41414 (N_41414,N_39632,N_39117);
or U41415 (N_41415,N_39044,N_38583);
or U41416 (N_41416,N_39005,N_38565);
nand U41417 (N_41417,N_39198,N_39185);
and U41418 (N_41418,N_39219,N_39198);
nand U41419 (N_41419,N_39027,N_39950);
nand U41420 (N_41420,N_39849,N_38278);
and U41421 (N_41421,N_39374,N_39284);
nand U41422 (N_41422,N_38615,N_38192);
nor U41423 (N_41423,N_39874,N_39226);
xor U41424 (N_41424,N_38982,N_38378);
or U41425 (N_41425,N_38267,N_39382);
nor U41426 (N_41426,N_39958,N_39921);
xnor U41427 (N_41427,N_38550,N_38144);
and U41428 (N_41428,N_38730,N_38473);
and U41429 (N_41429,N_39757,N_38228);
and U41430 (N_41430,N_39480,N_38450);
and U41431 (N_41431,N_38006,N_38279);
or U41432 (N_41432,N_38859,N_38482);
xnor U41433 (N_41433,N_38484,N_39043);
nand U41434 (N_41434,N_38548,N_39683);
or U41435 (N_41435,N_39014,N_38267);
xor U41436 (N_41436,N_39959,N_39874);
xor U41437 (N_41437,N_38520,N_38146);
xnor U41438 (N_41438,N_39290,N_39574);
nand U41439 (N_41439,N_39397,N_39840);
and U41440 (N_41440,N_38551,N_39303);
xnor U41441 (N_41441,N_39420,N_39887);
xor U41442 (N_41442,N_38525,N_39728);
nand U41443 (N_41443,N_39369,N_38569);
or U41444 (N_41444,N_39758,N_38899);
xnor U41445 (N_41445,N_38437,N_38560);
and U41446 (N_41446,N_38462,N_38791);
nand U41447 (N_41447,N_38322,N_38571);
nand U41448 (N_41448,N_39871,N_38869);
or U41449 (N_41449,N_38493,N_38059);
nand U41450 (N_41450,N_39584,N_38601);
xor U41451 (N_41451,N_39134,N_39977);
nor U41452 (N_41452,N_39062,N_39636);
and U41453 (N_41453,N_38764,N_38356);
nand U41454 (N_41454,N_38620,N_38250);
xor U41455 (N_41455,N_39967,N_39640);
xnor U41456 (N_41456,N_38236,N_38453);
or U41457 (N_41457,N_39414,N_39946);
and U41458 (N_41458,N_39002,N_38022);
and U41459 (N_41459,N_38805,N_39757);
xnor U41460 (N_41460,N_39561,N_39655);
or U41461 (N_41461,N_39133,N_39283);
nor U41462 (N_41462,N_39853,N_38645);
nand U41463 (N_41463,N_39669,N_38467);
nand U41464 (N_41464,N_38048,N_38385);
or U41465 (N_41465,N_39394,N_39605);
nor U41466 (N_41466,N_39940,N_39613);
xor U41467 (N_41467,N_39111,N_38353);
nor U41468 (N_41468,N_38432,N_38791);
nand U41469 (N_41469,N_39725,N_39305);
nor U41470 (N_41470,N_38234,N_39510);
and U41471 (N_41471,N_38277,N_39011);
and U41472 (N_41472,N_38827,N_39890);
nand U41473 (N_41473,N_38958,N_38043);
xor U41474 (N_41474,N_39597,N_39405);
nand U41475 (N_41475,N_39415,N_39185);
xor U41476 (N_41476,N_39499,N_39942);
or U41477 (N_41477,N_39983,N_39052);
nand U41478 (N_41478,N_39163,N_39583);
or U41479 (N_41479,N_38951,N_39312);
xor U41480 (N_41480,N_38325,N_39538);
and U41481 (N_41481,N_38789,N_38255);
xor U41482 (N_41482,N_39555,N_39897);
or U41483 (N_41483,N_38347,N_39477);
or U41484 (N_41484,N_38639,N_39313);
nand U41485 (N_41485,N_39256,N_39327);
nor U41486 (N_41486,N_39974,N_39535);
and U41487 (N_41487,N_39478,N_38927);
or U41488 (N_41488,N_38198,N_38913);
or U41489 (N_41489,N_39296,N_39923);
nor U41490 (N_41490,N_39882,N_38307);
xnor U41491 (N_41491,N_39235,N_39130);
or U41492 (N_41492,N_39284,N_39375);
xor U41493 (N_41493,N_38944,N_39424);
or U41494 (N_41494,N_38473,N_39095);
and U41495 (N_41495,N_38616,N_39924);
nand U41496 (N_41496,N_38072,N_39602);
xnor U41497 (N_41497,N_39343,N_39329);
nor U41498 (N_41498,N_39401,N_38042);
nand U41499 (N_41499,N_39193,N_39347);
xnor U41500 (N_41500,N_39308,N_38237);
nor U41501 (N_41501,N_39533,N_39086);
and U41502 (N_41502,N_38059,N_39537);
nor U41503 (N_41503,N_38576,N_38132);
and U41504 (N_41504,N_38875,N_39823);
nand U41505 (N_41505,N_38218,N_39531);
nor U41506 (N_41506,N_38045,N_39033);
and U41507 (N_41507,N_39060,N_39879);
xor U41508 (N_41508,N_38085,N_39982);
nand U41509 (N_41509,N_39275,N_38290);
or U41510 (N_41510,N_39584,N_38451);
nand U41511 (N_41511,N_38821,N_39708);
xnor U41512 (N_41512,N_39490,N_38331);
or U41513 (N_41513,N_38618,N_38872);
nor U41514 (N_41514,N_39140,N_39701);
xnor U41515 (N_41515,N_39268,N_39896);
or U41516 (N_41516,N_38553,N_38969);
or U41517 (N_41517,N_38570,N_39178);
nand U41518 (N_41518,N_39001,N_38495);
or U41519 (N_41519,N_38249,N_38767);
and U41520 (N_41520,N_39777,N_38427);
or U41521 (N_41521,N_38378,N_38673);
nor U41522 (N_41522,N_38275,N_38417);
xor U41523 (N_41523,N_39453,N_39297);
nor U41524 (N_41524,N_39176,N_38497);
xor U41525 (N_41525,N_38319,N_39806);
xor U41526 (N_41526,N_39734,N_39194);
nand U41527 (N_41527,N_38631,N_39517);
xor U41528 (N_41528,N_38661,N_38075);
and U41529 (N_41529,N_39681,N_39034);
nor U41530 (N_41530,N_39036,N_39556);
nand U41531 (N_41531,N_39521,N_38919);
xor U41532 (N_41532,N_39809,N_38676);
xnor U41533 (N_41533,N_38045,N_38209);
or U41534 (N_41534,N_39436,N_39391);
xnor U41535 (N_41535,N_38296,N_39300);
xor U41536 (N_41536,N_38259,N_38819);
xor U41537 (N_41537,N_39318,N_38985);
xor U41538 (N_41538,N_38442,N_38319);
or U41539 (N_41539,N_38533,N_38744);
nor U41540 (N_41540,N_38562,N_39792);
or U41541 (N_41541,N_39881,N_39094);
and U41542 (N_41542,N_39774,N_38875);
and U41543 (N_41543,N_39697,N_38942);
xnor U41544 (N_41544,N_39269,N_39460);
and U41545 (N_41545,N_39009,N_39751);
and U41546 (N_41546,N_38417,N_38069);
nor U41547 (N_41547,N_39146,N_39304);
and U41548 (N_41548,N_39580,N_38107);
xnor U41549 (N_41549,N_38004,N_38078);
xor U41550 (N_41550,N_39052,N_39461);
xor U41551 (N_41551,N_38436,N_39791);
nand U41552 (N_41552,N_39959,N_39060);
xnor U41553 (N_41553,N_39745,N_39114);
nor U41554 (N_41554,N_38762,N_39393);
or U41555 (N_41555,N_38765,N_39990);
nor U41556 (N_41556,N_38152,N_39399);
nand U41557 (N_41557,N_39611,N_39055);
nor U41558 (N_41558,N_39399,N_38837);
nand U41559 (N_41559,N_39390,N_39201);
xor U41560 (N_41560,N_39092,N_38091);
nand U41561 (N_41561,N_38404,N_39331);
nor U41562 (N_41562,N_39297,N_38154);
or U41563 (N_41563,N_38949,N_39782);
nand U41564 (N_41564,N_38805,N_38565);
xor U41565 (N_41565,N_38931,N_38705);
xnor U41566 (N_41566,N_38627,N_38456);
nand U41567 (N_41567,N_39828,N_38033);
xnor U41568 (N_41568,N_38865,N_39811);
and U41569 (N_41569,N_39367,N_39262);
xnor U41570 (N_41570,N_39065,N_39028);
nand U41571 (N_41571,N_39928,N_39743);
and U41572 (N_41572,N_38938,N_39596);
nor U41573 (N_41573,N_39358,N_38109);
or U41574 (N_41574,N_38369,N_38874);
or U41575 (N_41575,N_39495,N_39813);
nand U41576 (N_41576,N_39992,N_38354);
nor U41577 (N_41577,N_39031,N_39320);
nor U41578 (N_41578,N_39561,N_38665);
nor U41579 (N_41579,N_38117,N_38986);
or U41580 (N_41580,N_39770,N_39516);
or U41581 (N_41581,N_39306,N_38386);
nand U41582 (N_41582,N_39691,N_39729);
nand U41583 (N_41583,N_38213,N_38938);
xor U41584 (N_41584,N_38845,N_39483);
and U41585 (N_41585,N_38771,N_38944);
and U41586 (N_41586,N_38531,N_39359);
and U41587 (N_41587,N_39433,N_39024);
nor U41588 (N_41588,N_39265,N_38832);
nand U41589 (N_41589,N_39646,N_38732);
nand U41590 (N_41590,N_38737,N_38064);
and U41591 (N_41591,N_38179,N_38062);
or U41592 (N_41592,N_38200,N_38817);
xnor U41593 (N_41593,N_39649,N_39743);
or U41594 (N_41594,N_38469,N_38192);
nor U41595 (N_41595,N_39681,N_38932);
or U41596 (N_41596,N_39121,N_39277);
or U41597 (N_41597,N_39765,N_39166);
or U41598 (N_41598,N_38037,N_38627);
nor U41599 (N_41599,N_38237,N_38795);
xnor U41600 (N_41600,N_38145,N_38423);
nand U41601 (N_41601,N_39867,N_39836);
and U41602 (N_41602,N_38932,N_38988);
nor U41603 (N_41603,N_39220,N_39021);
nor U41604 (N_41604,N_39938,N_39907);
nand U41605 (N_41605,N_38732,N_39049);
nand U41606 (N_41606,N_39149,N_39184);
nand U41607 (N_41607,N_39967,N_38726);
nor U41608 (N_41608,N_39960,N_39376);
and U41609 (N_41609,N_39133,N_38356);
or U41610 (N_41610,N_38802,N_38645);
and U41611 (N_41611,N_38380,N_39372);
nor U41612 (N_41612,N_39966,N_38415);
nor U41613 (N_41613,N_38079,N_38709);
and U41614 (N_41614,N_39233,N_38990);
and U41615 (N_41615,N_38739,N_38218);
xor U41616 (N_41616,N_38771,N_38972);
and U41617 (N_41617,N_39906,N_39838);
xor U41618 (N_41618,N_38720,N_38920);
nor U41619 (N_41619,N_39305,N_38429);
and U41620 (N_41620,N_39203,N_39862);
nand U41621 (N_41621,N_39889,N_38738);
xor U41622 (N_41622,N_39732,N_39823);
xor U41623 (N_41623,N_38858,N_38422);
xnor U41624 (N_41624,N_39671,N_38884);
nor U41625 (N_41625,N_39795,N_38121);
and U41626 (N_41626,N_38951,N_38628);
xor U41627 (N_41627,N_39173,N_39988);
and U41628 (N_41628,N_39232,N_39098);
nor U41629 (N_41629,N_38521,N_39802);
nand U41630 (N_41630,N_39282,N_39298);
or U41631 (N_41631,N_39685,N_39981);
nor U41632 (N_41632,N_38935,N_38135);
xnor U41633 (N_41633,N_39372,N_38792);
xnor U41634 (N_41634,N_38148,N_39816);
nand U41635 (N_41635,N_38392,N_38950);
nand U41636 (N_41636,N_38439,N_39728);
and U41637 (N_41637,N_39452,N_38998);
or U41638 (N_41638,N_39883,N_38408);
xor U41639 (N_41639,N_39510,N_39662);
and U41640 (N_41640,N_38830,N_38245);
or U41641 (N_41641,N_39884,N_38612);
or U41642 (N_41642,N_39988,N_38873);
nor U41643 (N_41643,N_39652,N_39954);
nor U41644 (N_41644,N_38609,N_38614);
nand U41645 (N_41645,N_39876,N_38230);
nor U41646 (N_41646,N_39402,N_38555);
nand U41647 (N_41647,N_38528,N_39760);
xnor U41648 (N_41648,N_39861,N_39598);
or U41649 (N_41649,N_39354,N_39519);
nand U41650 (N_41650,N_38748,N_39879);
and U41651 (N_41651,N_39110,N_39273);
xor U41652 (N_41652,N_38274,N_38214);
or U41653 (N_41653,N_39261,N_39446);
nand U41654 (N_41654,N_39345,N_38957);
nor U41655 (N_41655,N_38537,N_38180);
nand U41656 (N_41656,N_38716,N_38938);
or U41657 (N_41657,N_39909,N_38133);
and U41658 (N_41658,N_39273,N_39675);
or U41659 (N_41659,N_38978,N_38506);
xor U41660 (N_41660,N_38568,N_39194);
or U41661 (N_41661,N_38870,N_39353);
nand U41662 (N_41662,N_39557,N_39310);
and U41663 (N_41663,N_38012,N_38355);
xnor U41664 (N_41664,N_39582,N_39506);
and U41665 (N_41665,N_39329,N_39950);
nand U41666 (N_41666,N_38765,N_39447);
or U41667 (N_41667,N_39741,N_38983);
xnor U41668 (N_41668,N_39011,N_39104);
nand U41669 (N_41669,N_39302,N_39010);
or U41670 (N_41670,N_39421,N_39998);
or U41671 (N_41671,N_39712,N_38669);
xor U41672 (N_41672,N_38294,N_38034);
and U41673 (N_41673,N_38646,N_38073);
nand U41674 (N_41674,N_39178,N_39742);
nor U41675 (N_41675,N_39155,N_39405);
and U41676 (N_41676,N_39484,N_39142);
or U41677 (N_41677,N_38467,N_39688);
or U41678 (N_41678,N_38858,N_39533);
xnor U41679 (N_41679,N_38136,N_38244);
and U41680 (N_41680,N_38341,N_38578);
and U41681 (N_41681,N_38114,N_38144);
and U41682 (N_41682,N_38126,N_38118);
or U41683 (N_41683,N_39273,N_38611);
nor U41684 (N_41684,N_39413,N_38154);
nand U41685 (N_41685,N_39876,N_38854);
and U41686 (N_41686,N_39505,N_38036);
xor U41687 (N_41687,N_39530,N_38395);
nand U41688 (N_41688,N_39253,N_39603);
or U41689 (N_41689,N_39089,N_38171);
nand U41690 (N_41690,N_39451,N_39607);
and U41691 (N_41691,N_39845,N_39831);
nand U41692 (N_41692,N_39706,N_38724);
xor U41693 (N_41693,N_38145,N_38367);
xor U41694 (N_41694,N_38506,N_38840);
and U41695 (N_41695,N_39580,N_38976);
or U41696 (N_41696,N_38530,N_39941);
xor U41697 (N_41697,N_38860,N_38671);
nand U41698 (N_41698,N_39662,N_39368);
xor U41699 (N_41699,N_38740,N_38039);
nand U41700 (N_41700,N_39248,N_39052);
nor U41701 (N_41701,N_39291,N_38331);
nand U41702 (N_41702,N_38248,N_39683);
or U41703 (N_41703,N_39128,N_38308);
nand U41704 (N_41704,N_38356,N_39891);
xnor U41705 (N_41705,N_38250,N_39363);
and U41706 (N_41706,N_38795,N_39557);
xor U41707 (N_41707,N_38389,N_39653);
nand U41708 (N_41708,N_38257,N_39182);
nor U41709 (N_41709,N_38905,N_38276);
xnor U41710 (N_41710,N_38137,N_39401);
xor U41711 (N_41711,N_39730,N_39350);
xnor U41712 (N_41712,N_38037,N_39118);
nand U41713 (N_41713,N_38723,N_38791);
or U41714 (N_41714,N_38238,N_39862);
or U41715 (N_41715,N_38895,N_38255);
xor U41716 (N_41716,N_39171,N_38167);
and U41717 (N_41717,N_38726,N_39096);
nand U41718 (N_41718,N_38846,N_39733);
nand U41719 (N_41719,N_38715,N_39338);
xor U41720 (N_41720,N_39259,N_39371);
nor U41721 (N_41721,N_39646,N_39413);
xnor U41722 (N_41722,N_39691,N_39611);
nor U41723 (N_41723,N_39579,N_39610);
nor U41724 (N_41724,N_38798,N_39315);
xor U41725 (N_41725,N_38927,N_39485);
nor U41726 (N_41726,N_38193,N_38444);
nor U41727 (N_41727,N_39532,N_38498);
nor U41728 (N_41728,N_38268,N_39434);
and U41729 (N_41729,N_39076,N_38975);
or U41730 (N_41730,N_39935,N_38967);
nor U41731 (N_41731,N_39228,N_38349);
or U41732 (N_41732,N_38422,N_38245);
and U41733 (N_41733,N_38541,N_39081);
xor U41734 (N_41734,N_39761,N_38964);
xnor U41735 (N_41735,N_38057,N_38061);
xnor U41736 (N_41736,N_39396,N_39478);
or U41737 (N_41737,N_39898,N_39835);
nor U41738 (N_41738,N_39139,N_38523);
or U41739 (N_41739,N_39859,N_38876);
nor U41740 (N_41740,N_39620,N_39810);
nand U41741 (N_41741,N_39327,N_38074);
nor U41742 (N_41742,N_38896,N_38029);
and U41743 (N_41743,N_38056,N_39284);
and U41744 (N_41744,N_39007,N_38796);
nor U41745 (N_41745,N_39917,N_39101);
and U41746 (N_41746,N_39500,N_38256);
nand U41747 (N_41747,N_39617,N_38609);
nor U41748 (N_41748,N_39284,N_39200);
nor U41749 (N_41749,N_39195,N_39326);
nand U41750 (N_41750,N_39773,N_39134);
or U41751 (N_41751,N_38351,N_39594);
nor U41752 (N_41752,N_39791,N_39376);
or U41753 (N_41753,N_39361,N_39921);
nor U41754 (N_41754,N_38100,N_38731);
nor U41755 (N_41755,N_38149,N_38534);
nand U41756 (N_41756,N_38254,N_39991);
and U41757 (N_41757,N_38925,N_39619);
and U41758 (N_41758,N_39161,N_39334);
and U41759 (N_41759,N_39905,N_39121);
nor U41760 (N_41760,N_39431,N_38910);
nand U41761 (N_41761,N_38572,N_38739);
xor U41762 (N_41762,N_39524,N_39561);
xnor U41763 (N_41763,N_38180,N_38142);
xnor U41764 (N_41764,N_38853,N_39836);
xor U41765 (N_41765,N_38269,N_39734);
nor U41766 (N_41766,N_39857,N_39988);
nor U41767 (N_41767,N_39669,N_39738);
nor U41768 (N_41768,N_39561,N_38312);
and U41769 (N_41769,N_38141,N_38088);
xnor U41770 (N_41770,N_39090,N_38240);
nor U41771 (N_41771,N_38852,N_39658);
and U41772 (N_41772,N_38251,N_38289);
or U41773 (N_41773,N_39426,N_39232);
nor U41774 (N_41774,N_39368,N_39367);
or U41775 (N_41775,N_39969,N_38560);
or U41776 (N_41776,N_38324,N_38294);
nor U41777 (N_41777,N_39483,N_39002);
xor U41778 (N_41778,N_38219,N_39609);
xor U41779 (N_41779,N_39289,N_39656);
nor U41780 (N_41780,N_39327,N_38288);
and U41781 (N_41781,N_39322,N_39023);
and U41782 (N_41782,N_39690,N_39600);
xor U41783 (N_41783,N_38988,N_39493);
and U41784 (N_41784,N_39020,N_38635);
and U41785 (N_41785,N_39635,N_39549);
nand U41786 (N_41786,N_39464,N_38240);
and U41787 (N_41787,N_39230,N_39051);
and U41788 (N_41788,N_39810,N_39285);
xor U41789 (N_41789,N_39374,N_38923);
or U41790 (N_41790,N_39561,N_39354);
nor U41791 (N_41791,N_39730,N_38959);
and U41792 (N_41792,N_38908,N_38430);
xnor U41793 (N_41793,N_39248,N_38022);
and U41794 (N_41794,N_38566,N_39910);
or U41795 (N_41795,N_38056,N_39697);
and U41796 (N_41796,N_38065,N_39160);
and U41797 (N_41797,N_39612,N_38990);
nand U41798 (N_41798,N_38900,N_39559);
nand U41799 (N_41799,N_39253,N_38686);
nor U41800 (N_41800,N_39291,N_38513);
xnor U41801 (N_41801,N_39560,N_38712);
xnor U41802 (N_41802,N_39633,N_39898);
nand U41803 (N_41803,N_38446,N_39812);
or U41804 (N_41804,N_39572,N_39790);
and U41805 (N_41805,N_39176,N_38994);
nand U41806 (N_41806,N_39931,N_38879);
and U41807 (N_41807,N_38362,N_39510);
xor U41808 (N_41808,N_38424,N_38594);
or U41809 (N_41809,N_39261,N_39502);
xnor U41810 (N_41810,N_39351,N_38603);
xor U41811 (N_41811,N_39283,N_39325);
or U41812 (N_41812,N_38261,N_39569);
and U41813 (N_41813,N_39451,N_39029);
xnor U41814 (N_41814,N_39108,N_38427);
xnor U41815 (N_41815,N_39031,N_38186);
nor U41816 (N_41816,N_38185,N_39661);
xor U41817 (N_41817,N_38740,N_39037);
or U41818 (N_41818,N_38632,N_39258);
and U41819 (N_41819,N_38348,N_39149);
nor U41820 (N_41820,N_38888,N_39826);
and U41821 (N_41821,N_39813,N_39141);
or U41822 (N_41822,N_38166,N_38915);
xnor U41823 (N_41823,N_39272,N_38326);
nor U41824 (N_41824,N_38493,N_38550);
nand U41825 (N_41825,N_38656,N_38971);
nand U41826 (N_41826,N_38512,N_39562);
nor U41827 (N_41827,N_39639,N_39723);
nor U41828 (N_41828,N_39875,N_39118);
or U41829 (N_41829,N_39536,N_39021);
nand U41830 (N_41830,N_38982,N_38482);
or U41831 (N_41831,N_38307,N_39901);
and U41832 (N_41832,N_39261,N_38093);
nand U41833 (N_41833,N_39190,N_39115);
nand U41834 (N_41834,N_38222,N_38925);
and U41835 (N_41835,N_38242,N_38244);
or U41836 (N_41836,N_39884,N_39172);
xnor U41837 (N_41837,N_38350,N_38385);
xnor U41838 (N_41838,N_38182,N_39160);
xnor U41839 (N_41839,N_39950,N_39604);
xor U41840 (N_41840,N_39065,N_38477);
or U41841 (N_41841,N_38647,N_39809);
nand U41842 (N_41842,N_39918,N_38668);
and U41843 (N_41843,N_39387,N_39907);
or U41844 (N_41844,N_38078,N_39355);
nand U41845 (N_41845,N_38649,N_38568);
nor U41846 (N_41846,N_39428,N_38751);
nand U41847 (N_41847,N_38591,N_39613);
or U41848 (N_41848,N_38236,N_38118);
nand U41849 (N_41849,N_38248,N_38234);
nor U41850 (N_41850,N_39468,N_38522);
xor U41851 (N_41851,N_38036,N_38978);
xor U41852 (N_41852,N_38454,N_39854);
or U41853 (N_41853,N_38352,N_38025);
or U41854 (N_41854,N_39260,N_39047);
nand U41855 (N_41855,N_38386,N_38030);
nor U41856 (N_41856,N_38013,N_38482);
or U41857 (N_41857,N_39739,N_39827);
and U41858 (N_41858,N_38317,N_38967);
or U41859 (N_41859,N_38617,N_39612);
and U41860 (N_41860,N_39720,N_38421);
xnor U41861 (N_41861,N_39791,N_39140);
nor U41862 (N_41862,N_39803,N_39800);
and U41863 (N_41863,N_39725,N_38718);
and U41864 (N_41864,N_39063,N_38407);
nor U41865 (N_41865,N_38468,N_38984);
xor U41866 (N_41866,N_38550,N_39225);
xnor U41867 (N_41867,N_38654,N_38914);
and U41868 (N_41868,N_39583,N_38827);
nand U41869 (N_41869,N_38643,N_39770);
nand U41870 (N_41870,N_39864,N_39143);
nand U41871 (N_41871,N_39146,N_39103);
and U41872 (N_41872,N_38963,N_39083);
nor U41873 (N_41873,N_39908,N_38724);
xnor U41874 (N_41874,N_39220,N_39664);
or U41875 (N_41875,N_39997,N_39790);
nor U41876 (N_41876,N_39695,N_39650);
and U41877 (N_41877,N_39983,N_39931);
nand U41878 (N_41878,N_39842,N_38463);
or U41879 (N_41879,N_39610,N_38932);
nand U41880 (N_41880,N_39437,N_38766);
or U41881 (N_41881,N_39328,N_39892);
xor U41882 (N_41882,N_39327,N_39727);
xor U41883 (N_41883,N_39726,N_39971);
nand U41884 (N_41884,N_38026,N_39833);
xnor U41885 (N_41885,N_38053,N_38167);
nand U41886 (N_41886,N_39803,N_39065);
or U41887 (N_41887,N_39440,N_39452);
nand U41888 (N_41888,N_38195,N_38768);
and U41889 (N_41889,N_39623,N_39620);
or U41890 (N_41890,N_38067,N_38813);
or U41891 (N_41891,N_39710,N_39756);
nand U41892 (N_41892,N_39158,N_38284);
and U41893 (N_41893,N_39569,N_38943);
and U41894 (N_41894,N_38375,N_38472);
nor U41895 (N_41895,N_38120,N_38365);
xnor U41896 (N_41896,N_39224,N_39135);
or U41897 (N_41897,N_39123,N_38513);
and U41898 (N_41898,N_38245,N_39283);
and U41899 (N_41899,N_38308,N_38466);
or U41900 (N_41900,N_39186,N_39728);
and U41901 (N_41901,N_39320,N_39819);
xor U41902 (N_41902,N_39515,N_39439);
xnor U41903 (N_41903,N_38417,N_39968);
nand U41904 (N_41904,N_38915,N_39920);
or U41905 (N_41905,N_39993,N_38304);
xnor U41906 (N_41906,N_39004,N_39372);
and U41907 (N_41907,N_38316,N_39535);
nand U41908 (N_41908,N_39354,N_39205);
xnor U41909 (N_41909,N_38570,N_38189);
nand U41910 (N_41910,N_38131,N_38152);
or U41911 (N_41911,N_39788,N_38321);
or U41912 (N_41912,N_39062,N_38960);
nor U41913 (N_41913,N_39566,N_39723);
or U41914 (N_41914,N_39219,N_39574);
nor U41915 (N_41915,N_38752,N_39025);
and U41916 (N_41916,N_39396,N_38917);
nor U41917 (N_41917,N_39838,N_38292);
and U41918 (N_41918,N_39620,N_38839);
nor U41919 (N_41919,N_38487,N_38053);
and U41920 (N_41920,N_39149,N_39737);
and U41921 (N_41921,N_39043,N_39583);
xor U41922 (N_41922,N_39117,N_39000);
xor U41923 (N_41923,N_38760,N_38261);
nand U41924 (N_41924,N_39141,N_39467);
and U41925 (N_41925,N_38873,N_38304);
and U41926 (N_41926,N_39388,N_38669);
nor U41927 (N_41927,N_38231,N_39140);
nand U41928 (N_41928,N_38953,N_39463);
xnor U41929 (N_41929,N_39651,N_38396);
xnor U41930 (N_41930,N_38246,N_39416);
or U41931 (N_41931,N_39977,N_38225);
nor U41932 (N_41932,N_38590,N_39924);
or U41933 (N_41933,N_38438,N_39340);
nand U41934 (N_41934,N_39416,N_38168);
nand U41935 (N_41935,N_39930,N_38422);
and U41936 (N_41936,N_38428,N_39702);
nor U41937 (N_41937,N_38478,N_38330);
xor U41938 (N_41938,N_38396,N_38681);
or U41939 (N_41939,N_39411,N_39476);
nand U41940 (N_41940,N_39478,N_39682);
nand U41941 (N_41941,N_38084,N_38904);
xnor U41942 (N_41942,N_39611,N_39143);
nand U41943 (N_41943,N_38157,N_39734);
xnor U41944 (N_41944,N_38975,N_39528);
nor U41945 (N_41945,N_38798,N_38153);
and U41946 (N_41946,N_38985,N_38809);
and U41947 (N_41947,N_38278,N_38479);
nand U41948 (N_41948,N_39028,N_38255);
and U41949 (N_41949,N_39958,N_38983);
or U41950 (N_41950,N_39142,N_38142);
or U41951 (N_41951,N_38668,N_38898);
xor U41952 (N_41952,N_39073,N_39313);
or U41953 (N_41953,N_39129,N_38906);
nand U41954 (N_41954,N_38243,N_38815);
nor U41955 (N_41955,N_39608,N_39347);
nor U41956 (N_41956,N_38840,N_38130);
or U41957 (N_41957,N_39511,N_38606);
and U41958 (N_41958,N_39554,N_38520);
xor U41959 (N_41959,N_38888,N_39190);
nor U41960 (N_41960,N_38469,N_39169);
or U41961 (N_41961,N_39824,N_39782);
or U41962 (N_41962,N_39734,N_38739);
nand U41963 (N_41963,N_39630,N_38136);
xnor U41964 (N_41964,N_39849,N_38384);
xnor U41965 (N_41965,N_38054,N_39484);
nor U41966 (N_41966,N_39577,N_39878);
or U41967 (N_41967,N_38309,N_39626);
nor U41968 (N_41968,N_39969,N_38114);
nand U41969 (N_41969,N_38706,N_38259);
or U41970 (N_41970,N_39190,N_38075);
or U41971 (N_41971,N_38323,N_38712);
nor U41972 (N_41972,N_39342,N_39565);
and U41973 (N_41973,N_38206,N_38835);
nor U41974 (N_41974,N_39687,N_38141);
and U41975 (N_41975,N_39343,N_39570);
xnor U41976 (N_41976,N_39823,N_38389);
or U41977 (N_41977,N_39090,N_38522);
nand U41978 (N_41978,N_38781,N_39968);
and U41979 (N_41979,N_39177,N_38593);
nand U41980 (N_41980,N_39989,N_38918);
xor U41981 (N_41981,N_39288,N_38768);
nand U41982 (N_41982,N_39656,N_38521);
or U41983 (N_41983,N_39193,N_39089);
or U41984 (N_41984,N_38540,N_39276);
and U41985 (N_41985,N_38220,N_38337);
and U41986 (N_41986,N_39636,N_38753);
and U41987 (N_41987,N_39763,N_38121);
and U41988 (N_41988,N_38316,N_39793);
and U41989 (N_41989,N_38796,N_38105);
or U41990 (N_41990,N_39618,N_38532);
or U41991 (N_41991,N_39383,N_39589);
nor U41992 (N_41992,N_38730,N_39844);
or U41993 (N_41993,N_39497,N_38993);
nand U41994 (N_41994,N_38344,N_39459);
and U41995 (N_41995,N_38386,N_38961);
or U41996 (N_41996,N_39047,N_38698);
nand U41997 (N_41997,N_39823,N_39149);
and U41998 (N_41998,N_38290,N_39994);
and U41999 (N_41999,N_39134,N_38370);
and U42000 (N_42000,N_40120,N_41362);
nand U42001 (N_42001,N_41448,N_41695);
nand U42002 (N_42002,N_41822,N_40730);
nor U42003 (N_42003,N_40649,N_40622);
and U42004 (N_42004,N_40435,N_40158);
nor U42005 (N_42005,N_40684,N_41838);
or U42006 (N_42006,N_40849,N_40045);
nor U42007 (N_42007,N_41542,N_40752);
nand U42008 (N_42008,N_40034,N_41901);
xnor U42009 (N_42009,N_40526,N_40431);
and U42010 (N_42010,N_40258,N_40966);
and U42011 (N_42011,N_41200,N_41507);
nand U42012 (N_42012,N_41475,N_40842);
or U42013 (N_42013,N_40825,N_40553);
nor U42014 (N_42014,N_40385,N_40074);
xor U42015 (N_42015,N_40169,N_41890);
or U42016 (N_42016,N_41461,N_40582);
and U42017 (N_42017,N_41817,N_41739);
nand U42018 (N_42018,N_41368,N_41498);
or U42019 (N_42019,N_40661,N_41968);
nor U42020 (N_42020,N_41298,N_41038);
nor U42021 (N_42021,N_40341,N_40065);
nor U42022 (N_42022,N_40038,N_40619);
xor U42023 (N_42023,N_40066,N_40519);
xnor U42024 (N_42024,N_41676,N_41066);
or U42025 (N_42025,N_41651,N_40240);
or U42026 (N_42026,N_40625,N_41563);
nor U42027 (N_42027,N_40122,N_41658);
or U42028 (N_42028,N_41440,N_41320);
and U42029 (N_42029,N_40010,N_41081);
xnor U42030 (N_42030,N_40837,N_40709);
nor U42031 (N_42031,N_40504,N_41694);
nand U42032 (N_42032,N_40404,N_41029);
or U42033 (N_42033,N_40474,N_41662);
and U42034 (N_42034,N_41574,N_41030);
and U42035 (N_42035,N_41585,N_40206);
and U42036 (N_42036,N_41364,N_40401);
or U42037 (N_42037,N_40182,N_41996);
nor U42038 (N_42038,N_41554,N_40803);
and U42039 (N_42039,N_40471,N_41823);
nand U42040 (N_42040,N_41270,N_41224);
xnor U42041 (N_42041,N_41677,N_41557);
nand U42042 (N_42042,N_41023,N_41580);
xor U42043 (N_42043,N_40561,N_40815);
xor U42044 (N_42044,N_40921,N_41025);
and U42045 (N_42045,N_41407,N_41700);
or U42046 (N_42046,N_41722,N_40807);
nand U42047 (N_42047,N_41210,N_41894);
nand U42048 (N_42048,N_41121,N_41887);
or U42049 (N_42049,N_41331,N_41741);
nand U42050 (N_42050,N_40745,N_40071);
xnor U42051 (N_42051,N_41184,N_40874);
nand U42052 (N_42052,N_41426,N_41047);
xor U42053 (N_42053,N_40953,N_40925);
and U42054 (N_42054,N_40779,N_41503);
and U42055 (N_42055,N_40718,N_41821);
nand U42056 (N_42056,N_41644,N_40774);
xor U42057 (N_42057,N_40928,N_40972);
nand U42058 (N_42058,N_41275,N_40156);
or U42059 (N_42059,N_41199,N_41683);
nor U42060 (N_42060,N_40390,N_40556);
and U42061 (N_42061,N_40729,N_41245);
nand U42062 (N_42062,N_41979,N_40562);
nor U42063 (N_42063,N_40734,N_41064);
nor U42064 (N_42064,N_41055,N_40545);
xnor U42065 (N_42065,N_40163,N_40941);
nand U42066 (N_42066,N_41451,N_40869);
xor U42067 (N_42067,N_41516,N_41036);
nor U42068 (N_42068,N_41975,N_40985);
or U42069 (N_42069,N_41246,N_40155);
nand U42070 (N_42070,N_41386,N_40129);
nor U42071 (N_42071,N_41022,N_40084);
and U42072 (N_42072,N_41005,N_41929);
nand U42073 (N_42073,N_40005,N_40466);
or U42074 (N_42074,N_40127,N_40114);
xnor U42075 (N_42075,N_41988,N_41450);
or U42076 (N_42076,N_41665,N_40975);
nand U42077 (N_42077,N_41434,N_40300);
nor U42078 (N_42078,N_40929,N_40805);
xnor U42079 (N_42079,N_40469,N_40472);
nor U42080 (N_42080,N_40133,N_41849);
nand U42081 (N_42081,N_40707,N_40688);
xor U42082 (N_42082,N_40678,N_40560);
or U42083 (N_42083,N_41203,N_40040);
or U42084 (N_42084,N_41202,N_41759);
and U42085 (N_42085,N_40783,N_41909);
nand U42086 (N_42086,N_40655,N_40213);
xor U42087 (N_42087,N_40047,N_41714);
or U42088 (N_42088,N_40420,N_41963);
and U42089 (N_42089,N_41619,N_41630);
nor U42090 (N_42090,N_40778,N_41396);
xnor U42091 (N_42091,N_41690,N_40682);
nand U42092 (N_42092,N_41835,N_41139);
nor U42093 (N_42093,N_41430,N_40824);
and U42094 (N_42094,N_40342,N_40876);
and U42095 (N_42095,N_40125,N_41089);
nor U42096 (N_42096,N_41462,N_40224);
nand U42097 (N_42097,N_41663,N_41325);
xor U42098 (N_42098,N_40376,N_40748);
nor U42099 (N_42099,N_41514,N_41708);
nor U42100 (N_42100,N_41073,N_40188);
xor U42101 (N_42101,N_41777,N_40836);
nor U42102 (N_42102,N_41871,N_40199);
nand U42103 (N_42103,N_41330,N_41416);
nand U42104 (N_42104,N_40676,N_40260);
nand U42105 (N_42105,N_41218,N_41295);
and U42106 (N_42106,N_40981,N_40489);
nand U42107 (N_42107,N_40360,N_40398);
or U42108 (N_42108,N_41208,N_41880);
or U42109 (N_42109,N_41457,N_41226);
and U42110 (N_42110,N_40605,N_40765);
or U42111 (N_42111,N_41276,N_40980);
nand U42112 (N_42112,N_41117,N_40830);
nand U42113 (N_42113,N_40136,N_41467);
and U42114 (N_42114,N_40712,N_41189);
xnor U42115 (N_42115,N_41806,N_40699);
nand U42116 (N_42116,N_40934,N_41950);
nand U42117 (N_42117,N_40381,N_41941);
nor U42118 (N_42118,N_41031,N_40723);
nor U42119 (N_42119,N_41054,N_40324);
or U42120 (N_42120,N_41102,N_41209);
nand U42121 (N_42121,N_40166,N_40701);
nor U42122 (N_42122,N_41789,N_40875);
or U42123 (N_42123,N_40256,N_40064);
nor U42124 (N_42124,N_40174,N_41687);
or U42125 (N_42125,N_41783,N_40895);
xnor U42126 (N_42126,N_41537,N_40440);
and U42127 (N_42127,N_40490,N_40202);
and U42128 (N_42128,N_41279,N_41405);
nand U42129 (N_42129,N_41414,N_40732);
xnor U42130 (N_42130,N_41755,N_41934);
xor U42131 (N_42131,N_40646,N_40116);
xor U42132 (N_42132,N_41671,N_40104);
or U42133 (N_42133,N_41911,N_41072);
and U42134 (N_42134,N_41422,N_41876);
and U42135 (N_42135,N_40069,N_41869);
or U42136 (N_42136,N_41341,N_41845);
nor U42137 (N_42137,N_40759,N_41425);
and U42138 (N_42138,N_41940,N_40184);
xor U42139 (N_42139,N_41281,N_41385);
nor U42140 (N_42140,N_40738,N_40677);
and U42141 (N_42141,N_40500,N_40578);
xor U42142 (N_42142,N_41088,N_41258);
xor U42143 (N_42143,N_41660,N_41427);
and U42144 (N_42144,N_41390,N_40464);
and U42145 (N_42145,N_41936,N_41985);
xnor U42146 (N_42146,N_40019,N_40549);
nor U42147 (N_42147,N_41858,N_41169);
xor U42148 (N_42148,N_40691,N_40534);
nor U42149 (N_42149,N_40354,N_41844);
nand U42150 (N_42150,N_41518,N_41626);
xnor U42151 (N_42151,N_41155,N_41327);
xnor U42152 (N_42152,N_41446,N_40742);
or U42153 (N_42153,N_41972,N_41253);
or U42154 (N_42154,N_41244,N_41346);
nand U42155 (N_42155,N_41052,N_40427);
xor U42156 (N_42156,N_40126,N_40329);
or U42157 (N_42157,N_40920,N_41361);
nor U42158 (N_42158,N_40667,N_40236);
and U42159 (N_42159,N_41681,N_40009);
nand U42160 (N_42160,N_41757,N_40516);
or U42161 (N_42161,N_40461,N_40105);
nor U42162 (N_42162,N_40580,N_41194);
and U42163 (N_42163,N_41527,N_40986);
or U42164 (N_42164,N_40444,N_40512);
nand U42165 (N_42165,N_41750,N_41540);
xor U42166 (N_42166,N_41198,N_41573);
xor U42167 (N_42167,N_41292,N_41381);
xor U42168 (N_42168,N_41302,N_41283);
xnor U42169 (N_42169,N_41277,N_41893);
and U42170 (N_42170,N_40450,N_40958);
nand U42171 (N_42171,N_40995,N_41534);
xnor U42172 (N_42172,N_41581,N_40608);
nor U42173 (N_42173,N_40072,N_40097);
nor U42174 (N_42174,N_41846,N_40901);
or U42175 (N_42175,N_40909,N_41696);
nor U42176 (N_42176,N_40770,N_40651);
and U42177 (N_42177,N_41884,N_40579);
or U42178 (N_42178,N_40772,N_40281);
xor U42179 (N_42179,N_41657,N_41753);
and U42180 (N_42180,N_41008,N_41832);
nand U42181 (N_42181,N_40724,N_40799);
and U42182 (N_42182,N_41485,N_41483);
or U42183 (N_42183,N_41191,N_41810);
xor U42184 (N_42184,N_41667,N_40755);
or U42185 (N_42185,N_41977,N_41267);
or U42186 (N_42186,N_40362,N_40261);
or U42187 (N_42187,N_40170,N_40657);
xor U42188 (N_42188,N_41261,N_40627);
nand U42189 (N_42189,N_41530,N_40250);
or U42190 (N_42190,N_41352,N_41284);
xnor U42191 (N_42191,N_40942,N_40477);
xor U42192 (N_42192,N_41032,N_41967);
nand U42193 (N_42193,N_41666,N_41603);
and U42194 (N_42194,N_40851,N_41595);
xnor U42195 (N_42195,N_41097,N_41829);
or U42196 (N_42196,N_40168,N_40621);
nand U42197 (N_42197,N_40101,N_41840);
or U42198 (N_42198,N_40343,N_41254);
nor U42199 (N_42199,N_41466,N_41920);
xor U42200 (N_42200,N_40023,N_40843);
or U42201 (N_42201,N_40103,N_41857);
and U42202 (N_42202,N_41016,N_41854);
xnor U42203 (N_42203,N_40673,N_40685);
nor U42204 (N_42204,N_41125,N_40983);
nand U42205 (N_42205,N_40082,N_40548);
nor U42206 (N_42206,N_41998,N_41924);
or U42207 (N_42207,N_41392,N_41365);
or U42208 (N_42208,N_40739,N_41307);
xnor U42209 (N_42209,N_41262,N_40547);
nand U42210 (N_42210,N_40115,N_40902);
and U42211 (N_42211,N_40460,N_40142);
nor U42212 (N_42212,N_40785,N_40539);
nand U42213 (N_42213,N_41148,N_41539);
and U42214 (N_42214,N_41227,N_41348);
and U42215 (N_42215,N_41098,N_41429);
nor U42216 (N_42216,N_41131,N_40639);
xnor U42217 (N_42217,N_41372,N_41009);
and U42218 (N_42218,N_40233,N_40607);
xnor U42219 (N_42219,N_40662,N_40429);
and U42220 (N_42220,N_40417,N_41956);
or U42221 (N_42221,N_41548,N_40971);
or U42222 (N_42222,N_41496,N_41515);
nand U42223 (N_42223,N_41176,N_41043);
xnor U42224 (N_42224,N_40977,N_40558);
nand U42225 (N_42225,N_41256,N_40510);
and U42226 (N_42226,N_40073,N_41536);
xnor U42227 (N_42227,N_41371,N_41670);
nand U42228 (N_42228,N_41899,N_41837);
and U42229 (N_42229,N_41553,N_40113);
xnor U42230 (N_42230,N_40248,N_41620);
and U42231 (N_42231,N_41965,N_41529);
nand U42232 (N_42232,N_41059,N_40861);
and U42233 (N_42233,N_41086,N_40346);
nor U42234 (N_42234,N_41797,N_41035);
nand U42235 (N_42235,N_41119,N_40829);
nand U42236 (N_42236,N_41373,N_40118);
or U42237 (N_42237,N_40674,N_40680);
nor U42238 (N_42238,N_40863,N_41492);
xor U42239 (N_42239,N_40918,N_41014);
and U42240 (N_42240,N_40181,N_40859);
and U42241 (N_42241,N_41981,N_41445);
or U42242 (N_42242,N_40823,N_41090);
nor U42243 (N_42243,N_40265,N_40092);
nand U42244 (N_42244,N_40271,N_41675);
or U42245 (N_42245,N_41178,N_40967);
and U42246 (N_42246,N_40232,N_40922);
xnor U42247 (N_42247,N_41653,N_40879);
xnor U42248 (N_42248,N_40523,N_40426);
nand U42249 (N_42249,N_41946,N_40838);
or U42250 (N_42250,N_40945,N_40744);
and U42251 (N_42251,N_41354,N_41624);
nand U42252 (N_42252,N_41494,N_41419);
and U42253 (N_42253,N_40784,N_40570);
or U42254 (N_42254,N_40997,N_40575);
xnor U42255 (N_42255,N_41674,N_40675);
nand U42256 (N_42256,N_41745,N_40349);
or U42257 (N_42257,N_41255,N_41351);
and U42258 (N_42258,N_40297,N_41509);
nand U42259 (N_42259,N_40303,N_40226);
or U42260 (N_42260,N_41685,N_40212);
and U42261 (N_42261,N_40200,N_40881);
xor U42262 (N_42262,N_41531,N_41217);
and U42263 (N_42263,N_40379,N_41400);
xnor U42264 (N_42264,N_41805,N_40004);
or U42265 (N_42265,N_40506,N_40892);
or U42266 (N_42266,N_40499,N_40230);
or U42267 (N_42267,N_41816,N_41775);
or U42268 (N_42268,N_41182,N_41294);
nand U42269 (N_42269,N_40436,N_41765);
or U42270 (N_42270,N_41538,N_40020);
xor U42271 (N_42271,N_40108,N_41010);
or U42272 (N_42272,N_40210,N_41421);
and U42273 (N_42273,N_41944,N_40315);
nor U42274 (N_42274,N_41980,N_40209);
xor U42275 (N_42275,N_41069,N_41411);
and U42276 (N_42276,N_40857,N_40318);
and U42277 (N_42277,N_40138,N_40217);
and U42278 (N_42278,N_41174,N_40832);
nand U42279 (N_42279,N_40386,N_41570);
or U42280 (N_42280,N_40810,N_40786);
nor U42281 (N_42281,N_41583,N_40481);
nor U42282 (N_42282,N_41146,N_41313);
or U42283 (N_42283,N_40228,N_41343);
xor U42284 (N_42284,N_41345,N_41037);
nand U42285 (N_42285,N_41597,N_40062);
and U42286 (N_42286,N_41406,N_40366);
and U42287 (N_42287,N_40624,N_40442);
xnor U42288 (N_42288,N_40957,N_40201);
xnor U42289 (N_42289,N_41769,N_40058);
and U42290 (N_42290,N_40036,N_41051);
and U42291 (N_42291,N_41549,N_41825);
and U42292 (N_42292,N_41642,N_40393);
nor U42293 (N_42293,N_41463,N_40352);
xor U42294 (N_42294,N_41617,N_41449);
or U42295 (N_42295,N_41964,N_41555);
nand U42296 (N_42296,N_41389,N_41007);
or U42297 (N_42297,N_41732,N_40294);
nand U42298 (N_42298,N_40797,N_40220);
xor U42299 (N_42299,N_41606,N_41136);
nand U42300 (N_42300,N_41593,N_40737);
nand U42301 (N_42301,N_41143,N_41391);
xor U42302 (N_42302,N_41018,N_40024);
and U42303 (N_42303,N_40447,N_40527);
nand U42304 (N_42304,N_40951,N_40495);
and U42305 (N_42305,N_41039,N_41288);
nand U42306 (N_42306,N_40486,N_41853);
xor U42307 (N_42307,N_41520,N_41228);
and U42308 (N_42308,N_41063,N_41773);
or U42309 (N_42309,N_40411,N_41635);
nor U42310 (N_42310,N_40291,N_41211);
nor U42311 (N_42311,N_40144,N_41071);
and U42312 (N_42312,N_41826,N_41616);
or U42313 (N_42313,N_40788,N_41094);
and U42314 (N_42314,N_40671,N_41152);
nor U42315 (N_42315,N_41874,N_41167);
or U42316 (N_42316,N_40021,N_40364);
xor U42317 (N_42317,N_40790,N_41060);
and U42318 (N_42318,N_40656,N_40333);
or U42319 (N_42319,N_41560,N_40190);
nor U42320 (N_42320,N_41955,N_41691);
nor U42321 (N_42321,N_40347,N_41689);
and U42322 (N_42322,N_41717,N_41339);
nand U42323 (N_42323,N_40160,N_40264);
nor U42324 (N_42324,N_40988,N_41360);
xnor U42325 (N_42325,N_41065,N_40095);
xor U42326 (N_42326,N_41710,N_40877);
or U42327 (N_42327,N_41096,N_41545);
or U42328 (N_42328,N_40776,N_40668);
or U42329 (N_42329,N_40239,N_41526);
xor U42330 (N_42330,N_41164,N_40974);
and U42331 (N_42331,N_41551,N_40728);
and U42332 (N_42332,N_40850,N_41382);
xor U42333 (N_42333,N_41692,N_41428);
nor U42334 (N_42334,N_40948,N_40344);
nor U42335 (N_42335,N_40868,N_41370);
nand U42336 (N_42336,N_40031,N_41013);
xor U42337 (N_42337,N_41966,N_40820);
xor U42338 (N_42338,N_41770,N_40377);
or U42339 (N_42339,N_41353,N_40848);
or U42340 (N_42340,N_40584,N_40695);
nor U42341 (N_42341,N_41586,N_41344);
or U42342 (N_42342,N_40270,N_41394);
nor U42343 (N_42343,N_41661,N_41974);
or U42344 (N_42344,N_41954,N_41075);
nor U42345 (N_42345,N_40669,N_41306);
and U42346 (N_42346,N_40269,N_41171);
or U42347 (N_42347,N_40310,N_41973);
nor U42348 (N_42348,N_40525,N_41235);
nand U42349 (N_42349,N_41786,N_41547);
xnor U42350 (N_42350,N_40099,N_41599);
xor U42351 (N_42351,N_40418,N_41324);
or U42352 (N_42352,N_41552,N_40106);
xnor U42353 (N_42353,N_41056,N_40367);
nor U42354 (N_42354,N_40339,N_40970);
or U42355 (N_42355,N_40086,N_40546);
and U42356 (N_42356,N_41535,N_40887);
xor U42357 (N_42357,N_40249,N_41868);
and U42358 (N_42358,N_41824,N_41395);
and U42359 (N_42359,N_41447,N_41106);
xnor U42360 (N_42360,N_41383,N_40493);
xnor U42361 (N_42361,N_41163,N_40611);
nand U42362 (N_42362,N_40596,N_40198);
nand U42363 (N_42363,N_41012,N_41623);
xor U42364 (N_42364,N_41308,N_41248);
nand U42365 (N_42365,N_40186,N_41144);
nor U42366 (N_42366,N_41633,N_41301);
or U42367 (N_42367,N_41044,N_40618);
or U42368 (N_42368,N_41519,N_40726);
or U42369 (N_42369,N_41495,N_41240);
xor U42370 (N_42370,N_40802,N_41177);
xnor U42371 (N_42371,N_40059,N_41282);
and U42372 (N_42372,N_41410,N_41356);
xnor U42373 (N_42373,N_40026,N_41150);
nor U42374 (N_42374,N_41656,N_40087);
and U42375 (N_42375,N_41237,N_41795);
and U42376 (N_42376,N_40369,N_41983);
xor U42377 (N_42377,N_40307,N_41834);
and U42378 (N_42378,N_41927,N_40497);
nor U42379 (N_42379,N_40904,N_40583);
nand U42380 (N_42380,N_40867,N_40211);
and U42381 (N_42381,N_41083,N_40704);
and U42382 (N_42382,N_41468,N_40392);
nor U42383 (N_42383,N_41165,N_41417);
nand U42384 (N_42384,N_40134,N_40402);
nand U42385 (N_42385,N_41471,N_40179);
xnor U42386 (N_42386,N_41225,N_41388);
nor U42387 (N_42387,N_40767,N_41349);
nor U42388 (N_42388,N_40008,N_41379);
xnor U42389 (N_42389,N_40777,N_40345);
and U42390 (N_42390,N_41318,N_41698);
and U42391 (N_42391,N_40162,N_41290);
xnor U42392 (N_42392,N_41913,N_40835);
or U42393 (N_42393,N_40912,N_40319);
and U42394 (N_42394,N_41149,N_40524);
nand U42395 (N_42395,N_41311,N_41484);
nor U42396 (N_42396,N_41409,N_40378);
nor U42397 (N_42397,N_40223,N_41742);
nand U42398 (N_42398,N_41172,N_40455);
nor U42399 (N_42399,N_40642,N_40245);
nand U42400 (N_42400,N_40154,N_40796);
nor U42401 (N_42401,N_41802,N_41730);
or U42402 (N_42402,N_40541,N_40808);
or U42403 (N_42403,N_40311,N_41758);
xor U42404 (N_42404,N_40979,N_40509);
and U42405 (N_42405,N_41612,N_40890);
or U42406 (N_42406,N_40374,N_40538);
and U42407 (N_42407,N_40987,N_41702);
and U42408 (N_42408,N_40462,N_40235);
or U42409 (N_42409,N_41020,N_40615);
nor U42410 (N_42410,N_41404,N_41828);
nand U42411 (N_42411,N_41334,N_41706);
and U42412 (N_42412,N_40242,N_41472);
and U42413 (N_42413,N_41465,N_40703);
xnor U42414 (N_42414,N_40171,N_41926);
or U42415 (N_42415,N_41092,N_40903);
nor U42416 (N_42416,N_41206,N_41239);
xor U42417 (N_42417,N_40930,N_41291);
xnor U42418 (N_42418,N_41648,N_40363);
and U42419 (N_42419,N_41843,N_40889);
or U42420 (N_42420,N_40017,N_41140);
xnor U42421 (N_42421,N_40111,N_40238);
or U42422 (N_42422,N_41576,N_40670);
nor U42423 (N_42423,N_40076,N_40722);
and U42424 (N_42424,N_41187,N_40964);
nor U42425 (N_42425,N_40801,N_41862);
nor U42426 (N_42426,N_40185,N_40032);
and U42427 (N_42427,N_40282,N_40992);
xnor U42428 (N_42428,N_40433,N_41002);
nor U42429 (N_42429,N_40834,N_40176);
nand U42430 (N_42430,N_41590,N_40821);
nor U42431 (N_42431,N_41704,N_41701);
or U42432 (N_42432,N_40976,N_40480);
nor U42433 (N_42433,N_41249,N_41487);
or U42434 (N_42434,N_41736,N_40070);
or U42435 (N_42435,N_41401,N_41310);
or U42436 (N_42436,N_40110,N_41566);
nand U42437 (N_42437,N_40043,N_41870);
nand U42438 (N_42438,N_40637,N_40425);
nor U42439 (N_42439,N_41234,N_40679);
xor U42440 (N_42440,N_40530,N_40888);
nor U42441 (N_42441,N_41567,N_41994);
and U42442 (N_42442,N_40394,N_41041);
or U42443 (N_42443,N_41491,N_41506);
and U42444 (N_42444,N_41376,N_41355);
or U42445 (N_42445,N_41333,N_40628);
and U42446 (N_42446,N_40130,N_40813);
nand U42447 (N_42447,N_41074,N_40629);
or U42448 (N_42448,N_40243,N_41575);
or U42449 (N_42449,N_41099,N_41393);
or U42450 (N_42450,N_41145,N_41269);
xor U42451 (N_42451,N_40806,N_41154);
nor U42452 (N_42452,N_40906,N_40914);
or U42453 (N_42453,N_40451,N_41921);
nand U42454 (N_42454,N_41836,N_40751);
and U42455 (N_42455,N_40370,N_40898);
nor U42456 (N_42456,N_41375,N_41902);
or U42457 (N_42457,N_41273,N_41918);
or U42458 (N_42458,N_40093,N_40996);
or U42459 (N_42459,N_40100,N_41752);
nor U42460 (N_42460,N_40022,N_41522);
xor U42461 (N_42461,N_41686,N_41889);
nand U42462 (N_42462,N_41505,N_41188);
xor U42463 (N_42463,N_41433,N_41546);
and U42464 (N_42464,N_41672,N_40614);
and U42465 (N_42465,N_40468,N_41367);
and U42466 (N_42466,N_41170,N_40193);
nor U42467 (N_42467,N_40632,N_41080);
and U42468 (N_42468,N_40692,N_40816);
nor U42469 (N_42469,N_41541,N_40153);
xor U42470 (N_42470,N_41631,N_40456);
nor U42471 (N_42471,N_41731,N_41872);
xnor U42472 (N_42472,N_41794,N_40478);
nor U42473 (N_42473,N_41160,N_40954);
xor U42474 (N_42474,N_41808,N_40445);
xnor U42475 (N_42475,N_40577,N_41727);
nand U42476 (N_42476,N_41912,N_41251);
xnor U42477 (N_42477,N_40192,N_41637);
nor U42478 (N_42478,N_41993,N_41439);
xor U42479 (N_42479,N_40085,N_40630);
and U42480 (N_42480,N_41161,N_40330);
and U42481 (N_42481,N_41321,N_41011);
nand U42482 (N_42482,N_41332,N_40862);
nand U42483 (N_42483,N_41109,N_40383);
or U42484 (N_42484,N_40756,N_40705);
nand U42485 (N_42485,N_40897,N_41067);
and U42486 (N_42486,N_41205,N_41923);
nor U42487 (N_42487,N_41919,N_41469);
and U42488 (N_42488,N_40331,N_40327);
nand U42489 (N_42489,N_40443,N_40873);
xor U42490 (N_42490,N_41733,N_40891);
nor U42491 (N_42491,N_41987,N_40222);
or U42492 (N_42492,N_41347,N_40537);
nand U42493 (N_42493,N_40531,N_41415);
xor U42494 (N_42494,N_41500,N_40295);
nand U42495 (N_42495,N_40077,N_40740);
nand U42496 (N_42496,N_40965,N_41992);
and U42497 (N_42497,N_40567,N_41982);
nand U42498 (N_42498,N_41336,N_41342);
nor U42499 (N_42499,N_41508,N_40518);
and U42500 (N_42500,N_41481,N_40854);
nor U42501 (N_42501,N_40079,N_40483);
nor U42502 (N_42502,N_40610,N_40663);
or U42503 (N_42503,N_40397,N_41122);
nand U42504 (N_42504,N_41079,N_40831);
xor U42505 (N_42505,N_41916,N_40773);
nand U42506 (N_42506,N_41123,N_41724);
or U42507 (N_42507,N_40312,N_40782);
and U42508 (N_42508,N_40473,N_40858);
xnor U42509 (N_42509,N_41278,N_41952);
nand U42510 (N_42510,N_40508,N_40588);
nand U42511 (N_42511,N_40494,N_40501);
and U42512 (N_42512,N_41104,N_40304);
nor U42513 (N_42513,N_41614,N_40492);
or U42514 (N_42514,N_41799,N_41779);
xnor U42515 (N_42515,N_41751,N_41168);
nand U42516 (N_42516,N_40602,N_40593);
xnor U42517 (N_42517,N_41726,N_41435);
nand U42518 (N_42518,N_40229,N_41314);
xnor U42519 (N_42519,N_40384,N_40189);
nor U42520 (N_42520,N_41436,N_41875);
nand U42521 (N_42521,N_41441,N_40117);
xnor U42522 (N_42522,N_40078,N_40780);
and U42523 (N_42523,N_41668,N_40140);
and U42524 (N_42524,N_40470,N_41113);
xnor U42525 (N_42525,N_41482,N_41420);
nor U42526 (N_42526,N_41784,N_41602);
and U42527 (N_42527,N_40416,N_41790);
or U42528 (N_42528,N_41556,N_40465);
and U42529 (N_42529,N_40399,N_41374);
xnor U42530 (N_42530,N_41850,N_41464);
nand U42531 (N_42531,N_41709,N_41721);
and U42532 (N_42532,N_41476,N_41377);
nand U42533 (N_42533,N_40091,N_41268);
xnor U42534 (N_42534,N_40758,N_41716);
and U42535 (N_42535,N_41673,N_40694);
nand U42536 (N_42536,N_41252,N_41737);
nand U42537 (N_42537,N_41437,N_41680);
nor U42538 (N_42538,N_41423,N_40913);
nand U42539 (N_42539,N_41309,N_40296);
and U42540 (N_42540,N_41524,N_40872);
xor U42541 (N_42541,N_41153,N_41510);
and U42542 (N_42542,N_40544,N_40761);
or U42543 (N_42543,N_40943,N_41578);
xnor U42544 (N_42544,N_41788,N_40035);
nor U42545 (N_42545,N_40254,N_40299);
or U42546 (N_42546,N_41562,N_40044);
and U42547 (N_42547,N_41319,N_41322);
and U42548 (N_42548,N_40221,N_41819);
xnor U42549 (N_42549,N_41247,N_40731);
or U42550 (N_42550,N_41118,N_41213);
and U42551 (N_42551,N_40214,N_41128);
or U42552 (N_42552,N_40284,N_40459);
and U42553 (N_42553,N_40749,N_41831);
and U42554 (N_42554,N_40847,N_40907);
xnor U42555 (N_42555,N_41222,N_41337);
xnor U42556 (N_42556,N_40263,N_41754);
and U42557 (N_42557,N_40947,N_40457);
nor U42558 (N_42558,N_40754,N_40911);
nand U42559 (N_42559,N_41147,N_41335);
nor U42560 (N_42560,N_40453,N_41632);
xor U42561 (N_42561,N_41999,N_41201);
and U42562 (N_42562,N_40090,N_40590);
xor U42563 (N_42563,N_41897,N_40827);
nor U42564 (N_42564,N_41166,N_41682);
or U42565 (N_42565,N_40380,N_40645);
or U42566 (N_42566,N_40900,N_41914);
nand U42567 (N_42567,N_41729,N_40309);
nor U42568 (N_42568,N_41180,N_41605);
and U42569 (N_42569,N_41898,N_41589);
nand U42570 (N_42570,N_41232,N_40050);
and U42571 (N_42571,N_41792,N_40735);
xor U42572 (N_42572,N_40030,N_41712);
xnor U42573 (N_42573,N_40382,N_40587);
nand U42574 (N_42574,N_40063,N_40746);
nand U42575 (N_42575,N_40573,N_40865);
nor U42576 (N_42576,N_40552,N_40325);
nor U42577 (N_42577,N_40219,N_40634);
and U42578 (N_42578,N_40648,N_40375);
and U42579 (N_42579,N_40081,N_41568);
xnor U42580 (N_42580,N_41749,N_40643);
nand U42581 (N_42581,N_40496,N_40141);
or U42582 (N_42582,N_41647,N_41625);
nor U42583 (N_42583,N_41049,N_41577);
or U42584 (N_42584,N_41001,N_41274);
and U42585 (N_42585,N_40540,N_41380);
xor U42586 (N_42586,N_40215,N_41438);
xnor U42587 (N_42587,N_41804,N_41713);
or U42588 (N_42588,N_41942,N_41271);
or U42589 (N_42589,N_41296,N_41774);
and U42590 (N_42590,N_41649,N_40388);
or U42591 (N_42591,N_41848,N_41791);
xnor U42592 (N_42592,N_41719,N_41579);
or U42593 (N_42593,N_40234,N_41101);
or U42594 (N_42594,N_40817,N_41947);
or U42595 (N_42595,N_41735,N_41861);
xor U42596 (N_42596,N_40990,N_40870);
and U42597 (N_42597,N_40368,N_40395);
or U42598 (N_42598,N_41896,N_40001);
nor U42599 (N_42599,N_40006,N_40438);
nand U42600 (N_42600,N_40789,N_40301);
nand U42601 (N_42601,N_41493,N_40145);
nand U42602 (N_42602,N_40884,N_40617);
nand U42603 (N_42603,N_41905,N_41317);
nor U42604 (N_42604,N_40165,N_40316);
nand U42605 (N_42605,N_41068,N_40335);
or U42606 (N_42606,N_40060,N_41460);
or U42607 (N_42607,N_41948,N_40439);
nor U42608 (N_42608,N_40505,N_41703);
nor U42609 (N_42609,N_40641,N_40794);
nand U42610 (N_42610,N_40348,N_41230);
nand U42611 (N_42611,N_40197,N_41006);
nor U42612 (N_42612,N_40616,N_40905);
or U42613 (N_42613,N_40532,N_41986);
nand U42614 (N_42614,N_41621,N_41141);
or U42615 (N_42615,N_41767,N_40195);
nor U42616 (N_42616,N_40102,N_41813);
nand U42617 (N_42617,N_41760,N_41771);
nor U42618 (N_42618,N_41960,N_40409);
or U42619 (N_42619,N_41190,N_40514);
nor U42620 (N_42620,N_41093,N_40683);
and U42621 (N_42621,N_41470,N_41903);
xnor U42622 (N_42622,N_41243,N_40415);
nand U42623 (N_42623,N_41513,N_40515);
xor U42624 (N_42624,N_40812,N_41350);
and U42625 (N_42625,N_40039,N_41820);
xor U42626 (N_42626,N_40218,N_40916);
or U42627 (N_42627,N_40267,N_41479);
nor U42628 (N_42628,N_40565,N_41272);
xor U42629 (N_42629,N_40283,N_41569);
xnor U42630 (N_42630,N_40991,N_41978);
nand U42631 (N_42631,N_41938,N_40048);
nand U42632 (N_42632,N_41780,N_41215);
and U42633 (N_42633,N_40644,N_40522);
xnor U42634 (N_42634,N_41664,N_40999);
nand U42635 (N_42635,N_41512,N_40855);
or U42636 (N_42636,N_41329,N_40372);
and U42637 (N_42637,N_40000,N_41766);
xnor U42638 (N_42638,N_41105,N_41598);
xnor U42639 (N_42639,N_40216,N_40589);
nand U42640 (N_42640,N_41718,N_41138);
nor U42641 (N_42641,N_40337,N_40960);
xor U42642 (N_42642,N_40246,N_41156);
xor U42643 (N_42643,N_41638,N_41369);
xnor U42644 (N_42644,N_40046,N_40428);
nand U42645 (N_42645,N_41646,N_41359);
xor U42646 (N_42646,N_41384,N_41815);
nand U42647 (N_42647,N_40503,N_40871);
nor U42648 (N_42648,N_40422,N_40716);
and U42649 (N_42649,N_41413,N_41162);
nor U42650 (N_42650,N_41565,N_40123);
and U42651 (N_42651,N_40720,N_40279);
and U42652 (N_42652,N_41867,N_40194);
nand U42653 (N_42653,N_40159,N_41110);
xor U42654 (N_42654,N_40528,N_40033);
or U42655 (N_42655,N_41236,N_40203);
nand U42656 (N_42656,N_40856,N_41796);
xor U42657 (N_42657,N_40498,N_40896);
nor U42658 (N_42658,N_41455,N_41812);
and U42659 (N_42659,N_40317,N_41939);
nand U42660 (N_42660,N_41935,N_40088);
and U42661 (N_42661,N_41265,N_41489);
and U42662 (N_42662,N_41111,N_41639);
or U42663 (N_42663,N_41521,N_41115);
nor U42664 (N_42664,N_41622,N_41725);
or U42665 (N_42665,N_41192,N_40052);
nor U42666 (N_42666,N_41910,N_41814);
xnor U42667 (N_42667,N_41473,N_40067);
nand U42668 (N_42668,N_40866,N_41442);
nand U42669 (N_42669,N_41312,N_41293);
nor U42670 (N_42670,N_41892,N_41501);
nor U42671 (N_42671,N_40178,N_40640);
and U42672 (N_42672,N_40603,N_41112);
nor U42673 (N_42673,N_40886,N_41550);
nor U42674 (N_42674,N_41859,N_41026);
or U42675 (N_42675,N_40157,N_40292);
nand U42676 (N_42676,N_41126,N_40574);
nor U42677 (N_42677,N_40939,N_40389);
and U42678 (N_42678,N_41316,N_41720);
and U42679 (N_42679,N_41743,N_40710);
or U42680 (N_42680,N_40846,N_40686);
nor U42681 (N_42681,N_40612,N_41017);
and U42682 (N_42682,N_40818,N_41915);
nand U42683 (N_42683,N_41961,N_41640);
xor U42684 (N_42684,N_41688,N_40419);
or U42685 (N_42685,N_40717,N_41403);
nand U42686 (N_42686,N_41502,N_40927);
xor U42687 (N_42687,N_40289,N_40148);
xor U42688 (N_42688,N_40741,N_40276);
or U42689 (N_42689,N_40454,N_40340);
nand U42690 (N_42690,N_41990,N_40237);
xor U42691 (N_42691,N_40013,N_40056);
or U42692 (N_42692,N_40391,N_41798);
xor U42693 (N_42693,N_41931,N_40766);
nor U42694 (N_42694,N_41229,N_41629);
nor U42695 (N_42695,N_40488,N_40350);
nor U42696 (N_42696,N_40598,N_40915);
nand U42697 (N_42697,N_40187,N_40620);
and U42698 (N_42698,N_40733,N_40041);
nor U42699 (N_42699,N_41042,N_41679);
or U42700 (N_42700,N_40878,N_41028);
nor U42701 (N_42701,N_41134,N_40273);
nand U42702 (N_42702,N_40191,N_41019);
and U42703 (N_42703,N_41456,N_40244);
nor U42704 (N_42704,N_40479,N_41408);
and U42705 (N_42705,N_40147,N_40571);
nand U42706 (N_42706,N_41158,N_41207);
or U42707 (N_42707,N_41204,N_40654);
nor U42708 (N_42708,N_41591,N_40529);
and U42709 (N_42709,N_41477,N_41723);
nand U42710 (N_42710,N_41497,N_41133);
and U42711 (N_42711,N_41596,N_41062);
nand U42712 (N_42712,N_40255,N_40652);
xor U42713 (N_42713,N_40586,N_41326);
xor U42714 (N_42714,N_40893,N_40109);
or U42715 (N_42715,N_40601,N_40083);
nor U42716 (N_42716,N_41855,N_40458);
or U42717 (N_42717,N_41387,N_40277);
or U42718 (N_42718,N_41627,N_40768);
or U42719 (N_42719,N_40949,N_41734);
nor U42720 (N_42720,N_40747,N_40681);
xor U42721 (N_42721,N_40581,N_40631);
xor U42722 (N_42722,N_41238,N_40328);
xnor U42723 (N_42723,N_40566,N_41669);
nand U42724 (N_42724,N_41906,N_40027);
and U42725 (N_42725,N_41655,N_40326);
or U42726 (N_42726,N_40594,N_40809);
or U42727 (N_42727,N_41928,N_40771);
nand U42728 (N_42728,N_41917,N_40288);
and U42729 (N_42729,N_40697,N_40196);
nor U42730 (N_42730,N_41478,N_40446);
xor U42731 (N_42731,N_41003,N_41564);
nor U42732 (N_42732,N_40713,N_40984);
nand U42733 (N_42733,N_40259,N_40882);
nand U42734 (N_42734,N_41185,N_41048);
nand U42735 (N_42735,N_40452,N_41841);
and U42736 (N_42736,N_40764,N_41748);
and U42737 (N_42737,N_40061,N_40750);
nor U42738 (N_42738,N_41611,N_40400);
or U42739 (N_42739,N_41091,N_40253);
and U42740 (N_42740,N_41108,N_40139);
nor U42741 (N_42741,N_40647,N_41378);
xor U42742 (N_42742,N_40094,N_41833);
nand U42743 (N_42743,N_40003,N_40952);
xor U42744 (N_42744,N_40533,N_41959);
or U42745 (N_42745,N_40696,N_41801);
nor U42746 (N_42746,N_41179,N_41587);
xor U42747 (N_42747,N_40161,N_41949);
or U42748 (N_42748,N_41040,N_40306);
or U42749 (N_42749,N_41604,N_41100);
or U42750 (N_42750,N_40653,N_41454);
or U42751 (N_42751,N_41214,N_40635);
nand U42752 (N_42752,N_40208,N_41459);
and U42753 (N_42753,N_40015,N_40487);
and U42754 (N_42754,N_41907,N_40792);
xor U42755 (N_42755,N_41705,N_40719);
or U42756 (N_42756,N_40332,N_40894);
or U42757 (N_42757,N_40414,N_41807);
nand U42758 (N_42758,N_40687,N_40421);
and U42759 (N_42759,N_41839,N_40923);
xnor U42760 (N_42760,N_40989,N_41781);
nand U42761 (N_42761,N_40924,N_41315);
nor U42762 (N_42762,N_41645,N_41873);
xnor U42763 (N_42763,N_40241,N_40959);
xor U42764 (N_42764,N_40715,N_41287);
and U42765 (N_42765,N_41654,N_40293);
and U42766 (N_42766,N_40963,N_40298);
nor U42767 (N_42767,N_41280,N_40068);
xor U42768 (N_42768,N_41778,N_41289);
nor U42769 (N_42769,N_40763,N_40373);
and U42770 (N_42770,N_41517,N_40396);
and U42771 (N_42771,N_41830,N_40841);
nand U42772 (N_42772,N_41842,N_41076);
nand U42773 (N_42773,N_41015,N_41338);
and U42774 (N_42774,N_41582,N_40795);
xnor U42775 (N_42775,N_40371,N_40359);
xor U42776 (N_42776,N_40323,N_41061);
nor U42777 (N_42777,N_41652,N_40137);
nor U42778 (N_42778,N_41399,N_41050);
xnor U42779 (N_42779,N_40543,N_40787);
xnor U42780 (N_42780,N_40336,N_40320);
xor U42781 (N_42781,N_41847,N_40278);
and U42782 (N_42782,N_40520,N_41764);
nor U42783 (N_42783,N_41803,N_41932);
or U42784 (N_42784,N_41811,N_41523);
nand U42785 (N_42785,N_41490,N_40164);
or U42786 (N_42786,N_40633,N_41021);
nor U42787 (N_42787,N_41151,N_41787);
or U42788 (N_42788,N_41818,N_41286);
or U42789 (N_42789,N_41763,N_40919);
or U42790 (N_42790,N_41904,N_40791);
nand U42791 (N_42791,N_41000,N_40025);
and U42792 (N_42792,N_41883,N_41544);
or U42793 (N_42793,N_40285,N_41525);
or U42794 (N_42794,N_40936,N_41260);
xor U42795 (N_42795,N_41738,N_41046);
or U42796 (N_42796,N_40268,N_40430);
nor U42797 (N_42797,N_41969,N_41558);
nand U42798 (N_42798,N_41607,N_40180);
xnor U42799 (N_42799,N_40080,N_41601);
or U42800 (N_42800,N_40484,N_40205);
or U42801 (N_42801,N_40476,N_41107);
nand U42802 (N_42802,N_41299,N_41340);
xnor U42803 (N_42803,N_41728,N_41103);
nor U42804 (N_42804,N_40962,N_40441);
nand U42805 (N_42805,N_40664,N_41250);
or U42806 (N_42806,N_40727,N_40693);
nor U42807 (N_42807,N_40011,N_41127);
and U42808 (N_42808,N_40932,N_41885);
nand U42809 (N_42809,N_41216,N_40623);
and U42810 (N_42810,N_40800,N_41285);
nor U42811 (N_42811,N_41323,N_41070);
and U42812 (N_42812,N_41263,N_40721);
xor U42813 (N_42813,N_40753,N_41962);
nand U42814 (N_42814,N_40860,N_41863);
nor U42815 (N_42815,N_40845,N_41300);
nand U42816 (N_42816,N_41114,N_41084);
or U42817 (N_42817,N_40946,N_41951);
and U42818 (N_42818,N_41711,N_41241);
nor U42819 (N_42819,N_40935,N_41528);
and U42820 (N_42820,N_41412,N_40568);
or U42821 (N_42821,N_40576,N_40407);
or U42822 (N_42822,N_41561,N_40225);
or U42823 (N_42823,N_41363,N_41129);
nor U42824 (N_42824,N_40736,N_41004);
or U42825 (N_42825,N_40650,N_41684);
nand U42826 (N_42826,N_40051,N_40361);
nand U42827 (N_42827,N_40146,N_41877);
or U42828 (N_42828,N_40536,N_40463);
xnor U42829 (N_42829,N_41159,N_41678);
and U42830 (N_42830,N_41135,N_40252);
or U42831 (N_42831,N_40356,N_40057);
xor U42832 (N_42832,N_41142,N_41358);
nand U42833 (N_42833,N_40262,N_41186);
nand U42834 (N_42834,N_40572,N_40135);
or U42835 (N_42835,N_40853,N_40128);
xor U42836 (N_42836,N_40910,N_40308);
nor U42837 (N_42837,N_41864,N_41881);
nand U42838 (N_42838,N_41397,N_41511);
or U42839 (N_42839,N_41559,N_40286);
nand U42840 (N_42840,N_41600,N_40626);
nor U42841 (N_42841,N_41608,N_41124);
and U42842 (N_42842,N_40266,N_40365);
or U42843 (N_42843,N_41641,N_41033);
nor U42844 (N_42844,N_41053,N_41933);
xnor U42845 (N_42845,N_41087,N_41175);
nand U42846 (N_42846,N_40151,N_41699);
or U42847 (N_42847,N_40334,N_41776);
nand U42848 (N_42848,N_40658,N_41543);
and U42849 (N_42849,N_40028,N_41958);
nor U42850 (N_42850,N_41922,N_40597);
nor U42851 (N_42851,N_41953,N_40698);
nor U42852 (N_42852,N_40482,N_41878);
nor U42853 (N_42853,N_40660,N_40551);
and U42854 (N_42854,N_40467,N_41045);
nand U42855 (N_42855,N_41304,N_40839);
nor U42856 (N_42856,N_40448,N_40089);
nand U42857 (N_42857,N_40423,N_41943);
nand U42858 (N_42858,N_41592,N_41891);
xnor U42859 (N_42859,N_40403,N_41634);
nor U42860 (N_42860,N_40517,N_40557);
xor U42861 (N_42861,N_41095,N_40852);
or U42862 (N_42862,N_41744,N_40569);
and U42863 (N_42863,N_41793,N_40257);
and U42864 (N_42864,N_40387,N_41504);
xor U42865 (N_42865,N_41183,N_40119);
xor U42866 (N_42866,N_40491,N_41984);
xor U42867 (N_42867,N_41707,N_41930);
nor U42868 (N_42868,N_41223,N_40950);
or U42869 (N_42869,N_41618,N_40826);
xor U42870 (N_42870,N_41297,N_40227);
xnor U42871 (N_42871,N_40507,N_40606);
and U42872 (N_42872,N_40314,N_41991);
nor U42873 (N_42873,N_40555,N_40819);
nand U42874 (N_42874,N_40955,N_40313);
or U42875 (N_42875,N_40124,N_40798);
or U42876 (N_42876,N_40112,N_40121);
or U42877 (N_42877,N_40132,N_41259);
xor U42878 (N_42878,N_41925,N_41443);
or U42879 (N_42879,N_41328,N_41196);
and U42880 (N_42880,N_41453,N_40149);
nor U42881 (N_42881,N_40743,N_40702);
nor U42882 (N_42882,N_40272,N_41995);
or U42883 (N_42883,N_40172,N_40405);
nor U42884 (N_42884,N_40714,N_40049);
and U42885 (N_42885,N_40521,N_40978);
and U42886 (N_42886,N_40007,N_40107);
xnor U42887 (N_42887,N_41989,N_41740);
nor U42888 (N_42888,N_40690,N_41078);
nor U42889 (N_42889,N_40485,N_40973);
nand U42890 (N_42890,N_41034,N_41024);
or U42891 (N_42891,N_41697,N_41772);
xnor U42892 (N_42892,N_40609,N_40998);
and U42893 (N_42893,N_40183,N_40604);
or U42894 (N_42894,N_41643,N_40969);
nor U42895 (N_42895,N_40880,N_40338);
and U42896 (N_42896,N_40968,N_40899);
and U42897 (N_42897,N_40833,N_40173);
nand U42898 (N_42898,N_40814,N_41458);
or U42899 (N_42899,N_40351,N_40665);
nand U42900 (N_42900,N_40037,N_41609);
xor U42901 (N_42901,N_41860,N_40885);
nor U42902 (N_42902,N_41264,N_40275);
nor U42903 (N_42903,N_40666,N_40994);
xnor U42904 (N_42904,N_41221,N_40513);
or U42905 (N_42905,N_41908,N_41116);
nor U42906 (N_42906,N_41636,N_41120);
nor U42907 (N_42907,N_41886,N_41970);
and U42908 (N_42908,N_40437,N_40689);
nor U42909 (N_42909,N_40781,N_40706);
or U42910 (N_42910,N_40542,N_41715);
xor U42911 (N_42911,N_41402,N_41895);
or U42912 (N_42912,N_40053,N_40152);
nor U42913 (N_42913,N_40054,N_40412);
nand U42914 (N_42914,N_41173,N_41800);
nor U42915 (N_42915,N_41197,N_41785);
nand U42916 (N_42916,N_41851,N_41761);
xnor U42917 (N_42917,N_40908,N_40096);
and U42918 (N_42918,N_40251,N_40700);
and U42919 (N_42919,N_40055,N_41532);
nand U42920 (N_42920,N_40636,N_40016);
or U42921 (N_42921,N_41488,N_41444);
and U42922 (N_42922,N_41432,N_41610);
nand U42923 (N_42923,N_41615,N_40828);
and U42924 (N_42924,N_40811,N_41584);
or U42925 (N_42925,N_41572,N_41474);
or U42926 (N_42926,N_40358,N_40613);
xor U42927 (N_42927,N_40131,N_41357);
nand U42928 (N_42928,N_40864,N_41747);
and U42929 (N_42929,N_40591,N_41193);
and U42930 (N_42930,N_40424,N_41231);
or U42931 (N_42931,N_40938,N_40231);
and U42932 (N_42932,N_40956,N_41650);
nand U42933 (N_42933,N_41305,N_41132);
and U42934 (N_42934,N_40098,N_41082);
nor U42935 (N_42935,N_41366,N_41879);
nand U42936 (N_42936,N_40012,N_40775);
nand U42937 (N_42937,N_40290,N_41756);
xor U42938 (N_42938,N_40075,N_41195);
or U42939 (N_42939,N_41424,N_41856);
nand U42940 (N_42940,N_40413,N_40432);
nor U42941 (N_42941,N_40449,N_40844);
or U42942 (N_42942,N_41431,N_41533);
or U42943 (N_42943,N_40592,N_41882);
xor U42944 (N_42944,N_40672,N_41865);
and U42945 (N_42945,N_41900,N_41157);
and U42946 (N_42946,N_41303,N_40595);
nand U42947 (N_42947,N_40280,N_41659);
or U42948 (N_42948,N_41057,N_40585);
and U42949 (N_42949,N_40840,N_41137);
xor U42950 (N_42950,N_40982,N_41762);
nand U42951 (N_42951,N_41242,N_40993);
or U42952 (N_42952,N_41220,N_41219);
nor U42953 (N_42953,N_40175,N_41480);
nor U42954 (N_42954,N_41233,N_41827);
xor U42955 (N_42955,N_40600,N_41130);
nand U42956 (N_42956,N_41628,N_40708);
and U42957 (N_42957,N_40357,N_41957);
nor U42958 (N_42958,N_40434,N_41693);
nor U42959 (N_42959,N_40564,N_41027);
and U42960 (N_42960,N_40822,N_41976);
or U42961 (N_42961,N_40769,N_40322);
nand U42962 (N_42962,N_40177,N_40804);
nor U42963 (N_42963,N_40014,N_40762);
or U42964 (N_42964,N_40204,N_40167);
or U42965 (N_42965,N_40760,N_40475);
xor U42966 (N_42966,N_41594,N_40535);
or U42967 (N_42967,N_40406,N_41266);
or U42968 (N_42968,N_40408,N_40917);
or U42969 (N_42969,N_41571,N_40353);
and U42970 (N_42970,N_40961,N_40926);
nor U42971 (N_42971,N_40931,N_40002);
nor U42972 (N_42972,N_40502,N_41418);
or U42973 (N_42973,N_40355,N_40559);
nand U42974 (N_42974,N_40883,N_40793);
or U42975 (N_42975,N_41613,N_41809);
or U42976 (N_42976,N_40940,N_40933);
nor U42977 (N_42977,N_41997,N_40143);
xnor U42978 (N_42978,N_41499,N_41852);
and U42979 (N_42979,N_41782,N_40511);
nor U42980 (N_42980,N_40944,N_40725);
or U42981 (N_42981,N_41937,N_40638);
nor U42982 (N_42982,N_40042,N_40302);
nand U42983 (N_42983,N_41768,N_40247);
or U42984 (N_42984,N_40563,N_41888);
nand U42985 (N_42985,N_40550,N_41212);
nand U42986 (N_42986,N_40554,N_41257);
nand U42987 (N_42987,N_40018,N_41398);
nand U42988 (N_42988,N_41746,N_41486);
nand U42989 (N_42989,N_40937,N_41085);
and U42990 (N_42990,N_40599,N_40711);
xnor U42991 (N_42991,N_40305,N_40207);
or U42992 (N_42992,N_41077,N_40150);
nor U42993 (N_42993,N_40029,N_41181);
nor U42994 (N_42994,N_40287,N_40757);
and U42995 (N_42995,N_41452,N_40321);
nand U42996 (N_42996,N_41058,N_40274);
or U42997 (N_42997,N_41588,N_41971);
and U42998 (N_42998,N_41945,N_40410);
nor U42999 (N_42999,N_41866,N_40659);
or U43000 (N_43000,N_41243,N_41101);
or U43001 (N_43001,N_41180,N_40049);
and U43002 (N_43002,N_40961,N_40188);
or U43003 (N_43003,N_41491,N_40721);
nor U43004 (N_43004,N_40767,N_41617);
and U43005 (N_43005,N_41877,N_40667);
xor U43006 (N_43006,N_41673,N_41797);
or U43007 (N_43007,N_40691,N_40903);
and U43008 (N_43008,N_40600,N_41072);
nor U43009 (N_43009,N_40204,N_41179);
xnor U43010 (N_43010,N_40359,N_40962);
nor U43011 (N_43011,N_41452,N_41286);
nand U43012 (N_43012,N_40250,N_41774);
nor U43013 (N_43013,N_40081,N_41112);
nor U43014 (N_43014,N_40302,N_40570);
and U43015 (N_43015,N_41593,N_40398);
nor U43016 (N_43016,N_40398,N_40946);
nor U43017 (N_43017,N_41177,N_41160);
and U43018 (N_43018,N_41415,N_40849);
nor U43019 (N_43019,N_40562,N_41967);
nand U43020 (N_43020,N_40139,N_41926);
nor U43021 (N_43021,N_41606,N_40236);
nand U43022 (N_43022,N_40200,N_41132);
nand U43023 (N_43023,N_40249,N_41061);
nor U43024 (N_43024,N_40132,N_40262);
nand U43025 (N_43025,N_40567,N_41677);
xor U43026 (N_43026,N_41405,N_41867);
nor U43027 (N_43027,N_40657,N_41267);
nand U43028 (N_43028,N_40189,N_41965);
or U43029 (N_43029,N_40495,N_40095);
nand U43030 (N_43030,N_41625,N_40130);
xor U43031 (N_43031,N_40340,N_40498);
nand U43032 (N_43032,N_40706,N_40122);
xor U43033 (N_43033,N_40584,N_41225);
xor U43034 (N_43034,N_40967,N_40490);
and U43035 (N_43035,N_41671,N_40403);
or U43036 (N_43036,N_40779,N_41849);
nor U43037 (N_43037,N_40180,N_40205);
xnor U43038 (N_43038,N_41720,N_40855);
nand U43039 (N_43039,N_40337,N_41761);
and U43040 (N_43040,N_41373,N_41431);
nor U43041 (N_43041,N_41909,N_41083);
nor U43042 (N_43042,N_41187,N_41767);
xor U43043 (N_43043,N_40738,N_40286);
or U43044 (N_43044,N_40508,N_40173);
or U43045 (N_43045,N_40597,N_41787);
or U43046 (N_43046,N_41896,N_41293);
nor U43047 (N_43047,N_41099,N_40736);
and U43048 (N_43048,N_41603,N_41992);
and U43049 (N_43049,N_40106,N_41030);
or U43050 (N_43050,N_40218,N_41328);
nand U43051 (N_43051,N_41725,N_40758);
nand U43052 (N_43052,N_41150,N_40941);
xnor U43053 (N_43053,N_40769,N_41509);
nand U43054 (N_43054,N_41461,N_40243);
xnor U43055 (N_43055,N_41119,N_41372);
xnor U43056 (N_43056,N_40548,N_41414);
nor U43057 (N_43057,N_40605,N_41837);
nand U43058 (N_43058,N_41039,N_41847);
or U43059 (N_43059,N_40968,N_41715);
nor U43060 (N_43060,N_40200,N_41838);
nor U43061 (N_43061,N_41625,N_40878);
xnor U43062 (N_43062,N_41908,N_41550);
and U43063 (N_43063,N_40547,N_41526);
nor U43064 (N_43064,N_41023,N_41803);
xor U43065 (N_43065,N_41967,N_40973);
and U43066 (N_43066,N_40052,N_40937);
nand U43067 (N_43067,N_40985,N_41602);
nand U43068 (N_43068,N_40636,N_41523);
nand U43069 (N_43069,N_41022,N_41246);
or U43070 (N_43070,N_40316,N_40688);
and U43071 (N_43071,N_40288,N_41085);
and U43072 (N_43072,N_41319,N_41668);
xor U43073 (N_43073,N_41757,N_41141);
nor U43074 (N_43074,N_40828,N_40031);
or U43075 (N_43075,N_40061,N_41678);
nor U43076 (N_43076,N_40247,N_41568);
or U43077 (N_43077,N_41260,N_40536);
nor U43078 (N_43078,N_40714,N_41507);
or U43079 (N_43079,N_41004,N_40533);
xor U43080 (N_43080,N_41871,N_40152);
nand U43081 (N_43081,N_41522,N_40127);
and U43082 (N_43082,N_41532,N_40591);
nand U43083 (N_43083,N_41443,N_41713);
nor U43084 (N_43084,N_40200,N_41142);
nand U43085 (N_43085,N_41566,N_40660);
nand U43086 (N_43086,N_40670,N_41074);
and U43087 (N_43087,N_41417,N_41495);
and U43088 (N_43088,N_41998,N_41878);
or U43089 (N_43089,N_40947,N_41478);
or U43090 (N_43090,N_41562,N_40863);
and U43091 (N_43091,N_40315,N_40653);
or U43092 (N_43092,N_40845,N_40667);
nand U43093 (N_43093,N_40608,N_40750);
and U43094 (N_43094,N_41844,N_40192);
and U43095 (N_43095,N_41191,N_40133);
nand U43096 (N_43096,N_40007,N_40584);
nand U43097 (N_43097,N_41304,N_40534);
and U43098 (N_43098,N_40469,N_41292);
nor U43099 (N_43099,N_41668,N_40530);
nor U43100 (N_43100,N_41221,N_41357);
xnor U43101 (N_43101,N_41005,N_41156);
xor U43102 (N_43102,N_40078,N_41344);
nand U43103 (N_43103,N_41648,N_41012);
xnor U43104 (N_43104,N_41703,N_41177);
xor U43105 (N_43105,N_41919,N_41348);
nand U43106 (N_43106,N_40055,N_40889);
or U43107 (N_43107,N_40811,N_40735);
or U43108 (N_43108,N_41759,N_41697);
and U43109 (N_43109,N_40801,N_40692);
or U43110 (N_43110,N_41761,N_41611);
nand U43111 (N_43111,N_41580,N_40270);
and U43112 (N_43112,N_40374,N_41008);
nor U43113 (N_43113,N_40729,N_40345);
xor U43114 (N_43114,N_40609,N_41270);
nor U43115 (N_43115,N_40931,N_41642);
nor U43116 (N_43116,N_41643,N_41924);
and U43117 (N_43117,N_40742,N_41637);
nor U43118 (N_43118,N_41459,N_40826);
and U43119 (N_43119,N_41806,N_40966);
nand U43120 (N_43120,N_40525,N_41884);
nor U43121 (N_43121,N_40615,N_40672);
and U43122 (N_43122,N_40457,N_41354);
xor U43123 (N_43123,N_41933,N_41126);
nand U43124 (N_43124,N_41419,N_40413);
or U43125 (N_43125,N_41460,N_41280);
or U43126 (N_43126,N_40382,N_41186);
or U43127 (N_43127,N_41570,N_40695);
nor U43128 (N_43128,N_41081,N_41055);
xnor U43129 (N_43129,N_41731,N_40273);
nor U43130 (N_43130,N_40005,N_41622);
nand U43131 (N_43131,N_40307,N_40329);
nor U43132 (N_43132,N_40542,N_40495);
xnor U43133 (N_43133,N_41284,N_40242);
and U43134 (N_43134,N_40484,N_40780);
and U43135 (N_43135,N_40157,N_41614);
nor U43136 (N_43136,N_40119,N_40457);
and U43137 (N_43137,N_41603,N_40506);
or U43138 (N_43138,N_40307,N_41720);
xnor U43139 (N_43139,N_40711,N_40852);
nand U43140 (N_43140,N_40903,N_40069);
nor U43141 (N_43141,N_40778,N_41083);
xnor U43142 (N_43142,N_40220,N_40911);
nand U43143 (N_43143,N_41470,N_40673);
and U43144 (N_43144,N_41416,N_40859);
and U43145 (N_43145,N_40167,N_40932);
and U43146 (N_43146,N_41222,N_41294);
or U43147 (N_43147,N_40641,N_40987);
nand U43148 (N_43148,N_41236,N_40390);
and U43149 (N_43149,N_41613,N_41808);
xnor U43150 (N_43150,N_41822,N_40427);
nand U43151 (N_43151,N_40816,N_40011);
nor U43152 (N_43152,N_40371,N_40790);
xor U43153 (N_43153,N_41348,N_41925);
and U43154 (N_43154,N_40686,N_40820);
nor U43155 (N_43155,N_40966,N_41835);
nand U43156 (N_43156,N_40668,N_41806);
xor U43157 (N_43157,N_40185,N_41378);
nor U43158 (N_43158,N_40683,N_40677);
nor U43159 (N_43159,N_41505,N_40304);
and U43160 (N_43160,N_41171,N_40705);
and U43161 (N_43161,N_40360,N_41528);
or U43162 (N_43162,N_41145,N_41391);
and U43163 (N_43163,N_40239,N_40718);
xor U43164 (N_43164,N_40904,N_41114);
or U43165 (N_43165,N_40567,N_41801);
nand U43166 (N_43166,N_40138,N_41955);
nor U43167 (N_43167,N_41628,N_41171);
nor U43168 (N_43168,N_40282,N_41843);
nand U43169 (N_43169,N_41297,N_40525);
nor U43170 (N_43170,N_40995,N_40903);
nand U43171 (N_43171,N_40750,N_40177);
or U43172 (N_43172,N_40873,N_40084);
xor U43173 (N_43173,N_41786,N_41622);
nand U43174 (N_43174,N_40916,N_41071);
or U43175 (N_43175,N_40158,N_40290);
nand U43176 (N_43176,N_41867,N_40802);
or U43177 (N_43177,N_41432,N_41450);
or U43178 (N_43178,N_41014,N_40471);
or U43179 (N_43179,N_41365,N_40719);
and U43180 (N_43180,N_41147,N_40873);
or U43181 (N_43181,N_41593,N_40553);
or U43182 (N_43182,N_41619,N_41361);
and U43183 (N_43183,N_41900,N_40290);
nand U43184 (N_43184,N_41986,N_40202);
nand U43185 (N_43185,N_41290,N_41093);
or U43186 (N_43186,N_40708,N_41842);
or U43187 (N_43187,N_41208,N_40592);
nand U43188 (N_43188,N_41263,N_40311);
xnor U43189 (N_43189,N_40512,N_41399);
nand U43190 (N_43190,N_41411,N_40422);
nor U43191 (N_43191,N_41847,N_40515);
nor U43192 (N_43192,N_41633,N_40659);
nand U43193 (N_43193,N_40760,N_40569);
or U43194 (N_43194,N_41213,N_41977);
xnor U43195 (N_43195,N_41668,N_41710);
or U43196 (N_43196,N_40641,N_40472);
or U43197 (N_43197,N_40701,N_40495);
xor U43198 (N_43198,N_41141,N_41942);
nand U43199 (N_43199,N_41834,N_41188);
and U43200 (N_43200,N_40020,N_41521);
xor U43201 (N_43201,N_41384,N_41757);
and U43202 (N_43202,N_41977,N_41953);
nand U43203 (N_43203,N_41183,N_40776);
nand U43204 (N_43204,N_40451,N_41091);
and U43205 (N_43205,N_40953,N_41987);
nand U43206 (N_43206,N_40767,N_41790);
and U43207 (N_43207,N_41032,N_40760);
and U43208 (N_43208,N_40808,N_40799);
xnor U43209 (N_43209,N_41654,N_41243);
nand U43210 (N_43210,N_40145,N_40722);
nor U43211 (N_43211,N_41539,N_40547);
or U43212 (N_43212,N_41079,N_40448);
xor U43213 (N_43213,N_40259,N_40875);
or U43214 (N_43214,N_40627,N_40459);
nand U43215 (N_43215,N_41557,N_40396);
xnor U43216 (N_43216,N_41611,N_41508);
xnor U43217 (N_43217,N_41793,N_40200);
xor U43218 (N_43218,N_40295,N_40095);
xnor U43219 (N_43219,N_40549,N_41321);
xnor U43220 (N_43220,N_40136,N_40995);
nand U43221 (N_43221,N_40481,N_41509);
nor U43222 (N_43222,N_40670,N_41144);
or U43223 (N_43223,N_40579,N_40340);
and U43224 (N_43224,N_41594,N_40001);
nor U43225 (N_43225,N_41508,N_40771);
nor U43226 (N_43226,N_40378,N_40229);
xnor U43227 (N_43227,N_40890,N_41118);
nand U43228 (N_43228,N_40673,N_40373);
nor U43229 (N_43229,N_40280,N_41409);
or U43230 (N_43230,N_40359,N_41267);
or U43231 (N_43231,N_41439,N_41407);
nand U43232 (N_43232,N_40654,N_40934);
nand U43233 (N_43233,N_41882,N_40871);
and U43234 (N_43234,N_40482,N_41260);
nand U43235 (N_43235,N_40425,N_40986);
xnor U43236 (N_43236,N_41595,N_40459);
and U43237 (N_43237,N_41273,N_40287);
or U43238 (N_43238,N_40378,N_40779);
nor U43239 (N_43239,N_41214,N_41294);
xor U43240 (N_43240,N_41769,N_40372);
xnor U43241 (N_43241,N_41010,N_41731);
nand U43242 (N_43242,N_40185,N_40765);
and U43243 (N_43243,N_40420,N_41385);
and U43244 (N_43244,N_40503,N_41673);
xnor U43245 (N_43245,N_41151,N_41691);
or U43246 (N_43246,N_40085,N_41090);
nand U43247 (N_43247,N_41484,N_40943);
nand U43248 (N_43248,N_40223,N_40456);
and U43249 (N_43249,N_40633,N_41511);
xnor U43250 (N_43250,N_40884,N_41198);
xnor U43251 (N_43251,N_40487,N_41317);
nor U43252 (N_43252,N_41498,N_40633);
nand U43253 (N_43253,N_40078,N_41975);
and U43254 (N_43254,N_40824,N_40935);
nand U43255 (N_43255,N_40205,N_40204);
or U43256 (N_43256,N_41241,N_41147);
xor U43257 (N_43257,N_40624,N_40256);
nand U43258 (N_43258,N_41738,N_40176);
nor U43259 (N_43259,N_40753,N_40900);
and U43260 (N_43260,N_40246,N_41450);
xor U43261 (N_43261,N_41200,N_41914);
nor U43262 (N_43262,N_40070,N_41455);
nand U43263 (N_43263,N_40273,N_40632);
and U43264 (N_43264,N_40983,N_41521);
or U43265 (N_43265,N_40937,N_40485);
or U43266 (N_43266,N_41187,N_40485);
xnor U43267 (N_43267,N_40919,N_41437);
or U43268 (N_43268,N_41461,N_41980);
xnor U43269 (N_43269,N_41849,N_40823);
xor U43270 (N_43270,N_40952,N_41755);
nand U43271 (N_43271,N_41436,N_41043);
or U43272 (N_43272,N_41367,N_41500);
nand U43273 (N_43273,N_41153,N_40444);
xor U43274 (N_43274,N_41076,N_40109);
nand U43275 (N_43275,N_41452,N_41199);
xor U43276 (N_43276,N_40434,N_40753);
or U43277 (N_43277,N_41594,N_41668);
and U43278 (N_43278,N_41167,N_40920);
nand U43279 (N_43279,N_41392,N_41975);
or U43280 (N_43280,N_41977,N_40661);
and U43281 (N_43281,N_41762,N_40145);
nor U43282 (N_43282,N_40614,N_40256);
or U43283 (N_43283,N_41484,N_40979);
xnor U43284 (N_43284,N_41436,N_40172);
nor U43285 (N_43285,N_41860,N_40327);
nor U43286 (N_43286,N_41855,N_41447);
nor U43287 (N_43287,N_40823,N_40671);
nor U43288 (N_43288,N_41214,N_40316);
or U43289 (N_43289,N_41133,N_40799);
xnor U43290 (N_43290,N_41900,N_41796);
or U43291 (N_43291,N_41436,N_40059);
and U43292 (N_43292,N_40013,N_41327);
nor U43293 (N_43293,N_40514,N_40372);
nor U43294 (N_43294,N_40399,N_40237);
nor U43295 (N_43295,N_41983,N_40131);
nor U43296 (N_43296,N_40942,N_40633);
xnor U43297 (N_43297,N_41340,N_40597);
or U43298 (N_43298,N_40455,N_40405);
or U43299 (N_43299,N_40132,N_40598);
or U43300 (N_43300,N_40724,N_41587);
nor U43301 (N_43301,N_41338,N_40026);
nand U43302 (N_43302,N_40519,N_41356);
xor U43303 (N_43303,N_41427,N_41001);
nor U43304 (N_43304,N_40937,N_40728);
nand U43305 (N_43305,N_40670,N_41301);
and U43306 (N_43306,N_40584,N_41041);
or U43307 (N_43307,N_40313,N_40985);
and U43308 (N_43308,N_41328,N_41049);
xor U43309 (N_43309,N_41100,N_40121);
nand U43310 (N_43310,N_41181,N_41172);
or U43311 (N_43311,N_41508,N_40990);
or U43312 (N_43312,N_41414,N_41399);
nor U43313 (N_43313,N_40185,N_41868);
and U43314 (N_43314,N_40035,N_40185);
and U43315 (N_43315,N_40820,N_40356);
xnor U43316 (N_43316,N_40752,N_40793);
nor U43317 (N_43317,N_41383,N_41623);
nor U43318 (N_43318,N_40469,N_40951);
nand U43319 (N_43319,N_41818,N_40051);
or U43320 (N_43320,N_41551,N_40926);
and U43321 (N_43321,N_41302,N_40562);
xor U43322 (N_43322,N_40725,N_40085);
nand U43323 (N_43323,N_41681,N_40750);
or U43324 (N_43324,N_41696,N_41497);
or U43325 (N_43325,N_41233,N_41923);
or U43326 (N_43326,N_40120,N_40735);
xnor U43327 (N_43327,N_41420,N_40779);
nor U43328 (N_43328,N_41181,N_41482);
xnor U43329 (N_43329,N_41836,N_41988);
nor U43330 (N_43330,N_40969,N_40721);
and U43331 (N_43331,N_41358,N_41208);
nand U43332 (N_43332,N_40005,N_41126);
nand U43333 (N_43333,N_40369,N_40164);
or U43334 (N_43334,N_41707,N_40387);
nand U43335 (N_43335,N_41272,N_41769);
nand U43336 (N_43336,N_41627,N_41937);
nand U43337 (N_43337,N_41784,N_40130);
nor U43338 (N_43338,N_41829,N_40862);
or U43339 (N_43339,N_41445,N_41819);
nor U43340 (N_43340,N_41701,N_41269);
or U43341 (N_43341,N_41631,N_41341);
nor U43342 (N_43342,N_41398,N_40427);
or U43343 (N_43343,N_40480,N_41056);
nor U43344 (N_43344,N_40586,N_40875);
xnor U43345 (N_43345,N_41107,N_41354);
and U43346 (N_43346,N_40241,N_40724);
or U43347 (N_43347,N_41223,N_41887);
nand U43348 (N_43348,N_40616,N_40538);
and U43349 (N_43349,N_40356,N_41622);
nand U43350 (N_43350,N_40849,N_41904);
nand U43351 (N_43351,N_40476,N_40265);
nand U43352 (N_43352,N_40276,N_40885);
nand U43353 (N_43353,N_41397,N_40704);
xnor U43354 (N_43354,N_41652,N_40828);
xnor U43355 (N_43355,N_41275,N_41855);
nor U43356 (N_43356,N_40112,N_40015);
nor U43357 (N_43357,N_40203,N_41196);
and U43358 (N_43358,N_41107,N_40144);
or U43359 (N_43359,N_41066,N_41773);
xor U43360 (N_43360,N_41540,N_41487);
and U43361 (N_43361,N_41446,N_41595);
or U43362 (N_43362,N_40495,N_40448);
nor U43363 (N_43363,N_40962,N_41711);
or U43364 (N_43364,N_40096,N_40356);
or U43365 (N_43365,N_40695,N_41889);
and U43366 (N_43366,N_41933,N_40340);
and U43367 (N_43367,N_40009,N_41232);
nand U43368 (N_43368,N_41577,N_41234);
nand U43369 (N_43369,N_40121,N_40435);
nor U43370 (N_43370,N_40689,N_40682);
or U43371 (N_43371,N_40753,N_41760);
nor U43372 (N_43372,N_40500,N_40107);
nand U43373 (N_43373,N_41184,N_40808);
nand U43374 (N_43374,N_41639,N_41617);
nor U43375 (N_43375,N_40143,N_41193);
and U43376 (N_43376,N_41241,N_40959);
or U43377 (N_43377,N_40479,N_41721);
xor U43378 (N_43378,N_41716,N_40869);
and U43379 (N_43379,N_41010,N_41178);
or U43380 (N_43380,N_41501,N_41076);
nor U43381 (N_43381,N_40425,N_41020);
nand U43382 (N_43382,N_41861,N_41061);
xnor U43383 (N_43383,N_40050,N_41807);
xor U43384 (N_43384,N_40291,N_40255);
nand U43385 (N_43385,N_40859,N_40817);
nand U43386 (N_43386,N_40055,N_41221);
or U43387 (N_43387,N_41467,N_40059);
xor U43388 (N_43388,N_40239,N_40982);
or U43389 (N_43389,N_40765,N_40665);
nor U43390 (N_43390,N_40280,N_41656);
or U43391 (N_43391,N_40029,N_40827);
or U43392 (N_43392,N_40121,N_41917);
or U43393 (N_43393,N_40230,N_41268);
xor U43394 (N_43394,N_41148,N_41567);
or U43395 (N_43395,N_40420,N_40689);
or U43396 (N_43396,N_40174,N_40747);
nor U43397 (N_43397,N_41761,N_41591);
nor U43398 (N_43398,N_40762,N_40909);
or U43399 (N_43399,N_40064,N_40370);
or U43400 (N_43400,N_41308,N_41687);
and U43401 (N_43401,N_41829,N_40526);
xnor U43402 (N_43402,N_40658,N_41481);
nor U43403 (N_43403,N_40766,N_40407);
nand U43404 (N_43404,N_40247,N_41144);
or U43405 (N_43405,N_41206,N_40750);
nand U43406 (N_43406,N_41941,N_41266);
nand U43407 (N_43407,N_40968,N_40681);
and U43408 (N_43408,N_41752,N_40435);
xnor U43409 (N_43409,N_41152,N_41008);
or U43410 (N_43410,N_40789,N_40286);
xor U43411 (N_43411,N_41907,N_41809);
or U43412 (N_43412,N_41587,N_40632);
xor U43413 (N_43413,N_41675,N_41787);
nand U43414 (N_43414,N_40546,N_40706);
nand U43415 (N_43415,N_41987,N_40739);
or U43416 (N_43416,N_40603,N_40269);
and U43417 (N_43417,N_41534,N_41696);
or U43418 (N_43418,N_41185,N_41517);
nor U43419 (N_43419,N_41599,N_41548);
xnor U43420 (N_43420,N_40193,N_41174);
nor U43421 (N_43421,N_40175,N_41916);
and U43422 (N_43422,N_41205,N_41339);
nor U43423 (N_43423,N_41674,N_40746);
xnor U43424 (N_43424,N_40720,N_41411);
or U43425 (N_43425,N_41055,N_40032);
nand U43426 (N_43426,N_40188,N_41805);
xnor U43427 (N_43427,N_41521,N_41920);
or U43428 (N_43428,N_41348,N_41875);
nor U43429 (N_43429,N_40237,N_40454);
nand U43430 (N_43430,N_41291,N_41978);
nor U43431 (N_43431,N_41615,N_41463);
xor U43432 (N_43432,N_40136,N_41085);
or U43433 (N_43433,N_41870,N_41160);
or U43434 (N_43434,N_40093,N_41968);
nor U43435 (N_43435,N_41564,N_40199);
nand U43436 (N_43436,N_41208,N_41776);
or U43437 (N_43437,N_41577,N_41056);
nand U43438 (N_43438,N_40250,N_41492);
or U43439 (N_43439,N_40788,N_40152);
and U43440 (N_43440,N_40758,N_40321);
xor U43441 (N_43441,N_40925,N_41037);
nor U43442 (N_43442,N_40995,N_40579);
nand U43443 (N_43443,N_41217,N_41703);
or U43444 (N_43444,N_41721,N_41951);
nor U43445 (N_43445,N_40965,N_41043);
and U43446 (N_43446,N_40608,N_40918);
xnor U43447 (N_43447,N_41092,N_40270);
nor U43448 (N_43448,N_40657,N_41184);
xnor U43449 (N_43449,N_40283,N_40937);
nor U43450 (N_43450,N_41107,N_41692);
and U43451 (N_43451,N_40543,N_40961);
and U43452 (N_43452,N_41050,N_40939);
and U43453 (N_43453,N_41371,N_41068);
nor U43454 (N_43454,N_40629,N_40361);
or U43455 (N_43455,N_40586,N_40869);
xnor U43456 (N_43456,N_40960,N_41474);
nor U43457 (N_43457,N_41549,N_41569);
nor U43458 (N_43458,N_40470,N_40169);
and U43459 (N_43459,N_41407,N_41327);
or U43460 (N_43460,N_41483,N_41945);
xnor U43461 (N_43461,N_40109,N_41858);
nor U43462 (N_43462,N_40721,N_41643);
nand U43463 (N_43463,N_41603,N_40278);
xor U43464 (N_43464,N_41752,N_41716);
and U43465 (N_43465,N_41239,N_40198);
nand U43466 (N_43466,N_41952,N_41919);
or U43467 (N_43467,N_41248,N_41536);
or U43468 (N_43468,N_41377,N_41028);
xor U43469 (N_43469,N_40071,N_41501);
nand U43470 (N_43470,N_40169,N_41114);
nor U43471 (N_43471,N_40958,N_41132);
nor U43472 (N_43472,N_40574,N_41553);
nor U43473 (N_43473,N_41968,N_40439);
and U43474 (N_43474,N_40771,N_41094);
or U43475 (N_43475,N_41737,N_41968);
xor U43476 (N_43476,N_41385,N_40892);
nor U43477 (N_43477,N_41927,N_41529);
nor U43478 (N_43478,N_40628,N_41761);
and U43479 (N_43479,N_41674,N_41039);
or U43480 (N_43480,N_40964,N_40003);
or U43481 (N_43481,N_41787,N_40638);
xnor U43482 (N_43482,N_40941,N_41320);
nor U43483 (N_43483,N_40944,N_40640);
or U43484 (N_43484,N_41360,N_40034);
or U43485 (N_43485,N_40842,N_40033);
nand U43486 (N_43486,N_41664,N_40312);
xnor U43487 (N_43487,N_41750,N_41913);
or U43488 (N_43488,N_41682,N_41593);
xor U43489 (N_43489,N_40826,N_40282);
or U43490 (N_43490,N_41434,N_40754);
xnor U43491 (N_43491,N_40687,N_40856);
nand U43492 (N_43492,N_40537,N_41452);
nor U43493 (N_43493,N_41973,N_41751);
xnor U43494 (N_43494,N_40592,N_40408);
nand U43495 (N_43495,N_40286,N_41211);
and U43496 (N_43496,N_41985,N_40504);
nor U43497 (N_43497,N_40708,N_41089);
or U43498 (N_43498,N_40404,N_40635);
nor U43499 (N_43499,N_40130,N_40206);
or U43500 (N_43500,N_41262,N_40938);
or U43501 (N_43501,N_40995,N_41650);
or U43502 (N_43502,N_40905,N_40306);
xor U43503 (N_43503,N_41295,N_41059);
xor U43504 (N_43504,N_41898,N_40453);
nand U43505 (N_43505,N_41558,N_41251);
xor U43506 (N_43506,N_40255,N_41673);
nand U43507 (N_43507,N_40340,N_40503);
nor U43508 (N_43508,N_40289,N_40388);
and U43509 (N_43509,N_41448,N_41518);
and U43510 (N_43510,N_41250,N_41228);
and U43511 (N_43511,N_40287,N_41479);
nor U43512 (N_43512,N_41449,N_40191);
nand U43513 (N_43513,N_40434,N_41071);
or U43514 (N_43514,N_40236,N_40889);
nor U43515 (N_43515,N_41910,N_40052);
nor U43516 (N_43516,N_41606,N_40787);
or U43517 (N_43517,N_41382,N_41762);
or U43518 (N_43518,N_40055,N_41123);
nand U43519 (N_43519,N_41263,N_41260);
and U43520 (N_43520,N_40159,N_41349);
nand U43521 (N_43521,N_40751,N_40521);
or U43522 (N_43522,N_41960,N_40424);
xnor U43523 (N_43523,N_41147,N_40379);
xnor U43524 (N_43524,N_41625,N_41214);
xor U43525 (N_43525,N_40330,N_40919);
or U43526 (N_43526,N_41050,N_41451);
and U43527 (N_43527,N_41096,N_41088);
and U43528 (N_43528,N_40079,N_41228);
and U43529 (N_43529,N_40227,N_41270);
nor U43530 (N_43530,N_40807,N_41393);
xnor U43531 (N_43531,N_41482,N_40842);
or U43532 (N_43532,N_41045,N_40119);
nand U43533 (N_43533,N_41995,N_41882);
nand U43534 (N_43534,N_41086,N_41015);
and U43535 (N_43535,N_40878,N_40713);
nor U43536 (N_43536,N_40512,N_40918);
xor U43537 (N_43537,N_41584,N_41287);
or U43538 (N_43538,N_40900,N_41363);
and U43539 (N_43539,N_41734,N_41316);
nand U43540 (N_43540,N_41163,N_41880);
nor U43541 (N_43541,N_41728,N_41661);
nand U43542 (N_43542,N_40885,N_40439);
and U43543 (N_43543,N_41739,N_40457);
nor U43544 (N_43544,N_40697,N_40430);
or U43545 (N_43545,N_41664,N_40387);
nor U43546 (N_43546,N_41806,N_41908);
xor U43547 (N_43547,N_40510,N_41168);
or U43548 (N_43548,N_41238,N_41476);
nor U43549 (N_43549,N_40579,N_40563);
and U43550 (N_43550,N_41475,N_40854);
nand U43551 (N_43551,N_40765,N_40456);
nand U43552 (N_43552,N_40099,N_41962);
xnor U43553 (N_43553,N_40365,N_41233);
and U43554 (N_43554,N_41166,N_40815);
and U43555 (N_43555,N_40833,N_40588);
or U43556 (N_43556,N_41221,N_40621);
xnor U43557 (N_43557,N_40214,N_41855);
and U43558 (N_43558,N_41582,N_41576);
nor U43559 (N_43559,N_40555,N_40057);
nor U43560 (N_43560,N_40455,N_41838);
nor U43561 (N_43561,N_40314,N_41181);
and U43562 (N_43562,N_41519,N_40054);
or U43563 (N_43563,N_41924,N_41462);
and U43564 (N_43564,N_40853,N_41017);
nand U43565 (N_43565,N_41049,N_41060);
or U43566 (N_43566,N_41348,N_41025);
nand U43567 (N_43567,N_40809,N_40868);
nand U43568 (N_43568,N_41315,N_40383);
xor U43569 (N_43569,N_41502,N_41226);
or U43570 (N_43570,N_40572,N_40529);
xor U43571 (N_43571,N_41190,N_41655);
and U43572 (N_43572,N_40853,N_40481);
nor U43573 (N_43573,N_41522,N_40404);
nor U43574 (N_43574,N_40358,N_41618);
nor U43575 (N_43575,N_41935,N_41424);
and U43576 (N_43576,N_40888,N_41354);
nor U43577 (N_43577,N_41571,N_41118);
nor U43578 (N_43578,N_40621,N_41980);
nor U43579 (N_43579,N_41759,N_41110);
or U43580 (N_43580,N_41878,N_41606);
nor U43581 (N_43581,N_41499,N_40844);
and U43582 (N_43582,N_40555,N_41379);
and U43583 (N_43583,N_41166,N_41997);
or U43584 (N_43584,N_41252,N_40610);
or U43585 (N_43585,N_40696,N_40358);
xor U43586 (N_43586,N_41654,N_41150);
xor U43587 (N_43587,N_40884,N_41309);
and U43588 (N_43588,N_40956,N_41581);
nor U43589 (N_43589,N_41115,N_41541);
or U43590 (N_43590,N_41673,N_41869);
or U43591 (N_43591,N_41845,N_40011);
nand U43592 (N_43592,N_40498,N_41825);
and U43593 (N_43593,N_40874,N_41015);
nand U43594 (N_43594,N_41242,N_40904);
or U43595 (N_43595,N_40223,N_41242);
xor U43596 (N_43596,N_41981,N_41822);
nor U43597 (N_43597,N_40964,N_41153);
or U43598 (N_43598,N_41668,N_40442);
or U43599 (N_43599,N_41352,N_41295);
and U43600 (N_43600,N_40324,N_40757);
and U43601 (N_43601,N_41443,N_40450);
nand U43602 (N_43602,N_40768,N_41401);
nand U43603 (N_43603,N_40594,N_41563);
nor U43604 (N_43604,N_40267,N_40519);
nor U43605 (N_43605,N_41169,N_40899);
nor U43606 (N_43606,N_41405,N_40672);
nor U43607 (N_43607,N_40451,N_40918);
xor U43608 (N_43608,N_40984,N_41196);
xnor U43609 (N_43609,N_40448,N_41654);
nor U43610 (N_43610,N_41750,N_41581);
nand U43611 (N_43611,N_41340,N_40388);
xor U43612 (N_43612,N_41335,N_40580);
and U43613 (N_43613,N_40324,N_40300);
and U43614 (N_43614,N_40842,N_40474);
nor U43615 (N_43615,N_41005,N_40704);
or U43616 (N_43616,N_40754,N_40534);
nand U43617 (N_43617,N_40599,N_41554);
xor U43618 (N_43618,N_41874,N_40182);
xor U43619 (N_43619,N_40018,N_40874);
xor U43620 (N_43620,N_40765,N_40615);
nand U43621 (N_43621,N_40524,N_41198);
nand U43622 (N_43622,N_41045,N_41582);
and U43623 (N_43623,N_40323,N_41664);
xnor U43624 (N_43624,N_40088,N_41623);
or U43625 (N_43625,N_41934,N_40856);
nand U43626 (N_43626,N_40409,N_40006);
or U43627 (N_43627,N_40068,N_41713);
nor U43628 (N_43628,N_40659,N_40623);
and U43629 (N_43629,N_40997,N_40831);
xor U43630 (N_43630,N_41140,N_41278);
and U43631 (N_43631,N_41004,N_41969);
nor U43632 (N_43632,N_40449,N_40853);
and U43633 (N_43633,N_41557,N_41721);
nor U43634 (N_43634,N_40261,N_41332);
nor U43635 (N_43635,N_40515,N_41566);
nand U43636 (N_43636,N_41646,N_40074);
or U43637 (N_43637,N_41780,N_41694);
and U43638 (N_43638,N_41088,N_40349);
or U43639 (N_43639,N_41727,N_41538);
and U43640 (N_43640,N_40790,N_41073);
nor U43641 (N_43641,N_41072,N_40574);
or U43642 (N_43642,N_40563,N_40330);
nand U43643 (N_43643,N_41468,N_41771);
xor U43644 (N_43644,N_40188,N_41777);
and U43645 (N_43645,N_40773,N_40952);
xnor U43646 (N_43646,N_41491,N_41125);
and U43647 (N_43647,N_40319,N_41227);
xnor U43648 (N_43648,N_41947,N_41209);
or U43649 (N_43649,N_41914,N_41000);
or U43650 (N_43650,N_41485,N_40798);
or U43651 (N_43651,N_41299,N_41451);
or U43652 (N_43652,N_40373,N_41987);
xor U43653 (N_43653,N_40640,N_40122);
nand U43654 (N_43654,N_40831,N_41634);
or U43655 (N_43655,N_40208,N_40566);
xor U43656 (N_43656,N_40552,N_41734);
nor U43657 (N_43657,N_40529,N_40708);
and U43658 (N_43658,N_41882,N_40448);
nand U43659 (N_43659,N_41572,N_40523);
and U43660 (N_43660,N_40439,N_40922);
xnor U43661 (N_43661,N_41749,N_40093);
nor U43662 (N_43662,N_41066,N_40689);
and U43663 (N_43663,N_41971,N_40777);
xor U43664 (N_43664,N_41623,N_41369);
and U43665 (N_43665,N_41608,N_41387);
and U43666 (N_43666,N_41611,N_40892);
nand U43667 (N_43667,N_40750,N_41640);
nand U43668 (N_43668,N_41080,N_41960);
and U43669 (N_43669,N_40998,N_41720);
nor U43670 (N_43670,N_41733,N_41065);
or U43671 (N_43671,N_40104,N_40210);
and U43672 (N_43672,N_41711,N_40520);
and U43673 (N_43673,N_40429,N_40475);
xnor U43674 (N_43674,N_41265,N_41576);
or U43675 (N_43675,N_41344,N_40885);
or U43676 (N_43676,N_40777,N_40329);
nor U43677 (N_43677,N_40664,N_41452);
nor U43678 (N_43678,N_40311,N_40886);
xnor U43679 (N_43679,N_41461,N_41696);
nor U43680 (N_43680,N_41440,N_41489);
nand U43681 (N_43681,N_40947,N_40747);
xnor U43682 (N_43682,N_40183,N_40690);
and U43683 (N_43683,N_40710,N_40968);
xnor U43684 (N_43684,N_41354,N_40826);
nor U43685 (N_43685,N_40336,N_40486);
xor U43686 (N_43686,N_40279,N_40287);
and U43687 (N_43687,N_41144,N_41662);
nor U43688 (N_43688,N_41001,N_41225);
nand U43689 (N_43689,N_41697,N_41332);
xor U43690 (N_43690,N_41743,N_41862);
nand U43691 (N_43691,N_41351,N_40500);
nand U43692 (N_43692,N_40904,N_40170);
or U43693 (N_43693,N_40046,N_40064);
and U43694 (N_43694,N_40764,N_40823);
nand U43695 (N_43695,N_41477,N_41942);
xnor U43696 (N_43696,N_41941,N_41255);
xor U43697 (N_43697,N_40537,N_40288);
xnor U43698 (N_43698,N_40824,N_41229);
nor U43699 (N_43699,N_41879,N_41059);
nor U43700 (N_43700,N_41234,N_40249);
nor U43701 (N_43701,N_40760,N_40089);
and U43702 (N_43702,N_40775,N_40741);
nor U43703 (N_43703,N_40323,N_40021);
nand U43704 (N_43704,N_41908,N_40868);
nand U43705 (N_43705,N_40955,N_41932);
and U43706 (N_43706,N_40972,N_41201);
or U43707 (N_43707,N_41176,N_41190);
and U43708 (N_43708,N_40630,N_41387);
and U43709 (N_43709,N_40573,N_41515);
nor U43710 (N_43710,N_40342,N_41977);
or U43711 (N_43711,N_40301,N_41425);
or U43712 (N_43712,N_41895,N_40810);
nor U43713 (N_43713,N_41479,N_41522);
xnor U43714 (N_43714,N_40964,N_40531);
and U43715 (N_43715,N_40868,N_41597);
xnor U43716 (N_43716,N_41574,N_41830);
and U43717 (N_43717,N_40045,N_41090);
nand U43718 (N_43718,N_40962,N_40147);
nor U43719 (N_43719,N_40337,N_40414);
or U43720 (N_43720,N_41668,N_40695);
or U43721 (N_43721,N_41938,N_41992);
xnor U43722 (N_43722,N_40448,N_40481);
nand U43723 (N_43723,N_41405,N_40533);
xor U43724 (N_43724,N_40622,N_40713);
or U43725 (N_43725,N_40761,N_40433);
xnor U43726 (N_43726,N_41968,N_40138);
and U43727 (N_43727,N_41699,N_40354);
nand U43728 (N_43728,N_40932,N_40392);
xor U43729 (N_43729,N_41081,N_41275);
nand U43730 (N_43730,N_41449,N_41288);
xnor U43731 (N_43731,N_40261,N_40416);
and U43732 (N_43732,N_40532,N_40804);
or U43733 (N_43733,N_40873,N_40004);
and U43734 (N_43734,N_40886,N_40653);
or U43735 (N_43735,N_41096,N_41028);
xor U43736 (N_43736,N_41616,N_41889);
nand U43737 (N_43737,N_41624,N_40093);
nor U43738 (N_43738,N_41146,N_41832);
xor U43739 (N_43739,N_40605,N_41775);
or U43740 (N_43740,N_40007,N_40327);
nor U43741 (N_43741,N_41302,N_40545);
nand U43742 (N_43742,N_41719,N_41695);
nor U43743 (N_43743,N_40482,N_41893);
nor U43744 (N_43744,N_41106,N_41842);
and U43745 (N_43745,N_41845,N_40463);
and U43746 (N_43746,N_41331,N_41754);
and U43747 (N_43747,N_41888,N_40452);
xor U43748 (N_43748,N_40011,N_41334);
nand U43749 (N_43749,N_40882,N_40742);
xor U43750 (N_43750,N_40169,N_41576);
or U43751 (N_43751,N_40504,N_41485);
or U43752 (N_43752,N_40892,N_41465);
nor U43753 (N_43753,N_40242,N_41183);
nand U43754 (N_43754,N_40501,N_40874);
nor U43755 (N_43755,N_40711,N_40080);
xnor U43756 (N_43756,N_40907,N_40949);
nand U43757 (N_43757,N_40465,N_41217);
nand U43758 (N_43758,N_41065,N_40705);
nand U43759 (N_43759,N_40205,N_41066);
and U43760 (N_43760,N_40999,N_41741);
nor U43761 (N_43761,N_40399,N_40640);
nor U43762 (N_43762,N_40079,N_40528);
nor U43763 (N_43763,N_41279,N_41309);
xnor U43764 (N_43764,N_41326,N_41192);
and U43765 (N_43765,N_40919,N_40993);
nor U43766 (N_43766,N_40454,N_41902);
nand U43767 (N_43767,N_40149,N_41669);
nor U43768 (N_43768,N_41038,N_40398);
and U43769 (N_43769,N_41763,N_40570);
nor U43770 (N_43770,N_41266,N_40448);
or U43771 (N_43771,N_40388,N_40394);
and U43772 (N_43772,N_41164,N_40614);
and U43773 (N_43773,N_40507,N_40258);
nor U43774 (N_43774,N_41587,N_40388);
xor U43775 (N_43775,N_40756,N_40650);
nand U43776 (N_43776,N_40460,N_40520);
nor U43777 (N_43777,N_40037,N_41876);
and U43778 (N_43778,N_40478,N_41378);
xnor U43779 (N_43779,N_40687,N_41793);
nand U43780 (N_43780,N_41496,N_41389);
nand U43781 (N_43781,N_40609,N_40016);
and U43782 (N_43782,N_41332,N_41136);
and U43783 (N_43783,N_40775,N_41097);
nor U43784 (N_43784,N_41749,N_40798);
nor U43785 (N_43785,N_40639,N_40894);
or U43786 (N_43786,N_40890,N_41396);
or U43787 (N_43787,N_41228,N_41145);
xor U43788 (N_43788,N_40672,N_40020);
nand U43789 (N_43789,N_41030,N_40436);
xor U43790 (N_43790,N_40468,N_41076);
nor U43791 (N_43791,N_41075,N_41823);
and U43792 (N_43792,N_41319,N_41358);
or U43793 (N_43793,N_41281,N_41814);
or U43794 (N_43794,N_41662,N_41766);
nor U43795 (N_43795,N_40264,N_40619);
or U43796 (N_43796,N_40202,N_41619);
and U43797 (N_43797,N_40928,N_41699);
and U43798 (N_43798,N_41997,N_40376);
and U43799 (N_43799,N_41563,N_40263);
nor U43800 (N_43800,N_41057,N_41781);
nand U43801 (N_43801,N_41463,N_41710);
and U43802 (N_43802,N_40719,N_41685);
and U43803 (N_43803,N_40155,N_41747);
xnor U43804 (N_43804,N_41564,N_40224);
or U43805 (N_43805,N_41798,N_41882);
xnor U43806 (N_43806,N_41437,N_41265);
xnor U43807 (N_43807,N_40951,N_40821);
and U43808 (N_43808,N_41986,N_41266);
or U43809 (N_43809,N_40594,N_40595);
nor U43810 (N_43810,N_40375,N_40438);
nand U43811 (N_43811,N_40325,N_41865);
nand U43812 (N_43812,N_40257,N_40726);
nand U43813 (N_43813,N_40284,N_40741);
and U43814 (N_43814,N_40846,N_41057);
xor U43815 (N_43815,N_41788,N_41057);
and U43816 (N_43816,N_40859,N_41998);
nor U43817 (N_43817,N_40726,N_41712);
or U43818 (N_43818,N_41580,N_40578);
nor U43819 (N_43819,N_40135,N_40830);
nor U43820 (N_43820,N_41488,N_41789);
or U43821 (N_43821,N_40974,N_40156);
and U43822 (N_43822,N_40325,N_40037);
nand U43823 (N_43823,N_41245,N_40712);
nor U43824 (N_43824,N_40023,N_40067);
and U43825 (N_43825,N_41924,N_40629);
and U43826 (N_43826,N_41823,N_40095);
or U43827 (N_43827,N_41110,N_41712);
nor U43828 (N_43828,N_40441,N_40865);
and U43829 (N_43829,N_40879,N_41729);
nand U43830 (N_43830,N_41463,N_40806);
nor U43831 (N_43831,N_41462,N_40679);
or U43832 (N_43832,N_41835,N_40928);
or U43833 (N_43833,N_41815,N_41675);
or U43834 (N_43834,N_40817,N_41863);
nand U43835 (N_43835,N_41247,N_41751);
nand U43836 (N_43836,N_40540,N_41778);
or U43837 (N_43837,N_41069,N_41431);
nor U43838 (N_43838,N_40759,N_40771);
nor U43839 (N_43839,N_40216,N_40645);
or U43840 (N_43840,N_40764,N_40421);
and U43841 (N_43841,N_41387,N_40154);
xor U43842 (N_43842,N_40354,N_40079);
nand U43843 (N_43843,N_40541,N_40701);
nor U43844 (N_43844,N_41111,N_40383);
and U43845 (N_43845,N_41084,N_41116);
nand U43846 (N_43846,N_40154,N_40601);
nand U43847 (N_43847,N_40364,N_40101);
nor U43848 (N_43848,N_40229,N_40657);
xor U43849 (N_43849,N_40926,N_40039);
nor U43850 (N_43850,N_40180,N_41230);
nand U43851 (N_43851,N_40721,N_41931);
or U43852 (N_43852,N_41101,N_40155);
and U43853 (N_43853,N_40344,N_41716);
or U43854 (N_43854,N_40796,N_40268);
and U43855 (N_43855,N_40542,N_40950);
and U43856 (N_43856,N_40345,N_40166);
nor U43857 (N_43857,N_41421,N_41318);
nand U43858 (N_43858,N_40561,N_40087);
or U43859 (N_43859,N_41846,N_41355);
or U43860 (N_43860,N_41650,N_41481);
nor U43861 (N_43861,N_40979,N_41175);
or U43862 (N_43862,N_41415,N_40962);
nand U43863 (N_43863,N_41991,N_41730);
xnor U43864 (N_43864,N_41155,N_41518);
nor U43865 (N_43865,N_41618,N_40325);
nor U43866 (N_43866,N_41294,N_41648);
nor U43867 (N_43867,N_40947,N_41896);
and U43868 (N_43868,N_40284,N_40044);
xor U43869 (N_43869,N_41795,N_41752);
and U43870 (N_43870,N_40775,N_41492);
xor U43871 (N_43871,N_40492,N_40331);
nand U43872 (N_43872,N_40799,N_41516);
and U43873 (N_43873,N_40992,N_40021);
xnor U43874 (N_43874,N_41210,N_40929);
or U43875 (N_43875,N_40298,N_40139);
or U43876 (N_43876,N_40088,N_41383);
nor U43877 (N_43877,N_40145,N_41975);
or U43878 (N_43878,N_40323,N_40031);
and U43879 (N_43879,N_41194,N_41043);
nand U43880 (N_43880,N_41797,N_40125);
and U43881 (N_43881,N_41859,N_41956);
nand U43882 (N_43882,N_41371,N_41705);
and U43883 (N_43883,N_41531,N_41524);
xnor U43884 (N_43884,N_41002,N_40690);
xor U43885 (N_43885,N_41274,N_40371);
and U43886 (N_43886,N_41362,N_41313);
xnor U43887 (N_43887,N_40326,N_41436);
nand U43888 (N_43888,N_40459,N_40475);
nor U43889 (N_43889,N_40639,N_40144);
nor U43890 (N_43890,N_41271,N_41297);
nand U43891 (N_43891,N_40302,N_40839);
xor U43892 (N_43892,N_40308,N_41556);
xor U43893 (N_43893,N_41280,N_41494);
nand U43894 (N_43894,N_41754,N_40833);
nand U43895 (N_43895,N_41163,N_41306);
nand U43896 (N_43896,N_40492,N_40507);
or U43897 (N_43897,N_40571,N_40277);
or U43898 (N_43898,N_41718,N_41133);
xnor U43899 (N_43899,N_41968,N_41045);
or U43900 (N_43900,N_40759,N_40797);
nor U43901 (N_43901,N_40645,N_41997);
and U43902 (N_43902,N_41000,N_40786);
nor U43903 (N_43903,N_41193,N_40101);
xor U43904 (N_43904,N_41790,N_40000);
nor U43905 (N_43905,N_41195,N_41991);
xnor U43906 (N_43906,N_41314,N_40675);
and U43907 (N_43907,N_40740,N_41961);
nand U43908 (N_43908,N_40198,N_40879);
nand U43909 (N_43909,N_40229,N_41349);
nand U43910 (N_43910,N_40432,N_41469);
nor U43911 (N_43911,N_40993,N_40415);
and U43912 (N_43912,N_41499,N_40094);
nor U43913 (N_43913,N_41193,N_41952);
xnor U43914 (N_43914,N_40428,N_41226);
or U43915 (N_43915,N_41874,N_41439);
nand U43916 (N_43916,N_41100,N_41160);
nand U43917 (N_43917,N_40028,N_41058);
nor U43918 (N_43918,N_40215,N_40385);
and U43919 (N_43919,N_40841,N_40260);
xnor U43920 (N_43920,N_41089,N_40351);
nor U43921 (N_43921,N_40428,N_40947);
xnor U43922 (N_43922,N_40642,N_41416);
xor U43923 (N_43923,N_40378,N_41132);
and U43924 (N_43924,N_40135,N_40194);
nand U43925 (N_43925,N_40381,N_41159);
xnor U43926 (N_43926,N_40050,N_41349);
xnor U43927 (N_43927,N_40325,N_41023);
or U43928 (N_43928,N_41892,N_40771);
nor U43929 (N_43929,N_41854,N_40912);
and U43930 (N_43930,N_40190,N_41648);
or U43931 (N_43931,N_40215,N_40634);
and U43932 (N_43932,N_41143,N_41964);
nand U43933 (N_43933,N_40955,N_41837);
nor U43934 (N_43934,N_40297,N_40082);
and U43935 (N_43935,N_40196,N_40383);
or U43936 (N_43936,N_40018,N_41773);
or U43937 (N_43937,N_40512,N_41943);
nor U43938 (N_43938,N_40190,N_41845);
nor U43939 (N_43939,N_40823,N_40899);
or U43940 (N_43940,N_40699,N_41108);
nand U43941 (N_43941,N_40139,N_40580);
xnor U43942 (N_43942,N_41454,N_41974);
and U43943 (N_43943,N_40355,N_40959);
nor U43944 (N_43944,N_40049,N_40179);
xnor U43945 (N_43945,N_41486,N_41184);
xnor U43946 (N_43946,N_41704,N_40203);
xor U43947 (N_43947,N_41621,N_40549);
and U43948 (N_43948,N_40816,N_40527);
xnor U43949 (N_43949,N_41062,N_41211);
and U43950 (N_43950,N_40436,N_41261);
and U43951 (N_43951,N_40752,N_40857);
or U43952 (N_43952,N_40683,N_40079);
nor U43953 (N_43953,N_40720,N_40740);
nor U43954 (N_43954,N_40659,N_40573);
and U43955 (N_43955,N_40240,N_41855);
xnor U43956 (N_43956,N_41712,N_41895);
and U43957 (N_43957,N_40339,N_40819);
xnor U43958 (N_43958,N_40928,N_41312);
xor U43959 (N_43959,N_40071,N_40882);
nor U43960 (N_43960,N_41874,N_41672);
and U43961 (N_43961,N_41543,N_40797);
nand U43962 (N_43962,N_40082,N_40777);
xnor U43963 (N_43963,N_41898,N_40579);
and U43964 (N_43964,N_40032,N_40221);
or U43965 (N_43965,N_41413,N_41902);
nand U43966 (N_43966,N_41201,N_40696);
nand U43967 (N_43967,N_41862,N_41181);
nand U43968 (N_43968,N_41543,N_40480);
or U43969 (N_43969,N_40612,N_40044);
nand U43970 (N_43970,N_40382,N_41464);
nor U43971 (N_43971,N_40599,N_40761);
nor U43972 (N_43972,N_40518,N_40005);
and U43973 (N_43973,N_40108,N_41645);
nand U43974 (N_43974,N_40971,N_41259);
or U43975 (N_43975,N_41026,N_40259);
xor U43976 (N_43976,N_40887,N_41681);
nor U43977 (N_43977,N_41119,N_41433);
nor U43978 (N_43978,N_40910,N_40741);
or U43979 (N_43979,N_41863,N_40731);
or U43980 (N_43980,N_40137,N_41352);
or U43981 (N_43981,N_40711,N_41271);
or U43982 (N_43982,N_40354,N_41148);
or U43983 (N_43983,N_41017,N_41613);
and U43984 (N_43984,N_40557,N_41037);
xor U43985 (N_43985,N_41251,N_40336);
nor U43986 (N_43986,N_40293,N_40555);
xor U43987 (N_43987,N_41924,N_40291);
and U43988 (N_43988,N_40076,N_41670);
xnor U43989 (N_43989,N_40572,N_41130);
nor U43990 (N_43990,N_41905,N_40216);
nor U43991 (N_43991,N_40689,N_41518);
nand U43992 (N_43992,N_40092,N_41280);
nand U43993 (N_43993,N_41774,N_40123);
and U43994 (N_43994,N_41107,N_40004);
and U43995 (N_43995,N_40979,N_40042);
nand U43996 (N_43996,N_40083,N_40992);
nor U43997 (N_43997,N_41754,N_40628);
nand U43998 (N_43998,N_40217,N_40748);
and U43999 (N_43999,N_40855,N_40163);
xnor U44000 (N_44000,N_43834,N_42196);
nor U44001 (N_44001,N_42409,N_42365);
nand U44002 (N_44002,N_43238,N_43245);
or U44003 (N_44003,N_43553,N_43389);
or U44004 (N_44004,N_42935,N_43848);
xor U44005 (N_44005,N_43923,N_43622);
nor U44006 (N_44006,N_43899,N_43631);
nand U44007 (N_44007,N_42502,N_43823);
or U44008 (N_44008,N_42452,N_42705);
nand U44009 (N_44009,N_43168,N_43390);
and U44010 (N_44010,N_43911,N_42340);
or U44011 (N_44011,N_43656,N_43675);
nor U44012 (N_44012,N_42082,N_42251);
nor U44013 (N_44013,N_42083,N_43567);
nand U44014 (N_44014,N_42779,N_43726);
and U44015 (N_44015,N_42938,N_42637);
and U44016 (N_44016,N_42173,N_42621);
xor U44017 (N_44017,N_43912,N_43134);
and U44018 (N_44018,N_43316,N_42035);
xnor U44019 (N_44019,N_43291,N_42649);
xnor U44020 (N_44020,N_43017,N_42027);
nor U44021 (N_44021,N_43585,N_42540);
and U44022 (N_44022,N_43318,N_43188);
nand U44023 (N_44023,N_43411,N_43840);
xnor U44024 (N_44024,N_43135,N_42530);
xor U44025 (N_44025,N_42740,N_43637);
nand U44026 (N_44026,N_42160,N_42494);
and U44027 (N_44027,N_43098,N_42104);
nor U44028 (N_44028,N_43597,N_42349);
or U44029 (N_44029,N_43375,N_43404);
xnor U44030 (N_44030,N_43261,N_43250);
or U44031 (N_44031,N_42119,N_42438);
or U44032 (N_44032,N_43505,N_43417);
and U44033 (N_44033,N_42516,N_42457);
xor U44034 (N_44034,N_43644,N_43229);
nand U44035 (N_44035,N_43594,N_43685);
and U44036 (N_44036,N_43486,N_43665);
nand U44037 (N_44037,N_43465,N_42469);
or U44038 (N_44038,N_42419,N_42967);
or U44039 (N_44039,N_42869,N_43497);
or U44040 (N_44040,N_42619,N_42575);
nand U44041 (N_44041,N_42741,N_43139);
nor U44042 (N_44042,N_43120,N_42958);
and U44043 (N_44043,N_42341,N_42262);
nand U44044 (N_44044,N_42029,N_43580);
nor U44045 (N_44045,N_42235,N_43921);
xor U44046 (N_44046,N_43716,N_43033);
nor U44047 (N_44047,N_42243,N_43147);
xnor U44048 (N_44048,N_42892,N_42272);
and U44049 (N_44049,N_43630,N_43066);
or U44050 (N_44050,N_43177,N_43997);
or U44051 (N_44051,N_42055,N_43640);
nor U44052 (N_44052,N_42204,N_42284);
and U44053 (N_44053,N_42988,N_43232);
and U44054 (N_44054,N_42695,N_43845);
and U44055 (N_44055,N_42057,N_43557);
nand U44056 (N_44056,N_42944,N_42248);
and U44057 (N_44057,N_43308,N_43795);
nand U44058 (N_44058,N_43555,N_43687);
nor U44059 (N_44059,N_42350,N_43180);
nor U44060 (N_44060,N_43895,N_43208);
nor U44061 (N_44061,N_42835,N_42887);
and U44062 (N_44062,N_42717,N_43020);
xor U44063 (N_44063,N_42022,N_43325);
nand U44064 (N_44064,N_43953,N_42023);
or U44065 (N_44065,N_42543,N_43666);
or U44066 (N_44066,N_42616,N_42846);
xor U44067 (N_44067,N_43545,N_43859);
and U44068 (N_44068,N_42845,N_43893);
nor U44069 (N_44069,N_42377,N_43565);
and U44070 (N_44070,N_43461,N_43200);
and U44071 (N_44071,N_42808,N_42586);
nand U44072 (N_44072,N_42482,N_43590);
xnor U44073 (N_44073,N_43045,N_43276);
or U44074 (N_44074,N_42965,N_42780);
nor U44075 (N_44075,N_43605,N_43056);
or U44076 (N_44076,N_43781,N_43560);
xor U44077 (N_44077,N_43937,N_42885);
and U44078 (N_44078,N_43544,N_42148);
nor U44079 (N_44079,N_43986,N_43549);
and U44080 (N_44080,N_42224,N_42982);
nand U44081 (N_44081,N_43538,N_42355);
nor U44082 (N_44082,N_43962,N_42607);
nand U44083 (N_44083,N_43492,N_42767);
nor U44084 (N_44084,N_42134,N_43998);
nand U44085 (N_44085,N_43889,N_42822);
xor U44086 (N_44086,N_42827,N_43430);
xnor U44087 (N_44087,N_43679,N_43697);
and U44088 (N_44088,N_43936,N_43743);
and U44089 (N_44089,N_43132,N_42283);
nor U44090 (N_44090,N_43927,N_42612);
and U44091 (N_44091,N_43830,N_43625);
nor U44092 (N_44092,N_43851,N_43803);
and U44093 (N_44093,N_43439,N_43429);
nand U44094 (N_44094,N_42901,N_43246);
or U44095 (N_44095,N_42477,N_43019);
or U44096 (N_44096,N_43365,N_43788);
nand U44097 (N_44097,N_43829,N_43877);
and U44098 (N_44098,N_43703,N_43143);
nor U44099 (N_44099,N_43535,N_43919);
nand U44100 (N_44100,N_42044,N_42598);
xnor U44101 (N_44101,N_43736,N_42026);
nor U44102 (N_44102,N_43901,N_43073);
nand U44103 (N_44103,N_43293,N_43582);
and U44104 (N_44104,N_42862,N_43519);
nand U44105 (N_44105,N_43612,N_43427);
nor U44106 (N_44106,N_42095,N_42094);
and U44107 (N_44107,N_43756,N_43265);
nand U44108 (N_44108,N_43052,N_43446);
xnor U44109 (N_44109,N_42990,N_42589);
or U44110 (N_44110,N_43623,N_42042);
nor U44111 (N_44111,N_43190,N_43213);
nor U44112 (N_44112,N_42445,N_42207);
nor U44113 (N_44113,N_42604,N_43797);
and U44114 (N_44114,N_42132,N_42289);
xor U44115 (N_44115,N_43347,N_43498);
nand U44116 (N_44116,N_43267,N_42868);
and U44117 (N_44117,N_42972,N_42379);
and U44118 (N_44118,N_43682,N_43460);
and U44119 (N_44119,N_43546,N_43882);
and U44120 (N_44120,N_43035,N_42410);
or U44121 (N_44121,N_43448,N_42194);
nor U44122 (N_44122,N_43271,N_42215);
and U44123 (N_44123,N_42680,N_43346);
xnor U44124 (N_44124,N_42246,N_42101);
nor U44125 (N_44125,N_43233,N_43214);
and U44126 (N_44126,N_43536,N_43332);
and U44127 (N_44127,N_43494,N_43686);
nor U44128 (N_44128,N_43857,N_43802);
and U44129 (N_44129,N_42781,N_42193);
or U44130 (N_44130,N_42713,N_43945);
nand U44131 (N_44131,N_42709,N_42858);
xnor U44132 (N_44132,N_42444,N_43202);
and U44133 (N_44133,N_43616,N_43632);
or U44134 (N_44134,N_43504,N_42345);
nor U44135 (N_44135,N_42925,N_42070);
nor U44136 (N_44136,N_42314,N_42150);
nor U44137 (N_44137,N_42963,N_42926);
xnor U44138 (N_44138,N_43678,N_42113);
and U44139 (N_44139,N_43279,N_43885);
xnor U44140 (N_44140,N_43022,N_42368);
and U44141 (N_44141,N_43138,N_42398);
nor U44142 (N_44142,N_43469,N_42447);
or U44143 (N_44143,N_42841,N_42127);
nor U44144 (N_44144,N_42499,N_42359);
xnor U44145 (N_44145,N_42508,N_42692);
xor U44146 (N_44146,N_43617,N_43776);
nand U44147 (N_44147,N_42242,N_43185);
or U44148 (N_44148,N_42613,N_43615);
or U44149 (N_44149,N_43345,N_43244);
nor U44150 (N_44150,N_42642,N_42372);
nor U44151 (N_44151,N_42573,N_42921);
or U44152 (N_44152,N_42747,N_42736);
and U44153 (N_44153,N_43521,N_42261);
nor U44154 (N_44154,N_43083,N_42665);
nor U44155 (N_44155,N_43051,N_42024);
nor U44156 (N_44156,N_43096,N_43161);
xnor U44157 (N_44157,N_43728,N_42959);
nor U44158 (N_44158,N_43146,N_43786);
and U44159 (N_44159,N_42899,N_43853);
nor U44160 (N_44160,N_42300,N_42125);
and U44161 (N_44161,N_42213,N_43892);
nor U44162 (N_44162,N_42080,N_43266);
nor U44163 (N_44163,N_43026,N_43210);
or U44164 (N_44164,N_42933,N_43760);
nor U44165 (N_44165,N_43558,N_42036);
xor U44166 (N_44166,N_43534,N_42673);
or U44167 (N_44167,N_43761,N_42567);
nand U44168 (N_44168,N_43916,N_42674);
or U44169 (N_44169,N_43330,N_42177);
and U44170 (N_44170,N_43248,N_43987);
nor U44171 (N_44171,N_43027,N_43993);
nor U44172 (N_44172,N_43217,N_43671);
xor U44173 (N_44173,N_43742,N_43262);
or U44174 (N_44174,N_43301,N_42249);
nand U44175 (N_44175,N_42762,N_42422);
xnor U44176 (N_44176,N_43194,N_43075);
nand U44177 (N_44177,N_42534,N_42800);
nor U44178 (N_44178,N_42323,N_42252);
xor U44179 (N_44179,N_42291,N_42545);
and U44180 (N_44180,N_42443,N_43974);
xor U44181 (N_44181,N_43110,N_43269);
nor U44182 (N_44182,N_43499,N_42253);
and U44183 (N_44183,N_43917,N_43516);
or U44184 (N_44184,N_42599,N_42299);
and U44185 (N_44185,N_42440,N_42946);
or U44186 (N_44186,N_42434,N_43991);
nand U44187 (N_44187,N_43394,N_42358);
nand U44188 (N_44188,N_43409,N_43981);
xnor U44189 (N_44189,N_42460,N_42608);
nand U44190 (N_44190,N_42495,N_42651);
and U44191 (N_44191,N_43924,N_42149);
nor U44192 (N_44192,N_43181,N_43136);
xnor U44193 (N_44193,N_43714,N_43285);
nand U44194 (N_44194,N_42656,N_43906);
xor U44195 (N_44195,N_42793,N_42819);
nor U44196 (N_44196,N_42784,N_42231);
and U44197 (N_44197,N_42511,N_43984);
nor U44198 (N_44198,N_43175,N_43350);
xnor U44199 (N_44199,N_42088,N_43996);
nand U44200 (N_44200,N_42049,N_42893);
xnor U44201 (N_44201,N_43137,N_42937);
xor U44202 (N_44202,N_43152,N_42244);
and U44203 (N_44203,N_42865,N_43782);
xnor U44204 (N_44204,N_43968,N_43774);
and U44205 (N_44205,N_43935,N_43176);
or U44206 (N_44206,N_42332,N_42572);
nand U44207 (N_44207,N_42518,N_42324);
or U44208 (N_44208,N_42704,N_43684);
or U44209 (N_44209,N_43903,N_42034);
nor U44210 (N_44210,N_43785,N_43282);
xnor U44211 (N_44211,N_43822,N_42075);
xnor U44212 (N_44212,N_43067,N_42334);
nand U44213 (N_44213,N_42484,N_42174);
and U44214 (N_44214,N_42128,N_42254);
and U44215 (N_44215,N_43408,N_43290);
and U44216 (N_44216,N_43807,N_42620);
nor U44217 (N_44217,N_43481,N_43057);
nand U44218 (N_44218,N_43995,N_43113);
xor U44219 (N_44219,N_43418,N_42617);
or U44220 (N_44220,N_42467,N_42752);
nand U44221 (N_44221,N_42542,N_42143);
nand U44222 (N_44222,N_43414,N_43746);
or U44223 (N_44223,N_42910,N_42165);
xor U44224 (N_44224,N_42896,N_42328);
xnor U44225 (N_44225,N_43435,N_42742);
nand U44226 (N_44226,N_42843,N_42754);
or U44227 (N_44227,N_43734,N_43681);
or U44228 (N_44228,N_43127,N_43541);
xor U44229 (N_44229,N_42370,N_42592);
or U44230 (N_44230,N_42900,N_43032);
xor U44231 (N_44231,N_43741,N_42367);
and U44232 (N_44232,N_42681,N_43235);
or U44233 (N_44233,N_43046,N_42090);
nand U44234 (N_44234,N_43596,N_43303);
or U44235 (N_44235,N_42924,N_43828);
nor U44236 (N_44236,N_42158,N_42319);
or U44237 (N_44237,N_42942,N_42428);
and U44238 (N_44238,N_43971,N_43377);
and U44239 (N_44239,N_43356,N_43798);
and U44240 (N_44240,N_42792,N_43664);
and U44241 (N_44241,N_43431,N_42219);
nand U44242 (N_44242,N_43989,N_43297);
nor U44243 (N_44243,N_42371,N_42473);
or U44244 (N_44244,N_43900,N_42555);
nand U44245 (N_44245,N_42363,N_43698);
and U44246 (N_44246,N_43854,N_42072);
nand U44247 (N_44247,N_43361,N_43566);
nand U44248 (N_44248,N_42954,N_42048);
nand U44249 (N_44249,N_43820,N_43349);
nand U44250 (N_44250,N_43328,N_43378);
or U44251 (N_44251,N_42668,N_43309);
nor U44252 (N_44252,N_43529,N_43362);
nand U44253 (N_44253,N_42050,N_42820);
xor U44254 (N_44254,N_43815,N_42003);
nand U44255 (N_44255,N_43500,N_42979);
and U44256 (N_44256,N_42645,N_42031);
nand U44257 (N_44257,N_42353,N_42821);
or U44258 (N_44258,N_43286,N_42487);
nor U44259 (N_44259,N_42774,N_43539);
nand U44260 (N_44260,N_43256,N_42514);
and U44261 (N_44261,N_43704,N_42977);
and U44262 (N_44262,N_43562,N_42533);
or U44263 (N_44263,N_43488,N_42163);
xnor U44264 (N_44264,N_43826,N_43072);
nor U44265 (N_44265,N_42015,N_43204);
xor U44266 (N_44266,N_42590,N_42804);
and U44267 (N_44267,N_42333,N_42585);
and U44268 (N_44268,N_42331,N_42888);
nor U44269 (N_44269,N_43321,N_42768);
nand U44270 (N_44270,N_42987,N_42994);
or U44271 (N_44271,N_43334,N_43197);
nor U44272 (N_44272,N_43359,N_43972);
or U44273 (N_44273,N_43095,N_42124);
or U44274 (N_44274,N_43241,N_43249);
nor U44275 (N_44275,N_43201,N_43568);
xnor U44276 (N_44276,N_43653,N_42907);
nand U44277 (N_44277,N_42200,N_43193);
and U44278 (N_44278,N_43485,N_43683);
and U44279 (N_44279,N_42810,N_43852);
nand U44280 (N_44280,N_43578,N_42574);
xor U44281 (N_44281,N_42288,N_42920);
and U44282 (N_44282,N_42004,N_42971);
and U44283 (N_44283,N_43865,N_43753);
xor U44284 (N_44284,N_42527,N_42303);
and U44285 (N_44285,N_43124,N_42690);
and U44286 (N_44286,N_42021,N_42632);
nand U44287 (N_44287,N_43647,N_42989);
or U44288 (N_44288,N_43457,N_42505);
nor U44289 (N_44289,N_42212,N_43940);
xor U44290 (N_44290,N_42884,N_43754);
nand U44291 (N_44291,N_42337,N_42571);
and U44292 (N_44292,N_43473,N_42292);
nor U44293 (N_44293,N_43357,N_42639);
nor U44294 (N_44294,N_42156,N_43164);
xnor U44295 (N_44295,N_42995,N_42582);
nand U44296 (N_44296,N_43367,N_43078);
or U44297 (N_44297,N_42818,N_43061);
or U44298 (N_44298,N_42797,N_43070);
nor U44299 (N_44299,N_42923,N_43341);
nor U44300 (N_44300,N_42264,N_43182);
nor U44301 (N_44301,N_43456,N_43455);
nand U44302 (N_44302,N_43107,N_43733);
and U44303 (N_44303,N_43231,N_42698);
nand U44304 (N_44304,N_42257,N_42622);
xor U44305 (N_44305,N_43844,N_43421);
xnor U44306 (N_44306,N_42828,N_42952);
nor U44307 (N_44307,N_42114,N_43978);
nor U44308 (N_44308,N_42276,N_43886);
and U44309 (N_44309,N_43620,N_43042);
nand U44310 (N_44310,N_42111,N_43926);
nor U44311 (N_44311,N_43464,N_43514);
nor U44312 (N_44312,N_42975,N_43482);
xnor U44313 (N_44313,N_42362,N_43012);
nand U44314 (N_44314,N_42435,N_43543);
nor U44315 (N_44315,N_42402,N_43272);
or U44316 (N_44316,N_42385,N_42138);
nor U44317 (N_44317,N_42964,N_42556);
nor U44318 (N_44318,N_42222,N_42208);
xnor U44319 (N_44319,N_42882,N_42730);
or U44320 (N_44320,N_43530,N_43619);
nor U44321 (N_44321,N_43510,N_43914);
or U44322 (N_44322,N_43125,N_42285);
or U44323 (N_44323,N_43478,N_43077);
nand U44324 (N_44324,N_42553,N_43260);
xnor U44325 (N_44325,N_42255,N_42183);
and U44326 (N_44326,N_43097,N_43988);
xnor U44327 (N_44327,N_43352,N_43651);
and U44328 (N_44328,N_42318,N_42356);
xnor U44329 (N_44329,N_43982,N_42738);
or U44330 (N_44330,N_42504,N_42525);
and U44331 (N_44331,N_43451,N_42197);
nand U44332 (N_44332,N_42378,N_42439);
nand U44333 (N_44333,N_43058,N_43099);
nand U44334 (N_44334,N_43159,N_43639);
or U44335 (N_44335,N_42547,N_42293);
and U44336 (N_44336,N_43192,N_43419);
and U44337 (N_44337,N_42190,N_42678);
and U44338 (N_44338,N_43842,N_42464);
and U44339 (N_44339,N_42198,N_43129);
nor U44340 (N_44340,N_42703,N_42169);
xnor U44341 (N_44341,N_43501,N_43720);
and U44342 (N_44342,N_43735,N_43677);
nor U44343 (N_44343,N_43230,N_43818);
nand U44344 (N_44344,N_42961,N_43021);
xnor U44345 (N_44345,N_42426,N_42765);
nand U44346 (N_44346,N_43385,N_42192);
or U44347 (N_44347,N_43918,N_43879);
nand U44348 (N_44348,N_42453,N_43205);
nor U44349 (N_44349,N_42915,N_42548);
nand U44350 (N_44350,N_43874,N_42528);
or U44351 (N_44351,N_42798,N_42305);
nor U44352 (N_44352,N_43477,N_42146);
and U44353 (N_44353,N_42463,N_43384);
xor U44354 (N_44354,N_42479,N_42100);
or U44355 (N_44355,N_42459,N_42315);
and U44356 (N_44356,N_42306,N_43695);
nand U44357 (N_44357,N_42561,N_42834);
or U44358 (N_44358,N_42056,N_42233);
or U44359 (N_44359,N_43858,N_42178);
nor U44360 (N_44360,N_42629,N_43283);
or U44361 (N_44361,N_43721,N_42700);
xnor U44362 (N_44362,N_43581,N_42316);
nand U44363 (N_44363,N_43115,N_43775);
and U44364 (N_44364,N_42610,N_43295);
nand U44365 (N_44365,N_42596,N_42140);
and U44366 (N_44366,N_43080,N_42170);
or U44367 (N_44367,N_43897,N_43976);
or U44368 (N_44368,N_43891,N_42570);
xor U44369 (N_44369,N_43709,N_43353);
nand U44370 (N_44370,N_42559,N_42809);
nand U44371 (N_44371,N_43471,N_42455);
xnor U44372 (N_44372,N_43824,N_43081);
nand U44373 (N_44373,N_42636,N_42664);
and U44374 (N_44374,N_42646,N_43225);
nand U44375 (N_44375,N_43195,N_42701);
nand U44376 (N_44376,N_42092,N_42702);
xnor U44377 (N_44377,N_43873,N_43397);
and U44378 (N_44378,N_43794,N_42856);
or U44379 (N_44379,N_43827,N_42129);
and U44380 (N_44380,N_42405,N_43843);
nor U44381 (N_44381,N_43944,N_42311);
nor U44382 (N_44382,N_42714,N_43575);
nand U44383 (N_44383,N_42870,N_43314);
or U44384 (N_44384,N_42181,N_43253);
or U44385 (N_44385,N_42205,N_42945);
and U44386 (N_44386,N_42273,N_43750);
and U44387 (N_44387,N_43730,N_43258);
or U44388 (N_44388,N_42040,N_43871);
nand U44389 (N_44389,N_43383,N_43688);
nor U44390 (N_44390,N_42223,N_42019);
xnor U44391 (N_44391,N_43329,N_43731);
and U44392 (N_44392,N_42670,N_42878);
nand U44393 (N_44393,N_42427,N_42853);
and U44394 (N_44394,N_43388,N_43793);
xor U44395 (N_44395,N_43315,N_42773);
and U44396 (N_44396,N_42594,N_43317);
xnor U44397 (N_44397,N_43662,N_43778);
nand U44398 (N_44398,N_42634,N_42451);
nand U44399 (N_44399,N_42551,N_42118);
xor U44400 (N_44400,N_43445,N_42325);
or U44401 (N_44401,N_43729,N_42776);
nand U44402 (N_44402,N_43273,N_43866);
or U44403 (N_44403,N_43128,N_43727);
nor U44404 (N_44404,N_42013,N_42338);
nand U44405 (N_44405,N_42322,N_42297);
nand U44406 (N_44406,N_43779,N_43509);
and U44407 (N_44407,N_42855,N_43219);
or U44408 (N_44408,N_42602,N_43173);
nor U44409 (N_44409,N_42580,N_42562);
nand U44410 (N_44410,N_42010,N_43552);
or U44411 (N_44411,N_42833,N_42541);
or U44412 (N_44412,N_43635,N_42201);
or U44413 (N_44413,N_42799,N_42756);
and U44414 (N_44414,N_43627,N_43186);
and U44415 (N_44415,N_42109,N_42184);
or U44416 (N_44416,N_43863,N_43592);
and U44417 (N_44417,N_43236,N_43490);
xnor U44418 (N_44418,N_43354,N_43207);
nor U44419 (N_44419,N_42941,N_43442);
nand U44420 (N_44420,N_42568,N_43513);
nor U44421 (N_44421,N_42006,N_42918);
nor U44422 (N_44422,N_43119,N_43480);
or U44423 (N_44423,N_42018,N_43992);
and U44424 (N_44424,N_42448,N_42860);
and U44425 (N_44425,N_42653,N_42815);
and U44426 (N_44426,N_42716,N_43013);
nand U44427 (N_44427,N_43031,N_42761);
xor U44428 (N_44428,N_43564,N_43368);
nand U44429 (N_44429,N_42051,N_43340);
and U44430 (N_44430,N_43495,N_43673);
nor U44431 (N_44431,N_43642,N_42216);
nand U44432 (N_44432,N_43018,N_42106);
xor U44433 (N_44433,N_42421,N_43343);
and U44434 (N_44434,N_43306,N_42817);
or U44435 (N_44435,N_42310,N_43668);
and U44436 (N_44436,N_42476,N_42641);
and U44437 (N_44437,N_43930,N_43449);
xor U44438 (N_44438,N_42515,N_42521);
or U44439 (N_44439,N_43811,N_42097);
nand U44440 (N_44440,N_43294,N_42507);
or U44441 (N_44441,N_42063,N_43327);
xor U44442 (N_44442,N_42266,N_43551);
nand U44443 (N_44443,N_43772,N_43239);
nor U44444 (N_44444,N_42232,N_42241);
and U44445 (N_44445,N_43890,N_43015);
and U44446 (N_44446,N_43082,N_42226);
nor U44447 (N_44447,N_43121,N_42258);
nor U44448 (N_44448,N_43108,N_42711);
nor U44449 (N_44449,N_42857,N_42526);
or U44450 (N_44450,N_43787,N_42456);
nor U44451 (N_44451,N_43382,N_43792);
nor U44452 (N_44452,N_42693,N_43748);
nor U44453 (N_44453,N_42011,N_43739);
xor U44454 (N_44454,N_43812,N_42795);
or U44455 (N_44455,N_43006,N_43595);
nand U44456 (N_44456,N_43037,N_42308);
and U44457 (N_44457,N_43255,N_43215);
xnor U44458 (N_44458,N_43715,N_43363);
xor U44459 (N_44459,N_43932,N_42116);
or U44460 (N_44460,N_43422,N_43089);
nor U44461 (N_44461,N_43718,N_42850);
nand U44462 (N_44462,N_43305,N_42352);
and U44463 (N_44463,N_42247,N_43878);
xnor U44464 (N_44464,N_43512,N_43613);
xor U44465 (N_44465,N_42005,N_43628);
nand U44466 (N_44466,N_43360,N_43508);
nor U44467 (N_44467,N_43770,N_42624);
xnor U44468 (N_44468,N_42579,N_43607);
or U44469 (N_44469,N_42191,N_43403);
and U44470 (N_44470,N_42278,N_43039);
nor U44471 (N_44471,N_42577,N_42060);
xor U44472 (N_44472,N_42836,N_42986);
nand U44473 (N_44473,N_42640,N_43206);
or U44474 (N_44474,N_42722,N_43453);
nor U44475 (N_44475,N_43894,N_43064);
xor U44476 (N_44476,N_42844,N_43708);
nand U44477 (N_44477,N_43980,N_42446);
xnor U44478 (N_44478,N_43040,N_42423);
nand U44479 (N_44479,N_42847,N_43771);
nor U44480 (N_44480,N_42108,N_42729);
xnor U44481 (N_44481,N_42218,N_43216);
nand U44482 (N_44482,N_42911,N_42466);
and U44483 (N_44483,N_43973,N_42211);
xor U44484 (N_44484,N_42563,N_43977);
or U44485 (N_44485,N_42472,N_43724);
or U44486 (N_44486,N_42864,N_42993);
or U44487 (N_44487,N_43157,N_43209);
xnor U44488 (N_44488,N_43983,N_43007);
nor U44489 (N_44489,N_42153,N_42852);
nand U44490 (N_44490,N_43570,N_42529);
nor U44491 (N_44491,N_42744,N_43657);
xor U44492 (N_44492,N_43148,N_42009);
nand U44493 (N_44493,N_42807,N_42260);
nor U44494 (N_44494,N_43010,N_42644);
nor U44495 (N_44495,N_43302,N_43841);
or U44496 (N_44496,N_43810,N_42032);
and U44497 (N_44497,N_43909,N_43904);
nor U44498 (N_44498,N_42889,N_43050);
and U44499 (N_44499,N_43416,N_42837);
nor U44500 (N_44500,N_43319,N_42386);
xor U44501 (N_44501,N_43949,N_43846);
nor U44502 (N_44502,N_42155,N_43626);
nor U44503 (N_44503,N_43963,N_43548);
or U44504 (N_44504,N_42643,N_43379);
xor U44505 (N_44505,N_43313,N_43275);
xnor U44506 (N_44506,N_42185,N_42470);
nor U44507 (N_44507,N_43447,N_43483);
nand U44508 (N_44508,N_43355,N_42152);
or U44509 (N_44509,N_43929,N_43079);
and U44510 (N_44510,N_42688,N_42718);
xor U44511 (N_44511,N_43268,N_43351);
and U44512 (N_44512,N_43090,N_43369);
and U44513 (N_44513,N_43034,N_42825);
nor U44514 (N_44514,N_42001,N_43410);
and U44515 (N_44515,N_42073,N_42803);
xor U44516 (N_44516,N_42007,N_43910);
nor U44517 (N_44517,N_42652,N_42710);
or U44518 (N_44518,N_42531,N_43187);
or U44519 (N_44519,N_43436,N_43780);
nor U44520 (N_44520,N_43141,N_42550);
nand U44521 (N_44521,N_43044,N_42814);
nand U44522 (N_44522,N_42102,N_43835);
xor U44523 (N_44523,N_43624,N_42298);
and U44524 (N_44524,N_43069,N_42905);
xnor U44525 (N_44525,N_42491,N_43970);
nor U44526 (N_44526,N_43946,N_43813);
nor U44527 (N_44527,N_43462,N_42801);
nor U44528 (N_44528,N_42361,N_42749);
and U44529 (N_44529,N_43170,N_43629);
nor U44530 (N_44530,N_43868,N_43598);
or U44531 (N_44531,N_42832,N_42560);
and U44532 (N_44532,N_42842,N_42949);
and U44533 (N_44533,N_43799,N_43593);
nand U44534 (N_44534,N_42676,N_43773);
nor U44535 (N_44535,N_43610,N_43413);
nor U44536 (N_44536,N_42829,N_42347);
nor U44537 (N_44537,N_42960,N_43693);
and U44538 (N_44538,N_42256,N_42983);
nand U44539 (N_44539,N_42112,N_42764);
xnor U44540 (N_44540,N_43339,N_43676);
nor U44541 (N_44541,N_43109,N_43958);
nor U44542 (N_44542,N_43169,N_42161);
or U44543 (N_44543,N_43608,N_42301);
nor U44544 (N_44544,N_42658,N_43459);
or U44545 (N_44545,N_43862,N_43062);
nand U44546 (N_44546,N_43669,N_42603);
and U44547 (N_44547,N_43226,N_43084);
nand U44548 (N_44548,N_42336,N_42390);
nand U44549 (N_44549,N_42538,N_42727);
xnor U44550 (N_44550,N_43747,N_42461);
nand U44551 (N_44551,N_43985,N_42724);
or U44552 (N_44552,N_42339,N_42290);
nor U44553 (N_44553,N_43001,N_43621);
xnor U44554 (N_44554,N_42766,N_42707);
nand U44555 (N_44555,N_43875,N_43614);
nor U44556 (N_44556,N_43049,N_42330);
nand U44557 (N_44557,N_43100,N_42916);
or U44558 (N_44558,N_43587,N_43837);
xnor U44559 (N_44559,N_42823,N_42880);
and U44560 (N_44560,N_43719,N_42745);
or U44561 (N_44561,N_42131,N_42045);
and U44562 (N_44562,N_43165,N_43130);
nand U44563 (N_44563,N_42873,N_43405);
xor U44564 (N_44564,N_43094,N_42351);
nand U44565 (N_44565,N_43415,N_43550);
nor U44566 (N_44566,N_42633,N_42566);
or U44567 (N_44567,N_42110,N_43705);
nor U44568 (N_44568,N_43423,N_42180);
nor U44569 (N_44569,N_42903,N_42731);
and U44570 (N_44570,N_42203,N_42406);
or U44571 (N_44571,N_43101,N_42601);
nand U44572 (N_44572,N_43024,N_43116);
nor U44573 (N_44573,N_42522,N_42008);
nor U44574 (N_44574,N_42712,N_43689);
or U44575 (N_44575,N_43563,N_42931);
or U44576 (N_44576,N_43133,N_42087);
xnor U44577 (N_44577,N_43398,N_42121);
and U44578 (N_44578,N_43104,N_42279);
or U44579 (N_44579,N_43864,N_42867);
and U44580 (N_44580,N_42493,N_42265);
or U44581 (N_44581,N_43470,N_43554);
xnor U44582 (N_44582,N_43331,N_43196);
or U44583 (N_44583,N_42984,N_42043);
nor U44584 (N_44584,N_42966,N_42955);
nor U44585 (N_44585,N_42512,N_42997);
xor U44586 (N_44586,N_43922,N_42917);
nor U44587 (N_44587,N_43376,N_42416);
xnor U44588 (N_44588,N_42411,N_43913);
and U44589 (N_44589,N_42117,N_43299);
nor U44590 (N_44590,N_43712,N_42786);
or U44591 (N_44591,N_43725,N_43491);
nor U44592 (N_44592,N_42628,N_43783);
xor U44593 (N_44593,N_42431,N_43433);
or U44594 (N_44594,N_42520,N_43573);
nand U44595 (N_44595,N_42228,N_42759);
or U44596 (N_44596,N_42879,N_42471);
or U44597 (N_44597,N_42544,N_42947);
nor U44598 (N_44598,N_43053,N_43584);
nand U44599 (N_44599,N_42430,N_42886);
or U44600 (N_44600,N_43652,N_43452);
and U44601 (N_44601,N_43126,N_42849);
xor U44602 (N_44602,N_42609,N_43140);
xor U44603 (N_44603,N_43591,N_42839);
and U44604 (N_44604,N_43713,N_43819);
or U44605 (N_44605,N_42875,N_43428);
xnor U44606 (N_44606,N_43322,N_42763);
nand U44607 (N_44607,N_43280,N_42501);
nand U44608 (N_44608,N_43221,N_43752);
xor U44609 (N_44609,N_43680,N_43387);
nor U44610 (N_44610,N_43659,N_43373);
nor U44611 (N_44611,N_43257,N_43738);
nor U44612 (N_44612,N_42771,N_42951);
xnor U44613 (N_44613,N_42195,N_42980);
and U44614 (N_44614,N_43335,N_43645);
nor U44615 (N_44615,N_43732,N_42891);
xnor U44616 (N_44616,N_42139,N_42675);
or U44617 (N_44617,N_42872,N_43825);
and U44618 (N_44618,N_43395,N_43412);
nor U44619 (N_44619,N_42250,N_42969);
xor U44620 (N_44620,N_42535,N_42654);
xor U44621 (N_44621,N_43211,N_43479);
or U44622 (N_44622,N_42237,N_43956);
nor U44623 (N_44623,N_42490,N_42953);
or U44624 (N_44624,N_42565,N_43304);
and U44625 (N_44625,N_43540,N_43005);
nand U44626 (N_44626,N_43234,N_42778);
or U44627 (N_44627,N_42239,N_42392);
nand U44628 (N_44628,N_43333,N_43528);
and U44629 (N_44629,N_42912,N_43518);
nor U44630 (N_44630,N_43284,N_43307);
nand U44631 (N_44631,N_42605,N_43142);
nor U44632 (N_44632,N_43223,N_42523);
and U44633 (N_44633,N_42666,N_43650);
nor U44634 (N_44634,N_42957,N_43931);
nor U44635 (N_44635,N_43008,N_42806);
nor U44636 (N_44636,N_42162,N_43951);
or U44637 (N_44637,N_42376,N_43074);
or U44638 (N_44638,N_43943,N_43432);
xor U44639 (N_44639,N_43336,N_43547);
nand U44640 (N_44640,N_42973,N_43183);
or U44641 (N_44641,N_43999,N_42267);
xor U44642 (N_44642,N_43723,N_42492);
and U44643 (N_44643,N_43264,N_42627);
or U44644 (N_44644,N_42304,N_43524);
nand U44645 (N_44645,N_43150,N_42757);
or U44646 (N_44646,N_42166,N_42655);
nor U44647 (N_44647,N_42569,N_43749);
nand U44648 (N_44648,N_43532,N_43762);
and U44649 (N_44649,N_43661,N_42769);
or U44650 (N_44650,N_42626,N_43338);
nor U44651 (N_44651,N_43179,N_42269);
and U44652 (N_44652,N_42238,N_43805);
nor U44653 (N_44653,N_43898,N_43961);
nor U44654 (N_44654,N_43699,N_43117);
nand U44655 (N_44655,N_42576,N_42326);
nand U44656 (N_44656,N_42475,N_43274);
and U44657 (N_44657,N_42047,N_43242);
xnor U44658 (N_44658,N_42375,N_43441);
xor U44659 (N_44659,N_43526,N_42136);
nand U44660 (N_44660,N_43870,N_42630);
nor U44661 (N_44661,N_43579,N_42739);
nand U44662 (N_44662,N_42234,N_43817);
nor U44663 (N_44663,N_42442,N_43833);
and U44664 (N_44664,N_42017,N_42142);
and U44665 (N_44665,N_43601,N_43472);
and U44666 (N_44666,N_43667,N_42928);
nand U44667 (N_44667,N_42122,N_43804);
nand U44668 (N_44668,N_43649,N_42851);
and U44669 (N_44669,N_43466,N_42016);
nand U44670 (N_44670,N_42179,N_42581);
nand U44671 (N_44671,N_42236,N_42760);
or U44672 (N_44672,N_42826,N_42513);
xor U44673 (N_44673,N_43086,N_43888);
nor U44674 (N_44674,N_42648,N_43401);
xor U44675 (N_44675,N_43806,N_42755);
xor U44676 (N_44676,N_42830,N_42098);
nor U44677 (N_44677,N_43358,N_43967);
or U44678 (N_44678,N_42898,N_43939);
or U44679 (N_44679,N_43312,N_43118);
and U44680 (N_44680,N_43836,N_43298);
and U44681 (N_44681,N_42229,N_42327);
nor U44682 (N_44682,N_42282,N_42066);
xnor U44683 (N_44683,N_43292,N_43496);
xor U44684 (N_44684,N_42425,N_42486);
nor U44685 (N_44685,N_43849,N_42071);
and U44686 (N_44686,N_43571,N_43757);
nor U44687 (N_44687,N_43281,N_43744);
or U44688 (N_44688,N_43691,N_42182);
or U44689 (N_44689,N_43531,N_43002);
or U44690 (N_44690,N_42274,N_42396);
and U44691 (N_44691,N_42081,N_42144);
xor U44692 (N_44692,N_43426,N_43252);
nand U44693 (N_44693,N_42578,N_43561);
nand U44694 (N_44694,N_43839,N_43717);
xor U44695 (N_44695,N_42751,N_42307);
nor U44696 (N_44696,N_42120,N_43320);
or U44697 (N_44697,N_42999,N_43288);
nand U44698 (N_44698,N_43392,N_43212);
nand U44699 (N_44699,N_42357,N_42956);
nor U44700 (N_44700,N_43572,N_43867);
nand U44701 (N_44701,N_43950,N_42746);
xnor U44702 (N_44702,N_43694,N_43278);
or U44703 (N_44703,N_42588,N_42014);
nor U44704 (N_44704,N_43092,N_43636);
or U44705 (N_44705,N_43861,N_43696);
nor U44706 (N_44706,N_43706,N_42489);
xnor U44707 (N_44707,N_43153,N_43149);
xor U44708 (N_44708,N_43172,N_42078);
nor U44709 (N_44709,N_42726,N_43816);
or U44710 (N_44710,N_43237,N_42805);
nor U44711 (N_44711,N_42432,N_42913);
xnor U44712 (N_44712,N_43990,N_43933);
or U44713 (N_44713,N_43583,N_42217);
nor U44714 (N_44714,N_42342,N_42039);
or U44715 (N_44715,N_42465,N_42052);
xnor U44716 (N_44716,N_42998,N_43767);
nand U44717 (N_44717,N_42772,N_43609);
or U44718 (N_44718,N_43556,N_42313);
and U44719 (N_44719,N_42939,N_43850);
xor U44720 (N_44720,N_42074,N_42468);
xnor U44721 (N_44721,N_42922,N_42481);
or U44722 (N_44722,N_42991,N_43502);
and U44723 (N_44723,N_43618,N_42859);
or U44724 (N_44724,N_43487,N_42783);
nand U44725 (N_44725,N_42059,N_42686);
xor U44726 (N_44726,N_42871,N_42414);
nand U44727 (N_44727,N_43574,N_43527);
nor U44728 (N_44728,N_42159,N_43658);
and U44729 (N_44729,N_42395,N_43957);
or U44730 (N_44730,N_43484,N_43199);
xor U44731 (N_44731,N_42697,N_43054);
nor U44732 (N_44732,N_43604,N_42202);
nand U44733 (N_44733,N_43954,N_42344);
nor U44734 (N_44734,N_42382,N_43576);
and U44735 (N_44735,N_43425,N_43220);
and U44736 (N_44736,N_43654,N_42597);
nand U44737 (N_44737,N_43396,N_42412);
or U44738 (N_44738,N_43174,N_42758);
nor U44739 (N_44739,N_42976,N_42962);
nand U44740 (N_44740,N_42611,N_43160);
nor U44741 (N_44741,N_43737,N_42894);
xnor U44742 (N_44742,N_42096,N_43243);
and U44743 (N_44743,N_43198,N_43821);
nand U44744 (N_44744,N_42187,N_43263);
and U44745 (N_44745,N_42787,N_42275);
nand U44746 (N_44746,N_43443,N_43122);
or U44747 (N_44747,N_43523,N_42329);
or U44748 (N_44748,N_42638,N_42948);
nor U44749 (N_44749,N_43745,N_42683);
nor U44750 (N_44750,N_43155,N_42794);
and U44751 (N_44751,N_43902,N_43048);
nand U44752 (N_44752,N_43337,N_42950);
nor U44753 (N_44753,N_43003,N_43758);
nand U44754 (N_44754,N_42206,N_42631);
and U44755 (N_44755,N_43701,N_42788);
and U44756 (N_44756,N_43191,N_43131);
nor U44757 (N_44757,N_42287,N_43386);
nor U44758 (N_44758,N_43111,N_42245);
nand U44759 (N_44759,N_43085,N_42775);
xor U44760 (N_44760,N_43768,N_42436);
xor U44761 (N_44761,N_42420,N_42320);
xnor U44762 (N_44762,N_43400,N_42785);
nand U44763 (N_44763,N_42408,N_43872);
and U44764 (N_44764,N_43920,N_43114);
xnor U44765 (N_44765,N_42554,N_43289);
nor U44766 (N_44766,N_43043,N_43088);
xor U44767 (N_44767,N_43569,N_42615);
nor U44768 (N_44768,N_43847,N_42354);
xor U44769 (N_44769,N_43151,N_43326);
or U44770 (N_44770,N_43751,N_42225);
xnor U44771 (N_44771,N_42777,N_42861);
or U44772 (N_44772,N_43876,N_43489);
nor U44773 (N_44773,N_43162,N_42719);
and U44774 (N_44774,N_43764,N_42263);
xnor U44775 (N_44775,N_43222,N_43218);
or U44776 (N_44776,N_43203,N_42417);
nand U44777 (N_44777,N_43600,N_43577);
or U44778 (N_44778,N_43517,N_42064);
and U44779 (N_44779,N_43450,N_43655);
or U44780 (N_44780,N_42037,N_42524);
nand U44781 (N_44781,N_42546,N_42904);
nand U44782 (N_44782,N_42210,N_43777);
nand U44783 (N_44783,N_43674,N_42220);
or U44784 (N_44784,N_42929,N_42661);
and U44785 (N_44785,N_42485,N_42635);
and U44786 (N_44786,N_42696,N_43144);
or U44787 (N_44787,N_43270,N_42068);
xor U44788 (N_44788,N_42789,N_43036);
or U44789 (N_44789,N_42141,N_42147);
or U44790 (N_44790,N_43960,N_43028);
nor U44791 (N_44791,N_42813,N_42046);
and U44792 (N_44792,N_43184,N_42373);
or U44793 (N_44793,N_42076,N_43784);
nor U44794 (N_44794,N_42462,N_42895);
nand U44795 (N_44795,N_42970,N_42286);
nand U44796 (N_44796,N_42227,N_42902);
or U44797 (N_44797,N_43896,N_42743);
nand U44798 (N_44798,N_42115,N_43881);
xnor U44799 (N_44799,N_43938,N_43634);
nand U44800 (N_44800,N_42732,N_42020);
nor U44801 (N_44801,N_42591,N_42424);
and U44802 (N_44802,N_42725,N_42312);
or U44803 (N_44803,N_42812,N_43511);
nand U44804 (N_44804,N_42908,N_43145);
nor U44805 (N_44805,N_42552,N_43171);
or U44806 (N_44806,N_42816,N_43801);
nand U44807 (N_44807,N_43966,N_42171);
nor U44808 (N_44808,N_42909,N_42897);
nand U44809 (N_44809,N_42478,N_42335);
nand U44810 (N_44810,N_42103,N_43158);
nand U44811 (N_44811,N_42667,N_42369);
and U44812 (N_44812,N_43522,N_42519);
xnor U44813 (N_44813,N_42280,N_42606);
xnor U44814 (N_44814,N_43065,N_42397);
or U44815 (N_44815,N_42145,N_42906);
xnor U44816 (N_44816,N_43364,N_42883);
nand U44817 (N_44817,N_43759,N_42374);
or U44818 (N_44818,N_43323,N_42126);
or U44819 (N_44819,N_42557,N_42927);
or U44820 (N_44820,N_42404,N_43178);
and U44821 (N_44821,N_43156,N_43766);
and U44822 (N_44822,N_43047,N_43163);
and U44823 (N_44823,N_43586,N_43831);
nor U44824 (N_44824,N_42811,N_42025);
xnor U44825 (N_44825,N_43102,N_42474);
or U44826 (N_44826,N_42137,N_42992);
nand U44827 (N_44827,N_42085,N_43402);
nand U44828 (N_44828,N_43520,N_43030);
nor U44829 (N_44829,N_43438,N_42699);
nor U44830 (N_44830,N_42093,N_43648);
nand U44831 (N_44831,N_43493,N_42978);
xor U44832 (N_44832,N_43740,N_42536);
xnor U44833 (N_44833,N_43374,N_42506);
or U44834 (N_44834,N_42107,N_42863);
and U44835 (N_44835,N_42854,N_42660);
nor U44836 (N_44836,N_42295,N_42791);
nand U44837 (N_44837,N_42831,N_42671);
and U44838 (N_44838,N_42657,N_42723);
and U44839 (N_44839,N_43611,N_43112);
nand U44840 (N_44840,N_42038,N_43860);
nand U44841 (N_44841,N_42176,N_43646);
nor U44842 (N_44842,N_43189,N_43093);
xor U44843 (N_44843,N_42498,N_43641);
xor U44844 (N_44844,N_42943,N_42399);
nand U44845 (N_44845,N_42214,N_42084);
or U44846 (N_44846,N_42735,N_42600);
or U44847 (N_44847,N_43942,N_43672);
nand U44848 (N_44848,N_43103,N_43941);
or U44849 (N_44849,N_43515,N_42062);
nor U44850 (N_44850,N_42595,N_43925);
nor U44851 (N_44851,N_42230,N_42012);
nor U44852 (N_44852,N_42672,N_42391);
xor U44853 (N_44853,N_43559,N_42848);
nand U44854 (N_44854,N_42647,N_42454);
nand U44855 (N_44855,N_42079,N_42458);
nand U44856 (N_44856,N_42281,N_43855);
xnor U44857 (N_44857,N_43300,N_42360);
nor U44858 (N_44858,N_42750,N_42890);
nand U44859 (N_44859,N_42383,N_42277);
xor U44860 (N_44860,N_42089,N_42387);
or U44861 (N_44861,N_42091,N_42914);
xnor U44862 (N_44862,N_43588,N_43602);
and U44863 (N_44863,N_42687,N_43399);
nor U44864 (N_44864,N_43537,N_42403);
or U44865 (N_44865,N_43071,N_43475);
nand U44866 (N_44866,N_43259,N_42770);
and U44867 (N_44867,N_42623,N_42734);
and U44868 (N_44868,N_43154,N_42877);
xnor U44869 (N_44869,N_42940,N_42033);
nand U44870 (N_44870,N_43311,N_42824);
xnor U44871 (N_44871,N_42240,N_43440);
and U44872 (N_44872,N_42985,N_43004);
and U44873 (N_44873,N_42105,N_42981);
nor U44874 (N_44874,N_42366,N_42175);
and U44875 (N_44875,N_43928,N_42932);
nand U44876 (N_44876,N_43905,N_43660);
nor U44877 (N_44877,N_42167,N_43068);
and U44878 (N_44878,N_43907,N_43011);
xor U44879 (N_44879,N_43406,N_43391);
nor U44880 (N_44880,N_42413,N_43710);
nor U44881 (N_44881,N_42065,N_42689);
nor U44882 (N_44882,N_43123,N_42564);
nand U44883 (N_44883,N_43014,N_43979);
xnor U44884 (N_44884,N_42030,N_42720);
nor U44885 (N_44885,N_42866,N_42321);
xor U44886 (N_44886,N_43542,N_42168);
or U44887 (N_44887,N_43476,N_43167);
nand U44888 (N_44888,N_43808,N_42790);
xnor U44889 (N_44889,N_42679,N_42041);
nand U44890 (N_44890,N_42271,N_42593);
xnor U44891 (N_44891,N_42157,N_43454);
nand U44892 (N_44892,N_42388,N_42682);
xnor U44893 (N_44893,N_42199,N_43908);
nand U44894 (N_44894,N_43952,N_42685);
xor U44895 (N_44895,N_42394,N_42294);
and U44896 (N_44896,N_42694,N_43809);
or U44897 (N_44897,N_43407,N_42028);
nand U44898 (N_44898,N_42364,N_42537);
and U44899 (N_44899,N_42067,N_42662);
and U44900 (N_44900,N_43009,N_42130);
or U44901 (N_44901,N_42209,N_42086);
or U44902 (N_44902,N_42401,N_42309);
xnor U44903 (N_44903,N_43393,N_43463);
or U44904 (N_44904,N_42221,N_42002);
or U44905 (N_44905,N_42733,N_43722);
and U44906 (N_44906,N_42133,N_43247);
xnor U44907 (N_44907,N_43251,N_42054);
nor U44908 (N_44908,N_42061,N_42840);
or U44909 (N_44909,N_42532,N_42708);
or U44910 (N_44910,N_43372,N_42968);
and U44911 (N_44911,N_42721,N_43227);
or U44912 (N_44912,N_42400,N_42259);
nor U44913 (N_44913,N_43690,N_42389);
and U44914 (N_44914,N_43643,N_42077);
nand U44915 (N_44915,N_43324,N_43769);
xnor U44916 (N_44916,N_42268,N_43029);
nand U44917 (N_44917,N_42930,N_42429);
and U44918 (N_44918,N_42737,N_43533);
and U44919 (N_44919,N_42488,N_43789);
xnor U44920 (N_44920,N_42433,N_43814);
and U44921 (N_44921,N_42802,N_43948);
nand U44922 (N_44922,N_43934,N_43884);
nand U44923 (N_44923,N_43060,N_43663);
nor U44924 (N_44924,N_42876,N_43700);
nand U44925 (N_44925,N_42796,N_43434);
nor U44926 (N_44926,N_42384,N_42172);
nand U44927 (N_44927,N_43105,N_43507);
and U44928 (N_44928,N_43800,N_42407);
and U44929 (N_44929,N_42874,N_43106);
xor U44930 (N_44930,N_43310,N_43994);
nor U44931 (N_44931,N_42584,N_42934);
and U44932 (N_44932,N_43087,N_43638);
and U44933 (N_44933,N_43444,N_43437);
and U44934 (N_44934,N_42123,N_43381);
or U44935 (N_44935,N_42497,N_43707);
xor U44936 (N_44936,N_42748,N_42517);
xnor U44937 (N_44937,N_43869,N_42381);
nand U44938 (N_44938,N_43603,N_43038);
xor U44939 (N_44939,N_43240,N_43763);
nor U44940 (N_44940,N_43964,N_43041);
nor U44941 (N_44941,N_43525,N_43791);
nor U44942 (N_44942,N_43467,N_43702);
nor U44943 (N_44943,N_42677,N_42691);
or U44944 (N_44944,N_43711,N_43589);
xor U44945 (N_44945,N_43277,N_42539);
xor U44946 (N_44946,N_43371,N_42480);
nor U44947 (N_44947,N_43692,N_43424);
nand U44948 (N_44948,N_43000,N_42343);
or U44949 (N_44949,N_42728,N_42099);
and U44950 (N_44950,N_43344,N_42881);
nor U44951 (N_44951,N_43790,N_42053);
nor U44952 (N_44952,N_43887,N_43059);
xnor U44953 (N_44953,N_42587,N_43254);
and U44954 (N_44954,N_42625,N_42549);
or U44955 (N_44955,N_43955,N_42483);
or U44956 (N_44956,N_42441,N_43959);
xnor U44957 (N_44957,N_43342,N_43969);
and U44958 (N_44958,N_43228,N_42583);
nand U44959 (N_44959,N_43458,N_42659);
or U44960 (N_44960,N_42684,N_43370);
nor U44961 (N_44961,N_42496,N_42450);
nor U44962 (N_44962,N_43975,N_42393);
and U44963 (N_44963,N_42437,N_42380);
xor U44964 (N_44964,N_43055,N_43420);
or U44965 (N_44965,N_43091,N_42936);
nand U44966 (N_44966,N_42000,N_42510);
and U44967 (N_44967,N_42069,N_43348);
and U44968 (N_44968,N_43670,N_43296);
nor U44969 (N_44969,N_43856,N_42418);
xnor U44970 (N_44970,N_43224,N_42189);
xnor U44971 (N_44971,N_42974,N_42415);
or U44972 (N_44972,N_43016,N_42618);
xor U44973 (N_44973,N_42348,N_42669);
and U44974 (N_44974,N_42151,N_42663);
and U44975 (N_44975,N_42838,N_43599);
or U44976 (N_44976,N_43883,N_43366);
nor U44977 (N_44977,N_42346,N_42302);
xnor U44978 (N_44978,N_43166,N_42509);
nor U44979 (N_44979,N_43832,N_43755);
xor U44980 (N_44980,N_43025,N_42186);
nand U44981 (N_44981,N_42449,N_43474);
and U44982 (N_44982,N_42188,N_43838);
or U44983 (N_44983,N_43063,N_42164);
nor U44984 (N_44984,N_43765,N_42135);
or U44985 (N_44985,N_43380,N_42558);
xor U44986 (N_44986,N_42503,N_43468);
xnor U44987 (N_44987,N_42782,N_43947);
nor U44988 (N_44988,N_43023,N_43880);
nor U44989 (N_44989,N_42500,N_43287);
or U44990 (N_44990,N_42650,N_43965);
or U44991 (N_44991,N_42317,N_43506);
or U44992 (N_44992,N_42058,N_43796);
or U44993 (N_44993,N_42270,N_42753);
nor U44994 (N_44994,N_43076,N_42614);
xor U44995 (N_44995,N_42996,N_42706);
or U44996 (N_44996,N_42296,N_43606);
nand U44997 (N_44997,N_42715,N_43503);
nor U44998 (N_44998,N_42154,N_42919);
xnor U44999 (N_44999,N_43915,N_43633);
and U45000 (N_45000,N_42393,N_42961);
or U45001 (N_45001,N_42169,N_43534);
or U45002 (N_45002,N_43544,N_43775);
nand U45003 (N_45003,N_42255,N_43617);
xnor U45004 (N_45004,N_43288,N_43268);
or U45005 (N_45005,N_43753,N_43822);
xnor U45006 (N_45006,N_43469,N_42807);
and U45007 (N_45007,N_42628,N_42989);
nand U45008 (N_45008,N_43854,N_42563);
nand U45009 (N_45009,N_43627,N_43987);
xor U45010 (N_45010,N_43471,N_43068);
nor U45011 (N_45011,N_42729,N_42080);
and U45012 (N_45012,N_43873,N_43530);
and U45013 (N_45013,N_43038,N_43383);
nand U45014 (N_45014,N_42226,N_42446);
nor U45015 (N_45015,N_43351,N_43238);
or U45016 (N_45016,N_43111,N_43507);
nor U45017 (N_45017,N_43493,N_43627);
xnor U45018 (N_45018,N_43122,N_43237);
xnor U45019 (N_45019,N_43180,N_43421);
xnor U45020 (N_45020,N_42299,N_42133);
nor U45021 (N_45021,N_43436,N_42440);
or U45022 (N_45022,N_42988,N_42742);
nor U45023 (N_45023,N_43741,N_42187);
xnor U45024 (N_45024,N_42689,N_43171);
nand U45025 (N_45025,N_43223,N_43876);
xor U45026 (N_45026,N_43514,N_43688);
xnor U45027 (N_45027,N_43007,N_42621);
and U45028 (N_45028,N_42415,N_43319);
or U45029 (N_45029,N_42374,N_43350);
xor U45030 (N_45030,N_43164,N_42314);
and U45031 (N_45031,N_42235,N_42176);
nor U45032 (N_45032,N_42119,N_43959);
or U45033 (N_45033,N_42152,N_43737);
xor U45034 (N_45034,N_42708,N_43428);
nand U45035 (N_45035,N_42756,N_43305);
xnor U45036 (N_45036,N_43440,N_42365);
nand U45037 (N_45037,N_43888,N_42921);
nand U45038 (N_45038,N_43492,N_42004);
nand U45039 (N_45039,N_43238,N_43205);
nand U45040 (N_45040,N_43177,N_42158);
xnor U45041 (N_45041,N_43100,N_43664);
and U45042 (N_45042,N_42467,N_43491);
or U45043 (N_45043,N_42295,N_42208);
xnor U45044 (N_45044,N_43107,N_43124);
nor U45045 (N_45045,N_42715,N_42502);
nand U45046 (N_45046,N_42829,N_42256);
and U45047 (N_45047,N_42535,N_42335);
or U45048 (N_45048,N_42018,N_43315);
and U45049 (N_45049,N_42054,N_43046);
nor U45050 (N_45050,N_42016,N_43735);
nand U45051 (N_45051,N_42046,N_43846);
or U45052 (N_45052,N_43150,N_42355);
nor U45053 (N_45053,N_42364,N_42800);
xnor U45054 (N_45054,N_43563,N_43109);
and U45055 (N_45055,N_43231,N_42251);
nand U45056 (N_45056,N_42438,N_42011);
or U45057 (N_45057,N_42871,N_43843);
or U45058 (N_45058,N_43923,N_42368);
or U45059 (N_45059,N_43390,N_43053);
nor U45060 (N_45060,N_42394,N_42984);
nor U45061 (N_45061,N_43859,N_43355);
or U45062 (N_45062,N_42849,N_43577);
or U45063 (N_45063,N_43653,N_43212);
nand U45064 (N_45064,N_43611,N_43543);
nor U45065 (N_45065,N_43709,N_43294);
xor U45066 (N_45066,N_43239,N_42501);
nand U45067 (N_45067,N_43896,N_43704);
and U45068 (N_45068,N_43939,N_42141);
nand U45069 (N_45069,N_43680,N_43803);
and U45070 (N_45070,N_42631,N_42627);
nand U45071 (N_45071,N_43823,N_42782);
nand U45072 (N_45072,N_43318,N_43730);
and U45073 (N_45073,N_43742,N_42128);
and U45074 (N_45074,N_43147,N_43493);
or U45075 (N_45075,N_43338,N_42641);
and U45076 (N_45076,N_42868,N_42175);
nand U45077 (N_45077,N_43950,N_42598);
nand U45078 (N_45078,N_42264,N_43757);
xnor U45079 (N_45079,N_42195,N_42563);
and U45080 (N_45080,N_43108,N_42570);
and U45081 (N_45081,N_42461,N_43125);
or U45082 (N_45082,N_42724,N_43927);
and U45083 (N_45083,N_43017,N_42829);
or U45084 (N_45084,N_43737,N_42595);
xnor U45085 (N_45085,N_42007,N_43839);
xor U45086 (N_45086,N_42155,N_42436);
and U45087 (N_45087,N_42329,N_42163);
nand U45088 (N_45088,N_43138,N_43315);
nor U45089 (N_45089,N_42067,N_42357);
and U45090 (N_45090,N_42626,N_43050);
and U45091 (N_45091,N_42046,N_42463);
and U45092 (N_45092,N_42365,N_42139);
and U45093 (N_45093,N_43781,N_43401);
and U45094 (N_45094,N_43783,N_43378);
and U45095 (N_45095,N_42727,N_42841);
nor U45096 (N_45096,N_43826,N_43958);
and U45097 (N_45097,N_43156,N_43580);
nor U45098 (N_45098,N_43768,N_42107);
nand U45099 (N_45099,N_42532,N_43820);
xor U45100 (N_45100,N_43791,N_43182);
xnor U45101 (N_45101,N_42361,N_42112);
nor U45102 (N_45102,N_42374,N_43389);
xor U45103 (N_45103,N_42300,N_42980);
and U45104 (N_45104,N_42719,N_43522);
or U45105 (N_45105,N_43357,N_43304);
nand U45106 (N_45106,N_43359,N_43966);
nor U45107 (N_45107,N_43484,N_42836);
or U45108 (N_45108,N_42494,N_43453);
and U45109 (N_45109,N_42079,N_42319);
xnor U45110 (N_45110,N_42878,N_43715);
nor U45111 (N_45111,N_43544,N_43434);
and U45112 (N_45112,N_43762,N_42421);
or U45113 (N_45113,N_42961,N_43190);
xnor U45114 (N_45114,N_42926,N_43296);
and U45115 (N_45115,N_43124,N_43783);
or U45116 (N_45116,N_42695,N_43906);
nand U45117 (N_45117,N_43799,N_42499);
or U45118 (N_45118,N_42124,N_42018);
and U45119 (N_45119,N_43906,N_42567);
or U45120 (N_45120,N_42373,N_43252);
and U45121 (N_45121,N_43837,N_42514);
nand U45122 (N_45122,N_42537,N_43726);
xnor U45123 (N_45123,N_42285,N_42601);
nor U45124 (N_45124,N_42279,N_42143);
xnor U45125 (N_45125,N_43675,N_42097);
or U45126 (N_45126,N_43162,N_42418);
and U45127 (N_45127,N_43103,N_42809);
or U45128 (N_45128,N_43769,N_43169);
and U45129 (N_45129,N_42646,N_42462);
nand U45130 (N_45130,N_42977,N_42607);
nand U45131 (N_45131,N_42629,N_42045);
nand U45132 (N_45132,N_43965,N_43001);
nand U45133 (N_45133,N_43873,N_43779);
or U45134 (N_45134,N_42372,N_43913);
nand U45135 (N_45135,N_42622,N_43579);
and U45136 (N_45136,N_43542,N_43750);
xor U45137 (N_45137,N_43738,N_42060);
or U45138 (N_45138,N_43225,N_42218);
nand U45139 (N_45139,N_43669,N_43218);
and U45140 (N_45140,N_43061,N_43130);
nor U45141 (N_45141,N_42815,N_42167);
or U45142 (N_45142,N_43121,N_42249);
nand U45143 (N_45143,N_43159,N_43236);
or U45144 (N_45144,N_42968,N_43226);
and U45145 (N_45145,N_42114,N_43572);
and U45146 (N_45146,N_42993,N_42283);
nand U45147 (N_45147,N_43977,N_42444);
nor U45148 (N_45148,N_42336,N_43907);
nor U45149 (N_45149,N_43069,N_43484);
or U45150 (N_45150,N_43265,N_42163);
xor U45151 (N_45151,N_42510,N_43887);
or U45152 (N_45152,N_42389,N_42390);
nor U45153 (N_45153,N_42333,N_42390);
nor U45154 (N_45154,N_43754,N_43452);
nand U45155 (N_45155,N_42723,N_43634);
and U45156 (N_45156,N_43492,N_43436);
or U45157 (N_45157,N_42713,N_42385);
nand U45158 (N_45158,N_42600,N_42228);
nand U45159 (N_45159,N_42331,N_43174);
nor U45160 (N_45160,N_43958,N_42318);
and U45161 (N_45161,N_42556,N_43645);
and U45162 (N_45162,N_42610,N_43764);
xor U45163 (N_45163,N_43844,N_43697);
and U45164 (N_45164,N_43521,N_42215);
xnor U45165 (N_45165,N_42543,N_43943);
nor U45166 (N_45166,N_42842,N_43317);
nor U45167 (N_45167,N_42483,N_43805);
nand U45168 (N_45168,N_43901,N_42900);
and U45169 (N_45169,N_42610,N_42005);
nand U45170 (N_45170,N_42915,N_42645);
and U45171 (N_45171,N_43924,N_42323);
or U45172 (N_45172,N_42290,N_43868);
nor U45173 (N_45173,N_43580,N_42984);
xor U45174 (N_45174,N_42759,N_42346);
xor U45175 (N_45175,N_43512,N_43039);
xor U45176 (N_45176,N_43454,N_43564);
xnor U45177 (N_45177,N_43906,N_42705);
or U45178 (N_45178,N_43451,N_43991);
or U45179 (N_45179,N_43750,N_42580);
nor U45180 (N_45180,N_42066,N_42301);
or U45181 (N_45181,N_43622,N_42635);
nor U45182 (N_45182,N_43126,N_43263);
nor U45183 (N_45183,N_42687,N_43329);
nand U45184 (N_45184,N_42941,N_42212);
and U45185 (N_45185,N_43564,N_42690);
nor U45186 (N_45186,N_42443,N_43242);
xor U45187 (N_45187,N_42890,N_43898);
nor U45188 (N_45188,N_43136,N_43402);
nand U45189 (N_45189,N_42263,N_42009);
and U45190 (N_45190,N_42850,N_42006);
nor U45191 (N_45191,N_42509,N_42004);
and U45192 (N_45192,N_42063,N_43508);
nand U45193 (N_45193,N_42760,N_42603);
or U45194 (N_45194,N_43475,N_43622);
nor U45195 (N_45195,N_43888,N_43506);
or U45196 (N_45196,N_43556,N_43786);
xnor U45197 (N_45197,N_43181,N_43208);
nor U45198 (N_45198,N_42157,N_43572);
or U45199 (N_45199,N_42089,N_43781);
nand U45200 (N_45200,N_42192,N_43381);
or U45201 (N_45201,N_43661,N_43453);
nor U45202 (N_45202,N_42690,N_43823);
nor U45203 (N_45203,N_42901,N_42563);
or U45204 (N_45204,N_43184,N_42109);
xnor U45205 (N_45205,N_42608,N_43583);
and U45206 (N_45206,N_42569,N_42131);
nor U45207 (N_45207,N_42651,N_43169);
and U45208 (N_45208,N_42412,N_43957);
or U45209 (N_45209,N_43959,N_42292);
nand U45210 (N_45210,N_42135,N_43501);
or U45211 (N_45211,N_43635,N_43032);
nor U45212 (N_45212,N_42129,N_43329);
or U45213 (N_45213,N_43481,N_42050);
nand U45214 (N_45214,N_43655,N_43931);
nor U45215 (N_45215,N_42274,N_42700);
or U45216 (N_45216,N_43203,N_43835);
nand U45217 (N_45217,N_43546,N_42676);
nor U45218 (N_45218,N_43495,N_43067);
nand U45219 (N_45219,N_42693,N_42397);
nand U45220 (N_45220,N_42543,N_43879);
nor U45221 (N_45221,N_42642,N_42912);
xor U45222 (N_45222,N_43891,N_43323);
or U45223 (N_45223,N_42831,N_43484);
and U45224 (N_45224,N_43715,N_42513);
xor U45225 (N_45225,N_42076,N_43477);
xor U45226 (N_45226,N_43972,N_42826);
and U45227 (N_45227,N_43338,N_43420);
xnor U45228 (N_45228,N_43101,N_42299);
nor U45229 (N_45229,N_43859,N_43117);
xor U45230 (N_45230,N_42864,N_42238);
or U45231 (N_45231,N_43343,N_43436);
nand U45232 (N_45232,N_43554,N_43990);
nor U45233 (N_45233,N_43199,N_43471);
nand U45234 (N_45234,N_42446,N_43451);
nand U45235 (N_45235,N_42616,N_42046);
xnor U45236 (N_45236,N_42187,N_43127);
nor U45237 (N_45237,N_43088,N_43743);
xor U45238 (N_45238,N_42781,N_43084);
nand U45239 (N_45239,N_43586,N_42488);
nor U45240 (N_45240,N_43155,N_43511);
nor U45241 (N_45241,N_43438,N_42922);
xor U45242 (N_45242,N_43628,N_43366);
nor U45243 (N_45243,N_43198,N_43135);
and U45244 (N_45244,N_42296,N_42513);
xor U45245 (N_45245,N_42480,N_42926);
or U45246 (N_45246,N_43011,N_43951);
nor U45247 (N_45247,N_43359,N_43676);
xor U45248 (N_45248,N_43361,N_42169);
xnor U45249 (N_45249,N_42118,N_42136);
or U45250 (N_45250,N_42461,N_43437);
or U45251 (N_45251,N_43458,N_42877);
nand U45252 (N_45252,N_42404,N_43738);
and U45253 (N_45253,N_42865,N_42582);
and U45254 (N_45254,N_42277,N_43790);
xnor U45255 (N_45255,N_42852,N_42224);
nand U45256 (N_45256,N_43993,N_42170);
nor U45257 (N_45257,N_42552,N_43847);
nor U45258 (N_45258,N_43757,N_42316);
and U45259 (N_45259,N_43496,N_42379);
or U45260 (N_45260,N_42166,N_43381);
nor U45261 (N_45261,N_43378,N_42137);
nand U45262 (N_45262,N_43986,N_42725);
nand U45263 (N_45263,N_43803,N_42159);
xnor U45264 (N_45264,N_43278,N_43793);
or U45265 (N_45265,N_43973,N_42136);
and U45266 (N_45266,N_42206,N_42434);
and U45267 (N_45267,N_43286,N_42038);
and U45268 (N_45268,N_42155,N_43534);
or U45269 (N_45269,N_42177,N_43091);
and U45270 (N_45270,N_43958,N_42237);
xnor U45271 (N_45271,N_42998,N_42865);
xnor U45272 (N_45272,N_42249,N_43229);
and U45273 (N_45273,N_42439,N_42915);
and U45274 (N_45274,N_43050,N_42678);
nand U45275 (N_45275,N_42186,N_43685);
nand U45276 (N_45276,N_43062,N_43121);
or U45277 (N_45277,N_43821,N_43621);
nand U45278 (N_45278,N_43845,N_42017);
or U45279 (N_45279,N_42628,N_42082);
nor U45280 (N_45280,N_42580,N_43016);
and U45281 (N_45281,N_43513,N_43271);
nor U45282 (N_45282,N_43876,N_43772);
nand U45283 (N_45283,N_42218,N_43535);
and U45284 (N_45284,N_43877,N_42764);
nor U45285 (N_45285,N_42471,N_43394);
and U45286 (N_45286,N_42545,N_43332);
and U45287 (N_45287,N_43390,N_42903);
nor U45288 (N_45288,N_42766,N_42227);
nand U45289 (N_45289,N_43963,N_43000);
or U45290 (N_45290,N_43490,N_42531);
xor U45291 (N_45291,N_42298,N_43491);
nand U45292 (N_45292,N_43807,N_43327);
and U45293 (N_45293,N_43669,N_42493);
nor U45294 (N_45294,N_42837,N_42385);
nand U45295 (N_45295,N_43349,N_43207);
nor U45296 (N_45296,N_43320,N_43595);
nor U45297 (N_45297,N_42823,N_42501);
xor U45298 (N_45298,N_43172,N_43212);
nand U45299 (N_45299,N_43817,N_43469);
or U45300 (N_45300,N_42224,N_43392);
nand U45301 (N_45301,N_42308,N_43045);
and U45302 (N_45302,N_42003,N_42582);
nor U45303 (N_45303,N_43945,N_42895);
xnor U45304 (N_45304,N_42052,N_43927);
xor U45305 (N_45305,N_42275,N_42421);
and U45306 (N_45306,N_42071,N_43538);
and U45307 (N_45307,N_42084,N_43175);
or U45308 (N_45308,N_43935,N_42993);
nor U45309 (N_45309,N_42442,N_43707);
nand U45310 (N_45310,N_43242,N_42742);
nor U45311 (N_45311,N_42245,N_42810);
or U45312 (N_45312,N_43308,N_42109);
and U45313 (N_45313,N_43341,N_42585);
nand U45314 (N_45314,N_42961,N_42735);
nor U45315 (N_45315,N_43407,N_42324);
nand U45316 (N_45316,N_42547,N_42919);
or U45317 (N_45317,N_43200,N_42787);
nor U45318 (N_45318,N_42037,N_43412);
nand U45319 (N_45319,N_42930,N_42944);
xor U45320 (N_45320,N_42326,N_43224);
nor U45321 (N_45321,N_43062,N_43225);
nand U45322 (N_45322,N_42745,N_43306);
xnor U45323 (N_45323,N_42992,N_42348);
nor U45324 (N_45324,N_42149,N_42607);
nand U45325 (N_45325,N_42796,N_42963);
nand U45326 (N_45326,N_42093,N_43634);
xnor U45327 (N_45327,N_43229,N_42874);
nand U45328 (N_45328,N_43831,N_42432);
xnor U45329 (N_45329,N_43811,N_42962);
and U45330 (N_45330,N_43538,N_43608);
nand U45331 (N_45331,N_42465,N_42102);
or U45332 (N_45332,N_43731,N_42999);
xnor U45333 (N_45333,N_43138,N_43319);
xor U45334 (N_45334,N_42178,N_43722);
xnor U45335 (N_45335,N_42761,N_43398);
nand U45336 (N_45336,N_42275,N_43118);
and U45337 (N_45337,N_42156,N_42221);
xnor U45338 (N_45338,N_42789,N_42481);
nand U45339 (N_45339,N_42838,N_42025);
nor U45340 (N_45340,N_43807,N_42333);
xor U45341 (N_45341,N_42763,N_43738);
nor U45342 (N_45342,N_42087,N_42999);
xnor U45343 (N_45343,N_42546,N_42001);
or U45344 (N_45344,N_42260,N_42983);
nand U45345 (N_45345,N_42761,N_43553);
and U45346 (N_45346,N_43094,N_42153);
and U45347 (N_45347,N_43467,N_42834);
xor U45348 (N_45348,N_42762,N_43375);
and U45349 (N_45349,N_42348,N_43359);
nand U45350 (N_45350,N_42046,N_43670);
and U45351 (N_45351,N_43040,N_43257);
nor U45352 (N_45352,N_43122,N_43832);
nand U45353 (N_45353,N_42401,N_42642);
xor U45354 (N_45354,N_43082,N_43256);
nand U45355 (N_45355,N_43663,N_42152);
and U45356 (N_45356,N_43328,N_43191);
or U45357 (N_45357,N_42813,N_42026);
nand U45358 (N_45358,N_42099,N_42928);
nor U45359 (N_45359,N_43428,N_43936);
nor U45360 (N_45360,N_42830,N_43196);
or U45361 (N_45361,N_42143,N_42947);
or U45362 (N_45362,N_43673,N_43414);
and U45363 (N_45363,N_42009,N_42674);
nor U45364 (N_45364,N_42771,N_42539);
and U45365 (N_45365,N_42420,N_43122);
and U45366 (N_45366,N_43162,N_43386);
or U45367 (N_45367,N_42680,N_42806);
or U45368 (N_45368,N_43065,N_42825);
and U45369 (N_45369,N_42264,N_43354);
nand U45370 (N_45370,N_42248,N_43928);
and U45371 (N_45371,N_43913,N_43338);
and U45372 (N_45372,N_42391,N_42188);
nor U45373 (N_45373,N_43180,N_42268);
nor U45374 (N_45374,N_43233,N_43039);
and U45375 (N_45375,N_42049,N_42202);
or U45376 (N_45376,N_43221,N_42383);
nand U45377 (N_45377,N_43093,N_43913);
or U45378 (N_45378,N_42007,N_42152);
nand U45379 (N_45379,N_42836,N_42277);
xor U45380 (N_45380,N_42459,N_43326);
xnor U45381 (N_45381,N_43478,N_42092);
and U45382 (N_45382,N_42889,N_43098);
or U45383 (N_45383,N_42113,N_42210);
or U45384 (N_45384,N_42999,N_43754);
or U45385 (N_45385,N_42767,N_43541);
nand U45386 (N_45386,N_42666,N_42669);
nand U45387 (N_45387,N_42698,N_42275);
and U45388 (N_45388,N_43100,N_43091);
nor U45389 (N_45389,N_43912,N_43227);
and U45390 (N_45390,N_43344,N_42495);
and U45391 (N_45391,N_42657,N_42739);
xnor U45392 (N_45392,N_43345,N_43058);
nor U45393 (N_45393,N_42376,N_42186);
nor U45394 (N_45394,N_42423,N_43354);
or U45395 (N_45395,N_42058,N_42356);
xor U45396 (N_45396,N_43968,N_43171);
nand U45397 (N_45397,N_42429,N_43745);
xor U45398 (N_45398,N_42744,N_42644);
nand U45399 (N_45399,N_43643,N_42825);
xor U45400 (N_45400,N_43184,N_42300);
or U45401 (N_45401,N_43518,N_42944);
and U45402 (N_45402,N_43776,N_42531);
nor U45403 (N_45403,N_42674,N_42851);
nand U45404 (N_45404,N_43066,N_42446);
nor U45405 (N_45405,N_42357,N_42470);
and U45406 (N_45406,N_42237,N_42545);
nor U45407 (N_45407,N_43525,N_43472);
nor U45408 (N_45408,N_43116,N_43420);
or U45409 (N_45409,N_42932,N_43354);
and U45410 (N_45410,N_42367,N_42407);
xnor U45411 (N_45411,N_43103,N_42168);
or U45412 (N_45412,N_42418,N_42731);
xor U45413 (N_45413,N_43313,N_43759);
and U45414 (N_45414,N_43688,N_42523);
nor U45415 (N_45415,N_42132,N_43010);
and U45416 (N_45416,N_42999,N_42235);
nand U45417 (N_45417,N_43818,N_43815);
or U45418 (N_45418,N_43371,N_43100);
and U45419 (N_45419,N_42614,N_42860);
and U45420 (N_45420,N_42619,N_43031);
or U45421 (N_45421,N_43215,N_42768);
or U45422 (N_45422,N_43207,N_42999);
or U45423 (N_45423,N_43802,N_43118);
or U45424 (N_45424,N_43474,N_42502);
or U45425 (N_45425,N_42891,N_43926);
nor U45426 (N_45426,N_43802,N_42442);
nor U45427 (N_45427,N_43110,N_42721);
nor U45428 (N_45428,N_43195,N_42173);
nor U45429 (N_45429,N_42178,N_43751);
xnor U45430 (N_45430,N_43255,N_42361);
and U45431 (N_45431,N_42868,N_43682);
xnor U45432 (N_45432,N_42611,N_42725);
and U45433 (N_45433,N_43312,N_43663);
nor U45434 (N_45434,N_43697,N_42106);
and U45435 (N_45435,N_43301,N_43395);
or U45436 (N_45436,N_42672,N_43162);
nor U45437 (N_45437,N_43638,N_42770);
xor U45438 (N_45438,N_42974,N_42989);
and U45439 (N_45439,N_43247,N_43920);
nor U45440 (N_45440,N_43901,N_42091);
and U45441 (N_45441,N_42195,N_42001);
and U45442 (N_45442,N_43431,N_42283);
xor U45443 (N_45443,N_42649,N_42872);
or U45444 (N_45444,N_43694,N_43959);
xor U45445 (N_45445,N_43835,N_42507);
or U45446 (N_45446,N_42901,N_42106);
nand U45447 (N_45447,N_43959,N_43875);
nand U45448 (N_45448,N_42141,N_43830);
or U45449 (N_45449,N_42838,N_42020);
nand U45450 (N_45450,N_42648,N_43610);
nor U45451 (N_45451,N_43034,N_43837);
nand U45452 (N_45452,N_42657,N_42815);
nor U45453 (N_45453,N_43874,N_43663);
nand U45454 (N_45454,N_43803,N_42998);
nor U45455 (N_45455,N_43662,N_42158);
nand U45456 (N_45456,N_42250,N_42711);
nand U45457 (N_45457,N_42702,N_42095);
and U45458 (N_45458,N_42317,N_43759);
nand U45459 (N_45459,N_42174,N_43182);
xnor U45460 (N_45460,N_42795,N_42701);
and U45461 (N_45461,N_43691,N_42975);
and U45462 (N_45462,N_42831,N_43965);
or U45463 (N_45463,N_42850,N_43671);
nand U45464 (N_45464,N_43366,N_42704);
and U45465 (N_45465,N_43675,N_43510);
nor U45466 (N_45466,N_42901,N_42766);
and U45467 (N_45467,N_43205,N_43882);
xor U45468 (N_45468,N_43119,N_43022);
or U45469 (N_45469,N_43517,N_43232);
xnor U45470 (N_45470,N_42929,N_43602);
nor U45471 (N_45471,N_43682,N_43247);
and U45472 (N_45472,N_43855,N_42377);
xor U45473 (N_45473,N_42024,N_43979);
or U45474 (N_45474,N_42948,N_42566);
and U45475 (N_45475,N_43727,N_42657);
and U45476 (N_45476,N_43128,N_42145);
or U45477 (N_45477,N_43931,N_43865);
nor U45478 (N_45478,N_43833,N_42297);
nor U45479 (N_45479,N_42960,N_43231);
nand U45480 (N_45480,N_43442,N_42028);
xor U45481 (N_45481,N_42324,N_43047);
nor U45482 (N_45482,N_43096,N_43418);
nor U45483 (N_45483,N_42996,N_43231);
or U45484 (N_45484,N_43531,N_43271);
and U45485 (N_45485,N_43862,N_42491);
and U45486 (N_45486,N_43440,N_42944);
nand U45487 (N_45487,N_43405,N_42526);
nand U45488 (N_45488,N_42442,N_43189);
nand U45489 (N_45489,N_43698,N_42182);
nand U45490 (N_45490,N_43598,N_42036);
nand U45491 (N_45491,N_42296,N_42102);
nor U45492 (N_45492,N_42927,N_43626);
nand U45493 (N_45493,N_43383,N_43106);
xor U45494 (N_45494,N_42076,N_42894);
nand U45495 (N_45495,N_42979,N_43942);
and U45496 (N_45496,N_42337,N_42999);
nand U45497 (N_45497,N_43316,N_42416);
xnor U45498 (N_45498,N_42333,N_43075);
and U45499 (N_45499,N_43079,N_42542);
and U45500 (N_45500,N_43101,N_42283);
or U45501 (N_45501,N_43055,N_43894);
xor U45502 (N_45502,N_42853,N_42336);
nand U45503 (N_45503,N_43320,N_43767);
nand U45504 (N_45504,N_43007,N_42987);
nor U45505 (N_45505,N_42544,N_43574);
nor U45506 (N_45506,N_42152,N_43861);
nor U45507 (N_45507,N_42400,N_42432);
or U45508 (N_45508,N_42034,N_42350);
nor U45509 (N_45509,N_43836,N_43143);
and U45510 (N_45510,N_42866,N_43240);
or U45511 (N_45511,N_43402,N_43763);
xor U45512 (N_45512,N_43721,N_42151);
nand U45513 (N_45513,N_42746,N_42369);
xnor U45514 (N_45514,N_43778,N_43265);
nor U45515 (N_45515,N_43614,N_43818);
nand U45516 (N_45516,N_43465,N_43431);
nor U45517 (N_45517,N_43287,N_42572);
and U45518 (N_45518,N_43030,N_42389);
xor U45519 (N_45519,N_43096,N_42297);
xnor U45520 (N_45520,N_42719,N_43563);
and U45521 (N_45521,N_43877,N_42955);
or U45522 (N_45522,N_42661,N_43878);
nor U45523 (N_45523,N_42361,N_42256);
nor U45524 (N_45524,N_43096,N_43646);
nand U45525 (N_45525,N_43161,N_42667);
and U45526 (N_45526,N_42822,N_43004);
nand U45527 (N_45527,N_42318,N_42550);
nor U45528 (N_45528,N_43977,N_42464);
or U45529 (N_45529,N_43122,N_42438);
or U45530 (N_45530,N_42351,N_42082);
or U45531 (N_45531,N_42945,N_43052);
nor U45532 (N_45532,N_43590,N_43408);
nor U45533 (N_45533,N_43404,N_43770);
nor U45534 (N_45534,N_42266,N_42554);
nor U45535 (N_45535,N_43388,N_43455);
nand U45536 (N_45536,N_43335,N_42024);
xnor U45537 (N_45537,N_43212,N_42986);
nor U45538 (N_45538,N_42629,N_43113);
nand U45539 (N_45539,N_43264,N_43828);
nand U45540 (N_45540,N_42048,N_42769);
xnor U45541 (N_45541,N_43523,N_42733);
nor U45542 (N_45542,N_42994,N_43354);
and U45543 (N_45543,N_42423,N_42684);
nor U45544 (N_45544,N_42359,N_42518);
xor U45545 (N_45545,N_43643,N_43210);
nor U45546 (N_45546,N_43567,N_43329);
xor U45547 (N_45547,N_42190,N_43873);
nor U45548 (N_45548,N_42613,N_43635);
and U45549 (N_45549,N_42590,N_42574);
or U45550 (N_45550,N_43156,N_42920);
or U45551 (N_45551,N_42227,N_42341);
nor U45552 (N_45552,N_42862,N_43344);
nor U45553 (N_45553,N_43307,N_43030);
nor U45554 (N_45554,N_43205,N_42368);
and U45555 (N_45555,N_43466,N_43908);
and U45556 (N_45556,N_43598,N_43858);
nor U45557 (N_45557,N_43251,N_42840);
nor U45558 (N_45558,N_43319,N_42150);
xor U45559 (N_45559,N_43669,N_43424);
or U45560 (N_45560,N_43308,N_42964);
xnor U45561 (N_45561,N_43337,N_43306);
nor U45562 (N_45562,N_43779,N_42827);
or U45563 (N_45563,N_43172,N_42136);
nand U45564 (N_45564,N_43712,N_43301);
nand U45565 (N_45565,N_43306,N_42036);
or U45566 (N_45566,N_43466,N_42428);
and U45567 (N_45567,N_42602,N_42581);
xor U45568 (N_45568,N_43036,N_42465);
or U45569 (N_45569,N_42261,N_43744);
xor U45570 (N_45570,N_42306,N_42687);
nor U45571 (N_45571,N_42742,N_42620);
nand U45572 (N_45572,N_43948,N_43466);
nand U45573 (N_45573,N_42251,N_43979);
xor U45574 (N_45574,N_43534,N_42370);
or U45575 (N_45575,N_42340,N_43791);
nor U45576 (N_45576,N_43287,N_43004);
nor U45577 (N_45577,N_43929,N_43463);
nor U45578 (N_45578,N_42492,N_42733);
or U45579 (N_45579,N_43886,N_43705);
nand U45580 (N_45580,N_43541,N_43356);
xor U45581 (N_45581,N_42506,N_42032);
nand U45582 (N_45582,N_43359,N_43824);
and U45583 (N_45583,N_42061,N_42960);
xor U45584 (N_45584,N_42382,N_43425);
nand U45585 (N_45585,N_43479,N_43629);
and U45586 (N_45586,N_42779,N_42195);
or U45587 (N_45587,N_43064,N_43855);
and U45588 (N_45588,N_43115,N_43079);
or U45589 (N_45589,N_43860,N_42074);
nor U45590 (N_45590,N_43707,N_43616);
xnor U45591 (N_45591,N_43893,N_42143);
and U45592 (N_45592,N_42876,N_43888);
and U45593 (N_45593,N_43288,N_43897);
xor U45594 (N_45594,N_43861,N_42012);
nor U45595 (N_45595,N_42900,N_42614);
nand U45596 (N_45596,N_42720,N_43983);
nor U45597 (N_45597,N_43061,N_42355);
xnor U45598 (N_45598,N_42348,N_43639);
nand U45599 (N_45599,N_42510,N_42641);
nand U45600 (N_45600,N_42300,N_43471);
nand U45601 (N_45601,N_43882,N_43260);
nand U45602 (N_45602,N_42831,N_42137);
nand U45603 (N_45603,N_43443,N_43352);
nor U45604 (N_45604,N_42483,N_42492);
and U45605 (N_45605,N_42418,N_43672);
nor U45606 (N_45606,N_43262,N_43071);
nor U45607 (N_45607,N_42938,N_43717);
nor U45608 (N_45608,N_42589,N_42035);
nand U45609 (N_45609,N_42304,N_42978);
or U45610 (N_45610,N_42323,N_42266);
and U45611 (N_45611,N_42260,N_42653);
nand U45612 (N_45612,N_43139,N_43243);
nand U45613 (N_45613,N_43378,N_43497);
or U45614 (N_45614,N_43750,N_42131);
and U45615 (N_45615,N_42920,N_42578);
or U45616 (N_45616,N_42965,N_42659);
nor U45617 (N_45617,N_42944,N_42183);
and U45618 (N_45618,N_43118,N_43808);
or U45619 (N_45619,N_42873,N_42414);
nor U45620 (N_45620,N_42233,N_43806);
nor U45621 (N_45621,N_43490,N_42728);
xnor U45622 (N_45622,N_42153,N_43995);
xnor U45623 (N_45623,N_43388,N_42895);
or U45624 (N_45624,N_42472,N_42861);
and U45625 (N_45625,N_42002,N_43472);
and U45626 (N_45626,N_42996,N_42663);
or U45627 (N_45627,N_42921,N_42241);
or U45628 (N_45628,N_43005,N_42880);
xor U45629 (N_45629,N_42887,N_43342);
or U45630 (N_45630,N_43791,N_42569);
and U45631 (N_45631,N_42530,N_43208);
nor U45632 (N_45632,N_43541,N_42822);
or U45633 (N_45633,N_43472,N_42569);
xor U45634 (N_45634,N_43556,N_43424);
nor U45635 (N_45635,N_42529,N_43280);
or U45636 (N_45636,N_42729,N_43805);
nand U45637 (N_45637,N_43200,N_42777);
or U45638 (N_45638,N_42664,N_42385);
nor U45639 (N_45639,N_42516,N_42090);
and U45640 (N_45640,N_43935,N_42231);
or U45641 (N_45641,N_43269,N_42650);
xnor U45642 (N_45642,N_43703,N_42419);
xnor U45643 (N_45643,N_43270,N_42806);
or U45644 (N_45644,N_42872,N_43139);
or U45645 (N_45645,N_42551,N_42236);
nand U45646 (N_45646,N_43838,N_42129);
nand U45647 (N_45647,N_43119,N_43990);
xor U45648 (N_45648,N_42533,N_42985);
xnor U45649 (N_45649,N_42481,N_43526);
or U45650 (N_45650,N_43525,N_43424);
nand U45651 (N_45651,N_43640,N_42719);
or U45652 (N_45652,N_43613,N_42030);
or U45653 (N_45653,N_42267,N_42439);
or U45654 (N_45654,N_43808,N_42362);
or U45655 (N_45655,N_42856,N_43353);
nand U45656 (N_45656,N_42235,N_42101);
xnor U45657 (N_45657,N_42294,N_42195);
nor U45658 (N_45658,N_43216,N_43688);
nand U45659 (N_45659,N_42992,N_42107);
xnor U45660 (N_45660,N_43009,N_43707);
or U45661 (N_45661,N_43555,N_42810);
nand U45662 (N_45662,N_43831,N_43105);
nand U45663 (N_45663,N_43958,N_42871);
and U45664 (N_45664,N_42996,N_43114);
nand U45665 (N_45665,N_43833,N_43092);
or U45666 (N_45666,N_42445,N_43988);
and U45667 (N_45667,N_43050,N_43286);
and U45668 (N_45668,N_42729,N_42944);
or U45669 (N_45669,N_42291,N_43728);
nand U45670 (N_45670,N_43239,N_43608);
or U45671 (N_45671,N_43200,N_43783);
or U45672 (N_45672,N_43543,N_43454);
nand U45673 (N_45673,N_42489,N_42987);
nor U45674 (N_45674,N_42986,N_43691);
and U45675 (N_45675,N_43164,N_43589);
and U45676 (N_45676,N_42573,N_42170);
nor U45677 (N_45677,N_42066,N_42722);
nor U45678 (N_45678,N_43004,N_42300);
nor U45679 (N_45679,N_42014,N_42281);
and U45680 (N_45680,N_43945,N_42358);
and U45681 (N_45681,N_43538,N_43146);
xor U45682 (N_45682,N_43940,N_42832);
nor U45683 (N_45683,N_42912,N_43020);
nor U45684 (N_45684,N_42638,N_43561);
or U45685 (N_45685,N_42558,N_42466);
or U45686 (N_45686,N_42889,N_43189);
or U45687 (N_45687,N_42245,N_42603);
xnor U45688 (N_45688,N_42762,N_43438);
xor U45689 (N_45689,N_43451,N_43005);
xor U45690 (N_45690,N_42790,N_43730);
xnor U45691 (N_45691,N_42176,N_43351);
xnor U45692 (N_45692,N_42867,N_43119);
nand U45693 (N_45693,N_43074,N_42468);
nand U45694 (N_45694,N_42001,N_43400);
nor U45695 (N_45695,N_43548,N_43650);
xor U45696 (N_45696,N_43439,N_42035);
or U45697 (N_45697,N_42986,N_43892);
xnor U45698 (N_45698,N_42569,N_43764);
and U45699 (N_45699,N_42012,N_43092);
xor U45700 (N_45700,N_43383,N_43497);
xnor U45701 (N_45701,N_43777,N_43335);
or U45702 (N_45702,N_43249,N_42709);
and U45703 (N_45703,N_42777,N_43850);
nor U45704 (N_45704,N_42914,N_42412);
nor U45705 (N_45705,N_43042,N_42568);
or U45706 (N_45706,N_43311,N_43727);
nand U45707 (N_45707,N_43227,N_43157);
and U45708 (N_45708,N_42047,N_42050);
nor U45709 (N_45709,N_43076,N_43912);
and U45710 (N_45710,N_43966,N_42890);
xor U45711 (N_45711,N_43051,N_42811);
nor U45712 (N_45712,N_42425,N_42562);
nand U45713 (N_45713,N_42747,N_42593);
nand U45714 (N_45714,N_43583,N_42845);
xnor U45715 (N_45715,N_42843,N_43290);
nand U45716 (N_45716,N_42806,N_42690);
nand U45717 (N_45717,N_43430,N_42870);
and U45718 (N_45718,N_42711,N_43136);
xnor U45719 (N_45719,N_43678,N_43776);
or U45720 (N_45720,N_43725,N_42057);
nand U45721 (N_45721,N_43895,N_42383);
nor U45722 (N_45722,N_43119,N_43092);
or U45723 (N_45723,N_42953,N_42332);
xor U45724 (N_45724,N_43700,N_43168);
nand U45725 (N_45725,N_42078,N_43272);
nand U45726 (N_45726,N_43405,N_43256);
or U45727 (N_45727,N_43275,N_42959);
nand U45728 (N_45728,N_43940,N_42153);
xor U45729 (N_45729,N_43152,N_42607);
nand U45730 (N_45730,N_43802,N_42716);
nand U45731 (N_45731,N_42392,N_42422);
xor U45732 (N_45732,N_42472,N_42162);
xor U45733 (N_45733,N_42396,N_43632);
and U45734 (N_45734,N_43375,N_43600);
and U45735 (N_45735,N_43480,N_42336);
and U45736 (N_45736,N_42452,N_42279);
and U45737 (N_45737,N_43247,N_43592);
nor U45738 (N_45738,N_43134,N_43067);
or U45739 (N_45739,N_42631,N_42641);
xnor U45740 (N_45740,N_43316,N_43857);
and U45741 (N_45741,N_42845,N_42996);
nor U45742 (N_45742,N_43793,N_42411);
xor U45743 (N_45743,N_43628,N_43735);
nor U45744 (N_45744,N_43904,N_43577);
nand U45745 (N_45745,N_42903,N_42804);
nor U45746 (N_45746,N_42429,N_43014);
xnor U45747 (N_45747,N_43195,N_43760);
and U45748 (N_45748,N_42109,N_43667);
or U45749 (N_45749,N_42280,N_43449);
and U45750 (N_45750,N_42313,N_42118);
and U45751 (N_45751,N_42104,N_43933);
nor U45752 (N_45752,N_42994,N_42935);
or U45753 (N_45753,N_43737,N_42316);
nor U45754 (N_45754,N_42530,N_43423);
nand U45755 (N_45755,N_42996,N_42432);
nand U45756 (N_45756,N_43044,N_42829);
nand U45757 (N_45757,N_43084,N_43776);
nand U45758 (N_45758,N_42131,N_43067);
or U45759 (N_45759,N_43890,N_43499);
and U45760 (N_45760,N_42433,N_42027);
and U45761 (N_45761,N_42003,N_43605);
nand U45762 (N_45762,N_42525,N_43371);
xnor U45763 (N_45763,N_42995,N_42573);
or U45764 (N_45764,N_43090,N_42022);
or U45765 (N_45765,N_43466,N_43046);
nand U45766 (N_45766,N_42755,N_42765);
nor U45767 (N_45767,N_42757,N_42102);
and U45768 (N_45768,N_42542,N_43624);
and U45769 (N_45769,N_42201,N_43414);
nor U45770 (N_45770,N_42292,N_43026);
xor U45771 (N_45771,N_42682,N_43908);
nand U45772 (N_45772,N_42074,N_42276);
nand U45773 (N_45773,N_42228,N_42234);
xnor U45774 (N_45774,N_42086,N_42734);
xor U45775 (N_45775,N_42274,N_43242);
nand U45776 (N_45776,N_42119,N_43257);
xor U45777 (N_45777,N_42624,N_42035);
nor U45778 (N_45778,N_43089,N_42531);
and U45779 (N_45779,N_42698,N_42847);
or U45780 (N_45780,N_43410,N_43873);
nor U45781 (N_45781,N_43926,N_43828);
nand U45782 (N_45782,N_42610,N_42484);
or U45783 (N_45783,N_43453,N_43728);
nor U45784 (N_45784,N_43483,N_43337);
and U45785 (N_45785,N_43000,N_42922);
and U45786 (N_45786,N_42319,N_42184);
and U45787 (N_45787,N_42511,N_42719);
xnor U45788 (N_45788,N_43340,N_42941);
and U45789 (N_45789,N_42647,N_42645);
nor U45790 (N_45790,N_43360,N_43499);
nand U45791 (N_45791,N_42855,N_43340);
or U45792 (N_45792,N_42186,N_42761);
nor U45793 (N_45793,N_43604,N_42537);
nor U45794 (N_45794,N_42098,N_42584);
and U45795 (N_45795,N_42207,N_43869);
or U45796 (N_45796,N_43979,N_42821);
nand U45797 (N_45797,N_42757,N_43547);
nand U45798 (N_45798,N_43022,N_42934);
or U45799 (N_45799,N_42513,N_43340);
and U45800 (N_45800,N_43310,N_42273);
xor U45801 (N_45801,N_43329,N_42744);
xnor U45802 (N_45802,N_42826,N_42028);
xnor U45803 (N_45803,N_43661,N_43830);
and U45804 (N_45804,N_43121,N_42194);
nor U45805 (N_45805,N_42872,N_42017);
or U45806 (N_45806,N_42727,N_43901);
xnor U45807 (N_45807,N_43389,N_43501);
or U45808 (N_45808,N_42945,N_43346);
xnor U45809 (N_45809,N_43251,N_42511);
xnor U45810 (N_45810,N_43167,N_42913);
nor U45811 (N_45811,N_42226,N_42200);
and U45812 (N_45812,N_42101,N_42754);
nand U45813 (N_45813,N_43217,N_42484);
and U45814 (N_45814,N_42364,N_43302);
nor U45815 (N_45815,N_42129,N_43525);
xnor U45816 (N_45816,N_42248,N_43304);
nor U45817 (N_45817,N_42176,N_43944);
nor U45818 (N_45818,N_42820,N_42314);
nor U45819 (N_45819,N_43344,N_43950);
xor U45820 (N_45820,N_42890,N_42285);
and U45821 (N_45821,N_42513,N_42120);
nand U45822 (N_45822,N_42712,N_42081);
nand U45823 (N_45823,N_43695,N_43219);
xor U45824 (N_45824,N_43396,N_43192);
nand U45825 (N_45825,N_43457,N_42161);
xnor U45826 (N_45826,N_43694,N_43755);
xor U45827 (N_45827,N_42800,N_42397);
nand U45828 (N_45828,N_42029,N_42062);
xnor U45829 (N_45829,N_43095,N_42537);
xor U45830 (N_45830,N_42074,N_43017);
and U45831 (N_45831,N_42296,N_43507);
nor U45832 (N_45832,N_42897,N_42284);
xnor U45833 (N_45833,N_43387,N_42805);
nor U45834 (N_45834,N_42666,N_42641);
xor U45835 (N_45835,N_43111,N_43452);
xor U45836 (N_45836,N_42540,N_42683);
or U45837 (N_45837,N_43659,N_42862);
nor U45838 (N_45838,N_42111,N_43445);
and U45839 (N_45839,N_42637,N_42812);
or U45840 (N_45840,N_43363,N_43844);
and U45841 (N_45841,N_43740,N_42173);
and U45842 (N_45842,N_42953,N_42464);
nor U45843 (N_45843,N_43821,N_42327);
or U45844 (N_45844,N_42332,N_42771);
or U45845 (N_45845,N_43675,N_43591);
nand U45846 (N_45846,N_43357,N_43684);
nor U45847 (N_45847,N_43446,N_42354);
and U45848 (N_45848,N_42036,N_43789);
nand U45849 (N_45849,N_42994,N_43295);
or U45850 (N_45850,N_43486,N_43036);
or U45851 (N_45851,N_43012,N_43754);
nor U45852 (N_45852,N_43694,N_43604);
nor U45853 (N_45853,N_42539,N_42914);
xor U45854 (N_45854,N_43166,N_43828);
and U45855 (N_45855,N_43311,N_42616);
or U45856 (N_45856,N_42867,N_43929);
nor U45857 (N_45857,N_42846,N_43090);
nor U45858 (N_45858,N_43013,N_43363);
xor U45859 (N_45859,N_43414,N_42754);
nor U45860 (N_45860,N_43928,N_42998);
nor U45861 (N_45861,N_42676,N_43332);
and U45862 (N_45862,N_43889,N_42977);
xnor U45863 (N_45863,N_42143,N_42727);
and U45864 (N_45864,N_43810,N_43519);
and U45865 (N_45865,N_43975,N_43144);
and U45866 (N_45866,N_42560,N_43160);
xnor U45867 (N_45867,N_43708,N_43860);
xor U45868 (N_45868,N_42804,N_42991);
nand U45869 (N_45869,N_42584,N_42342);
and U45870 (N_45870,N_42908,N_43095);
nor U45871 (N_45871,N_43419,N_43706);
or U45872 (N_45872,N_42830,N_42946);
nand U45873 (N_45873,N_43841,N_42546);
nor U45874 (N_45874,N_43361,N_43029);
and U45875 (N_45875,N_43355,N_42975);
nand U45876 (N_45876,N_42543,N_42321);
nand U45877 (N_45877,N_43637,N_43240);
and U45878 (N_45878,N_42362,N_43344);
nand U45879 (N_45879,N_42009,N_42626);
and U45880 (N_45880,N_42882,N_43760);
or U45881 (N_45881,N_43190,N_43693);
and U45882 (N_45882,N_43919,N_43313);
nor U45883 (N_45883,N_42799,N_43090);
xnor U45884 (N_45884,N_43063,N_43820);
or U45885 (N_45885,N_43721,N_42619);
nor U45886 (N_45886,N_42132,N_42516);
xor U45887 (N_45887,N_43522,N_43094);
nand U45888 (N_45888,N_43433,N_42574);
nor U45889 (N_45889,N_42942,N_43328);
or U45890 (N_45890,N_42498,N_43606);
or U45891 (N_45891,N_42119,N_42782);
nor U45892 (N_45892,N_43486,N_43387);
or U45893 (N_45893,N_42067,N_42700);
or U45894 (N_45894,N_43775,N_42918);
nor U45895 (N_45895,N_42591,N_43843);
xor U45896 (N_45896,N_42920,N_42945);
nand U45897 (N_45897,N_42282,N_43033);
xor U45898 (N_45898,N_42462,N_43481);
or U45899 (N_45899,N_42433,N_42669);
nor U45900 (N_45900,N_42146,N_42599);
and U45901 (N_45901,N_43972,N_42798);
nand U45902 (N_45902,N_42880,N_42943);
xor U45903 (N_45903,N_43010,N_42252);
xor U45904 (N_45904,N_43787,N_43213);
or U45905 (N_45905,N_43799,N_42555);
and U45906 (N_45906,N_43846,N_42643);
and U45907 (N_45907,N_43909,N_42933);
xor U45908 (N_45908,N_42322,N_43716);
or U45909 (N_45909,N_42716,N_42670);
and U45910 (N_45910,N_42039,N_43886);
and U45911 (N_45911,N_43224,N_43746);
and U45912 (N_45912,N_42893,N_42692);
or U45913 (N_45913,N_43853,N_42135);
or U45914 (N_45914,N_43394,N_42127);
and U45915 (N_45915,N_43940,N_42461);
nand U45916 (N_45916,N_42097,N_43162);
xor U45917 (N_45917,N_42602,N_43182);
or U45918 (N_45918,N_43528,N_42035);
xnor U45919 (N_45919,N_43850,N_42938);
or U45920 (N_45920,N_42713,N_42965);
xor U45921 (N_45921,N_42987,N_43889);
or U45922 (N_45922,N_43675,N_43157);
or U45923 (N_45923,N_42216,N_43714);
xnor U45924 (N_45924,N_43865,N_42402);
or U45925 (N_45925,N_43197,N_43928);
or U45926 (N_45926,N_42208,N_42759);
xnor U45927 (N_45927,N_42205,N_43296);
and U45928 (N_45928,N_42027,N_43965);
nand U45929 (N_45929,N_43474,N_42016);
xor U45930 (N_45930,N_42566,N_42354);
or U45931 (N_45931,N_43169,N_43594);
nand U45932 (N_45932,N_43665,N_42819);
nand U45933 (N_45933,N_42288,N_42570);
and U45934 (N_45934,N_42402,N_42978);
or U45935 (N_45935,N_42977,N_43355);
nor U45936 (N_45936,N_43575,N_42107);
nor U45937 (N_45937,N_43849,N_43330);
or U45938 (N_45938,N_42396,N_43260);
nor U45939 (N_45939,N_42803,N_43009);
xnor U45940 (N_45940,N_43322,N_43811);
nand U45941 (N_45941,N_42540,N_42378);
nor U45942 (N_45942,N_42548,N_43925);
xor U45943 (N_45943,N_43034,N_43876);
nand U45944 (N_45944,N_43025,N_42942);
or U45945 (N_45945,N_42791,N_43163);
or U45946 (N_45946,N_43607,N_43759);
xnor U45947 (N_45947,N_42543,N_43367);
and U45948 (N_45948,N_43644,N_43466);
nand U45949 (N_45949,N_42764,N_43471);
nand U45950 (N_45950,N_42228,N_43720);
xor U45951 (N_45951,N_42879,N_42951);
or U45952 (N_45952,N_43232,N_42850);
nor U45953 (N_45953,N_43699,N_42494);
xor U45954 (N_45954,N_42064,N_43201);
nor U45955 (N_45955,N_43981,N_42450);
and U45956 (N_45956,N_42342,N_42077);
xor U45957 (N_45957,N_43995,N_42985);
or U45958 (N_45958,N_42366,N_42127);
or U45959 (N_45959,N_42704,N_43777);
or U45960 (N_45960,N_43771,N_42365);
or U45961 (N_45961,N_43119,N_43544);
and U45962 (N_45962,N_42850,N_42549);
nor U45963 (N_45963,N_43656,N_42439);
or U45964 (N_45964,N_43431,N_42381);
or U45965 (N_45965,N_43169,N_42882);
or U45966 (N_45966,N_43244,N_42515);
xnor U45967 (N_45967,N_42526,N_43534);
or U45968 (N_45968,N_42768,N_43720);
and U45969 (N_45969,N_42657,N_43067);
and U45970 (N_45970,N_43992,N_42291);
nand U45971 (N_45971,N_43789,N_42855);
nand U45972 (N_45972,N_43880,N_42752);
nand U45973 (N_45973,N_43740,N_43927);
and U45974 (N_45974,N_42244,N_43458);
nor U45975 (N_45975,N_42193,N_42636);
nor U45976 (N_45976,N_43136,N_43759);
nor U45977 (N_45977,N_43850,N_43683);
and U45978 (N_45978,N_42260,N_43100);
and U45979 (N_45979,N_43131,N_43351);
nand U45980 (N_45980,N_43738,N_43895);
xnor U45981 (N_45981,N_42243,N_43609);
nand U45982 (N_45982,N_43275,N_43729);
and U45983 (N_45983,N_43145,N_43574);
and U45984 (N_45984,N_42279,N_43462);
and U45985 (N_45985,N_43290,N_42218);
nor U45986 (N_45986,N_42167,N_43367);
nand U45987 (N_45987,N_42469,N_42481);
xnor U45988 (N_45988,N_42363,N_42315);
or U45989 (N_45989,N_43390,N_42389);
nor U45990 (N_45990,N_43870,N_43749);
or U45991 (N_45991,N_42733,N_43504);
or U45992 (N_45992,N_42794,N_42569);
xnor U45993 (N_45993,N_43552,N_42059);
nor U45994 (N_45994,N_43449,N_43882);
and U45995 (N_45995,N_43512,N_42259);
xor U45996 (N_45996,N_43210,N_42915);
nand U45997 (N_45997,N_42869,N_43369);
and U45998 (N_45998,N_43971,N_42325);
nand U45999 (N_45999,N_43808,N_42111);
xor U46000 (N_46000,N_45559,N_44363);
xnor U46001 (N_46001,N_44793,N_45448);
xnor U46002 (N_46002,N_44509,N_45461);
nand U46003 (N_46003,N_44535,N_45647);
and U46004 (N_46004,N_44506,N_45710);
nand U46005 (N_46005,N_45832,N_45373);
nand U46006 (N_46006,N_45189,N_44142);
nand U46007 (N_46007,N_45483,N_44634);
and U46008 (N_46008,N_45631,N_45219);
xor U46009 (N_46009,N_44338,N_45503);
or U46010 (N_46010,N_44359,N_45689);
or U46011 (N_46011,N_45825,N_44252);
nor U46012 (N_46012,N_45978,N_44273);
or U46013 (N_46013,N_44976,N_45768);
nand U46014 (N_46014,N_45520,N_45255);
or U46015 (N_46015,N_44556,N_44477);
nor U46016 (N_46016,N_44092,N_44456);
or U46017 (N_46017,N_45963,N_44182);
xnor U46018 (N_46018,N_45338,N_44345);
or U46019 (N_46019,N_45034,N_45927);
and U46020 (N_46020,N_44179,N_44137);
xor U46021 (N_46021,N_44451,N_44813);
or U46022 (N_46022,N_45014,N_45252);
nor U46023 (N_46023,N_45551,N_44545);
and U46024 (N_46024,N_44406,N_45964);
nor U46025 (N_46025,N_45342,N_44340);
xor U46026 (N_46026,N_45104,N_45542);
nor U46027 (N_46027,N_44757,N_44081);
nand U46028 (N_46028,N_45755,N_45835);
nand U46029 (N_46029,N_44669,N_44730);
nor U46030 (N_46030,N_45114,N_44377);
nor U46031 (N_46031,N_44573,N_44581);
nor U46032 (N_46032,N_44411,N_45350);
and U46033 (N_46033,N_44471,N_44143);
xnor U46034 (N_46034,N_45422,N_45567);
and U46035 (N_46035,N_44693,N_45327);
and U46036 (N_46036,N_45848,N_44957);
nand U46037 (N_46037,N_45119,N_44498);
and U46038 (N_46038,N_45495,N_44438);
xor U46039 (N_46039,N_44020,N_45696);
and U46040 (N_46040,N_45596,N_45188);
nand U46041 (N_46041,N_44098,N_44825);
and U46042 (N_46042,N_45013,N_45180);
nand U46043 (N_46043,N_44915,N_45721);
nand U46044 (N_46044,N_45820,N_44246);
xor U46045 (N_46045,N_45929,N_44880);
or U46046 (N_46046,N_44871,N_44970);
nand U46047 (N_46047,N_45836,N_45815);
nand U46048 (N_46048,N_45008,N_45377);
nor U46049 (N_46049,N_44741,N_45829);
or U46050 (N_46050,N_44085,N_45256);
or U46051 (N_46051,N_45749,N_44572);
or U46052 (N_46052,N_44433,N_44938);
nand U46053 (N_46053,N_45995,N_45310);
or U46054 (N_46054,N_45068,N_44313);
nor U46055 (N_46055,N_44155,N_45365);
nand U46056 (N_46056,N_45867,N_44106);
xor U46057 (N_46057,N_45385,N_45282);
or U46058 (N_46058,N_44758,N_45741);
nand U46059 (N_46059,N_44360,N_45702);
or U46060 (N_46060,N_44470,N_44718);
nor U46061 (N_46061,N_44019,N_45799);
nor U46062 (N_46062,N_45692,N_44689);
or U46063 (N_46063,N_45113,N_44474);
xor U46064 (N_46064,N_45878,N_45270);
xor U46065 (N_46065,N_45415,N_45630);
nand U46066 (N_46066,N_45445,N_44251);
or U46067 (N_46067,N_45807,N_44427);
nor U46068 (N_46068,N_44337,N_45881);
xor U46069 (N_46069,N_44074,N_45475);
nor U46070 (N_46070,N_44479,N_45744);
nand U46071 (N_46071,N_45145,N_45213);
nor U46072 (N_46072,N_44888,N_45913);
or U46073 (N_46073,N_44962,N_44829);
and U46074 (N_46074,N_45683,N_44589);
nand U46075 (N_46075,N_44401,N_44692);
nor U46076 (N_46076,N_44435,N_44442);
or U46077 (N_46077,N_44512,N_44141);
and U46078 (N_46078,N_44196,N_45165);
or U46079 (N_46079,N_44705,N_45044);
nor U46080 (N_46080,N_44980,N_45439);
xnor U46081 (N_46081,N_44995,N_44950);
nor U46082 (N_46082,N_44253,N_45552);
xor U46083 (N_46083,N_45306,N_44817);
and U46084 (N_46084,N_45223,N_45750);
nor U46085 (N_46085,N_44316,N_44090);
or U46086 (N_46086,N_45039,N_44447);
xor U46087 (N_46087,N_45061,N_45684);
and U46088 (N_46088,N_44408,N_44744);
and U46089 (N_46089,N_45669,N_45970);
nand U46090 (N_46090,N_45981,N_44868);
xor U46091 (N_46091,N_45915,N_45833);
nand U46092 (N_46092,N_45923,N_44002);
or U46093 (N_46093,N_44102,N_44886);
and U46094 (N_46094,N_45147,N_44862);
xor U46095 (N_46095,N_45328,N_44614);
xnor U46096 (N_46096,N_44563,N_44358);
nor U46097 (N_46097,N_44462,N_45257);
and U46098 (N_46098,N_44894,N_44844);
or U46099 (N_46099,N_44169,N_44079);
or U46100 (N_46100,N_44985,N_45058);
and U46101 (N_46101,N_44336,N_45758);
xnor U46102 (N_46102,N_44680,N_44655);
nand U46103 (N_46103,N_45419,N_44603);
nor U46104 (N_46104,N_45616,N_44561);
or U46105 (N_46105,N_44626,N_44518);
and U46106 (N_46106,N_45183,N_44230);
and U46107 (N_46107,N_44071,N_44217);
nor U46108 (N_46108,N_44500,N_45731);
or U46109 (N_46109,N_45679,N_44224);
xnor U46110 (N_46110,N_44089,N_44211);
nor U46111 (N_46111,N_44875,N_44769);
nor U46112 (N_46112,N_45378,N_44931);
or U46113 (N_46113,N_45850,N_45229);
xnor U46114 (N_46114,N_44028,N_45046);
nand U46115 (N_46115,N_44575,N_45421);
nand U46116 (N_46116,N_44215,N_45688);
or U46117 (N_46117,N_45837,N_44147);
or U46118 (N_46118,N_44440,N_45716);
nand U46119 (N_46119,N_45018,N_45776);
nor U46120 (N_46120,N_45124,N_45813);
xor U46121 (N_46121,N_44299,N_44233);
nor U46122 (N_46122,N_44391,N_45116);
xor U46123 (N_46123,N_45239,N_45091);
xor U46124 (N_46124,N_44870,N_45766);
and U46125 (N_46125,N_44944,N_44134);
xor U46126 (N_46126,N_45979,N_45621);
xnor U46127 (N_46127,N_44084,N_44538);
nand U46128 (N_46128,N_45823,N_44181);
or U46129 (N_46129,N_45737,N_44428);
nand U46130 (N_46130,N_44667,N_45198);
nor U46131 (N_46131,N_45764,N_44052);
nand U46132 (N_46132,N_45759,N_44854);
xnor U46133 (N_46133,N_44687,N_45957);
xor U46134 (N_46134,N_45700,N_45535);
and U46135 (N_46135,N_44012,N_45901);
and U46136 (N_46136,N_45537,N_45889);
nor U46137 (N_46137,N_44262,N_45109);
or U46138 (N_46138,N_44178,N_44135);
nand U46139 (N_46139,N_44612,N_44986);
xor U46140 (N_46140,N_44530,N_44108);
and U46141 (N_46141,N_45747,N_44000);
nand U46142 (N_46142,N_44896,N_45990);
xnor U46143 (N_46143,N_44170,N_44841);
nor U46144 (N_46144,N_45453,N_44367);
or U46145 (N_46145,N_44180,N_45938);
nor U46146 (N_46146,N_45222,N_45397);
xnor U46147 (N_46147,N_45356,N_45292);
and U46148 (N_46148,N_45101,N_45316);
nand U46149 (N_46149,N_44790,N_44908);
or U46150 (N_46150,N_45612,N_45676);
or U46151 (N_46151,N_45548,N_45933);
or U46152 (N_46152,N_44984,N_45406);
or U46153 (N_46153,N_44963,N_44992);
or U46154 (N_46154,N_45089,N_44587);
xnor U46155 (N_46155,N_44704,N_44569);
xnor U46156 (N_46156,N_44752,N_44192);
nand U46157 (N_46157,N_45886,N_45900);
or U46158 (N_46158,N_44907,N_44925);
or U46159 (N_46159,N_44959,N_45863);
or U46160 (N_46160,N_44505,N_44328);
or U46161 (N_46161,N_44370,N_45462);
xnor U46162 (N_46162,N_44499,N_44786);
or U46163 (N_46163,N_44241,N_44351);
xor U46164 (N_46164,N_45481,N_44623);
and U46165 (N_46165,N_44651,N_44111);
nand U46166 (N_46166,N_45125,N_44808);
nor U46167 (N_46167,N_44866,N_45795);
nand U46168 (N_46168,N_44945,N_44318);
nor U46169 (N_46169,N_44076,N_44026);
nand U46170 (N_46170,N_45533,N_44759);
and U46171 (N_46171,N_44195,N_44383);
xnor U46172 (N_46172,N_45059,N_45278);
nor U46173 (N_46173,N_44240,N_44777);
nor U46174 (N_46174,N_44812,N_44403);
and U46175 (N_46175,N_44782,N_45589);
nand U46176 (N_46176,N_44099,N_44014);
nor U46177 (N_46177,N_44172,N_44764);
nand U46178 (N_46178,N_45617,N_44625);
xor U46179 (N_46179,N_45186,N_45505);
xor U46180 (N_46180,N_45479,N_44835);
xor U46181 (N_46181,N_44128,N_44123);
xnor U46182 (N_46182,N_44309,N_45335);
and U46183 (N_46183,N_45429,N_44225);
or U46184 (N_46184,N_45580,N_45975);
nor U46185 (N_46185,N_45959,N_44784);
nand U46186 (N_46186,N_44465,N_45530);
xor U46187 (N_46187,N_45088,N_44158);
nor U46188 (N_46188,N_45332,N_44577);
nand U46189 (N_46189,N_45137,N_44642);
and U46190 (N_46190,N_45494,N_45296);
and U46191 (N_46191,N_45723,N_44036);
and U46192 (N_46192,N_44469,N_45802);
or U46193 (N_46193,N_45396,N_45334);
and U46194 (N_46194,N_45674,N_44672);
xor U46195 (N_46195,N_44326,N_45910);
and U46196 (N_46196,N_44308,N_44130);
nor U46197 (N_46197,N_44031,N_44413);
nand U46198 (N_46198,N_45115,N_45940);
or U46199 (N_46199,N_44348,N_44046);
xnor U46200 (N_46200,N_45469,N_45887);
nand U46201 (N_46201,N_45809,N_44657);
and U46202 (N_46202,N_44549,N_45320);
and U46203 (N_46203,N_44867,N_45062);
xor U46204 (N_46204,N_45380,N_45038);
or U46205 (N_46205,N_45681,N_45553);
nor U46206 (N_46206,N_44724,N_44293);
nand U46207 (N_46207,N_44366,N_45499);
and U46208 (N_46208,N_45288,N_44912);
nand U46209 (N_46209,N_45425,N_45171);
or U46210 (N_46210,N_44885,N_44901);
nand U46211 (N_46211,N_45030,N_44390);
nor U46212 (N_46212,N_45295,N_45208);
and U46213 (N_46213,N_44231,N_45403);
and U46214 (N_46214,N_45247,N_45591);
nand U46215 (N_46215,N_45740,N_45751);
nand U46216 (N_46216,N_45660,N_45563);
nand U46217 (N_46217,N_45917,N_44774);
xor U46218 (N_46218,N_44503,N_45491);
nand U46219 (N_46219,N_44117,N_44703);
or U46220 (N_46220,N_44124,N_44558);
or U46221 (N_46221,N_44480,N_45374);
nor U46222 (N_46222,N_44132,N_44668);
nor U46223 (N_46223,N_44942,N_44746);
xor U46224 (N_46224,N_44616,N_44039);
or U46225 (N_46225,N_45321,N_44576);
nand U46226 (N_46226,N_44062,N_45950);
xnor U46227 (N_46227,N_45080,N_44017);
xnor U46228 (N_46228,N_45426,N_45642);
xor U46229 (N_46229,N_45918,N_44087);
nor U46230 (N_46230,N_45644,N_45160);
nand U46231 (N_46231,N_44997,N_44260);
nand U46232 (N_46232,N_45811,N_45906);
nand U46233 (N_46233,N_44740,N_45523);
nand U46234 (N_46234,N_45201,N_45339);
nor U46235 (N_46235,N_44156,N_44802);
or U46236 (N_46236,N_44965,N_45845);
and U46237 (N_46237,N_45128,N_45271);
and U46238 (N_46238,N_44727,N_44795);
or U46239 (N_46239,N_44129,N_44484);
and U46240 (N_46240,N_44537,N_45476);
nor U46241 (N_46241,N_44315,N_44638);
or U46242 (N_46242,N_44362,N_45251);
nand U46243 (N_46243,N_45079,N_44635);
or U46244 (N_46244,N_45007,N_44464);
or U46245 (N_46245,N_45036,N_45955);
and U46246 (N_46246,N_45844,N_44881);
nor U46247 (N_46247,N_44785,N_45760);
nor U46248 (N_46248,N_44787,N_45827);
and U46249 (N_46249,N_45985,N_44685);
xnor U46250 (N_46250,N_44374,N_45178);
and U46251 (N_46251,N_44199,N_45191);
xor U46252 (N_46252,N_44991,N_44415);
and U46253 (N_46253,N_45680,N_44566);
or U46254 (N_46254,N_45055,N_44522);
nor U46255 (N_46255,N_44323,N_45389);
xor U46256 (N_46256,N_45690,N_45362);
or U46257 (N_46257,N_44726,N_44977);
or U46258 (N_46258,N_45797,N_45947);
xor U46259 (N_46259,N_44275,N_44475);
nor U46260 (N_46260,N_44996,N_44119);
xnor U46261 (N_46261,N_44792,N_44357);
xnor U46262 (N_46262,N_45440,N_44677);
nor U46263 (N_46263,N_44654,N_45211);
or U46264 (N_46264,N_45607,N_45071);
xnor U46265 (N_46265,N_44443,N_45383);
or U46266 (N_46266,N_44906,N_44204);
nor U46267 (N_46267,N_44399,N_45218);
nor U46268 (N_46268,N_44698,N_44206);
nand U46269 (N_46269,N_44828,N_45333);
or U46270 (N_46270,N_45808,N_44463);
or U46271 (N_46271,N_45077,N_44482);
nor U46272 (N_46272,N_45122,N_45216);
or U46273 (N_46273,N_45274,N_44640);
and U46274 (N_46274,N_44734,N_44183);
nand U46275 (N_46275,N_45942,N_45875);
or U46276 (N_46276,N_45199,N_44096);
nand U46277 (N_46277,N_45769,N_45926);
nand U46278 (N_46278,N_44524,N_44218);
nand U46279 (N_46279,N_45965,N_44115);
nand U46280 (N_46280,N_45595,N_44882);
nor U46281 (N_46281,N_44521,N_44534);
or U46282 (N_46282,N_44565,N_44059);
or U46283 (N_46283,N_44053,N_45694);
and U46284 (N_46284,N_44816,N_44139);
nand U46285 (N_46285,N_45574,N_44619);
and U46286 (N_46286,N_45347,N_44420);
xor U46287 (N_46287,N_45463,N_45883);
nor U46288 (N_46288,N_45516,N_44258);
xnor U46289 (N_46289,N_44045,N_45245);
or U46290 (N_46290,N_45118,N_45381);
nor U46291 (N_46291,N_45614,N_44571);
xor U46292 (N_46292,N_44259,N_44686);
or U46293 (N_46293,N_44822,N_44305);
nand U46294 (N_46294,N_44282,N_45096);
nand U46295 (N_46295,N_45562,N_45279);
xnor U46296 (N_46296,N_44617,N_45954);
and U46297 (N_46297,N_45106,N_44319);
nand U46298 (N_46298,N_44653,N_45572);
xnor U46299 (N_46299,N_44818,N_45675);
nor U46300 (N_46300,N_44520,N_44583);
or U46301 (N_46301,N_44335,N_44244);
xor U46302 (N_46302,N_45063,N_44922);
nor U46303 (N_46303,N_44780,N_45816);
and U46304 (N_46304,N_44320,N_45914);
or U46305 (N_46305,N_45443,N_44903);
or U46306 (N_46306,N_44389,N_44030);
xor U46307 (N_46307,N_44820,N_44437);
nand U46308 (N_46308,N_44298,N_44238);
or U46309 (N_46309,N_44941,N_45051);
and U46310 (N_46310,N_44037,N_45961);
or U46311 (N_46311,N_45507,N_44051);
nand U46312 (N_46312,N_45812,N_45531);
xor U46313 (N_46313,N_44673,N_44765);
and U46314 (N_46314,N_45163,N_44212);
and U46315 (N_46315,N_44064,N_45485);
or U46316 (N_46316,N_44190,N_44201);
nand U46317 (N_46317,N_44890,N_44150);
nand U46318 (N_46318,N_44250,N_44656);
or U46319 (N_46319,N_44519,N_44236);
nand U46320 (N_46320,N_45538,N_44112);
nand U46321 (N_46321,N_44398,N_44879);
and U46322 (N_46322,N_44690,N_45635);
or U46323 (N_46323,N_45015,N_44277);
xor U46324 (N_46324,N_45289,N_44494);
nor U46325 (N_46325,N_44376,N_44436);
nor U46326 (N_46326,N_44666,N_44781);
xor U46327 (N_46327,N_44618,N_45130);
nor U46328 (N_46328,N_44501,N_45800);
and U46329 (N_46329,N_45040,N_45301);
and U46330 (N_46330,N_45772,N_45922);
and U46331 (N_46331,N_45801,N_45496);
and U46332 (N_46332,N_45949,N_45127);
and U46333 (N_46333,N_44833,N_45826);
nor U46334 (N_46334,N_44314,N_45952);
nor U46335 (N_46335,N_45262,N_45539);
nand U46336 (N_46336,N_45739,N_44193);
or U46337 (N_46337,N_45637,N_44956);
nor U46338 (N_46338,N_44968,N_45204);
or U46339 (N_46339,N_45509,N_45154);
xor U46340 (N_46340,N_44060,N_44184);
nand U46341 (N_46341,N_44173,N_44900);
nand U46342 (N_46342,N_44247,N_44773);
or U46343 (N_46343,N_45187,N_45623);
nand U46344 (N_46344,N_45341,N_44859);
and U46345 (N_46345,N_45956,N_44550);
nand U46346 (N_46346,N_44738,N_45012);
nand U46347 (N_46347,N_45597,N_45110);
and U46348 (N_46348,N_45546,N_45627);
or U46349 (N_46349,N_45451,N_44902);
xnor U46350 (N_46350,N_44473,N_45794);
nand U46351 (N_46351,N_45578,N_44929);
xor U46352 (N_46352,N_44707,N_44272);
and U46353 (N_46353,N_45076,N_45212);
or U46354 (N_46354,N_45624,N_45100);
nor U46355 (N_46355,N_44160,N_45065);
nand U46356 (N_46356,N_45558,N_44432);
xor U46357 (N_46357,N_45294,N_45930);
xnor U46358 (N_46358,N_45151,N_44557);
xnor U46359 (N_46359,N_45131,N_44861);
or U46360 (N_46360,N_44801,N_45010);
nor U46361 (N_46361,N_44009,N_44049);
and U46362 (N_46362,N_44600,N_44761);
or U46363 (N_46363,N_44989,N_45515);
xnor U46364 (N_46364,N_44610,N_45763);
nand U46365 (N_46365,N_45444,N_45277);
and U46366 (N_46366,N_45474,N_44836);
and U46367 (N_46367,N_45142,N_44189);
and U46368 (N_46368,N_44267,N_44283);
and U46369 (N_46369,N_44865,N_44485);
or U46370 (N_46370,N_45220,N_45756);
or U46371 (N_46371,N_45659,N_45242);
nand U46372 (N_46372,N_44013,N_44416);
nor U46373 (N_46373,N_45235,N_45898);
xnor U46374 (N_46374,N_44466,N_45719);
and U46375 (N_46375,N_44453,N_44152);
nor U46376 (N_46376,N_45035,N_44120);
nor U46377 (N_46377,N_44307,N_44756);
xor U46378 (N_46378,N_45579,N_44384);
and U46379 (N_46379,N_45911,N_45093);
nor U46380 (N_46380,N_44203,N_45330);
xor U46381 (N_46381,N_45784,N_44213);
and U46382 (N_46382,N_44636,N_44927);
nor U46383 (N_46383,N_44100,N_45632);
nand U46384 (N_46384,N_45518,N_44332);
or U46385 (N_46385,N_44716,N_44797);
and U46386 (N_46386,N_44011,N_44597);
nor U46387 (N_46387,N_44033,N_45004);
nor U46388 (N_46388,N_45384,N_44921);
xor U46389 (N_46389,N_44527,N_45834);
nor U46390 (N_46390,N_44632,N_45770);
nand U46391 (N_46391,N_44091,N_44385);
and U46392 (N_46392,N_45028,N_45874);
nand U46393 (N_46393,N_44732,N_45584);
nor U46394 (N_46394,N_44819,N_44711);
xnor U46395 (N_46395,N_45796,N_44850);
or U46396 (N_46396,N_45701,N_45896);
or U46397 (N_46397,N_45753,N_44257);
xor U46398 (N_46398,N_45715,N_44973);
or U46399 (N_46399,N_44719,N_45798);
or U46400 (N_46400,N_44895,N_45268);
xor U46401 (N_46401,N_45438,N_45042);
xor U46402 (N_46402,N_45117,N_45728);
nand U46403 (N_46403,N_44429,N_44864);
nand U46404 (N_46404,N_45661,N_45522);
xor U46405 (N_46405,N_45905,N_45904);
and U46406 (N_46406,N_45138,N_44198);
nor U46407 (N_46407,N_44271,N_45067);
or U46408 (N_46408,N_45454,N_45746);
xor U46409 (N_46409,N_45269,N_45236);
and U46410 (N_46410,N_45169,N_45312);
xor U46411 (N_46411,N_45907,N_45313);
xnor U46412 (N_46412,N_45738,N_44960);
nand U46413 (N_46413,N_44486,N_45394);
nand U46414 (N_46414,N_45276,N_44953);
and U46415 (N_46415,N_44419,N_45792);
and U46416 (N_46416,N_45785,N_45555);
or U46417 (N_46417,N_44776,N_44729);
or U46418 (N_46418,N_44842,N_45167);
nand U46419 (N_46419,N_45969,N_44721);
or U46420 (N_46420,N_45317,N_45407);
or U46421 (N_46421,N_44916,N_45166);
nand U46422 (N_46422,N_44266,N_45363);
nor U46423 (N_46423,N_45032,N_45678);
and U46424 (N_46424,N_45500,N_45576);
nand U46425 (N_46425,N_45240,N_45273);
nor U46426 (N_46426,N_45023,N_44426);
nor U46427 (N_46427,N_44609,N_44523);
and U46428 (N_46428,N_44015,N_45105);
nand U46429 (N_46429,N_44811,N_45361);
nor U46430 (N_46430,N_45243,N_45983);
nand U46431 (N_46431,N_45937,N_45078);
and U46432 (N_46432,N_44167,N_44884);
nor U46433 (N_46433,N_45634,N_44388);
xnor U46434 (N_46434,N_45368,N_44676);
xor U46435 (N_46435,N_45549,N_45090);
and U46436 (N_46436,N_44932,N_44430);
nand U46437 (N_46437,N_45254,N_44994);
nor U46438 (N_46438,N_44660,N_44110);
nand U46439 (N_46439,N_45352,N_44274);
and U46440 (N_46440,N_45082,N_45314);
or U46441 (N_46441,N_45976,N_44736);
or U46442 (N_46442,N_45250,N_44449);
nor U46443 (N_46443,N_45309,N_44291);
or U46444 (N_46444,N_44683,N_44295);
and U46445 (N_46445,N_44939,N_45893);
and U46446 (N_46446,N_45851,N_44967);
nor U46447 (N_46447,N_45490,N_45121);
nor U46448 (N_46448,N_45604,N_44745);
or U46449 (N_46449,N_45852,N_45666);
or U46450 (N_46450,N_44094,N_44688);
or U46451 (N_46451,N_45311,N_44659);
nand U46452 (N_46452,N_45541,N_45876);
xor U46453 (N_46453,N_44754,N_44439);
xnor U46454 (N_46454,N_45944,N_44005);
and U46455 (N_46455,N_45967,N_45050);
nand U46456 (N_46456,N_45217,N_45416);
nor U46457 (N_46457,N_45966,N_44590);
or U46458 (N_46458,N_45399,N_44472);
nor U46459 (N_46459,N_44254,N_45550);
and U46460 (N_46460,N_44947,N_44528);
or U46461 (N_46461,N_45290,N_44508);
xor U46462 (N_46462,N_44568,N_45457);
xnor U46463 (N_46463,N_44214,N_45265);
nor U46464 (N_46464,N_45771,N_45935);
nand U46465 (N_46465,N_45720,N_44940);
nor U46466 (N_46466,N_45971,N_44814);
nand U46467 (N_46467,N_44375,N_44007);
nand U46468 (N_46468,N_45497,N_45297);
xor U46469 (N_46469,N_45083,N_45564);
nand U46470 (N_46470,N_45074,N_44604);
xor U46471 (N_46471,N_45506,N_44431);
and U46472 (N_46472,N_44993,N_45467);
xor U46473 (N_46473,N_44424,N_44905);
or U46474 (N_46474,N_45258,N_44234);
or U46475 (N_46475,N_45691,N_44845);
nand U46476 (N_46476,N_44974,N_44027);
nand U46477 (N_46477,N_45951,N_44652);
nor U46478 (N_46478,N_44460,N_44481);
xnor U46479 (N_46479,N_45711,N_44622);
or U46480 (N_46480,N_44446,N_45434);
xor U46481 (N_46481,N_45318,N_44559);
nor U46482 (N_46482,N_44872,N_44760);
nor U46483 (N_46483,N_45645,N_45566);
nand U46484 (N_46484,N_45980,N_44101);
nor U46485 (N_46485,N_45858,N_45354);
nand U46486 (N_46486,N_45962,N_45184);
xor U46487 (N_46487,N_45909,N_44713);
nand U46488 (N_46488,N_44798,N_44306);
nand U46489 (N_46489,N_44047,N_44333);
nor U46490 (N_46490,N_44560,N_44114);
or U46491 (N_46491,N_45355,N_45471);
xor U46492 (N_46492,N_44006,N_45838);
nor U46493 (N_46493,N_45307,N_44001);
nor U46494 (N_46494,N_44961,N_45185);
xor U46495 (N_46495,N_45215,N_45478);
or U46496 (N_46496,N_44457,N_44770);
nor U46497 (N_46497,N_45281,N_45112);
and U46498 (N_46498,N_45323,N_45427);
nor U46499 (N_46499,N_45757,N_45388);
nor U46500 (N_46500,N_44382,N_45441);
or U46501 (N_46501,N_44564,N_45775);
or U46502 (N_46502,N_44067,N_45968);
or U46503 (N_46503,N_44645,N_44422);
xor U46504 (N_46504,N_44934,N_45646);
and U46505 (N_46505,N_44018,N_45141);
xor U46506 (N_46506,N_44159,N_45779);
and U46507 (N_46507,N_45284,N_45103);
nor U46508 (N_46508,N_45417,N_44300);
nor U46509 (N_46509,N_44830,N_45026);
xor U46510 (N_46510,N_44596,N_45094);
or U46511 (N_46511,N_45987,N_45302);
and U46512 (N_46512,N_44526,N_44983);
nand U46513 (N_46513,N_45366,N_45897);
nand U46514 (N_46514,N_45123,N_45400);
nor U46515 (N_46515,N_44138,N_44517);
or U46516 (N_46516,N_44441,N_45369);
nor U46517 (N_46517,N_44136,N_45272);
xor U46518 (N_46518,N_45590,N_44022);
and U46519 (N_46519,N_45871,N_44856);
or U46520 (N_46520,N_44343,N_45859);
or U46521 (N_46521,N_44088,N_45864);
or U46522 (N_46522,N_44725,N_44848);
nand U46523 (N_46523,N_45392,N_45280);
xor U46524 (N_46524,N_45993,N_44361);
nand U46525 (N_46525,N_45070,N_45371);
and U46526 (N_46526,N_44086,N_45345);
nand U46527 (N_46527,N_45598,N_45214);
xor U46528 (N_46528,N_44296,N_44407);
nor U46529 (N_46529,N_45393,N_44342);
nor U46530 (N_46530,N_44324,N_44372);
xor U46531 (N_46531,N_44630,N_44665);
nor U46532 (N_46532,N_44873,N_45919);
nand U46533 (N_46533,N_44171,N_45654);
and U46534 (N_46534,N_44514,N_44352);
and U46535 (N_46535,N_45736,N_45207);
nand U46536 (N_46536,N_44551,N_45402);
xor U46537 (N_46537,N_44548,N_45504);
or U46538 (N_46538,N_44321,N_45465);
xor U46539 (N_46539,N_44988,N_45587);
nand U46540 (N_46540,N_45846,N_45560);
or U46541 (N_46541,N_44177,N_45882);
xnor U46542 (N_46542,N_45888,N_44346);
or U46543 (N_46543,N_45508,N_44029);
nand U46544 (N_46544,N_45570,N_44536);
and U46545 (N_46545,N_44380,N_45525);
or U46546 (N_46546,N_45673,N_45638);
nor U46547 (N_46547,N_45027,N_44418);
and U46548 (N_46548,N_44552,N_45787);
or U46549 (N_46549,N_45636,N_45743);
xor U46550 (N_46550,N_45197,N_44855);
xor U46551 (N_46551,N_44126,N_45041);
xor U46552 (N_46552,N_45781,N_44948);
and U46553 (N_46553,N_44113,N_45872);
nand U46554 (N_46554,N_44131,N_44919);
xor U46555 (N_46555,N_44735,N_44631);
nand U46556 (N_46556,N_44851,N_44396);
or U46557 (N_46557,N_44368,N_45622);
nand U46558 (N_46558,N_45565,N_45351);
nand U46559 (N_46559,N_45657,N_45568);
or U46560 (N_46560,N_44237,N_44601);
nor U46561 (N_46561,N_45134,N_45618);
and U46562 (N_46562,N_45275,N_44349);
or U46563 (N_46563,N_45011,N_44369);
nand U46564 (N_46564,N_45873,N_45605);
xor U46565 (N_46565,N_45860,N_44904);
nor U46566 (N_46566,N_44068,N_44289);
nand U46567 (N_46567,N_44731,N_45890);
or U46568 (N_46568,N_45176,N_45266);
xnor U46569 (N_46569,N_44010,N_44292);
and U46570 (N_46570,N_45583,N_44926);
or U46571 (N_46571,N_44174,N_45821);
nor U46572 (N_46572,N_44290,N_45626);
xor U46573 (N_46573,N_44284,N_44297);
nand U46574 (N_46574,N_44355,N_44082);
or U46575 (N_46575,N_44602,N_44699);
and U46576 (N_46576,N_45658,N_45725);
xor U46577 (N_46577,N_44393,N_44897);
nor U46578 (N_46578,N_45047,N_44701);
xnor U46579 (N_46579,N_44910,N_45732);
nand U46580 (N_46580,N_45401,N_44235);
xnor U46581 (N_46581,N_44853,N_45582);
nor U46582 (N_46582,N_44330,N_44525);
nand U46583 (N_46583,N_45708,N_45994);
nand U46584 (N_46584,N_45810,N_44400);
and U46585 (N_46585,N_44834,N_44467);
nor U46586 (N_46586,N_45581,N_44643);
nand U46587 (N_46587,N_44691,N_45020);
nand U46588 (N_46588,N_44809,N_44365);
xor U46589 (N_46589,N_45423,N_45175);
and U46590 (N_46590,N_44706,N_44048);
and U46591 (N_46591,N_44476,N_44806);
and U46592 (N_46592,N_44621,N_44341);
and U46593 (N_46593,N_45726,N_44887);
nand U46594 (N_46594,N_45037,N_45754);
or U46595 (N_46595,N_44728,N_44280);
nand U46596 (N_46596,N_44662,N_44869);
or U46597 (N_46597,N_45002,N_44971);
nor U46598 (N_46598,N_45226,N_45428);
nand U46599 (N_46599,N_45891,N_45953);
or U46600 (N_46600,N_45843,N_44205);
xnor U46601 (N_46601,N_44531,N_44070);
xor U46602 (N_46602,N_44347,N_45652);
nand U46603 (N_46603,N_45510,N_45016);
or U46604 (N_46604,N_44496,N_44924);
and U46605 (N_46605,N_45655,N_45899);
and U46606 (N_46606,N_44301,N_44043);
nand U46607 (N_46607,N_44788,N_44826);
nor U46608 (N_46608,N_44220,N_45724);
xnor U46609 (N_46609,N_45298,N_44946);
xnor U46610 (N_46610,N_44543,N_45432);
or U46611 (N_46611,N_45231,N_44981);
and U46612 (N_46612,N_44423,N_44796);
xor U46613 (N_46613,N_44107,N_44849);
xor U46614 (N_46614,N_44952,N_44185);
nor U46615 (N_46615,N_45557,N_44743);
or U46616 (N_46616,N_44075,N_45486);
or U46617 (N_46617,N_44857,N_44317);
nor U46618 (N_46618,N_44145,N_44878);
or U46619 (N_46619,N_45129,N_44458);
nand U46620 (N_46620,N_44495,N_44387);
or U46621 (N_46621,N_44574,N_45611);
nor U46622 (N_46622,N_44595,N_44344);
nand U46623 (N_46623,N_44216,N_44539);
nand U46624 (N_46624,N_44133,N_44186);
nand U46625 (N_46625,N_45409,N_44935);
or U46626 (N_46626,N_45477,N_44288);
xnor U46627 (N_46627,N_44371,N_44491);
nand U46628 (N_46628,N_45865,N_44302);
nand U46629 (N_46629,N_45870,N_45085);
nand U46630 (N_46630,N_44709,N_45326);
or U46631 (N_46631,N_44151,N_44846);
or U46632 (N_46632,N_44261,N_44414);
nor U46633 (N_46633,N_45228,N_45999);
and U46634 (N_46634,N_45466,N_44570);
xnor U46635 (N_46635,N_45482,N_45346);
or U46636 (N_46636,N_44584,N_45806);
and U46637 (N_46637,N_44444,N_44620);
nor U46638 (N_46638,N_45161,N_44483);
or U46639 (N_46639,N_45603,N_44154);
nand U46640 (N_46640,N_44116,N_44327);
and U46641 (N_46641,N_45149,N_45536);
or U46642 (N_46642,N_44546,N_44165);
or U46643 (N_46643,N_44737,N_45936);
xnor U46644 (N_46644,N_44930,N_45609);
and U46645 (N_46645,N_44035,N_45649);
and U46646 (N_46646,N_45305,N_45502);
and U46647 (N_46647,N_45722,N_44805);
nand U46648 (N_46648,N_44807,N_44647);
nor U46649 (N_46649,N_45672,N_44242);
and U46650 (N_46650,N_45945,N_45487);
nand U46651 (N_46651,N_44840,N_45585);
nand U46652 (N_46652,N_45903,N_45547);
nor U46653 (N_46653,N_45248,N_45224);
nand U46654 (N_46654,N_44594,N_45375);
xor U46655 (N_46655,N_45519,N_45348);
or U46656 (N_46656,N_45249,N_44937);
xnor U46657 (N_46657,N_44078,N_44755);
and U46658 (N_46658,N_45267,N_45600);
or U46659 (N_46659,N_44207,N_45000);
nand U46660 (N_46660,N_45493,N_44386);
xor U46661 (N_46661,N_45343,N_45991);
and U46662 (N_46662,N_45158,N_44162);
nor U46663 (N_46663,N_44334,N_45643);
nor U46664 (N_46664,N_45073,N_44717);
nor U46665 (N_46665,N_44544,N_44733);
nor U46666 (N_46666,N_45285,N_45822);
nand U46667 (N_46667,N_45379,N_45430);
nor U46668 (N_46668,N_45748,N_45592);
xor U46669 (N_46669,N_45468,N_45264);
nand U46670 (N_46670,N_45005,N_45641);
and U46671 (N_46671,N_45237,N_44628);
nand U46672 (N_46672,N_44789,N_45190);
and U46673 (N_46673,N_45856,N_44516);
xnor U46674 (N_46674,N_45286,N_44061);
nor U46675 (N_46675,N_45048,N_44489);
nand U46676 (N_46676,N_45620,N_45594);
xnor U46677 (N_46677,N_44379,N_45029);
xor U46678 (N_46678,N_45625,N_44219);
nor U46679 (N_46679,N_44459,N_44268);
or U46680 (N_46680,N_45452,N_45304);
or U46681 (N_46681,N_45608,N_45412);
or U46682 (N_46682,N_44109,N_45752);
and U46683 (N_46683,N_45569,N_45916);
and U46684 (N_46684,N_45705,N_44753);
nand U46685 (N_46685,N_45144,N_45060);
xor U46686 (N_46686,N_44394,N_45733);
nand U46687 (N_46687,N_45033,N_45436);
xor U46688 (N_46688,N_44883,N_44540);
nor U46689 (N_46689,N_44354,N_45984);
and U46690 (N_46690,N_44256,N_45447);
xor U46691 (N_46691,N_44056,N_45706);
nand U46692 (N_46692,N_45238,N_45168);
nor U46693 (N_46693,N_44125,N_44492);
xor U46694 (N_46694,N_45988,N_45413);
xor U46695 (N_46695,N_44402,N_44964);
nor U46696 (N_46696,N_45449,N_45411);
nand U46697 (N_46697,N_44339,N_45619);
and U46698 (N_46698,N_45606,N_45717);
xnor U46699 (N_46699,N_44800,N_45824);
nand U46700 (N_46700,N_45671,N_44695);
or U46701 (N_46701,N_44228,N_44032);
xor U46702 (N_46702,N_44751,N_45472);
xnor U46703 (N_46703,N_44933,N_44913);
xnor U46704 (N_46704,N_44767,N_45908);
or U46705 (N_46705,N_44050,N_44679);
or U46706 (N_46706,N_44990,N_45790);
xor U46707 (N_46707,N_45610,N_45765);
xor U46708 (N_46708,N_44194,N_45948);
xnor U46709 (N_46709,N_45545,N_44200);
or U46710 (N_46710,N_45892,N_45712);
nand U46711 (N_46711,N_45331,N_45941);
xor U46712 (N_46712,N_44077,N_44004);
or U46713 (N_46713,N_45767,N_45200);
or U46714 (N_46714,N_44507,N_45081);
nor U46715 (N_46715,N_45524,N_45098);
nor U46716 (N_46716,N_45227,N_44763);
xnor U46717 (N_46717,N_45571,N_44448);
and U46718 (N_46718,N_45804,N_44898);
nand U46719 (N_46719,N_45202,N_45958);
or U46720 (N_46720,N_45849,N_44409);
and U46721 (N_46721,N_44712,N_44294);
nor U46722 (N_46722,N_44421,N_45205);
and U46723 (N_46723,N_45177,N_45513);
or U46724 (N_46724,N_45853,N_45868);
or U46725 (N_46725,N_45925,N_44541);
nor U46726 (N_46726,N_45932,N_44649);
xnor U46727 (N_46727,N_44255,N_44281);
nor U46728 (N_46728,N_45066,N_45287);
or U46729 (N_46729,N_44264,N_45006);
nor U46730 (N_46730,N_44768,N_44891);
xor U46731 (N_46731,N_45783,N_45360);
and U46732 (N_46732,N_44226,N_44972);
and U46733 (N_46733,N_45456,N_44663);
and U46734 (N_46734,N_44003,N_45450);
nor U46735 (N_46735,N_45291,N_44187);
and U46736 (N_46736,N_45157,N_45132);
xor U46737 (N_46737,N_44608,N_44410);
and U46738 (N_46738,N_44310,N_44304);
nor U46739 (N_46739,N_45774,N_44815);
and U46740 (N_46740,N_44696,N_45172);
nor U46741 (N_46741,N_44069,N_44877);
nand U46742 (N_46742,N_45556,N_45126);
and U46743 (N_46743,N_44127,N_45260);
and U46744 (N_46744,N_44779,N_44063);
nand U46745 (N_46745,N_45152,N_45862);
or U46746 (N_46746,N_44502,N_44148);
and U46747 (N_46747,N_44949,N_45102);
nand U46748 (N_46748,N_44708,N_44747);
or U46749 (N_46749,N_44762,N_44831);
xnor U46750 (N_46750,N_45195,N_45470);
xor U46751 (N_46751,N_45839,N_44658);
xor U46752 (N_46752,N_45593,N_45857);
and U46753 (N_46753,N_45424,N_45069);
xor U46754 (N_46754,N_45001,N_45727);
nand U46755 (N_46755,N_44248,N_45075);
nand U46756 (N_46756,N_45931,N_45140);
xnor U46757 (N_46757,N_44176,N_45458);
or U46758 (N_46758,N_44555,N_45639);
and U46759 (N_46759,N_45107,N_44105);
xnor U46760 (N_46760,N_44454,N_44923);
nor U46761 (N_46761,N_44714,N_44852);
xnor U46762 (N_46762,N_45025,N_45133);
nand U46763 (N_46763,N_44876,N_44331);
nand U46764 (N_46764,N_45996,N_44263);
and U46765 (N_46765,N_45884,N_45805);
xor U46766 (N_46766,N_44080,N_44287);
nor U46767 (N_46767,N_45376,N_45773);
nor U46768 (N_46768,N_44661,N_45340);
nor U46769 (N_46769,N_45232,N_44243);
xor U46770 (N_46770,N_45293,N_45554);
nor U46771 (N_46771,N_45484,N_45283);
xnor U46772 (N_46772,N_45729,N_44468);
nor U46773 (N_46773,N_44582,N_44627);
xnor U46774 (N_46774,N_44221,N_45819);
xor U46775 (N_46775,N_44153,N_44095);
xnor U46776 (N_46776,N_44839,N_44038);
xnor U46777 (N_46777,N_45651,N_44395);
or U46778 (N_46778,N_45511,N_45344);
nor U46779 (N_46779,N_44593,N_44412);
nand U46780 (N_46780,N_44425,N_44392);
nor U46781 (N_46781,N_45253,N_45150);
or U46782 (N_46782,N_44356,N_45599);
or U46783 (N_46783,N_44821,N_45761);
or U46784 (N_46784,N_45687,N_45446);
nand U46785 (N_46785,N_45387,N_44311);
nor U46786 (N_46786,N_45745,N_45540);
or U46787 (N_46787,N_45367,N_44682);
or U46788 (N_46788,N_45322,N_45517);
xnor U46789 (N_46789,N_44513,N_45885);
or U46790 (N_46790,N_44073,N_44715);
xor U46791 (N_46791,N_45442,N_45629);
and U46792 (N_46792,N_45788,N_45939);
and U46793 (N_46793,N_45529,N_45698);
xor U46794 (N_46794,N_44325,N_44223);
or U46795 (N_46795,N_45390,N_45973);
nand U46796 (N_46796,N_45372,N_45512);
nand U46797 (N_46797,N_45992,N_45364);
xor U46798 (N_46798,N_44598,N_44588);
nor U46799 (N_46799,N_44847,N_45977);
xor U46800 (N_46800,N_44918,N_44208);
and U46801 (N_46801,N_44097,N_45532);
nand U46802 (N_46802,N_45841,N_45686);
nor U46803 (N_46803,N_45193,N_45847);
and U46804 (N_46804,N_45049,N_45814);
or U46805 (N_46805,N_45241,N_44586);
and U46806 (N_46806,N_45489,N_44312);
nor U46807 (N_46807,N_45398,N_45668);
nor U46808 (N_46808,N_44700,N_44766);
or U46809 (N_46809,N_44269,N_45695);
nor U46810 (N_46810,N_45086,N_44585);
or U46811 (N_46811,N_44911,N_45209);
nor U46812 (N_46812,N_45464,N_44804);
nand U46813 (N_46813,N_44547,N_44794);
xor U46814 (N_46814,N_45043,N_45182);
or U46815 (N_46815,N_45780,N_44748);
xor U46816 (N_46816,N_45924,N_44232);
and U46817 (N_46817,N_44674,N_45210);
xor U46818 (N_46818,N_45817,N_45386);
xor U46819 (N_46819,N_45246,N_45714);
nand U46820 (N_46820,N_44648,N_44975);
nand U46821 (N_46821,N_44042,N_45943);
xnor U46822 (N_46822,N_44276,N_44533);
xnor U46823 (N_46823,N_44197,N_45206);
nor U46824 (N_46824,N_45986,N_45056);
xnor U46825 (N_46825,N_44605,N_44860);
or U46826 (N_46826,N_44592,N_45418);
and U46827 (N_46827,N_44008,N_45433);
nand U46828 (N_46828,N_44055,N_45174);
xnor U46829 (N_46829,N_45960,N_44044);
nand U46830 (N_46830,N_44710,N_45455);
xor U46831 (N_46831,N_45640,N_44373);
nor U46832 (N_46832,N_44720,N_45017);
nand U46833 (N_46833,N_44065,N_45382);
nand U46834 (N_46834,N_44943,N_45778);
nand U46835 (N_46835,N_44810,N_44646);
or U46836 (N_46836,N_45713,N_44510);
nand U46837 (N_46837,N_45156,N_44529);
and U46838 (N_46838,N_44149,N_45358);
nor U46839 (N_46839,N_44493,N_44562);
nand U46840 (N_46840,N_44553,N_45734);
or U46841 (N_46841,N_45791,N_44863);
or U46842 (N_46842,N_44611,N_44771);
or U46843 (N_46843,N_44103,N_45325);
nor U46844 (N_46844,N_45019,N_45633);
nor U46845 (N_46845,N_45982,N_45677);
or U46846 (N_46846,N_44858,N_44664);
or U46847 (N_46847,N_44675,N_45003);
nand U46848 (N_46848,N_44161,N_45912);
nand U46849 (N_46849,N_44778,N_45704);
nand U46850 (N_46850,N_45742,N_45087);
or U46851 (N_46851,N_44697,N_44054);
and U46852 (N_46852,N_45414,N_45064);
nor U46853 (N_46853,N_44278,N_44966);
and U46854 (N_46854,N_45097,N_45707);
and U46855 (N_46855,N_44874,N_45664);
nor U46856 (N_46856,N_44982,N_45009);
and U46857 (N_46857,N_45699,N_44969);
xnor U46858 (N_46858,N_45492,N_44121);
xor U46859 (N_46859,N_44144,N_45300);
and U46860 (N_46860,N_45173,N_44265);
and U46861 (N_46861,N_44381,N_44772);
and U46862 (N_46862,N_45601,N_45586);
nand U46863 (N_46863,N_45998,N_45244);
nand U46864 (N_46864,N_45072,N_44364);
and U46865 (N_46865,N_45920,N_45934);
and U46866 (N_46866,N_44227,N_45135);
and U46867 (N_46867,N_45588,N_45179);
xor U46868 (N_46868,N_44920,N_44058);
nor U46869 (N_46869,N_45120,N_45053);
nand U46870 (N_46870,N_45842,N_45308);
nor U46871 (N_46871,N_44554,N_45139);
or U46872 (N_46872,N_44578,N_44515);
xor U46873 (N_46873,N_44670,N_45895);
and U46874 (N_46874,N_45840,N_45391);
nand U46875 (N_46875,N_45024,N_44249);
nor U46876 (N_46876,N_44580,N_44742);
nor U46877 (N_46877,N_45703,N_44567);
and U46878 (N_46878,N_45359,N_45682);
and U46879 (N_46879,N_45946,N_44951);
nand U46880 (N_46880,N_44057,N_45315);
xnor U46881 (N_46881,N_45880,N_44955);
and U46882 (N_46882,N_44025,N_44914);
nand U46883 (N_46883,N_45789,N_45303);
and U46884 (N_46884,N_44791,N_44824);
xor U46885 (N_46885,N_44450,N_45902);
xnor U46886 (N_46886,N_44461,N_45861);
or U46887 (N_46887,N_44633,N_44021);
nand U46888 (N_46888,N_45099,N_45561);
or U46889 (N_46889,N_45437,N_45498);
xnor U46890 (N_46890,N_44999,N_44532);
and U46891 (N_46891,N_44629,N_45777);
nor U46892 (N_46892,N_44639,N_45111);
and U46893 (N_46893,N_44749,N_44093);
xnor U46894 (N_46894,N_45057,N_45196);
nor U46895 (N_46895,N_45573,N_44163);
nor U46896 (N_46896,N_44040,N_45663);
xnor U46897 (N_46897,N_45735,N_45473);
and U46898 (N_46898,N_45460,N_44202);
nor U46899 (N_46899,N_44329,N_45997);
or U46900 (N_46900,N_45337,N_45162);
nand U46901 (N_46901,N_45718,N_44405);
nand U46902 (N_46902,N_44893,N_45225);
nor U46903 (N_46903,N_45782,N_44239);
xor U46904 (N_46904,N_44285,N_45408);
nor U46905 (N_46905,N_45974,N_44209);
nor U46906 (N_46906,N_45431,N_44445);
xor U46907 (N_46907,N_45084,N_45527);
nand U46908 (N_46908,N_45155,N_45543);
nor U46909 (N_46909,N_45170,N_45855);
xor U46910 (N_46910,N_45762,N_44229);
xnor U46911 (N_46911,N_45615,N_45866);
xor U46912 (N_46912,N_44455,N_45793);
nand U46913 (N_46913,N_45092,N_44838);
nand U46914 (N_46914,N_45665,N_45052);
or U46915 (N_46915,N_44417,N_44397);
or U46916 (N_46916,N_45667,N_45420);
and U46917 (N_46917,N_45685,N_44591);
or U46918 (N_46918,N_45299,N_45528);
nor U46919 (N_46919,N_44650,N_45628);
or U46920 (N_46920,N_45234,N_45324);
nor U46921 (N_46921,N_45670,N_44024);
nor U46922 (N_46922,N_45319,N_45146);
nand U46923 (N_46923,N_45021,N_44579);
and U46924 (N_46924,N_44799,N_44958);
or U46925 (N_46925,N_44353,N_45730);
nand U46926 (N_46926,N_44140,N_44641);
xor U46927 (N_46927,N_45869,N_45830);
or U46928 (N_46928,N_45410,N_45230);
nor U46929 (N_46929,N_44998,N_45192);
and U46930 (N_46930,N_44624,N_45159);
nor U46931 (N_46931,N_44889,N_45194);
nand U46932 (N_46932,N_45404,N_44615);
or U46933 (N_46933,N_45349,N_45164);
and U46934 (N_46934,N_44637,N_45693);
nor U46935 (N_46935,N_44434,N_44511);
and U46936 (N_46936,N_45045,N_44488);
or U46937 (N_46937,N_45648,N_44322);
xnor U46938 (N_46938,N_44175,N_45263);
nand U46939 (N_46939,N_45575,N_44542);
nor U46940 (N_46940,N_44210,N_45697);
nor U46941 (N_46941,N_44490,N_44452);
or U46942 (N_46942,N_44504,N_45577);
nor U46943 (N_46943,N_44909,N_44164);
or U46944 (N_46944,N_45709,N_44606);
or U46945 (N_46945,N_45544,N_44613);
and U46946 (N_46946,N_44750,N_45329);
or U46947 (N_46947,N_45031,N_44684);
nor U46948 (N_46948,N_44899,N_45357);
nand U46949 (N_46949,N_44644,N_45989);
xnor U46950 (N_46950,N_45928,N_45514);
nor U46951 (N_46951,N_45662,N_45353);
nand U46952 (N_46952,N_45972,N_44083);
nand U46953 (N_46953,N_45108,N_45613);
nor U46954 (N_46954,N_44723,N_45203);
and U46955 (N_46955,N_44122,N_45921);
nand U46956 (N_46956,N_44279,N_44832);
nand U46957 (N_46957,N_44378,N_44478);
nor U46958 (N_46958,N_44350,N_45054);
and U46959 (N_46959,N_45526,N_45405);
xnor U46960 (N_46960,N_45459,N_44803);
or U46961 (N_46961,N_44739,N_44286);
and U46962 (N_46962,N_45153,N_45879);
xor U46963 (N_46963,N_44843,N_45831);
nand U46964 (N_46964,N_44671,N_44245);
and U46965 (N_46965,N_45854,N_44270);
or U46966 (N_46966,N_45233,N_45650);
xor U46967 (N_46967,N_45803,N_44487);
nand U46968 (N_46968,N_44404,N_45435);
and U46969 (N_46969,N_45521,N_45261);
nor U46970 (N_46970,N_44607,N_44837);
nor U46971 (N_46971,N_45181,N_45602);
or U46972 (N_46972,N_44016,N_45022);
nor U46973 (N_46973,N_45259,N_45877);
or U46974 (N_46974,N_44694,N_44827);
nor U46975 (N_46975,N_44978,N_44023);
nor U46976 (N_46976,N_44191,N_44157);
nand U46977 (N_46977,N_45501,N_44166);
and U46978 (N_46978,N_44979,N_45818);
xnor U46979 (N_46979,N_44917,N_45395);
xnor U46980 (N_46980,N_44072,N_44303);
xnor U46981 (N_46981,N_44823,N_45370);
xor U46982 (N_46982,N_45828,N_44775);
nor U46983 (N_46983,N_44146,N_44928);
or U46984 (N_46984,N_44104,N_44892);
xnor U46985 (N_46985,N_44722,N_45894);
or U46986 (N_46986,N_45148,N_45221);
nand U46987 (N_46987,N_45143,N_45488);
nor U46988 (N_46988,N_45136,N_45786);
nand U46989 (N_46989,N_45095,N_45656);
xor U46990 (N_46990,N_45480,N_44034);
nor U46991 (N_46991,N_44954,N_44188);
nand U46992 (N_46992,N_45653,N_44681);
xnor U46993 (N_46993,N_44599,N_44168);
and U46994 (N_46994,N_44987,N_44783);
nand U46995 (N_46995,N_44118,N_44678);
nand U46996 (N_46996,N_44222,N_44497);
and U46997 (N_46997,N_44936,N_44066);
nor U46998 (N_46998,N_45534,N_45336);
or U46999 (N_46999,N_44702,N_44041);
and U47000 (N_47000,N_44511,N_44929);
and U47001 (N_47001,N_45769,N_45683);
or U47002 (N_47002,N_44293,N_45450);
or U47003 (N_47003,N_44682,N_44044);
and U47004 (N_47004,N_45502,N_44366);
xor U47005 (N_47005,N_45718,N_44000);
nand U47006 (N_47006,N_45305,N_44740);
or U47007 (N_47007,N_45068,N_45245);
nand U47008 (N_47008,N_44783,N_44800);
nand U47009 (N_47009,N_45912,N_45329);
or U47010 (N_47010,N_45390,N_44302);
nand U47011 (N_47011,N_44258,N_44722);
nand U47012 (N_47012,N_45017,N_45877);
nor U47013 (N_47013,N_44467,N_44100);
nand U47014 (N_47014,N_44898,N_45994);
nor U47015 (N_47015,N_45026,N_44175);
nor U47016 (N_47016,N_45020,N_44037);
nand U47017 (N_47017,N_45456,N_44952);
nor U47018 (N_47018,N_44770,N_44961);
nand U47019 (N_47019,N_45682,N_45747);
xor U47020 (N_47020,N_44578,N_44002);
or U47021 (N_47021,N_44891,N_45603);
nor U47022 (N_47022,N_44715,N_45528);
or U47023 (N_47023,N_45362,N_45809);
nor U47024 (N_47024,N_45735,N_45831);
or U47025 (N_47025,N_45355,N_44199);
and U47026 (N_47026,N_44628,N_45264);
xor U47027 (N_47027,N_45666,N_45776);
nand U47028 (N_47028,N_45486,N_44928);
or U47029 (N_47029,N_44207,N_45230);
and U47030 (N_47030,N_45103,N_44877);
nor U47031 (N_47031,N_44511,N_45229);
nand U47032 (N_47032,N_44939,N_44657);
and U47033 (N_47033,N_44998,N_45556);
nand U47034 (N_47034,N_45412,N_45629);
nand U47035 (N_47035,N_45259,N_44732);
nor U47036 (N_47036,N_44851,N_45117);
xnor U47037 (N_47037,N_44362,N_44487);
and U47038 (N_47038,N_44678,N_45658);
xnor U47039 (N_47039,N_44434,N_44573);
nand U47040 (N_47040,N_44940,N_45470);
and U47041 (N_47041,N_44719,N_44599);
and U47042 (N_47042,N_44294,N_44398);
xnor U47043 (N_47043,N_45509,N_45735);
and U47044 (N_47044,N_45030,N_44473);
xor U47045 (N_47045,N_45730,N_44412);
xnor U47046 (N_47046,N_44879,N_44409);
and U47047 (N_47047,N_44804,N_44501);
and U47048 (N_47048,N_45445,N_44676);
xnor U47049 (N_47049,N_45343,N_45113);
and U47050 (N_47050,N_44890,N_45347);
and U47051 (N_47051,N_44526,N_44582);
xor U47052 (N_47052,N_44397,N_44804);
and U47053 (N_47053,N_45212,N_44067);
or U47054 (N_47054,N_44063,N_45041);
or U47055 (N_47055,N_45930,N_44434);
nor U47056 (N_47056,N_44588,N_45705);
nor U47057 (N_47057,N_45692,N_45536);
or U47058 (N_47058,N_45444,N_44062);
and U47059 (N_47059,N_45758,N_45585);
nor U47060 (N_47060,N_44030,N_44031);
nand U47061 (N_47061,N_45410,N_44126);
or U47062 (N_47062,N_45524,N_45665);
and U47063 (N_47063,N_45970,N_45603);
and U47064 (N_47064,N_44155,N_45204);
xor U47065 (N_47065,N_45977,N_45515);
or U47066 (N_47066,N_44638,N_45233);
xor U47067 (N_47067,N_45000,N_44831);
nor U47068 (N_47068,N_45232,N_44326);
xnor U47069 (N_47069,N_45049,N_45420);
xor U47070 (N_47070,N_44125,N_44530);
and U47071 (N_47071,N_45271,N_44173);
nand U47072 (N_47072,N_44417,N_45777);
xnor U47073 (N_47073,N_45045,N_45723);
and U47074 (N_47074,N_44577,N_45484);
nor U47075 (N_47075,N_44747,N_44371);
or U47076 (N_47076,N_44609,N_44588);
nand U47077 (N_47077,N_45163,N_45823);
xnor U47078 (N_47078,N_44328,N_44494);
and U47079 (N_47079,N_44789,N_45447);
or U47080 (N_47080,N_44968,N_44090);
and U47081 (N_47081,N_44951,N_45572);
nand U47082 (N_47082,N_44870,N_44428);
nor U47083 (N_47083,N_44742,N_44698);
or U47084 (N_47084,N_44403,N_44144);
nand U47085 (N_47085,N_45361,N_45861);
and U47086 (N_47086,N_44418,N_45547);
and U47087 (N_47087,N_45514,N_44166);
and U47088 (N_47088,N_45022,N_44841);
and U47089 (N_47089,N_45277,N_44089);
xor U47090 (N_47090,N_45875,N_45075);
nor U47091 (N_47091,N_45195,N_45277);
nand U47092 (N_47092,N_45917,N_44022);
xor U47093 (N_47093,N_45782,N_45294);
nor U47094 (N_47094,N_44665,N_45227);
and U47095 (N_47095,N_44617,N_44020);
or U47096 (N_47096,N_45488,N_44790);
or U47097 (N_47097,N_44666,N_44905);
xnor U47098 (N_47098,N_45568,N_45061);
xnor U47099 (N_47099,N_44272,N_44746);
nor U47100 (N_47100,N_44144,N_45673);
and U47101 (N_47101,N_44640,N_45204);
and U47102 (N_47102,N_45983,N_44267);
xnor U47103 (N_47103,N_44842,N_44624);
xor U47104 (N_47104,N_45109,N_44353);
or U47105 (N_47105,N_44498,N_44831);
and U47106 (N_47106,N_45110,N_45828);
xnor U47107 (N_47107,N_44875,N_45230);
and U47108 (N_47108,N_44751,N_45509);
xnor U47109 (N_47109,N_45426,N_44614);
and U47110 (N_47110,N_45261,N_45437);
and U47111 (N_47111,N_45197,N_45677);
xnor U47112 (N_47112,N_45400,N_45827);
nor U47113 (N_47113,N_45714,N_45354);
or U47114 (N_47114,N_45440,N_45525);
nand U47115 (N_47115,N_44177,N_44287);
nor U47116 (N_47116,N_45908,N_44258);
nor U47117 (N_47117,N_45089,N_45305);
or U47118 (N_47118,N_44128,N_45833);
xnor U47119 (N_47119,N_44488,N_44309);
and U47120 (N_47120,N_45566,N_44016);
or U47121 (N_47121,N_44390,N_44610);
nor U47122 (N_47122,N_44113,N_45586);
and U47123 (N_47123,N_44230,N_45882);
or U47124 (N_47124,N_44009,N_44563);
xor U47125 (N_47125,N_44653,N_45943);
and U47126 (N_47126,N_44223,N_44153);
nand U47127 (N_47127,N_44253,N_44415);
and U47128 (N_47128,N_44610,N_44502);
xnor U47129 (N_47129,N_44363,N_45067);
or U47130 (N_47130,N_45388,N_45665);
nor U47131 (N_47131,N_45709,N_45100);
nand U47132 (N_47132,N_44750,N_44055);
and U47133 (N_47133,N_44046,N_45956);
xnor U47134 (N_47134,N_44380,N_45356);
or U47135 (N_47135,N_44961,N_44035);
nand U47136 (N_47136,N_45486,N_44051);
and U47137 (N_47137,N_44857,N_45717);
xor U47138 (N_47138,N_45062,N_44546);
or U47139 (N_47139,N_45683,N_45546);
xor U47140 (N_47140,N_44104,N_45492);
or U47141 (N_47141,N_44369,N_45851);
xor U47142 (N_47142,N_44034,N_45154);
nand U47143 (N_47143,N_44087,N_44621);
and U47144 (N_47144,N_45172,N_45020);
nor U47145 (N_47145,N_44581,N_44879);
or U47146 (N_47146,N_45313,N_44918);
and U47147 (N_47147,N_45704,N_44374);
xnor U47148 (N_47148,N_44902,N_45716);
and U47149 (N_47149,N_44604,N_45517);
and U47150 (N_47150,N_44353,N_45126);
xnor U47151 (N_47151,N_44089,N_45964);
or U47152 (N_47152,N_45505,N_45788);
nor U47153 (N_47153,N_44500,N_45021);
and U47154 (N_47154,N_44838,N_44370);
xor U47155 (N_47155,N_45028,N_44977);
nand U47156 (N_47156,N_44998,N_44817);
nor U47157 (N_47157,N_45335,N_45713);
xor U47158 (N_47158,N_44392,N_45210);
nand U47159 (N_47159,N_44475,N_44327);
and U47160 (N_47160,N_44682,N_44151);
or U47161 (N_47161,N_45655,N_45153);
or U47162 (N_47162,N_45569,N_44796);
and U47163 (N_47163,N_44480,N_45154);
nor U47164 (N_47164,N_45572,N_44763);
or U47165 (N_47165,N_45303,N_45371);
and U47166 (N_47166,N_45736,N_45139);
or U47167 (N_47167,N_45760,N_45459);
nor U47168 (N_47168,N_44732,N_44765);
nor U47169 (N_47169,N_45328,N_44413);
nor U47170 (N_47170,N_45061,N_44314);
or U47171 (N_47171,N_45560,N_45150);
or U47172 (N_47172,N_45776,N_45246);
nor U47173 (N_47173,N_44111,N_44993);
nor U47174 (N_47174,N_45403,N_44527);
and U47175 (N_47175,N_45416,N_45992);
xnor U47176 (N_47176,N_45998,N_44386);
nor U47177 (N_47177,N_44979,N_45880);
nand U47178 (N_47178,N_44046,N_44780);
xor U47179 (N_47179,N_44171,N_45297);
nor U47180 (N_47180,N_45493,N_45340);
nand U47181 (N_47181,N_45785,N_45200);
nand U47182 (N_47182,N_45807,N_45387);
xor U47183 (N_47183,N_44026,N_44863);
xor U47184 (N_47184,N_45102,N_44382);
xnor U47185 (N_47185,N_44999,N_44989);
or U47186 (N_47186,N_44255,N_44794);
xor U47187 (N_47187,N_44627,N_45073);
xnor U47188 (N_47188,N_45810,N_44160);
nand U47189 (N_47189,N_45701,N_45599);
nand U47190 (N_47190,N_45686,N_44522);
and U47191 (N_47191,N_45594,N_44343);
and U47192 (N_47192,N_45500,N_44124);
nand U47193 (N_47193,N_44673,N_45677);
nor U47194 (N_47194,N_44045,N_45653);
nand U47195 (N_47195,N_44868,N_45134);
and U47196 (N_47196,N_44535,N_45465);
nor U47197 (N_47197,N_44902,N_44503);
nor U47198 (N_47198,N_44928,N_45038);
nand U47199 (N_47199,N_44155,N_45494);
or U47200 (N_47200,N_45225,N_45543);
or U47201 (N_47201,N_45574,N_45527);
and U47202 (N_47202,N_44516,N_44780);
xor U47203 (N_47203,N_45337,N_45579);
or U47204 (N_47204,N_44364,N_44182);
and U47205 (N_47205,N_45409,N_44841);
xnor U47206 (N_47206,N_44868,N_44690);
and U47207 (N_47207,N_45961,N_44047);
nand U47208 (N_47208,N_45654,N_45582);
xnor U47209 (N_47209,N_45795,N_45364);
nand U47210 (N_47210,N_44975,N_45750);
xnor U47211 (N_47211,N_45930,N_44819);
nand U47212 (N_47212,N_45029,N_44341);
nand U47213 (N_47213,N_44126,N_45690);
xnor U47214 (N_47214,N_44240,N_44844);
nor U47215 (N_47215,N_45219,N_45417);
nand U47216 (N_47216,N_44433,N_44678);
nor U47217 (N_47217,N_44247,N_44938);
nor U47218 (N_47218,N_45545,N_45303);
nor U47219 (N_47219,N_44917,N_44203);
or U47220 (N_47220,N_44759,N_44181);
nand U47221 (N_47221,N_44398,N_44091);
nor U47222 (N_47222,N_44736,N_44083);
nand U47223 (N_47223,N_45274,N_45205);
or U47224 (N_47224,N_45187,N_44960);
nor U47225 (N_47225,N_45512,N_45505);
and U47226 (N_47226,N_45277,N_45920);
xnor U47227 (N_47227,N_45605,N_45578);
and U47228 (N_47228,N_45622,N_44869);
nand U47229 (N_47229,N_44412,N_44209);
nand U47230 (N_47230,N_44932,N_44012);
or U47231 (N_47231,N_45508,N_44794);
and U47232 (N_47232,N_45140,N_45733);
and U47233 (N_47233,N_45262,N_45978);
or U47234 (N_47234,N_44052,N_44861);
nor U47235 (N_47235,N_45681,N_45279);
or U47236 (N_47236,N_44176,N_44855);
and U47237 (N_47237,N_44685,N_45320);
xor U47238 (N_47238,N_44076,N_45507);
xor U47239 (N_47239,N_44691,N_44324);
xor U47240 (N_47240,N_45524,N_44186);
nor U47241 (N_47241,N_45709,N_45789);
and U47242 (N_47242,N_45890,N_44329);
nor U47243 (N_47243,N_45197,N_45027);
nand U47244 (N_47244,N_45887,N_45715);
and U47245 (N_47245,N_44658,N_45377);
and U47246 (N_47246,N_44542,N_45680);
nor U47247 (N_47247,N_44578,N_45333);
and U47248 (N_47248,N_45647,N_44253);
nand U47249 (N_47249,N_45084,N_45105);
nand U47250 (N_47250,N_45293,N_45402);
nand U47251 (N_47251,N_45981,N_45980);
nand U47252 (N_47252,N_45185,N_45694);
nand U47253 (N_47253,N_44005,N_44012);
and U47254 (N_47254,N_45307,N_45577);
xor U47255 (N_47255,N_45170,N_44642);
nor U47256 (N_47256,N_45526,N_45628);
or U47257 (N_47257,N_44034,N_45719);
and U47258 (N_47258,N_44682,N_45976);
nand U47259 (N_47259,N_45049,N_45288);
or U47260 (N_47260,N_45724,N_45725);
xor U47261 (N_47261,N_45569,N_44177);
and U47262 (N_47262,N_44933,N_44437);
xnor U47263 (N_47263,N_44760,N_45344);
nand U47264 (N_47264,N_44492,N_45124);
or U47265 (N_47265,N_45559,N_45997);
nand U47266 (N_47266,N_44774,N_45271);
xor U47267 (N_47267,N_44486,N_45186);
nand U47268 (N_47268,N_45435,N_44523);
nand U47269 (N_47269,N_45088,N_44587);
xor U47270 (N_47270,N_44641,N_44991);
nor U47271 (N_47271,N_44507,N_45240);
nor U47272 (N_47272,N_45110,N_44246);
and U47273 (N_47273,N_44842,N_45503);
or U47274 (N_47274,N_45029,N_44845);
xnor U47275 (N_47275,N_44193,N_44223);
or U47276 (N_47276,N_45120,N_44108);
or U47277 (N_47277,N_44658,N_45942);
xnor U47278 (N_47278,N_45867,N_45946);
xnor U47279 (N_47279,N_44618,N_45874);
nor U47280 (N_47280,N_45901,N_44928);
nor U47281 (N_47281,N_45488,N_44936);
and U47282 (N_47282,N_44596,N_45319);
nand U47283 (N_47283,N_45533,N_44205);
xor U47284 (N_47284,N_44563,N_44196);
xnor U47285 (N_47285,N_45450,N_45739);
and U47286 (N_47286,N_45987,N_44441);
nand U47287 (N_47287,N_44002,N_45531);
xnor U47288 (N_47288,N_44403,N_44132);
and U47289 (N_47289,N_44541,N_44789);
xor U47290 (N_47290,N_44496,N_45320);
nor U47291 (N_47291,N_44617,N_45953);
xnor U47292 (N_47292,N_45645,N_45873);
and U47293 (N_47293,N_45170,N_44513);
nand U47294 (N_47294,N_44759,N_45319);
xor U47295 (N_47295,N_45632,N_44095);
nand U47296 (N_47296,N_44928,N_44603);
and U47297 (N_47297,N_45918,N_45781);
and U47298 (N_47298,N_45600,N_45094);
or U47299 (N_47299,N_45560,N_45476);
nand U47300 (N_47300,N_44001,N_45311);
and U47301 (N_47301,N_44403,N_44582);
nand U47302 (N_47302,N_44211,N_45430);
nor U47303 (N_47303,N_44770,N_45905);
and U47304 (N_47304,N_45713,N_45898);
xnor U47305 (N_47305,N_44573,N_45286);
or U47306 (N_47306,N_44006,N_45485);
nand U47307 (N_47307,N_44792,N_44697);
and U47308 (N_47308,N_44729,N_45010);
and U47309 (N_47309,N_44356,N_45313);
nor U47310 (N_47310,N_44713,N_45326);
nand U47311 (N_47311,N_45463,N_44374);
nor U47312 (N_47312,N_45688,N_45159);
nor U47313 (N_47313,N_44549,N_44836);
or U47314 (N_47314,N_44670,N_44782);
and U47315 (N_47315,N_44246,N_44602);
and U47316 (N_47316,N_44098,N_44500);
xor U47317 (N_47317,N_44664,N_45744);
nand U47318 (N_47318,N_44066,N_44997);
or U47319 (N_47319,N_44616,N_45197);
nor U47320 (N_47320,N_44656,N_44470);
nor U47321 (N_47321,N_45534,N_45607);
or U47322 (N_47322,N_44916,N_45140);
or U47323 (N_47323,N_44291,N_44330);
or U47324 (N_47324,N_44772,N_45626);
or U47325 (N_47325,N_45001,N_44261);
or U47326 (N_47326,N_45489,N_45474);
nand U47327 (N_47327,N_45203,N_44105);
or U47328 (N_47328,N_45333,N_44846);
nand U47329 (N_47329,N_44078,N_45645);
nand U47330 (N_47330,N_45510,N_44013);
and U47331 (N_47331,N_44905,N_44064);
xor U47332 (N_47332,N_44990,N_44282);
and U47333 (N_47333,N_45993,N_44432);
and U47334 (N_47334,N_45233,N_44206);
and U47335 (N_47335,N_45125,N_44471);
xor U47336 (N_47336,N_45483,N_44615);
xnor U47337 (N_47337,N_45783,N_45868);
nor U47338 (N_47338,N_45105,N_45930);
nand U47339 (N_47339,N_45521,N_45124);
nand U47340 (N_47340,N_44934,N_44987);
xor U47341 (N_47341,N_45295,N_44904);
or U47342 (N_47342,N_44829,N_45095);
nor U47343 (N_47343,N_45845,N_44317);
nor U47344 (N_47344,N_44639,N_44698);
or U47345 (N_47345,N_45424,N_45191);
nor U47346 (N_47346,N_45049,N_44876);
or U47347 (N_47347,N_44348,N_44617);
xnor U47348 (N_47348,N_45551,N_44821);
or U47349 (N_47349,N_45781,N_44608);
or U47350 (N_47350,N_44756,N_45408);
nand U47351 (N_47351,N_44400,N_45918);
xor U47352 (N_47352,N_44809,N_44022);
or U47353 (N_47353,N_44555,N_44307);
or U47354 (N_47354,N_44499,N_44819);
nand U47355 (N_47355,N_44184,N_45016);
nor U47356 (N_47356,N_44853,N_45785);
nor U47357 (N_47357,N_44345,N_44096);
xnor U47358 (N_47358,N_44633,N_44531);
nand U47359 (N_47359,N_45041,N_44877);
and U47360 (N_47360,N_44311,N_45370);
or U47361 (N_47361,N_44120,N_44104);
nand U47362 (N_47362,N_44834,N_45841);
or U47363 (N_47363,N_45115,N_45612);
and U47364 (N_47364,N_45258,N_45941);
xor U47365 (N_47365,N_44454,N_45894);
nor U47366 (N_47366,N_44703,N_45873);
nand U47367 (N_47367,N_44874,N_44527);
xnor U47368 (N_47368,N_45287,N_44419);
nor U47369 (N_47369,N_45118,N_44681);
or U47370 (N_47370,N_44614,N_44341);
nor U47371 (N_47371,N_44795,N_44696);
xor U47372 (N_47372,N_45225,N_45776);
nand U47373 (N_47373,N_45437,N_44499);
or U47374 (N_47374,N_45250,N_45197);
xor U47375 (N_47375,N_45547,N_44905);
xor U47376 (N_47376,N_44527,N_44478);
xor U47377 (N_47377,N_45504,N_45361);
or U47378 (N_47378,N_44474,N_44786);
nand U47379 (N_47379,N_45533,N_45196);
nor U47380 (N_47380,N_44616,N_45340);
nand U47381 (N_47381,N_45470,N_45795);
nand U47382 (N_47382,N_44820,N_44694);
and U47383 (N_47383,N_45003,N_45921);
xnor U47384 (N_47384,N_44312,N_45330);
nand U47385 (N_47385,N_45477,N_44184);
or U47386 (N_47386,N_44765,N_45606);
and U47387 (N_47387,N_45800,N_45319);
xor U47388 (N_47388,N_45509,N_45294);
or U47389 (N_47389,N_44551,N_45974);
or U47390 (N_47390,N_44957,N_44655);
nand U47391 (N_47391,N_45862,N_45866);
or U47392 (N_47392,N_44632,N_44497);
nor U47393 (N_47393,N_44843,N_44041);
or U47394 (N_47394,N_45781,N_44332);
nor U47395 (N_47395,N_45418,N_44304);
xor U47396 (N_47396,N_44408,N_44178);
nand U47397 (N_47397,N_45750,N_44034);
or U47398 (N_47398,N_45126,N_45391);
nor U47399 (N_47399,N_44547,N_44514);
or U47400 (N_47400,N_44175,N_45354);
and U47401 (N_47401,N_44885,N_44906);
or U47402 (N_47402,N_44143,N_45769);
nand U47403 (N_47403,N_44908,N_44957);
xor U47404 (N_47404,N_45529,N_45132);
xor U47405 (N_47405,N_44325,N_44259);
xor U47406 (N_47406,N_44918,N_45524);
or U47407 (N_47407,N_44823,N_44278);
xor U47408 (N_47408,N_44337,N_44715);
xor U47409 (N_47409,N_44348,N_45987);
nand U47410 (N_47410,N_44816,N_45956);
xor U47411 (N_47411,N_44117,N_44913);
xor U47412 (N_47412,N_45501,N_45883);
nor U47413 (N_47413,N_44742,N_44243);
and U47414 (N_47414,N_44964,N_45026);
xnor U47415 (N_47415,N_44005,N_44452);
or U47416 (N_47416,N_45272,N_44599);
xnor U47417 (N_47417,N_44958,N_44256);
xor U47418 (N_47418,N_45090,N_44943);
nor U47419 (N_47419,N_44010,N_44970);
or U47420 (N_47420,N_44281,N_45071);
xor U47421 (N_47421,N_45737,N_44866);
or U47422 (N_47422,N_44710,N_45090);
nor U47423 (N_47423,N_45798,N_44688);
xor U47424 (N_47424,N_44861,N_44169);
nand U47425 (N_47425,N_45895,N_44862);
and U47426 (N_47426,N_44001,N_45467);
nor U47427 (N_47427,N_45044,N_45082);
nand U47428 (N_47428,N_44565,N_44722);
xor U47429 (N_47429,N_44058,N_44203);
nor U47430 (N_47430,N_45331,N_45581);
or U47431 (N_47431,N_45045,N_44138);
xor U47432 (N_47432,N_44490,N_45166);
nor U47433 (N_47433,N_44252,N_45772);
nand U47434 (N_47434,N_45484,N_44724);
or U47435 (N_47435,N_45453,N_45480);
or U47436 (N_47436,N_45028,N_44775);
xnor U47437 (N_47437,N_45878,N_45356);
and U47438 (N_47438,N_44991,N_45735);
nor U47439 (N_47439,N_44263,N_45131);
xor U47440 (N_47440,N_45070,N_44950);
nor U47441 (N_47441,N_44949,N_44592);
xnor U47442 (N_47442,N_45629,N_44783);
or U47443 (N_47443,N_44703,N_45614);
nor U47444 (N_47444,N_45751,N_45124);
nand U47445 (N_47445,N_44098,N_44709);
nor U47446 (N_47446,N_44935,N_44820);
xor U47447 (N_47447,N_44719,N_45663);
xor U47448 (N_47448,N_44424,N_45492);
and U47449 (N_47449,N_44101,N_44816);
xnor U47450 (N_47450,N_45314,N_44495);
nor U47451 (N_47451,N_44398,N_45746);
and U47452 (N_47452,N_45291,N_44560);
and U47453 (N_47453,N_45254,N_45632);
and U47454 (N_47454,N_45867,N_45178);
xor U47455 (N_47455,N_45311,N_45615);
nor U47456 (N_47456,N_45713,N_45029);
and U47457 (N_47457,N_44089,N_44792);
nor U47458 (N_47458,N_45420,N_45205);
and U47459 (N_47459,N_45225,N_45399);
nor U47460 (N_47460,N_45469,N_45047);
and U47461 (N_47461,N_45789,N_44564);
and U47462 (N_47462,N_45346,N_44573);
xnor U47463 (N_47463,N_45397,N_44383);
nor U47464 (N_47464,N_45635,N_45808);
nor U47465 (N_47465,N_44125,N_44313);
and U47466 (N_47466,N_45545,N_44336);
and U47467 (N_47467,N_44555,N_45845);
xor U47468 (N_47468,N_45609,N_44271);
or U47469 (N_47469,N_44299,N_45963);
nor U47470 (N_47470,N_44580,N_44165);
nor U47471 (N_47471,N_44625,N_45517);
nor U47472 (N_47472,N_44924,N_44687);
and U47473 (N_47473,N_44158,N_44390);
nor U47474 (N_47474,N_45942,N_44485);
and U47475 (N_47475,N_45548,N_44995);
or U47476 (N_47476,N_45341,N_44863);
or U47477 (N_47477,N_44580,N_45804);
nor U47478 (N_47478,N_44487,N_44199);
and U47479 (N_47479,N_45605,N_44447);
or U47480 (N_47480,N_44763,N_45598);
nor U47481 (N_47481,N_45395,N_44048);
and U47482 (N_47482,N_45754,N_45023);
nor U47483 (N_47483,N_44963,N_45139);
xnor U47484 (N_47484,N_44117,N_44657);
or U47485 (N_47485,N_45966,N_45209);
xnor U47486 (N_47486,N_44792,N_44199);
nor U47487 (N_47487,N_44234,N_44769);
and U47488 (N_47488,N_45815,N_45420);
and U47489 (N_47489,N_45978,N_45938);
and U47490 (N_47490,N_44373,N_45373);
and U47491 (N_47491,N_45561,N_45514);
nor U47492 (N_47492,N_44809,N_44862);
nand U47493 (N_47493,N_44632,N_45905);
xnor U47494 (N_47494,N_44834,N_45017);
nor U47495 (N_47495,N_44137,N_45738);
nor U47496 (N_47496,N_45788,N_45244);
nor U47497 (N_47497,N_45751,N_44784);
xnor U47498 (N_47498,N_44680,N_44183);
or U47499 (N_47499,N_45570,N_44054);
nor U47500 (N_47500,N_44467,N_44760);
and U47501 (N_47501,N_45351,N_44188);
and U47502 (N_47502,N_45342,N_45964);
nand U47503 (N_47503,N_44180,N_45436);
and U47504 (N_47504,N_44101,N_44014);
and U47505 (N_47505,N_45443,N_44200);
xnor U47506 (N_47506,N_44733,N_44270);
nand U47507 (N_47507,N_45365,N_45931);
or U47508 (N_47508,N_45077,N_45909);
and U47509 (N_47509,N_44373,N_45436);
and U47510 (N_47510,N_45950,N_45833);
nor U47511 (N_47511,N_44659,N_44737);
nor U47512 (N_47512,N_45532,N_45500);
xor U47513 (N_47513,N_45543,N_44355);
and U47514 (N_47514,N_45047,N_44361);
and U47515 (N_47515,N_44260,N_45778);
or U47516 (N_47516,N_44826,N_44917);
nand U47517 (N_47517,N_45427,N_45892);
or U47518 (N_47518,N_45925,N_44146);
xor U47519 (N_47519,N_44787,N_44624);
nand U47520 (N_47520,N_45144,N_45351);
nand U47521 (N_47521,N_45561,N_45377);
nand U47522 (N_47522,N_44112,N_45197);
nand U47523 (N_47523,N_44802,N_45129);
nor U47524 (N_47524,N_45315,N_44983);
or U47525 (N_47525,N_45628,N_44909);
xnor U47526 (N_47526,N_44595,N_44447);
and U47527 (N_47527,N_44661,N_44694);
xor U47528 (N_47528,N_45320,N_45350);
and U47529 (N_47529,N_44909,N_45664);
or U47530 (N_47530,N_44454,N_45868);
nand U47531 (N_47531,N_44382,N_44202);
nand U47532 (N_47532,N_45351,N_44125);
and U47533 (N_47533,N_44193,N_44567);
nor U47534 (N_47534,N_44009,N_44330);
xnor U47535 (N_47535,N_44460,N_44080);
nand U47536 (N_47536,N_44129,N_44101);
nor U47537 (N_47537,N_45199,N_44765);
or U47538 (N_47538,N_45309,N_44060);
nand U47539 (N_47539,N_45586,N_44865);
nand U47540 (N_47540,N_45405,N_44533);
nor U47541 (N_47541,N_45881,N_45855);
nor U47542 (N_47542,N_44251,N_45113);
nand U47543 (N_47543,N_45649,N_44168);
or U47544 (N_47544,N_45150,N_45895);
or U47545 (N_47545,N_44608,N_45898);
or U47546 (N_47546,N_44230,N_44552);
nand U47547 (N_47547,N_45026,N_45537);
or U47548 (N_47548,N_44108,N_45634);
or U47549 (N_47549,N_45120,N_45125);
nor U47550 (N_47550,N_45457,N_45629);
or U47551 (N_47551,N_44341,N_45234);
and U47552 (N_47552,N_45405,N_45449);
xor U47553 (N_47553,N_45175,N_44139);
or U47554 (N_47554,N_44479,N_44599);
xor U47555 (N_47555,N_44995,N_45765);
and U47556 (N_47556,N_45341,N_45964);
nand U47557 (N_47557,N_44830,N_44210);
or U47558 (N_47558,N_44648,N_45449);
xnor U47559 (N_47559,N_45255,N_44066);
xor U47560 (N_47560,N_45915,N_45313);
nor U47561 (N_47561,N_45596,N_45014);
xor U47562 (N_47562,N_44786,N_44624);
xor U47563 (N_47563,N_44782,N_44889);
xnor U47564 (N_47564,N_45358,N_45070);
nand U47565 (N_47565,N_45997,N_45046);
xnor U47566 (N_47566,N_44277,N_44841);
nor U47567 (N_47567,N_44828,N_45801);
nand U47568 (N_47568,N_44109,N_44712);
or U47569 (N_47569,N_45424,N_44889);
nor U47570 (N_47570,N_45646,N_44611);
and U47571 (N_47571,N_44907,N_44309);
or U47572 (N_47572,N_44014,N_45116);
nand U47573 (N_47573,N_45213,N_45631);
nor U47574 (N_47574,N_45827,N_44121);
xor U47575 (N_47575,N_45437,N_44228);
and U47576 (N_47576,N_45133,N_45306);
nand U47577 (N_47577,N_45384,N_44132);
nor U47578 (N_47578,N_45913,N_45246);
and U47579 (N_47579,N_44997,N_45738);
xnor U47580 (N_47580,N_45773,N_44953);
or U47581 (N_47581,N_44964,N_45194);
nand U47582 (N_47582,N_45274,N_44873);
nand U47583 (N_47583,N_44206,N_45592);
nand U47584 (N_47584,N_44934,N_44678);
xor U47585 (N_47585,N_45389,N_44987);
nand U47586 (N_47586,N_45201,N_45579);
xnor U47587 (N_47587,N_45402,N_45314);
xor U47588 (N_47588,N_44877,N_44879);
nand U47589 (N_47589,N_45237,N_44247);
xor U47590 (N_47590,N_44808,N_44508);
xor U47591 (N_47591,N_45557,N_44052);
and U47592 (N_47592,N_44307,N_44584);
and U47593 (N_47593,N_44945,N_44064);
nand U47594 (N_47594,N_44107,N_44260);
nor U47595 (N_47595,N_44592,N_44511);
or U47596 (N_47596,N_45563,N_44212);
nand U47597 (N_47597,N_44260,N_44676);
nand U47598 (N_47598,N_44070,N_45573);
nor U47599 (N_47599,N_44463,N_45264);
nor U47600 (N_47600,N_45246,N_44898);
and U47601 (N_47601,N_45544,N_45280);
nand U47602 (N_47602,N_45343,N_44929);
and U47603 (N_47603,N_44884,N_44750);
nand U47604 (N_47604,N_44346,N_45294);
and U47605 (N_47605,N_45903,N_44072);
nor U47606 (N_47606,N_44664,N_44354);
nand U47607 (N_47607,N_44601,N_45452);
xnor U47608 (N_47608,N_44792,N_45730);
nand U47609 (N_47609,N_44076,N_44436);
and U47610 (N_47610,N_44206,N_45100);
xor U47611 (N_47611,N_44359,N_44829);
xor U47612 (N_47612,N_45644,N_44516);
nand U47613 (N_47613,N_45383,N_44058);
nand U47614 (N_47614,N_44259,N_45285);
and U47615 (N_47615,N_44157,N_44866);
xor U47616 (N_47616,N_44555,N_45138);
nand U47617 (N_47617,N_44891,N_44527);
nand U47618 (N_47618,N_44103,N_45912);
xnor U47619 (N_47619,N_45622,N_44631);
nor U47620 (N_47620,N_44831,N_45349);
and U47621 (N_47621,N_45203,N_44059);
and U47622 (N_47622,N_44203,N_45891);
nor U47623 (N_47623,N_44552,N_44953);
xor U47624 (N_47624,N_44245,N_45254);
nand U47625 (N_47625,N_44615,N_44760);
nand U47626 (N_47626,N_45079,N_45204);
nand U47627 (N_47627,N_45694,N_44110);
xnor U47628 (N_47628,N_45575,N_44919);
or U47629 (N_47629,N_45746,N_45196);
nand U47630 (N_47630,N_44328,N_44620);
xnor U47631 (N_47631,N_45669,N_45097);
nor U47632 (N_47632,N_44866,N_44102);
nor U47633 (N_47633,N_45980,N_45214);
nor U47634 (N_47634,N_44903,N_44448);
xor U47635 (N_47635,N_44578,N_45719);
nor U47636 (N_47636,N_44069,N_44913);
xor U47637 (N_47637,N_44339,N_44255);
and U47638 (N_47638,N_45837,N_44341);
or U47639 (N_47639,N_45531,N_45509);
nand U47640 (N_47640,N_44300,N_44796);
xor U47641 (N_47641,N_44318,N_45659);
and U47642 (N_47642,N_44637,N_44011);
or U47643 (N_47643,N_45576,N_45302);
or U47644 (N_47644,N_44722,N_44748);
nand U47645 (N_47645,N_45565,N_44275);
nor U47646 (N_47646,N_45098,N_45143);
nor U47647 (N_47647,N_45084,N_45339);
and U47648 (N_47648,N_44796,N_45601);
or U47649 (N_47649,N_45540,N_44786);
nor U47650 (N_47650,N_45846,N_44788);
nor U47651 (N_47651,N_45033,N_44530);
and U47652 (N_47652,N_44654,N_45938);
nor U47653 (N_47653,N_44059,N_44736);
and U47654 (N_47654,N_45698,N_45904);
xnor U47655 (N_47655,N_45460,N_45297);
or U47656 (N_47656,N_44563,N_45719);
nor U47657 (N_47657,N_45915,N_45922);
and U47658 (N_47658,N_44410,N_45939);
and U47659 (N_47659,N_44079,N_45104);
nor U47660 (N_47660,N_45690,N_44831);
xnor U47661 (N_47661,N_44996,N_44334);
nor U47662 (N_47662,N_44656,N_45681);
and U47663 (N_47663,N_45579,N_44468);
or U47664 (N_47664,N_44592,N_45536);
nor U47665 (N_47665,N_44538,N_45430);
xor U47666 (N_47666,N_45378,N_44026);
nand U47667 (N_47667,N_45892,N_45088);
and U47668 (N_47668,N_45585,N_45431);
or U47669 (N_47669,N_45498,N_44131);
or U47670 (N_47670,N_44494,N_45422);
or U47671 (N_47671,N_44470,N_44752);
and U47672 (N_47672,N_44192,N_44218);
and U47673 (N_47673,N_45956,N_45077);
or U47674 (N_47674,N_44842,N_44604);
or U47675 (N_47675,N_45487,N_45874);
xor U47676 (N_47676,N_44296,N_45528);
xnor U47677 (N_47677,N_44484,N_44137);
nand U47678 (N_47678,N_44506,N_45603);
xor U47679 (N_47679,N_44141,N_45186);
nand U47680 (N_47680,N_45908,N_44051);
nand U47681 (N_47681,N_44730,N_45412);
xor U47682 (N_47682,N_45727,N_45060);
xor U47683 (N_47683,N_45847,N_45026);
xor U47684 (N_47684,N_44849,N_44133);
or U47685 (N_47685,N_44350,N_44468);
xor U47686 (N_47686,N_44217,N_45530);
or U47687 (N_47687,N_45400,N_44459);
nor U47688 (N_47688,N_44091,N_45359);
nand U47689 (N_47689,N_45415,N_44484);
and U47690 (N_47690,N_44527,N_44313);
nand U47691 (N_47691,N_45253,N_44481);
and U47692 (N_47692,N_44993,N_44489);
or U47693 (N_47693,N_45089,N_45515);
nor U47694 (N_47694,N_45653,N_45756);
nor U47695 (N_47695,N_45595,N_45621);
or U47696 (N_47696,N_45592,N_45797);
xnor U47697 (N_47697,N_45892,N_45734);
and U47698 (N_47698,N_44364,N_44060);
or U47699 (N_47699,N_45451,N_44385);
xor U47700 (N_47700,N_44313,N_44598);
and U47701 (N_47701,N_44679,N_44462);
xor U47702 (N_47702,N_45053,N_44748);
xor U47703 (N_47703,N_44830,N_45287);
and U47704 (N_47704,N_44502,N_45307);
nand U47705 (N_47705,N_45588,N_44064);
or U47706 (N_47706,N_44455,N_45152);
and U47707 (N_47707,N_44871,N_45676);
xor U47708 (N_47708,N_44610,N_44828);
and U47709 (N_47709,N_44953,N_45576);
and U47710 (N_47710,N_44000,N_45792);
or U47711 (N_47711,N_44978,N_45421);
and U47712 (N_47712,N_45273,N_45247);
nand U47713 (N_47713,N_44331,N_45185);
nand U47714 (N_47714,N_45650,N_44849);
nor U47715 (N_47715,N_44796,N_44096);
nand U47716 (N_47716,N_45482,N_44383);
or U47717 (N_47717,N_44502,N_45194);
nand U47718 (N_47718,N_45773,N_44232);
or U47719 (N_47719,N_45152,N_45362);
or U47720 (N_47720,N_44964,N_44609);
nor U47721 (N_47721,N_45650,N_44696);
nor U47722 (N_47722,N_44138,N_45758);
or U47723 (N_47723,N_45327,N_44692);
nand U47724 (N_47724,N_44522,N_45406);
or U47725 (N_47725,N_45087,N_45966);
nor U47726 (N_47726,N_45664,N_45670);
and U47727 (N_47727,N_45564,N_45964);
xnor U47728 (N_47728,N_44517,N_44955);
nor U47729 (N_47729,N_44064,N_45097);
nor U47730 (N_47730,N_44168,N_44617);
xor U47731 (N_47731,N_45403,N_45524);
nor U47732 (N_47732,N_44642,N_45959);
nand U47733 (N_47733,N_44301,N_45003);
nor U47734 (N_47734,N_44784,N_44850);
and U47735 (N_47735,N_44543,N_44821);
nor U47736 (N_47736,N_44371,N_44011);
nand U47737 (N_47737,N_44656,N_45854);
or U47738 (N_47738,N_44262,N_45195);
or U47739 (N_47739,N_44405,N_44317);
nand U47740 (N_47740,N_45227,N_45313);
nand U47741 (N_47741,N_45968,N_44779);
nand U47742 (N_47742,N_45754,N_45316);
and U47743 (N_47743,N_45096,N_45596);
nand U47744 (N_47744,N_44032,N_44219);
or U47745 (N_47745,N_45000,N_44979);
xnor U47746 (N_47746,N_44235,N_45975);
nand U47747 (N_47747,N_45017,N_45762);
xnor U47748 (N_47748,N_45285,N_45785);
or U47749 (N_47749,N_44417,N_45383);
and U47750 (N_47750,N_45641,N_45079);
nand U47751 (N_47751,N_45261,N_44887);
nand U47752 (N_47752,N_44158,N_45176);
or U47753 (N_47753,N_45379,N_45671);
nor U47754 (N_47754,N_45412,N_45182);
nor U47755 (N_47755,N_44204,N_45810);
and U47756 (N_47756,N_45470,N_44159);
nand U47757 (N_47757,N_44500,N_45805);
xnor U47758 (N_47758,N_45686,N_45510);
xnor U47759 (N_47759,N_44046,N_45536);
nor U47760 (N_47760,N_44595,N_44713);
nand U47761 (N_47761,N_44877,N_44322);
and U47762 (N_47762,N_44012,N_45549);
nor U47763 (N_47763,N_44479,N_44023);
nand U47764 (N_47764,N_44811,N_44855);
nand U47765 (N_47765,N_45275,N_45708);
xor U47766 (N_47766,N_44518,N_45512);
nand U47767 (N_47767,N_44399,N_45708);
or U47768 (N_47768,N_44778,N_45415);
or U47769 (N_47769,N_44693,N_45115);
nand U47770 (N_47770,N_45856,N_45186);
and U47771 (N_47771,N_45851,N_45856);
nand U47772 (N_47772,N_45317,N_45498);
or U47773 (N_47773,N_44299,N_45649);
xor U47774 (N_47774,N_44049,N_44218);
nor U47775 (N_47775,N_45575,N_45309);
or U47776 (N_47776,N_45067,N_44435);
and U47777 (N_47777,N_44434,N_45533);
xnor U47778 (N_47778,N_45308,N_45632);
and U47779 (N_47779,N_45150,N_45606);
nand U47780 (N_47780,N_44920,N_45985);
and U47781 (N_47781,N_45701,N_44856);
xor U47782 (N_47782,N_45553,N_45473);
xnor U47783 (N_47783,N_45741,N_44969);
nor U47784 (N_47784,N_44810,N_45862);
nor U47785 (N_47785,N_44017,N_44655);
and U47786 (N_47786,N_45332,N_44266);
or U47787 (N_47787,N_45863,N_44340);
nand U47788 (N_47788,N_45826,N_45174);
and U47789 (N_47789,N_44140,N_44960);
or U47790 (N_47790,N_44392,N_44721);
xor U47791 (N_47791,N_45255,N_44141);
or U47792 (N_47792,N_44193,N_44993);
and U47793 (N_47793,N_44121,N_45680);
or U47794 (N_47794,N_44487,N_45126);
xnor U47795 (N_47795,N_44796,N_44831);
or U47796 (N_47796,N_44633,N_45781);
nor U47797 (N_47797,N_45908,N_44023);
nor U47798 (N_47798,N_44545,N_44929);
nand U47799 (N_47799,N_44656,N_44175);
xnor U47800 (N_47800,N_45222,N_45751);
nor U47801 (N_47801,N_45411,N_44037);
xnor U47802 (N_47802,N_44859,N_44371);
nor U47803 (N_47803,N_44220,N_45312);
xnor U47804 (N_47804,N_45471,N_44699);
or U47805 (N_47805,N_45848,N_45628);
xnor U47806 (N_47806,N_45512,N_44792);
and U47807 (N_47807,N_45802,N_44510);
or U47808 (N_47808,N_44183,N_45671);
and U47809 (N_47809,N_44899,N_44032);
nor U47810 (N_47810,N_45601,N_45732);
nand U47811 (N_47811,N_45290,N_44754);
nor U47812 (N_47812,N_45128,N_45207);
xor U47813 (N_47813,N_44567,N_44376);
xor U47814 (N_47814,N_44126,N_45848);
and U47815 (N_47815,N_44226,N_45104);
nor U47816 (N_47816,N_44376,N_44659);
or U47817 (N_47817,N_45050,N_44814);
xor U47818 (N_47818,N_45174,N_44673);
nand U47819 (N_47819,N_44264,N_45396);
and U47820 (N_47820,N_44324,N_45078);
nor U47821 (N_47821,N_45056,N_44849);
nand U47822 (N_47822,N_44039,N_45043);
or U47823 (N_47823,N_45987,N_44749);
nand U47824 (N_47824,N_44197,N_45581);
nand U47825 (N_47825,N_44653,N_44217);
or U47826 (N_47826,N_44705,N_45318);
nand U47827 (N_47827,N_45787,N_45049);
nor U47828 (N_47828,N_45636,N_44391);
nor U47829 (N_47829,N_44894,N_45586);
nor U47830 (N_47830,N_45810,N_44977);
xor U47831 (N_47831,N_45353,N_45541);
xnor U47832 (N_47832,N_44435,N_44319);
nand U47833 (N_47833,N_44829,N_44616);
or U47834 (N_47834,N_44033,N_45008);
or U47835 (N_47835,N_44411,N_45382);
or U47836 (N_47836,N_44390,N_44219);
nor U47837 (N_47837,N_44614,N_45347);
nand U47838 (N_47838,N_44622,N_44049);
nor U47839 (N_47839,N_45223,N_45252);
and U47840 (N_47840,N_44668,N_44455);
nor U47841 (N_47841,N_45770,N_44727);
xor U47842 (N_47842,N_45565,N_45839);
nand U47843 (N_47843,N_44350,N_44830);
xor U47844 (N_47844,N_45863,N_44147);
or U47845 (N_47845,N_45739,N_44708);
or U47846 (N_47846,N_44683,N_44834);
xnor U47847 (N_47847,N_44813,N_44001);
or U47848 (N_47848,N_44017,N_45540);
nand U47849 (N_47849,N_45887,N_45520);
and U47850 (N_47850,N_44229,N_45020);
xor U47851 (N_47851,N_45531,N_45561);
nand U47852 (N_47852,N_45576,N_45930);
nor U47853 (N_47853,N_45625,N_45522);
nand U47854 (N_47854,N_44960,N_45494);
and U47855 (N_47855,N_45137,N_44656);
and U47856 (N_47856,N_44769,N_45818);
or U47857 (N_47857,N_44954,N_45492);
xor U47858 (N_47858,N_45699,N_44147);
and U47859 (N_47859,N_45506,N_44970);
xor U47860 (N_47860,N_45570,N_45807);
or U47861 (N_47861,N_45578,N_44414);
nor U47862 (N_47862,N_44896,N_45689);
xor U47863 (N_47863,N_44413,N_45060);
nor U47864 (N_47864,N_45237,N_44390);
or U47865 (N_47865,N_45816,N_44567);
xor U47866 (N_47866,N_45224,N_44614);
xnor U47867 (N_47867,N_45418,N_45692);
xor U47868 (N_47868,N_45740,N_45985);
xnor U47869 (N_47869,N_45858,N_44899);
nand U47870 (N_47870,N_44237,N_45967);
xor U47871 (N_47871,N_44137,N_45815);
nand U47872 (N_47872,N_44234,N_45030);
nor U47873 (N_47873,N_44970,N_45834);
and U47874 (N_47874,N_44487,N_44663);
nor U47875 (N_47875,N_45451,N_45570);
and U47876 (N_47876,N_45501,N_44873);
and U47877 (N_47877,N_44724,N_44931);
nor U47878 (N_47878,N_45138,N_44429);
and U47879 (N_47879,N_44583,N_44745);
xnor U47880 (N_47880,N_45642,N_44214);
or U47881 (N_47881,N_45134,N_45097);
nand U47882 (N_47882,N_44689,N_44470);
xnor U47883 (N_47883,N_45858,N_45841);
and U47884 (N_47884,N_45843,N_44333);
nor U47885 (N_47885,N_45480,N_44546);
and U47886 (N_47886,N_45982,N_44110);
nand U47887 (N_47887,N_44685,N_45153);
nand U47888 (N_47888,N_44613,N_45232);
xor U47889 (N_47889,N_44057,N_44454);
and U47890 (N_47890,N_44211,N_44167);
xor U47891 (N_47891,N_45857,N_44822);
nand U47892 (N_47892,N_45038,N_44240);
nand U47893 (N_47893,N_45500,N_45735);
or U47894 (N_47894,N_45465,N_44742);
and U47895 (N_47895,N_45646,N_45840);
nand U47896 (N_47896,N_45355,N_44449);
nor U47897 (N_47897,N_44495,N_44373);
nor U47898 (N_47898,N_44632,N_45229);
and U47899 (N_47899,N_45228,N_44063);
nand U47900 (N_47900,N_44111,N_44831);
nor U47901 (N_47901,N_44639,N_45294);
and U47902 (N_47902,N_45095,N_45288);
nor U47903 (N_47903,N_44041,N_45007);
nand U47904 (N_47904,N_45612,N_44048);
nor U47905 (N_47905,N_45853,N_45838);
nand U47906 (N_47906,N_45264,N_45307);
or U47907 (N_47907,N_44786,N_44439);
xor U47908 (N_47908,N_45281,N_45958);
and U47909 (N_47909,N_44088,N_44490);
nand U47910 (N_47910,N_45224,N_44064);
nor U47911 (N_47911,N_44356,N_45486);
xnor U47912 (N_47912,N_45035,N_45230);
or U47913 (N_47913,N_45349,N_45048);
nand U47914 (N_47914,N_44115,N_45494);
and U47915 (N_47915,N_44912,N_44441);
xnor U47916 (N_47916,N_45374,N_44660);
or U47917 (N_47917,N_45187,N_45941);
nand U47918 (N_47918,N_45959,N_45147);
xor U47919 (N_47919,N_44586,N_45626);
nor U47920 (N_47920,N_45659,N_44648);
nor U47921 (N_47921,N_45092,N_45998);
nor U47922 (N_47922,N_45715,N_44674);
or U47923 (N_47923,N_44065,N_45965);
nand U47924 (N_47924,N_44326,N_44564);
nand U47925 (N_47925,N_44563,N_44259);
xnor U47926 (N_47926,N_44572,N_45087);
nor U47927 (N_47927,N_44948,N_45315);
nand U47928 (N_47928,N_45560,N_44021);
nand U47929 (N_47929,N_44028,N_45325);
nand U47930 (N_47930,N_45797,N_45162);
nand U47931 (N_47931,N_44484,N_44026);
nand U47932 (N_47932,N_45565,N_45043);
nand U47933 (N_47933,N_44055,N_44186);
nand U47934 (N_47934,N_45768,N_45348);
nor U47935 (N_47935,N_45509,N_44324);
xnor U47936 (N_47936,N_45303,N_45648);
or U47937 (N_47937,N_44935,N_44853);
and U47938 (N_47938,N_44936,N_44713);
or U47939 (N_47939,N_44338,N_45788);
and U47940 (N_47940,N_45385,N_44516);
and U47941 (N_47941,N_44279,N_45922);
or U47942 (N_47942,N_45490,N_44881);
nor U47943 (N_47943,N_45898,N_45163);
or U47944 (N_47944,N_45256,N_45827);
and U47945 (N_47945,N_44129,N_44176);
and U47946 (N_47946,N_44105,N_44011);
nand U47947 (N_47947,N_45226,N_45712);
and U47948 (N_47948,N_44107,N_45703);
nor U47949 (N_47949,N_44653,N_45363);
nand U47950 (N_47950,N_45258,N_44558);
and U47951 (N_47951,N_45756,N_45248);
or U47952 (N_47952,N_45032,N_45226);
or U47953 (N_47953,N_45362,N_44459);
or U47954 (N_47954,N_45542,N_44836);
nor U47955 (N_47955,N_45006,N_45333);
nand U47956 (N_47956,N_45344,N_44128);
xnor U47957 (N_47957,N_44396,N_44319);
or U47958 (N_47958,N_44346,N_44018);
xor U47959 (N_47959,N_45285,N_44214);
nand U47960 (N_47960,N_44688,N_44169);
or U47961 (N_47961,N_45322,N_45238);
and U47962 (N_47962,N_45749,N_45478);
or U47963 (N_47963,N_45764,N_45769);
nor U47964 (N_47964,N_44845,N_44025);
or U47965 (N_47965,N_45734,N_45073);
or U47966 (N_47966,N_44597,N_44610);
and U47967 (N_47967,N_44600,N_45364);
or U47968 (N_47968,N_44398,N_44401);
xnor U47969 (N_47969,N_45319,N_45877);
or U47970 (N_47970,N_45952,N_45925);
nor U47971 (N_47971,N_44637,N_44707);
or U47972 (N_47972,N_45053,N_45703);
nand U47973 (N_47973,N_44522,N_45464);
or U47974 (N_47974,N_44143,N_45545);
xnor U47975 (N_47975,N_45280,N_44423);
nand U47976 (N_47976,N_44435,N_44070);
xnor U47977 (N_47977,N_44405,N_45002);
xnor U47978 (N_47978,N_44509,N_44505);
or U47979 (N_47979,N_45703,N_44532);
xor U47980 (N_47980,N_45744,N_44229);
nor U47981 (N_47981,N_44256,N_44251);
xor U47982 (N_47982,N_44915,N_45887);
nand U47983 (N_47983,N_45315,N_45478);
nand U47984 (N_47984,N_45345,N_45632);
and U47985 (N_47985,N_45887,N_45021);
nor U47986 (N_47986,N_45136,N_45023);
and U47987 (N_47987,N_45300,N_45292);
xor U47988 (N_47988,N_44143,N_44536);
nor U47989 (N_47989,N_44099,N_45802);
nor U47990 (N_47990,N_44531,N_44635);
and U47991 (N_47991,N_44724,N_44575);
xor U47992 (N_47992,N_45148,N_44805);
nand U47993 (N_47993,N_45786,N_45538);
or U47994 (N_47994,N_44612,N_44377);
nor U47995 (N_47995,N_44410,N_45563);
nand U47996 (N_47996,N_44451,N_44591);
or U47997 (N_47997,N_44637,N_44153);
nand U47998 (N_47998,N_45269,N_44159);
and U47999 (N_47999,N_44222,N_45120);
nand U48000 (N_48000,N_47626,N_46004);
and U48001 (N_48001,N_46494,N_46829);
or U48002 (N_48002,N_47448,N_47007);
nor U48003 (N_48003,N_46242,N_47386);
or U48004 (N_48004,N_47667,N_46845);
nor U48005 (N_48005,N_47244,N_47812);
xor U48006 (N_48006,N_47500,N_46312);
xnor U48007 (N_48007,N_46558,N_46692);
xnor U48008 (N_48008,N_47375,N_47327);
nand U48009 (N_48009,N_47921,N_47475);
nand U48010 (N_48010,N_46455,N_46405);
xor U48011 (N_48011,N_46086,N_46870);
and U48012 (N_48012,N_46489,N_46419);
nand U48013 (N_48013,N_46787,N_47277);
nand U48014 (N_48014,N_47847,N_47395);
nor U48015 (N_48015,N_46580,N_47035);
and U48016 (N_48016,N_47903,N_46612);
or U48017 (N_48017,N_47433,N_47490);
xnor U48018 (N_48018,N_46183,N_47341);
xnor U48019 (N_48019,N_47225,N_46487);
nand U48020 (N_48020,N_46745,N_46036);
and U48021 (N_48021,N_47021,N_47907);
nand U48022 (N_48022,N_47464,N_47407);
nor U48023 (N_48023,N_46142,N_46576);
and U48024 (N_48024,N_46880,N_46114);
nor U48025 (N_48025,N_46181,N_47821);
xor U48026 (N_48026,N_46951,N_47227);
or U48027 (N_48027,N_46848,N_47278);
nor U48028 (N_48028,N_46407,N_46983);
and U48029 (N_48029,N_47182,N_46621);
nor U48030 (N_48030,N_47250,N_47671);
and U48031 (N_48031,N_47852,N_47460);
nand U48032 (N_48032,N_47934,N_46477);
or U48033 (N_48033,N_46055,N_46457);
or U48034 (N_48034,N_46480,N_47684);
or U48035 (N_48035,N_46384,N_47749);
or U48036 (N_48036,N_47185,N_46875);
and U48037 (N_48037,N_47158,N_47930);
nor U48038 (N_48038,N_47222,N_46273);
xor U48039 (N_48039,N_46145,N_46740);
nand U48040 (N_48040,N_47195,N_47027);
and U48041 (N_48041,N_46902,N_46328);
or U48042 (N_48042,N_47703,N_46015);
nand U48043 (N_48043,N_46435,N_47226);
xnor U48044 (N_48044,N_46675,N_46700);
and U48045 (N_48045,N_46473,N_47177);
xor U48046 (N_48046,N_47493,N_46199);
or U48047 (N_48047,N_47036,N_47335);
nor U48048 (N_48048,N_47659,N_46097);
xor U48049 (N_48049,N_46041,N_46826);
or U48050 (N_48050,N_46536,N_46859);
xnor U48051 (N_48051,N_47442,N_46561);
nand U48052 (N_48052,N_47510,N_47496);
and U48053 (N_48053,N_46193,N_46288);
and U48054 (N_48054,N_46661,N_46044);
xnor U48055 (N_48055,N_47048,N_47108);
nor U48056 (N_48056,N_46757,N_46638);
xor U48057 (N_48057,N_46838,N_47274);
nor U48058 (N_48058,N_47113,N_47658);
or U48059 (N_48059,N_46802,N_46235);
xor U48060 (N_48060,N_46581,N_47162);
nor U48061 (N_48061,N_47075,N_46828);
and U48062 (N_48062,N_47254,N_46831);
nor U48063 (N_48063,N_47874,N_47529);
nor U48064 (N_48064,N_47023,N_46202);
xnor U48065 (N_48065,N_47466,N_46393);
nor U48066 (N_48066,N_47209,N_47573);
nand U48067 (N_48067,N_46942,N_46538);
nor U48068 (N_48068,N_46395,N_47926);
and U48069 (N_48069,N_47008,N_47423);
xor U48070 (N_48070,N_46557,N_46377);
xor U48071 (N_48071,N_47791,N_46468);
and U48072 (N_48072,N_47371,N_46450);
xor U48073 (N_48073,N_46894,N_46436);
nor U48074 (N_48074,N_46132,N_47831);
nand U48075 (N_48075,N_47649,N_46192);
nand U48076 (N_48076,N_46998,N_47757);
xor U48077 (N_48077,N_47869,N_47815);
nor U48078 (N_48078,N_47217,N_46529);
xnor U48079 (N_48079,N_47196,N_46754);
and U48080 (N_48080,N_47987,N_47774);
nor U48081 (N_48081,N_47619,N_47031);
and U48082 (N_48082,N_47688,N_47894);
nor U48083 (N_48083,N_47977,N_46355);
or U48084 (N_48084,N_46185,N_46440);
or U48085 (N_48085,N_46175,N_47288);
nor U48086 (N_48086,N_47727,N_46492);
nand U48087 (N_48087,N_46146,N_47611);
and U48088 (N_48088,N_47692,N_46897);
xor U48089 (N_48089,N_46148,N_47319);
nand U48090 (N_48090,N_46263,N_47854);
nand U48091 (N_48091,N_47176,N_46807);
nand U48092 (N_48092,N_47419,N_47236);
or U48093 (N_48093,N_46043,N_47875);
nor U48094 (N_48094,N_46153,N_46048);
or U48095 (N_48095,N_46216,N_47102);
xor U48096 (N_48096,N_47194,N_46840);
nand U48097 (N_48097,N_47302,N_46766);
or U48098 (N_48098,N_46399,N_46720);
nand U48099 (N_48099,N_46070,N_47439);
xnor U48100 (N_48100,N_47437,N_47775);
nand U48101 (N_48101,N_47893,N_46987);
nor U48102 (N_48102,N_46873,N_47342);
and U48103 (N_48103,N_46630,N_46750);
or U48104 (N_48104,N_46472,N_47586);
nor U48105 (N_48105,N_46311,N_46849);
nor U48106 (N_48106,N_47802,N_47268);
or U48107 (N_48107,N_46844,N_47426);
and U48108 (N_48108,N_47693,N_47050);
and U48109 (N_48109,N_46375,N_47279);
nand U48110 (N_48110,N_47404,N_47032);
nor U48111 (N_48111,N_47382,N_46151);
nand U48112 (N_48112,N_47465,N_47932);
nand U48113 (N_48113,N_46304,N_46843);
nand U48114 (N_48114,N_46247,N_46644);
and U48115 (N_48115,N_47920,N_47340);
nand U48116 (N_48116,N_47537,N_46356);
and U48117 (N_48117,N_46491,N_46636);
or U48118 (N_48118,N_47840,N_47306);
xnor U48119 (N_48119,N_46194,N_46915);
nor U48120 (N_48120,N_47741,N_46308);
and U48121 (N_48121,N_46496,N_46103);
nor U48122 (N_48122,N_47374,N_46508);
xor U48123 (N_48123,N_47047,N_46079);
or U48124 (N_48124,N_46486,N_47512);
and U48125 (N_48125,N_46751,N_46299);
nor U48126 (N_48126,N_46954,N_47785);
and U48127 (N_48127,N_47314,N_47432);
or U48128 (N_48128,N_46591,N_46542);
xor U48129 (N_48129,N_47685,N_47730);
or U48130 (N_48130,N_47579,N_46735);
and U48131 (N_48131,N_46825,N_46137);
nor U48132 (N_48132,N_46085,N_46075);
or U48133 (N_48133,N_47294,N_47083);
nand U48134 (N_48134,N_47914,N_46364);
nor U48135 (N_48135,N_46539,N_46819);
nand U48136 (N_48136,N_46526,N_46546);
nor U48137 (N_48137,N_46686,N_46068);
xor U48138 (N_48138,N_47181,N_46470);
xnor U48139 (N_48139,N_47830,N_46764);
xnor U48140 (N_48140,N_46232,N_47180);
nand U48141 (N_48141,N_47845,N_46238);
and U48142 (N_48142,N_46669,N_46369);
nor U48143 (N_48143,N_47017,N_47892);
and U48144 (N_48144,N_46101,N_46748);
nand U48145 (N_48145,N_47249,N_47208);
xnor U48146 (N_48146,N_46275,N_47644);
and U48147 (N_48147,N_47834,N_47015);
xor U48148 (N_48148,N_46280,N_47801);
xnor U48149 (N_48149,N_46276,N_46615);
xor U48150 (N_48150,N_47729,N_47780);
nand U48151 (N_48151,N_46960,N_47555);
nor U48152 (N_48152,N_46417,N_46303);
nand U48153 (N_48153,N_46903,N_46379);
xor U48154 (N_48154,N_46523,N_47993);
and U48155 (N_48155,N_46882,N_47119);
xnor U48156 (N_48156,N_46483,N_46279);
or U48157 (N_48157,N_47642,N_47811);
nand U48158 (N_48158,N_46810,N_46078);
and U48159 (N_48159,N_47410,N_47469);
nor U48160 (N_48160,N_47515,N_46241);
nor U48161 (N_48161,N_46966,N_46033);
and U48162 (N_48162,N_46712,N_47878);
or U48163 (N_48163,N_47298,N_47485);
nand U48164 (N_48164,N_47711,N_47049);
nor U48165 (N_48165,N_46025,N_47985);
and U48166 (N_48166,N_47309,N_47440);
xnor U48167 (N_48167,N_46429,N_46290);
and U48168 (N_48168,N_47584,N_47558);
xnor U48169 (N_48169,N_46448,N_46909);
and U48170 (N_48170,N_46166,N_47415);
xor U48171 (N_48171,N_47098,N_46603);
and U48172 (N_48172,N_46673,N_46578);
nand U48173 (N_48173,N_46830,N_47848);
and U48174 (N_48174,N_47480,N_47166);
nand U48175 (N_48175,N_46991,N_46406);
nand U48176 (N_48176,N_47043,N_46530);
and U48177 (N_48177,N_47782,N_46818);
xor U48178 (N_48178,N_46045,N_47908);
xor U48179 (N_48179,N_47936,N_46133);
and U48180 (N_48180,N_46098,N_47056);
or U48181 (N_48181,N_46511,N_46518);
nand U48182 (N_48182,N_46214,N_47240);
nor U48183 (N_48183,N_46034,N_47165);
xnor U48184 (N_48184,N_47418,N_47184);
xor U48185 (N_48185,N_46198,N_46234);
and U48186 (N_48186,N_47494,N_46274);
nand U48187 (N_48187,N_46365,N_46560);
nand U48188 (N_48188,N_47428,N_47383);
xor U48189 (N_48189,N_47221,N_47100);
nor U48190 (N_48190,N_46459,N_47479);
or U48191 (N_48191,N_46864,N_46442);
or U48192 (N_48192,N_46527,N_47600);
and U48193 (N_48193,N_47486,N_46126);
nand U48194 (N_48194,N_47518,N_47273);
or U48195 (N_48195,N_47927,N_47458);
nand U48196 (N_48196,N_46236,N_46475);
nand U48197 (N_48197,N_46378,N_47147);
xor U48198 (N_48198,N_46462,N_47389);
nor U48199 (N_48199,N_46599,N_47096);
xnor U48200 (N_48200,N_46458,N_46123);
nand U48201 (N_48201,N_47805,N_46069);
or U48202 (N_48202,N_46352,N_47962);
xnor U48203 (N_48203,N_46794,N_47623);
xnor U48204 (N_48204,N_46167,N_46727);
and U48205 (N_48205,N_46189,N_46503);
nor U48206 (N_48206,N_47149,N_46090);
nor U48207 (N_48207,N_47939,N_47417);
nor U48208 (N_48208,N_46115,N_46382);
and U48209 (N_48209,N_47063,N_46037);
xnor U48210 (N_48210,N_47753,N_46590);
nand U48211 (N_48211,N_47593,N_46792);
nor U48212 (N_48212,N_47354,N_46402);
or U48213 (N_48213,N_47204,N_47723);
and U48214 (N_48214,N_47451,N_46583);
nand U48215 (N_48215,N_46310,N_46593);
and U48216 (N_48216,N_46704,N_47495);
xor U48217 (N_48217,N_46208,N_46143);
xor U48218 (N_48218,N_46451,N_46698);
xor U48219 (N_48219,N_47059,N_46656);
and U48220 (N_48220,N_47813,N_46923);
xor U48221 (N_48221,N_47369,N_46484);
and U48222 (N_48222,N_47797,N_46891);
and U48223 (N_48223,N_47614,N_46959);
and U48224 (N_48224,N_47427,N_47997);
xor U48225 (N_48225,N_46002,N_47164);
and U48226 (N_48226,N_46556,N_46327);
xnor U48227 (N_48227,N_46040,N_46980);
or U48228 (N_48228,N_47715,N_46622);
and U48229 (N_48229,N_47077,N_47540);
nor U48230 (N_48230,N_46774,N_46400);
nor U48231 (N_48231,N_46598,N_46338);
and U48232 (N_48232,N_47257,N_47259);
xnor U48233 (N_48233,N_46376,N_46808);
xor U48234 (N_48234,N_46282,N_47533);
or U48235 (N_48235,N_46067,N_47959);
or U48236 (N_48236,N_47473,N_46705);
nand U48237 (N_48237,N_47393,N_47981);
nor U48238 (N_48238,N_47890,N_47039);
nor U48239 (N_48239,N_46449,N_46482);
nor U48240 (N_48240,N_47139,N_46568);
nor U48241 (N_48241,N_47541,N_47950);
xor U48242 (N_48242,N_47054,N_47795);
xnor U48243 (N_48243,N_47357,N_46551);
nor U48244 (N_48244,N_47942,N_47148);
xor U48245 (N_48245,N_47991,N_47322);
nor U48246 (N_48246,N_46390,N_46767);
nand U48247 (N_48247,N_47312,N_47067);
and U48248 (N_48248,N_46747,N_47258);
nor U48249 (N_48249,N_47636,N_47676);
or U48250 (N_48250,N_46566,N_47436);
nor U48251 (N_48251,N_47514,N_46076);
and U48252 (N_48252,N_46267,N_46413);
nor U48253 (N_48253,N_47001,N_46089);
and U48254 (N_48254,N_47560,N_46373);
nand U48255 (N_48255,N_46962,N_47153);
and U48256 (N_48256,N_46061,N_46485);
and U48257 (N_48257,N_47502,N_46682);
xnor U48258 (N_48258,N_46018,N_46456);
and U48259 (N_48259,N_46052,N_47728);
nor U48260 (N_48260,N_47186,N_47680);
and U48261 (N_48261,N_46722,N_47948);
nor U48262 (N_48262,N_46618,N_47046);
and U48263 (N_48263,N_46269,N_47694);
nand U48264 (N_48264,N_46935,N_47712);
or U48265 (N_48265,N_47755,N_46296);
xnor U48266 (N_48266,N_46982,N_47045);
xor U48267 (N_48267,N_47632,N_47958);
and U48268 (N_48268,N_47669,N_46926);
or U48269 (N_48269,N_46995,N_46380);
xnor U48270 (N_48270,N_47005,N_47951);
nand U48271 (N_48271,N_46865,N_47989);
nor U48272 (N_48272,N_47122,N_46605);
xor U48273 (N_48273,N_46936,N_47899);
or U48274 (N_48274,N_47138,N_47980);
and U48275 (N_48275,N_46889,N_47324);
or U48276 (N_48276,N_47606,N_46180);
nor U48277 (N_48277,N_46761,N_46127);
nor U48278 (N_48278,N_46277,N_46822);
or U48279 (N_48279,N_47197,N_47116);
nor U48280 (N_48280,N_46424,N_46213);
xnor U48281 (N_48281,N_47707,N_46649);
nand U48282 (N_48282,N_47362,N_47722);
xnor U48283 (N_48283,N_47858,N_47356);
nor U48284 (N_48284,N_47234,N_46077);
nor U48285 (N_48285,N_46662,N_46677);
or U48286 (N_48286,N_46878,N_46841);
or U48287 (N_48287,N_46914,N_47999);
xnor U48288 (N_48288,N_46737,N_46988);
or U48289 (N_48289,N_46119,N_46339);
xor U48290 (N_48290,N_46083,N_47935);
nand U48291 (N_48291,N_47863,N_46349);
xnor U48292 (N_48292,N_46266,N_47976);
and U48293 (N_48293,N_47477,N_46651);
nand U48294 (N_48294,N_47866,N_47992);
nor U48295 (N_48295,N_46879,N_46857);
or U48296 (N_48296,N_47781,N_47124);
and U48297 (N_48297,N_47613,N_46949);
xor U48298 (N_48298,N_46620,N_46871);
or U48299 (N_48299,N_46361,N_47912);
and U48300 (N_48300,N_46427,N_47702);
xor U48301 (N_48301,N_46782,N_47873);
and U48302 (N_48302,N_46138,N_47624);
or U48303 (N_48303,N_46798,N_46717);
nor U48304 (N_48304,N_46021,N_46813);
xor U48305 (N_48305,N_47161,N_46803);
or U48306 (N_48306,N_47996,N_46362);
nor U48307 (N_48307,N_47704,N_47542);
and U48308 (N_48308,N_46504,N_46804);
and U48309 (N_48309,N_46801,N_47968);
nand U48310 (N_48310,N_46188,N_46158);
and U48311 (N_48311,N_46421,N_46577);
or U48312 (N_48312,N_46348,N_47776);
and U48313 (N_48313,N_47822,N_47343);
nor U48314 (N_48314,N_47175,N_46139);
xnor U48315 (N_48315,N_46001,N_47476);
or U48316 (N_48316,N_47123,N_47378);
or U48317 (N_48317,N_47708,N_46370);
nor U48318 (N_48318,N_47751,N_46324);
and U48319 (N_48319,N_46159,N_46931);
nand U48320 (N_48320,N_47489,N_47889);
or U48321 (N_48321,N_46051,N_46224);
or U48322 (N_48322,N_46921,N_46701);
and U48323 (N_48323,N_46898,N_46610);
nand U48324 (N_48324,N_46817,N_46855);
nand U48325 (N_48325,N_47762,N_47429);
xor U48326 (N_48326,N_46149,N_47504);
nor U48327 (N_48327,N_46938,N_47548);
and U48328 (N_48328,N_47901,N_47397);
and U48329 (N_48329,N_47638,N_46209);
nor U48330 (N_48330,N_46331,N_46094);
or U48331 (N_48331,N_47870,N_47617);
nand U48332 (N_48332,N_47524,N_47607);
nor U48333 (N_48333,N_46010,N_47768);
nor U48334 (N_48334,N_46031,N_47328);
xor U48335 (N_48335,N_47453,N_46336);
and U48336 (N_48336,N_46625,N_47527);
xor U48337 (N_48337,N_47672,N_46904);
nor U48338 (N_48338,N_47013,N_46107);
or U48339 (N_48339,N_47986,N_46883);
or U48340 (N_48340,N_46659,N_47773);
and U48341 (N_48341,N_47145,N_47655);
and U48342 (N_48342,N_46755,N_46297);
nor U48343 (N_48343,N_46329,N_46706);
or U48344 (N_48344,N_47699,N_46999);
nor U48345 (N_48345,N_47264,N_46555);
and U48346 (N_48346,N_46081,N_46796);
and U48347 (N_48347,N_47169,N_47499);
nand U48348 (N_48348,N_46809,N_47660);
and U48349 (N_48349,N_47062,N_46358);
and U48350 (N_48350,N_47092,N_46746);
and U48351 (N_48351,N_47945,N_46478);
nand U48352 (N_48352,N_47344,N_47424);
nor U48353 (N_48353,N_47943,N_47082);
nand U48354 (N_48354,N_47631,N_46912);
nor U48355 (N_48355,N_46301,N_46154);
nand U48356 (N_48356,N_47871,N_46552);
or U48357 (N_48357,N_46385,N_47550);
nand U48358 (N_48358,N_46685,N_47804);
and U48359 (N_48359,N_47745,N_46467);
or U48360 (N_48360,N_47006,N_47783);
nand U48361 (N_48361,N_46009,N_47070);
xor U48362 (N_48362,N_46286,N_46326);
xor U48363 (N_48363,N_46933,N_46237);
nor U48364 (N_48364,N_46423,N_46690);
or U48365 (N_48365,N_47135,N_47482);
nand U48366 (N_48366,N_47587,N_47849);
nor U48367 (N_48367,N_46658,N_47117);
nand U48368 (N_48368,N_47615,N_47364);
or U48369 (N_48369,N_47744,N_46587);
xor U48370 (N_48370,N_46490,N_47020);
nand U48371 (N_48371,N_46000,N_46093);
nor U48372 (N_48372,N_47242,N_47207);
xnor U48373 (N_48373,N_46753,N_47025);
nor U48374 (N_48374,N_47026,N_47630);
nor U48375 (N_48375,N_47561,N_46291);
or U48376 (N_48376,N_47060,N_47530);
nor U48377 (N_48377,N_46643,N_47305);
nor U48378 (N_48378,N_46760,N_47311);
nor U48379 (N_48379,N_46631,N_46298);
nand U48380 (N_48380,N_47718,N_47091);
nor U48381 (N_48381,N_47832,N_46606);
and U48382 (N_48382,N_47851,N_46847);
or U48383 (N_48383,N_46919,N_47756);
xnor U48384 (N_48384,N_47545,N_46640);
and U48385 (N_48385,N_47933,N_47174);
or U48386 (N_48386,N_47329,N_46799);
and U48387 (N_48387,N_47069,N_46901);
nor U48388 (N_48388,N_46863,N_46688);
or U48389 (N_48389,N_47403,N_47752);
xor U48390 (N_48390,N_46836,N_46162);
or U48391 (N_48391,N_46200,N_47150);
xnor U48392 (N_48392,N_46833,N_46674);
xnor U48393 (N_48393,N_47009,N_47778);
nor U48394 (N_48394,N_46397,N_47839);
or U48395 (N_48395,N_47041,N_46695);
xor U48396 (N_48396,N_47183,N_47095);
xor U48397 (N_48397,N_46113,N_46318);
xnor U48398 (N_48398,N_47235,N_46082);
or U48399 (N_48399,N_47733,N_46354);
nor U48400 (N_48400,N_47301,N_47097);
or U48401 (N_48401,N_47154,N_46899);
nand U48402 (N_48402,N_47736,N_47074);
and U48403 (N_48403,N_46289,N_46763);
nand U48404 (N_48404,N_47777,N_47982);
xnor U48405 (N_48405,N_47897,N_46634);
nor U48406 (N_48406,N_46479,N_47764);
or U48407 (N_48407,N_46135,N_47080);
and U48408 (N_48408,N_46363,N_47528);
xor U48409 (N_48409,N_46515,N_46295);
and U48410 (N_48410,N_47238,N_46602);
nand U48411 (N_48411,N_47979,N_46812);
and U48412 (N_48412,N_46736,N_47970);
nand U48413 (N_48413,N_46854,N_47066);
nor U48414 (N_48414,N_47902,N_46258);
or U48415 (N_48415,N_46220,N_47260);
nand U48416 (N_48416,N_47585,N_46768);
or U48417 (N_48417,N_47336,N_47519);
xnor U48418 (N_48418,N_46514,N_46657);
xnor U48419 (N_48419,N_47697,N_46869);
nand U48420 (N_48420,N_46038,N_47739);
and U48421 (N_48421,N_47525,N_46582);
nor U48422 (N_48422,N_46956,N_47019);
nand U48423 (N_48423,N_46409,N_46707);
or U48424 (N_48424,N_46654,N_46171);
and U48425 (N_48425,N_46244,N_46928);
and U48426 (N_48426,N_47334,N_47106);
and U48427 (N_48427,N_47665,N_46832);
nor U48428 (N_48428,N_47915,N_46383);
xor U48429 (N_48429,N_46471,N_46493);
and U48430 (N_48430,N_46716,N_47438);
nand U48431 (N_48431,N_46565,N_46474);
nor U48432 (N_48432,N_47916,N_46650);
or U48433 (N_48433,N_46549,N_47705);
and U48434 (N_48434,N_47232,N_47131);
xnor U48435 (N_48435,N_46262,N_47881);
and U48436 (N_48436,N_46431,N_47798);
nand U48437 (N_48437,N_46510,N_46203);
and U48438 (N_48438,N_47720,N_47352);
xnor U48439 (N_48439,N_46520,N_47443);
xor U48440 (N_48440,N_46343,N_47478);
nand U48441 (N_48441,N_46432,N_46965);
and U48442 (N_48442,N_47919,N_46014);
nand U48443 (N_48443,N_47168,N_46206);
or U48444 (N_48444,N_46368,N_47929);
xor U48445 (N_48445,N_47570,N_46059);
nand U48446 (N_48446,N_47366,N_47957);
xor U48447 (N_48447,N_46795,N_46885);
nand U48448 (N_48448,N_47964,N_47230);
nor U48449 (N_48449,N_46333,N_46758);
and U48450 (N_48450,N_46911,N_47900);
nor U48451 (N_48451,N_47099,N_47474);
xnor U48452 (N_48452,N_47323,N_47520);
nand U48453 (N_48453,N_47747,N_47596);
xor U48454 (N_48454,N_47963,N_46042);
and U48455 (N_48455,N_47351,N_47212);
nor U48456 (N_48456,N_47549,N_46533);
nand U48457 (N_48457,N_46439,N_47506);
xor U48458 (N_48458,N_47406,N_47171);
nor U48459 (N_48459,N_47205,N_46786);
nand U48460 (N_48460,N_46752,N_47178);
and U48461 (N_48461,N_47492,N_46430);
or U48462 (N_48462,N_46228,N_46574);
nor U48463 (N_48463,N_46117,N_47841);
nor U48464 (N_48464,N_47370,N_47193);
nor U48465 (N_48465,N_47882,N_47826);
and U48466 (N_48466,N_46416,N_46080);
nand U48467 (N_48467,N_46667,N_46924);
nor U48468 (N_48468,N_47621,N_47405);
or U48469 (N_48469,N_46394,N_46195);
nand U48470 (N_48470,N_47190,N_47983);
or U48471 (N_48471,N_46645,N_46152);
nor U48472 (N_48472,N_46866,N_46253);
nand U48473 (N_48473,N_47136,N_46895);
nor U48474 (N_48474,N_46488,N_46218);
nand U48475 (N_48475,N_47159,N_46762);
and U48476 (N_48476,N_47719,N_47656);
xnor U48477 (N_48477,N_47975,N_46283);
xnor U48478 (N_48478,N_46734,N_46943);
xnor U48479 (N_48479,N_46941,N_47944);
nand U48480 (N_48480,N_46334,N_47239);
and U48481 (N_48481,N_47865,N_46102);
xor U48482 (N_48482,N_47125,N_47673);
and U48483 (N_48483,N_46392,N_46547);
and U48484 (N_48484,N_46824,N_46302);
or U48485 (N_48485,N_46011,N_46250);
and U48486 (N_48486,N_47079,N_46481);
and U48487 (N_48487,N_47118,N_46872);
and U48488 (N_48488,N_46939,N_47716);
or U48489 (N_48489,N_47856,N_46927);
or U48490 (N_48490,N_46120,N_46222);
and U48491 (N_48491,N_46210,N_46594);
nor U48492 (N_48492,N_47895,N_47661);
and U48493 (N_48493,N_46715,N_46505);
nor U48494 (N_48494,N_47201,N_47300);
nor U48495 (N_48495,N_46422,N_47835);
nor U48496 (N_48496,N_47618,N_47461);
nand U48497 (N_48497,N_46961,N_47953);
nand U48498 (N_48498,N_46541,N_47029);
nand U48499 (N_48499,N_46062,N_47683);
and U48500 (N_48500,N_47891,N_46229);
and U48501 (N_48501,N_47228,N_46721);
or U48502 (N_48502,N_47040,N_46834);
nand U48503 (N_48503,N_46968,N_47107);
nand U48504 (N_48504,N_46315,N_47002);
nand U48505 (N_48505,N_46619,N_46313);
or U48506 (N_48506,N_46559,N_47952);
nor U48507 (N_48507,N_47779,N_47931);
xor U48508 (N_48508,N_47668,N_47387);
and U48509 (N_48509,N_47608,N_47954);
nand U48510 (N_48510,N_47068,N_47604);
and U48511 (N_48511,N_47320,N_47167);
nor U48512 (N_48512,N_47450,N_46346);
nor U48513 (N_48513,N_46460,N_47140);
nor U48514 (N_48514,N_46441,N_47678);
and U48515 (N_48515,N_47559,N_46248);
and U48516 (N_48516,N_46501,N_47876);
xor U48517 (N_48517,N_46699,N_46785);
nand U48518 (N_48518,N_46749,N_46595);
or U48519 (N_48519,N_47906,N_47513);
nand U48520 (N_48520,N_46791,N_46668);
nor U48521 (N_48521,N_47843,N_46800);
nor U48522 (N_48522,N_47269,N_47114);
xor U48523 (N_48523,N_46071,N_46020);
xnor U48524 (N_48524,N_46007,N_47972);
and U48525 (N_48525,N_47956,N_47682);
and U48526 (N_48526,N_46784,N_47634);
nand U48527 (N_48527,N_46512,N_46420);
or U48528 (N_48528,N_46434,N_46437);
xor U48529 (N_48529,N_46255,N_47084);
and U48530 (N_48530,N_47321,N_47296);
or U48531 (N_48531,N_46732,N_46613);
or U48532 (N_48532,N_47332,N_46411);
or U48533 (N_48533,N_46341,N_46499);
nor U48534 (N_48534,N_46738,N_46215);
nor U48535 (N_48535,N_47400,N_47111);
xor U48536 (N_48536,N_46655,N_47110);
and U48537 (N_48537,N_47554,N_46609);
nand U48538 (N_48538,N_47552,N_46337);
nor U48539 (N_48539,N_47640,N_46506);
xor U48540 (N_48540,N_47345,N_47690);
xnor U48541 (N_48541,N_47128,N_47546);
and U48542 (N_48542,N_47051,N_46165);
and U48543 (N_48543,N_46708,N_47748);
and U48544 (N_48544,N_47855,N_47192);
or U48545 (N_48545,N_46049,N_47285);
or U48546 (N_48546,N_47152,N_47566);
nor U48547 (N_48547,N_47203,N_47452);
xnor U48548 (N_48548,N_46563,N_47248);
nand U48549 (N_48549,N_47155,N_47689);
nor U48550 (N_48550,N_47252,N_46016);
xor U48551 (N_48551,N_46876,N_46122);
xnor U48552 (N_48552,N_46554,N_47861);
and U48553 (N_48553,N_47501,N_47016);
xor U48554 (N_48554,N_47717,N_46072);
xnor U48555 (N_48555,N_46816,N_46781);
nand U48556 (N_48556,N_47544,N_46130);
or U48557 (N_48557,N_47141,N_47674);
nor U48558 (N_48558,N_47887,N_46095);
nand U48559 (N_48559,N_46967,N_47918);
xor U48560 (N_48560,N_46465,N_47898);
nand U48561 (N_48561,N_46443,N_47271);
xor U48562 (N_48562,N_47333,N_47011);
and U48563 (N_48563,N_47971,N_47094);
and U48564 (N_48564,N_46319,N_46013);
xor U48565 (N_48565,N_46065,N_46683);
nand U48566 (N_48566,N_46916,N_47647);
and U48567 (N_48567,N_46466,N_46948);
or U48568 (N_48568,N_47567,N_46678);
nor U48569 (N_48569,N_47065,N_47078);
nand U48570 (N_48570,N_46163,N_47837);
or U48571 (N_48571,N_47923,N_46433);
and U48572 (N_48572,N_47353,N_46271);
or U48573 (N_48573,N_47557,N_46681);
nand U48574 (N_48574,N_46172,N_47978);
nand U48575 (N_48575,N_47471,N_46345);
xor U48576 (N_48576,N_46106,N_47629);
xnor U48577 (N_48577,N_47272,N_46330);
and U48578 (N_48578,N_46190,N_47838);
and U48579 (N_48579,N_47399,N_46261);
xnor U48580 (N_48580,N_46272,N_47170);
nor U48581 (N_48581,N_47580,N_47218);
and U48582 (N_48582,N_46993,N_46012);
and U48583 (N_48583,N_46453,N_46779);
nor U48584 (N_48584,N_47828,N_46131);
nand U48585 (N_48585,N_46893,N_46759);
or U48586 (N_48586,N_47053,N_47994);
nor U48587 (N_48587,N_47654,N_46186);
nor U48588 (N_48588,N_47827,N_46281);
nand U48589 (N_48589,N_46711,N_46806);
xor U48590 (N_48590,N_46170,N_47338);
nand U48591 (N_48591,N_47535,N_46562);
nor U48592 (N_48592,N_47787,N_46976);
nor U48593 (N_48593,N_47380,N_47024);
nand U48594 (N_48594,N_47965,N_47829);
and U48595 (N_48595,N_46217,N_46105);
and U48596 (N_48596,N_47818,N_47028);
and U48597 (N_48597,N_47732,N_47646);
nand U48598 (N_48598,N_46513,N_46335);
nand U48599 (N_48599,N_46981,N_46689);
and U48600 (N_48600,N_47430,N_47313);
and U48601 (N_48601,N_47012,N_46309);
and U48602 (N_48602,N_47565,N_46805);
or U48603 (N_48603,N_47904,N_47358);
and U48604 (N_48604,N_46907,N_46387);
or U48605 (N_48605,N_46814,N_47071);
and U48606 (N_48606,N_46322,N_46996);
xor U48607 (N_48607,N_46985,N_47368);
xnor U48608 (N_48608,N_47713,N_46461);
or U48609 (N_48609,N_47879,N_46543);
nand U48610 (N_48610,N_46412,N_47913);
nand U48611 (N_48611,N_46626,N_46989);
and U48612 (N_48612,N_47547,N_46950);
nor U48613 (N_48613,N_46196,N_47004);
nand U48614 (N_48614,N_46860,N_46092);
xnor U48615 (N_48615,N_46452,N_47859);
xnor U48616 (N_48616,N_46403,N_47973);
nor U48617 (N_48617,N_46846,N_46332);
or U48618 (N_48618,N_46099,N_46589);
nor U48619 (N_48619,N_46386,N_47384);
xnor U48620 (N_48620,N_46223,N_46868);
nand U48621 (N_48621,N_47735,N_46978);
xor U48622 (N_48622,N_47058,N_47846);
or U48623 (N_48623,N_47792,N_47784);
or U48624 (N_48624,N_46788,N_46952);
or U48625 (N_48625,N_46066,N_47522);
or U48626 (N_48626,N_46940,N_47809);
or U48627 (N_48627,N_47955,N_46225);
xnor U48628 (N_48628,N_47291,N_47241);
or U48629 (N_48629,N_46256,N_47609);
nor U48630 (N_48630,N_47088,N_47924);
xnor U48631 (N_48631,N_46797,N_46544);
or U48632 (N_48632,N_46702,N_46687);
xnor U48633 (N_48633,N_46932,N_47769);
xnor U48634 (N_48634,N_46129,N_47538);
and U48635 (N_48635,N_47998,N_46270);
xor U48636 (N_48636,N_46672,N_46314);
and U48637 (N_48637,N_47765,N_47616);
and U48638 (N_48638,N_46600,N_46884);
or U48639 (N_48639,N_46028,N_47657);
or U48640 (N_48640,N_46125,N_47014);
nor U48641 (N_48641,N_46278,N_47044);
and U48642 (N_48642,N_46670,N_46886);
nor U48643 (N_48643,N_46964,N_46633);
or U48644 (N_48644,N_47883,N_47691);
nand U48645 (N_48645,N_47701,N_47662);
and U48646 (N_48646,N_47219,N_47599);
xnor U48647 (N_48647,N_46024,N_46294);
xnor U48648 (N_48648,N_46741,N_46906);
nor U48649 (N_48649,N_46564,N_47725);
nand U48650 (N_48650,N_46005,N_47280);
xnor U48651 (N_48651,N_46837,N_47568);
or U48652 (N_48652,N_46073,N_47266);
nand U48653 (N_48653,N_47434,N_46997);
nor U48654 (N_48654,N_47577,N_47652);
nand U48655 (N_48655,N_47721,N_46823);
nor U48656 (N_48656,N_46922,N_47133);
or U48657 (N_48657,N_47698,N_47526);
nand U48658 (N_48658,N_47304,N_47842);
xor U48659 (N_48659,N_47297,N_47365);
and U48660 (N_48660,N_47146,N_47030);
nor U48661 (N_48661,N_46694,N_46321);
and U48662 (N_48662,N_47299,N_47337);
and U48663 (N_48663,N_46744,N_47444);
or U48664 (N_48664,N_46398,N_46359);
xnor U48665 (N_48665,N_47808,N_47648);
xor U48666 (N_48666,N_47622,N_47543);
or U48667 (N_48667,N_46026,N_46827);
and U48668 (N_48668,N_46531,N_46691);
nor U48669 (N_48669,N_47574,N_46890);
and U48670 (N_48670,N_46006,N_46347);
nor U48671 (N_48671,N_47157,N_47850);
xor U48672 (N_48672,N_46204,N_47251);
nand U48673 (N_48673,N_46003,N_46671);
or U48674 (N_48674,N_47653,N_46252);
or U48675 (N_48675,N_47686,N_46632);
nor U48676 (N_48676,N_46790,N_46990);
nand U48677 (N_48677,N_46254,N_47886);
nor U48678 (N_48678,N_47598,N_46179);
xnor U48679 (N_48679,N_47003,N_47937);
nand U48680 (N_48680,N_47758,N_47635);
or U48681 (N_48681,N_47385,N_47695);
or U48682 (N_48682,N_47740,N_47738);
and U48683 (N_48683,N_47210,N_47416);
and U48684 (N_48684,N_47431,N_47104);
or U48685 (N_48685,N_46444,N_47824);
and U48686 (N_48686,N_46032,N_46519);
nand U48687 (N_48687,N_46047,N_47396);
xnor U48688 (N_48688,N_47884,N_46391);
and U48689 (N_48689,N_47868,N_47663);
and U48690 (N_48690,N_47409,N_46284);
or U48691 (N_48691,N_47457,N_47488);
nor U48692 (N_48692,N_47603,N_46858);
xnor U48693 (N_48693,N_47270,N_46793);
or U48694 (N_48694,N_46867,N_46627);
xor U48695 (N_48695,N_46743,N_46946);
xnor U48696 (N_48696,N_47275,N_47394);
xnor U48697 (N_48697,N_46703,N_46596);
nor U48698 (N_48698,N_46570,N_46614);
and U48699 (N_48699,N_47372,N_46264);
or U48700 (N_48700,N_47243,N_46285);
and U48701 (N_48701,N_46550,N_46842);
xor U48702 (N_48702,N_46696,N_47819);
and U48703 (N_48703,N_47772,N_47229);
nand U48704 (N_48704,N_46516,N_46464);
or U48705 (N_48705,N_47134,N_46783);
nand U48706 (N_48706,N_46091,N_47188);
xnor U48707 (N_48707,N_47799,N_47675);
and U48708 (N_48708,N_46765,N_47441);
or U48709 (N_48709,N_47583,N_47817);
nor U48710 (N_48710,N_47988,N_47326);
or U48711 (N_48711,N_46230,N_47928);
nand U48712 (N_48712,N_47536,N_47508);
and U48713 (N_48713,N_46584,N_47625);
and U48714 (N_48714,N_46724,N_46316);
and U48715 (N_48715,N_47087,N_46713);
or U48716 (N_48716,N_47810,N_46944);
xnor U48717 (N_48717,N_47462,N_46775);
or U48718 (N_48718,N_46896,N_46164);
and U48719 (N_48719,N_47880,N_47398);
or U48720 (N_48720,N_47917,N_47974);
and U48721 (N_48721,N_46060,N_46320);
nor U48722 (N_48722,N_46534,N_47388);
nor U48723 (N_48723,N_47076,N_46389);
and U48724 (N_48724,N_46969,N_46553);
nor U48725 (N_48725,N_46035,N_46776);
or U48726 (N_48726,N_47246,N_46739);
nand U48727 (N_48727,N_47163,N_46623);
nor U48728 (N_48728,N_46046,N_46396);
and U48729 (N_48729,N_46913,N_47220);
xor U48730 (N_48730,N_47645,N_46653);
nor U48731 (N_48731,N_46293,N_47491);
and U48732 (N_48732,N_47572,N_46360);
nand U48733 (N_48733,N_47569,N_46053);
and U48734 (N_48734,N_46426,N_46476);
xnor U48735 (N_48735,N_47664,N_47911);
or U48736 (N_48736,N_47940,N_47349);
and U48737 (N_48737,N_46905,N_47022);
and U48738 (N_48738,N_47551,N_47539);
nand U48739 (N_48739,N_47612,N_47127);
nand U48740 (N_48740,N_47709,N_47137);
nor U48741 (N_48741,N_47734,N_46934);
and U48742 (N_48742,N_46772,N_46157);
nand U48743 (N_48743,N_47633,N_47760);
xor U48744 (N_48744,N_47793,N_47348);
xor U48745 (N_48745,N_46023,N_47677);
nand U48746 (N_48746,N_46572,N_47034);
and U48747 (N_48747,N_46548,N_47449);
nor U48748 (N_48748,N_46410,N_47532);
nand U48749 (N_48749,N_47055,N_47081);
and U48750 (N_48750,N_47263,N_46446);
or U48751 (N_48751,N_46161,N_46756);
and U48752 (N_48752,N_47823,N_46726);
or U48753 (N_48753,N_46174,N_47331);
xnor U48754 (N_48754,N_47293,N_47472);
xor U48755 (N_48755,N_47770,N_47318);
nand U48756 (N_48756,N_46226,N_46665);
xor U48757 (N_48757,N_47553,N_46084);
or U48758 (N_48758,N_47037,N_46569);
nor U48759 (N_48759,N_46191,N_46287);
or U48760 (N_48760,N_46522,N_46910);
nor U48761 (N_48761,N_47350,N_46050);
xor U48762 (N_48762,N_47262,N_47206);
or U48763 (N_48763,N_46221,N_47651);
and U48764 (N_48764,N_47276,N_46729);
xor U48765 (N_48765,N_46109,N_46265);
xnor U48766 (N_48766,N_46585,N_46601);
nand U48767 (N_48767,N_46575,N_47390);
xnor U48768 (N_48768,N_46469,N_47995);
nand U48769 (N_48769,N_47347,N_47857);
and U48770 (N_48770,N_46769,N_47459);
or U48771 (N_48771,N_46680,N_46888);
or U48772 (N_48772,N_47129,N_47367);
and U48773 (N_48773,N_46979,N_46971);
nand U48774 (N_48774,N_46239,N_46342);
xor U48775 (N_48775,N_47109,N_47726);
nor U48776 (N_48776,N_46124,N_46205);
nor U48777 (N_48777,N_47949,N_47265);
nor U48778 (N_48778,N_47455,N_46182);
and U48779 (N_48779,N_46371,N_46243);
and U48780 (N_48780,N_47315,N_47905);
xor U48781 (N_48781,N_47581,N_46134);
nand U48782 (N_48782,N_47941,N_46604);
nor U48783 (N_48783,N_46528,N_46447);
nand U48784 (N_48784,N_47018,N_47307);
xnor U48785 (N_48785,N_47556,N_47143);
or U48786 (N_48786,N_46660,N_46540);
and U48787 (N_48787,N_46502,N_47173);
nand U48788 (N_48788,N_46588,N_47000);
nor U48789 (N_48789,N_47414,N_46160);
xor U48790 (N_48790,N_47126,N_47767);
nand U48791 (N_48791,N_47563,N_46509);
nor U48792 (N_48792,N_46628,N_46323);
nor U48793 (N_48793,N_46325,N_47355);
nand U48794 (N_48794,N_46963,N_47346);
and U48795 (N_48795,N_47422,N_47085);
and U48796 (N_48796,N_46714,N_46545);
xnor U48797 (N_48797,N_46087,N_46495);
and U48798 (N_48798,N_47960,N_47938);
nor U48799 (N_48799,N_47516,N_47454);
nand U48800 (N_48800,N_46917,N_46777);
or U48801 (N_48801,N_46096,N_47295);
nand U48802 (N_48802,N_46063,N_47790);
xnor U48803 (N_48803,N_47290,N_46646);
or U48804 (N_48804,N_47681,N_46257);
or U48805 (N_48805,N_47381,N_47316);
or U48806 (N_48806,N_47833,N_46064);
nand U48807 (N_48807,N_46500,N_47292);
nand U48808 (N_48808,N_46173,N_46742);
nand U48809 (N_48809,N_47497,N_46351);
or U48810 (N_48810,N_46307,N_47373);
and U48811 (N_48811,N_47468,N_47910);
nor U48812 (N_48812,N_47594,N_46027);
and U48813 (N_48813,N_46731,N_46187);
nor U48814 (N_48814,N_46573,N_46497);
nor U48815 (N_48815,N_46245,N_46920);
or U48816 (N_48816,N_47820,N_46947);
and U48817 (N_48817,N_47308,N_47282);
xnor U48818 (N_48818,N_46973,N_47287);
xor U48819 (N_48819,N_46945,N_46317);
nand U48820 (N_48820,N_47151,N_47706);
xor U48821 (N_48821,N_46147,N_46177);
nor U48822 (N_48822,N_47112,N_47435);
nand U48823 (N_48823,N_47597,N_47289);
xor U48824 (N_48824,N_46128,N_47408);
or U48825 (N_48825,N_46211,N_47411);
nor U48826 (N_48826,N_47696,N_47401);
and U48827 (N_48827,N_46579,N_46908);
nand U48828 (N_48828,N_47223,N_47700);
nand U48829 (N_48829,N_47484,N_47420);
nor U48830 (N_48830,N_46608,N_47836);
nor U48831 (N_48831,N_46629,N_46111);
xnor U48832 (N_48832,N_46438,N_47202);
xor U48833 (N_48833,N_46030,N_47261);
nand U48834 (N_48834,N_46029,N_47731);
nor U48835 (N_48835,N_47800,N_47073);
and U48836 (N_48836,N_46372,N_47853);
nand U48837 (N_48837,N_47679,N_46201);
xnor U48838 (N_48838,N_46176,N_46259);
or U48839 (N_48839,N_47121,N_46088);
nand U48840 (N_48840,N_47867,N_47224);
or U48841 (N_48841,N_47666,N_46778);
or U48842 (N_48842,N_46141,N_47172);
and U48843 (N_48843,N_46773,N_47402);
xor U48844 (N_48844,N_46984,N_47038);
nor U48845 (N_48845,N_46381,N_47456);
or U48846 (N_48846,N_47803,N_46249);
xnor U48847 (N_48847,N_46197,N_47984);
and U48848 (N_48848,N_47256,N_47521);
nor U48849 (N_48849,N_47233,N_46535);
xor U48850 (N_48850,N_47794,N_46240);
and U48851 (N_48851,N_47806,N_46607);
nand U48852 (N_48852,N_46925,N_46730);
xor U48853 (N_48853,N_47967,N_47179);
xnor U48854 (N_48854,N_46353,N_47766);
nand U48855 (N_48855,N_46268,N_47639);
xnor U48856 (N_48856,N_47578,N_47946);
and U48857 (N_48857,N_47511,N_47763);
nand U48858 (N_48858,N_46676,N_47628);
nor U48859 (N_48859,N_46445,N_47267);
nor U48860 (N_48860,N_46414,N_46054);
and U48861 (N_48861,N_46937,N_47093);
xnor U48862 (N_48862,N_46340,N_46647);
nor U48863 (N_48863,N_47253,N_47214);
xnor U48864 (N_48864,N_47130,N_47284);
nor U48865 (N_48865,N_46861,N_46733);
and U48866 (N_48866,N_47947,N_47592);
or U48867 (N_48867,N_46428,N_46401);
nor U48868 (N_48868,N_47216,N_47237);
and U48869 (N_48869,N_46771,N_46637);
xor U48870 (N_48870,N_47330,N_47191);
and U48871 (N_48871,N_46156,N_47213);
and U48872 (N_48872,N_46770,N_46212);
and U48873 (N_48873,N_47590,N_47483);
nor U48874 (N_48874,N_47359,N_46811);
or U48875 (N_48875,N_47445,N_47057);
nand U48876 (N_48876,N_47255,N_46136);
xor U48877 (N_48877,N_47199,N_47281);
or U48878 (N_48878,N_47737,N_46887);
and U48879 (N_48879,N_46977,N_46008);
and U48880 (N_48880,N_47754,N_46019);
xnor U48881 (N_48881,N_47391,N_47376);
or U48882 (N_48882,N_47620,N_46684);
or U48883 (N_48883,N_46616,N_46571);
or U48884 (N_48884,N_47360,N_47103);
and U48885 (N_48885,N_46697,N_46852);
xnor U48886 (N_48886,N_46617,N_47286);
nand U48887 (N_48887,N_46207,N_46116);
nor U48888 (N_48888,N_47575,N_46017);
and U48889 (N_48889,N_46532,N_46524);
and U48890 (N_48890,N_47198,N_46056);
and U48891 (N_48891,N_47160,N_47961);
nor U48892 (N_48892,N_46404,N_47576);
and U48893 (N_48893,N_46892,N_46169);
xor U48894 (N_48894,N_47105,N_46710);
and U48895 (N_48895,N_47142,N_46231);
nor U48896 (N_48896,N_46663,N_47885);
and U48897 (N_48897,N_46986,N_47888);
xnor U48898 (N_48898,N_47101,N_46100);
nand U48899 (N_48899,N_46521,N_46155);
nor U48900 (N_48900,N_47990,N_46227);
and U48901 (N_48901,N_46664,N_47470);
or U48902 (N_48902,N_46874,N_47090);
or U48903 (N_48903,N_47339,N_46611);
xnor U48904 (N_48904,N_47564,N_46835);
or U48905 (N_48905,N_47602,N_46862);
and U48906 (N_48906,N_47582,N_47534);
and U48907 (N_48907,N_47189,N_47392);
or U48908 (N_48908,N_47215,N_46815);
xnor U48909 (N_48909,N_47650,N_47789);
nor U48910 (N_48910,N_46877,N_46953);
nor U48911 (N_48911,N_46300,N_46728);
xor U48912 (N_48912,N_46839,N_46586);
or U48913 (N_48913,N_46970,N_46652);
and U48914 (N_48914,N_46719,N_47061);
and U48915 (N_48915,N_46057,N_46641);
or U48916 (N_48916,N_47487,N_47505);
or U48917 (N_48917,N_46958,N_46144);
xnor U48918 (N_48918,N_47283,N_47759);
or U48919 (N_48919,N_46306,N_46219);
or U48920 (N_48920,N_47969,N_47643);
nor U48921 (N_48921,N_46367,N_47814);
or U48922 (N_48922,N_46168,N_46357);
and U48923 (N_48923,N_47042,N_46292);
or U48924 (N_48924,N_47200,N_46039);
nand U48925 (N_48925,N_47247,N_47447);
nand U48926 (N_48926,N_47517,N_47446);
nand U48927 (N_48927,N_47925,N_47589);
and U48928 (N_48928,N_46074,N_46955);
nand U48929 (N_48929,N_46666,N_46454);
or U48930 (N_48930,N_46994,N_47010);
or U48931 (N_48931,N_47325,N_46972);
nand U48932 (N_48932,N_47303,N_47864);
nand U48933 (N_48933,N_47724,N_47641);
and U48934 (N_48934,N_46639,N_46592);
nand U48935 (N_48935,N_47531,N_47771);
nand U48936 (N_48936,N_46184,N_46918);
xnor U48937 (N_48937,N_47710,N_46853);
nand U48938 (N_48938,N_47750,N_46305);
and U48939 (N_48939,N_46975,N_47086);
nor U48940 (N_48940,N_47498,N_46251);
or U48941 (N_48941,N_47610,N_47743);
or U48942 (N_48942,N_47796,N_46820);
nor U48943 (N_48943,N_46679,N_47187);
nand U48944 (N_48944,N_47601,N_46498);
nor U48945 (N_48945,N_47714,N_46567);
nor U48946 (N_48946,N_47523,N_47072);
nor U48947 (N_48947,N_47412,N_46112);
nor U48948 (N_48948,N_46121,N_47033);
or U48949 (N_48949,N_46642,N_47132);
and U48950 (N_48950,N_47670,N_47463);
nor U48951 (N_48951,N_47816,N_47788);
nand U48952 (N_48952,N_47922,N_46058);
and U48953 (N_48953,N_47807,N_46344);
xor U48954 (N_48954,N_46789,N_47786);
or U48955 (N_48955,N_46418,N_46260);
xor U48956 (N_48956,N_47591,N_47317);
xor U48957 (N_48957,N_46725,N_47571);
nor U48958 (N_48958,N_46118,N_46463);
nor U48959 (N_48959,N_47052,N_47507);
and U48960 (N_48960,N_47896,N_47120);
nor U48961 (N_48961,N_47503,N_46408);
xor U48962 (N_48962,N_46900,N_46957);
xnor U48963 (N_48963,N_46635,N_46624);
nand U48964 (N_48964,N_46140,N_46929);
and U48965 (N_48965,N_46350,N_46415);
or U48966 (N_48966,N_46693,N_46718);
nand U48967 (N_48967,N_47844,N_47156);
nand U48968 (N_48968,N_47377,N_47637);
or U48969 (N_48969,N_47877,N_47687);
nor U48970 (N_48970,N_47742,N_46507);
nor U48971 (N_48971,N_47605,N_47860);
or U48972 (N_48972,N_47089,N_46366);
nand U48973 (N_48973,N_46709,N_47425);
nand U48974 (N_48974,N_47595,N_46525);
nor U48975 (N_48975,N_46110,N_46537);
xnor U48976 (N_48976,N_46022,N_47627);
and U48977 (N_48977,N_47379,N_47115);
nand U48978 (N_48978,N_47064,N_46104);
xor U48979 (N_48979,N_46150,N_47144);
and U48980 (N_48980,N_47245,N_47211);
xor U48981 (N_48981,N_46851,N_47761);
or U48982 (N_48982,N_47966,N_46821);
nand U48983 (N_48983,N_46246,N_47363);
and U48984 (N_48984,N_46425,N_46974);
xor U48985 (N_48985,N_46780,N_46930);
or U48986 (N_48986,N_47872,N_46881);
or U48987 (N_48987,N_46856,N_46723);
and U48988 (N_48988,N_47588,N_46517);
or U48989 (N_48989,N_47421,N_46374);
xor U48990 (N_48990,N_47467,N_47481);
nor U48991 (N_48991,N_46178,N_47509);
nor U48992 (N_48992,N_47909,N_47746);
xnor U48993 (N_48993,N_46388,N_46233);
nor U48994 (N_48994,N_46850,N_47862);
xor U48995 (N_48995,N_46597,N_46992);
or U48996 (N_48996,N_46648,N_47231);
xor U48997 (N_48997,N_47310,N_47413);
xor U48998 (N_48998,N_46108,N_47562);
nand U48999 (N_48999,N_47361,N_47825);
nand U49000 (N_49000,N_46114,N_47966);
nand U49001 (N_49001,N_46552,N_46351);
or U49002 (N_49002,N_47517,N_47630);
xnor U49003 (N_49003,N_46615,N_46286);
and U49004 (N_49004,N_46807,N_47149);
and U49005 (N_49005,N_47296,N_46021);
xor U49006 (N_49006,N_46949,N_46049);
or U49007 (N_49007,N_47053,N_47530);
and U49008 (N_49008,N_47930,N_47029);
nor U49009 (N_49009,N_47367,N_47895);
nor U49010 (N_49010,N_47395,N_47260);
and U49011 (N_49011,N_47824,N_47099);
and U49012 (N_49012,N_46495,N_46459);
xnor U49013 (N_49013,N_47125,N_47524);
and U49014 (N_49014,N_46836,N_46653);
or U49015 (N_49015,N_47846,N_46349);
xor U49016 (N_49016,N_47590,N_47420);
or U49017 (N_49017,N_46258,N_47605);
or U49018 (N_49018,N_47549,N_47053);
nor U49019 (N_49019,N_47336,N_46323);
nor U49020 (N_49020,N_47463,N_47341);
xnor U49021 (N_49021,N_47245,N_47301);
nand U49022 (N_49022,N_46497,N_47353);
or U49023 (N_49023,N_47429,N_47084);
or U49024 (N_49024,N_47160,N_47380);
nand U49025 (N_49025,N_47288,N_47633);
or U49026 (N_49026,N_47107,N_46061);
or U49027 (N_49027,N_47881,N_46524);
or U49028 (N_49028,N_47569,N_46015);
xor U49029 (N_49029,N_47325,N_47519);
or U49030 (N_49030,N_46252,N_46571);
nand U49031 (N_49031,N_47853,N_47613);
nor U49032 (N_49032,N_46103,N_46951);
nor U49033 (N_49033,N_46836,N_47120);
nand U49034 (N_49034,N_46618,N_47201);
or U49035 (N_49035,N_47930,N_46851);
nand U49036 (N_49036,N_46806,N_47746);
nor U49037 (N_49037,N_47538,N_46168);
nor U49038 (N_49038,N_46122,N_47318);
nand U49039 (N_49039,N_46396,N_46706);
nor U49040 (N_49040,N_46960,N_46787);
or U49041 (N_49041,N_47323,N_46879);
and U49042 (N_49042,N_46251,N_47234);
nand U49043 (N_49043,N_47114,N_46268);
nand U49044 (N_49044,N_47410,N_46857);
and U49045 (N_49045,N_46806,N_46036);
and U49046 (N_49046,N_47315,N_47574);
xnor U49047 (N_49047,N_47865,N_46088);
nor U49048 (N_49048,N_47689,N_46719);
or U49049 (N_49049,N_46541,N_47668);
xnor U49050 (N_49050,N_46783,N_47803);
or U49051 (N_49051,N_47667,N_46882);
or U49052 (N_49052,N_47306,N_46055);
nand U49053 (N_49053,N_47797,N_46116);
or U49054 (N_49054,N_46345,N_47494);
xor U49055 (N_49055,N_46985,N_47312);
or U49056 (N_49056,N_47365,N_47239);
and U49057 (N_49057,N_46126,N_46546);
and U49058 (N_49058,N_47475,N_46784);
and U49059 (N_49059,N_47999,N_46251);
and U49060 (N_49060,N_46257,N_47073);
and U49061 (N_49061,N_46660,N_47584);
nor U49062 (N_49062,N_46175,N_46218);
or U49063 (N_49063,N_46054,N_47558);
xnor U49064 (N_49064,N_46790,N_46048);
nor U49065 (N_49065,N_47840,N_46326);
or U49066 (N_49066,N_46571,N_47788);
nor U49067 (N_49067,N_47485,N_47287);
nand U49068 (N_49068,N_46221,N_46794);
xor U49069 (N_49069,N_46229,N_47895);
nor U49070 (N_49070,N_47972,N_46061);
or U49071 (N_49071,N_46311,N_47466);
nor U49072 (N_49072,N_46461,N_46107);
xor U49073 (N_49073,N_47301,N_46943);
nand U49074 (N_49074,N_47097,N_46803);
or U49075 (N_49075,N_46529,N_46430);
nor U49076 (N_49076,N_46598,N_47528);
and U49077 (N_49077,N_47679,N_47582);
or U49078 (N_49078,N_46927,N_47044);
or U49079 (N_49079,N_46389,N_47498);
xnor U49080 (N_49080,N_46117,N_47898);
nand U49081 (N_49081,N_47009,N_46697);
xnor U49082 (N_49082,N_46213,N_46060);
or U49083 (N_49083,N_46174,N_47403);
nor U49084 (N_49084,N_47567,N_47406);
xnor U49085 (N_49085,N_47879,N_47582);
or U49086 (N_49086,N_47559,N_47492);
xor U49087 (N_49087,N_46067,N_47143);
or U49088 (N_49088,N_47376,N_46658);
xor U49089 (N_49089,N_46351,N_46762);
nand U49090 (N_49090,N_47919,N_47951);
and U49091 (N_49091,N_47097,N_46396);
or U49092 (N_49092,N_46473,N_47583);
and U49093 (N_49093,N_47008,N_46773);
xor U49094 (N_49094,N_47107,N_47532);
and U49095 (N_49095,N_47885,N_46867);
xor U49096 (N_49096,N_46541,N_46564);
nand U49097 (N_49097,N_47274,N_46906);
xor U49098 (N_49098,N_46202,N_47298);
xor U49099 (N_49099,N_46334,N_47156);
or U49100 (N_49100,N_46081,N_47427);
or U49101 (N_49101,N_47861,N_47830);
nor U49102 (N_49102,N_47676,N_47124);
nand U49103 (N_49103,N_46690,N_46983);
xnor U49104 (N_49104,N_47463,N_46395);
xor U49105 (N_49105,N_46189,N_47030);
xor U49106 (N_49106,N_47172,N_47413);
nor U49107 (N_49107,N_46214,N_46104);
nor U49108 (N_49108,N_47239,N_47089);
nor U49109 (N_49109,N_47043,N_46732);
xor U49110 (N_49110,N_46073,N_47167);
and U49111 (N_49111,N_46101,N_47098);
nor U49112 (N_49112,N_46799,N_46318);
nor U49113 (N_49113,N_46388,N_47836);
and U49114 (N_49114,N_47277,N_46424);
nand U49115 (N_49115,N_46023,N_47234);
and U49116 (N_49116,N_46530,N_46703);
and U49117 (N_49117,N_47900,N_46713);
xnor U49118 (N_49118,N_46954,N_46044);
nor U49119 (N_49119,N_47089,N_46400);
xnor U49120 (N_49120,N_46828,N_46673);
xnor U49121 (N_49121,N_46361,N_46046);
or U49122 (N_49122,N_46917,N_46965);
and U49123 (N_49123,N_46798,N_46780);
and U49124 (N_49124,N_46684,N_46748);
nand U49125 (N_49125,N_46059,N_47521);
nand U49126 (N_49126,N_47234,N_46081);
nor U49127 (N_49127,N_46502,N_46104);
and U49128 (N_49128,N_46850,N_46065);
and U49129 (N_49129,N_46104,N_47309);
nor U49130 (N_49130,N_47510,N_46504);
and U49131 (N_49131,N_47749,N_47027);
or U49132 (N_49132,N_47645,N_47010);
and U49133 (N_49133,N_47842,N_46979);
nand U49134 (N_49134,N_47966,N_47729);
nand U49135 (N_49135,N_47687,N_47107);
nor U49136 (N_49136,N_47504,N_47019);
or U49137 (N_49137,N_46910,N_46169);
and U49138 (N_49138,N_47131,N_47088);
and U49139 (N_49139,N_47602,N_47346);
xnor U49140 (N_49140,N_47157,N_46577);
and U49141 (N_49141,N_46181,N_47511);
and U49142 (N_49142,N_47923,N_46428);
nand U49143 (N_49143,N_47079,N_46350);
nand U49144 (N_49144,N_47063,N_47659);
xnor U49145 (N_49145,N_46561,N_47214);
nor U49146 (N_49146,N_46240,N_46840);
nor U49147 (N_49147,N_46843,N_46217);
and U49148 (N_49148,N_46336,N_47603);
nand U49149 (N_49149,N_46879,N_47902);
or U49150 (N_49150,N_47969,N_46994);
or U49151 (N_49151,N_46993,N_47831);
or U49152 (N_49152,N_46378,N_47400);
nand U49153 (N_49153,N_46145,N_47379);
nand U49154 (N_49154,N_46481,N_47257);
nand U49155 (N_49155,N_47090,N_47983);
nor U49156 (N_49156,N_46653,N_46620);
xor U49157 (N_49157,N_46524,N_46263);
xnor U49158 (N_49158,N_46653,N_47315);
xnor U49159 (N_49159,N_46981,N_47851);
and U49160 (N_49160,N_47680,N_47764);
or U49161 (N_49161,N_46188,N_47131);
or U49162 (N_49162,N_47362,N_46068);
xnor U49163 (N_49163,N_47025,N_46408);
and U49164 (N_49164,N_47394,N_46897);
xor U49165 (N_49165,N_46682,N_47431);
or U49166 (N_49166,N_47991,N_46750);
and U49167 (N_49167,N_46506,N_47881);
nor U49168 (N_49168,N_47137,N_47500);
nand U49169 (N_49169,N_46563,N_47432);
xnor U49170 (N_49170,N_47340,N_46946);
and U49171 (N_49171,N_47433,N_47080);
nand U49172 (N_49172,N_46313,N_47205);
nand U49173 (N_49173,N_47872,N_46322);
nand U49174 (N_49174,N_47550,N_46959);
nand U49175 (N_49175,N_47019,N_47390);
xnor U49176 (N_49176,N_47267,N_47518);
and U49177 (N_49177,N_47540,N_46536);
nand U49178 (N_49178,N_47494,N_47798);
nor U49179 (N_49179,N_46153,N_47802);
xor U49180 (N_49180,N_46300,N_46424);
nand U49181 (N_49181,N_47653,N_47499);
or U49182 (N_49182,N_46413,N_46717);
or U49183 (N_49183,N_46938,N_47579);
xor U49184 (N_49184,N_47833,N_46179);
and U49185 (N_49185,N_47154,N_47566);
nor U49186 (N_49186,N_46056,N_46461);
nor U49187 (N_49187,N_47472,N_46489);
and U49188 (N_49188,N_46784,N_47624);
and U49189 (N_49189,N_47085,N_47654);
xor U49190 (N_49190,N_47742,N_47415);
xor U49191 (N_49191,N_46020,N_46628);
nor U49192 (N_49192,N_47624,N_46031);
or U49193 (N_49193,N_46223,N_47507);
nand U49194 (N_49194,N_47346,N_46596);
xor U49195 (N_49195,N_47643,N_46445);
and U49196 (N_49196,N_47123,N_47649);
and U49197 (N_49197,N_46154,N_47113);
or U49198 (N_49198,N_46832,N_46164);
xor U49199 (N_49199,N_47259,N_47605);
and U49200 (N_49200,N_46347,N_47440);
and U49201 (N_49201,N_46834,N_46577);
nand U49202 (N_49202,N_47383,N_47026);
nand U49203 (N_49203,N_46157,N_46135);
nor U49204 (N_49204,N_46794,N_47737);
and U49205 (N_49205,N_46405,N_46015);
nand U49206 (N_49206,N_47294,N_46223);
nor U49207 (N_49207,N_46350,N_46417);
or U49208 (N_49208,N_46721,N_47637);
nor U49209 (N_49209,N_47289,N_46550);
xnor U49210 (N_49210,N_46470,N_47718);
nor U49211 (N_49211,N_47015,N_47310);
and U49212 (N_49212,N_46625,N_47061);
and U49213 (N_49213,N_47422,N_47278);
and U49214 (N_49214,N_46180,N_47622);
nand U49215 (N_49215,N_47154,N_47535);
nand U49216 (N_49216,N_46641,N_46346);
xnor U49217 (N_49217,N_47618,N_46500);
and U49218 (N_49218,N_47705,N_46460);
and U49219 (N_49219,N_47201,N_46298);
and U49220 (N_49220,N_47259,N_47084);
or U49221 (N_49221,N_47866,N_47700);
and U49222 (N_49222,N_47791,N_46959);
xnor U49223 (N_49223,N_47402,N_46291);
nor U49224 (N_49224,N_46283,N_46847);
or U49225 (N_49225,N_47893,N_47535);
and U49226 (N_49226,N_47750,N_47351);
and U49227 (N_49227,N_47555,N_46380);
and U49228 (N_49228,N_47755,N_47487);
xnor U49229 (N_49229,N_46069,N_47702);
and U49230 (N_49230,N_47305,N_46614);
nor U49231 (N_49231,N_46311,N_47563);
and U49232 (N_49232,N_46488,N_47696);
nand U49233 (N_49233,N_46852,N_47450);
nand U49234 (N_49234,N_47821,N_47921);
and U49235 (N_49235,N_46665,N_46454);
nor U49236 (N_49236,N_46523,N_47857);
xnor U49237 (N_49237,N_47312,N_46846);
xnor U49238 (N_49238,N_47327,N_46389);
and U49239 (N_49239,N_47025,N_47178);
nor U49240 (N_49240,N_47615,N_47983);
or U49241 (N_49241,N_47214,N_47627);
xnor U49242 (N_49242,N_46821,N_46277);
or U49243 (N_49243,N_47426,N_47185);
nand U49244 (N_49244,N_46498,N_46566);
or U49245 (N_49245,N_46477,N_47295);
or U49246 (N_49246,N_46844,N_46442);
nand U49247 (N_49247,N_46793,N_47947);
or U49248 (N_49248,N_46596,N_47544);
and U49249 (N_49249,N_46467,N_46224);
xnor U49250 (N_49250,N_46106,N_47095);
or U49251 (N_49251,N_46791,N_46148);
xnor U49252 (N_49252,N_47931,N_47842);
nand U49253 (N_49253,N_47209,N_47786);
or U49254 (N_49254,N_47831,N_47089);
and U49255 (N_49255,N_47084,N_46657);
or U49256 (N_49256,N_47010,N_47781);
or U49257 (N_49257,N_46971,N_46429);
xor U49258 (N_49258,N_47241,N_47769);
or U49259 (N_49259,N_47903,N_47819);
xor U49260 (N_49260,N_47304,N_47827);
nor U49261 (N_49261,N_46657,N_47328);
and U49262 (N_49262,N_46921,N_46691);
nor U49263 (N_49263,N_47205,N_46554);
or U49264 (N_49264,N_47862,N_47273);
xor U49265 (N_49265,N_47705,N_47720);
and U49266 (N_49266,N_47685,N_46136);
nor U49267 (N_49267,N_47808,N_47800);
xor U49268 (N_49268,N_47710,N_47034);
xor U49269 (N_49269,N_47737,N_47532);
and U49270 (N_49270,N_46668,N_46920);
and U49271 (N_49271,N_47963,N_47814);
nand U49272 (N_49272,N_47118,N_46556);
xor U49273 (N_49273,N_46453,N_47406);
or U49274 (N_49274,N_47497,N_47271);
and U49275 (N_49275,N_46169,N_47030);
xor U49276 (N_49276,N_46741,N_47387);
nor U49277 (N_49277,N_47028,N_46722);
and U49278 (N_49278,N_47614,N_46654);
xor U49279 (N_49279,N_47951,N_46848);
and U49280 (N_49280,N_47896,N_46358);
or U49281 (N_49281,N_47673,N_47742);
xnor U49282 (N_49282,N_46250,N_46803);
nand U49283 (N_49283,N_46964,N_47870);
and U49284 (N_49284,N_46328,N_47048);
xor U49285 (N_49285,N_46663,N_46809);
xor U49286 (N_49286,N_46634,N_46166);
and U49287 (N_49287,N_47760,N_46034);
or U49288 (N_49288,N_47174,N_47286);
and U49289 (N_49289,N_47884,N_47244);
nor U49290 (N_49290,N_47946,N_47382);
xor U49291 (N_49291,N_46803,N_46369);
nand U49292 (N_49292,N_46478,N_46115);
nand U49293 (N_49293,N_47707,N_47732);
nor U49294 (N_49294,N_46035,N_47909);
nor U49295 (N_49295,N_47976,N_46997);
and U49296 (N_49296,N_46499,N_46501);
xnor U49297 (N_49297,N_46292,N_47092);
nand U49298 (N_49298,N_47530,N_46553);
and U49299 (N_49299,N_46002,N_47408);
or U49300 (N_49300,N_46820,N_46291);
nor U49301 (N_49301,N_46420,N_46008);
nand U49302 (N_49302,N_46301,N_47323);
nor U49303 (N_49303,N_46379,N_47019);
nor U49304 (N_49304,N_47165,N_47798);
nand U49305 (N_49305,N_47248,N_46370);
nor U49306 (N_49306,N_46608,N_46661);
or U49307 (N_49307,N_47854,N_46355);
nor U49308 (N_49308,N_46908,N_47566);
xnor U49309 (N_49309,N_46085,N_47410);
xor U49310 (N_49310,N_47941,N_46055);
xor U49311 (N_49311,N_46040,N_47132);
or U49312 (N_49312,N_46966,N_46275);
and U49313 (N_49313,N_47448,N_46283);
nand U49314 (N_49314,N_47331,N_46512);
or U49315 (N_49315,N_47560,N_46443);
xnor U49316 (N_49316,N_47096,N_47454);
and U49317 (N_49317,N_47449,N_47418);
nand U49318 (N_49318,N_46811,N_46171);
nand U49319 (N_49319,N_46139,N_47072);
nor U49320 (N_49320,N_46164,N_47443);
xnor U49321 (N_49321,N_47483,N_47379);
and U49322 (N_49322,N_47650,N_46649);
nand U49323 (N_49323,N_46257,N_47683);
xor U49324 (N_49324,N_47586,N_46747);
nor U49325 (N_49325,N_47922,N_47382);
and U49326 (N_49326,N_46197,N_47105);
and U49327 (N_49327,N_46222,N_46256);
and U49328 (N_49328,N_46468,N_46519);
or U49329 (N_49329,N_46905,N_47822);
xnor U49330 (N_49330,N_46776,N_46778);
xnor U49331 (N_49331,N_47814,N_46991);
nand U49332 (N_49332,N_47188,N_46112);
or U49333 (N_49333,N_46343,N_47007);
nor U49334 (N_49334,N_46502,N_46648);
and U49335 (N_49335,N_46279,N_47267);
nand U49336 (N_49336,N_46206,N_47061);
xnor U49337 (N_49337,N_46074,N_46528);
xnor U49338 (N_49338,N_47116,N_46781);
xor U49339 (N_49339,N_46147,N_47951);
xor U49340 (N_49340,N_46615,N_46733);
or U49341 (N_49341,N_47507,N_46816);
or U49342 (N_49342,N_47899,N_46904);
or U49343 (N_49343,N_47585,N_47906);
xnor U49344 (N_49344,N_47235,N_46813);
nor U49345 (N_49345,N_46926,N_47913);
nand U49346 (N_49346,N_46285,N_46109);
nor U49347 (N_49347,N_46475,N_46349);
nor U49348 (N_49348,N_46759,N_46105);
xor U49349 (N_49349,N_46392,N_47042);
nor U49350 (N_49350,N_46388,N_47455);
nor U49351 (N_49351,N_47390,N_47968);
nor U49352 (N_49352,N_47106,N_46257);
nand U49353 (N_49353,N_46247,N_46169);
nand U49354 (N_49354,N_46088,N_46756);
nand U49355 (N_49355,N_46982,N_46102);
xnor U49356 (N_49356,N_46729,N_47384);
nand U49357 (N_49357,N_47174,N_46543);
and U49358 (N_49358,N_46006,N_46515);
xnor U49359 (N_49359,N_47855,N_47561);
or U49360 (N_49360,N_46798,N_46726);
or U49361 (N_49361,N_46230,N_47017);
nor U49362 (N_49362,N_47624,N_47682);
nor U49363 (N_49363,N_46891,N_47746);
nand U49364 (N_49364,N_46524,N_46827);
xor U49365 (N_49365,N_47598,N_46971);
or U49366 (N_49366,N_47050,N_47852);
or U49367 (N_49367,N_47074,N_47019);
nor U49368 (N_49368,N_47490,N_46559);
xor U49369 (N_49369,N_47216,N_46170);
nand U49370 (N_49370,N_47966,N_46768);
xor U49371 (N_49371,N_46424,N_46647);
or U49372 (N_49372,N_47965,N_47558);
xor U49373 (N_49373,N_46032,N_47776);
nor U49374 (N_49374,N_47860,N_46501);
nor U49375 (N_49375,N_46975,N_47908);
nor U49376 (N_49376,N_47058,N_46957);
nor U49377 (N_49377,N_47407,N_47077);
nor U49378 (N_49378,N_46577,N_47011);
and U49379 (N_49379,N_47149,N_47080);
xnor U49380 (N_49380,N_47958,N_46142);
or U49381 (N_49381,N_47449,N_46608);
nor U49382 (N_49382,N_47213,N_46400);
and U49383 (N_49383,N_46652,N_47636);
or U49384 (N_49384,N_46194,N_46813);
xor U49385 (N_49385,N_46405,N_46721);
nand U49386 (N_49386,N_46300,N_46042);
xor U49387 (N_49387,N_46316,N_47794);
nor U49388 (N_49388,N_46948,N_47904);
xnor U49389 (N_49389,N_46214,N_47454);
xor U49390 (N_49390,N_46244,N_46422);
nand U49391 (N_49391,N_46985,N_46965);
and U49392 (N_49392,N_47907,N_46043);
or U49393 (N_49393,N_47878,N_46860);
nand U49394 (N_49394,N_46142,N_47286);
xor U49395 (N_49395,N_46391,N_46873);
nand U49396 (N_49396,N_47003,N_47186);
nand U49397 (N_49397,N_46136,N_46702);
nand U49398 (N_49398,N_47307,N_46213);
or U49399 (N_49399,N_47588,N_46750);
and U49400 (N_49400,N_46380,N_46352);
nor U49401 (N_49401,N_46361,N_47394);
xnor U49402 (N_49402,N_46515,N_46883);
or U49403 (N_49403,N_46289,N_46121);
nor U49404 (N_49404,N_47838,N_46975);
or U49405 (N_49405,N_47991,N_47002);
or U49406 (N_49406,N_46657,N_46490);
or U49407 (N_49407,N_47313,N_47603);
nand U49408 (N_49408,N_46829,N_47676);
and U49409 (N_49409,N_46171,N_47047);
xnor U49410 (N_49410,N_47292,N_47132);
and U49411 (N_49411,N_47594,N_46940);
xor U49412 (N_49412,N_46896,N_46813);
and U49413 (N_49413,N_46474,N_46699);
nor U49414 (N_49414,N_47875,N_47723);
or U49415 (N_49415,N_47105,N_46941);
or U49416 (N_49416,N_47476,N_47055);
or U49417 (N_49417,N_47437,N_47500);
or U49418 (N_49418,N_47141,N_46180);
and U49419 (N_49419,N_47536,N_47274);
nor U49420 (N_49420,N_46459,N_47309);
nand U49421 (N_49421,N_47397,N_46926);
or U49422 (N_49422,N_47257,N_46466);
nor U49423 (N_49423,N_47876,N_47197);
nor U49424 (N_49424,N_46834,N_46890);
nand U49425 (N_49425,N_46861,N_47784);
nor U49426 (N_49426,N_46247,N_47243);
xnor U49427 (N_49427,N_46786,N_46680);
or U49428 (N_49428,N_47184,N_47724);
or U49429 (N_49429,N_46977,N_46785);
nor U49430 (N_49430,N_47327,N_46832);
nor U49431 (N_49431,N_46452,N_46208);
xnor U49432 (N_49432,N_46117,N_46244);
xor U49433 (N_49433,N_46697,N_46666);
nand U49434 (N_49434,N_46371,N_47020);
nand U49435 (N_49435,N_47585,N_46743);
nand U49436 (N_49436,N_47565,N_46258);
and U49437 (N_49437,N_46002,N_47316);
nand U49438 (N_49438,N_46401,N_47793);
nor U49439 (N_49439,N_46228,N_47341);
and U49440 (N_49440,N_47116,N_47211);
and U49441 (N_49441,N_46024,N_46329);
or U49442 (N_49442,N_46168,N_47942);
or U49443 (N_49443,N_47858,N_46043);
nand U49444 (N_49444,N_46093,N_46747);
xnor U49445 (N_49445,N_47300,N_46041);
or U49446 (N_49446,N_47114,N_47926);
xor U49447 (N_49447,N_47923,N_47813);
nand U49448 (N_49448,N_46782,N_46229);
and U49449 (N_49449,N_47022,N_46423);
nor U49450 (N_49450,N_46550,N_46052);
nor U49451 (N_49451,N_47399,N_47161);
xor U49452 (N_49452,N_46343,N_46049);
or U49453 (N_49453,N_46090,N_46237);
xnor U49454 (N_49454,N_47266,N_46901);
or U49455 (N_49455,N_46603,N_46790);
and U49456 (N_49456,N_47708,N_46064);
nand U49457 (N_49457,N_46934,N_46404);
or U49458 (N_49458,N_47542,N_46485);
and U49459 (N_49459,N_46885,N_47777);
or U49460 (N_49460,N_46871,N_47094);
xnor U49461 (N_49461,N_47875,N_46508);
and U49462 (N_49462,N_47745,N_47799);
nor U49463 (N_49463,N_47515,N_46897);
xnor U49464 (N_49464,N_47221,N_47474);
nand U49465 (N_49465,N_46728,N_46052);
or U49466 (N_49466,N_46417,N_46559);
nand U49467 (N_49467,N_47543,N_46433);
and U49468 (N_49468,N_46852,N_47458);
or U49469 (N_49469,N_47285,N_46369);
and U49470 (N_49470,N_47834,N_46603);
and U49471 (N_49471,N_46043,N_46267);
xor U49472 (N_49472,N_47905,N_46040);
nor U49473 (N_49473,N_46141,N_46723);
and U49474 (N_49474,N_47147,N_46138);
nor U49475 (N_49475,N_47135,N_46335);
nand U49476 (N_49476,N_47422,N_47542);
nor U49477 (N_49477,N_46991,N_47100);
or U49478 (N_49478,N_47441,N_46869);
or U49479 (N_49479,N_47041,N_46859);
xnor U49480 (N_49480,N_47203,N_46701);
and U49481 (N_49481,N_47530,N_47634);
xnor U49482 (N_49482,N_47090,N_46262);
nand U49483 (N_49483,N_47053,N_46306);
nand U49484 (N_49484,N_46176,N_47695);
or U49485 (N_49485,N_47433,N_46126);
and U49486 (N_49486,N_47820,N_46173);
and U49487 (N_49487,N_46455,N_46744);
nand U49488 (N_49488,N_47904,N_46630);
and U49489 (N_49489,N_46069,N_46143);
and U49490 (N_49490,N_46930,N_47597);
xor U49491 (N_49491,N_47878,N_46683);
nor U49492 (N_49492,N_47588,N_47725);
nor U49493 (N_49493,N_46642,N_47479);
and U49494 (N_49494,N_47682,N_46917);
nor U49495 (N_49495,N_46844,N_46736);
or U49496 (N_49496,N_46868,N_47375);
xor U49497 (N_49497,N_47827,N_46722);
xor U49498 (N_49498,N_47436,N_46254);
nor U49499 (N_49499,N_46973,N_46355);
or U49500 (N_49500,N_46855,N_46803);
and U49501 (N_49501,N_47366,N_46406);
and U49502 (N_49502,N_46504,N_47805);
nand U49503 (N_49503,N_46706,N_46898);
and U49504 (N_49504,N_46976,N_47830);
or U49505 (N_49505,N_46595,N_46631);
or U49506 (N_49506,N_46378,N_46676);
or U49507 (N_49507,N_46461,N_46172);
nand U49508 (N_49508,N_47659,N_46541);
or U49509 (N_49509,N_46469,N_46655);
or U49510 (N_49510,N_47943,N_46883);
nor U49511 (N_49511,N_46843,N_47284);
nor U49512 (N_49512,N_47726,N_46338);
and U49513 (N_49513,N_46383,N_47230);
xnor U49514 (N_49514,N_47036,N_47546);
xnor U49515 (N_49515,N_46932,N_47442);
or U49516 (N_49516,N_46388,N_47958);
and U49517 (N_49517,N_46970,N_46810);
nor U49518 (N_49518,N_47237,N_46191);
or U49519 (N_49519,N_46864,N_46377);
and U49520 (N_49520,N_47036,N_46930);
or U49521 (N_49521,N_46132,N_47823);
or U49522 (N_49522,N_46403,N_47428);
xnor U49523 (N_49523,N_47599,N_46313);
nor U49524 (N_49524,N_46899,N_47484);
xor U49525 (N_49525,N_46848,N_46940);
and U49526 (N_49526,N_47597,N_47587);
nand U49527 (N_49527,N_47269,N_47292);
and U49528 (N_49528,N_46266,N_47959);
nor U49529 (N_49529,N_46883,N_47617);
xnor U49530 (N_49530,N_47156,N_47379);
xnor U49531 (N_49531,N_46163,N_46250);
and U49532 (N_49532,N_47451,N_46780);
xor U49533 (N_49533,N_46289,N_47956);
or U49534 (N_49534,N_47149,N_47722);
or U49535 (N_49535,N_46336,N_47489);
and U49536 (N_49536,N_47602,N_47522);
xnor U49537 (N_49537,N_46981,N_46993);
xor U49538 (N_49538,N_46243,N_46187);
nand U49539 (N_49539,N_46879,N_46154);
nand U49540 (N_49540,N_46965,N_47493);
nand U49541 (N_49541,N_47107,N_47845);
nor U49542 (N_49542,N_47998,N_46732);
and U49543 (N_49543,N_47718,N_46501);
xor U49544 (N_49544,N_46511,N_47138);
and U49545 (N_49545,N_47985,N_47133);
xnor U49546 (N_49546,N_46978,N_47802);
or U49547 (N_49547,N_47658,N_46019);
xor U49548 (N_49548,N_47889,N_46520);
nor U49549 (N_49549,N_47066,N_46616);
and U49550 (N_49550,N_46236,N_47289);
and U49551 (N_49551,N_46777,N_47258);
or U49552 (N_49552,N_46632,N_46328);
nor U49553 (N_49553,N_47518,N_46709);
nor U49554 (N_49554,N_46537,N_47431);
and U49555 (N_49555,N_47593,N_46529);
nand U49556 (N_49556,N_47502,N_47070);
nand U49557 (N_49557,N_46017,N_46058);
xnor U49558 (N_49558,N_47080,N_47257);
xor U49559 (N_49559,N_47799,N_46823);
nand U49560 (N_49560,N_46958,N_47163);
xnor U49561 (N_49561,N_46769,N_46519);
and U49562 (N_49562,N_46151,N_46760);
and U49563 (N_49563,N_46788,N_47533);
or U49564 (N_49564,N_47289,N_47531);
nand U49565 (N_49565,N_46124,N_47266);
and U49566 (N_49566,N_47577,N_46603);
nand U49567 (N_49567,N_46193,N_47324);
or U49568 (N_49568,N_47116,N_47284);
nand U49569 (N_49569,N_46527,N_46583);
xnor U49570 (N_49570,N_46551,N_46728);
xnor U49571 (N_49571,N_47394,N_47647);
nor U49572 (N_49572,N_46911,N_46569);
xnor U49573 (N_49573,N_46966,N_46945);
or U49574 (N_49574,N_47148,N_47733);
or U49575 (N_49575,N_47776,N_46506);
and U49576 (N_49576,N_47559,N_47655);
xor U49577 (N_49577,N_47498,N_47729);
and U49578 (N_49578,N_46657,N_47099);
or U49579 (N_49579,N_47038,N_47636);
or U49580 (N_49580,N_46889,N_47764);
nand U49581 (N_49581,N_47524,N_46486);
and U49582 (N_49582,N_47483,N_46440);
nor U49583 (N_49583,N_47273,N_47433);
xnor U49584 (N_49584,N_47965,N_47332);
or U49585 (N_49585,N_46891,N_46030);
or U49586 (N_49586,N_46989,N_46105);
and U49587 (N_49587,N_46595,N_47961);
nand U49588 (N_49588,N_47085,N_47811);
nand U49589 (N_49589,N_47754,N_46739);
xnor U49590 (N_49590,N_46540,N_46412);
or U49591 (N_49591,N_47443,N_47811);
and U49592 (N_49592,N_46122,N_46668);
nand U49593 (N_49593,N_46043,N_47640);
nand U49594 (N_49594,N_47912,N_47784);
nand U49595 (N_49595,N_47220,N_47773);
nor U49596 (N_49596,N_47476,N_47495);
or U49597 (N_49597,N_47542,N_47600);
nor U49598 (N_49598,N_46974,N_47066);
nand U49599 (N_49599,N_46961,N_46161);
nor U49600 (N_49600,N_47079,N_46449);
xnor U49601 (N_49601,N_47298,N_46983);
nor U49602 (N_49602,N_47007,N_47065);
nand U49603 (N_49603,N_47141,N_47103);
nor U49604 (N_49604,N_46362,N_47602);
nor U49605 (N_49605,N_47766,N_47755);
and U49606 (N_49606,N_46032,N_47285);
nor U49607 (N_49607,N_46517,N_47229);
nor U49608 (N_49608,N_47172,N_47654);
and U49609 (N_49609,N_46836,N_46006);
and U49610 (N_49610,N_47728,N_47155);
or U49611 (N_49611,N_46279,N_47914);
nor U49612 (N_49612,N_46491,N_47299);
or U49613 (N_49613,N_46535,N_47575);
and U49614 (N_49614,N_46684,N_47338);
and U49615 (N_49615,N_47600,N_46192);
or U49616 (N_49616,N_46228,N_46163);
and U49617 (N_49617,N_47317,N_46395);
xnor U49618 (N_49618,N_46839,N_46555);
and U49619 (N_49619,N_46330,N_46980);
nor U49620 (N_49620,N_46558,N_46428);
and U49621 (N_49621,N_47305,N_47711);
and U49622 (N_49622,N_46620,N_47525);
nand U49623 (N_49623,N_47196,N_46684);
nor U49624 (N_49624,N_46095,N_47948);
xor U49625 (N_49625,N_47609,N_47659);
or U49626 (N_49626,N_46688,N_46419);
nand U49627 (N_49627,N_46117,N_47269);
xor U49628 (N_49628,N_47593,N_46241);
xor U49629 (N_49629,N_46684,N_47974);
nand U49630 (N_49630,N_46608,N_46986);
xnor U49631 (N_49631,N_47105,N_47862);
nand U49632 (N_49632,N_46402,N_46117);
xnor U49633 (N_49633,N_46041,N_47320);
nor U49634 (N_49634,N_47226,N_47842);
and U49635 (N_49635,N_46525,N_47352);
nand U49636 (N_49636,N_46021,N_46861);
or U49637 (N_49637,N_47116,N_46588);
or U49638 (N_49638,N_47596,N_46775);
nor U49639 (N_49639,N_47009,N_47986);
and U49640 (N_49640,N_46565,N_47734);
and U49641 (N_49641,N_47648,N_47338);
or U49642 (N_49642,N_46585,N_47056);
xnor U49643 (N_49643,N_46513,N_47869);
nor U49644 (N_49644,N_46188,N_46751);
and U49645 (N_49645,N_47791,N_47453);
and U49646 (N_49646,N_46654,N_46058);
nand U49647 (N_49647,N_47042,N_47586);
or U49648 (N_49648,N_46948,N_46707);
nand U49649 (N_49649,N_46601,N_46881);
xor U49650 (N_49650,N_47016,N_47502);
and U49651 (N_49651,N_47964,N_46914);
nand U49652 (N_49652,N_47268,N_46868);
and U49653 (N_49653,N_47671,N_47247);
and U49654 (N_49654,N_47479,N_47800);
nand U49655 (N_49655,N_46477,N_46528);
xor U49656 (N_49656,N_47240,N_46885);
and U49657 (N_49657,N_46501,N_46982);
or U49658 (N_49658,N_47877,N_46690);
xor U49659 (N_49659,N_47675,N_46079);
xor U49660 (N_49660,N_46306,N_46513);
nand U49661 (N_49661,N_46496,N_46875);
xor U49662 (N_49662,N_47344,N_46799);
nor U49663 (N_49663,N_47447,N_47116);
or U49664 (N_49664,N_46435,N_46314);
or U49665 (N_49665,N_47696,N_46478);
nor U49666 (N_49666,N_47752,N_47919);
and U49667 (N_49667,N_46637,N_47525);
or U49668 (N_49668,N_47969,N_47301);
or U49669 (N_49669,N_47362,N_46308);
and U49670 (N_49670,N_46226,N_46555);
nor U49671 (N_49671,N_46300,N_47975);
nor U49672 (N_49672,N_46252,N_47970);
and U49673 (N_49673,N_47007,N_47918);
nor U49674 (N_49674,N_47797,N_46847);
or U49675 (N_49675,N_47024,N_46091);
xor U49676 (N_49676,N_46046,N_47980);
or U49677 (N_49677,N_47894,N_47151);
nand U49678 (N_49678,N_47655,N_46708);
and U49679 (N_49679,N_46108,N_47483);
or U49680 (N_49680,N_46016,N_46980);
nand U49681 (N_49681,N_46091,N_46524);
or U49682 (N_49682,N_47483,N_47425);
and U49683 (N_49683,N_46630,N_46520);
and U49684 (N_49684,N_47797,N_46484);
nand U49685 (N_49685,N_46600,N_46674);
and U49686 (N_49686,N_46703,N_47443);
or U49687 (N_49687,N_46143,N_46527);
xor U49688 (N_49688,N_46149,N_46408);
xnor U49689 (N_49689,N_46486,N_46618);
and U49690 (N_49690,N_47477,N_46334);
nand U49691 (N_49691,N_47197,N_47645);
and U49692 (N_49692,N_46234,N_47238);
or U49693 (N_49693,N_46504,N_47309);
or U49694 (N_49694,N_47353,N_46328);
nand U49695 (N_49695,N_46909,N_46787);
xnor U49696 (N_49696,N_46263,N_47179);
nand U49697 (N_49697,N_46199,N_47447);
and U49698 (N_49698,N_46627,N_47425);
and U49699 (N_49699,N_47364,N_46271);
nor U49700 (N_49700,N_46002,N_47237);
and U49701 (N_49701,N_46998,N_46944);
nand U49702 (N_49702,N_46321,N_46719);
nor U49703 (N_49703,N_47254,N_46738);
nor U49704 (N_49704,N_47976,N_46300);
nor U49705 (N_49705,N_46488,N_47199);
or U49706 (N_49706,N_46368,N_46309);
or U49707 (N_49707,N_47784,N_47918);
and U49708 (N_49708,N_46879,N_46523);
xor U49709 (N_49709,N_47909,N_47976);
xnor U49710 (N_49710,N_46327,N_47166);
nor U49711 (N_49711,N_46626,N_47137);
and U49712 (N_49712,N_46813,N_47347);
or U49713 (N_49713,N_46453,N_47073);
xor U49714 (N_49714,N_47273,N_47470);
nand U49715 (N_49715,N_47888,N_47382);
and U49716 (N_49716,N_46032,N_47877);
nor U49717 (N_49717,N_46992,N_47044);
nor U49718 (N_49718,N_47297,N_46433);
nand U49719 (N_49719,N_47482,N_47304);
or U49720 (N_49720,N_46934,N_47305);
xnor U49721 (N_49721,N_47268,N_47887);
nor U49722 (N_49722,N_47665,N_47750);
xor U49723 (N_49723,N_47972,N_47315);
or U49724 (N_49724,N_46438,N_46174);
xnor U49725 (N_49725,N_47294,N_47284);
or U49726 (N_49726,N_46889,N_46010);
or U49727 (N_49727,N_47678,N_46886);
nand U49728 (N_49728,N_47282,N_46013);
or U49729 (N_49729,N_47569,N_46940);
and U49730 (N_49730,N_47533,N_46882);
xor U49731 (N_49731,N_46997,N_47735);
or U49732 (N_49732,N_46596,N_46714);
nor U49733 (N_49733,N_46593,N_47879);
xor U49734 (N_49734,N_46551,N_47994);
or U49735 (N_49735,N_47291,N_46244);
xor U49736 (N_49736,N_46635,N_47079);
and U49737 (N_49737,N_47411,N_46517);
and U49738 (N_49738,N_46619,N_46948);
nand U49739 (N_49739,N_47180,N_47022);
xor U49740 (N_49740,N_47651,N_47822);
or U49741 (N_49741,N_47471,N_47965);
and U49742 (N_49742,N_47752,N_46433);
nor U49743 (N_49743,N_47786,N_47626);
nand U49744 (N_49744,N_46472,N_46826);
or U49745 (N_49745,N_46673,N_47836);
nand U49746 (N_49746,N_46116,N_47460);
and U49747 (N_49747,N_47102,N_46959);
and U49748 (N_49748,N_47915,N_47143);
and U49749 (N_49749,N_47950,N_46025);
nand U49750 (N_49750,N_47931,N_46156);
xor U49751 (N_49751,N_47348,N_47770);
or U49752 (N_49752,N_46721,N_46525);
xnor U49753 (N_49753,N_47023,N_46949);
nand U49754 (N_49754,N_46659,N_46234);
xor U49755 (N_49755,N_47578,N_47513);
nand U49756 (N_49756,N_46590,N_46774);
nor U49757 (N_49757,N_46508,N_47426);
nor U49758 (N_49758,N_47878,N_46779);
or U49759 (N_49759,N_46231,N_46261);
nand U49760 (N_49760,N_47907,N_47321);
nand U49761 (N_49761,N_47082,N_47833);
xor U49762 (N_49762,N_47527,N_47969);
xnor U49763 (N_49763,N_46685,N_47164);
and U49764 (N_49764,N_47213,N_47381);
and U49765 (N_49765,N_46680,N_47952);
and U49766 (N_49766,N_47342,N_47776);
nor U49767 (N_49767,N_47428,N_47577);
or U49768 (N_49768,N_47293,N_46010);
nand U49769 (N_49769,N_47054,N_46295);
xor U49770 (N_49770,N_46521,N_46056);
xor U49771 (N_49771,N_46136,N_47089);
xor U49772 (N_49772,N_47279,N_46657);
xor U49773 (N_49773,N_47584,N_46062);
and U49774 (N_49774,N_47330,N_46573);
nor U49775 (N_49775,N_46590,N_46639);
xnor U49776 (N_49776,N_47228,N_47591);
nand U49777 (N_49777,N_47951,N_46919);
xor U49778 (N_49778,N_46125,N_47878);
nand U49779 (N_49779,N_47662,N_46268);
or U49780 (N_49780,N_47994,N_46994);
xnor U49781 (N_49781,N_47759,N_46271);
xnor U49782 (N_49782,N_47618,N_46931);
or U49783 (N_49783,N_47252,N_46935);
or U49784 (N_49784,N_46090,N_47168);
or U49785 (N_49785,N_47420,N_46952);
xnor U49786 (N_49786,N_47115,N_47598);
nand U49787 (N_49787,N_46421,N_46360);
and U49788 (N_49788,N_46170,N_47305);
and U49789 (N_49789,N_46552,N_47875);
or U49790 (N_49790,N_47360,N_47560);
nand U49791 (N_49791,N_47513,N_46701);
xor U49792 (N_49792,N_46752,N_46431);
nor U49793 (N_49793,N_46550,N_47500);
nand U49794 (N_49794,N_47915,N_47812);
nand U49795 (N_49795,N_46421,N_47321);
nor U49796 (N_49796,N_47573,N_46123);
nand U49797 (N_49797,N_47285,N_47777);
and U49798 (N_49798,N_47611,N_46886);
nor U49799 (N_49799,N_46193,N_47336);
or U49800 (N_49800,N_46899,N_46408);
nor U49801 (N_49801,N_47411,N_47138);
nor U49802 (N_49802,N_46251,N_46895);
nor U49803 (N_49803,N_47931,N_47418);
xor U49804 (N_49804,N_47681,N_46683);
and U49805 (N_49805,N_47387,N_46368);
xnor U49806 (N_49806,N_46549,N_46024);
nor U49807 (N_49807,N_46928,N_47911);
nand U49808 (N_49808,N_47380,N_46136);
nor U49809 (N_49809,N_46659,N_46956);
or U49810 (N_49810,N_47843,N_47451);
and U49811 (N_49811,N_47187,N_46155);
xnor U49812 (N_49812,N_47158,N_46562);
and U49813 (N_49813,N_46785,N_46623);
and U49814 (N_49814,N_46945,N_46721);
nand U49815 (N_49815,N_47029,N_46916);
or U49816 (N_49816,N_46648,N_46828);
and U49817 (N_49817,N_47554,N_47438);
xnor U49818 (N_49818,N_46257,N_47715);
nand U49819 (N_49819,N_46363,N_47584);
nor U49820 (N_49820,N_47838,N_47395);
or U49821 (N_49821,N_47440,N_46724);
xor U49822 (N_49822,N_46926,N_46177);
nor U49823 (N_49823,N_46702,N_46708);
nand U49824 (N_49824,N_46881,N_47007);
xnor U49825 (N_49825,N_46082,N_47599);
nor U49826 (N_49826,N_46507,N_46538);
xor U49827 (N_49827,N_47840,N_46207);
xnor U49828 (N_49828,N_47021,N_47062);
nor U49829 (N_49829,N_47280,N_47805);
and U49830 (N_49830,N_46062,N_47705);
nor U49831 (N_49831,N_46385,N_46254);
nor U49832 (N_49832,N_47289,N_46343);
and U49833 (N_49833,N_47797,N_46628);
nor U49834 (N_49834,N_47337,N_47294);
or U49835 (N_49835,N_46389,N_47099);
and U49836 (N_49836,N_46506,N_47943);
nand U49837 (N_49837,N_46390,N_46765);
xnor U49838 (N_49838,N_46498,N_47766);
xor U49839 (N_49839,N_47800,N_46405);
or U49840 (N_49840,N_47021,N_47586);
or U49841 (N_49841,N_47629,N_46808);
xor U49842 (N_49842,N_46774,N_46967);
xor U49843 (N_49843,N_47914,N_47747);
or U49844 (N_49844,N_46772,N_46288);
and U49845 (N_49845,N_47782,N_46704);
or U49846 (N_49846,N_46648,N_47367);
nand U49847 (N_49847,N_46962,N_46191);
and U49848 (N_49848,N_47204,N_47334);
or U49849 (N_49849,N_46745,N_46827);
xor U49850 (N_49850,N_47036,N_47181);
or U49851 (N_49851,N_46551,N_47683);
xnor U49852 (N_49852,N_47629,N_47348);
xnor U49853 (N_49853,N_46807,N_46081);
and U49854 (N_49854,N_47800,N_46739);
xnor U49855 (N_49855,N_47851,N_47581);
nor U49856 (N_49856,N_46830,N_46665);
nor U49857 (N_49857,N_47208,N_47902);
xnor U49858 (N_49858,N_47335,N_46549);
nand U49859 (N_49859,N_47481,N_47706);
nand U49860 (N_49860,N_47054,N_46912);
and U49861 (N_49861,N_47558,N_47072);
xor U49862 (N_49862,N_47801,N_47229);
xor U49863 (N_49863,N_46085,N_46600);
nor U49864 (N_49864,N_47289,N_47340);
xnor U49865 (N_49865,N_46318,N_46763);
or U49866 (N_49866,N_47021,N_46791);
and U49867 (N_49867,N_47363,N_47536);
nand U49868 (N_49868,N_46293,N_47385);
xor U49869 (N_49869,N_47087,N_46640);
nand U49870 (N_49870,N_47388,N_47690);
nor U49871 (N_49871,N_46168,N_46603);
or U49872 (N_49872,N_46207,N_47854);
and U49873 (N_49873,N_47679,N_46264);
and U49874 (N_49874,N_46346,N_47162);
nand U49875 (N_49875,N_46284,N_46604);
xor U49876 (N_49876,N_46119,N_46732);
xor U49877 (N_49877,N_46638,N_47361);
xor U49878 (N_49878,N_47202,N_46520);
nand U49879 (N_49879,N_46171,N_47946);
nand U49880 (N_49880,N_46825,N_47559);
xor U49881 (N_49881,N_46640,N_46193);
nor U49882 (N_49882,N_47828,N_46072);
and U49883 (N_49883,N_46293,N_46093);
xor U49884 (N_49884,N_46398,N_46636);
nor U49885 (N_49885,N_46734,N_47014);
nand U49886 (N_49886,N_47278,N_46760);
and U49887 (N_49887,N_46089,N_47604);
and U49888 (N_49888,N_46893,N_46550);
or U49889 (N_49889,N_47848,N_47766);
or U49890 (N_49890,N_47422,N_47544);
or U49891 (N_49891,N_47674,N_46691);
xor U49892 (N_49892,N_47461,N_47168);
nand U49893 (N_49893,N_46614,N_46460);
and U49894 (N_49894,N_46524,N_46370);
or U49895 (N_49895,N_46300,N_46810);
and U49896 (N_49896,N_46119,N_46149);
nor U49897 (N_49897,N_47016,N_47405);
or U49898 (N_49898,N_47684,N_47950);
nor U49899 (N_49899,N_47137,N_47202);
or U49900 (N_49900,N_47137,N_46407);
or U49901 (N_49901,N_47568,N_46938);
xnor U49902 (N_49902,N_47199,N_46754);
or U49903 (N_49903,N_47994,N_46713);
or U49904 (N_49904,N_46236,N_47265);
nor U49905 (N_49905,N_47436,N_46479);
xor U49906 (N_49906,N_47810,N_47090);
nor U49907 (N_49907,N_46272,N_46913);
xnor U49908 (N_49908,N_47446,N_46067);
or U49909 (N_49909,N_47718,N_46636);
nor U49910 (N_49910,N_46474,N_46246);
and U49911 (N_49911,N_46013,N_47880);
and U49912 (N_49912,N_46903,N_47613);
nand U49913 (N_49913,N_47201,N_46858);
nor U49914 (N_49914,N_46453,N_47066);
and U49915 (N_49915,N_47292,N_46435);
nand U49916 (N_49916,N_46778,N_46132);
nor U49917 (N_49917,N_46347,N_47797);
nor U49918 (N_49918,N_46100,N_46579);
and U49919 (N_49919,N_47186,N_47817);
nand U49920 (N_49920,N_47694,N_46909);
or U49921 (N_49921,N_47835,N_46413);
or U49922 (N_49922,N_47607,N_47755);
nand U49923 (N_49923,N_46171,N_47898);
and U49924 (N_49924,N_46163,N_47778);
xor U49925 (N_49925,N_47663,N_47999);
or U49926 (N_49926,N_47624,N_47840);
or U49927 (N_49927,N_46415,N_47942);
nand U49928 (N_49928,N_46170,N_46535);
nor U49929 (N_49929,N_46042,N_46062);
nor U49930 (N_49930,N_47490,N_46562);
and U49931 (N_49931,N_47324,N_46830);
xnor U49932 (N_49932,N_47410,N_47669);
xor U49933 (N_49933,N_46801,N_46235);
nand U49934 (N_49934,N_47599,N_46913);
xor U49935 (N_49935,N_47219,N_46701);
or U49936 (N_49936,N_46138,N_47882);
and U49937 (N_49937,N_46228,N_47936);
nand U49938 (N_49938,N_46290,N_46819);
nor U49939 (N_49939,N_47440,N_47342);
nand U49940 (N_49940,N_46716,N_47474);
or U49941 (N_49941,N_47760,N_46584);
nor U49942 (N_49942,N_46343,N_46548);
nand U49943 (N_49943,N_47993,N_46498);
xnor U49944 (N_49944,N_46694,N_46276);
xnor U49945 (N_49945,N_46916,N_47952);
nand U49946 (N_49946,N_47572,N_46204);
xor U49947 (N_49947,N_46763,N_47930);
nand U49948 (N_49948,N_47377,N_46308);
xnor U49949 (N_49949,N_46610,N_47307);
and U49950 (N_49950,N_47894,N_46016);
nor U49951 (N_49951,N_47433,N_47308);
xor U49952 (N_49952,N_47550,N_46721);
nor U49953 (N_49953,N_47351,N_47588);
xnor U49954 (N_49954,N_46319,N_47770);
nor U49955 (N_49955,N_46144,N_47213);
xnor U49956 (N_49956,N_46075,N_46545);
xor U49957 (N_49957,N_47323,N_47413);
or U49958 (N_49958,N_46368,N_46638);
and U49959 (N_49959,N_47784,N_46862);
and U49960 (N_49960,N_46713,N_46002);
nand U49961 (N_49961,N_46165,N_46732);
nor U49962 (N_49962,N_47166,N_46845);
or U49963 (N_49963,N_46750,N_46235);
xor U49964 (N_49964,N_46939,N_46407);
nor U49965 (N_49965,N_47414,N_46343);
nand U49966 (N_49966,N_46004,N_47466);
or U49967 (N_49967,N_46830,N_46110);
or U49968 (N_49968,N_46688,N_46273);
xor U49969 (N_49969,N_47681,N_47909);
nand U49970 (N_49970,N_47710,N_46110);
nand U49971 (N_49971,N_47204,N_46929);
or U49972 (N_49972,N_47464,N_46194);
and U49973 (N_49973,N_47050,N_47109);
nand U49974 (N_49974,N_46851,N_47456);
and U49975 (N_49975,N_47739,N_46300);
or U49976 (N_49976,N_47223,N_46890);
nand U49977 (N_49977,N_47761,N_46015);
nor U49978 (N_49978,N_47872,N_47041);
and U49979 (N_49979,N_47417,N_47004);
nor U49980 (N_49980,N_47085,N_46711);
nand U49981 (N_49981,N_46402,N_46850);
xnor U49982 (N_49982,N_47346,N_47857);
xor U49983 (N_49983,N_46365,N_46857);
and U49984 (N_49984,N_47314,N_46187);
nand U49985 (N_49985,N_46859,N_47918);
nor U49986 (N_49986,N_47362,N_46736);
or U49987 (N_49987,N_46403,N_46810);
nand U49988 (N_49988,N_46816,N_47889);
or U49989 (N_49989,N_47414,N_46742);
or U49990 (N_49990,N_46245,N_47318);
xor U49991 (N_49991,N_47810,N_46025);
or U49992 (N_49992,N_46907,N_46608);
nand U49993 (N_49993,N_47918,N_47958);
nand U49994 (N_49994,N_46176,N_47058);
and U49995 (N_49995,N_46416,N_46134);
or U49996 (N_49996,N_46322,N_46956);
nor U49997 (N_49997,N_47536,N_47253);
xor U49998 (N_49998,N_46739,N_47702);
nand U49999 (N_49999,N_47271,N_47800);
nor UO_0 (O_0,N_49669,N_49703);
nand UO_1 (O_1,N_48713,N_49149);
xnor UO_2 (O_2,N_49325,N_48623);
or UO_3 (O_3,N_49462,N_48900);
or UO_4 (O_4,N_49518,N_48437);
xor UO_5 (O_5,N_48467,N_48994);
and UO_6 (O_6,N_49015,N_49282);
xor UO_7 (O_7,N_49562,N_49289);
or UO_8 (O_8,N_48884,N_49117);
nand UO_9 (O_9,N_48554,N_49083);
or UO_10 (O_10,N_48950,N_49308);
nor UO_11 (O_11,N_49391,N_48400);
xor UO_12 (O_12,N_48429,N_48225);
and UO_13 (O_13,N_48911,N_48822);
nand UO_14 (O_14,N_48439,N_49121);
xor UO_15 (O_15,N_48552,N_49965);
xnor UO_16 (O_16,N_49489,N_48710);
or UO_17 (O_17,N_48798,N_48540);
nor UO_18 (O_18,N_49850,N_48396);
or UO_19 (O_19,N_49789,N_48243);
or UO_20 (O_20,N_49095,N_48779);
nand UO_21 (O_21,N_48919,N_48344);
nand UO_22 (O_22,N_48522,N_48685);
xnor UO_23 (O_23,N_49376,N_49655);
xor UO_24 (O_24,N_49947,N_49682);
nand UO_25 (O_25,N_48741,N_48062);
and UO_26 (O_26,N_49998,N_48456);
and UO_27 (O_27,N_49649,N_48935);
nor UO_28 (O_28,N_48416,N_48244);
and UO_29 (O_29,N_49700,N_49480);
nor UO_30 (O_30,N_48667,N_48515);
and UO_31 (O_31,N_48765,N_49260);
and UO_32 (O_32,N_48715,N_49668);
xnor UO_33 (O_33,N_48252,N_49296);
nor UO_34 (O_34,N_49973,N_49805);
nand UO_35 (O_35,N_48378,N_48510);
and UO_36 (O_36,N_48938,N_49370);
nand UO_37 (O_37,N_48991,N_48732);
nand UO_38 (O_38,N_48721,N_48015);
xor UO_39 (O_39,N_49096,N_48695);
or UO_40 (O_40,N_49999,N_49497);
xnor UO_41 (O_41,N_48035,N_49092);
and UO_42 (O_42,N_49544,N_49596);
nand UO_43 (O_43,N_48782,N_49016);
nor UO_44 (O_44,N_49206,N_48292);
or UO_45 (O_45,N_49113,N_49635);
xnor UO_46 (O_46,N_49283,N_48356);
nor UO_47 (O_47,N_49127,N_49255);
nand UO_48 (O_48,N_48983,N_48608);
nor UO_49 (O_49,N_49483,N_49560);
and UO_50 (O_50,N_48574,N_48915);
nand UO_51 (O_51,N_49890,N_49458);
xnor UO_52 (O_52,N_49392,N_48187);
nand UO_53 (O_53,N_48219,N_49464);
and UO_54 (O_54,N_49258,N_48113);
and UO_55 (O_55,N_48290,N_48431);
nor UO_56 (O_56,N_48004,N_49160);
nand UO_57 (O_57,N_49532,N_49443);
nand UO_58 (O_58,N_49214,N_48230);
nor UO_59 (O_59,N_49666,N_49374);
nand UO_60 (O_60,N_49387,N_49050);
nor UO_61 (O_61,N_49102,N_48382);
nand UO_62 (O_62,N_49781,N_49119);
nand UO_63 (O_63,N_48310,N_48862);
xnor UO_64 (O_64,N_48912,N_49447);
or UO_65 (O_65,N_49995,N_49234);
and UO_66 (O_66,N_49075,N_48160);
or UO_67 (O_67,N_48955,N_49424);
nor UO_68 (O_68,N_49077,N_48897);
and UO_69 (O_69,N_48235,N_49974);
nand UO_70 (O_70,N_48642,N_49369);
nor UO_71 (O_71,N_49902,N_48261);
nor UO_72 (O_72,N_48363,N_48968);
nor UO_73 (O_73,N_49826,N_49907);
and UO_74 (O_74,N_48211,N_48253);
or UO_75 (O_75,N_49247,N_48568);
or UO_76 (O_76,N_48750,N_48107);
nor UO_77 (O_77,N_49870,N_48240);
nor UO_78 (O_78,N_49082,N_48156);
and UO_79 (O_79,N_49660,N_49626);
nor UO_80 (O_80,N_48829,N_48943);
nor UO_81 (O_81,N_48877,N_49768);
and UO_82 (O_82,N_49802,N_48996);
nor UO_83 (O_83,N_49719,N_48179);
or UO_84 (O_84,N_49909,N_48098);
or UO_85 (O_85,N_49548,N_48759);
nand UO_86 (O_86,N_49963,N_48631);
or UO_87 (O_87,N_48360,N_48946);
or UO_88 (O_88,N_49236,N_49257);
nor UO_89 (O_89,N_49949,N_49344);
xor UO_90 (O_90,N_49832,N_48327);
xor UO_91 (O_91,N_49526,N_48508);
nor UO_92 (O_92,N_49593,N_48802);
or UO_93 (O_93,N_49686,N_49295);
xor UO_94 (O_94,N_48890,N_49294);
nor UO_95 (O_95,N_49120,N_49100);
xor UO_96 (O_96,N_48742,N_49776);
and UO_97 (O_97,N_48628,N_48135);
xnor UO_98 (O_98,N_49453,N_49499);
and UO_99 (O_99,N_49473,N_49767);
xor UO_100 (O_100,N_48982,N_49908);
or UO_101 (O_101,N_48720,N_49905);
nand UO_102 (O_102,N_49208,N_49863);
nor UO_103 (O_103,N_49601,N_48293);
and UO_104 (O_104,N_48056,N_49235);
xnor UO_105 (O_105,N_49403,N_49530);
nand UO_106 (O_106,N_49381,N_48579);
and UO_107 (O_107,N_48743,N_49617);
or UO_108 (O_108,N_49492,N_49290);
xor UO_109 (O_109,N_49709,N_49270);
or UO_110 (O_110,N_49068,N_49089);
and UO_111 (O_111,N_49419,N_49031);
nand UO_112 (O_112,N_48825,N_49272);
nor UO_113 (O_113,N_49036,N_49969);
nand UO_114 (O_114,N_49239,N_48347);
nand UO_115 (O_115,N_48975,N_49051);
xnor UO_116 (O_116,N_48899,N_49181);
nand UO_117 (O_117,N_48154,N_49972);
or UO_118 (O_118,N_49529,N_49074);
nand UO_119 (O_119,N_48415,N_48972);
nand UO_120 (O_120,N_49631,N_49343);
xor UO_121 (O_121,N_48881,N_48678);
or UO_122 (O_122,N_49506,N_48419);
and UO_123 (O_123,N_49538,N_48316);
xnor UO_124 (O_124,N_49306,N_49007);
or UO_125 (O_125,N_48397,N_49689);
and UO_126 (O_126,N_48538,N_48161);
xnor UO_127 (O_127,N_48085,N_49049);
or UO_128 (O_128,N_48818,N_49612);
xnor UO_129 (O_129,N_49494,N_48158);
and UO_130 (O_130,N_48859,N_48236);
or UO_131 (O_131,N_48755,N_48521);
or UO_132 (O_132,N_49345,N_48573);
and UO_133 (O_133,N_48973,N_48242);
nor UO_134 (O_134,N_49903,N_49211);
or UO_135 (O_135,N_48557,N_49542);
xor UO_136 (O_136,N_48686,N_48263);
xnor UO_137 (O_137,N_49503,N_48927);
or UO_138 (O_138,N_49076,N_49812);
and UO_139 (O_139,N_48426,N_48934);
and UO_140 (O_140,N_49845,N_49365);
xor UO_141 (O_141,N_48599,N_49558);
xnor UO_142 (O_142,N_48998,N_49399);
xnor UO_143 (O_143,N_48902,N_48339);
and UO_144 (O_144,N_48365,N_48016);
and UO_145 (O_145,N_49001,N_49070);
nand UO_146 (O_146,N_49157,N_48870);
xnor UO_147 (O_147,N_48485,N_48793);
nand UO_148 (O_148,N_48030,N_49749);
nor UO_149 (O_149,N_48335,N_49440);
and UO_150 (O_150,N_48479,N_49245);
and UO_151 (O_151,N_48848,N_48851);
xnor UO_152 (O_152,N_48895,N_49733);
nor UO_153 (O_153,N_49913,N_49069);
and UO_154 (O_154,N_49755,N_48957);
nand UO_155 (O_155,N_48550,N_49607);
xnor UO_156 (O_156,N_48379,N_49196);
nand UO_157 (O_157,N_48644,N_48398);
and UO_158 (O_158,N_48860,N_49303);
and UO_159 (O_159,N_48372,N_49271);
nand UO_160 (O_160,N_49982,N_48208);
xnor UO_161 (O_161,N_49977,N_48639);
and UO_162 (O_162,N_49004,N_49348);
nor UO_163 (O_163,N_48115,N_48455);
nand UO_164 (O_164,N_49524,N_48120);
and UO_165 (O_165,N_48952,N_49991);
xnor UO_166 (O_166,N_49843,N_49279);
and UO_167 (O_167,N_49167,N_49528);
nand UO_168 (O_168,N_49860,N_49823);
nor UO_169 (O_169,N_49925,N_48032);
nand UO_170 (O_170,N_48979,N_49638);
or UO_171 (O_171,N_49411,N_49984);
xor UO_172 (O_172,N_48254,N_48764);
nand UO_173 (O_173,N_48110,N_48108);
and UO_174 (O_174,N_49468,N_49109);
xnor UO_175 (O_175,N_48931,N_48215);
nand UO_176 (O_176,N_48509,N_48487);
or UO_177 (O_177,N_49501,N_48141);
xnor UO_178 (O_178,N_49861,N_49414);
or UO_179 (O_179,N_49899,N_48852);
xor UO_180 (O_180,N_48704,N_48441);
xor UO_181 (O_181,N_48925,N_49441);
nor UO_182 (O_182,N_48582,N_48100);
and UO_183 (O_183,N_48696,N_49243);
xnor UO_184 (O_184,N_49652,N_49418);
and UO_185 (O_185,N_48993,N_48638);
nor UO_186 (O_186,N_48505,N_49293);
and UO_187 (O_187,N_49624,N_49135);
and UO_188 (O_188,N_48780,N_48662);
or UO_189 (O_189,N_49107,N_49675);
xnor UO_190 (O_190,N_49372,N_49207);
xnor UO_191 (O_191,N_49807,N_49922);
xor UO_192 (O_192,N_48036,N_49757);
nand UO_193 (O_193,N_48178,N_48361);
nand UO_194 (O_194,N_49362,N_49531);
xnor UO_195 (O_195,N_48130,N_48025);
nand UO_196 (O_196,N_48346,N_48393);
nor UO_197 (O_197,N_48525,N_48207);
xor UO_198 (O_198,N_48893,N_49151);
or UO_199 (O_199,N_48082,N_49246);
nor UO_200 (O_200,N_48280,N_49831);
nand UO_201 (O_201,N_48116,N_49536);
xor UO_202 (O_202,N_48921,N_49305);
or UO_203 (O_203,N_48733,N_48204);
and UO_204 (O_204,N_48808,N_48420);
xnor UO_205 (O_205,N_49307,N_49620);
and UO_206 (O_206,N_48433,N_48997);
nand UO_207 (O_207,N_48708,N_49046);
xnor UO_208 (O_208,N_48237,N_49364);
nand UO_209 (O_209,N_48677,N_49882);
and UO_210 (O_210,N_49192,N_48812);
nor UO_211 (O_211,N_49734,N_49093);
nor UO_212 (O_212,N_49793,N_48326);
xor UO_213 (O_213,N_48145,N_48387);
or UO_214 (O_214,N_49797,N_48071);
nand UO_215 (O_215,N_48806,N_49985);
and UO_216 (O_216,N_48754,N_49566);
and UO_217 (O_217,N_48033,N_49367);
xnor UO_218 (O_218,N_49934,N_49912);
or UO_219 (O_219,N_49152,N_48435);
nand UO_220 (O_220,N_49729,N_48049);
or UO_221 (O_221,N_49815,N_48267);
nand UO_222 (O_222,N_49375,N_48665);
and UO_223 (O_223,N_48556,N_49926);
or UO_224 (O_224,N_48362,N_49401);
nor UO_225 (O_225,N_49397,N_48588);
nor UO_226 (O_226,N_48513,N_49487);
nor UO_227 (O_227,N_48453,N_48184);
xor UO_228 (O_228,N_49302,N_49130);
and UO_229 (O_229,N_48432,N_48101);
or UO_230 (O_230,N_48930,N_49516);
nand UO_231 (O_231,N_48039,N_48059);
or UO_232 (O_232,N_48007,N_48080);
and UO_233 (O_233,N_48641,N_49361);
or UO_234 (O_234,N_48675,N_49030);
nand UO_235 (O_235,N_48700,N_48121);
xor UO_236 (O_236,N_49554,N_49339);
or UO_237 (O_237,N_49939,N_48447);
and UO_238 (O_238,N_49433,N_49416);
or UO_239 (O_239,N_48804,N_48132);
and UO_240 (O_240,N_48606,N_48969);
nand UO_241 (O_241,N_48923,N_49654);
or UO_242 (O_242,N_49262,N_48868);
or UO_243 (O_243,N_48180,N_49980);
xnor UO_244 (O_244,N_49047,N_49696);
nand UO_245 (O_245,N_49502,N_49975);
xor UO_246 (O_246,N_48916,N_48451);
and UO_247 (O_247,N_48034,N_49604);
nand UO_248 (O_248,N_48268,N_48075);
xnor UO_249 (O_249,N_48773,N_49485);
or UO_250 (O_250,N_48601,N_49616);
xor UO_251 (O_251,N_49818,N_49880);
or UO_252 (O_252,N_49436,N_49780);
nor UO_253 (O_253,N_49563,N_49978);
nor UO_254 (O_254,N_49849,N_48459);
nor UO_255 (O_255,N_49058,N_48289);
and UO_256 (O_256,N_49968,N_48664);
nand UO_257 (O_257,N_48707,N_48257);
and UO_258 (O_258,N_49929,N_49210);
and UO_259 (O_259,N_48216,N_48645);
nor UO_260 (O_260,N_49123,N_48711);
xor UO_261 (O_261,N_49546,N_49814);
nor UO_262 (O_262,N_49966,N_48443);
nor UO_263 (O_263,N_49432,N_48724);
and UO_264 (O_264,N_48234,N_49013);
and UO_265 (O_265,N_49280,N_49162);
xor UO_266 (O_266,N_49565,N_48112);
and UO_267 (O_267,N_49273,N_48649);
xnor UO_268 (O_268,N_48152,N_48618);
nor UO_269 (O_269,N_49088,N_48694);
and UO_270 (O_270,N_49000,N_49512);
xnor UO_271 (O_271,N_49352,N_48144);
or UO_272 (O_272,N_48669,N_49628);
nand UO_273 (O_273,N_48408,N_49856);
or UO_274 (O_274,N_48373,N_49541);
and UO_275 (O_275,N_48679,N_48600);
nand UO_276 (O_276,N_48507,N_49037);
nand UO_277 (O_277,N_49324,N_49510);
xnor UO_278 (O_278,N_48406,N_48567);
nand UO_279 (O_279,N_49571,N_48102);
or UO_280 (O_280,N_49382,N_48321);
nor UO_281 (O_281,N_49263,N_49938);
nand UO_282 (O_282,N_49569,N_48846);
nand UO_283 (O_283,N_49952,N_49951);
or UO_284 (O_284,N_49062,N_49222);
xor UO_285 (O_285,N_49646,N_49932);
nand UO_286 (O_286,N_48496,N_48084);
nand UO_287 (O_287,N_49836,N_49317);
or UO_288 (O_288,N_49378,N_48264);
xnor UO_289 (O_289,N_48587,N_49958);
or UO_290 (O_290,N_49390,N_48723);
and UO_291 (O_291,N_49924,N_49131);
and UO_292 (O_292,N_49170,N_49828);
nand UO_293 (O_293,N_48570,N_48519);
nand UO_294 (O_294,N_49105,N_48622);
nand UO_295 (O_295,N_49981,N_49261);
nand UO_296 (O_296,N_48605,N_49987);
or UO_297 (O_297,N_49479,N_48248);
nor UO_298 (O_298,N_49163,N_49347);
xor UO_299 (O_299,N_48005,N_49681);
xnor UO_300 (O_300,N_48562,N_49786);
or UO_301 (O_301,N_48886,N_48183);
xnor UO_302 (O_302,N_49629,N_48046);
or UO_303 (O_303,N_49385,N_48218);
and UO_304 (O_304,N_48962,N_48474);
and UO_305 (O_305,N_49720,N_48539);
nor UO_306 (O_306,N_48729,N_48330);
nand UO_307 (O_307,N_49971,N_48091);
xnor UO_308 (O_308,N_48936,N_48630);
or UO_309 (O_309,N_49673,N_49314);
nor UO_310 (O_310,N_49758,N_49683);
nor UO_311 (O_311,N_48559,N_48551);
or UO_312 (O_312,N_49901,N_48809);
and UO_313 (O_313,N_49388,N_48146);
and UO_314 (O_314,N_49085,N_49622);
nor UO_315 (O_315,N_49227,N_48576);
nor UO_316 (O_316,N_49841,N_49064);
and UO_317 (O_317,N_48528,N_48546);
and UO_318 (O_318,N_48865,N_49379);
nor UO_319 (O_319,N_48027,N_48652);
xor UO_320 (O_320,N_49623,N_49816);
and UO_321 (O_321,N_49108,N_48635);
nor UO_322 (O_322,N_48625,N_48399);
nand UO_323 (O_323,N_48555,N_48749);
nor UO_324 (O_324,N_48309,N_48634);
xnor UO_325 (O_325,N_49943,N_48872);
or UO_326 (O_326,N_49900,N_49745);
or UO_327 (O_327,N_48853,N_48947);
or UO_328 (O_328,N_49481,N_48910);
nand UO_329 (O_329,N_48940,N_49034);
nor UO_330 (O_330,N_49886,N_49155);
nand UO_331 (O_331,N_48355,N_48295);
nand UO_332 (O_332,N_49773,N_49664);
or UO_333 (O_333,N_48125,N_48799);
and UO_334 (O_334,N_48527,N_48908);
nand UO_335 (O_335,N_49421,N_48195);
xnor UO_336 (O_336,N_49523,N_49876);
nor UO_337 (O_337,N_49360,N_49663);
nand UO_338 (O_338,N_48718,N_48409);
nand UO_339 (O_339,N_48864,N_49422);
nand UO_340 (O_340,N_49463,N_48055);
and UO_341 (O_341,N_48383,N_48746);
nand UO_342 (O_342,N_49126,N_48045);
and UO_343 (O_343,N_48029,N_48315);
nor UO_344 (O_344,N_48022,N_48772);
xnor UO_345 (O_345,N_49410,N_49389);
nand UO_346 (O_346,N_49318,N_49241);
xor UO_347 (O_347,N_48421,N_48756);
nand UO_348 (O_348,N_49368,N_48354);
nor UO_349 (O_349,N_48122,N_49825);
and UO_350 (O_350,N_49630,N_48709);
or UO_351 (O_351,N_48461,N_49790);
xor UO_352 (O_352,N_49430,N_48970);
nor UO_353 (O_353,N_49132,N_49930);
nor UO_354 (O_354,N_48739,N_48514);
xor UO_355 (O_355,N_48768,N_49509);
or UO_356 (O_356,N_49237,N_49285);
nor UO_357 (O_357,N_49642,N_48963);
xnor UO_358 (O_358,N_48980,N_48604);
and UO_359 (O_359,N_49619,N_48698);
nand UO_360 (O_360,N_49471,N_49465);
and UO_361 (O_361,N_49704,N_49099);
nor UO_362 (O_362,N_49967,N_48942);
nand UO_363 (O_363,N_48735,N_49573);
nor UO_364 (O_364,N_49752,N_49184);
and UO_365 (O_365,N_48123,N_49041);
or UO_366 (O_366,N_49976,N_48444);
and UO_367 (O_367,N_48212,N_48815);
or UO_368 (O_368,N_49060,N_49110);
nand UO_369 (O_369,N_48270,N_49459);
or UO_370 (O_370,N_48014,N_49787);
xor UO_371 (O_371,N_48291,N_49919);
nand UO_372 (O_372,N_49676,N_49835);
and UO_373 (O_373,N_49627,N_49784);
nand UO_374 (O_374,N_49803,N_49201);
nor UO_375 (O_375,N_49396,N_49687);
xnor UO_376 (O_376,N_48480,N_49026);
or UO_377 (O_377,N_49104,N_49144);
nand UO_378 (O_378,N_48151,N_49645);
or UO_379 (O_379,N_49625,N_49817);
xor UO_380 (O_380,N_48182,N_48563);
nor UO_381 (O_381,N_48838,N_48048);
or UO_382 (O_382,N_48840,N_48358);
or UO_383 (O_383,N_49173,N_49274);
or UO_384 (O_384,N_49002,N_48428);
or UO_385 (O_385,N_49953,N_49840);
nor UO_386 (O_386,N_48438,N_49553);
nand UO_387 (O_387,N_49266,N_48308);
nor UO_388 (O_388,N_48352,N_49640);
and UO_389 (O_389,N_48651,N_48299);
or UO_390 (O_390,N_49839,N_48671);
xnor UO_391 (O_391,N_49848,N_49986);
and UO_392 (O_392,N_49819,N_48464);
nand UO_393 (O_393,N_48850,N_48092);
or UO_394 (O_394,N_48659,N_48117);
nor UO_395 (O_395,N_49042,N_49508);
nor UO_396 (O_396,N_49587,N_48589);
or UO_397 (O_397,N_49714,N_49288);
xor UO_398 (O_398,N_49993,N_48894);
xor UO_399 (O_399,N_48164,N_49224);
xnor UO_400 (O_400,N_49496,N_48757);
or UO_401 (O_401,N_49732,N_48458);
xnor UO_402 (O_402,N_48405,N_48560);
or UO_403 (O_403,N_48073,N_49721);
nand UO_404 (O_404,N_48167,N_49177);
xnor UO_405 (O_405,N_49128,N_48534);
or UO_406 (O_406,N_48227,N_48281);
or UO_407 (O_407,N_49338,N_48127);
nor UO_408 (O_408,N_48078,N_48325);
and UO_409 (O_409,N_48484,N_48826);
xor UO_410 (O_410,N_49086,N_48901);
and UO_411 (O_411,N_49159,N_48909);
nand UO_412 (O_412,N_49012,N_49188);
and UO_413 (O_413,N_49024,N_49568);
nand UO_414 (O_414,N_49961,N_48767);
nand UO_415 (O_415,N_48914,N_49810);
and UO_416 (O_416,N_49864,N_48465);
nor UO_417 (O_417,N_49738,N_48319);
or UO_418 (O_418,N_49543,N_48186);
and UO_419 (O_419,N_49218,N_49168);
xor UO_420 (O_420,N_48386,N_49754);
and UO_421 (O_421,N_49634,N_49021);
or UO_422 (O_422,N_48828,N_49112);
and UO_423 (O_423,N_49599,N_49500);
nor UO_424 (O_424,N_49498,N_49923);
or UO_425 (O_425,N_49442,N_48265);
xor UO_426 (O_426,N_49641,N_48333);
and UO_427 (O_427,N_48964,N_48811);
nand UO_428 (O_428,N_49467,N_49723);
or UO_429 (O_429,N_49346,N_48857);
or UO_430 (O_430,N_49588,N_49847);
xnor UO_431 (O_431,N_49935,N_48418);
or UO_432 (O_432,N_49190,N_48136);
or UO_433 (O_433,N_48626,N_48607);
or UO_434 (O_434,N_48021,N_48329);
nor UO_435 (O_435,N_48401,N_49292);
xor UO_436 (O_436,N_48760,N_48904);
or UO_437 (O_437,N_48954,N_49281);
and UO_438 (O_438,N_48512,N_48486);
nand UO_439 (O_439,N_49320,N_49028);
xnor UO_440 (O_440,N_48462,N_48803);
and UO_441 (O_441,N_49040,N_48371);
nand UO_442 (O_442,N_49079,N_48017);
nor UO_443 (O_443,N_49697,N_48200);
and UO_444 (O_444,N_48673,N_49595);
nand UO_445 (O_445,N_48882,N_48226);
or UO_446 (O_446,N_49373,N_48932);
or UO_447 (O_447,N_49022,N_48198);
or UO_448 (O_448,N_49006,N_48390);
and UO_449 (O_449,N_48341,N_48181);
xnor UO_450 (O_450,N_48874,N_49765);
or UO_451 (O_451,N_49897,N_49896);
or UO_452 (O_452,N_49066,N_49778);
xnor UO_453 (O_453,N_48959,N_49834);
nand UO_454 (O_454,N_48770,N_49065);
nand UO_455 (O_455,N_48504,N_49194);
or UO_456 (O_456,N_48883,N_49098);
or UO_457 (O_457,N_49232,N_49078);
xnor UO_458 (O_458,N_49122,N_49517);
or UO_459 (O_459,N_49106,N_48222);
nor UO_460 (O_460,N_48585,N_49337);
nand UO_461 (O_461,N_49670,N_49353);
or UO_462 (O_462,N_48984,N_49942);
or UO_463 (O_463,N_49514,N_48469);
nor UO_464 (O_464,N_49142,N_49063);
nor UO_465 (O_465,N_49695,N_48369);
nor UO_466 (O_466,N_48611,N_49470);
or UO_467 (O_467,N_48047,N_48670);
and UO_468 (O_468,N_49858,N_48561);
nand UO_469 (O_469,N_49685,N_49165);
or UO_470 (O_470,N_48572,N_49888);
nand UO_471 (O_471,N_48821,N_48043);
nor UO_472 (O_472,N_49591,N_48201);
xor UO_473 (O_473,N_48238,N_48873);
nor UO_474 (O_474,N_48300,N_49796);
xor UO_475 (O_475,N_48758,N_49753);
nand UO_476 (O_476,N_49231,N_49872);
nand UO_477 (O_477,N_49877,N_48658);
xnor UO_478 (O_478,N_48896,N_48747);
or UO_479 (O_479,N_49651,N_48637);
nor UO_480 (O_480,N_48068,N_48976);
or UO_481 (O_481,N_49252,N_49647);
and UO_482 (O_482,N_48624,N_48924);
nor UO_483 (O_483,N_48577,N_48357);
nand UO_484 (O_484,N_48377,N_49186);
and UO_485 (O_485,N_48569,N_49774);
nand UO_486 (O_486,N_48394,N_49688);
nand UO_487 (O_487,N_48636,N_49989);
nor UO_488 (O_488,N_49116,N_48610);
xnor UO_489 (O_489,N_49435,N_48109);
or UO_490 (O_490,N_48978,N_49713);
xor UO_491 (O_491,N_49851,N_49712);
or UO_492 (O_492,N_49643,N_49091);
nand UO_493 (O_493,N_49478,N_48191);
and UO_494 (O_494,N_48282,N_49747);
or UO_495 (O_495,N_48072,N_49025);
and UO_496 (O_496,N_48999,N_48699);
nor UO_497 (O_497,N_48596,N_49141);
and UO_498 (O_498,N_49609,N_49366);
or UO_499 (O_499,N_48981,N_48956);
nor UO_500 (O_500,N_49763,N_49472);
and UO_501 (O_501,N_49114,N_49087);
or UO_502 (O_502,N_49310,N_49862);
or UO_503 (O_503,N_48026,N_49889);
or UO_504 (O_504,N_49312,N_49229);
xnor UO_505 (O_505,N_48482,N_49035);
xor UO_506 (O_506,N_48199,N_48285);
or UO_507 (O_507,N_49240,N_48627);
or UO_508 (O_508,N_48661,N_48087);
or UO_509 (O_509,N_49584,N_49594);
and UO_510 (O_510,N_49171,N_49610);
and UO_511 (O_511,N_49043,N_48580);
xor UO_512 (O_512,N_48807,N_48586);
and UO_513 (O_513,N_49434,N_48920);
nand UO_514 (O_514,N_49315,N_48717);
nand UO_515 (O_515,N_49739,N_49313);
xnor UO_516 (O_516,N_48847,N_48543);
nand UO_517 (O_517,N_48816,N_48621);
or UO_518 (O_518,N_49736,N_49150);
xnor UO_519 (O_519,N_49937,N_49865);
xor UO_520 (O_520,N_48176,N_48163);
and UO_521 (O_521,N_49547,N_48824);
nor UO_522 (O_522,N_48575,N_49693);
and UO_523 (O_523,N_49567,N_48088);
or UO_524 (O_524,N_48531,N_49444);
nand UO_525 (O_525,N_48977,N_48448);
nor UO_526 (O_526,N_49866,N_48497);
nand UO_527 (O_527,N_49055,N_48171);
xor UO_528 (O_528,N_49597,N_49761);
xnor UO_529 (O_529,N_48761,N_49722);
and UO_530 (O_530,N_49202,N_49800);
nor UO_531 (O_531,N_48210,N_49057);
xor UO_532 (O_532,N_48375,N_48832);
xnor UO_533 (O_533,N_48781,N_48106);
nor UO_534 (O_534,N_48247,N_49829);
nor UO_535 (O_535,N_48213,N_49854);
xnor UO_536 (O_536,N_49504,N_49710);
nand UO_537 (O_537,N_49244,N_48331);
and UO_538 (O_538,N_48205,N_49445);
nor UO_539 (O_539,N_49166,N_48524);
or UO_540 (O_540,N_48617,N_49251);
and UO_541 (O_541,N_49193,N_49488);
nand UO_542 (O_542,N_49852,N_49505);
xor UO_543 (O_543,N_48302,N_49475);
nand UO_544 (O_544,N_49895,N_48031);
and UO_545 (O_545,N_48789,N_49894);
nor UO_546 (O_546,N_49992,N_49794);
nor UO_547 (O_547,N_48958,N_49744);
and UO_548 (O_548,N_49054,N_49881);
or UO_549 (O_549,N_49960,N_48277);
xor UO_550 (O_550,N_48702,N_48012);
and UO_551 (O_551,N_48680,N_48775);
nand UO_552 (O_552,N_48042,N_49941);
xnor UO_553 (O_553,N_48105,N_48745);
nand UO_554 (O_554,N_49533,N_48311);
nor UO_555 (O_555,N_48737,N_49694);
or UO_556 (O_556,N_48274,N_49600);
nor UO_557 (O_557,N_48468,N_49145);
nand UO_558 (O_558,N_48165,N_48545);
nand UO_559 (O_559,N_49253,N_49357);
or UO_560 (O_560,N_48907,N_49115);
nand UO_561 (O_561,N_49783,N_49535);
nand UO_562 (O_562,N_49005,N_48633);
xnor UO_563 (O_563,N_49979,N_49139);
nand UO_564 (O_564,N_48057,N_48436);
and UO_565 (O_565,N_48714,N_48093);
or UO_566 (O_566,N_49195,N_48547);
xnor UO_567 (O_567,N_48214,N_48876);
xnor UO_568 (O_568,N_49429,N_48490);
and UO_569 (O_569,N_49639,N_48298);
nand UO_570 (O_570,N_49838,N_49550);
nor UO_571 (O_571,N_49080,N_49164);
or UO_572 (O_572,N_48992,N_49259);
nor UO_573 (O_573,N_48148,N_49534);
or UO_574 (O_574,N_48209,N_49301);
and UO_575 (O_575,N_49545,N_48050);
or UO_576 (O_576,N_49185,N_49044);
or UO_577 (O_577,N_48692,N_48194);
nor UO_578 (O_578,N_48424,N_49017);
or UO_579 (O_579,N_49990,N_48359);
and UO_580 (O_580,N_48672,N_49581);
and UO_581 (O_581,N_48239,N_48830);
or UO_582 (O_582,N_49997,N_49883);
or UO_583 (O_583,N_49189,N_49417);
or UO_584 (O_584,N_49608,N_48384);
or UO_585 (O_585,N_48583,N_48837);
or UO_586 (O_586,N_48609,N_49906);
or UO_587 (O_587,N_48612,N_48067);
xor UO_588 (O_588,N_48712,N_49706);
xnor UO_589 (O_589,N_49705,N_48306);
or UO_590 (O_590,N_48414,N_48217);
xor UO_591 (O_591,N_48477,N_49084);
nand UO_592 (O_592,N_48425,N_49808);
nor UO_593 (O_593,N_48196,N_48023);
and UO_594 (O_594,N_49799,N_48166);
or UO_595 (O_595,N_49537,N_48153);
and UO_596 (O_596,N_49449,N_48537);
xnor UO_597 (O_597,N_48643,N_48653);
or UO_598 (O_598,N_49354,N_49944);
and UO_599 (O_599,N_49648,N_48097);
nand UO_600 (O_600,N_48389,N_48233);
xor UO_601 (O_601,N_48558,N_49316);
and UO_602 (O_602,N_49437,N_48450);
and UO_603 (O_603,N_49611,N_49329);
xor UO_604 (O_604,N_48065,N_49097);
and UO_605 (O_605,N_49023,N_48077);
or UO_606 (O_606,N_48143,N_48913);
or UO_607 (O_607,N_49129,N_49291);
and UO_608 (O_608,N_48190,N_49658);
and UO_609 (O_609,N_49801,N_49667);
xnor UO_610 (O_610,N_48722,N_49936);
and UO_611 (O_611,N_48603,N_49711);
nor UO_612 (O_612,N_49964,N_48616);
nand UO_613 (O_613,N_49191,N_48987);
nor UO_614 (O_614,N_49319,N_48241);
and UO_615 (O_615,N_49209,N_48324);
nand UO_616 (O_616,N_48256,N_48269);
xnor UO_617 (O_617,N_49598,N_49701);
nand UO_618 (O_618,N_48061,N_48953);
and UO_619 (O_619,N_49679,N_48951);
and UO_620 (O_620,N_49742,N_49134);
nand UO_621 (O_621,N_49383,N_48351);
xor UO_622 (O_622,N_49576,N_49632);
and UO_623 (O_623,N_48086,N_48348);
or UO_624 (O_624,N_48752,N_48276);
nand UO_625 (O_625,N_49331,N_48831);
nor UO_626 (O_626,N_49351,N_48989);
or UO_627 (O_627,N_48619,N_49921);
nor UO_628 (O_628,N_48466,N_49522);
nor UO_629 (O_629,N_49748,N_48008);
or UO_630 (O_630,N_48118,N_48013);
and UO_631 (O_631,N_49559,N_48869);
nor UO_632 (O_632,N_49557,N_48937);
nand UO_633 (O_633,N_49039,N_49743);
xnor UO_634 (O_634,N_49572,N_48040);
nor UO_635 (O_635,N_49153,N_48595);
or UO_636 (O_636,N_48529,N_49111);
nor UO_637 (O_637,N_49323,N_48800);
nor UO_638 (O_638,N_48368,N_48332);
or UO_639 (O_639,N_48338,N_49822);
and UO_640 (O_640,N_48251,N_48845);
nand UO_641 (O_641,N_49052,N_49161);
xnor UO_642 (O_642,N_48703,N_48523);
and UO_643 (O_643,N_48705,N_48498);
xnor UO_644 (O_644,N_48009,N_49751);
or UO_645 (O_645,N_49917,N_48342);
and UO_646 (O_646,N_48314,N_48452);
and UO_647 (O_647,N_48819,N_48168);
or UO_648 (O_648,N_49474,N_48249);
nand UO_649 (O_649,N_49456,N_49515);
and UO_650 (O_650,N_49350,N_49395);
xnor UO_651 (O_651,N_48301,N_49495);
and UO_652 (O_652,N_48278,N_49008);
nand UO_653 (O_653,N_48792,N_49867);
and UO_654 (O_654,N_49406,N_48391);
nand UO_655 (O_655,N_49813,N_49408);
or UO_656 (O_656,N_48367,N_49398);
nand UO_657 (O_657,N_49791,N_48296);
nor UO_658 (O_658,N_48323,N_48961);
and UO_659 (O_659,N_48844,N_49072);
and UO_660 (O_660,N_48037,N_49197);
nand UO_661 (O_661,N_49073,N_49413);
or UO_662 (O_662,N_48193,N_48366);
or UO_663 (O_663,N_49525,N_48119);
and UO_664 (O_664,N_48417,N_49770);
or UO_665 (O_665,N_48839,N_49915);
and UO_666 (O_666,N_49766,N_48676);
or UO_667 (O_667,N_49521,N_48155);
xnor UO_668 (O_668,N_49661,N_48271);
or UO_669 (O_669,N_48590,N_48052);
and UO_670 (O_670,N_49003,N_49212);
nand UO_671 (O_671,N_48126,N_48791);
or UO_672 (O_672,N_48449,N_49230);
xnor UO_673 (O_673,N_49665,N_49140);
or UO_674 (O_674,N_48553,N_48795);
nand UO_675 (O_675,N_49955,N_48175);
xor UO_676 (O_676,N_49677,N_49564);
nand UO_677 (O_677,N_48312,N_49657);
xor UO_678 (O_678,N_48784,N_48500);
or UO_679 (O_679,N_48138,N_49678);
or UO_680 (O_680,N_49220,N_49371);
nor UO_681 (O_681,N_48689,N_49090);
and UO_682 (O_682,N_49460,N_49691);
and UO_683 (O_683,N_49415,N_48255);
nand UO_684 (O_684,N_49267,N_48147);
nand UO_685 (O_685,N_48402,N_49455);
and UO_686 (O_686,N_48855,N_49893);
xnor UO_687 (O_687,N_48823,N_49724);
xor UO_688 (O_688,N_48726,N_48472);
xnor UO_689 (O_689,N_49359,N_49027);
or UO_690 (O_690,N_49561,N_48258);
or UO_691 (O_691,N_49715,N_49869);
xnor UO_692 (O_692,N_48748,N_49914);
nand UO_693 (O_693,N_49225,N_48024);
xnor UO_694 (O_694,N_49918,N_49741);
or UO_695 (O_695,N_48740,N_49213);
nor UO_696 (O_696,N_49779,N_49334);
xor UO_697 (O_697,N_49174,N_49412);
or UO_698 (O_698,N_48094,N_49717);
nor UO_699 (O_699,N_49071,N_49887);
xor UO_700 (O_700,N_49539,N_48889);
and UO_701 (O_701,N_48849,N_48423);
nand UO_702 (O_702,N_48079,N_48473);
nor UO_703 (O_703,N_48949,N_48751);
and UO_704 (O_704,N_48871,N_49309);
and UO_705 (O_705,N_49552,N_49583);
and UO_706 (O_706,N_48794,N_49910);
and UO_707 (O_707,N_48177,N_49059);
nand UO_708 (O_708,N_48805,N_48262);
nor UO_709 (O_709,N_48104,N_48470);
xor UO_710 (O_710,N_48985,N_49284);
nor UO_711 (O_711,N_49874,N_48427);
or UO_712 (O_712,N_48140,N_48762);
and UO_713 (O_713,N_49795,N_48297);
or UO_714 (O_714,N_49457,N_48944);
or UO_715 (O_715,N_48584,N_48693);
nor UO_716 (O_716,N_49898,N_49200);
xor UO_717 (O_717,N_49183,N_49010);
nand UO_718 (O_718,N_49945,N_48284);
and UO_719 (O_719,N_48288,N_49287);
xnor UO_720 (O_720,N_48683,N_49133);
or UO_721 (O_721,N_48303,N_48499);
nand UO_722 (O_722,N_48891,N_49420);
nor UO_723 (O_723,N_49575,N_49405);
nand UO_724 (O_724,N_49311,N_49871);
nand UO_725 (O_725,N_48471,N_49592);
nor UO_726 (O_726,N_48051,N_48434);
and UO_727 (O_727,N_48488,N_49996);
nand UO_728 (O_728,N_49957,N_48381);
and UO_729 (O_729,N_48220,N_49032);
nand UO_730 (O_730,N_49824,N_49698);
xnor UO_731 (O_731,N_49855,N_49788);
or UO_732 (O_732,N_48948,N_49491);
xor UO_733 (O_733,N_49853,N_49175);
nand UO_734 (O_734,N_48044,N_49580);
or UO_735 (O_735,N_49920,N_48727);
nor UO_736 (O_736,N_49764,N_49053);
nor UO_737 (O_737,N_49423,N_49298);
xor UO_738 (O_738,N_48413,N_48858);
or UO_739 (O_739,N_48096,N_49452);
xnor UO_740 (O_740,N_49837,N_48922);
nor UO_741 (O_741,N_48986,N_48460);
and UO_742 (O_742,N_48813,N_48530);
and UO_743 (O_743,N_48615,N_48203);
or UO_744 (O_744,N_49328,N_49454);
or UO_745 (O_745,N_49426,N_48725);
or UO_746 (O_746,N_48275,N_48657);
or UO_747 (O_747,N_48159,N_49511);
xnor UO_748 (O_748,N_49172,N_49804);
nor UO_749 (O_749,N_49394,N_48192);
nand UO_750 (O_750,N_49158,N_49431);
or UO_751 (O_751,N_49771,N_48629);
or UO_752 (O_752,N_49199,N_48542);
or UO_753 (O_753,N_49340,N_49879);
xor UO_754 (O_754,N_49377,N_49249);
nor UO_755 (O_755,N_49606,N_48738);
and UO_756 (O_756,N_48602,N_49233);
nor UO_757 (O_757,N_49950,N_49446);
and UO_758 (O_758,N_49821,N_48646);
or UO_759 (O_759,N_49217,N_48260);
xnor UO_760 (O_760,N_49927,N_48656);
xnor UO_761 (O_761,N_49507,N_49138);
or UO_762 (O_762,N_49342,N_49009);
nor UO_763 (O_763,N_49928,N_48385);
and UO_764 (O_764,N_48169,N_48650);
or UO_765 (O_765,N_48549,N_48149);
or UO_766 (O_766,N_48294,N_49493);
nand UO_767 (O_767,N_48003,N_48681);
nor UO_768 (O_768,N_48139,N_49692);
and UO_769 (O_769,N_48019,N_49154);
and UO_770 (O_770,N_49578,N_49248);
or UO_771 (O_771,N_48834,N_48492);
and UO_772 (O_772,N_49402,N_48613);
or UO_773 (O_773,N_49326,N_48010);
nand UO_774 (O_774,N_48928,N_49911);
nand UO_775 (O_775,N_48903,N_49527);
or UO_776 (O_776,N_49425,N_48197);
and UO_777 (O_777,N_49556,N_48407);
xor UO_778 (O_778,N_48753,N_48173);
and UO_779 (O_779,N_49933,N_48422);
nor UO_780 (O_780,N_48070,N_49690);
or UO_781 (O_781,N_49203,N_49011);
xor UO_782 (O_782,N_49884,N_49228);
or UO_783 (O_783,N_48388,N_49585);
nor UO_784 (O_784,N_49242,N_49605);
nor UO_785 (O_785,N_48945,N_48502);
or UO_786 (O_786,N_48836,N_48801);
nor UO_787 (O_787,N_49762,N_48137);
nor UO_788 (O_788,N_49707,N_48457);
nand UO_789 (O_789,N_49304,N_49590);
and UO_790 (O_790,N_48287,N_48403);
or UO_791 (O_791,N_48185,N_48783);
nand UO_792 (O_792,N_48888,N_48286);
and UO_793 (O_793,N_48189,N_48246);
nor UO_794 (O_794,N_48089,N_48716);
nand UO_795 (O_795,N_49428,N_48172);
nand UO_796 (O_796,N_49540,N_48620);
nand UO_797 (O_797,N_49264,N_49653);
xnor UO_798 (O_798,N_48103,N_49603);
xor UO_799 (O_799,N_48128,N_49056);
and UO_800 (O_800,N_48272,N_49355);
nor UO_801 (O_801,N_48223,N_48597);
nand UO_802 (O_802,N_48150,N_48133);
and UO_803 (O_803,N_49579,N_48967);
xnor UO_804 (O_804,N_48820,N_49380);
and UO_805 (O_805,N_49409,N_48898);
and UO_806 (O_806,N_48283,N_48440);
xor UO_807 (O_807,N_48259,N_48917);
and UO_808 (O_808,N_48517,N_49702);
nand UO_809 (O_809,N_48648,N_49868);
and UO_810 (O_810,N_48350,N_48965);
and UO_811 (O_811,N_48392,N_49358);
or UO_812 (O_812,N_49061,N_48001);
and UO_813 (O_813,N_48503,N_49988);
nand UO_814 (O_814,N_48328,N_48231);
nor UO_815 (O_815,N_49892,N_48157);
nand UO_816 (O_816,N_49708,N_48124);
nor UO_817 (O_817,N_49954,N_48343);
nor UO_818 (O_818,N_49400,N_48719);
xnor UO_819 (O_819,N_48006,N_49726);
or UO_820 (O_820,N_49045,N_49846);
nor UO_821 (O_821,N_48766,N_48337);
and UO_822 (O_822,N_49349,N_49484);
and UO_823 (O_823,N_48776,N_49769);
or UO_824 (O_824,N_48744,N_48533);
or UO_825 (O_825,N_49275,N_48827);
nor UO_826 (O_826,N_49469,N_49033);
or UO_827 (O_827,N_48536,N_48541);
xor UO_828 (O_828,N_48410,N_48697);
xnor UO_829 (O_829,N_48380,N_48446);
or UO_830 (O_830,N_48131,N_48786);
or UO_831 (O_831,N_49519,N_48682);
nand UO_832 (O_832,N_48349,N_49746);
xnor UO_833 (O_833,N_49959,N_48054);
or UO_834 (O_834,N_48111,N_49341);
nand UO_835 (O_835,N_48966,N_48374);
and UO_836 (O_836,N_48495,N_48565);
or UO_837 (O_837,N_48591,N_49276);
and UO_838 (O_838,N_48066,N_49486);
xnor UO_839 (O_839,N_48229,N_49940);
and UO_840 (O_840,N_48511,N_48861);
and UO_841 (O_841,N_49833,N_49931);
nand UO_842 (O_842,N_48885,N_48867);
nand UO_843 (O_843,N_48081,N_48769);
nand UO_844 (O_844,N_49451,N_49019);
nand UO_845 (O_845,N_49169,N_49265);
and UO_846 (O_846,N_48083,N_49873);
and UO_847 (O_847,N_49384,N_48706);
nor UO_848 (O_848,N_48307,N_48000);
xor UO_849 (O_849,N_49067,N_48053);
or UO_850 (O_850,N_49577,N_48774);
nand UO_851 (O_851,N_48095,N_49637);
and UO_852 (O_852,N_49859,N_48995);
and UO_853 (O_853,N_48647,N_49333);
xor UO_854 (O_854,N_49143,N_48064);
xnor UO_855 (O_855,N_49614,N_48090);
xor UO_856 (O_856,N_49756,N_49238);
xnor UO_857 (O_857,N_49662,N_48279);
nor UO_858 (O_858,N_49269,N_48506);
or UO_859 (O_859,N_49613,N_48778);
nor UO_860 (O_860,N_49461,N_49254);
and UO_861 (O_861,N_49148,N_49268);
and UO_862 (O_862,N_49407,N_48797);
or UO_863 (O_863,N_49223,N_49300);
nand UO_864 (O_864,N_49439,N_49216);
nor UO_865 (O_865,N_48489,N_49322);
nor UO_866 (O_866,N_48483,N_48763);
and UO_867 (O_867,N_48578,N_49363);
xor UO_868 (O_868,N_49482,N_49404);
and UO_869 (O_869,N_48011,N_48304);
nor UO_870 (O_870,N_49671,N_49187);
xor UO_871 (O_871,N_49277,N_49699);
and UO_872 (O_872,N_48516,N_48566);
or UO_873 (O_873,N_49582,N_48817);
xnor UO_874 (O_874,N_48592,N_49490);
nor UO_875 (O_875,N_48445,N_48640);
nand UO_876 (O_876,N_48114,N_48250);
or UO_877 (O_877,N_48478,N_48790);
xor UO_878 (O_878,N_49948,N_49221);
or UO_879 (O_879,N_49555,N_48320);
and UO_880 (O_880,N_49332,N_49650);
nand UO_881 (O_881,N_48887,N_49327);
and UO_882 (O_882,N_48002,N_49020);
and UO_883 (O_883,N_49759,N_48535);
nand UO_884 (O_884,N_48463,N_49146);
nand UO_885 (O_885,N_48322,N_48221);
and UO_886 (O_886,N_49811,N_49081);
nor UO_887 (O_887,N_48454,N_48370);
nand UO_888 (O_888,N_48063,N_49857);
nor UO_889 (O_889,N_48691,N_49477);
nand UO_890 (O_890,N_49782,N_48734);
or UO_891 (O_891,N_48038,N_49785);
and UO_892 (O_892,N_49226,N_48796);
nor UO_893 (O_893,N_49750,N_49844);
and UO_894 (O_894,N_48412,N_49737);
nand UO_895 (O_895,N_49182,N_49730);
or UO_896 (O_896,N_48305,N_48632);
or UO_897 (O_897,N_49137,N_49994);
or UO_898 (O_898,N_49672,N_49777);
or UO_899 (O_899,N_48777,N_48663);
nand UO_900 (O_900,N_49775,N_49427);
nand UO_901 (O_901,N_48518,N_48593);
xor UO_902 (O_902,N_48866,N_48687);
nand UO_903 (O_903,N_48833,N_49725);
nand UO_904 (O_904,N_48654,N_48843);
or UO_905 (O_905,N_49956,N_49735);
nor UO_906 (O_906,N_48188,N_48771);
or UO_907 (O_907,N_49278,N_48475);
or UO_908 (O_908,N_48974,N_49659);
and UO_909 (O_909,N_48564,N_49101);
nand UO_910 (O_910,N_48660,N_49147);
xnor UO_911 (O_911,N_49962,N_49727);
xor UO_912 (O_912,N_49299,N_49250);
or UO_913 (O_913,N_48353,N_49680);
nor UO_914 (O_914,N_49830,N_48933);
nor UO_915 (O_915,N_48174,N_48875);
and UO_916 (O_916,N_49125,N_48906);
or UO_917 (O_917,N_48788,N_49204);
or UO_918 (O_918,N_48905,N_48134);
xnor UO_919 (O_919,N_48318,N_49513);
xor UO_920 (O_920,N_49438,N_49256);
or UO_921 (O_921,N_49891,N_49574);
nor UO_922 (O_922,N_48842,N_49885);
nand UO_923 (O_923,N_48526,N_48404);
nand UO_924 (O_924,N_49728,N_48020);
and UO_925 (O_925,N_48655,N_49618);
or UO_926 (O_926,N_48785,N_48224);
or UO_927 (O_927,N_48345,N_48491);
and UO_928 (O_928,N_48668,N_49589);
nor UO_929 (O_929,N_49335,N_49644);
nor UO_930 (O_930,N_48990,N_49615);
nand UO_931 (O_931,N_48736,N_48364);
xor UO_932 (O_932,N_48856,N_49018);
and UO_933 (O_933,N_48598,N_49156);
nor UO_934 (O_934,N_48376,N_49586);
or UO_935 (O_935,N_48481,N_48878);
nor UO_936 (O_936,N_49809,N_48688);
nor UO_937 (O_937,N_49983,N_49330);
xor UO_938 (O_938,N_49716,N_48971);
xor UO_939 (O_939,N_48701,N_49205);
nand UO_940 (O_940,N_48684,N_48142);
or UO_941 (O_941,N_48941,N_49386);
nand UO_942 (O_942,N_49038,N_48334);
nor UO_943 (O_943,N_49916,N_48069);
xor UO_944 (O_944,N_49806,N_48202);
or UO_945 (O_945,N_48814,N_49476);
and UO_946 (O_946,N_48863,N_49336);
nor UO_947 (O_947,N_49731,N_49970);
nor UO_948 (O_948,N_49215,N_48395);
and UO_949 (O_949,N_49878,N_48273);
nand UO_950 (O_950,N_49798,N_49286);
and UO_951 (O_951,N_48880,N_48544);
nand UO_952 (O_952,N_49118,N_48787);
xnor UO_953 (O_953,N_48594,N_49772);
nor UO_954 (O_954,N_49827,N_48929);
xnor UO_955 (O_955,N_49520,N_48810);
or UO_956 (O_956,N_49740,N_48690);
nand UO_957 (O_957,N_49904,N_48170);
nand UO_958 (O_958,N_48336,N_49570);
nand UO_959 (O_959,N_48129,N_48841);
and UO_960 (O_960,N_48532,N_48571);
xor UO_961 (O_961,N_48581,N_48340);
nor UO_962 (O_962,N_49760,N_48614);
nor UO_963 (O_963,N_48494,N_48018);
nor UO_964 (O_964,N_48266,N_48548);
xor UO_965 (O_965,N_49029,N_48493);
or UO_966 (O_966,N_48162,N_48430);
nor UO_967 (O_967,N_49842,N_48411);
nand UO_968 (O_968,N_49602,N_48060);
xnor UO_969 (O_969,N_48879,N_49549);
nor UO_970 (O_970,N_49448,N_48099);
xnor UO_971 (O_971,N_49875,N_48232);
or UO_972 (O_972,N_48520,N_49450);
nor UO_973 (O_973,N_49946,N_49820);
and UO_974 (O_974,N_48442,N_48313);
nor UO_975 (O_975,N_49176,N_48988);
nand UO_976 (O_976,N_49674,N_49178);
nor UO_977 (O_977,N_48918,N_48666);
xnor UO_978 (O_978,N_49321,N_49792);
or UO_979 (O_979,N_48854,N_48074);
or UO_980 (O_980,N_49048,N_49684);
or UO_981 (O_981,N_49636,N_49656);
nor UO_982 (O_982,N_49179,N_49718);
nor UO_983 (O_983,N_48730,N_49466);
xnor UO_984 (O_984,N_49124,N_49633);
nand UO_985 (O_985,N_48731,N_48835);
xor UO_986 (O_986,N_48892,N_49551);
or UO_987 (O_987,N_48939,N_49621);
and UO_988 (O_988,N_48028,N_48317);
nand UO_989 (O_989,N_48206,N_48728);
and UO_990 (O_990,N_49103,N_49014);
and UO_991 (O_991,N_48960,N_49297);
or UO_992 (O_992,N_49198,N_49393);
nand UO_993 (O_993,N_49136,N_48058);
or UO_994 (O_994,N_48228,N_48041);
xnor UO_995 (O_995,N_49356,N_49219);
nor UO_996 (O_996,N_48476,N_48076);
or UO_997 (O_997,N_49094,N_49180);
xnor UO_998 (O_998,N_48245,N_48926);
or UO_999 (O_999,N_48674,N_48501);
and UO_1000 (O_1000,N_49291,N_49105);
xnor UO_1001 (O_1001,N_49127,N_49504);
and UO_1002 (O_1002,N_49099,N_48868);
nand UO_1003 (O_1003,N_48034,N_49463);
or UO_1004 (O_1004,N_48037,N_48199);
nor UO_1005 (O_1005,N_49132,N_48733);
xnor UO_1006 (O_1006,N_49514,N_48888);
nor UO_1007 (O_1007,N_49173,N_48105);
and UO_1008 (O_1008,N_48170,N_49835);
xor UO_1009 (O_1009,N_48489,N_49401);
nand UO_1010 (O_1010,N_49417,N_49029);
nor UO_1011 (O_1011,N_48043,N_48199);
and UO_1012 (O_1012,N_49175,N_49187);
xnor UO_1013 (O_1013,N_49243,N_48101);
nand UO_1014 (O_1014,N_49785,N_48715);
and UO_1015 (O_1015,N_48364,N_48901);
and UO_1016 (O_1016,N_49309,N_49840);
and UO_1017 (O_1017,N_48576,N_49918);
xnor UO_1018 (O_1018,N_49997,N_48061);
or UO_1019 (O_1019,N_48294,N_48643);
and UO_1020 (O_1020,N_49866,N_49234);
or UO_1021 (O_1021,N_49174,N_49630);
nor UO_1022 (O_1022,N_48422,N_48963);
or UO_1023 (O_1023,N_48932,N_48209);
nand UO_1024 (O_1024,N_49510,N_49426);
xnor UO_1025 (O_1025,N_49235,N_49118);
xor UO_1026 (O_1026,N_48876,N_49924);
xnor UO_1027 (O_1027,N_48747,N_48255);
nand UO_1028 (O_1028,N_48136,N_49892);
xnor UO_1029 (O_1029,N_48815,N_48460);
nor UO_1030 (O_1030,N_48677,N_48653);
xnor UO_1031 (O_1031,N_49944,N_48000);
nor UO_1032 (O_1032,N_49230,N_48363);
xor UO_1033 (O_1033,N_48365,N_49809);
or UO_1034 (O_1034,N_49599,N_48206);
or UO_1035 (O_1035,N_48749,N_48186);
and UO_1036 (O_1036,N_48483,N_49820);
nor UO_1037 (O_1037,N_48322,N_48497);
nand UO_1038 (O_1038,N_49299,N_48885);
nor UO_1039 (O_1039,N_48987,N_49897);
and UO_1040 (O_1040,N_48285,N_49014);
nor UO_1041 (O_1041,N_48210,N_48743);
nor UO_1042 (O_1042,N_48863,N_48726);
or UO_1043 (O_1043,N_48565,N_49599);
nor UO_1044 (O_1044,N_49257,N_48779);
nor UO_1045 (O_1045,N_48964,N_48032);
and UO_1046 (O_1046,N_49143,N_49908);
or UO_1047 (O_1047,N_48853,N_49302);
or UO_1048 (O_1048,N_48044,N_49099);
nor UO_1049 (O_1049,N_49456,N_49399);
nand UO_1050 (O_1050,N_48855,N_49223);
or UO_1051 (O_1051,N_49301,N_48203);
xnor UO_1052 (O_1052,N_48002,N_48042);
nor UO_1053 (O_1053,N_49192,N_48227);
and UO_1054 (O_1054,N_48650,N_49370);
or UO_1055 (O_1055,N_48191,N_48955);
and UO_1056 (O_1056,N_49427,N_48053);
nor UO_1057 (O_1057,N_48700,N_48090);
nor UO_1058 (O_1058,N_49834,N_49658);
xor UO_1059 (O_1059,N_48172,N_49954);
xor UO_1060 (O_1060,N_48769,N_49594);
and UO_1061 (O_1061,N_48471,N_48322);
nand UO_1062 (O_1062,N_48854,N_49199);
nor UO_1063 (O_1063,N_48344,N_49890);
nand UO_1064 (O_1064,N_49502,N_49037);
nand UO_1065 (O_1065,N_49781,N_49267);
or UO_1066 (O_1066,N_48001,N_49084);
nand UO_1067 (O_1067,N_49680,N_49279);
xor UO_1068 (O_1068,N_49570,N_49274);
xnor UO_1069 (O_1069,N_49507,N_49633);
nor UO_1070 (O_1070,N_48826,N_48607);
xor UO_1071 (O_1071,N_48138,N_48143);
nand UO_1072 (O_1072,N_49521,N_48008);
or UO_1073 (O_1073,N_49580,N_48479);
xnor UO_1074 (O_1074,N_48530,N_48328);
or UO_1075 (O_1075,N_49278,N_49169);
nor UO_1076 (O_1076,N_49648,N_48956);
nor UO_1077 (O_1077,N_48899,N_49663);
and UO_1078 (O_1078,N_48314,N_48072);
xnor UO_1079 (O_1079,N_49355,N_49710);
xnor UO_1080 (O_1080,N_48469,N_48823);
nand UO_1081 (O_1081,N_48937,N_48691);
and UO_1082 (O_1082,N_48473,N_48456);
nand UO_1083 (O_1083,N_48898,N_49829);
nor UO_1084 (O_1084,N_49508,N_48590);
or UO_1085 (O_1085,N_48230,N_48217);
and UO_1086 (O_1086,N_48932,N_48900);
or UO_1087 (O_1087,N_48564,N_49749);
nand UO_1088 (O_1088,N_48038,N_48601);
xnor UO_1089 (O_1089,N_48923,N_49851);
and UO_1090 (O_1090,N_49710,N_48982);
xor UO_1091 (O_1091,N_49814,N_48398);
or UO_1092 (O_1092,N_49543,N_48525);
nor UO_1093 (O_1093,N_48540,N_49509);
nand UO_1094 (O_1094,N_49843,N_48937);
nor UO_1095 (O_1095,N_49702,N_49069);
or UO_1096 (O_1096,N_49420,N_49754);
nor UO_1097 (O_1097,N_49665,N_49777);
or UO_1098 (O_1098,N_48377,N_49680);
xor UO_1099 (O_1099,N_48563,N_48772);
xor UO_1100 (O_1100,N_49040,N_49465);
nor UO_1101 (O_1101,N_48613,N_48926);
and UO_1102 (O_1102,N_49428,N_49375);
nand UO_1103 (O_1103,N_48436,N_48969);
nor UO_1104 (O_1104,N_48025,N_48769);
nor UO_1105 (O_1105,N_49128,N_49668);
nand UO_1106 (O_1106,N_49780,N_49675);
or UO_1107 (O_1107,N_48793,N_48164);
and UO_1108 (O_1108,N_48398,N_48103);
xor UO_1109 (O_1109,N_49747,N_48492);
xnor UO_1110 (O_1110,N_49609,N_49407);
and UO_1111 (O_1111,N_49202,N_48541);
nor UO_1112 (O_1112,N_48027,N_48249);
and UO_1113 (O_1113,N_49417,N_48793);
or UO_1114 (O_1114,N_48117,N_49382);
xnor UO_1115 (O_1115,N_49378,N_49568);
nor UO_1116 (O_1116,N_48221,N_49871);
xnor UO_1117 (O_1117,N_48860,N_49315);
and UO_1118 (O_1118,N_48900,N_49704);
nor UO_1119 (O_1119,N_48573,N_48235);
nor UO_1120 (O_1120,N_48218,N_49305);
and UO_1121 (O_1121,N_49651,N_49196);
xor UO_1122 (O_1122,N_49767,N_49517);
or UO_1123 (O_1123,N_49292,N_49037);
nand UO_1124 (O_1124,N_49178,N_49018);
xor UO_1125 (O_1125,N_49017,N_49041);
nand UO_1126 (O_1126,N_48872,N_49185);
xnor UO_1127 (O_1127,N_49872,N_48347);
nand UO_1128 (O_1128,N_49499,N_48556);
and UO_1129 (O_1129,N_49990,N_48037);
xor UO_1130 (O_1130,N_48217,N_48447);
xnor UO_1131 (O_1131,N_49147,N_48890);
or UO_1132 (O_1132,N_49606,N_49956);
and UO_1133 (O_1133,N_49273,N_48725);
or UO_1134 (O_1134,N_49458,N_48012);
nor UO_1135 (O_1135,N_49204,N_48863);
xor UO_1136 (O_1136,N_48358,N_48318);
nor UO_1137 (O_1137,N_49380,N_49133);
nand UO_1138 (O_1138,N_49258,N_49657);
and UO_1139 (O_1139,N_48871,N_48178);
nor UO_1140 (O_1140,N_48277,N_48410);
or UO_1141 (O_1141,N_49935,N_49598);
xor UO_1142 (O_1142,N_49173,N_49175);
and UO_1143 (O_1143,N_49023,N_49359);
nand UO_1144 (O_1144,N_49915,N_49162);
or UO_1145 (O_1145,N_49712,N_48322);
or UO_1146 (O_1146,N_49448,N_48888);
nor UO_1147 (O_1147,N_48990,N_48722);
and UO_1148 (O_1148,N_49556,N_48062);
nand UO_1149 (O_1149,N_48527,N_48661);
nand UO_1150 (O_1150,N_48588,N_48565);
nor UO_1151 (O_1151,N_48679,N_48182);
nand UO_1152 (O_1152,N_48403,N_48981);
xnor UO_1153 (O_1153,N_48266,N_49563);
nor UO_1154 (O_1154,N_48526,N_48741);
nand UO_1155 (O_1155,N_48563,N_49922);
nand UO_1156 (O_1156,N_49756,N_49510);
or UO_1157 (O_1157,N_48346,N_48955);
nand UO_1158 (O_1158,N_48086,N_48101);
xor UO_1159 (O_1159,N_49420,N_48892);
and UO_1160 (O_1160,N_49926,N_49049);
xor UO_1161 (O_1161,N_48000,N_49008);
xnor UO_1162 (O_1162,N_49067,N_49470);
nand UO_1163 (O_1163,N_48817,N_49781);
and UO_1164 (O_1164,N_48662,N_48164);
or UO_1165 (O_1165,N_49028,N_48544);
nor UO_1166 (O_1166,N_49191,N_48486);
nor UO_1167 (O_1167,N_48328,N_49951);
or UO_1168 (O_1168,N_49398,N_48818);
nor UO_1169 (O_1169,N_49105,N_49985);
or UO_1170 (O_1170,N_48908,N_48101);
and UO_1171 (O_1171,N_48743,N_49483);
nand UO_1172 (O_1172,N_48307,N_48220);
xor UO_1173 (O_1173,N_49581,N_49216);
nor UO_1174 (O_1174,N_49969,N_48874);
and UO_1175 (O_1175,N_48754,N_49357);
nor UO_1176 (O_1176,N_49205,N_49178);
and UO_1177 (O_1177,N_49858,N_48860);
nand UO_1178 (O_1178,N_49911,N_48149);
nor UO_1179 (O_1179,N_48394,N_49527);
or UO_1180 (O_1180,N_48537,N_48493);
or UO_1181 (O_1181,N_48745,N_49148);
and UO_1182 (O_1182,N_48489,N_48560);
or UO_1183 (O_1183,N_49261,N_48782);
nor UO_1184 (O_1184,N_49521,N_48588);
or UO_1185 (O_1185,N_49679,N_49097);
and UO_1186 (O_1186,N_49110,N_49874);
nor UO_1187 (O_1187,N_48507,N_49951);
nand UO_1188 (O_1188,N_48601,N_49412);
nor UO_1189 (O_1189,N_48552,N_49945);
and UO_1190 (O_1190,N_48182,N_49803);
nor UO_1191 (O_1191,N_49032,N_48526);
or UO_1192 (O_1192,N_48203,N_49497);
nor UO_1193 (O_1193,N_48835,N_49761);
nor UO_1194 (O_1194,N_49993,N_48629);
and UO_1195 (O_1195,N_49323,N_49866);
nor UO_1196 (O_1196,N_48336,N_48130);
or UO_1197 (O_1197,N_48289,N_49512);
and UO_1198 (O_1198,N_48271,N_49724);
and UO_1199 (O_1199,N_49924,N_49810);
nor UO_1200 (O_1200,N_49412,N_49217);
and UO_1201 (O_1201,N_48778,N_49785);
nand UO_1202 (O_1202,N_49988,N_48241);
nand UO_1203 (O_1203,N_48531,N_49307);
nor UO_1204 (O_1204,N_48375,N_48622);
nand UO_1205 (O_1205,N_48154,N_48631);
xor UO_1206 (O_1206,N_49870,N_48145);
or UO_1207 (O_1207,N_48412,N_49666);
nand UO_1208 (O_1208,N_48857,N_49750);
and UO_1209 (O_1209,N_49635,N_49277);
xnor UO_1210 (O_1210,N_49930,N_48786);
and UO_1211 (O_1211,N_48832,N_49656);
xor UO_1212 (O_1212,N_49149,N_48914);
nand UO_1213 (O_1213,N_48453,N_48327);
nand UO_1214 (O_1214,N_49553,N_48669);
xor UO_1215 (O_1215,N_49129,N_48391);
nor UO_1216 (O_1216,N_48769,N_49863);
xor UO_1217 (O_1217,N_49358,N_48045);
xnor UO_1218 (O_1218,N_48771,N_48318);
or UO_1219 (O_1219,N_49428,N_49802);
nor UO_1220 (O_1220,N_49008,N_48578);
or UO_1221 (O_1221,N_49438,N_49506);
xor UO_1222 (O_1222,N_49701,N_49510);
nand UO_1223 (O_1223,N_48872,N_48340);
nor UO_1224 (O_1224,N_49734,N_48630);
nor UO_1225 (O_1225,N_48714,N_48633);
or UO_1226 (O_1226,N_48948,N_48743);
nor UO_1227 (O_1227,N_49373,N_48317);
and UO_1228 (O_1228,N_49736,N_48338);
nand UO_1229 (O_1229,N_49790,N_48262);
or UO_1230 (O_1230,N_48484,N_48576);
xor UO_1231 (O_1231,N_48141,N_49809);
and UO_1232 (O_1232,N_48672,N_49378);
nor UO_1233 (O_1233,N_48521,N_49114);
or UO_1234 (O_1234,N_48255,N_48230);
nand UO_1235 (O_1235,N_48096,N_49922);
and UO_1236 (O_1236,N_48123,N_49541);
nor UO_1237 (O_1237,N_48450,N_49065);
nand UO_1238 (O_1238,N_48866,N_48926);
and UO_1239 (O_1239,N_49652,N_48656);
nand UO_1240 (O_1240,N_48564,N_48377);
nor UO_1241 (O_1241,N_48682,N_49695);
nand UO_1242 (O_1242,N_48697,N_49444);
nor UO_1243 (O_1243,N_49555,N_48712);
or UO_1244 (O_1244,N_49112,N_49926);
xnor UO_1245 (O_1245,N_48727,N_49314);
nor UO_1246 (O_1246,N_49452,N_49070);
xor UO_1247 (O_1247,N_49816,N_49474);
or UO_1248 (O_1248,N_48258,N_48327);
nand UO_1249 (O_1249,N_49534,N_49199);
nand UO_1250 (O_1250,N_49698,N_48195);
or UO_1251 (O_1251,N_48343,N_49873);
nor UO_1252 (O_1252,N_48336,N_48709);
and UO_1253 (O_1253,N_49144,N_48134);
nand UO_1254 (O_1254,N_48403,N_48334);
and UO_1255 (O_1255,N_49904,N_48471);
and UO_1256 (O_1256,N_49113,N_48304);
and UO_1257 (O_1257,N_48897,N_49409);
nand UO_1258 (O_1258,N_49224,N_48696);
xnor UO_1259 (O_1259,N_49403,N_49451);
nor UO_1260 (O_1260,N_48190,N_49747);
nand UO_1261 (O_1261,N_49545,N_48818);
or UO_1262 (O_1262,N_49192,N_48882);
xor UO_1263 (O_1263,N_49611,N_49510);
xor UO_1264 (O_1264,N_48635,N_48514);
nand UO_1265 (O_1265,N_49560,N_48291);
and UO_1266 (O_1266,N_48231,N_49972);
and UO_1267 (O_1267,N_48438,N_48886);
nor UO_1268 (O_1268,N_48882,N_49450);
and UO_1269 (O_1269,N_49773,N_48605);
and UO_1270 (O_1270,N_48612,N_48760);
and UO_1271 (O_1271,N_48176,N_48687);
and UO_1272 (O_1272,N_48315,N_49241);
and UO_1273 (O_1273,N_48699,N_49504);
and UO_1274 (O_1274,N_48180,N_49781);
nor UO_1275 (O_1275,N_49653,N_48093);
nor UO_1276 (O_1276,N_48565,N_49233);
nor UO_1277 (O_1277,N_48564,N_48259);
nand UO_1278 (O_1278,N_48445,N_49145);
xnor UO_1279 (O_1279,N_49108,N_49598);
xor UO_1280 (O_1280,N_48211,N_48403);
xor UO_1281 (O_1281,N_49767,N_49787);
nor UO_1282 (O_1282,N_49280,N_48346);
nand UO_1283 (O_1283,N_49667,N_49033);
or UO_1284 (O_1284,N_49490,N_49390);
nand UO_1285 (O_1285,N_49506,N_49967);
nand UO_1286 (O_1286,N_48444,N_48676);
nand UO_1287 (O_1287,N_48779,N_49406);
nor UO_1288 (O_1288,N_49589,N_48309);
nand UO_1289 (O_1289,N_49245,N_49516);
xnor UO_1290 (O_1290,N_49534,N_48963);
nand UO_1291 (O_1291,N_49588,N_49458);
nand UO_1292 (O_1292,N_48534,N_49604);
or UO_1293 (O_1293,N_49670,N_48911);
or UO_1294 (O_1294,N_48827,N_48148);
or UO_1295 (O_1295,N_48585,N_49342);
xor UO_1296 (O_1296,N_49421,N_49891);
xor UO_1297 (O_1297,N_48831,N_49757);
nand UO_1298 (O_1298,N_49006,N_49287);
and UO_1299 (O_1299,N_48251,N_48892);
and UO_1300 (O_1300,N_49892,N_48552);
nor UO_1301 (O_1301,N_48738,N_49666);
xor UO_1302 (O_1302,N_48412,N_49425);
xnor UO_1303 (O_1303,N_48081,N_48065);
nand UO_1304 (O_1304,N_48589,N_48629);
xnor UO_1305 (O_1305,N_48075,N_49443);
or UO_1306 (O_1306,N_48601,N_49706);
xor UO_1307 (O_1307,N_48719,N_48456);
nor UO_1308 (O_1308,N_49081,N_49117);
nand UO_1309 (O_1309,N_48284,N_49048);
and UO_1310 (O_1310,N_49751,N_48912);
nand UO_1311 (O_1311,N_48327,N_49881);
and UO_1312 (O_1312,N_48681,N_48491);
nor UO_1313 (O_1313,N_48594,N_49587);
and UO_1314 (O_1314,N_48185,N_49845);
nor UO_1315 (O_1315,N_49079,N_49286);
or UO_1316 (O_1316,N_48954,N_48970);
xnor UO_1317 (O_1317,N_48876,N_49830);
or UO_1318 (O_1318,N_49696,N_48230);
xnor UO_1319 (O_1319,N_49443,N_49650);
xnor UO_1320 (O_1320,N_48644,N_49116);
nor UO_1321 (O_1321,N_49302,N_49210);
nand UO_1322 (O_1322,N_49261,N_48259);
nor UO_1323 (O_1323,N_48238,N_49700);
and UO_1324 (O_1324,N_48807,N_48311);
xnor UO_1325 (O_1325,N_49307,N_49898);
nand UO_1326 (O_1326,N_48160,N_48066);
nor UO_1327 (O_1327,N_49521,N_48592);
nor UO_1328 (O_1328,N_48212,N_48956);
and UO_1329 (O_1329,N_48592,N_48471);
nand UO_1330 (O_1330,N_49431,N_48961);
or UO_1331 (O_1331,N_48822,N_49545);
nand UO_1332 (O_1332,N_48595,N_49702);
nand UO_1333 (O_1333,N_48021,N_49141);
xnor UO_1334 (O_1334,N_48013,N_48147);
or UO_1335 (O_1335,N_49941,N_49670);
or UO_1336 (O_1336,N_48903,N_49325);
or UO_1337 (O_1337,N_48657,N_49867);
nor UO_1338 (O_1338,N_48526,N_48701);
xnor UO_1339 (O_1339,N_48652,N_49455);
nand UO_1340 (O_1340,N_48284,N_48513);
nor UO_1341 (O_1341,N_48223,N_48574);
or UO_1342 (O_1342,N_48676,N_49759);
nor UO_1343 (O_1343,N_49699,N_49123);
nor UO_1344 (O_1344,N_48525,N_48092);
or UO_1345 (O_1345,N_48401,N_48862);
xnor UO_1346 (O_1346,N_48862,N_48185);
nor UO_1347 (O_1347,N_49453,N_49631);
or UO_1348 (O_1348,N_48137,N_49754);
nand UO_1349 (O_1349,N_48023,N_48004);
xor UO_1350 (O_1350,N_49640,N_48757);
or UO_1351 (O_1351,N_48500,N_49010);
nand UO_1352 (O_1352,N_48801,N_49526);
and UO_1353 (O_1353,N_48397,N_48922);
nand UO_1354 (O_1354,N_49916,N_49608);
nor UO_1355 (O_1355,N_49963,N_48377);
nor UO_1356 (O_1356,N_48928,N_48500);
nor UO_1357 (O_1357,N_48605,N_48420);
or UO_1358 (O_1358,N_49029,N_49133);
nand UO_1359 (O_1359,N_48839,N_48426);
nand UO_1360 (O_1360,N_48167,N_49168);
nor UO_1361 (O_1361,N_49108,N_48893);
or UO_1362 (O_1362,N_49339,N_48782);
nor UO_1363 (O_1363,N_48563,N_49055);
nand UO_1364 (O_1364,N_48403,N_48481);
or UO_1365 (O_1365,N_49048,N_49784);
nor UO_1366 (O_1366,N_49412,N_49574);
or UO_1367 (O_1367,N_48112,N_48314);
and UO_1368 (O_1368,N_49963,N_48118);
xnor UO_1369 (O_1369,N_49066,N_48816);
nor UO_1370 (O_1370,N_49575,N_49868);
nand UO_1371 (O_1371,N_49409,N_48800);
and UO_1372 (O_1372,N_49424,N_49327);
and UO_1373 (O_1373,N_49172,N_49047);
or UO_1374 (O_1374,N_48156,N_49134);
or UO_1375 (O_1375,N_48605,N_49099);
and UO_1376 (O_1376,N_48161,N_48213);
and UO_1377 (O_1377,N_48077,N_48921);
or UO_1378 (O_1378,N_49107,N_49707);
xnor UO_1379 (O_1379,N_48130,N_49643);
nor UO_1380 (O_1380,N_48683,N_48549);
nand UO_1381 (O_1381,N_48406,N_49490);
or UO_1382 (O_1382,N_48877,N_48738);
xor UO_1383 (O_1383,N_49913,N_49262);
nor UO_1384 (O_1384,N_48928,N_48014);
and UO_1385 (O_1385,N_49580,N_48143);
and UO_1386 (O_1386,N_48877,N_48594);
or UO_1387 (O_1387,N_49478,N_48412);
or UO_1388 (O_1388,N_49365,N_49254);
xnor UO_1389 (O_1389,N_49337,N_48578);
nor UO_1390 (O_1390,N_48824,N_48471);
and UO_1391 (O_1391,N_48193,N_48811);
nor UO_1392 (O_1392,N_49648,N_48017);
and UO_1393 (O_1393,N_48855,N_48779);
xor UO_1394 (O_1394,N_48176,N_49785);
nor UO_1395 (O_1395,N_49421,N_49231);
or UO_1396 (O_1396,N_48751,N_48507);
nand UO_1397 (O_1397,N_48558,N_48526);
nor UO_1398 (O_1398,N_48736,N_48694);
and UO_1399 (O_1399,N_49244,N_48576);
nor UO_1400 (O_1400,N_48299,N_48458);
or UO_1401 (O_1401,N_49500,N_49656);
xor UO_1402 (O_1402,N_49113,N_49329);
nor UO_1403 (O_1403,N_49821,N_49766);
or UO_1404 (O_1404,N_48392,N_48246);
or UO_1405 (O_1405,N_48622,N_48876);
nand UO_1406 (O_1406,N_48412,N_48169);
xnor UO_1407 (O_1407,N_49380,N_48486);
or UO_1408 (O_1408,N_48380,N_49966);
nor UO_1409 (O_1409,N_48034,N_48496);
nor UO_1410 (O_1410,N_48238,N_48821);
and UO_1411 (O_1411,N_48608,N_49474);
nor UO_1412 (O_1412,N_49078,N_48472);
xnor UO_1413 (O_1413,N_49623,N_48976);
and UO_1414 (O_1414,N_49406,N_48624);
xor UO_1415 (O_1415,N_48857,N_49856);
xnor UO_1416 (O_1416,N_48438,N_48820);
nand UO_1417 (O_1417,N_48157,N_49897);
nor UO_1418 (O_1418,N_48920,N_49747);
or UO_1419 (O_1419,N_49680,N_48390);
nand UO_1420 (O_1420,N_48086,N_49321);
nor UO_1421 (O_1421,N_49894,N_48930);
or UO_1422 (O_1422,N_49791,N_49756);
or UO_1423 (O_1423,N_49526,N_49068);
xor UO_1424 (O_1424,N_49679,N_48405);
nand UO_1425 (O_1425,N_48440,N_49060);
or UO_1426 (O_1426,N_49854,N_48548);
or UO_1427 (O_1427,N_49601,N_49498);
and UO_1428 (O_1428,N_49231,N_49958);
xnor UO_1429 (O_1429,N_49623,N_48226);
and UO_1430 (O_1430,N_49322,N_49453);
or UO_1431 (O_1431,N_48991,N_48188);
xor UO_1432 (O_1432,N_49714,N_49848);
nor UO_1433 (O_1433,N_48270,N_49929);
and UO_1434 (O_1434,N_48306,N_49740);
or UO_1435 (O_1435,N_49106,N_48856);
or UO_1436 (O_1436,N_48606,N_49791);
and UO_1437 (O_1437,N_48242,N_49378);
nor UO_1438 (O_1438,N_48071,N_48537);
or UO_1439 (O_1439,N_49413,N_48356);
nor UO_1440 (O_1440,N_49022,N_48175);
nand UO_1441 (O_1441,N_48368,N_48446);
xor UO_1442 (O_1442,N_49261,N_48341);
nand UO_1443 (O_1443,N_49893,N_48360);
and UO_1444 (O_1444,N_49753,N_49824);
nand UO_1445 (O_1445,N_49458,N_48418);
nand UO_1446 (O_1446,N_48313,N_48255);
or UO_1447 (O_1447,N_49463,N_48383);
and UO_1448 (O_1448,N_48673,N_48756);
and UO_1449 (O_1449,N_49997,N_49341);
nand UO_1450 (O_1450,N_49168,N_49387);
and UO_1451 (O_1451,N_48104,N_48534);
nand UO_1452 (O_1452,N_49292,N_49151);
nand UO_1453 (O_1453,N_48144,N_49441);
nand UO_1454 (O_1454,N_48875,N_48003);
nor UO_1455 (O_1455,N_49960,N_49491);
nand UO_1456 (O_1456,N_48491,N_48408);
nor UO_1457 (O_1457,N_49057,N_49577);
nand UO_1458 (O_1458,N_49485,N_49231);
and UO_1459 (O_1459,N_49011,N_48037);
and UO_1460 (O_1460,N_49772,N_49889);
nor UO_1461 (O_1461,N_48111,N_48371);
nor UO_1462 (O_1462,N_48125,N_49732);
or UO_1463 (O_1463,N_49244,N_49474);
and UO_1464 (O_1464,N_49869,N_48458);
nor UO_1465 (O_1465,N_48344,N_49813);
nor UO_1466 (O_1466,N_48899,N_49414);
nor UO_1467 (O_1467,N_49334,N_48554);
nor UO_1468 (O_1468,N_49671,N_49745);
nand UO_1469 (O_1469,N_48298,N_48148);
xor UO_1470 (O_1470,N_48754,N_49804);
xnor UO_1471 (O_1471,N_48923,N_49545);
or UO_1472 (O_1472,N_49091,N_49722);
or UO_1473 (O_1473,N_49407,N_49870);
nor UO_1474 (O_1474,N_49706,N_49937);
nand UO_1475 (O_1475,N_49783,N_48735);
or UO_1476 (O_1476,N_49735,N_48957);
and UO_1477 (O_1477,N_48579,N_48679);
nor UO_1478 (O_1478,N_48815,N_48987);
nand UO_1479 (O_1479,N_49618,N_49751);
nand UO_1480 (O_1480,N_49996,N_49897);
nor UO_1481 (O_1481,N_49884,N_48762);
xor UO_1482 (O_1482,N_48966,N_49823);
nand UO_1483 (O_1483,N_48354,N_49274);
or UO_1484 (O_1484,N_49619,N_48541);
and UO_1485 (O_1485,N_49261,N_48002);
xor UO_1486 (O_1486,N_48585,N_48774);
xor UO_1487 (O_1487,N_49246,N_48979);
and UO_1488 (O_1488,N_48638,N_49165);
or UO_1489 (O_1489,N_49005,N_48081);
nor UO_1490 (O_1490,N_49089,N_49840);
xor UO_1491 (O_1491,N_49220,N_49932);
nor UO_1492 (O_1492,N_48634,N_48806);
and UO_1493 (O_1493,N_48070,N_48614);
or UO_1494 (O_1494,N_49892,N_48238);
nand UO_1495 (O_1495,N_49230,N_48156);
xnor UO_1496 (O_1496,N_48446,N_48228);
nor UO_1497 (O_1497,N_49751,N_48116);
xor UO_1498 (O_1498,N_49502,N_49394);
and UO_1499 (O_1499,N_49813,N_49096);
or UO_1500 (O_1500,N_48808,N_49687);
and UO_1501 (O_1501,N_49331,N_48699);
or UO_1502 (O_1502,N_48778,N_48297);
nor UO_1503 (O_1503,N_48913,N_49476);
xor UO_1504 (O_1504,N_49156,N_49719);
and UO_1505 (O_1505,N_48524,N_48068);
nor UO_1506 (O_1506,N_48950,N_48392);
xor UO_1507 (O_1507,N_49363,N_49551);
nor UO_1508 (O_1508,N_49247,N_48043);
xor UO_1509 (O_1509,N_49260,N_48079);
nand UO_1510 (O_1510,N_48178,N_49347);
nand UO_1511 (O_1511,N_48649,N_49676);
and UO_1512 (O_1512,N_48830,N_48050);
xor UO_1513 (O_1513,N_49265,N_49264);
and UO_1514 (O_1514,N_48704,N_48983);
nor UO_1515 (O_1515,N_48056,N_48070);
xor UO_1516 (O_1516,N_48531,N_48962);
or UO_1517 (O_1517,N_49557,N_49027);
xor UO_1518 (O_1518,N_48794,N_49899);
nor UO_1519 (O_1519,N_49708,N_48954);
nand UO_1520 (O_1520,N_48584,N_49038);
or UO_1521 (O_1521,N_48173,N_48052);
and UO_1522 (O_1522,N_48804,N_48699);
and UO_1523 (O_1523,N_49832,N_49268);
and UO_1524 (O_1524,N_49856,N_48423);
nor UO_1525 (O_1525,N_49946,N_48682);
nand UO_1526 (O_1526,N_49591,N_48088);
nand UO_1527 (O_1527,N_49433,N_49693);
and UO_1528 (O_1528,N_48761,N_49231);
nor UO_1529 (O_1529,N_49290,N_48686);
xnor UO_1530 (O_1530,N_49081,N_49590);
or UO_1531 (O_1531,N_49669,N_48092);
or UO_1532 (O_1532,N_49556,N_48143);
or UO_1533 (O_1533,N_48804,N_48457);
and UO_1534 (O_1534,N_49621,N_48960);
and UO_1535 (O_1535,N_48555,N_49742);
nand UO_1536 (O_1536,N_48336,N_49649);
or UO_1537 (O_1537,N_48591,N_49397);
or UO_1538 (O_1538,N_49751,N_48620);
and UO_1539 (O_1539,N_48103,N_49936);
nand UO_1540 (O_1540,N_48862,N_49998);
and UO_1541 (O_1541,N_49776,N_49589);
and UO_1542 (O_1542,N_48780,N_48496);
nor UO_1543 (O_1543,N_48612,N_49758);
xnor UO_1544 (O_1544,N_48520,N_48546);
nand UO_1545 (O_1545,N_48010,N_48878);
or UO_1546 (O_1546,N_49995,N_49775);
and UO_1547 (O_1547,N_49085,N_49983);
nor UO_1548 (O_1548,N_48374,N_48553);
xnor UO_1549 (O_1549,N_49694,N_49426);
nor UO_1550 (O_1550,N_49362,N_48948);
or UO_1551 (O_1551,N_48170,N_49268);
or UO_1552 (O_1552,N_49986,N_48607);
nor UO_1553 (O_1553,N_49197,N_48769);
nand UO_1554 (O_1554,N_49419,N_48049);
nor UO_1555 (O_1555,N_48007,N_48748);
nand UO_1556 (O_1556,N_49584,N_49524);
nand UO_1557 (O_1557,N_49809,N_48803);
xnor UO_1558 (O_1558,N_49340,N_48470);
nor UO_1559 (O_1559,N_49360,N_48948);
or UO_1560 (O_1560,N_49253,N_49527);
nor UO_1561 (O_1561,N_49408,N_48311);
nor UO_1562 (O_1562,N_49967,N_49163);
or UO_1563 (O_1563,N_49513,N_49056);
xnor UO_1564 (O_1564,N_49355,N_49322);
and UO_1565 (O_1565,N_48574,N_49550);
nand UO_1566 (O_1566,N_48418,N_49521);
nand UO_1567 (O_1567,N_48333,N_49116);
and UO_1568 (O_1568,N_48572,N_49819);
xor UO_1569 (O_1569,N_48835,N_48352);
and UO_1570 (O_1570,N_48618,N_49035);
nand UO_1571 (O_1571,N_49817,N_48824);
nor UO_1572 (O_1572,N_48965,N_49500);
nor UO_1573 (O_1573,N_48933,N_49730);
or UO_1574 (O_1574,N_49729,N_48246);
xnor UO_1575 (O_1575,N_48119,N_49074);
xor UO_1576 (O_1576,N_48531,N_49592);
xor UO_1577 (O_1577,N_49358,N_49952);
or UO_1578 (O_1578,N_49496,N_48012);
or UO_1579 (O_1579,N_49679,N_49287);
or UO_1580 (O_1580,N_49478,N_48745);
nand UO_1581 (O_1581,N_48575,N_49842);
xor UO_1582 (O_1582,N_49012,N_49654);
xnor UO_1583 (O_1583,N_49069,N_48324);
or UO_1584 (O_1584,N_49116,N_48533);
or UO_1585 (O_1585,N_48681,N_49399);
nor UO_1586 (O_1586,N_49029,N_48333);
nand UO_1587 (O_1587,N_48737,N_49015);
nor UO_1588 (O_1588,N_49003,N_48831);
xnor UO_1589 (O_1589,N_48010,N_48564);
nand UO_1590 (O_1590,N_49509,N_49464);
xor UO_1591 (O_1591,N_48142,N_48102);
xnor UO_1592 (O_1592,N_49762,N_49387);
xnor UO_1593 (O_1593,N_49197,N_49036);
nand UO_1594 (O_1594,N_48022,N_49298);
nor UO_1595 (O_1595,N_49772,N_48102);
nor UO_1596 (O_1596,N_49119,N_49666);
and UO_1597 (O_1597,N_48783,N_49503);
xnor UO_1598 (O_1598,N_49436,N_48834);
xnor UO_1599 (O_1599,N_49314,N_49118);
nor UO_1600 (O_1600,N_49608,N_49569);
xnor UO_1601 (O_1601,N_49499,N_49429);
nand UO_1602 (O_1602,N_48233,N_49653);
and UO_1603 (O_1603,N_49420,N_49431);
or UO_1604 (O_1604,N_49306,N_48276);
nand UO_1605 (O_1605,N_49690,N_49698);
and UO_1606 (O_1606,N_49106,N_49100);
nor UO_1607 (O_1607,N_48601,N_48795);
xnor UO_1608 (O_1608,N_48200,N_49580);
nor UO_1609 (O_1609,N_49081,N_49074);
nor UO_1610 (O_1610,N_49569,N_48347);
nand UO_1611 (O_1611,N_48550,N_48111);
nand UO_1612 (O_1612,N_49441,N_49503);
and UO_1613 (O_1613,N_49194,N_49468);
nand UO_1614 (O_1614,N_48941,N_48196);
xor UO_1615 (O_1615,N_48933,N_49094);
nand UO_1616 (O_1616,N_49149,N_48684);
nor UO_1617 (O_1617,N_49994,N_49576);
nor UO_1618 (O_1618,N_49040,N_48752);
and UO_1619 (O_1619,N_49877,N_48164);
xnor UO_1620 (O_1620,N_48787,N_49192);
nor UO_1621 (O_1621,N_49965,N_48359);
xor UO_1622 (O_1622,N_48863,N_48888);
xnor UO_1623 (O_1623,N_48394,N_49805);
and UO_1624 (O_1624,N_49861,N_48964);
nand UO_1625 (O_1625,N_49520,N_48394);
nand UO_1626 (O_1626,N_48333,N_49862);
nand UO_1627 (O_1627,N_49552,N_49791);
nor UO_1628 (O_1628,N_49573,N_48972);
nor UO_1629 (O_1629,N_48624,N_49151);
or UO_1630 (O_1630,N_49318,N_49385);
or UO_1631 (O_1631,N_48398,N_48328);
nand UO_1632 (O_1632,N_49553,N_49515);
and UO_1633 (O_1633,N_48094,N_49503);
and UO_1634 (O_1634,N_48407,N_49731);
nand UO_1635 (O_1635,N_48677,N_48349);
and UO_1636 (O_1636,N_49050,N_49932);
and UO_1637 (O_1637,N_48521,N_48202);
or UO_1638 (O_1638,N_48911,N_48402);
and UO_1639 (O_1639,N_49705,N_48102);
and UO_1640 (O_1640,N_48205,N_49736);
or UO_1641 (O_1641,N_49514,N_48354);
nand UO_1642 (O_1642,N_49272,N_48676);
nand UO_1643 (O_1643,N_49803,N_48272);
xnor UO_1644 (O_1644,N_48164,N_49543);
xor UO_1645 (O_1645,N_49648,N_48249);
or UO_1646 (O_1646,N_49373,N_49673);
nand UO_1647 (O_1647,N_48586,N_48775);
nor UO_1648 (O_1648,N_49065,N_48350);
nor UO_1649 (O_1649,N_48311,N_48671);
xor UO_1650 (O_1650,N_49510,N_49332);
or UO_1651 (O_1651,N_48142,N_48129);
xnor UO_1652 (O_1652,N_48088,N_48397);
and UO_1653 (O_1653,N_49100,N_48202);
and UO_1654 (O_1654,N_49343,N_48672);
and UO_1655 (O_1655,N_49573,N_48527);
nand UO_1656 (O_1656,N_49052,N_48083);
or UO_1657 (O_1657,N_49372,N_48700);
nand UO_1658 (O_1658,N_48302,N_48161);
or UO_1659 (O_1659,N_48156,N_49439);
xor UO_1660 (O_1660,N_48394,N_49718);
nand UO_1661 (O_1661,N_48427,N_49278);
xnor UO_1662 (O_1662,N_48420,N_48274);
and UO_1663 (O_1663,N_48504,N_49999);
xor UO_1664 (O_1664,N_49518,N_49408);
or UO_1665 (O_1665,N_49730,N_49092);
xor UO_1666 (O_1666,N_48636,N_48761);
nor UO_1667 (O_1667,N_49206,N_48486);
or UO_1668 (O_1668,N_48484,N_48524);
xnor UO_1669 (O_1669,N_48861,N_48245);
xor UO_1670 (O_1670,N_48292,N_48106);
or UO_1671 (O_1671,N_48968,N_48244);
or UO_1672 (O_1672,N_49712,N_48249);
xor UO_1673 (O_1673,N_49945,N_49058);
xor UO_1674 (O_1674,N_48193,N_48241);
or UO_1675 (O_1675,N_49853,N_49070);
nand UO_1676 (O_1676,N_48574,N_48208);
and UO_1677 (O_1677,N_49526,N_48625);
nor UO_1678 (O_1678,N_49817,N_49245);
xor UO_1679 (O_1679,N_48362,N_49732);
nor UO_1680 (O_1680,N_49457,N_49633);
or UO_1681 (O_1681,N_48544,N_48306);
and UO_1682 (O_1682,N_48649,N_48622);
nor UO_1683 (O_1683,N_49799,N_48375);
xor UO_1684 (O_1684,N_48731,N_48852);
xnor UO_1685 (O_1685,N_49450,N_48759);
nand UO_1686 (O_1686,N_49299,N_48748);
and UO_1687 (O_1687,N_48819,N_49089);
xor UO_1688 (O_1688,N_49753,N_49894);
nor UO_1689 (O_1689,N_49418,N_49900);
xor UO_1690 (O_1690,N_48358,N_49694);
or UO_1691 (O_1691,N_49324,N_49210);
xor UO_1692 (O_1692,N_49105,N_48881);
xor UO_1693 (O_1693,N_48937,N_49943);
and UO_1694 (O_1694,N_48284,N_49955);
xor UO_1695 (O_1695,N_48755,N_48423);
xnor UO_1696 (O_1696,N_49178,N_49262);
nor UO_1697 (O_1697,N_48725,N_49625);
and UO_1698 (O_1698,N_48695,N_48272);
or UO_1699 (O_1699,N_49641,N_48945);
xnor UO_1700 (O_1700,N_49209,N_48511);
nand UO_1701 (O_1701,N_49507,N_48750);
xnor UO_1702 (O_1702,N_49979,N_49891);
and UO_1703 (O_1703,N_48654,N_49716);
nor UO_1704 (O_1704,N_49279,N_48211);
nand UO_1705 (O_1705,N_49428,N_49174);
and UO_1706 (O_1706,N_48822,N_48713);
xnor UO_1707 (O_1707,N_49973,N_49900);
nand UO_1708 (O_1708,N_49025,N_49115);
nand UO_1709 (O_1709,N_48824,N_48218);
nand UO_1710 (O_1710,N_48257,N_48085);
nor UO_1711 (O_1711,N_48994,N_49882);
nand UO_1712 (O_1712,N_48297,N_48348);
nor UO_1713 (O_1713,N_48022,N_48409);
nor UO_1714 (O_1714,N_48710,N_48242);
or UO_1715 (O_1715,N_49116,N_49551);
or UO_1716 (O_1716,N_49731,N_48546);
and UO_1717 (O_1717,N_49696,N_48698);
nor UO_1718 (O_1718,N_48598,N_49941);
and UO_1719 (O_1719,N_48808,N_49537);
nor UO_1720 (O_1720,N_49265,N_49206);
nor UO_1721 (O_1721,N_48559,N_48931);
and UO_1722 (O_1722,N_48088,N_49894);
and UO_1723 (O_1723,N_49855,N_49401);
or UO_1724 (O_1724,N_49057,N_48324);
nand UO_1725 (O_1725,N_48632,N_48881);
xnor UO_1726 (O_1726,N_48124,N_48973);
nor UO_1727 (O_1727,N_49709,N_48033);
and UO_1728 (O_1728,N_48237,N_48770);
or UO_1729 (O_1729,N_49368,N_49790);
nor UO_1730 (O_1730,N_49389,N_49159);
xor UO_1731 (O_1731,N_48531,N_49415);
nor UO_1732 (O_1732,N_48790,N_48003);
or UO_1733 (O_1733,N_49135,N_48607);
and UO_1734 (O_1734,N_48594,N_49508);
xor UO_1735 (O_1735,N_49437,N_49469);
and UO_1736 (O_1736,N_49465,N_48041);
nor UO_1737 (O_1737,N_49995,N_49269);
xnor UO_1738 (O_1738,N_49148,N_49853);
xor UO_1739 (O_1739,N_48291,N_49759);
or UO_1740 (O_1740,N_48267,N_48230);
nor UO_1741 (O_1741,N_49117,N_49806);
nor UO_1742 (O_1742,N_49733,N_49819);
or UO_1743 (O_1743,N_49478,N_49143);
and UO_1744 (O_1744,N_48609,N_49939);
and UO_1745 (O_1745,N_48061,N_49677);
nand UO_1746 (O_1746,N_49453,N_48816);
nand UO_1747 (O_1747,N_48033,N_49333);
xor UO_1748 (O_1748,N_48565,N_48916);
and UO_1749 (O_1749,N_49145,N_49358);
nor UO_1750 (O_1750,N_49688,N_49227);
or UO_1751 (O_1751,N_49049,N_49738);
nor UO_1752 (O_1752,N_48501,N_48258);
or UO_1753 (O_1753,N_49782,N_48045);
xor UO_1754 (O_1754,N_49924,N_48297);
or UO_1755 (O_1755,N_48028,N_48733);
or UO_1756 (O_1756,N_48090,N_49993);
or UO_1757 (O_1757,N_48817,N_48025);
xnor UO_1758 (O_1758,N_49634,N_49451);
xnor UO_1759 (O_1759,N_49797,N_48508);
or UO_1760 (O_1760,N_49124,N_48583);
nand UO_1761 (O_1761,N_48320,N_49626);
nand UO_1762 (O_1762,N_48054,N_48403);
nand UO_1763 (O_1763,N_48722,N_49560);
and UO_1764 (O_1764,N_49194,N_49771);
nand UO_1765 (O_1765,N_49423,N_48294);
and UO_1766 (O_1766,N_48667,N_49887);
nor UO_1767 (O_1767,N_49349,N_48693);
nor UO_1768 (O_1768,N_49730,N_48384);
xor UO_1769 (O_1769,N_49721,N_48043);
xnor UO_1770 (O_1770,N_48874,N_49137);
xnor UO_1771 (O_1771,N_48384,N_49612);
nor UO_1772 (O_1772,N_49382,N_48955);
or UO_1773 (O_1773,N_48364,N_48401);
or UO_1774 (O_1774,N_49792,N_49121);
xnor UO_1775 (O_1775,N_48591,N_49640);
nand UO_1776 (O_1776,N_48339,N_48323);
nand UO_1777 (O_1777,N_49895,N_48837);
and UO_1778 (O_1778,N_48997,N_49402);
and UO_1779 (O_1779,N_49201,N_49936);
xnor UO_1780 (O_1780,N_48327,N_48170);
nand UO_1781 (O_1781,N_48757,N_49902);
nand UO_1782 (O_1782,N_48905,N_48606);
xor UO_1783 (O_1783,N_48053,N_49733);
and UO_1784 (O_1784,N_49690,N_49076);
nor UO_1785 (O_1785,N_49734,N_49676);
and UO_1786 (O_1786,N_49973,N_49244);
or UO_1787 (O_1787,N_49714,N_49797);
xnor UO_1788 (O_1788,N_49112,N_49173);
and UO_1789 (O_1789,N_48348,N_49637);
nor UO_1790 (O_1790,N_49271,N_48262);
and UO_1791 (O_1791,N_48355,N_48064);
or UO_1792 (O_1792,N_48028,N_48948);
and UO_1793 (O_1793,N_48416,N_48078);
and UO_1794 (O_1794,N_48890,N_48287);
and UO_1795 (O_1795,N_49938,N_49766);
or UO_1796 (O_1796,N_49119,N_48380);
nor UO_1797 (O_1797,N_49500,N_49352);
nand UO_1798 (O_1798,N_49434,N_48400);
and UO_1799 (O_1799,N_48932,N_49737);
and UO_1800 (O_1800,N_48714,N_48237);
nand UO_1801 (O_1801,N_49395,N_49870);
nor UO_1802 (O_1802,N_48336,N_48610);
nand UO_1803 (O_1803,N_48713,N_49215);
nor UO_1804 (O_1804,N_49907,N_49253);
nor UO_1805 (O_1805,N_49847,N_48221);
xor UO_1806 (O_1806,N_48007,N_49560);
or UO_1807 (O_1807,N_49499,N_49335);
nor UO_1808 (O_1808,N_49585,N_49426);
or UO_1809 (O_1809,N_48053,N_48836);
nand UO_1810 (O_1810,N_49171,N_49308);
nand UO_1811 (O_1811,N_49152,N_48422);
xor UO_1812 (O_1812,N_48895,N_49326);
nand UO_1813 (O_1813,N_48534,N_49253);
nor UO_1814 (O_1814,N_49632,N_48978);
nand UO_1815 (O_1815,N_49989,N_49176);
nand UO_1816 (O_1816,N_48852,N_49719);
or UO_1817 (O_1817,N_48899,N_49150);
nand UO_1818 (O_1818,N_49912,N_48467);
nand UO_1819 (O_1819,N_48975,N_48905);
xor UO_1820 (O_1820,N_48663,N_48201);
and UO_1821 (O_1821,N_48503,N_48401);
and UO_1822 (O_1822,N_48041,N_48160);
nand UO_1823 (O_1823,N_49527,N_48083);
xnor UO_1824 (O_1824,N_48102,N_48491);
or UO_1825 (O_1825,N_48090,N_49186);
xnor UO_1826 (O_1826,N_48369,N_48129);
nor UO_1827 (O_1827,N_48181,N_48827);
nor UO_1828 (O_1828,N_49624,N_48421);
xnor UO_1829 (O_1829,N_49847,N_48191);
and UO_1830 (O_1830,N_48581,N_48145);
or UO_1831 (O_1831,N_48127,N_48087);
nand UO_1832 (O_1832,N_49020,N_49602);
and UO_1833 (O_1833,N_49321,N_48309);
or UO_1834 (O_1834,N_49147,N_48655);
nand UO_1835 (O_1835,N_48687,N_49946);
and UO_1836 (O_1836,N_48949,N_48638);
nand UO_1837 (O_1837,N_49068,N_48272);
nor UO_1838 (O_1838,N_48148,N_49743);
nor UO_1839 (O_1839,N_48281,N_49066);
nor UO_1840 (O_1840,N_48953,N_49077);
and UO_1841 (O_1841,N_48787,N_48768);
and UO_1842 (O_1842,N_48125,N_49334);
or UO_1843 (O_1843,N_49246,N_49806);
nand UO_1844 (O_1844,N_48088,N_49946);
nor UO_1845 (O_1845,N_49718,N_48904);
xnor UO_1846 (O_1846,N_48424,N_48032);
xor UO_1847 (O_1847,N_48064,N_49451);
nor UO_1848 (O_1848,N_48124,N_49004);
and UO_1849 (O_1849,N_49613,N_49944);
or UO_1850 (O_1850,N_49811,N_48113);
nor UO_1851 (O_1851,N_48279,N_48358);
or UO_1852 (O_1852,N_49739,N_49749);
or UO_1853 (O_1853,N_48517,N_49561);
nor UO_1854 (O_1854,N_49503,N_48507);
xnor UO_1855 (O_1855,N_49878,N_49419);
nor UO_1856 (O_1856,N_48496,N_48533);
nor UO_1857 (O_1857,N_48543,N_48164);
nand UO_1858 (O_1858,N_48351,N_48807);
and UO_1859 (O_1859,N_48467,N_48585);
or UO_1860 (O_1860,N_48425,N_49008);
nand UO_1861 (O_1861,N_49388,N_49731);
xor UO_1862 (O_1862,N_49222,N_49919);
and UO_1863 (O_1863,N_48405,N_48356);
nand UO_1864 (O_1864,N_48918,N_49354);
nand UO_1865 (O_1865,N_48276,N_49122);
and UO_1866 (O_1866,N_49030,N_49367);
nand UO_1867 (O_1867,N_49443,N_48938);
nand UO_1868 (O_1868,N_48811,N_48151);
and UO_1869 (O_1869,N_49015,N_48138);
nand UO_1870 (O_1870,N_49440,N_48935);
or UO_1871 (O_1871,N_49484,N_48322);
or UO_1872 (O_1872,N_49915,N_49207);
xor UO_1873 (O_1873,N_48949,N_48055);
xor UO_1874 (O_1874,N_48607,N_48059);
nand UO_1875 (O_1875,N_48444,N_49016);
or UO_1876 (O_1876,N_49805,N_48220);
or UO_1877 (O_1877,N_48648,N_48880);
nor UO_1878 (O_1878,N_48715,N_48075);
nand UO_1879 (O_1879,N_49522,N_48570);
xnor UO_1880 (O_1880,N_49222,N_48486);
nand UO_1881 (O_1881,N_49556,N_48561);
or UO_1882 (O_1882,N_49010,N_49024);
or UO_1883 (O_1883,N_48142,N_49514);
nand UO_1884 (O_1884,N_49245,N_48876);
nand UO_1885 (O_1885,N_49501,N_48748);
xor UO_1886 (O_1886,N_49093,N_49225);
nor UO_1887 (O_1887,N_48905,N_49187);
nand UO_1888 (O_1888,N_49473,N_49827);
and UO_1889 (O_1889,N_48349,N_49006);
nand UO_1890 (O_1890,N_49013,N_49487);
or UO_1891 (O_1891,N_48960,N_48232);
and UO_1892 (O_1892,N_48808,N_48028);
and UO_1893 (O_1893,N_49885,N_49315);
and UO_1894 (O_1894,N_48985,N_48776);
nand UO_1895 (O_1895,N_49283,N_49729);
xnor UO_1896 (O_1896,N_48100,N_49164);
or UO_1897 (O_1897,N_48350,N_49850);
nand UO_1898 (O_1898,N_49228,N_49288);
or UO_1899 (O_1899,N_48841,N_48731);
nor UO_1900 (O_1900,N_48069,N_48968);
xor UO_1901 (O_1901,N_49377,N_49813);
nand UO_1902 (O_1902,N_48363,N_49423);
xor UO_1903 (O_1903,N_48241,N_48526);
nand UO_1904 (O_1904,N_48118,N_49430);
xnor UO_1905 (O_1905,N_48834,N_48176);
xor UO_1906 (O_1906,N_49615,N_48273);
xnor UO_1907 (O_1907,N_48487,N_49878);
nor UO_1908 (O_1908,N_48605,N_49196);
xnor UO_1909 (O_1909,N_49324,N_48292);
nor UO_1910 (O_1910,N_48828,N_49025);
nand UO_1911 (O_1911,N_49151,N_49497);
and UO_1912 (O_1912,N_49713,N_48220);
nor UO_1913 (O_1913,N_48050,N_49679);
and UO_1914 (O_1914,N_49137,N_49603);
or UO_1915 (O_1915,N_48514,N_48405);
or UO_1916 (O_1916,N_48676,N_48559);
nand UO_1917 (O_1917,N_48732,N_48061);
or UO_1918 (O_1918,N_48359,N_49334);
or UO_1919 (O_1919,N_49246,N_48161);
nor UO_1920 (O_1920,N_49266,N_49140);
or UO_1921 (O_1921,N_49317,N_48905);
or UO_1922 (O_1922,N_49760,N_48152);
xnor UO_1923 (O_1923,N_48942,N_48441);
nand UO_1924 (O_1924,N_48052,N_48814);
nand UO_1925 (O_1925,N_48771,N_49859);
xor UO_1926 (O_1926,N_49031,N_48635);
or UO_1927 (O_1927,N_49879,N_48882);
nor UO_1928 (O_1928,N_48014,N_49247);
and UO_1929 (O_1929,N_49202,N_48994);
xnor UO_1930 (O_1930,N_49002,N_49273);
nor UO_1931 (O_1931,N_49736,N_48695);
nor UO_1932 (O_1932,N_48685,N_48398);
nand UO_1933 (O_1933,N_49154,N_49309);
xnor UO_1934 (O_1934,N_48494,N_49629);
nor UO_1935 (O_1935,N_48852,N_49854);
and UO_1936 (O_1936,N_49154,N_48268);
or UO_1937 (O_1937,N_49509,N_49782);
or UO_1938 (O_1938,N_48449,N_49449);
xnor UO_1939 (O_1939,N_49812,N_49804);
nor UO_1940 (O_1940,N_49985,N_49014);
nor UO_1941 (O_1941,N_48898,N_48178);
nor UO_1942 (O_1942,N_48188,N_48627);
nand UO_1943 (O_1943,N_48343,N_48833);
nor UO_1944 (O_1944,N_49653,N_49445);
nor UO_1945 (O_1945,N_48364,N_49984);
xnor UO_1946 (O_1946,N_48310,N_49769);
and UO_1947 (O_1947,N_48375,N_49635);
nor UO_1948 (O_1948,N_49203,N_48910);
and UO_1949 (O_1949,N_48251,N_48565);
and UO_1950 (O_1950,N_48063,N_48848);
xor UO_1951 (O_1951,N_48489,N_49725);
nor UO_1952 (O_1952,N_48030,N_48770);
and UO_1953 (O_1953,N_48544,N_48257);
xnor UO_1954 (O_1954,N_49528,N_49493);
xnor UO_1955 (O_1955,N_48169,N_48339);
and UO_1956 (O_1956,N_49867,N_48366);
nand UO_1957 (O_1957,N_48142,N_49768);
nand UO_1958 (O_1958,N_49410,N_48250);
or UO_1959 (O_1959,N_49755,N_48871);
xor UO_1960 (O_1960,N_49077,N_49837);
xnor UO_1961 (O_1961,N_48014,N_48345);
xnor UO_1962 (O_1962,N_48854,N_49268);
nand UO_1963 (O_1963,N_49084,N_48360);
and UO_1964 (O_1964,N_48634,N_48594);
nand UO_1965 (O_1965,N_48442,N_48409);
or UO_1966 (O_1966,N_49174,N_48773);
or UO_1967 (O_1967,N_49977,N_48837);
and UO_1968 (O_1968,N_49959,N_49461);
or UO_1969 (O_1969,N_48739,N_49350);
nor UO_1970 (O_1970,N_48329,N_48010);
or UO_1971 (O_1971,N_48844,N_48637);
or UO_1972 (O_1972,N_49159,N_48092);
and UO_1973 (O_1973,N_48399,N_49540);
and UO_1974 (O_1974,N_49936,N_49878);
or UO_1975 (O_1975,N_49663,N_49331);
and UO_1976 (O_1976,N_48048,N_49521);
and UO_1977 (O_1977,N_48709,N_49566);
xnor UO_1978 (O_1978,N_49237,N_48115);
or UO_1979 (O_1979,N_48183,N_49526);
nand UO_1980 (O_1980,N_49303,N_49802);
or UO_1981 (O_1981,N_48190,N_48933);
xor UO_1982 (O_1982,N_48685,N_48214);
xnor UO_1983 (O_1983,N_48466,N_49089);
nand UO_1984 (O_1984,N_49181,N_48161);
xor UO_1985 (O_1985,N_48300,N_48451);
xnor UO_1986 (O_1986,N_48544,N_48526);
or UO_1987 (O_1987,N_49759,N_49569);
or UO_1988 (O_1988,N_49479,N_48089);
and UO_1989 (O_1989,N_49001,N_48276);
and UO_1990 (O_1990,N_49618,N_48279);
nand UO_1991 (O_1991,N_48872,N_48639);
or UO_1992 (O_1992,N_49770,N_49165);
nor UO_1993 (O_1993,N_48451,N_49760);
or UO_1994 (O_1994,N_49690,N_48413);
nor UO_1995 (O_1995,N_48136,N_48742);
nor UO_1996 (O_1996,N_48034,N_49141);
xor UO_1997 (O_1997,N_49795,N_48400);
nor UO_1998 (O_1998,N_49908,N_49634);
xor UO_1999 (O_1999,N_49290,N_48516);
and UO_2000 (O_2000,N_49707,N_49525);
and UO_2001 (O_2001,N_49806,N_49539);
and UO_2002 (O_2002,N_49356,N_48756);
or UO_2003 (O_2003,N_49085,N_48836);
nand UO_2004 (O_2004,N_48414,N_48618);
nor UO_2005 (O_2005,N_48139,N_49394);
xnor UO_2006 (O_2006,N_49598,N_48288);
xor UO_2007 (O_2007,N_49443,N_48841);
and UO_2008 (O_2008,N_49370,N_48688);
xor UO_2009 (O_2009,N_49454,N_49988);
or UO_2010 (O_2010,N_49920,N_49136);
or UO_2011 (O_2011,N_48733,N_48460);
xnor UO_2012 (O_2012,N_49173,N_49360);
or UO_2013 (O_2013,N_48951,N_49630);
and UO_2014 (O_2014,N_49079,N_49542);
nand UO_2015 (O_2015,N_49486,N_48576);
nand UO_2016 (O_2016,N_49880,N_48598);
nand UO_2017 (O_2017,N_48814,N_49848);
nor UO_2018 (O_2018,N_48396,N_48737);
nor UO_2019 (O_2019,N_48373,N_49010);
and UO_2020 (O_2020,N_49585,N_48047);
xor UO_2021 (O_2021,N_49737,N_49897);
nand UO_2022 (O_2022,N_49050,N_48732);
or UO_2023 (O_2023,N_49062,N_48002);
xnor UO_2024 (O_2024,N_48579,N_49045);
xnor UO_2025 (O_2025,N_49759,N_48543);
nor UO_2026 (O_2026,N_48800,N_49115);
and UO_2027 (O_2027,N_49044,N_49262);
and UO_2028 (O_2028,N_49859,N_49068);
and UO_2029 (O_2029,N_48054,N_48906);
and UO_2030 (O_2030,N_48120,N_49869);
xor UO_2031 (O_2031,N_48969,N_49212);
and UO_2032 (O_2032,N_48834,N_49900);
nor UO_2033 (O_2033,N_49906,N_48768);
or UO_2034 (O_2034,N_48350,N_48612);
xnor UO_2035 (O_2035,N_49497,N_49120);
or UO_2036 (O_2036,N_48309,N_48818);
or UO_2037 (O_2037,N_48801,N_48776);
nor UO_2038 (O_2038,N_49782,N_48465);
xnor UO_2039 (O_2039,N_49632,N_48025);
xor UO_2040 (O_2040,N_48794,N_49638);
and UO_2041 (O_2041,N_48234,N_48267);
xor UO_2042 (O_2042,N_49893,N_49553);
nand UO_2043 (O_2043,N_48062,N_48070);
xnor UO_2044 (O_2044,N_49142,N_48180);
and UO_2045 (O_2045,N_48274,N_48187);
and UO_2046 (O_2046,N_48198,N_49502);
xor UO_2047 (O_2047,N_48752,N_48388);
and UO_2048 (O_2048,N_48216,N_49290);
nor UO_2049 (O_2049,N_48018,N_48900);
nor UO_2050 (O_2050,N_48424,N_48363);
nor UO_2051 (O_2051,N_49800,N_48826);
or UO_2052 (O_2052,N_48861,N_48794);
nand UO_2053 (O_2053,N_49351,N_48463);
and UO_2054 (O_2054,N_48667,N_49970);
nand UO_2055 (O_2055,N_49350,N_49770);
xor UO_2056 (O_2056,N_48528,N_49706);
nor UO_2057 (O_2057,N_48632,N_49055);
nand UO_2058 (O_2058,N_49360,N_49538);
nor UO_2059 (O_2059,N_48137,N_49735);
xor UO_2060 (O_2060,N_48162,N_49044);
xnor UO_2061 (O_2061,N_49791,N_49001);
xnor UO_2062 (O_2062,N_48408,N_48972);
nand UO_2063 (O_2063,N_48397,N_48097);
or UO_2064 (O_2064,N_49215,N_49185);
nand UO_2065 (O_2065,N_48141,N_49574);
nor UO_2066 (O_2066,N_49214,N_48413);
xnor UO_2067 (O_2067,N_49023,N_48456);
xnor UO_2068 (O_2068,N_49477,N_49183);
nand UO_2069 (O_2069,N_49268,N_48970);
xnor UO_2070 (O_2070,N_48048,N_49531);
or UO_2071 (O_2071,N_49714,N_48791);
and UO_2072 (O_2072,N_48288,N_48999);
or UO_2073 (O_2073,N_49409,N_49518);
nand UO_2074 (O_2074,N_49384,N_49219);
xnor UO_2075 (O_2075,N_49687,N_48289);
and UO_2076 (O_2076,N_48503,N_48330);
xor UO_2077 (O_2077,N_49556,N_49065);
xnor UO_2078 (O_2078,N_48487,N_48732);
nor UO_2079 (O_2079,N_48473,N_48245);
nor UO_2080 (O_2080,N_49452,N_49338);
and UO_2081 (O_2081,N_48264,N_48671);
nand UO_2082 (O_2082,N_48332,N_49262);
and UO_2083 (O_2083,N_49962,N_48886);
nor UO_2084 (O_2084,N_48244,N_49013);
or UO_2085 (O_2085,N_48941,N_48412);
nor UO_2086 (O_2086,N_49274,N_49367);
and UO_2087 (O_2087,N_49932,N_48601);
nand UO_2088 (O_2088,N_49443,N_49680);
or UO_2089 (O_2089,N_49175,N_48193);
and UO_2090 (O_2090,N_49675,N_49185);
nand UO_2091 (O_2091,N_49305,N_48553);
or UO_2092 (O_2092,N_48841,N_49686);
and UO_2093 (O_2093,N_49828,N_48572);
or UO_2094 (O_2094,N_48091,N_49955);
xor UO_2095 (O_2095,N_49137,N_48087);
xnor UO_2096 (O_2096,N_48565,N_48311);
or UO_2097 (O_2097,N_48790,N_48015);
xor UO_2098 (O_2098,N_48960,N_49492);
xor UO_2099 (O_2099,N_49166,N_49718);
and UO_2100 (O_2100,N_48760,N_49193);
xor UO_2101 (O_2101,N_49825,N_49163);
nor UO_2102 (O_2102,N_49932,N_48828);
nor UO_2103 (O_2103,N_49821,N_48854);
or UO_2104 (O_2104,N_48762,N_48020);
and UO_2105 (O_2105,N_49423,N_49048);
nand UO_2106 (O_2106,N_49632,N_49710);
or UO_2107 (O_2107,N_48127,N_48491);
nor UO_2108 (O_2108,N_48767,N_48580);
nor UO_2109 (O_2109,N_48551,N_48262);
or UO_2110 (O_2110,N_48304,N_48013);
nor UO_2111 (O_2111,N_48057,N_49751);
or UO_2112 (O_2112,N_49638,N_49309);
nand UO_2113 (O_2113,N_49719,N_48153);
nand UO_2114 (O_2114,N_48136,N_48917);
or UO_2115 (O_2115,N_49191,N_48193);
and UO_2116 (O_2116,N_48633,N_49090);
or UO_2117 (O_2117,N_49785,N_48946);
nor UO_2118 (O_2118,N_49835,N_49020);
xnor UO_2119 (O_2119,N_48495,N_49270);
nor UO_2120 (O_2120,N_48250,N_49071);
xor UO_2121 (O_2121,N_48928,N_49946);
nand UO_2122 (O_2122,N_49835,N_48929);
and UO_2123 (O_2123,N_49594,N_49034);
and UO_2124 (O_2124,N_49884,N_48755);
nand UO_2125 (O_2125,N_48280,N_49177);
or UO_2126 (O_2126,N_49808,N_48321);
nand UO_2127 (O_2127,N_48591,N_49295);
and UO_2128 (O_2128,N_49880,N_49238);
nand UO_2129 (O_2129,N_48227,N_49752);
and UO_2130 (O_2130,N_49397,N_49171);
nand UO_2131 (O_2131,N_49954,N_48386);
xor UO_2132 (O_2132,N_49109,N_49093);
xnor UO_2133 (O_2133,N_48395,N_49486);
or UO_2134 (O_2134,N_48078,N_48493);
nor UO_2135 (O_2135,N_48476,N_49003);
and UO_2136 (O_2136,N_49089,N_49807);
nand UO_2137 (O_2137,N_49496,N_49732);
nand UO_2138 (O_2138,N_48047,N_48433);
or UO_2139 (O_2139,N_49391,N_49648);
or UO_2140 (O_2140,N_48045,N_48631);
xnor UO_2141 (O_2141,N_49485,N_48230);
or UO_2142 (O_2142,N_49505,N_48647);
nand UO_2143 (O_2143,N_48605,N_48780);
nor UO_2144 (O_2144,N_48489,N_48460);
nor UO_2145 (O_2145,N_49908,N_49321);
and UO_2146 (O_2146,N_48608,N_49226);
nand UO_2147 (O_2147,N_49423,N_49806);
and UO_2148 (O_2148,N_48275,N_48231);
nand UO_2149 (O_2149,N_48556,N_48642);
nand UO_2150 (O_2150,N_49575,N_48943);
nand UO_2151 (O_2151,N_49397,N_49702);
nand UO_2152 (O_2152,N_48561,N_49934);
nand UO_2153 (O_2153,N_48673,N_48972);
xnor UO_2154 (O_2154,N_49045,N_49936);
nor UO_2155 (O_2155,N_48775,N_49507);
and UO_2156 (O_2156,N_48262,N_49634);
xnor UO_2157 (O_2157,N_49296,N_49373);
and UO_2158 (O_2158,N_48764,N_49016);
xnor UO_2159 (O_2159,N_49952,N_49872);
nor UO_2160 (O_2160,N_48734,N_48911);
nor UO_2161 (O_2161,N_48132,N_49860);
and UO_2162 (O_2162,N_48268,N_48907);
and UO_2163 (O_2163,N_49900,N_48603);
or UO_2164 (O_2164,N_48068,N_49439);
nor UO_2165 (O_2165,N_48693,N_49696);
xnor UO_2166 (O_2166,N_48337,N_48988);
xor UO_2167 (O_2167,N_48044,N_48207);
and UO_2168 (O_2168,N_49616,N_48550);
and UO_2169 (O_2169,N_49539,N_48926);
nand UO_2170 (O_2170,N_49966,N_49050);
xor UO_2171 (O_2171,N_49530,N_48542);
or UO_2172 (O_2172,N_49473,N_48360);
or UO_2173 (O_2173,N_48014,N_49857);
nor UO_2174 (O_2174,N_48412,N_48612);
xnor UO_2175 (O_2175,N_49510,N_48830);
xnor UO_2176 (O_2176,N_48953,N_48418);
nand UO_2177 (O_2177,N_48179,N_49693);
nor UO_2178 (O_2178,N_48618,N_49244);
and UO_2179 (O_2179,N_48084,N_49571);
or UO_2180 (O_2180,N_49376,N_48625);
xor UO_2181 (O_2181,N_49534,N_49819);
and UO_2182 (O_2182,N_49705,N_49558);
nor UO_2183 (O_2183,N_49871,N_49295);
nor UO_2184 (O_2184,N_49142,N_48969);
nor UO_2185 (O_2185,N_49500,N_49065);
nor UO_2186 (O_2186,N_49627,N_48535);
nand UO_2187 (O_2187,N_48082,N_48318);
nor UO_2188 (O_2188,N_49242,N_49513);
nor UO_2189 (O_2189,N_48636,N_48677);
and UO_2190 (O_2190,N_49623,N_48119);
nor UO_2191 (O_2191,N_48547,N_49587);
nand UO_2192 (O_2192,N_48766,N_48914);
nor UO_2193 (O_2193,N_49926,N_49453);
and UO_2194 (O_2194,N_49571,N_49607);
and UO_2195 (O_2195,N_49078,N_48718);
nor UO_2196 (O_2196,N_48765,N_49075);
or UO_2197 (O_2197,N_49061,N_49357);
and UO_2198 (O_2198,N_48694,N_48822);
nor UO_2199 (O_2199,N_49165,N_48061);
nand UO_2200 (O_2200,N_48682,N_48553);
or UO_2201 (O_2201,N_48494,N_49211);
nor UO_2202 (O_2202,N_48216,N_49474);
and UO_2203 (O_2203,N_48520,N_49385);
nand UO_2204 (O_2204,N_49336,N_48565);
and UO_2205 (O_2205,N_48970,N_48502);
and UO_2206 (O_2206,N_48671,N_49248);
or UO_2207 (O_2207,N_49946,N_48225);
or UO_2208 (O_2208,N_49817,N_48941);
or UO_2209 (O_2209,N_49655,N_49984);
nand UO_2210 (O_2210,N_48883,N_49165);
or UO_2211 (O_2211,N_49865,N_49994);
or UO_2212 (O_2212,N_49130,N_49637);
xor UO_2213 (O_2213,N_48852,N_48381);
and UO_2214 (O_2214,N_49484,N_48796);
nand UO_2215 (O_2215,N_48090,N_49844);
nand UO_2216 (O_2216,N_48880,N_48868);
xnor UO_2217 (O_2217,N_48874,N_48120);
or UO_2218 (O_2218,N_48849,N_49381);
nand UO_2219 (O_2219,N_49230,N_49786);
nand UO_2220 (O_2220,N_49761,N_48656);
or UO_2221 (O_2221,N_48016,N_49182);
and UO_2222 (O_2222,N_48051,N_48130);
or UO_2223 (O_2223,N_49075,N_49230);
nor UO_2224 (O_2224,N_48407,N_49161);
nand UO_2225 (O_2225,N_49144,N_49339);
nor UO_2226 (O_2226,N_49867,N_48589);
nand UO_2227 (O_2227,N_48290,N_48810);
nor UO_2228 (O_2228,N_49197,N_48953);
nor UO_2229 (O_2229,N_48199,N_48901);
nor UO_2230 (O_2230,N_49977,N_49143);
nor UO_2231 (O_2231,N_48168,N_48221);
xnor UO_2232 (O_2232,N_48363,N_49863);
nor UO_2233 (O_2233,N_49304,N_48887);
xor UO_2234 (O_2234,N_49406,N_48518);
nor UO_2235 (O_2235,N_49026,N_48443);
or UO_2236 (O_2236,N_48772,N_48462);
nand UO_2237 (O_2237,N_49900,N_48412);
nor UO_2238 (O_2238,N_49437,N_48190);
nand UO_2239 (O_2239,N_49811,N_49181);
xnor UO_2240 (O_2240,N_49912,N_49564);
and UO_2241 (O_2241,N_49366,N_48459);
xnor UO_2242 (O_2242,N_48881,N_49338);
nor UO_2243 (O_2243,N_48306,N_49622);
xnor UO_2244 (O_2244,N_48748,N_48940);
nor UO_2245 (O_2245,N_49789,N_49250);
nand UO_2246 (O_2246,N_48792,N_48627);
or UO_2247 (O_2247,N_48893,N_48025);
xor UO_2248 (O_2248,N_49208,N_49892);
nand UO_2249 (O_2249,N_49948,N_48812);
xor UO_2250 (O_2250,N_48042,N_48560);
and UO_2251 (O_2251,N_49240,N_49477);
or UO_2252 (O_2252,N_48909,N_48491);
or UO_2253 (O_2253,N_49424,N_48647);
and UO_2254 (O_2254,N_49806,N_49171);
nand UO_2255 (O_2255,N_48904,N_48936);
or UO_2256 (O_2256,N_48771,N_49393);
and UO_2257 (O_2257,N_48024,N_49297);
xor UO_2258 (O_2258,N_48033,N_49563);
nor UO_2259 (O_2259,N_49403,N_48773);
and UO_2260 (O_2260,N_48323,N_48156);
xor UO_2261 (O_2261,N_48482,N_48297);
or UO_2262 (O_2262,N_48021,N_49434);
and UO_2263 (O_2263,N_48972,N_48281);
xnor UO_2264 (O_2264,N_49022,N_49795);
xor UO_2265 (O_2265,N_49072,N_49720);
nand UO_2266 (O_2266,N_49940,N_48277);
xor UO_2267 (O_2267,N_49609,N_49531);
nand UO_2268 (O_2268,N_48466,N_48971);
nand UO_2269 (O_2269,N_48387,N_48885);
nor UO_2270 (O_2270,N_48317,N_49239);
xnor UO_2271 (O_2271,N_49770,N_49196);
nor UO_2272 (O_2272,N_48663,N_48796);
and UO_2273 (O_2273,N_48413,N_48986);
nand UO_2274 (O_2274,N_49095,N_49917);
nand UO_2275 (O_2275,N_48428,N_49251);
xor UO_2276 (O_2276,N_49467,N_48449);
and UO_2277 (O_2277,N_49587,N_48530);
nand UO_2278 (O_2278,N_49572,N_48881);
nand UO_2279 (O_2279,N_48846,N_48516);
and UO_2280 (O_2280,N_48812,N_49861);
and UO_2281 (O_2281,N_49942,N_48709);
or UO_2282 (O_2282,N_48314,N_48032);
nand UO_2283 (O_2283,N_49793,N_48278);
or UO_2284 (O_2284,N_48595,N_49312);
or UO_2285 (O_2285,N_48233,N_48374);
and UO_2286 (O_2286,N_49209,N_48259);
and UO_2287 (O_2287,N_48487,N_48475);
or UO_2288 (O_2288,N_49627,N_48062);
xor UO_2289 (O_2289,N_48933,N_49634);
xor UO_2290 (O_2290,N_48601,N_48487);
nand UO_2291 (O_2291,N_49494,N_49686);
or UO_2292 (O_2292,N_49548,N_48604);
xor UO_2293 (O_2293,N_49810,N_49016);
nand UO_2294 (O_2294,N_49672,N_48892);
nand UO_2295 (O_2295,N_49874,N_49561);
xnor UO_2296 (O_2296,N_48841,N_48059);
and UO_2297 (O_2297,N_49199,N_49050);
nand UO_2298 (O_2298,N_49952,N_48642);
xnor UO_2299 (O_2299,N_49156,N_48735);
xor UO_2300 (O_2300,N_48854,N_48616);
or UO_2301 (O_2301,N_48372,N_48715);
xor UO_2302 (O_2302,N_49103,N_49417);
or UO_2303 (O_2303,N_48865,N_48690);
and UO_2304 (O_2304,N_49407,N_49024);
xnor UO_2305 (O_2305,N_48250,N_48582);
nor UO_2306 (O_2306,N_49325,N_49418);
xnor UO_2307 (O_2307,N_49110,N_48185);
or UO_2308 (O_2308,N_48569,N_49327);
and UO_2309 (O_2309,N_48131,N_49245);
nor UO_2310 (O_2310,N_48323,N_48218);
and UO_2311 (O_2311,N_49766,N_48714);
nand UO_2312 (O_2312,N_48363,N_48494);
nand UO_2313 (O_2313,N_48266,N_49704);
and UO_2314 (O_2314,N_48329,N_49670);
nand UO_2315 (O_2315,N_49945,N_48915);
xor UO_2316 (O_2316,N_48273,N_48034);
or UO_2317 (O_2317,N_49812,N_48424);
xor UO_2318 (O_2318,N_49434,N_48554);
nor UO_2319 (O_2319,N_49874,N_48197);
xnor UO_2320 (O_2320,N_48868,N_48820);
nor UO_2321 (O_2321,N_49399,N_49998);
or UO_2322 (O_2322,N_48250,N_48941);
and UO_2323 (O_2323,N_48228,N_48169);
or UO_2324 (O_2324,N_49341,N_48547);
and UO_2325 (O_2325,N_49242,N_49046);
xor UO_2326 (O_2326,N_48132,N_49474);
and UO_2327 (O_2327,N_49533,N_49148);
xor UO_2328 (O_2328,N_49066,N_49117);
xor UO_2329 (O_2329,N_49469,N_49411);
xor UO_2330 (O_2330,N_48557,N_49094);
and UO_2331 (O_2331,N_49244,N_49606);
nand UO_2332 (O_2332,N_49220,N_49051);
xor UO_2333 (O_2333,N_49995,N_49492);
or UO_2334 (O_2334,N_49353,N_48468);
and UO_2335 (O_2335,N_48111,N_48829);
nor UO_2336 (O_2336,N_48880,N_48336);
and UO_2337 (O_2337,N_48464,N_48422);
nor UO_2338 (O_2338,N_48109,N_48675);
and UO_2339 (O_2339,N_49863,N_48144);
or UO_2340 (O_2340,N_49893,N_49524);
or UO_2341 (O_2341,N_49530,N_48031);
nand UO_2342 (O_2342,N_49748,N_48862);
nand UO_2343 (O_2343,N_49247,N_49018);
and UO_2344 (O_2344,N_49202,N_49427);
xor UO_2345 (O_2345,N_48069,N_49266);
nand UO_2346 (O_2346,N_48448,N_48724);
nand UO_2347 (O_2347,N_48561,N_48078);
nor UO_2348 (O_2348,N_49074,N_48734);
xnor UO_2349 (O_2349,N_48307,N_49877);
and UO_2350 (O_2350,N_49267,N_48764);
and UO_2351 (O_2351,N_48090,N_49836);
xnor UO_2352 (O_2352,N_48615,N_48832);
or UO_2353 (O_2353,N_48121,N_49201);
xnor UO_2354 (O_2354,N_49900,N_49775);
nor UO_2355 (O_2355,N_48955,N_49071);
or UO_2356 (O_2356,N_49702,N_48853);
and UO_2357 (O_2357,N_49010,N_48656);
nand UO_2358 (O_2358,N_49884,N_49639);
nand UO_2359 (O_2359,N_48338,N_48141);
xnor UO_2360 (O_2360,N_48950,N_48884);
nand UO_2361 (O_2361,N_48731,N_48318);
or UO_2362 (O_2362,N_49311,N_48439);
or UO_2363 (O_2363,N_48886,N_49882);
nor UO_2364 (O_2364,N_48309,N_49093);
or UO_2365 (O_2365,N_49564,N_48052);
nand UO_2366 (O_2366,N_49012,N_49325);
and UO_2367 (O_2367,N_49114,N_49909);
and UO_2368 (O_2368,N_48379,N_48144);
and UO_2369 (O_2369,N_49018,N_49887);
and UO_2370 (O_2370,N_48946,N_48214);
and UO_2371 (O_2371,N_49227,N_48900);
xor UO_2372 (O_2372,N_49920,N_49689);
and UO_2373 (O_2373,N_48625,N_49482);
or UO_2374 (O_2374,N_49331,N_48792);
and UO_2375 (O_2375,N_49037,N_49359);
nand UO_2376 (O_2376,N_49750,N_49678);
nor UO_2377 (O_2377,N_49836,N_48913);
nor UO_2378 (O_2378,N_48746,N_48105);
xnor UO_2379 (O_2379,N_48300,N_48203);
and UO_2380 (O_2380,N_49330,N_48651);
or UO_2381 (O_2381,N_49406,N_49065);
or UO_2382 (O_2382,N_49566,N_49412);
and UO_2383 (O_2383,N_49701,N_49485);
nand UO_2384 (O_2384,N_48067,N_49227);
or UO_2385 (O_2385,N_48641,N_49874);
nand UO_2386 (O_2386,N_48967,N_48610);
xnor UO_2387 (O_2387,N_48346,N_48604);
nand UO_2388 (O_2388,N_48013,N_49214);
nor UO_2389 (O_2389,N_48473,N_48664);
nor UO_2390 (O_2390,N_49597,N_49820);
nor UO_2391 (O_2391,N_49300,N_48656);
or UO_2392 (O_2392,N_48444,N_49594);
and UO_2393 (O_2393,N_48956,N_48058);
nor UO_2394 (O_2394,N_49379,N_49224);
nand UO_2395 (O_2395,N_49552,N_48591);
and UO_2396 (O_2396,N_49786,N_48659);
nor UO_2397 (O_2397,N_49191,N_48867);
xnor UO_2398 (O_2398,N_48679,N_49567);
or UO_2399 (O_2399,N_48463,N_48178);
or UO_2400 (O_2400,N_48997,N_49033);
or UO_2401 (O_2401,N_48543,N_49140);
and UO_2402 (O_2402,N_49407,N_48794);
and UO_2403 (O_2403,N_48043,N_48207);
and UO_2404 (O_2404,N_49332,N_48877);
nor UO_2405 (O_2405,N_48630,N_49748);
nor UO_2406 (O_2406,N_49380,N_49740);
nand UO_2407 (O_2407,N_48153,N_49477);
and UO_2408 (O_2408,N_49274,N_48771);
nor UO_2409 (O_2409,N_48677,N_49871);
and UO_2410 (O_2410,N_48473,N_49887);
nor UO_2411 (O_2411,N_49206,N_49674);
nand UO_2412 (O_2412,N_49562,N_48129);
nand UO_2413 (O_2413,N_48944,N_49631);
or UO_2414 (O_2414,N_48398,N_49374);
or UO_2415 (O_2415,N_49866,N_48417);
xor UO_2416 (O_2416,N_48210,N_48237);
or UO_2417 (O_2417,N_49892,N_49495);
xnor UO_2418 (O_2418,N_49383,N_49738);
and UO_2419 (O_2419,N_48088,N_49968);
nor UO_2420 (O_2420,N_48364,N_48562);
xnor UO_2421 (O_2421,N_49154,N_49364);
nand UO_2422 (O_2422,N_48844,N_49147);
xor UO_2423 (O_2423,N_48619,N_48940);
xor UO_2424 (O_2424,N_49768,N_49233);
and UO_2425 (O_2425,N_49540,N_48214);
nor UO_2426 (O_2426,N_49672,N_48424);
or UO_2427 (O_2427,N_49643,N_49182);
nor UO_2428 (O_2428,N_48457,N_49264);
nor UO_2429 (O_2429,N_49233,N_48892);
xor UO_2430 (O_2430,N_49525,N_48459);
nor UO_2431 (O_2431,N_48776,N_48722);
nand UO_2432 (O_2432,N_49770,N_48044);
or UO_2433 (O_2433,N_48364,N_49815);
nor UO_2434 (O_2434,N_49428,N_49181);
nor UO_2435 (O_2435,N_48851,N_49466);
or UO_2436 (O_2436,N_48625,N_48730);
nor UO_2437 (O_2437,N_48993,N_49027);
nor UO_2438 (O_2438,N_49596,N_49024);
and UO_2439 (O_2439,N_48355,N_48403);
nor UO_2440 (O_2440,N_49882,N_48466);
or UO_2441 (O_2441,N_49182,N_48814);
xnor UO_2442 (O_2442,N_48353,N_48331);
or UO_2443 (O_2443,N_49611,N_48945);
and UO_2444 (O_2444,N_48960,N_49553);
and UO_2445 (O_2445,N_49882,N_48042);
or UO_2446 (O_2446,N_49713,N_49917);
or UO_2447 (O_2447,N_49868,N_49302);
and UO_2448 (O_2448,N_49480,N_49079);
and UO_2449 (O_2449,N_49849,N_48610);
or UO_2450 (O_2450,N_48752,N_48102);
or UO_2451 (O_2451,N_48146,N_48076);
xnor UO_2452 (O_2452,N_48761,N_49576);
nor UO_2453 (O_2453,N_49082,N_48496);
nand UO_2454 (O_2454,N_49591,N_49478);
or UO_2455 (O_2455,N_49482,N_48731);
nand UO_2456 (O_2456,N_48743,N_49505);
or UO_2457 (O_2457,N_49839,N_49709);
and UO_2458 (O_2458,N_49776,N_49587);
xnor UO_2459 (O_2459,N_49927,N_48247);
xor UO_2460 (O_2460,N_48785,N_48798);
or UO_2461 (O_2461,N_48088,N_48641);
nor UO_2462 (O_2462,N_49019,N_49867);
or UO_2463 (O_2463,N_48170,N_49085);
nand UO_2464 (O_2464,N_49627,N_48216);
nand UO_2465 (O_2465,N_48174,N_49904);
and UO_2466 (O_2466,N_48249,N_48255);
or UO_2467 (O_2467,N_48461,N_49751);
nor UO_2468 (O_2468,N_48774,N_48956);
or UO_2469 (O_2469,N_48180,N_48656);
or UO_2470 (O_2470,N_49065,N_48215);
and UO_2471 (O_2471,N_48557,N_48622);
nand UO_2472 (O_2472,N_48445,N_48700);
nor UO_2473 (O_2473,N_48462,N_49807);
nor UO_2474 (O_2474,N_48887,N_48639);
nor UO_2475 (O_2475,N_48699,N_49472);
or UO_2476 (O_2476,N_49080,N_48529);
nand UO_2477 (O_2477,N_49578,N_48010);
or UO_2478 (O_2478,N_48151,N_49532);
nor UO_2479 (O_2479,N_48839,N_48911);
and UO_2480 (O_2480,N_49674,N_48011);
or UO_2481 (O_2481,N_49025,N_49634);
and UO_2482 (O_2482,N_48678,N_48706);
nor UO_2483 (O_2483,N_49340,N_49362);
or UO_2484 (O_2484,N_49625,N_48464);
xnor UO_2485 (O_2485,N_48774,N_48812);
and UO_2486 (O_2486,N_49880,N_48179);
nand UO_2487 (O_2487,N_49362,N_49592);
or UO_2488 (O_2488,N_48619,N_48467);
nand UO_2489 (O_2489,N_48000,N_49079);
nand UO_2490 (O_2490,N_49719,N_48726);
nor UO_2491 (O_2491,N_49028,N_49008);
or UO_2492 (O_2492,N_48585,N_49354);
nor UO_2493 (O_2493,N_49777,N_48291);
nor UO_2494 (O_2494,N_49699,N_49151);
or UO_2495 (O_2495,N_49938,N_48510);
nand UO_2496 (O_2496,N_49641,N_48645);
nand UO_2497 (O_2497,N_48158,N_49371);
xor UO_2498 (O_2498,N_49613,N_48147);
and UO_2499 (O_2499,N_49415,N_49321);
nand UO_2500 (O_2500,N_48959,N_48044);
nand UO_2501 (O_2501,N_48229,N_48053);
and UO_2502 (O_2502,N_49945,N_49711);
xor UO_2503 (O_2503,N_48740,N_49685);
nor UO_2504 (O_2504,N_49994,N_48379);
nor UO_2505 (O_2505,N_49923,N_49548);
and UO_2506 (O_2506,N_48859,N_49169);
or UO_2507 (O_2507,N_48721,N_48256);
or UO_2508 (O_2508,N_49949,N_48181);
xor UO_2509 (O_2509,N_49673,N_49829);
xnor UO_2510 (O_2510,N_49877,N_48777);
nor UO_2511 (O_2511,N_49639,N_48940);
xnor UO_2512 (O_2512,N_49065,N_49368);
and UO_2513 (O_2513,N_48423,N_49418);
and UO_2514 (O_2514,N_49103,N_48661);
or UO_2515 (O_2515,N_48437,N_49281);
or UO_2516 (O_2516,N_48707,N_48401);
xor UO_2517 (O_2517,N_48938,N_49438);
xnor UO_2518 (O_2518,N_48929,N_48739);
xnor UO_2519 (O_2519,N_49280,N_49705);
nand UO_2520 (O_2520,N_49313,N_49601);
and UO_2521 (O_2521,N_49594,N_48042);
nor UO_2522 (O_2522,N_49097,N_49736);
and UO_2523 (O_2523,N_49226,N_48472);
nor UO_2524 (O_2524,N_48197,N_48078);
or UO_2525 (O_2525,N_49318,N_48442);
and UO_2526 (O_2526,N_49625,N_48063);
nor UO_2527 (O_2527,N_48721,N_48496);
and UO_2528 (O_2528,N_48938,N_49850);
nor UO_2529 (O_2529,N_48333,N_48959);
xor UO_2530 (O_2530,N_49314,N_49057);
nand UO_2531 (O_2531,N_48882,N_48486);
xnor UO_2532 (O_2532,N_49781,N_48175);
and UO_2533 (O_2533,N_48767,N_49938);
or UO_2534 (O_2534,N_48548,N_49501);
xnor UO_2535 (O_2535,N_48105,N_49601);
nand UO_2536 (O_2536,N_48613,N_49999);
xor UO_2537 (O_2537,N_49505,N_49328);
and UO_2538 (O_2538,N_48359,N_48091);
and UO_2539 (O_2539,N_48981,N_49342);
and UO_2540 (O_2540,N_49763,N_48534);
nand UO_2541 (O_2541,N_48327,N_49386);
nand UO_2542 (O_2542,N_48576,N_48984);
or UO_2543 (O_2543,N_48218,N_49960);
and UO_2544 (O_2544,N_49980,N_48451);
and UO_2545 (O_2545,N_49473,N_49521);
nor UO_2546 (O_2546,N_48667,N_48054);
and UO_2547 (O_2547,N_48860,N_48906);
nand UO_2548 (O_2548,N_48633,N_48667);
or UO_2549 (O_2549,N_49332,N_49786);
nand UO_2550 (O_2550,N_48715,N_48929);
or UO_2551 (O_2551,N_48094,N_48277);
nand UO_2552 (O_2552,N_48861,N_48249);
and UO_2553 (O_2553,N_48624,N_48063);
or UO_2554 (O_2554,N_48378,N_49214);
and UO_2555 (O_2555,N_49492,N_49507);
or UO_2556 (O_2556,N_49205,N_48882);
xor UO_2557 (O_2557,N_48414,N_49427);
xor UO_2558 (O_2558,N_49075,N_48546);
xnor UO_2559 (O_2559,N_49572,N_49478);
nand UO_2560 (O_2560,N_48573,N_49874);
xnor UO_2561 (O_2561,N_49797,N_48774);
nand UO_2562 (O_2562,N_49194,N_48987);
xnor UO_2563 (O_2563,N_49193,N_49214);
and UO_2564 (O_2564,N_49632,N_48115);
nand UO_2565 (O_2565,N_49682,N_49974);
or UO_2566 (O_2566,N_49750,N_48045);
and UO_2567 (O_2567,N_48553,N_49985);
nand UO_2568 (O_2568,N_48984,N_48608);
or UO_2569 (O_2569,N_48800,N_48940);
nor UO_2570 (O_2570,N_49984,N_48320);
nand UO_2571 (O_2571,N_48178,N_48291);
or UO_2572 (O_2572,N_48776,N_49828);
or UO_2573 (O_2573,N_49519,N_49368);
or UO_2574 (O_2574,N_49930,N_49220);
xor UO_2575 (O_2575,N_49030,N_48526);
xnor UO_2576 (O_2576,N_48954,N_49300);
or UO_2577 (O_2577,N_48820,N_49564);
xor UO_2578 (O_2578,N_49710,N_49946);
or UO_2579 (O_2579,N_48428,N_49425);
nor UO_2580 (O_2580,N_48126,N_48380);
nor UO_2581 (O_2581,N_48454,N_48585);
or UO_2582 (O_2582,N_48411,N_48158);
nand UO_2583 (O_2583,N_48636,N_48494);
nand UO_2584 (O_2584,N_48838,N_49372);
nor UO_2585 (O_2585,N_49997,N_48646);
or UO_2586 (O_2586,N_49485,N_48952);
xor UO_2587 (O_2587,N_48216,N_49462);
and UO_2588 (O_2588,N_49037,N_49960);
xnor UO_2589 (O_2589,N_48615,N_48538);
nand UO_2590 (O_2590,N_48576,N_49170);
and UO_2591 (O_2591,N_49645,N_48768);
and UO_2592 (O_2592,N_48571,N_48539);
nor UO_2593 (O_2593,N_49495,N_49035);
and UO_2594 (O_2594,N_49391,N_49488);
and UO_2595 (O_2595,N_48595,N_49408);
nand UO_2596 (O_2596,N_48369,N_49576);
nand UO_2597 (O_2597,N_48891,N_49402);
or UO_2598 (O_2598,N_49620,N_48281);
or UO_2599 (O_2599,N_48724,N_49868);
xor UO_2600 (O_2600,N_48973,N_48720);
and UO_2601 (O_2601,N_48246,N_49794);
nand UO_2602 (O_2602,N_49164,N_49223);
xor UO_2603 (O_2603,N_49814,N_49625);
and UO_2604 (O_2604,N_48659,N_48818);
nand UO_2605 (O_2605,N_49822,N_48237);
nor UO_2606 (O_2606,N_49843,N_48892);
xor UO_2607 (O_2607,N_48904,N_49986);
nor UO_2608 (O_2608,N_48831,N_48384);
nor UO_2609 (O_2609,N_49307,N_49105);
nor UO_2610 (O_2610,N_49021,N_49864);
xor UO_2611 (O_2611,N_49797,N_49741);
xor UO_2612 (O_2612,N_49974,N_49978);
nor UO_2613 (O_2613,N_49967,N_48427);
nand UO_2614 (O_2614,N_49095,N_48042);
nor UO_2615 (O_2615,N_48920,N_49524);
and UO_2616 (O_2616,N_49451,N_48614);
or UO_2617 (O_2617,N_48209,N_49742);
nand UO_2618 (O_2618,N_49415,N_48198);
or UO_2619 (O_2619,N_49901,N_48131);
nand UO_2620 (O_2620,N_49042,N_48266);
and UO_2621 (O_2621,N_48596,N_49398);
or UO_2622 (O_2622,N_49977,N_49771);
or UO_2623 (O_2623,N_48832,N_48117);
or UO_2624 (O_2624,N_49531,N_48458);
xor UO_2625 (O_2625,N_49528,N_48956);
nand UO_2626 (O_2626,N_48112,N_48631);
and UO_2627 (O_2627,N_48282,N_49596);
nor UO_2628 (O_2628,N_49816,N_49350);
or UO_2629 (O_2629,N_49705,N_48581);
or UO_2630 (O_2630,N_49306,N_48981);
and UO_2631 (O_2631,N_48125,N_49900);
nor UO_2632 (O_2632,N_49417,N_49474);
xor UO_2633 (O_2633,N_48395,N_49303);
xor UO_2634 (O_2634,N_49710,N_49059);
nor UO_2635 (O_2635,N_49652,N_48555);
nand UO_2636 (O_2636,N_48774,N_48201);
and UO_2637 (O_2637,N_49297,N_49167);
nand UO_2638 (O_2638,N_48237,N_49629);
and UO_2639 (O_2639,N_48132,N_48095);
xor UO_2640 (O_2640,N_48165,N_48464);
nor UO_2641 (O_2641,N_48522,N_49524);
xnor UO_2642 (O_2642,N_48527,N_48178);
nand UO_2643 (O_2643,N_49132,N_49400);
xor UO_2644 (O_2644,N_48344,N_49365);
and UO_2645 (O_2645,N_49350,N_48460);
xnor UO_2646 (O_2646,N_48996,N_49873);
nor UO_2647 (O_2647,N_48043,N_49281);
and UO_2648 (O_2648,N_49929,N_48833);
or UO_2649 (O_2649,N_48878,N_49437);
nor UO_2650 (O_2650,N_49856,N_49651);
or UO_2651 (O_2651,N_48623,N_48761);
or UO_2652 (O_2652,N_49103,N_48627);
nor UO_2653 (O_2653,N_48554,N_48261);
xor UO_2654 (O_2654,N_48924,N_49565);
and UO_2655 (O_2655,N_48493,N_48466);
nor UO_2656 (O_2656,N_48406,N_49185);
nand UO_2657 (O_2657,N_49415,N_48985);
nor UO_2658 (O_2658,N_49734,N_48051);
or UO_2659 (O_2659,N_48094,N_48333);
nand UO_2660 (O_2660,N_49917,N_48636);
xor UO_2661 (O_2661,N_48574,N_49190);
xnor UO_2662 (O_2662,N_48629,N_48218);
and UO_2663 (O_2663,N_49326,N_48020);
and UO_2664 (O_2664,N_49568,N_48150);
nand UO_2665 (O_2665,N_49112,N_48369);
nand UO_2666 (O_2666,N_48245,N_48277);
xnor UO_2667 (O_2667,N_48046,N_48079);
and UO_2668 (O_2668,N_48524,N_49384);
and UO_2669 (O_2669,N_49524,N_48953);
nand UO_2670 (O_2670,N_49114,N_48418);
nor UO_2671 (O_2671,N_48742,N_49783);
xnor UO_2672 (O_2672,N_49188,N_48518);
xor UO_2673 (O_2673,N_48286,N_48101);
xor UO_2674 (O_2674,N_49200,N_49333);
xnor UO_2675 (O_2675,N_48288,N_48823);
nand UO_2676 (O_2676,N_49848,N_48476);
nand UO_2677 (O_2677,N_49565,N_48846);
nor UO_2678 (O_2678,N_48415,N_49550);
nand UO_2679 (O_2679,N_48336,N_49141);
and UO_2680 (O_2680,N_49765,N_49578);
nand UO_2681 (O_2681,N_49702,N_48965);
or UO_2682 (O_2682,N_49188,N_48820);
or UO_2683 (O_2683,N_49028,N_48744);
xnor UO_2684 (O_2684,N_49542,N_48271);
or UO_2685 (O_2685,N_48367,N_48776);
or UO_2686 (O_2686,N_48867,N_48191);
nand UO_2687 (O_2687,N_48367,N_49150);
nor UO_2688 (O_2688,N_49139,N_49032);
nand UO_2689 (O_2689,N_49671,N_48516);
xnor UO_2690 (O_2690,N_49194,N_48855);
xor UO_2691 (O_2691,N_49085,N_48433);
nand UO_2692 (O_2692,N_49846,N_49518);
or UO_2693 (O_2693,N_48035,N_48621);
nor UO_2694 (O_2694,N_48253,N_48487);
nand UO_2695 (O_2695,N_49607,N_49698);
nand UO_2696 (O_2696,N_48197,N_49171);
xnor UO_2697 (O_2697,N_48846,N_48326);
and UO_2698 (O_2698,N_48953,N_48239);
and UO_2699 (O_2699,N_49576,N_49890);
and UO_2700 (O_2700,N_49525,N_48602);
nand UO_2701 (O_2701,N_48139,N_48975);
nand UO_2702 (O_2702,N_48526,N_49895);
and UO_2703 (O_2703,N_49404,N_49672);
and UO_2704 (O_2704,N_48657,N_49871);
and UO_2705 (O_2705,N_48114,N_48561);
nand UO_2706 (O_2706,N_49746,N_49975);
nor UO_2707 (O_2707,N_49372,N_48911);
nand UO_2708 (O_2708,N_49768,N_49343);
and UO_2709 (O_2709,N_48813,N_48937);
nor UO_2710 (O_2710,N_49945,N_49182);
xnor UO_2711 (O_2711,N_49898,N_49935);
xor UO_2712 (O_2712,N_48586,N_49451);
xnor UO_2713 (O_2713,N_48494,N_49663);
nor UO_2714 (O_2714,N_49640,N_48134);
nand UO_2715 (O_2715,N_49083,N_49024);
nand UO_2716 (O_2716,N_48306,N_49340);
xor UO_2717 (O_2717,N_48816,N_48235);
nor UO_2718 (O_2718,N_49866,N_49562);
xor UO_2719 (O_2719,N_49307,N_48274);
nand UO_2720 (O_2720,N_49181,N_48077);
xnor UO_2721 (O_2721,N_49551,N_48712);
nand UO_2722 (O_2722,N_48199,N_49646);
nand UO_2723 (O_2723,N_49241,N_49541);
or UO_2724 (O_2724,N_48504,N_48639);
or UO_2725 (O_2725,N_49097,N_48424);
xnor UO_2726 (O_2726,N_48296,N_48849);
nor UO_2727 (O_2727,N_49882,N_48102);
xnor UO_2728 (O_2728,N_49021,N_48811);
nand UO_2729 (O_2729,N_49098,N_49788);
nand UO_2730 (O_2730,N_48395,N_48440);
xnor UO_2731 (O_2731,N_48159,N_49350);
nor UO_2732 (O_2732,N_48305,N_49939);
nand UO_2733 (O_2733,N_49361,N_48175);
nand UO_2734 (O_2734,N_49629,N_48692);
nor UO_2735 (O_2735,N_49782,N_49130);
xor UO_2736 (O_2736,N_49676,N_49749);
xor UO_2737 (O_2737,N_49268,N_48239);
or UO_2738 (O_2738,N_49835,N_49413);
nand UO_2739 (O_2739,N_48236,N_49047);
nand UO_2740 (O_2740,N_48734,N_48128);
and UO_2741 (O_2741,N_48004,N_49477);
and UO_2742 (O_2742,N_49075,N_49092);
or UO_2743 (O_2743,N_48515,N_49299);
or UO_2744 (O_2744,N_49205,N_48177);
and UO_2745 (O_2745,N_49568,N_48411);
xor UO_2746 (O_2746,N_49844,N_49739);
and UO_2747 (O_2747,N_48409,N_48636);
nor UO_2748 (O_2748,N_48897,N_48887);
nand UO_2749 (O_2749,N_49549,N_48125);
xnor UO_2750 (O_2750,N_49934,N_48629);
and UO_2751 (O_2751,N_49919,N_49795);
and UO_2752 (O_2752,N_49360,N_49498);
xor UO_2753 (O_2753,N_49852,N_48523);
and UO_2754 (O_2754,N_49631,N_48158);
and UO_2755 (O_2755,N_49047,N_49698);
nor UO_2756 (O_2756,N_48794,N_49172);
or UO_2757 (O_2757,N_49557,N_49493);
nand UO_2758 (O_2758,N_48995,N_48864);
nand UO_2759 (O_2759,N_49609,N_48705);
xnor UO_2760 (O_2760,N_49582,N_48560);
and UO_2761 (O_2761,N_48413,N_48509);
xor UO_2762 (O_2762,N_48759,N_48709);
nor UO_2763 (O_2763,N_48359,N_49785);
or UO_2764 (O_2764,N_49401,N_48073);
nor UO_2765 (O_2765,N_49386,N_49049);
or UO_2766 (O_2766,N_49648,N_48328);
nor UO_2767 (O_2767,N_49563,N_49886);
nand UO_2768 (O_2768,N_49410,N_49309);
nor UO_2769 (O_2769,N_48718,N_48849);
and UO_2770 (O_2770,N_49608,N_48719);
nand UO_2771 (O_2771,N_49567,N_49319);
nor UO_2772 (O_2772,N_49258,N_49275);
nand UO_2773 (O_2773,N_48682,N_49186);
and UO_2774 (O_2774,N_48458,N_49692);
nand UO_2775 (O_2775,N_49553,N_48094);
xor UO_2776 (O_2776,N_49262,N_49490);
and UO_2777 (O_2777,N_48986,N_49328);
and UO_2778 (O_2778,N_49967,N_49724);
and UO_2779 (O_2779,N_49662,N_48099);
xor UO_2780 (O_2780,N_49999,N_49076);
nor UO_2781 (O_2781,N_49009,N_48857);
nand UO_2782 (O_2782,N_48853,N_49265);
and UO_2783 (O_2783,N_48085,N_49662);
or UO_2784 (O_2784,N_48487,N_49998);
and UO_2785 (O_2785,N_49252,N_49079);
nand UO_2786 (O_2786,N_49559,N_49131);
nand UO_2787 (O_2787,N_49157,N_49473);
and UO_2788 (O_2788,N_48935,N_48388);
or UO_2789 (O_2789,N_49770,N_49316);
and UO_2790 (O_2790,N_49992,N_49398);
and UO_2791 (O_2791,N_49002,N_49145);
or UO_2792 (O_2792,N_48851,N_48739);
xor UO_2793 (O_2793,N_48254,N_49639);
nor UO_2794 (O_2794,N_49141,N_49092);
or UO_2795 (O_2795,N_49022,N_48078);
nand UO_2796 (O_2796,N_49304,N_48434);
and UO_2797 (O_2797,N_49410,N_49745);
or UO_2798 (O_2798,N_49825,N_49025);
xnor UO_2799 (O_2799,N_48150,N_49229);
nor UO_2800 (O_2800,N_48274,N_49968);
nand UO_2801 (O_2801,N_48537,N_49029);
or UO_2802 (O_2802,N_48256,N_48804);
nand UO_2803 (O_2803,N_49984,N_48024);
and UO_2804 (O_2804,N_49598,N_49972);
nor UO_2805 (O_2805,N_49373,N_49337);
and UO_2806 (O_2806,N_48605,N_48593);
or UO_2807 (O_2807,N_49765,N_48759);
xor UO_2808 (O_2808,N_49579,N_48067);
xor UO_2809 (O_2809,N_48784,N_49848);
nand UO_2810 (O_2810,N_49541,N_48934);
xnor UO_2811 (O_2811,N_49395,N_48822);
nor UO_2812 (O_2812,N_48626,N_48555);
or UO_2813 (O_2813,N_48586,N_49578);
and UO_2814 (O_2814,N_48557,N_49748);
and UO_2815 (O_2815,N_49480,N_48353);
and UO_2816 (O_2816,N_49171,N_48936);
nor UO_2817 (O_2817,N_49774,N_48641);
or UO_2818 (O_2818,N_49338,N_49230);
xor UO_2819 (O_2819,N_48326,N_48348);
or UO_2820 (O_2820,N_49406,N_49021);
or UO_2821 (O_2821,N_49839,N_48392);
nand UO_2822 (O_2822,N_49528,N_48685);
nand UO_2823 (O_2823,N_49147,N_48144);
nor UO_2824 (O_2824,N_49420,N_48946);
nand UO_2825 (O_2825,N_48229,N_49495);
xor UO_2826 (O_2826,N_49766,N_48581);
nor UO_2827 (O_2827,N_48973,N_49884);
xor UO_2828 (O_2828,N_49293,N_48038);
xor UO_2829 (O_2829,N_49272,N_48170);
and UO_2830 (O_2830,N_49272,N_49043);
nand UO_2831 (O_2831,N_48944,N_48703);
or UO_2832 (O_2832,N_48893,N_48482);
nand UO_2833 (O_2833,N_49133,N_48313);
xnor UO_2834 (O_2834,N_49358,N_49894);
or UO_2835 (O_2835,N_49693,N_48739);
xnor UO_2836 (O_2836,N_49395,N_49208);
nand UO_2837 (O_2837,N_49991,N_49361);
or UO_2838 (O_2838,N_48603,N_48595);
or UO_2839 (O_2839,N_49220,N_49106);
nor UO_2840 (O_2840,N_48713,N_48305);
xnor UO_2841 (O_2841,N_49897,N_48093);
nor UO_2842 (O_2842,N_48369,N_49670);
nand UO_2843 (O_2843,N_49237,N_48372);
or UO_2844 (O_2844,N_49330,N_49243);
or UO_2845 (O_2845,N_49252,N_48649);
and UO_2846 (O_2846,N_48947,N_49473);
or UO_2847 (O_2847,N_48961,N_49032);
xnor UO_2848 (O_2848,N_49052,N_48902);
xor UO_2849 (O_2849,N_49662,N_49797);
nor UO_2850 (O_2850,N_48742,N_49565);
nor UO_2851 (O_2851,N_48013,N_48384);
nand UO_2852 (O_2852,N_48017,N_48231);
or UO_2853 (O_2853,N_48947,N_48138);
nand UO_2854 (O_2854,N_49550,N_49632);
nor UO_2855 (O_2855,N_49841,N_49693);
nand UO_2856 (O_2856,N_48108,N_48691);
and UO_2857 (O_2857,N_48511,N_49794);
and UO_2858 (O_2858,N_48765,N_48795);
xor UO_2859 (O_2859,N_48454,N_49399);
nor UO_2860 (O_2860,N_48432,N_49143);
nor UO_2861 (O_2861,N_48785,N_48386);
nor UO_2862 (O_2862,N_49605,N_48518);
xnor UO_2863 (O_2863,N_48033,N_49668);
nand UO_2864 (O_2864,N_48192,N_48313);
xnor UO_2865 (O_2865,N_48687,N_48215);
nor UO_2866 (O_2866,N_49910,N_49283);
and UO_2867 (O_2867,N_49978,N_48577);
xor UO_2868 (O_2868,N_49119,N_49980);
xnor UO_2869 (O_2869,N_48648,N_49978);
xor UO_2870 (O_2870,N_49619,N_49280);
nand UO_2871 (O_2871,N_49625,N_49556);
nor UO_2872 (O_2872,N_49937,N_48581);
nor UO_2873 (O_2873,N_48709,N_48323);
nor UO_2874 (O_2874,N_48422,N_48260);
nand UO_2875 (O_2875,N_48748,N_49172);
nand UO_2876 (O_2876,N_49900,N_48800);
and UO_2877 (O_2877,N_48421,N_48167);
nand UO_2878 (O_2878,N_49753,N_49168);
xor UO_2879 (O_2879,N_48997,N_48866);
or UO_2880 (O_2880,N_49754,N_49582);
and UO_2881 (O_2881,N_48247,N_48544);
nor UO_2882 (O_2882,N_49021,N_49140);
nand UO_2883 (O_2883,N_48801,N_49480);
xor UO_2884 (O_2884,N_49000,N_49758);
or UO_2885 (O_2885,N_48316,N_49683);
xnor UO_2886 (O_2886,N_49640,N_48340);
nand UO_2887 (O_2887,N_48019,N_49406);
xor UO_2888 (O_2888,N_49348,N_48709);
nand UO_2889 (O_2889,N_48573,N_49733);
nor UO_2890 (O_2890,N_48528,N_49103);
or UO_2891 (O_2891,N_49691,N_49510);
nor UO_2892 (O_2892,N_49698,N_48029);
xor UO_2893 (O_2893,N_49317,N_49339);
xor UO_2894 (O_2894,N_48999,N_49596);
nand UO_2895 (O_2895,N_49604,N_48605);
and UO_2896 (O_2896,N_48484,N_48448);
nor UO_2897 (O_2897,N_49311,N_48289);
xor UO_2898 (O_2898,N_48321,N_49113);
or UO_2899 (O_2899,N_49306,N_48458);
or UO_2900 (O_2900,N_49356,N_48167);
nor UO_2901 (O_2901,N_48520,N_49832);
or UO_2902 (O_2902,N_48771,N_49998);
nor UO_2903 (O_2903,N_49364,N_48491);
and UO_2904 (O_2904,N_48059,N_49570);
nand UO_2905 (O_2905,N_49418,N_48514);
nor UO_2906 (O_2906,N_48792,N_49594);
xnor UO_2907 (O_2907,N_49616,N_49581);
nand UO_2908 (O_2908,N_49111,N_48400);
nor UO_2909 (O_2909,N_48017,N_48979);
nor UO_2910 (O_2910,N_48656,N_49427);
nor UO_2911 (O_2911,N_48835,N_48966);
and UO_2912 (O_2912,N_48015,N_49608);
nand UO_2913 (O_2913,N_48655,N_49340);
nand UO_2914 (O_2914,N_48904,N_49263);
xor UO_2915 (O_2915,N_48539,N_48299);
xor UO_2916 (O_2916,N_48661,N_48956);
and UO_2917 (O_2917,N_49349,N_48990);
and UO_2918 (O_2918,N_49392,N_48684);
and UO_2919 (O_2919,N_49767,N_49307);
nor UO_2920 (O_2920,N_48462,N_49984);
xnor UO_2921 (O_2921,N_48331,N_49438);
nor UO_2922 (O_2922,N_48105,N_48306);
xor UO_2923 (O_2923,N_48471,N_48774);
nand UO_2924 (O_2924,N_49301,N_48629);
nand UO_2925 (O_2925,N_49935,N_48164);
or UO_2926 (O_2926,N_48292,N_48044);
xor UO_2927 (O_2927,N_48348,N_48627);
xnor UO_2928 (O_2928,N_48709,N_49819);
nor UO_2929 (O_2929,N_49586,N_48995);
nor UO_2930 (O_2930,N_49765,N_48141);
nor UO_2931 (O_2931,N_49235,N_48422);
and UO_2932 (O_2932,N_48674,N_48533);
and UO_2933 (O_2933,N_49915,N_48660);
xor UO_2934 (O_2934,N_49115,N_49277);
or UO_2935 (O_2935,N_49191,N_49328);
xor UO_2936 (O_2936,N_49883,N_48461);
and UO_2937 (O_2937,N_48016,N_49939);
or UO_2938 (O_2938,N_48419,N_49667);
nand UO_2939 (O_2939,N_48589,N_48194);
or UO_2940 (O_2940,N_48649,N_48633);
or UO_2941 (O_2941,N_48986,N_48947);
nand UO_2942 (O_2942,N_48944,N_49870);
and UO_2943 (O_2943,N_48746,N_49177);
and UO_2944 (O_2944,N_48694,N_49872);
or UO_2945 (O_2945,N_49433,N_49413);
xor UO_2946 (O_2946,N_49362,N_48713);
and UO_2947 (O_2947,N_49848,N_48218);
xor UO_2948 (O_2948,N_49106,N_48679);
nand UO_2949 (O_2949,N_48047,N_49431);
nand UO_2950 (O_2950,N_48865,N_48055);
nand UO_2951 (O_2951,N_48383,N_49189);
nor UO_2952 (O_2952,N_48338,N_49663);
xnor UO_2953 (O_2953,N_49716,N_48557);
xnor UO_2954 (O_2954,N_48785,N_49770);
xor UO_2955 (O_2955,N_49972,N_48003);
or UO_2956 (O_2956,N_48845,N_48394);
xor UO_2957 (O_2957,N_48625,N_48415);
and UO_2958 (O_2958,N_49127,N_48787);
nand UO_2959 (O_2959,N_48091,N_48613);
or UO_2960 (O_2960,N_49749,N_48228);
or UO_2961 (O_2961,N_48805,N_49814);
and UO_2962 (O_2962,N_49652,N_48563);
or UO_2963 (O_2963,N_49553,N_48947);
nor UO_2964 (O_2964,N_49567,N_49410);
xor UO_2965 (O_2965,N_48587,N_48717);
xor UO_2966 (O_2966,N_48699,N_49066);
nor UO_2967 (O_2967,N_49921,N_49745);
nor UO_2968 (O_2968,N_49041,N_49767);
xor UO_2969 (O_2969,N_49466,N_48573);
or UO_2970 (O_2970,N_49168,N_49984);
nand UO_2971 (O_2971,N_48668,N_48549);
nor UO_2972 (O_2972,N_48220,N_48091);
xor UO_2973 (O_2973,N_48448,N_48061);
nor UO_2974 (O_2974,N_48336,N_48536);
xor UO_2975 (O_2975,N_48823,N_48863);
xnor UO_2976 (O_2976,N_48034,N_48250);
or UO_2977 (O_2977,N_48983,N_49266);
nand UO_2978 (O_2978,N_49727,N_49045);
nor UO_2979 (O_2979,N_48136,N_49921);
nor UO_2980 (O_2980,N_48923,N_49719);
and UO_2981 (O_2981,N_49119,N_49599);
nand UO_2982 (O_2982,N_49714,N_49324);
nor UO_2983 (O_2983,N_48229,N_49114);
and UO_2984 (O_2984,N_49286,N_48138);
xor UO_2985 (O_2985,N_48762,N_49063);
nor UO_2986 (O_2986,N_48563,N_49524);
or UO_2987 (O_2987,N_48692,N_49506);
xor UO_2988 (O_2988,N_48380,N_48704);
or UO_2989 (O_2989,N_49168,N_48947);
and UO_2990 (O_2990,N_49241,N_49526);
and UO_2991 (O_2991,N_49693,N_49607);
nor UO_2992 (O_2992,N_48477,N_48460);
nor UO_2993 (O_2993,N_49498,N_48530);
nor UO_2994 (O_2994,N_49279,N_49366);
nand UO_2995 (O_2995,N_49423,N_49248);
nand UO_2996 (O_2996,N_48812,N_49111);
xnor UO_2997 (O_2997,N_48165,N_48146);
and UO_2998 (O_2998,N_48218,N_48808);
nand UO_2999 (O_2999,N_49610,N_49065);
xnor UO_3000 (O_3000,N_48176,N_49051);
and UO_3001 (O_3001,N_48101,N_48201);
nand UO_3002 (O_3002,N_48322,N_48508);
nor UO_3003 (O_3003,N_49700,N_49197);
nand UO_3004 (O_3004,N_48677,N_49405);
xnor UO_3005 (O_3005,N_49323,N_49229);
nor UO_3006 (O_3006,N_48726,N_48324);
nand UO_3007 (O_3007,N_49178,N_48376);
xor UO_3008 (O_3008,N_48008,N_49879);
nor UO_3009 (O_3009,N_48536,N_49830);
xnor UO_3010 (O_3010,N_48101,N_49260);
nand UO_3011 (O_3011,N_48350,N_49575);
or UO_3012 (O_3012,N_49771,N_48859);
xor UO_3013 (O_3013,N_49935,N_49406);
xnor UO_3014 (O_3014,N_48338,N_49333);
xor UO_3015 (O_3015,N_48971,N_49553);
and UO_3016 (O_3016,N_49047,N_48144);
nand UO_3017 (O_3017,N_49857,N_48698);
nor UO_3018 (O_3018,N_48133,N_49728);
or UO_3019 (O_3019,N_48885,N_48163);
xnor UO_3020 (O_3020,N_49815,N_48478);
and UO_3021 (O_3021,N_48192,N_49011);
xor UO_3022 (O_3022,N_48693,N_48736);
nand UO_3023 (O_3023,N_48552,N_48089);
or UO_3024 (O_3024,N_48542,N_48124);
nand UO_3025 (O_3025,N_48276,N_48589);
nand UO_3026 (O_3026,N_49754,N_48914);
xor UO_3027 (O_3027,N_48338,N_48490);
or UO_3028 (O_3028,N_49331,N_49363);
or UO_3029 (O_3029,N_48261,N_48296);
and UO_3030 (O_3030,N_48682,N_49959);
nor UO_3031 (O_3031,N_49069,N_48686);
or UO_3032 (O_3032,N_49744,N_49982);
and UO_3033 (O_3033,N_48025,N_49336);
nor UO_3034 (O_3034,N_48299,N_49558);
and UO_3035 (O_3035,N_49153,N_49180);
xnor UO_3036 (O_3036,N_48843,N_48483);
or UO_3037 (O_3037,N_48265,N_48864);
or UO_3038 (O_3038,N_49977,N_48678);
nand UO_3039 (O_3039,N_49961,N_48934);
xnor UO_3040 (O_3040,N_48606,N_48086);
or UO_3041 (O_3041,N_48448,N_48405);
nor UO_3042 (O_3042,N_48355,N_48760);
nor UO_3043 (O_3043,N_48621,N_49640);
nand UO_3044 (O_3044,N_49233,N_49870);
nand UO_3045 (O_3045,N_48542,N_48561);
or UO_3046 (O_3046,N_48898,N_48837);
nor UO_3047 (O_3047,N_48970,N_48389);
nand UO_3048 (O_3048,N_48407,N_49078);
nor UO_3049 (O_3049,N_48366,N_48152);
nand UO_3050 (O_3050,N_49828,N_49826);
and UO_3051 (O_3051,N_48374,N_49425);
nor UO_3052 (O_3052,N_49866,N_48617);
or UO_3053 (O_3053,N_48243,N_48658);
and UO_3054 (O_3054,N_48719,N_48175);
or UO_3055 (O_3055,N_49638,N_48472);
nand UO_3056 (O_3056,N_49066,N_49667);
nand UO_3057 (O_3057,N_49121,N_49187);
nand UO_3058 (O_3058,N_49647,N_49653);
or UO_3059 (O_3059,N_49969,N_49039);
xnor UO_3060 (O_3060,N_49942,N_48090);
nand UO_3061 (O_3061,N_48273,N_49286);
and UO_3062 (O_3062,N_48278,N_49875);
or UO_3063 (O_3063,N_49865,N_49570);
or UO_3064 (O_3064,N_48564,N_49630);
or UO_3065 (O_3065,N_49938,N_49256);
xor UO_3066 (O_3066,N_49813,N_48100);
xor UO_3067 (O_3067,N_48160,N_48289);
or UO_3068 (O_3068,N_49671,N_48930);
and UO_3069 (O_3069,N_48731,N_49726);
xor UO_3070 (O_3070,N_49769,N_48929);
nor UO_3071 (O_3071,N_48617,N_48538);
nand UO_3072 (O_3072,N_48942,N_48220);
xnor UO_3073 (O_3073,N_48010,N_49030);
xnor UO_3074 (O_3074,N_48059,N_48480);
and UO_3075 (O_3075,N_48865,N_48802);
nor UO_3076 (O_3076,N_49282,N_48389);
xor UO_3077 (O_3077,N_49367,N_49403);
or UO_3078 (O_3078,N_48444,N_49201);
or UO_3079 (O_3079,N_48693,N_48702);
nor UO_3080 (O_3080,N_49560,N_48719);
or UO_3081 (O_3081,N_49697,N_49698);
nor UO_3082 (O_3082,N_48806,N_49203);
nor UO_3083 (O_3083,N_48295,N_48219);
nor UO_3084 (O_3084,N_49995,N_48778);
or UO_3085 (O_3085,N_49297,N_49915);
xor UO_3086 (O_3086,N_48323,N_49631);
xor UO_3087 (O_3087,N_49525,N_49722);
nor UO_3088 (O_3088,N_48852,N_48569);
nand UO_3089 (O_3089,N_49340,N_49593);
nand UO_3090 (O_3090,N_49140,N_48237);
xnor UO_3091 (O_3091,N_48782,N_48318);
xor UO_3092 (O_3092,N_48073,N_48928);
or UO_3093 (O_3093,N_48110,N_49555);
and UO_3094 (O_3094,N_48924,N_49955);
xor UO_3095 (O_3095,N_48629,N_48178);
nor UO_3096 (O_3096,N_48132,N_49880);
or UO_3097 (O_3097,N_48793,N_49852);
xnor UO_3098 (O_3098,N_48940,N_48685);
nor UO_3099 (O_3099,N_48325,N_49801);
and UO_3100 (O_3100,N_49395,N_49228);
nand UO_3101 (O_3101,N_49005,N_49545);
or UO_3102 (O_3102,N_48880,N_49048);
xnor UO_3103 (O_3103,N_48120,N_48116);
xor UO_3104 (O_3104,N_49546,N_48641);
or UO_3105 (O_3105,N_49097,N_48850);
nand UO_3106 (O_3106,N_49006,N_48054);
nor UO_3107 (O_3107,N_48682,N_48257);
nor UO_3108 (O_3108,N_48167,N_48724);
and UO_3109 (O_3109,N_48651,N_48150);
xnor UO_3110 (O_3110,N_49132,N_48528);
xnor UO_3111 (O_3111,N_49550,N_48111);
or UO_3112 (O_3112,N_49395,N_49935);
xnor UO_3113 (O_3113,N_48172,N_49260);
xor UO_3114 (O_3114,N_48530,N_48610);
xor UO_3115 (O_3115,N_48577,N_48955);
xnor UO_3116 (O_3116,N_48430,N_49516);
nor UO_3117 (O_3117,N_48826,N_48462);
and UO_3118 (O_3118,N_49370,N_48773);
nor UO_3119 (O_3119,N_49268,N_49218);
xnor UO_3120 (O_3120,N_48262,N_48276);
nor UO_3121 (O_3121,N_49082,N_49390);
xnor UO_3122 (O_3122,N_49900,N_49020);
nand UO_3123 (O_3123,N_48621,N_48029);
nand UO_3124 (O_3124,N_49808,N_49653);
or UO_3125 (O_3125,N_49161,N_48005);
nor UO_3126 (O_3126,N_48469,N_49251);
and UO_3127 (O_3127,N_49329,N_48930);
nand UO_3128 (O_3128,N_48229,N_49606);
nand UO_3129 (O_3129,N_48523,N_49624);
nor UO_3130 (O_3130,N_48274,N_48506);
nand UO_3131 (O_3131,N_49523,N_49334);
and UO_3132 (O_3132,N_49831,N_49582);
xor UO_3133 (O_3133,N_48691,N_49801);
nand UO_3134 (O_3134,N_48249,N_48480);
or UO_3135 (O_3135,N_49056,N_48329);
and UO_3136 (O_3136,N_49791,N_49977);
xor UO_3137 (O_3137,N_48287,N_48383);
xnor UO_3138 (O_3138,N_49714,N_49265);
xnor UO_3139 (O_3139,N_49803,N_49478);
and UO_3140 (O_3140,N_49368,N_49847);
xor UO_3141 (O_3141,N_49191,N_49983);
nor UO_3142 (O_3142,N_49993,N_49584);
nor UO_3143 (O_3143,N_48802,N_48112);
xnor UO_3144 (O_3144,N_49877,N_48273);
or UO_3145 (O_3145,N_48688,N_49651);
or UO_3146 (O_3146,N_49341,N_49026);
nor UO_3147 (O_3147,N_48408,N_48537);
or UO_3148 (O_3148,N_48152,N_48197);
nor UO_3149 (O_3149,N_49877,N_48595);
nor UO_3150 (O_3150,N_49700,N_48503);
nand UO_3151 (O_3151,N_48392,N_49439);
or UO_3152 (O_3152,N_49273,N_49090);
xor UO_3153 (O_3153,N_49501,N_49426);
nor UO_3154 (O_3154,N_49815,N_48357);
or UO_3155 (O_3155,N_49825,N_48979);
nor UO_3156 (O_3156,N_48420,N_49277);
and UO_3157 (O_3157,N_48819,N_48271);
nor UO_3158 (O_3158,N_49190,N_48065);
and UO_3159 (O_3159,N_48037,N_48994);
nor UO_3160 (O_3160,N_49875,N_48196);
nand UO_3161 (O_3161,N_49973,N_49902);
nand UO_3162 (O_3162,N_49776,N_49736);
nand UO_3163 (O_3163,N_49684,N_48073);
nor UO_3164 (O_3164,N_48525,N_49224);
nor UO_3165 (O_3165,N_48238,N_49164);
nand UO_3166 (O_3166,N_49106,N_49319);
xnor UO_3167 (O_3167,N_49364,N_49007);
nand UO_3168 (O_3168,N_49229,N_48340);
nand UO_3169 (O_3169,N_48625,N_49397);
nand UO_3170 (O_3170,N_49004,N_49268);
xnor UO_3171 (O_3171,N_48645,N_49936);
and UO_3172 (O_3172,N_48825,N_48080);
nand UO_3173 (O_3173,N_48638,N_48760);
nand UO_3174 (O_3174,N_48664,N_48649);
and UO_3175 (O_3175,N_48171,N_48052);
or UO_3176 (O_3176,N_48131,N_49858);
and UO_3177 (O_3177,N_49206,N_48267);
or UO_3178 (O_3178,N_48035,N_48597);
or UO_3179 (O_3179,N_49920,N_49669);
nor UO_3180 (O_3180,N_48875,N_48815);
or UO_3181 (O_3181,N_48917,N_48476);
xor UO_3182 (O_3182,N_48751,N_49485);
nor UO_3183 (O_3183,N_49622,N_48735);
xnor UO_3184 (O_3184,N_48079,N_48795);
and UO_3185 (O_3185,N_49316,N_48375);
nand UO_3186 (O_3186,N_49376,N_48908);
or UO_3187 (O_3187,N_48839,N_49879);
nand UO_3188 (O_3188,N_48489,N_48556);
or UO_3189 (O_3189,N_48135,N_49064);
nor UO_3190 (O_3190,N_49242,N_49722);
and UO_3191 (O_3191,N_48704,N_49841);
xnor UO_3192 (O_3192,N_49394,N_49036);
nor UO_3193 (O_3193,N_49411,N_48068);
or UO_3194 (O_3194,N_49640,N_49347);
or UO_3195 (O_3195,N_49406,N_49297);
or UO_3196 (O_3196,N_49559,N_48261);
xnor UO_3197 (O_3197,N_49453,N_48402);
nor UO_3198 (O_3198,N_49694,N_49138);
nor UO_3199 (O_3199,N_48561,N_49007);
xor UO_3200 (O_3200,N_49427,N_49280);
or UO_3201 (O_3201,N_48063,N_48847);
or UO_3202 (O_3202,N_49511,N_48757);
nand UO_3203 (O_3203,N_48596,N_49301);
and UO_3204 (O_3204,N_49237,N_49594);
or UO_3205 (O_3205,N_48671,N_48037);
xnor UO_3206 (O_3206,N_48584,N_49199);
nor UO_3207 (O_3207,N_48107,N_48751);
nor UO_3208 (O_3208,N_48590,N_49734);
nor UO_3209 (O_3209,N_49588,N_49526);
and UO_3210 (O_3210,N_49915,N_48545);
xor UO_3211 (O_3211,N_48324,N_49356);
and UO_3212 (O_3212,N_48025,N_49214);
nor UO_3213 (O_3213,N_49637,N_49048);
nor UO_3214 (O_3214,N_49643,N_49090);
or UO_3215 (O_3215,N_49070,N_48472);
nand UO_3216 (O_3216,N_48027,N_48162);
and UO_3217 (O_3217,N_48107,N_48281);
and UO_3218 (O_3218,N_48796,N_48031);
nand UO_3219 (O_3219,N_49687,N_49503);
xnor UO_3220 (O_3220,N_49734,N_48168);
and UO_3221 (O_3221,N_48979,N_49333);
nand UO_3222 (O_3222,N_48748,N_48146);
xor UO_3223 (O_3223,N_48145,N_48602);
nand UO_3224 (O_3224,N_49123,N_48827);
and UO_3225 (O_3225,N_48205,N_48000);
or UO_3226 (O_3226,N_48197,N_49875);
xor UO_3227 (O_3227,N_48745,N_48764);
or UO_3228 (O_3228,N_49191,N_49511);
nand UO_3229 (O_3229,N_49688,N_48795);
or UO_3230 (O_3230,N_49114,N_48581);
xnor UO_3231 (O_3231,N_49853,N_49255);
or UO_3232 (O_3232,N_49272,N_49122);
or UO_3233 (O_3233,N_49866,N_49016);
nand UO_3234 (O_3234,N_49968,N_49426);
or UO_3235 (O_3235,N_49860,N_49324);
nor UO_3236 (O_3236,N_48396,N_49029);
xor UO_3237 (O_3237,N_49882,N_49606);
nor UO_3238 (O_3238,N_48751,N_49581);
xor UO_3239 (O_3239,N_49491,N_48618);
xor UO_3240 (O_3240,N_49503,N_49122);
nand UO_3241 (O_3241,N_48317,N_48612);
and UO_3242 (O_3242,N_48697,N_49941);
nand UO_3243 (O_3243,N_48275,N_48036);
or UO_3244 (O_3244,N_49375,N_48583);
or UO_3245 (O_3245,N_48597,N_48919);
xor UO_3246 (O_3246,N_48346,N_49284);
xor UO_3247 (O_3247,N_48748,N_48191);
and UO_3248 (O_3248,N_48110,N_49691);
or UO_3249 (O_3249,N_49860,N_48735);
nor UO_3250 (O_3250,N_48944,N_49539);
xor UO_3251 (O_3251,N_48616,N_49109);
and UO_3252 (O_3252,N_48705,N_48567);
xor UO_3253 (O_3253,N_49930,N_48549);
nand UO_3254 (O_3254,N_48120,N_48172);
and UO_3255 (O_3255,N_49675,N_48011);
xor UO_3256 (O_3256,N_48709,N_49184);
nand UO_3257 (O_3257,N_48750,N_49541);
and UO_3258 (O_3258,N_48527,N_48433);
or UO_3259 (O_3259,N_48008,N_48861);
xnor UO_3260 (O_3260,N_48322,N_48005);
and UO_3261 (O_3261,N_48277,N_48212);
xnor UO_3262 (O_3262,N_48847,N_48851);
or UO_3263 (O_3263,N_49432,N_48240);
nand UO_3264 (O_3264,N_49373,N_49911);
and UO_3265 (O_3265,N_48937,N_48481);
or UO_3266 (O_3266,N_49225,N_48261);
or UO_3267 (O_3267,N_49387,N_49652);
or UO_3268 (O_3268,N_48026,N_48110);
nand UO_3269 (O_3269,N_49701,N_49410);
or UO_3270 (O_3270,N_48625,N_49102);
and UO_3271 (O_3271,N_48352,N_48311);
nand UO_3272 (O_3272,N_48871,N_49169);
nor UO_3273 (O_3273,N_48368,N_49607);
nand UO_3274 (O_3274,N_48216,N_49238);
nand UO_3275 (O_3275,N_48184,N_48002);
nand UO_3276 (O_3276,N_48147,N_48502);
nand UO_3277 (O_3277,N_49352,N_48522);
and UO_3278 (O_3278,N_49713,N_48492);
or UO_3279 (O_3279,N_48356,N_48365);
xnor UO_3280 (O_3280,N_48389,N_49642);
and UO_3281 (O_3281,N_48976,N_48865);
and UO_3282 (O_3282,N_48432,N_48007);
and UO_3283 (O_3283,N_49360,N_49576);
or UO_3284 (O_3284,N_49487,N_49091);
or UO_3285 (O_3285,N_48634,N_48322);
nand UO_3286 (O_3286,N_48177,N_49319);
nand UO_3287 (O_3287,N_48865,N_48529);
or UO_3288 (O_3288,N_48391,N_49948);
and UO_3289 (O_3289,N_48376,N_49773);
nor UO_3290 (O_3290,N_49764,N_49732);
nand UO_3291 (O_3291,N_48485,N_49242);
or UO_3292 (O_3292,N_48426,N_49445);
nor UO_3293 (O_3293,N_48149,N_49320);
nor UO_3294 (O_3294,N_49230,N_49260);
xnor UO_3295 (O_3295,N_49057,N_48227);
or UO_3296 (O_3296,N_49410,N_48797);
or UO_3297 (O_3297,N_49771,N_49176);
nand UO_3298 (O_3298,N_49501,N_49456);
and UO_3299 (O_3299,N_49546,N_48394);
and UO_3300 (O_3300,N_49823,N_49769);
xor UO_3301 (O_3301,N_48459,N_49596);
or UO_3302 (O_3302,N_48590,N_49580);
or UO_3303 (O_3303,N_48187,N_48160);
or UO_3304 (O_3304,N_49230,N_49917);
and UO_3305 (O_3305,N_49476,N_49937);
or UO_3306 (O_3306,N_49017,N_49037);
nor UO_3307 (O_3307,N_48931,N_48331);
nand UO_3308 (O_3308,N_49765,N_48223);
xor UO_3309 (O_3309,N_49495,N_48539);
xor UO_3310 (O_3310,N_49732,N_48563);
xnor UO_3311 (O_3311,N_48852,N_49400);
nor UO_3312 (O_3312,N_48171,N_48639);
and UO_3313 (O_3313,N_48549,N_49111);
or UO_3314 (O_3314,N_48959,N_48193);
nand UO_3315 (O_3315,N_48631,N_49067);
nand UO_3316 (O_3316,N_49860,N_49545);
or UO_3317 (O_3317,N_48410,N_48110);
nor UO_3318 (O_3318,N_48648,N_48952);
nor UO_3319 (O_3319,N_48630,N_48893);
xor UO_3320 (O_3320,N_49108,N_49404);
nor UO_3321 (O_3321,N_48952,N_48984);
xor UO_3322 (O_3322,N_48500,N_48214);
xor UO_3323 (O_3323,N_49635,N_49310);
or UO_3324 (O_3324,N_49744,N_48055);
xor UO_3325 (O_3325,N_49780,N_48550);
nor UO_3326 (O_3326,N_48304,N_49041);
xor UO_3327 (O_3327,N_48769,N_49314);
nor UO_3328 (O_3328,N_48993,N_49945);
nor UO_3329 (O_3329,N_48668,N_48025);
and UO_3330 (O_3330,N_48543,N_49396);
nand UO_3331 (O_3331,N_48345,N_48513);
and UO_3332 (O_3332,N_49896,N_49959);
nand UO_3333 (O_3333,N_48198,N_49567);
nor UO_3334 (O_3334,N_49304,N_48046);
and UO_3335 (O_3335,N_48490,N_48002);
xnor UO_3336 (O_3336,N_49252,N_49658);
nor UO_3337 (O_3337,N_49103,N_48968);
or UO_3338 (O_3338,N_49873,N_49238);
nor UO_3339 (O_3339,N_49452,N_48625);
nor UO_3340 (O_3340,N_49900,N_49948);
or UO_3341 (O_3341,N_49800,N_49580);
and UO_3342 (O_3342,N_48342,N_49858);
nand UO_3343 (O_3343,N_48669,N_48351);
nand UO_3344 (O_3344,N_48948,N_48501);
nand UO_3345 (O_3345,N_49173,N_49687);
nor UO_3346 (O_3346,N_48712,N_49773);
nor UO_3347 (O_3347,N_48747,N_49477);
or UO_3348 (O_3348,N_49425,N_49102);
nor UO_3349 (O_3349,N_48955,N_49966);
or UO_3350 (O_3350,N_48272,N_49097);
xor UO_3351 (O_3351,N_49468,N_48148);
nor UO_3352 (O_3352,N_48182,N_48083);
nor UO_3353 (O_3353,N_49497,N_48110);
or UO_3354 (O_3354,N_48870,N_49330);
and UO_3355 (O_3355,N_49283,N_49522);
nor UO_3356 (O_3356,N_49336,N_48723);
or UO_3357 (O_3357,N_48821,N_48970);
xnor UO_3358 (O_3358,N_48105,N_49928);
or UO_3359 (O_3359,N_48934,N_48487);
nand UO_3360 (O_3360,N_49915,N_49527);
and UO_3361 (O_3361,N_48722,N_48130);
nand UO_3362 (O_3362,N_49366,N_48707);
and UO_3363 (O_3363,N_48257,N_48467);
nor UO_3364 (O_3364,N_49913,N_48299);
nand UO_3365 (O_3365,N_48141,N_49650);
and UO_3366 (O_3366,N_49965,N_49913);
and UO_3367 (O_3367,N_49171,N_49282);
nor UO_3368 (O_3368,N_48384,N_49705);
nor UO_3369 (O_3369,N_48506,N_48286);
nand UO_3370 (O_3370,N_49818,N_48167);
and UO_3371 (O_3371,N_49242,N_48215);
xor UO_3372 (O_3372,N_49747,N_49426);
or UO_3373 (O_3373,N_49141,N_48334);
and UO_3374 (O_3374,N_48950,N_48179);
nand UO_3375 (O_3375,N_48439,N_49986);
nor UO_3376 (O_3376,N_48679,N_48036);
or UO_3377 (O_3377,N_48374,N_48995);
or UO_3378 (O_3378,N_49712,N_49838);
and UO_3379 (O_3379,N_49022,N_48432);
and UO_3380 (O_3380,N_49160,N_48657);
nor UO_3381 (O_3381,N_49765,N_49349);
or UO_3382 (O_3382,N_48780,N_48978);
xnor UO_3383 (O_3383,N_48452,N_48664);
xor UO_3384 (O_3384,N_49903,N_49506);
and UO_3385 (O_3385,N_48832,N_49886);
nor UO_3386 (O_3386,N_48394,N_49386);
nand UO_3387 (O_3387,N_49160,N_48216);
and UO_3388 (O_3388,N_48862,N_48425);
nor UO_3389 (O_3389,N_49057,N_49917);
nand UO_3390 (O_3390,N_48628,N_48380);
and UO_3391 (O_3391,N_49845,N_48641);
nor UO_3392 (O_3392,N_49372,N_49279);
and UO_3393 (O_3393,N_48164,N_49986);
nor UO_3394 (O_3394,N_48688,N_48612);
xor UO_3395 (O_3395,N_49319,N_48715);
and UO_3396 (O_3396,N_49526,N_48533);
or UO_3397 (O_3397,N_49858,N_49074);
or UO_3398 (O_3398,N_48159,N_49917);
nand UO_3399 (O_3399,N_48193,N_48405);
xor UO_3400 (O_3400,N_49206,N_49987);
or UO_3401 (O_3401,N_48171,N_48816);
nand UO_3402 (O_3402,N_48362,N_48965);
or UO_3403 (O_3403,N_48362,N_48676);
or UO_3404 (O_3404,N_49200,N_48805);
xor UO_3405 (O_3405,N_48562,N_48539);
or UO_3406 (O_3406,N_49636,N_48850);
nand UO_3407 (O_3407,N_49989,N_48003);
and UO_3408 (O_3408,N_49290,N_49546);
and UO_3409 (O_3409,N_48683,N_49984);
or UO_3410 (O_3410,N_49455,N_49225);
or UO_3411 (O_3411,N_49045,N_49235);
xor UO_3412 (O_3412,N_48438,N_49954);
nor UO_3413 (O_3413,N_48668,N_49233);
or UO_3414 (O_3414,N_48306,N_49477);
xor UO_3415 (O_3415,N_48724,N_49645);
nand UO_3416 (O_3416,N_49798,N_49786);
xnor UO_3417 (O_3417,N_48014,N_49889);
nor UO_3418 (O_3418,N_48566,N_48127);
and UO_3419 (O_3419,N_49997,N_49753);
nand UO_3420 (O_3420,N_48769,N_49712);
and UO_3421 (O_3421,N_49949,N_49020);
nand UO_3422 (O_3422,N_48643,N_48801);
nor UO_3423 (O_3423,N_48514,N_48287);
xnor UO_3424 (O_3424,N_48468,N_48662);
or UO_3425 (O_3425,N_48871,N_49137);
or UO_3426 (O_3426,N_48044,N_48391);
xnor UO_3427 (O_3427,N_48182,N_48937);
and UO_3428 (O_3428,N_48115,N_48748);
or UO_3429 (O_3429,N_49121,N_49655);
nor UO_3430 (O_3430,N_48353,N_49510);
nor UO_3431 (O_3431,N_49633,N_48024);
xnor UO_3432 (O_3432,N_49072,N_49785);
nor UO_3433 (O_3433,N_48444,N_49705);
nand UO_3434 (O_3434,N_48232,N_48500);
and UO_3435 (O_3435,N_49018,N_49677);
or UO_3436 (O_3436,N_49956,N_48384);
nor UO_3437 (O_3437,N_49010,N_48779);
or UO_3438 (O_3438,N_49173,N_48506);
or UO_3439 (O_3439,N_49484,N_48513);
and UO_3440 (O_3440,N_49589,N_48099);
xnor UO_3441 (O_3441,N_48266,N_49195);
xnor UO_3442 (O_3442,N_48678,N_48658);
or UO_3443 (O_3443,N_48898,N_48187);
and UO_3444 (O_3444,N_49691,N_48621);
nand UO_3445 (O_3445,N_49530,N_49177);
nand UO_3446 (O_3446,N_48822,N_48315);
or UO_3447 (O_3447,N_49273,N_49646);
nor UO_3448 (O_3448,N_49592,N_48595);
and UO_3449 (O_3449,N_48210,N_49218);
nand UO_3450 (O_3450,N_49584,N_48601);
nor UO_3451 (O_3451,N_48416,N_48457);
nand UO_3452 (O_3452,N_49966,N_49156);
nor UO_3453 (O_3453,N_48157,N_49437);
nand UO_3454 (O_3454,N_49690,N_48158);
and UO_3455 (O_3455,N_48317,N_49578);
and UO_3456 (O_3456,N_48693,N_48887);
xor UO_3457 (O_3457,N_49763,N_48545);
nand UO_3458 (O_3458,N_49207,N_48575);
or UO_3459 (O_3459,N_49611,N_48266);
nor UO_3460 (O_3460,N_49569,N_48991);
nand UO_3461 (O_3461,N_48173,N_49325);
xor UO_3462 (O_3462,N_48347,N_49013);
or UO_3463 (O_3463,N_48952,N_49860);
nand UO_3464 (O_3464,N_48981,N_49557);
or UO_3465 (O_3465,N_49433,N_49938);
and UO_3466 (O_3466,N_48467,N_48138);
nor UO_3467 (O_3467,N_49938,N_49961);
nand UO_3468 (O_3468,N_49268,N_49352);
nor UO_3469 (O_3469,N_48425,N_48204);
and UO_3470 (O_3470,N_49722,N_49299);
nor UO_3471 (O_3471,N_49889,N_49157);
nand UO_3472 (O_3472,N_48462,N_49862);
xor UO_3473 (O_3473,N_49970,N_48573);
or UO_3474 (O_3474,N_49837,N_48530);
xor UO_3475 (O_3475,N_48327,N_48025);
nand UO_3476 (O_3476,N_49887,N_48074);
nand UO_3477 (O_3477,N_48342,N_48925);
nor UO_3478 (O_3478,N_49037,N_48136);
nor UO_3479 (O_3479,N_49524,N_49498);
nand UO_3480 (O_3480,N_49581,N_48774);
nor UO_3481 (O_3481,N_49002,N_49054);
nand UO_3482 (O_3482,N_49080,N_48257);
nand UO_3483 (O_3483,N_49504,N_48806);
nand UO_3484 (O_3484,N_48504,N_48511);
or UO_3485 (O_3485,N_48806,N_49079);
xnor UO_3486 (O_3486,N_49025,N_49966);
xnor UO_3487 (O_3487,N_49356,N_49024);
nor UO_3488 (O_3488,N_49607,N_48783);
nand UO_3489 (O_3489,N_49703,N_48924);
nor UO_3490 (O_3490,N_49032,N_48356);
or UO_3491 (O_3491,N_48977,N_48262);
nor UO_3492 (O_3492,N_48386,N_48727);
or UO_3493 (O_3493,N_48416,N_49918);
nor UO_3494 (O_3494,N_48716,N_48636);
xor UO_3495 (O_3495,N_48734,N_49100);
xnor UO_3496 (O_3496,N_49776,N_48181);
and UO_3497 (O_3497,N_49016,N_48711);
nand UO_3498 (O_3498,N_49290,N_48150);
or UO_3499 (O_3499,N_48094,N_49772);
or UO_3500 (O_3500,N_48937,N_48948);
xnor UO_3501 (O_3501,N_49100,N_48784);
xnor UO_3502 (O_3502,N_49345,N_48145);
or UO_3503 (O_3503,N_48865,N_48518);
nor UO_3504 (O_3504,N_48791,N_49155);
nor UO_3505 (O_3505,N_49824,N_49791);
nor UO_3506 (O_3506,N_49521,N_48224);
xnor UO_3507 (O_3507,N_49911,N_48809);
or UO_3508 (O_3508,N_48333,N_48575);
nand UO_3509 (O_3509,N_48971,N_48270);
xor UO_3510 (O_3510,N_48301,N_49137);
and UO_3511 (O_3511,N_48006,N_48546);
or UO_3512 (O_3512,N_48352,N_49520);
nor UO_3513 (O_3513,N_49978,N_48746);
nor UO_3514 (O_3514,N_49836,N_49837);
xnor UO_3515 (O_3515,N_48794,N_49505);
nand UO_3516 (O_3516,N_48324,N_48298);
and UO_3517 (O_3517,N_49890,N_49462);
xor UO_3518 (O_3518,N_49310,N_49178);
nand UO_3519 (O_3519,N_49281,N_49121);
xor UO_3520 (O_3520,N_48567,N_49444);
and UO_3521 (O_3521,N_48328,N_49787);
nand UO_3522 (O_3522,N_49076,N_49297);
or UO_3523 (O_3523,N_49728,N_49260);
nor UO_3524 (O_3524,N_48405,N_48036);
and UO_3525 (O_3525,N_48745,N_48217);
nand UO_3526 (O_3526,N_48703,N_49412);
xnor UO_3527 (O_3527,N_48459,N_48947);
xor UO_3528 (O_3528,N_48609,N_49844);
nand UO_3529 (O_3529,N_48205,N_49100);
nor UO_3530 (O_3530,N_48458,N_48775);
nand UO_3531 (O_3531,N_48133,N_49241);
nor UO_3532 (O_3532,N_48406,N_49524);
nand UO_3533 (O_3533,N_48681,N_48213);
nand UO_3534 (O_3534,N_48132,N_48235);
xnor UO_3535 (O_3535,N_49717,N_48630);
and UO_3536 (O_3536,N_48540,N_49622);
xor UO_3537 (O_3537,N_48038,N_48881);
or UO_3538 (O_3538,N_49297,N_49829);
nor UO_3539 (O_3539,N_49259,N_49355);
nand UO_3540 (O_3540,N_49728,N_48750);
or UO_3541 (O_3541,N_48779,N_48387);
and UO_3542 (O_3542,N_49474,N_48871);
nor UO_3543 (O_3543,N_48322,N_49935);
nor UO_3544 (O_3544,N_48239,N_48572);
and UO_3545 (O_3545,N_48253,N_48899);
xnor UO_3546 (O_3546,N_48751,N_49656);
or UO_3547 (O_3547,N_49562,N_48818);
and UO_3548 (O_3548,N_48483,N_49255);
or UO_3549 (O_3549,N_49345,N_49377);
nor UO_3550 (O_3550,N_49663,N_49232);
xnor UO_3551 (O_3551,N_48119,N_49870);
xnor UO_3552 (O_3552,N_49670,N_49096);
and UO_3553 (O_3553,N_48533,N_49979);
xor UO_3554 (O_3554,N_49702,N_49571);
nor UO_3555 (O_3555,N_49850,N_48251);
xnor UO_3556 (O_3556,N_48977,N_48237);
nand UO_3557 (O_3557,N_48104,N_48992);
nand UO_3558 (O_3558,N_48303,N_49201);
nor UO_3559 (O_3559,N_49461,N_48222);
and UO_3560 (O_3560,N_49264,N_49559);
or UO_3561 (O_3561,N_48180,N_49055);
nand UO_3562 (O_3562,N_49001,N_49614);
and UO_3563 (O_3563,N_48465,N_49755);
and UO_3564 (O_3564,N_48150,N_48636);
and UO_3565 (O_3565,N_49397,N_48391);
and UO_3566 (O_3566,N_48736,N_48494);
xor UO_3567 (O_3567,N_49721,N_48971);
nor UO_3568 (O_3568,N_48271,N_49169);
and UO_3569 (O_3569,N_49143,N_49276);
or UO_3570 (O_3570,N_48080,N_48396);
nor UO_3571 (O_3571,N_49897,N_49064);
xor UO_3572 (O_3572,N_48651,N_48104);
nand UO_3573 (O_3573,N_49394,N_49656);
or UO_3574 (O_3574,N_49222,N_48415);
nand UO_3575 (O_3575,N_49673,N_48901);
or UO_3576 (O_3576,N_49389,N_49858);
or UO_3577 (O_3577,N_48210,N_49617);
xor UO_3578 (O_3578,N_48677,N_49975);
xnor UO_3579 (O_3579,N_49779,N_48068);
nand UO_3580 (O_3580,N_48005,N_49508);
and UO_3581 (O_3581,N_49678,N_49592);
and UO_3582 (O_3582,N_48561,N_48001);
xor UO_3583 (O_3583,N_48516,N_49148);
or UO_3584 (O_3584,N_49083,N_48927);
or UO_3585 (O_3585,N_49624,N_48753);
nor UO_3586 (O_3586,N_48485,N_49608);
nor UO_3587 (O_3587,N_49651,N_49138);
nor UO_3588 (O_3588,N_48567,N_49974);
nand UO_3589 (O_3589,N_49610,N_49476);
and UO_3590 (O_3590,N_48931,N_49507);
xor UO_3591 (O_3591,N_48800,N_48534);
and UO_3592 (O_3592,N_48056,N_48977);
xor UO_3593 (O_3593,N_48601,N_48390);
and UO_3594 (O_3594,N_49313,N_49588);
nor UO_3595 (O_3595,N_49055,N_48493);
xnor UO_3596 (O_3596,N_48321,N_48058);
nand UO_3597 (O_3597,N_49713,N_49237);
and UO_3598 (O_3598,N_48727,N_48064);
or UO_3599 (O_3599,N_48666,N_49378);
nor UO_3600 (O_3600,N_48951,N_49820);
xnor UO_3601 (O_3601,N_49878,N_49714);
nor UO_3602 (O_3602,N_49178,N_48206);
nand UO_3603 (O_3603,N_49756,N_48932);
and UO_3604 (O_3604,N_48803,N_48911);
nand UO_3605 (O_3605,N_49393,N_48895);
and UO_3606 (O_3606,N_48379,N_49054);
xnor UO_3607 (O_3607,N_48539,N_48503);
and UO_3608 (O_3608,N_49418,N_48374);
xnor UO_3609 (O_3609,N_48356,N_49264);
and UO_3610 (O_3610,N_48672,N_48069);
and UO_3611 (O_3611,N_48109,N_49694);
or UO_3612 (O_3612,N_49055,N_49016);
xnor UO_3613 (O_3613,N_49235,N_49226);
nor UO_3614 (O_3614,N_49768,N_48597);
nor UO_3615 (O_3615,N_48097,N_49513);
xor UO_3616 (O_3616,N_49833,N_49065);
and UO_3617 (O_3617,N_48496,N_49089);
nor UO_3618 (O_3618,N_49355,N_48058);
nand UO_3619 (O_3619,N_48826,N_48174);
or UO_3620 (O_3620,N_48159,N_48840);
xnor UO_3621 (O_3621,N_48393,N_49285);
or UO_3622 (O_3622,N_48457,N_49657);
nor UO_3623 (O_3623,N_48035,N_48521);
or UO_3624 (O_3624,N_49251,N_49706);
nor UO_3625 (O_3625,N_48191,N_49570);
xnor UO_3626 (O_3626,N_49923,N_49748);
nand UO_3627 (O_3627,N_49492,N_48589);
xor UO_3628 (O_3628,N_48190,N_48837);
nor UO_3629 (O_3629,N_49831,N_48356);
and UO_3630 (O_3630,N_48484,N_48437);
xnor UO_3631 (O_3631,N_48670,N_49478);
nand UO_3632 (O_3632,N_48093,N_48839);
or UO_3633 (O_3633,N_49674,N_48711);
and UO_3634 (O_3634,N_49306,N_48520);
and UO_3635 (O_3635,N_48489,N_48009);
and UO_3636 (O_3636,N_48815,N_48511);
and UO_3637 (O_3637,N_49665,N_48495);
or UO_3638 (O_3638,N_49589,N_49460);
nand UO_3639 (O_3639,N_48383,N_48201);
xnor UO_3640 (O_3640,N_49372,N_48728);
or UO_3641 (O_3641,N_48345,N_48747);
xnor UO_3642 (O_3642,N_49657,N_49923);
nand UO_3643 (O_3643,N_49969,N_48169);
and UO_3644 (O_3644,N_48463,N_48977);
or UO_3645 (O_3645,N_48897,N_48592);
or UO_3646 (O_3646,N_48168,N_49891);
nor UO_3647 (O_3647,N_49945,N_49555);
or UO_3648 (O_3648,N_48285,N_48975);
xnor UO_3649 (O_3649,N_48255,N_48879);
nor UO_3650 (O_3650,N_48937,N_49001);
nor UO_3651 (O_3651,N_49600,N_48088);
nand UO_3652 (O_3652,N_48806,N_49153);
nand UO_3653 (O_3653,N_48050,N_49889);
xor UO_3654 (O_3654,N_48031,N_48827);
xnor UO_3655 (O_3655,N_49873,N_48310);
and UO_3656 (O_3656,N_48246,N_49751);
or UO_3657 (O_3657,N_49421,N_48507);
and UO_3658 (O_3658,N_49382,N_49972);
and UO_3659 (O_3659,N_48153,N_49459);
xor UO_3660 (O_3660,N_48813,N_49754);
and UO_3661 (O_3661,N_48890,N_49162);
nor UO_3662 (O_3662,N_48944,N_48057);
nor UO_3663 (O_3663,N_48798,N_49025);
nor UO_3664 (O_3664,N_48418,N_48728);
nor UO_3665 (O_3665,N_49959,N_48542);
nor UO_3666 (O_3666,N_48022,N_49219);
nand UO_3667 (O_3667,N_48767,N_49045);
nand UO_3668 (O_3668,N_49211,N_48571);
nor UO_3669 (O_3669,N_49515,N_49219);
nor UO_3670 (O_3670,N_49559,N_49025);
xor UO_3671 (O_3671,N_49178,N_49669);
nor UO_3672 (O_3672,N_49998,N_48580);
xor UO_3673 (O_3673,N_49549,N_48325);
xor UO_3674 (O_3674,N_48856,N_49314);
nor UO_3675 (O_3675,N_48837,N_48135);
and UO_3676 (O_3676,N_48161,N_49594);
or UO_3677 (O_3677,N_48007,N_48357);
xor UO_3678 (O_3678,N_48510,N_49585);
nand UO_3679 (O_3679,N_49500,N_48412);
xnor UO_3680 (O_3680,N_48353,N_49849);
or UO_3681 (O_3681,N_49579,N_48633);
nor UO_3682 (O_3682,N_48970,N_48204);
nor UO_3683 (O_3683,N_48930,N_48572);
nand UO_3684 (O_3684,N_49841,N_48235);
nand UO_3685 (O_3685,N_49366,N_48044);
and UO_3686 (O_3686,N_49345,N_48427);
nor UO_3687 (O_3687,N_49381,N_48008);
and UO_3688 (O_3688,N_48926,N_48167);
or UO_3689 (O_3689,N_48593,N_49469);
or UO_3690 (O_3690,N_49094,N_48884);
xor UO_3691 (O_3691,N_48220,N_48612);
or UO_3692 (O_3692,N_49390,N_49750);
xnor UO_3693 (O_3693,N_48773,N_48356);
or UO_3694 (O_3694,N_49422,N_49465);
nor UO_3695 (O_3695,N_48113,N_48319);
nor UO_3696 (O_3696,N_48309,N_48927);
and UO_3697 (O_3697,N_49350,N_49220);
nor UO_3698 (O_3698,N_49370,N_49254);
nand UO_3699 (O_3699,N_49887,N_48332);
xnor UO_3700 (O_3700,N_48933,N_49018);
xnor UO_3701 (O_3701,N_48569,N_48073);
xor UO_3702 (O_3702,N_49735,N_48172);
xor UO_3703 (O_3703,N_48370,N_49619);
nor UO_3704 (O_3704,N_49662,N_49398);
xnor UO_3705 (O_3705,N_49978,N_49531);
nand UO_3706 (O_3706,N_48523,N_48890);
xor UO_3707 (O_3707,N_48806,N_48459);
nand UO_3708 (O_3708,N_48937,N_49196);
nor UO_3709 (O_3709,N_49215,N_48111);
nor UO_3710 (O_3710,N_48658,N_48416);
nand UO_3711 (O_3711,N_49635,N_48651);
nand UO_3712 (O_3712,N_48995,N_49459);
nor UO_3713 (O_3713,N_48729,N_49958);
or UO_3714 (O_3714,N_49576,N_48522);
nor UO_3715 (O_3715,N_48973,N_49806);
or UO_3716 (O_3716,N_48302,N_49708);
or UO_3717 (O_3717,N_49739,N_49969);
nor UO_3718 (O_3718,N_48144,N_48551);
and UO_3719 (O_3719,N_49724,N_49740);
and UO_3720 (O_3720,N_48324,N_49704);
and UO_3721 (O_3721,N_48728,N_49208);
and UO_3722 (O_3722,N_48226,N_49014);
xnor UO_3723 (O_3723,N_48178,N_49483);
and UO_3724 (O_3724,N_49338,N_48119);
or UO_3725 (O_3725,N_48000,N_48562);
nand UO_3726 (O_3726,N_48351,N_49656);
nor UO_3727 (O_3727,N_48522,N_49146);
or UO_3728 (O_3728,N_49812,N_49132);
and UO_3729 (O_3729,N_48190,N_48196);
nor UO_3730 (O_3730,N_48383,N_48556);
xor UO_3731 (O_3731,N_49119,N_48192);
nor UO_3732 (O_3732,N_48267,N_49230);
or UO_3733 (O_3733,N_48819,N_49875);
or UO_3734 (O_3734,N_49379,N_48916);
xor UO_3735 (O_3735,N_48014,N_49551);
nor UO_3736 (O_3736,N_48927,N_49435);
xor UO_3737 (O_3737,N_49943,N_49050);
or UO_3738 (O_3738,N_48135,N_48161);
nor UO_3739 (O_3739,N_49799,N_48591);
and UO_3740 (O_3740,N_48664,N_48985);
nor UO_3741 (O_3741,N_48838,N_49380);
xor UO_3742 (O_3742,N_48847,N_48184);
xnor UO_3743 (O_3743,N_48013,N_48171);
xnor UO_3744 (O_3744,N_49577,N_48191);
nor UO_3745 (O_3745,N_48813,N_48447);
nor UO_3746 (O_3746,N_49281,N_48885);
and UO_3747 (O_3747,N_49124,N_48991);
nand UO_3748 (O_3748,N_49366,N_49147);
nor UO_3749 (O_3749,N_48857,N_48766);
and UO_3750 (O_3750,N_49270,N_48691);
nor UO_3751 (O_3751,N_48080,N_49538);
or UO_3752 (O_3752,N_49996,N_48578);
or UO_3753 (O_3753,N_48119,N_49179);
and UO_3754 (O_3754,N_48947,N_48052);
nor UO_3755 (O_3755,N_48041,N_49593);
nand UO_3756 (O_3756,N_49954,N_49565);
nand UO_3757 (O_3757,N_48481,N_49753);
nand UO_3758 (O_3758,N_48823,N_49384);
xor UO_3759 (O_3759,N_48319,N_49862);
nand UO_3760 (O_3760,N_49911,N_48374);
nand UO_3761 (O_3761,N_48333,N_48737);
xnor UO_3762 (O_3762,N_49227,N_49682);
nor UO_3763 (O_3763,N_49243,N_48548);
xnor UO_3764 (O_3764,N_49646,N_49443);
and UO_3765 (O_3765,N_48941,N_48536);
or UO_3766 (O_3766,N_48067,N_48174);
xnor UO_3767 (O_3767,N_49844,N_49103);
nor UO_3768 (O_3768,N_49771,N_49727);
xor UO_3769 (O_3769,N_48422,N_49461);
nor UO_3770 (O_3770,N_49052,N_49853);
and UO_3771 (O_3771,N_48802,N_49886);
nand UO_3772 (O_3772,N_48971,N_49003);
nand UO_3773 (O_3773,N_48972,N_48774);
xnor UO_3774 (O_3774,N_48931,N_49423);
nor UO_3775 (O_3775,N_48075,N_48981);
nor UO_3776 (O_3776,N_48897,N_49284);
and UO_3777 (O_3777,N_49748,N_49720);
nand UO_3778 (O_3778,N_48027,N_48323);
xor UO_3779 (O_3779,N_48440,N_49422);
and UO_3780 (O_3780,N_49462,N_48948);
nand UO_3781 (O_3781,N_48864,N_48201);
nand UO_3782 (O_3782,N_49644,N_48444);
xnor UO_3783 (O_3783,N_49471,N_49542);
nor UO_3784 (O_3784,N_49245,N_48621);
and UO_3785 (O_3785,N_49443,N_49344);
and UO_3786 (O_3786,N_49141,N_49236);
or UO_3787 (O_3787,N_48430,N_49209);
nand UO_3788 (O_3788,N_49217,N_48913);
xor UO_3789 (O_3789,N_49647,N_48411);
xnor UO_3790 (O_3790,N_49094,N_49610);
and UO_3791 (O_3791,N_49654,N_48444);
and UO_3792 (O_3792,N_49974,N_49752);
and UO_3793 (O_3793,N_48046,N_48980);
or UO_3794 (O_3794,N_49242,N_48514);
nor UO_3795 (O_3795,N_49736,N_49328);
and UO_3796 (O_3796,N_49909,N_48050);
or UO_3797 (O_3797,N_49423,N_49406);
or UO_3798 (O_3798,N_48797,N_48006);
or UO_3799 (O_3799,N_49297,N_49314);
nor UO_3800 (O_3800,N_48302,N_48432);
nand UO_3801 (O_3801,N_48599,N_49161);
nor UO_3802 (O_3802,N_48118,N_48534);
nand UO_3803 (O_3803,N_49092,N_48967);
xor UO_3804 (O_3804,N_49614,N_49533);
or UO_3805 (O_3805,N_49674,N_49802);
or UO_3806 (O_3806,N_48899,N_49578);
nand UO_3807 (O_3807,N_49530,N_49105);
or UO_3808 (O_3808,N_49347,N_49674);
nor UO_3809 (O_3809,N_48430,N_48802);
xnor UO_3810 (O_3810,N_49757,N_48174);
nand UO_3811 (O_3811,N_49332,N_49157);
nand UO_3812 (O_3812,N_49998,N_49343);
xnor UO_3813 (O_3813,N_48813,N_48805);
nand UO_3814 (O_3814,N_49973,N_48483);
nand UO_3815 (O_3815,N_48128,N_48495);
and UO_3816 (O_3816,N_48923,N_49642);
nand UO_3817 (O_3817,N_49408,N_49689);
nor UO_3818 (O_3818,N_49164,N_49920);
xnor UO_3819 (O_3819,N_48733,N_48156);
nand UO_3820 (O_3820,N_48751,N_48181);
or UO_3821 (O_3821,N_48398,N_49593);
nor UO_3822 (O_3822,N_49143,N_48051);
and UO_3823 (O_3823,N_49275,N_49549);
xor UO_3824 (O_3824,N_49097,N_49436);
nor UO_3825 (O_3825,N_49018,N_48065);
or UO_3826 (O_3826,N_48925,N_48874);
nor UO_3827 (O_3827,N_49127,N_49515);
nor UO_3828 (O_3828,N_49095,N_49472);
or UO_3829 (O_3829,N_49996,N_48463);
and UO_3830 (O_3830,N_49661,N_48591);
and UO_3831 (O_3831,N_49190,N_48949);
nor UO_3832 (O_3832,N_48635,N_49885);
and UO_3833 (O_3833,N_49776,N_49611);
nand UO_3834 (O_3834,N_48721,N_49370);
nand UO_3835 (O_3835,N_49264,N_48334);
xor UO_3836 (O_3836,N_48510,N_48431);
or UO_3837 (O_3837,N_49382,N_48131);
and UO_3838 (O_3838,N_48019,N_49483);
xnor UO_3839 (O_3839,N_48649,N_48902);
nand UO_3840 (O_3840,N_48132,N_48059);
nand UO_3841 (O_3841,N_49054,N_48700);
xnor UO_3842 (O_3842,N_49534,N_49641);
nor UO_3843 (O_3843,N_48920,N_48429);
and UO_3844 (O_3844,N_49862,N_48606);
nor UO_3845 (O_3845,N_49993,N_48393);
and UO_3846 (O_3846,N_49616,N_48835);
or UO_3847 (O_3847,N_49684,N_48553);
xnor UO_3848 (O_3848,N_49898,N_49821);
and UO_3849 (O_3849,N_49303,N_48339);
nor UO_3850 (O_3850,N_48415,N_48801);
or UO_3851 (O_3851,N_49274,N_48659);
and UO_3852 (O_3852,N_48052,N_48624);
and UO_3853 (O_3853,N_48909,N_49365);
nand UO_3854 (O_3854,N_48365,N_49946);
nor UO_3855 (O_3855,N_48748,N_48659);
or UO_3856 (O_3856,N_49568,N_48167);
nor UO_3857 (O_3857,N_48005,N_49872);
and UO_3858 (O_3858,N_48793,N_48135);
nand UO_3859 (O_3859,N_48082,N_49630);
or UO_3860 (O_3860,N_49862,N_49445);
xor UO_3861 (O_3861,N_48829,N_49071);
and UO_3862 (O_3862,N_49327,N_49926);
and UO_3863 (O_3863,N_48789,N_49163);
nand UO_3864 (O_3864,N_48006,N_49890);
nand UO_3865 (O_3865,N_49795,N_49740);
and UO_3866 (O_3866,N_49603,N_49269);
xnor UO_3867 (O_3867,N_49671,N_49011);
or UO_3868 (O_3868,N_49737,N_48222);
or UO_3869 (O_3869,N_48458,N_49004);
nand UO_3870 (O_3870,N_48584,N_49287);
nor UO_3871 (O_3871,N_49802,N_49512);
xor UO_3872 (O_3872,N_49905,N_49951);
and UO_3873 (O_3873,N_49330,N_48028);
nor UO_3874 (O_3874,N_49048,N_49719);
xnor UO_3875 (O_3875,N_49783,N_49902);
or UO_3876 (O_3876,N_48893,N_49389);
nand UO_3877 (O_3877,N_48456,N_48867);
and UO_3878 (O_3878,N_49115,N_48944);
and UO_3879 (O_3879,N_48328,N_48170);
nor UO_3880 (O_3880,N_49167,N_49565);
xor UO_3881 (O_3881,N_48656,N_48582);
xnor UO_3882 (O_3882,N_48904,N_49472);
or UO_3883 (O_3883,N_48775,N_48058);
nand UO_3884 (O_3884,N_48951,N_48997);
nor UO_3885 (O_3885,N_48532,N_49300);
nor UO_3886 (O_3886,N_49793,N_48899);
or UO_3887 (O_3887,N_49268,N_48238);
nand UO_3888 (O_3888,N_48308,N_49853);
nor UO_3889 (O_3889,N_48969,N_49008);
nor UO_3890 (O_3890,N_49213,N_49770);
or UO_3891 (O_3891,N_49266,N_49351);
or UO_3892 (O_3892,N_49054,N_49638);
nand UO_3893 (O_3893,N_48634,N_49746);
and UO_3894 (O_3894,N_49900,N_49296);
nand UO_3895 (O_3895,N_48963,N_48900);
or UO_3896 (O_3896,N_48944,N_48265);
and UO_3897 (O_3897,N_48457,N_48338);
and UO_3898 (O_3898,N_49822,N_48766);
and UO_3899 (O_3899,N_49538,N_49308);
nand UO_3900 (O_3900,N_48361,N_48831);
or UO_3901 (O_3901,N_49498,N_48913);
or UO_3902 (O_3902,N_48229,N_49635);
or UO_3903 (O_3903,N_48845,N_49422);
nor UO_3904 (O_3904,N_49872,N_48675);
xor UO_3905 (O_3905,N_49214,N_48596);
and UO_3906 (O_3906,N_49206,N_48183);
or UO_3907 (O_3907,N_48553,N_49152);
or UO_3908 (O_3908,N_49089,N_48003);
nand UO_3909 (O_3909,N_49057,N_48585);
xnor UO_3910 (O_3910,N_48391,N_49788);
nand UO_3911 (O_3911,N_49189,N_48541);
nand UO_3912 (O_3912,N_49685,N_49686);
or UO_3913 (O_3913,N_48428,N_49906);
nor UO_3914 (O_3914,N_48376,N_49497);
xor UO_3915 (O_3915,N_49059,N_49021);
and UO_3916 (O_3916,N_48170,N_49153);
or UO_3917 (O_3917,N_49219,N_48439);
or UO_3918 (O_3918,N_49750,N_49503);
xnor UO_3919 (O_3919,N_49929,N_48610);
nor UO_3920 (O_3920,N_49713,N_49626);
or UO_3921 (O_3921,N_48903,N_48357);
nand UO_3922 (O_3922,N_48297,N_49352);
nor UO_3923 (O_3923,N_49795,N_48622);
and UO_3924 (O_3924,N_48532,N_48254);
nand UO_3925 (O_3925,N_49982,N_49476);
and UO_3926 (O_3926,N_49458,N_49683);
and UO_3927 (O_3927,N_49794,N_48398);
and UO_3928 (O_3928,N_49668,N_49142);
and UO_3929 (O_3929,N_49877,N_48524);
and UO_3930 (O_3930,N_48878,N_49733);
or UO_3931 (O_3931,N_49101,N_49231);
or UO_3932 (O_3932,N_49084,N_48779);
or UO_3933 (O_3933,N_48800,N_48706);
or UO_3934 (O_3934,N_48716,N_49664);
nand UO_3935 (O_3935,N_49065,N_48525);
nor UO_3936 (O_3936,N_49510,N_49286);
xnor UO_3937 (O_3937,N_49782,N_49768);
and UO_3938 (O_3938,N_48563,N_48237);
and UO_3939 (O_3939,N_48776,N_49332);
and UO_3940 (O_3940,N_49501,N_49105);
and UO_3941 (O_3941,N_48953,N_49773);
or UO_3942 (O_3942,N_48812,N_49340);
and UO_3943 (O_3943,N_48895,N_49212);
xor UO_3944 (O_3944,N_49779,N_48654);
or UO_3945 (O_3945,N_49715,N_49587);
and UO_3946 (O_3946,N_48684,N_48180);
nor UO_3947 (O_3947,N_48361,N_48994);
xnor UO_3948 (O_3948,N_48391,N_49325);
xor UO_3949 (O_3949,N_48263,N_48391);
or UO_3950 (O_3950,N_49171,N_49929);
nand UO_3951 (O_3951,N_48910,N_48084);
xnor UO_3952 (O_3952,N_49528,N_48334);
nor UO_3953 (O_3953,N_48889,N_48544);
nor UO_3954 (O_3954,N_49224,N_48720);
and UO_3955 (O_3955,N_48481,N_49338);
or UO_3956 (O_3956,N_48716,N_48324);
and UO_3957 (O_3957,N_49048,N_48897);
nor UO_3958 (O_3958,N_48336,N_48089);
and UO_3959 (O_3959,N_48029,N_49507);
xnor UO_3960 (O_3960,N_48145,N_49763);
and UO_3961 (O_3961,N_49368,N_48445);
and UO_3962 (O_3962,N_48277,N_48766);
nor UO_3963 (O_3963,N_48582,N_48015);
nand UO_3964 (O_3964,N_48964,N_49603);
and UO_3965 (O_3965,N_48553,N_48023);
and UO_3966 (O_3966,N_48461,N_49472);
nand UO_3967 (O_3967,N_49262,N_49360);
or UO_3968 (O_3968,N_49577,N_49673);
xnor UO_3969 (O_3969,N_49688,N_49933);
and UO_3970 (O_3970,N_49775,N_48449);
or UO_3971 (O_3971,N_49819,N_49335);
xnor UO_3972 (O_3972,N_48562,N_48244);
and UO_3973 (O_3973,N_48052,N_49959);
nand UO_3974 (O_3974,N_48893,N_48556);
nand UO_3975 (O_3975,N_49937,N_49784);
or UO_3976 (O_3976,N_49706,N_49747);
and UO_3977 (O_3977,N_48649,N_49691);
nand UO_3978 (O_3978,N_49666,N_49159);
nor UO_3979 (O_3979,N_49860,N_48238);
xor UO_3980 (O_3980,N_49659,N_49153);
xnor UO_3981 (O_3981,N_48433,N_48055);
and UO_3982 (O_3982,N_49653,N_48236);
nand UO_3983 (O_3983,N_48108,N_49129);
nand UO_3984 (O_3984,N_48666,N_49908);
or UO_3985 (O_3985,N_48584,N_48018);
and UO_3986 (O_3986,N_48258,N_49370);
xor UO_3987 (O_3987,N_48898,N_48882);
or UO_3988 (O_3988,N_48137,N_49160);
xor UO_3989 (O_3989,N_49413,N_49255);
nand UO_3990 (O_3990,N_49028,N_48682);
nand UO_3991 (O_3991,N_49155,N_49800);
nor UO_3992 (O_3992,N_49354,N_48444);
xor UO_3993 (O_3993,N_48866,N_49161);
or UO_3994 (O_3994,N_48182,N_48942);
nor UO_3995 (O_3995,N_49848,N_48316);
xor UO_3996 (O_3996,N_48506,N_49907);
and UO_3997 (O_3997,N_48174,N_48575);
nor UO_3998 (O_3998,N_49615,N_48866);
and UO_3999 (O_3999,N_49391,N_48264);
xnor UO_4000 (O_4000,N_49165,N_49341);
and UO_4001 (O_4001,N_49178,N_48817);
xor UO_4002 (O_4002,N_48076,N_48281);
nor UO_4003 (O_4003,N_48597,N_49066);
or UO_4004 (O_4004,N_48469,N_49831);
xnor UO_4005 (O_4005,N_49341,N_49209);
xnor UO_4006 (O_4006,N_48665,N_49160);
or UO_4007 (O_4007,N_48317,N_49153);
xor UO_4008 (O_4008,N_48979,N_48677);
nor UO_4009 (O_4009,N_48502,N_49416);
or UO_4010 (O_4010,N_49878,N_49787);
xnor UO_4011 (O_4011,N_49294,N_49538);
nand UO_4012 (O_4012,N_49856,N_49686);
and UO_4013 (O_4013,N_49466,N_49168);
xor UO_4014 (O_4014,N_49230,N_49645);
xor UO_4015 (O_4015,N_49090,N_48180);
nor UO_4016 (O_4016,N_48649,N_48630);
or UO_4017 (O_4017,N_48774,N_49918);
nor UO_4018 (O_4018,N_48097,N_49009);
nor UO_4019 (O_4019,N_48626,N_49311);
nand UO_4020 (O_4020,N_48285,N_49110);
or UO_4021 (O_4021,N_48422,N_48377);
xor UO_4022 (O_4022,N_49865,N_48622);
or UO_4023 (O_4023,N_49433,N_49060);
or UO_4024 (O_4024,N_49410,N_48032);
and UO_4025 (O_4025,N_48731,N_48186);
nand UO_4026 (O_4026,N_48995,N_49552);
and UO_4027 (O_4027,N_49023,N_48792);
or UO_4028 (O_4028,N_48598,N_49761);
or UO_4029 (O_4029,N_48996,N_48780);
nand UO_4030 (O_4030,N_49483,N_48205);
or UO_4031 (O_4031,N_48165,N_48274);
xnor UO_4032 (O_4032,N_48951,N_49719);
or UO_4033 (O_4033,N_49292,N_48805);
xor UO_4034 (O_4034,N_49875,N_48096);
or UO_4035 (O_4035,N_49433,N_49424);
xnor UO_4036 (O_4036,N_48665,N_49756);
nand UO_4037 (O_4037,N_49500,N_49089);
nor UO_4038 (O_4038,N_48403,N_49795);
nand UO_4039 (O_4039,N_48308,N_49399);
nor UO_4040 (O_4040,N_48141,N_49785);
xnor UO_4041 (O_4041,N_48863,N_48174);
nor UO_4042 (O_4042,N_49660,N_49204);
xnor UO_4043 (O_4043,N_48758,N_48816);
or UO_4044 (O_4044,N_48093,N_48250);
or UO_4045 (O_4045,N_49043,N_49814);
or UO_4046 (O_4046,N_49185,N_49383);
or UO_4047 (O_4047,N_49202,N_49106);
and UO_4048 (O_4048,N_48500,N_49431);
xor UO_4049 (O_4049,N_49002,N_48174);
xnor UO_4050 (O_4050,N_49834,N_49729);
nor UO_4051 (O_4051,N_49238,N_48184);
nand UO_4052 (O_4052,N_48120,N_48498);
or UO_4053 (O_4053,N_49960,N_48093);
xor UO_4054 (O_4054,N_48387,N_49007);
and UO_4055 (O_4055,N_49229,N_49041);
or UO_4056 (O_4056,N_49083,N_48367);
xnor UO_4057 (O_4057,N_49835,N_48492);
xor UO_4058 (O_4058,N_49894,N_49587);
and UO_4059 (O_4059,N_48142,N_49360);
and UO_4060 (O_4060,N_48925,N_48037);
nand UO_4061 (O_4061,N_49066,N_49084);
and UO_4062 (O_4062,N_49069,N_49601);
or UO_4063 (O_4063,N_48496,N_48360);
xor UO_4064 (O_4064,N_49215,N_48172);
or UO_4065 (O_4065,N_49299,N_49984);
nand UO_4066 (O_4066,N_48311,N_49547);
and UO_4067 (O_4067,N_49354,N_49101);
and UO_4068 (O_4068,N_49430,N_48654);
nor UO_4069 (O_4069,N_49014,N_48079);
nor UO_4070 (O_4070,N_49113,N_49932);
nor UO_4071 (O_4071,N_48807,N_48925);
or UO_4072 (O_4072,N_49162,N_49863);
xnor UO_4073 (O_4073,N_49948,N_49263);
or UO_4074 (O_4074,N_48213,N_49417);
xor UO_4075 (O_4075,N_49604,N_48937);
or UO_4076 (O_4076,N_48260,N_49137);
nor UO_4077 (O_4077,N_49333,N_49982);
nand UO_4078 (O_4078,N_48864,N_48915);
and UO_4079 (O_4079,N_48310,N_49040);
or UO_4080 (O_4080,N_48209,N_49898);
nor UO_4081 (O_4081,N_49273,N_48137);
or UO_4082 (O_4082,N_49996,N_48580);
nand UO_4083 (O_4083,N_48081,N_49047);
and UO_4084 (O_4084,N_49770,N_48096);
and UO_4085 (O_4085,N_48645,N_49649);
or UO_4086 (O_4086,N_48932,N_49603);
nor UO_4087 (O_4087,N_48173,N_48213);
nand UO_4088 (O_4088,N_49091,N_49752);
and UO_4089 (O_4089,N_48990,N_49276);
nor UO_4090 (O_4090,N_49625,N_48501);
nor UO_4091 (O_4091,N_48604,N_48654);
or UO_4092 (O_4092,N_48383,N_49611);
and UO_4093 (O_4093,N_48781,N_48675);
and UO_4094 (O_4094,N_48739,N_48825);
nor UO_4095 (O_4095,N_48940,N_48446);
nor UO_4096 (O_4096,N_49253,N_48222);
nand UO_4097 (O_4097,N_48657,N_49410);
and UO_4098 (O_4098,N_48316,N_49112);
nand UO_4099 (O_4099,N_49807,N_49234);
nand UO_4100 (O_4100,N_49210,N_49055);
or UO_4101 (O_4101,N_48754,N_48985);
and UO_4102 (O_4102,N_48737,N_49888);
or UO_4103 (O_4103,N_48209,N_48599);
or UO_4104 (O_4104,N_49236,N_48078);
or UO_4105 (O_4105,N_49401,N_48714);
and UO_4106 (O_4106,N_49653,N_48033);
nor UO_4107 (O_4107,N_49995,N_48421);
xnor UO_4108 (O_4108,N_49872,N_48133);
nor UO_4109 (O_4109,N_48648,N_48280);
xnor UO_4110 (O_4110,N_49631,N_49280);
and UO_4111 (O_4111,N_48991,N_48024);
or UO_4112 (O_4112,N_48207,N_48465);
nor UO_4113 (O_4113,N_48065,N_49585);
and UO_4114 (O_4114,N_49329,N_49586);
nand UO_4115 (O_4115,N_49384,N_48780);
and UO_4116 (O_4116,N_49741,N_48554);
nor UO_4117 (O_4117,N_48870,N_49593);
nand UO_4118 (O_4118,N_49231,N_48830);
nand UO_4119 (O_4119,N_48717,N_49096);
nand UO_4120 (O_4120,N_48271,N_49941);
nand UO_4121 (O_4121,N_49920,N_49720);
nor UO_4122 (O_4122,N_48322,N_48421);
and UO_4123 (O_4123,N_49196,N_48238);
and UO_4124 (O_4124,N_49957,N_49074);
nor UO_4125 (O_4125,N_49350,N_48926);
and UO_4126 (O_4126,N_49796,N_49695);
or UO_4127 (O_4127,N_49875,N_48971);
nor UO_4128 (O_4128,N_49644,N_48891);
nand UO_4129 (O_4129,N_48167,N_48334);
nand UO_4130 (O_4130,N_49965,N_48953);
nand UO_4131 (O_4131,N_48964,N_48039);
nand UO_4132 (O_4132,N_49659,N_48590);
xor UO_4133 (O_4133,N_49389,N_48058);
and UO_4134 (O_4134,N_49718,N_49121);
and UO_4135 (O_4135,N_49053,N_49743);
nor UO_4136 (O_4136,N_48256,N_49127);
and UO_4137 (O_4137,N_49395,N_49043);
nor UO_4138 (O_4138,N_49410,N_49688);
xnor UO_4139 (O_4139,N_49492,N_48017);
xnor UO_4140 (O_4140,N_49068,N_48182);
xnor UO_4141 (O_4141,N_49483,N_49640);
xnor UO_4142 (O_4142,N_48076,N_49028);
nand UO_4143 (O_4143,N_49625,N_49020);
nor UO_4144 (O_4144,N_48208,N_48776);
nand UO_4145 (O_4145,N_48210,N_49108);
nand UO_4146 (O_4146,N_48858,N_48478);
nand UO_4147 (O_4147,N_48481,N_49783);
nand UO_4148 (O_4148,N_49926,N_48505);
and UO_4149 (O_4149,N_48819,N_48274);
nor UO_4150 (O_4150,N_49152,N_48198);
and UO_4151 (O_4151,N_49972,N_48885);
xor UO_4152 (O_4152,N_48738,N_48252);
xor UO_4153 (O_4153,N_48060,N_48379);
and UO_4154 (O_4154,N_49336,N_49951);
nand UO_4155 (O_4155,N_49697,N_48450);
and UO_4156 (O_4156,N_48478,N_49341);
or UO_4157 (O_4157,N_48979,N_48244);
nand UO_4158 (O_4158,N_48587,N_48631);
or UO_4159 (O_4159,N_48522,N_48839);
nand UO_4160 (O_4160,N_48514,N_48392);
xor UO_4161 (O_4161,N_48393,N_48135);
nand UO_4162 (O_4162,N_48229,N_49133);
and UO_4163 (O_4163,N_48040,N_49865);
nor UO_4164 (O_4164,N_48268,N_48906);
nor UO_4165 (O_4165,N_49345,N_49467);
xnor UO_4166 (O_4166,N_49709,N_48018);
nand UO_4167 (O_4167,N_49971,N_48755);
xnor UO_4168 (O_4168,N_49516,N_49856);
and UO_4169 (O_4169,N_48824,N_48618);
xor UO_4170 (O_4170,N_49882,N_49912);
nand UO_4171 (O_4171,N_49657,N_49615);
nor UO_4172 (O_4172,N_49535,N_48708);
nor UO_4173 (O_4173,N_48159,N_48646);
xor UO_4174 (O_4174,N_48993,N_48670);
nor UO_4175 (O_4175,N_48247,N_49472);
or UO_4176 (O_4176,N_48499,N_49105);
nor UO_4177 (O_4177,N_49606,N_48086);
nor UO_4178 (O_4178,N_49760,N_48869);
or UO_4179 (O_4179,N_49648,N_48315);
or UO_4180 (O_4180,N_49171,N_49631);
nand UO_4181 (O_4181,N_49273,N_48691);
nor UO_4182 (O_4182,N_48382,N_48389);
and UO_4183 (O_4183,N_48066,N_48254);
and UO_4184 (O_4184,N_48878,N_49442);
nor UO_4185 (O_4185,N_49774,N_48436);
nor UO_4186 (O_4186,N_48726,N_49821);
nor UO_4187 (O_4187,N_48531,N_49990);
nor UO_4188 (O_4188,N_48861,N_49604);
nand UO_4189 (O_4189,N_49517,N_48306);
and UO_4190 (O_4190,N_49616,N_49872);
nor UO_4191 (O_4191,N_48014,N_49336);
nand UO_4192 (O_4192,N_48941,N_48580);
nor UO_4193 (O_4193,N_48244,N_48421);
nand UO_4194 (O_4194,N_48156,N_49298);
or UO_4195 (O_4195,N_49889,N_49666);
or UO_4196 (O_4196,N_49397,N_48237);
or UO_4197 (O_4197,N_48923,N_49953);
and UO_4198 (O_4198,N_48051,N_48410);
nor UO_4199 (O_4199,N_48089,N_48054);
nand UO_4200 (O_4200,N_48524,N_48071);
xor UO_4201 (O_4201,N_48350,N_48408);
xor UO_4202 (O_4202,N_48308,N_48433);
and UO_4203 (O_4203,N_49458,N_48799);
nor UO_4204 (O_4204,N_49723,N_48403);
xnor UO_4205 (O_4205,N_48219,N_49063);
xnor UO_4206 (O_4206,N_48091,N_49402);
nand UO_4207 (O_4207,N_49613,N_48256);
or UO_4208 (O_4208,N_49295,N_49977);
nand UO_4209 (O_4209,N_48736,N_49728);
nand UO_4210 (O_4210,N_49670,N_48063);
xnor UO_4211 (O_4211,N_49291,N_48543);
nor UO_4212 (O_4212,N_48836,N_48537);
and UO_4213 (O_4213,N_48253,N_49881);
xor UO_4214 (O_4214,N_49205,N_49229);
xnor UO_4215 (O_4215,N_49865,N_49567);
xnor UO_4216 (O_4216,N_49715,N_49331);
and UO_4217 (O_4217,N_49030,N_49983);
xor UO_4218 (O_4218,N_49506,N_49627);
nor UO_4219 (O_4219,N_49447,N_48884);
or UO_4220 (O_4220,N_49192,N_48620);
and UO_4221 (O_4221,N_49965,N_49592);
xnor UO_4222 (O_4222,N_48610,N_48204);
and UO_4223 (O_4223,N_48304,N_49313);
nor UO_4224 (O_4224,N_49479,N_48643);
nor UO_4225 (O_4225,N_48692,N_48001);
and UO_4226 (O_4226,N_48733,N_49233);
and UO_4227 (O_4227,N_49548,N_49140);
nor UO_4228 (O_4228,N_48787,N_48715);
nand UO_4229 (O_4229,N_48283,N_49782);
xnor UO_4230 (O_4230,N_48886,N_49398);
or UO_4231 (O_4231,N_49695,N_49073);
nand UO_4232 (O_4232,N_49172,N_49785);
and UO_4233 (O_4233,N_49531,N_49517);
nor UO_4234 (O_4234,N_48117,N_48183);
or UO_4235 (O_4235,N_49534,N_49144);
nor UO_4236 (O_4236,N_49880,N_49437);
and UO_4237 (O_4237,N_48488,N_49086);
nor UO_4238 (O_4238,N_49962,N_49137);
xnor UO_4239 (O_4239,N_49323,N_48928);
nand UO_4240 (O_4240,N_48800,N_49876);
or UO_4241 (O_4241,N_49587,N_48253);
and UO_4242 (O_4242,N_49346,N_49934);
xnor UO_4243 (O_4243,N_48220,N_49622);
and UO_4244 (O_4244,N_49006,N_49410);
nand UO_4245 (O_4245,N_48633,N_49248);
or UO_4246 (O_4246,N_49222,N_49238);
nor UO_4247 (O_4247,N_49983,N_48047);
and UO_4248 (O_4248,N_49081,N_48774);
nand UO_4249 (O_4249,N_48921,N_49581);
or UO_4250 (O_4250,N_49219,N_49419);
nor UO_4251 (O_4251,N_48211,N_48148);
and UO_4252 (O_4252,N_49481,N_49269);
nand UO_4253 (O_4253,N_48452,N_48364);
and UO_4254 (O_4254,N_49103,N_48812);
and UO_4255 (O_4255,N_48122,N_48357);
nor UO_4256 (O_4256,N_49817,N_49360);
xnor UO_4257 (O_4257,N_48935,N_49932);
or UO_4258 (O_4258,N_48142,N_48139);
or UO_4259 (O_4259,N_49804,N_48385);
nor UO_4260 (O_4260,N_48740,N_48728);
or UO_4261 (O_4261,N_49544,N_48792);
nand UO_4262 (O_4262,N_49054,N_48309);
and UO_4263 (O_4263,N_49022,N_49821);
nor UO_4264 (O_4264,N_48211,N_49694);
and UO_4265 (O_4265,N_48648,N_49443);
nor UO_4266 (O_4266,N_48196,N_49119);
nor UO_4267 (O_4267,N_49723,N_48147);
and UO_4268 (O_4268,N_49354,N_49091);
or UO_4269 (O_4269,N_49545,N_48361);
xnor UO_4270 (O_4270,N_48095,N_48881);
and UO_4271 (O_4271,N_48461,N_49990);
nor UO_4272 (O_4272,N_48167,N_49744);
nand UO_4273 (O_4273,N_48256,N_49940);
or UO_4274 (O_4274,N_48302,N_49890);
nand UO_4275 (O_4275,N_49097,N_48724);
xor UO_4276 (O_4276,N_48224,N_48995);
and UO_4277 (O_4277,N_48918,N_49623);
xor UO_4278 (O_4278,N_49883,N_49938);
nand UO_4279 (O_4279,N_48002,N_48368);
and UO_4280 (O_4280,N_48751,N_48846);
nor UO_4281 (O_4281,N_48955,N_49030);
nand UO_4282 (O_4282,N_49516,N_49061);
and UO_4283 (O_4283,N_48767,N_48245);
and UO_4284 (O_4284,N_49209,N_48361);
and UO_4285 (O_4285,N_49388,N_49249);
or UO_4286 (O_4286,N_49089,N_48746);
or UO_4287 (O_4287,N_48425,N_49013);
nand UO_4288 (O_4288,N_49248,N_48382);
xor UO_4289 (O_4289,N_49465,N_49865);
or UO_4290 (O_4290,N_48107,N_49960);
xnor UO_4291 (O_4291,N_49534,N_48289);
nand UO_4292 (O_4292,N_48664,N_49824);
xnor UO_4293 (O_4293,N_48045,N_49572);
xor UO_4294 (O_4294,N_49797,N_49976);
xnor UO_4295 (O_4295,N_49126,N_49965);
xnor UO_4296 (O_4296,N_48100,N_49151);
xor UO_4297 (O_4297,N_48505,N_48057);
xnor UO_4298 (O_4298,N_49042,N_49750);
nand UO_4299 (O_4299,N_49535,N_48422);
nand UO_4300 (O_4300,N_49835,N_48964);
xnor UO_4301 (O_4301,N_49266,N_49133);
nand UO_4302 (O_4302,N_48186,N_49803);
and UO_4303 (O_4303,N_48974,N_48227);
or UO_4304 (O_4304,N_48273,N_49630);
nand UO_4305 (O_4305,N_49668,N_49156);
nand UO_4306 (O_4306,N_49048,N_48438);
xor UO_4307 (O_4307,N_48526,N_49829);
nor UO_4308 (O_4308,N_49224,N_49045);
or UO_4309 (O_4309,N_49269,N_49980);
xor UO_4310 (O_4310,N_49302,N_48994);
and UO_4311 (O_4311,N_49950,N_48999);
and UO_4312 (O_4312,N_49602,N_48633);
nor UO_4313 (O_4313,N_48693,N_48607);
or UO_4314 (O_4314,N_48764,N_48408);
xor UO_4315 (O_4315,N_48730,N_48433);
and UO_4316 (O_4316,N_49695,N_48563);
nor UO_4317 (O_4317,N_48054,N_49780);
and UO_4318 (O_4318,N_49053,N_48918);
xor UO_4319 (O_4319,N_48006,N_48928);
nand UO_4320 (O_4320,N_48952,N_48715);
and UO_4321 (O_4321,N_49299,N_48321);
xor UO_4322 (O_4322,N_48410,N_48052);
nand UO_4323 (O_4323,N_48544,N_49229);
nor UO_4324 (O_4324,N_49957,N_48456);
nand UO_4325 (O_4325,N_49085,N_49818);
and UO_4326 (O_4326,N_48280,N_49117);
and UO_4327 (O_4327,N_48124,N_49162);
nor UO_4328 (O_4328,N_48930,N_49024);
and UO_4329 (O_4329,N_48521,N_48356);
xnor UO_4330 (O_4330,N_48937,N_49792);
or UO_4331 (O_4331,N_49133,N_49908);
or UO_4332 (O_4332,N_48934,N_49407);
or UO_4333 (O_4333,N_48464,N_48069);
xor UO_4334 (O_4334,N_49778,N_49890);
and UO_4335 (O_4335,N_48239,N_48598);
or UO_4336 (O_4336,N_48896,N_49683);
nand UO_4337 (O_4337,N_48526,N_48189);
nand UO_4338 (O_4338,N_48192,N_48796);
or UO_4339 (O_4339,N_49036,N_49195);
nor UO_4340 (O_4340,N_49719,N_48159);
nand UO_4341 (O_4341,N_49157,N_49359);
xor UO_4342 (O_4342,N_48578,N_49858);
xor UO_4343 (O_4343,N_48826,N_48910);
and UO_4344 (O_4344,N_48637,N_49415);
nor UO_4345 (O_4345,N_49012,N_48222);
or UO_4346 (O_4346,N_49568,N_49580);
nand UO_4347 (O_4347,N_49474,N_48455);
nor UO_4348 (O_4348,N_49195,N_48267);
nand UO_4349 (O_4349,N_48900,N_49687);
nor UO_4350 (O_4350,N_48122,N_48205);
nor UO_4351 (O_4351,N_49472,N_48873);
and UO_4352 (O_4352,N_48695,N_49257);
xor UO_4353 (O_4353,N_49354,N_49281);
nor UO_4354 (O_4354,N_48141,N_48928);
nor UO_4355 (O_4355,N_49366,N_49512);
or UO_4356 (O_4356,N_48085,N_48075);
nand UO_4357 (O_4357,N_48437,N_48003);
or UO_4358 (O_4358,N_48025,N_48138);
nand UO_4359 (O_4359,N_49833,N_49116);
or UO_4360 (O_4360,N_49249,N_49161);
and UO_4361 (O_4361,N_49361,N_49635);
nor UO_4362 (O_4362,N_49246,N_48589);
nand UO_4363 (O_4363,N_49094,N_48601);
or UO_4364 (O_4364,N_49189,N_49209);
xnor UO_4365 (O_4365,N_49768,N_48133);
xor UO_4366 (O_4366,N_49397,N_49012);
or UO_4367 (O_4367,N_48856,N_49816);
nor UO_4368 (O_4368,N_48644,N_49476);
xnor UO_4369 (O_4369,N_49449,N_48382);
nand UO_4370 (O_4370,N_49620,N_49920);
or UO_4371 (O_4371,N_49944,N_49539);
nor UO_4372 (O_4372,N_49633,N_48591);
nor UO_4373 (O_4373,N_48440,N_48030);
or UO_4374 (O_4374,N_48319,N_48091);
or UO_4375 (O_4375,N_49570,N_48207);
and UO_4376 (O_4376,N_49009,N_49974);
xor UO_4377 (O_4377,N_48216,N_48908);
and UO_4378 (O_4378,N_48302,N_48166);
nor UO_4379 (O_4379,N_49001,N_48794);
or UO_4380 (O_4380,N_49012,N_49839);
xnor UO_4381 (O_4381,N_48185,N_49718);
nor UO_4382 (O_4382,N_48782,N_49359);
and UO_4383 (O_4383,N_49264,N_48749);
or UO_4384 (O_4384,N_49343,N_48193);
or UO_4385 (O_4385,N_48681,N_49186);
or UO_4386 (O_4386,N_48267,N_49371);
nor UO_4387 (O_4387,N_49090,N_48169);
nand UO_4388 (O_4388,N_49253,N_49562);
xor UO_4389 (O_4389,N_48186,N_49304);
nor UO_4390 (O_4390,N_49589,N_49090);
and UO_4391 (O_4391,N_49306,N_49824);
xnor UO_4392 (O_4392,N_48392,N_49778);
nand UO_4393 (O_4393,N_49499,N_48305);
or UO_4394 (O_4394,N_49505,N_49053);
or UO_4395 (O_4395,N_48482,N_48582);
or UO_4396 (O_4396,N_48808,N_48188);
and UO_4397 (O_4397,N_49738,N_48874);
xnor UO_4398 (O_4398,N_48967,N_49233);
xor UO_4399 (O_4399,N_49247,N_49200);
or UO_4400 (O_4400,N_48648,N_49488);
nand UO_4401 (O_4401,N_49998,N_49773);
xor UO_4402 (O_4402,N_48120,N_49234);
and UO_4403 (O_4403,N_48144,N_49981);
or UO_4404 (O_4404,N_48843,N_49462);
or UO_4405 (O_4405,N_48765,N_48701);
or UO_4406 (O_4406,N_48059,N_49768);
or UO_4407 (O_4407,N_48906,N_48826);
nor UO_4408 (O_4408,N_48773,N_48604);
xnor UO_4409 (O_4409,N_49419,N_48363);
nor UO_4410 (O_4410,N_49854,N_49783);
or UO_4411 (O_4411,N_48982,N_49461);
nand UO_4412 (O_4412,N_49736,N_49939);
nor UO_4413 (O_4413,N_49899,N_48876);
nand UO_4414 (O_4414,N_48015,N_48244);
nor UO_4415 (O_4415,N_48239,N_48115);
and UO_4416 (O_4416,N_48089,N_49567);
or UO_4417 (O_4417,N_48450,N_49836);
xnor UO_4418 (O_4418,N_49960,N_49897);
nand UO_4419 (O_4419,N_49345,N_49607);
nand UO_4420 (O_4420,N_48572,N_49035);
and UO_4421 (O_4421,N_48300,N_49589);
and UO_4422 (O_4422,N_48401,N_48771);
and UO_4423 (O_4423,N_48011,N_49011);
xnor UO_4424 (O_4424,N_48776,N_48714);
or UO_4425 (O_4425,N_49855,N_49857);
nor UO_4426 (O_4426,N_49310,N_48160);
nand UO_4427 (O_4427,N_48598,N_48110);
or UO_4428 (O_4428,N_49945,N_48480);
and UO_4429 (O_4429,N_49390,N_49540);
and UO_4430 (O_4430,N_49181,N_48360);
or UO_4431 (O_4431,N_49867,N_48150);
or UO_4432 (O_4432,N_48323,N_48091);
nand UO_4433 (O_4433,N_48627,N_49784);
and UO_4434 (O_4434,N_49678,N_49692);
and UO_4435 (O_4435,N_48840,N_49413);
or UO_4436 (O_4436,N_49570,N_49107);
xor UO_4437 (O_4437,N_49835,N_48832);
xor UO_4438 (O_4438,N_49390,N_48333);
or UO_4439 (O_4439,N_49368,N_48094);
or UO_4440 (O_4440,N_48471,N_49280);
nand UO_4441 (O_4441,N_49005,N_49648);
or UO_4442 (O_4442,N_49146,N_49770);
nor UO_4443 (O_4443,N_49797,N_48707);
nor UO_4444 (O_4444,N_49866,N_49269);
nor UO_4445 (O_4445,N_49123,N_49222);
xnor UO_4446 (O_4446,N_48714,N_49646);
or UO_4447 (O_4447,N_48221,N_48690);
xor UO_4448 (O_4448,N_48532,N_48383);
xor UO_4449 (O_4449,N_49584,N_48465);
and UO_4450 (O_4450,N_49890,N_49014);
nand UO_4451 (O_4451,N_48072,N_48884);
xnor UO_4452 (O_4452,N_49495,N_49077);
and UO_4453 (O_4453,N_49273,N_49715);
nand UO_4454 (O_4454,N_48231,N_49761);
and UO_4455 (O_4455,N_48977,N_48440);
and UO_4456 (O_4456,N_48644,N_48295);
nor UO_4457 (O_4457,N_48441,N_48644);
nand UO_4458 (O_4458,N_49775,N_49970);
nand UO_4459 (O_4459,N_48109,N_49640);
nand UO_4460 (O_4460,N_49097,N_49744);
and UO_4461 (O_4461,N_49761,N_49861);
nor UO_4462 (O_4462,N_48855,N_49280);
nand UO_4463 (O_4463,N_48228,N_49153);
xor UO_4464 (O_4464,N_48417,N_48160);
nor UO_4465 (O_4465,N_49920,N_49500);
xnor UO_4466 (O_4466,N_48209,N_49093);
nand UO_4467 (O_4467,N_48007,N_49507);
and UO_4468 (O_4468,N_48165,N_48600);
nor UO_4469 (O_4469,N_49303,N_48359);
or UO_4470 (O_4470,N_48232,N_48287);
nand UO_4471 (O_4471,N_49551,N_48507);
or UO_4472 (O_4472,N_48628,N_48474);
nand UO_4473 (O_4473,N_49065,N_49805);
nor UO_4474 (O_4474,N_49110,N_49983);
and UO_4475 (O_4475,N_49589,N_49908);
nor UO_4476 (O_4476,N_49983,N_49035);
nor UO_4477 (O_4477,N_48602,N_48474);
nor UO_4478 (O_4478,N_48689,N_49718);
or UO_4479 (O_4479,N_48252,N_49671);
and UO_4480 (O_4480,N_48876,N_48724);
nand UO_4481 (O_4481,N_49322,N_48113);
nor UO_4482 (O_4482,N_48200,N_49537);
nor UO_4483 (O_4483,N_48013,N_48299);
nor UO_4484 (O_4484,N_48485,N_49659);
nor UO_4485 (O_4485,N_48143,N_49145);
xnor UO_4486 (O_4486,N_49454,N_48864);
xnor UO_4487 (O_4487,N_49974,N_49498);
and UO_4488 (O_4488,N_48396,N_48472);
or UO_4489 (O_4489,N_48727,N_49596);
nor UO_4490 (O_4490,N_48188,N_48270);
xor UO_4491 (O_4491,N_49003,N_48058);
and UO_4492 (O_4492,N_49621,N_49063);
nor UO_4493 (O_4493,N_48212,N_49254);
nand UO_4494 (O_4494,N_49142,N_49521);
nor UO_4495 (O_4495,N_49362,N_48501);
and UO_4496 (O_4496,N_48134,N_49904);
or UO_4497 (O_4497,N_49842,N_49534);
nand UO_4498 (O_4498,N_48164,N_48661);
xnor UO_4499 (O_4499,N_49618,N_48096);
xnor UO_4500 (O_4500,N_48625,N_49310);
nand UO_4501 (O_4501,N_48884,N_49621);
or UO_4502 (O_4502,N_49477,N_49490);
xnor UO_4503 (O_4503,N_49638,N_48625);
or UO_4504 (O_4504,N_48299,N_48500);
nand UO_4505 (O_4505,N_48256,N_48104);
xnor UO_4506 (O_4506,N_48579,N_48447);
and UO_4507 (O_4507,N_49837,N_49193);
or UO_4508 (O_4508,N_49783,N_49251);
and UO_4509 (O_4509,N_48995,N_48722);
and UO_4510 (O_4510,N_48504,N_49988);
nor UO_4511 (O_4511,N_49989,N_48838);
and UO_4512 (O_4512,N_48202,N_49588);
and UO_4513 (O_4513,N_49912,N_48210);
nand UO_4514 (O_4514,N_48630,N_48642);
nor UO_4515 (O_4515,N_48762,N_48479);
and UO_4516 (O_4516,N_49360,N_48868);
or UO_4517 (O_4517,N_48023,N_49547);
nand UO_4518 (O_4518,N_49424,N_49747);
xnor UO_4519 (O_4519,N_48169,N_48594);
and UO_4520 (O_4520,N_48441,N_49403);
or UO_4521 (O_4521,N_48524,N_48606);
nor UO_4522 (O_4522,N_48662,N_48477);
or UO_4523 (O_4523,N_48312,N_49870);
xor UO_4524 (O_4524,N_48410,N_49870);
xnor UO_4525 (O_4525,N_49704,N_49726);
nor UO_4526 (O_4526,N_49694,N_49559);
nor UO_4527 (O_4527,N_49606,N_48333);
xnor UO_4528 (O_4528,N_49781,N_49785);
and UO_4529 (O_4529,N_49606,N_48815);
nand UO_4530 (O_4530,N_48039,N_49623);
nand UO_4531 (O_4531,N_48242,N_49966);
nand UO_4532 (O_4532,N_49077,N_49926);
or UO_4533 (O_4533,N_48363,N_48119);
nand UO_4534 (O_4534,N_48350,N_49018);
nand UO_4535 (O_4535,N_48574,N_48212);
or UO_4536 (O_4536,N_48961,N_48954);
nor UO_4537 (O_4537,N_49309,N_49040);
nor UO_4538 (O_4538,N_49605,N_49836);
nor UO_4539 (O_4539,N_48464,N_49012);
and UO_4540 (O_4540,N_48960,N_49674);
and UO_4541 (O_4541,N_48804,N_49025);
nor UO_4542 (O_4542,N_49497,N_48197);
xor UO_4543 (O_4543,N_48092,N_48457);
nand UO_4544 (O_4544,N_49417,N_49543);
and UO_4545 (O_4545,N_49171,N_48785);
or UO_4546 (O_4546,N_48201,N_49003);
or UO_4547 (O_4547,N_48864,N_48243);
and UO_4548 (O_4548,N_48946,N_48316);
or UO_4549 (O_4549,N_48331,N_49410);
nand UO_4550 (O_4550,N_49455,N_48135);
and UO_4551 (O_4551,N_48302,N_48656);
nand UO_4552 (O_4552,N_48431,N_49341);
nor UO_4553 (O_4553,N_48925,N_49127);
and UO_4554 (O_4554,N_48757,N_49036);
or UO_4555 (O_4555,N_49252,N_48543);
xor UO_4556 (O_4556,N_48224,N_49546);
nor UO_4557 (O_4557,N_49910,N_49984);
xor UO_4558 (O_4558,N_48776,N_49954);
xnor UO_4559 (O_4559,N_48232,N_49141);
nor UO_4560 (O_4560,N_49339,N_49224);
nand UO_4561 (O_4561,N_48767,N_49309);
xnor UO_4562 (O_4562,N_48982,N_49462);
nand UO_4563 (O_4563,N_49524,N_48816);
xor UO_4564 (O_4564,N_49983,N_49411);
xnor UO_4565 (O_4565,N_49494,N_48876);
nand UO_4566 (O_4566,N_49137,N_48236);
xor UO_4567 (O_4567,N_48032,N_48139);
nand UO_4568 (O_4568,N_49296,N_48320);
nand UO_4569 (O_4569,N_48106,N_49928);
nand UO_4570 (O_4570,N_49064,N_49524);
nor UO_4571 (O_4571,N_49599,N_49165);
or UO_4572 (O_4572,N_49333,N_49929);
nor UO_4573 (O_4573,N_48740,N_48225);
and UO_4574 (O_4574,N_49363,N_48038);
or UO_4575 (O_4575,N_48780,N_49188);
and UO_4576 (O_4576,N_49053,N_48764);
xnor UO_4577 (O_4577,N_49171,N_49008);
nor UO_4578 (O_4578,N_49280,N_49493);
xnor UO_4579 (O_4579,N_49700,N_48683);
or UO_4580 (O_4580,N_48062,N_48871);
and UO_4581 (O_4581,N_48300,N_49858);
nor UO_4582 (O_4582,N_48472,N_49908);
xor UO_4583 (O_4583,N_49867,N_49345);
and UO_4584 (O_4584,N_48081,N_48891);
and UO_4585 (O_4585,N_49195,N_48090);
and UO_4586 (O_4586,N_49524,N_48383);
and UO_4587 (O_4587,N_49449,N_49007);
and UO_4588 (O_4588,N_49524,N_49699);
xor UO_4589 (O_4589,N_48498,N_48664);
and UO_4590 (O_4590,N_48117,N_48313);
nor UO_4591 (O_4591,N_48796,N_49340);
xnor UO_4592 (O_4592,N_49770,N_49166);
xnor UO_4593 (O_4593,N_49783,N_48267);
xnor UO_4594 (O_4594,N_48361,N_49266);
nand UO_4595 (O_4595,N_49781,N_48143);
nor UO_4596 (O_4596,N_49888,N_49726);
xnor UO_4597 (O_4597,N_48883,N_48869);
or UO_4598 (O_4598,N_49714,N_48583);
xnor UO_4599 (O_4599,N_49805,N_48079);
or UO_4600 (O_4600,N_49672,N_48708);
or UO_4601 (O_4601,N_48193,N_49631);
xor UO_4602 (O_4602,N_48743,N_48896);
xor UO_4603 (O_4603,N_49361,N_48707);
and UO_4604 (O_4604,N_48742,N_49149);
nor UO_4605 (O_4605,N_49276,N_48611);
nor UO_4606 (O_4606,N_48080,N_49051);
xor UO_4607 (O_4607,N_49928,N_48621);
nand UO_4608 (O_4608,N_48623,N_48479);
xnor UO_4609 (O_4609,N_49797,N_49904);
nor UO_4610 (O_4610,N_48190,N_48801);
nand UO_4611 (O_4611,N_49086,N_48074);
nor UO_4612 (O_4612,N_48462,N_49481);
xor UO_4613 (O_4613,N_48618,N_49732);
nand UO_4614 (O_4614,N_49455,N_48405);
nor UO_4615 (O_4615,N_49609,N_49566);
and UO_4616 (O_4616,N_49964,N_48962);
or UO_4617 (O_4617,N_48557,N_49332);
nor UO_4618 (O_4618,N_48805,N_48181);
and UO_4619 (O_4619,N_48066,N_48789);
xnor UO_4620 (O_4620,N_49884,N_48032);
or UO_4621 (O_4621,N_48495,N_49661);
nand UO_4622 (O_4622,N_49979,N_48822);
and UO_4623 (O_4623,N_48929,N_48872);
or UO_4624 (O_4624,N_49071,N_49366);
xnor UO_4625 (O_4625,N_48940,N_49454);
xor UO_4626 (O_4626,N_49767,N_48684);
and UO_4627 (O_4627,N_48652,N_49397);
xnor UO_4628 (O_4628,N_48925,N_48379);
nand UO_4629 (O_4629,N_49935,N_49859);
nor UO_4630 (O_4630,N_49814,N_48251);
nand UO_4631 (O_4631,N_49703,N_49795);
xnor UO_4632 (O_4632,N_49675,N_49951);
xor UO_4633 (O_4633,N_49010,N_48845);
nor UO_4634 (O_4634,N_48232,N_48235);
xor UO_4635 (O_4635,N_48122,N_49693);
nand UO_4636 (O_4636,N_48418,N_49977);
nand UO_4637 (O_4637,N_49076,N_49706);
nand UO_4638 (O_4638,N_48046,N_49139);
or UO_4639 (O_4639,N_48949,N_48992);
nand UO_4640 (O_4640,N_48448,N_49174);
xnor UO_4641 (O_4641,N_49742,N_48999);
or UO_4642 (O_4642,N_48485,N_49774);
nor UO_4643 (O_4643,N_49555,N_49155);
or UO_4644 (O_4644,N_48556,N_49237);
nor UO_4645 (O_4645,N_49694,N_48113);
nand UO_4646 (O_4646,N_49311,N_48178);
nor UO_4647 (O_4647,N_49099,N_49271);
xor UO_4648 (O_4648,N_49733,N_49807);
nand UO_4649 (O_4649,N_48408,N_49016);
nor UO_4650 (O_4650,N_48719,N_49039);
nor UO_4651 (O_4651,N_49944,N_49625);
xor UO_4652 (O_4652,N_48295,N_49669);
and UO_4653 (O_4653,N_49400,N_49434);
nor UO_4654 (O_4654,N_48573,N_49461);
or UO_4655 (O_4655,N_48430,N_49804);
and UO_4656 (O_4656,N_49870,N_48694);
xor UO_4657 (O_4657,N_49085,N_49362);
nand UO_4658 (O_4658,N_48681,N_49814);
and UO_4659 (O_4659,N_48895,N_49841);
or UO_4660 (O_4660,N_48317,N_48242);
and UO_4661 (O_4661,N_49493,N_49512);
nand UO_4662 (O_4662,N_49877,N_48082);
nand UO_4663 (O_4663,N_48312,N_49157);
or UO_4664 (O_4664,N_49128,N_49985);
xor UO_4665 (O_4665,N_49844,N_49945);
and UO_4666 (O_4666,N_48917,N_49763);
or UO_4667 (O_4667,N_49502,N_49340);
or UO_4668 (O_4668,N_48771,N_48730);
and UO_4669 (O_4669,N_49367,N_49497);
xor UO_4670 (O_4670,N_49184,N_49583);
xor UO_4671 (O_4671,N_48977,N_49272);
and UO_4672 (O_4672,N_49810,N_48160);
xor UO_4673 (O_4673,N_48960,N_49684);
nand UO_4674 (O_4674,N_48108,N_48694);
or UO_4675 (O_4675,N_49204,N_48438);
or UO_4676 (O_4676,N_49999,N_49743);
nor UO_4677 (O_4677,N_48387,N_49953);
and UO_4678 (O_4678,N_48571,N_48228);
and UO_4679 (O_4679,N_49853,N_49532);
nor UO_4680 (O_4680,N_48348,N_49620);
xnor UO_4681 (O_4681,N_49349,N_48869);
and UO_4682 (O_4682,N_48617,N_48946);
nor UO_4683 (O_4683,N_48810,N_48771);
or UO_4684 (O_4684,N_48857,N_49501);
nor UO_4685 (O_4685,N_49050,N_48151);
nand UO_4686 (O_4686,N_48298,N_48624);
nand UO_4687 (O_4687,N_49320,N_48726);
nand UO_4688 (O_4688,N_48504,N_49574);
or UO_4689 (O_4689,N_49552,N_48761);
xor UO_4690 (O_4690,N_48585,N_48448);
xor UO_4691 (O_4691,N_49121,N_49876);
or UO_4692 (O_4692,N_48989,N_48522);
and UO_4693 (O_4693,N_49359,N_49748);
or UO_4694 (O_4694,N_49155,N_49904);
nand UO_4695 (O_4695,N_49255,N_49356);
nand UO_4696 (O_4696,N_49214,N_49020);
nor UO_4697 (O_4697,N_49260,N_49835);
xor UO_4698 (O_4698,N_49902,N_48170);
nand UO_4699 (O_4699,N_49298,N_48365);
nand UO_4700 (O_4700,N_48165,N_48300);
nand UO_4701 (O_4701,N_49148,N_48301);
xor UO_4702 (O_4702,N_49660,N_48496);
xnor UO_4703 (O_4703,N_48665,N_48796);
nor UO_4704 (O_4704,N_49131,N_49639);
xor UO_4705 (O_4705,N_48257,N_48405);
and UO_4706 (O_4706,N_49599,N_48851);
and UO_4707 (O_4707,N_48010,N_48790);
nand UO_4708 (O_4708,N_48897,N_48843);
or UO_4709 (O_4709,N_49957,N_48625);
nand UO_4710 (O_4710,N_49050,N_48759);
or UO_4711 (O_4711,N_48831,N_48054);
or UO_4712 (O_4712,N_49157,N_49919);
or UO_4713 (O_4713,N_49547,N_49702);
xor UO_4714 (O_4714,N_48390,N_48795);
nor UO_4715 (O_4715,N_48031,N_49312);
or UO_4716 (O_4716,N_48559,N_49741);
nor UO_4717 (O_4717,N_48378,N_49403);
nor UO_4718 (O_4718,N_48129,N_49527);
or UO_4719 (O_4719,N_48400,N_48603);
xor UO_4720 (O_4720,N_49916,N_49433);
or UO_4721 (O_4721,N_48711,N_49104);
xor UO_4722 (O_4722,N_48676,N_49331);
xnor UO_4723 (O_4723,N_49060,N_48659);
nand UO_4724 (O_4724,N_48493,N_49698);
and UO_4725 (O_4725,N_49772,N_48840);
xor UO_4726 (O_4726,N_49621,N_49943);
and UO_4727 (O_4727,N_49291,N_49108);
xor UO_4728 (O_4728,N_49496,N_48553);
nand UO_4729 (O_4729,N_48776,N_48141);
or UO_4730 (O_4730,N_48258,N_48077);
and UO_4731 (O_4731,N_48615,N_48186);
or UO_4732 (O_4732,N_49325,N_49997);
nand UO_4733 (O_4733,N_48022,N_49426);
nor UO_4734 (O_4734,N_48092,N_48142);
nor UO_4735 (O_4735,N_48365,N_49192);
nand UO_4736 (O_4736,N_49152,N_48273);
nor UO_4737 (O_4737,N_48941,N_48205);
xor UO_4738 (O_4738,N_49994,N_48607);
xor UO_4739 (O_4739,N_49807,N_48652);
and UO_4740 (O_4740,N_48829,N_48135);
nor UO_4741 (O_4741,N_48796,N_48547);
nand UO_4742 (O_4742,N_48143,N_49017);
nor UO_4743 (O_4743,N_48388,N_49487);
xor UO_4744 (O_4744,N_48412,N_48822);
or UO_4745 (O_4745,N_49066,N_49502);
and UO_4746 (O_4746,N_49175,N_49458);
or UO_4747 (O_4747,N_49327,N_48826);
nor UO_4748 (O_4748,N_48176,N_48222);
or UO_4749 (O_4749,N_48044,N_49465);
nand UO_4750 (O_4750,N_49801,N_48748);
xor UO_4751 (O_4751,N_48990,N_49086);
nand UO_4752 (O_4752,N_49449,N_49811);
or UO_4753 (O_4753,N_48514,N_49470);
xor UO_4754 (O_4754,N_48604,N_49914);
nor UO_4755 (O_4755,N_49445,N_48183);
or UO_4756 (O_4756,N_49743,N_48998);
xnor UO_4757 (O_4757,N_49459,N_48554);
xor UO_4758 (O_4758,N_49509,N_49834);
or UO_4759 (O_4759,N_49387,N_48823);
nor UO_4760 (O_4760,N_48121,N_49737);
or UO_4761 (O_4761,N_48151,N_49138);
nand UO_4762 (O_4762,N_48735,N_49328);
or UO_4763 (O_4763,N_48024,N_48093);
nand UO_4764 (O_4764,N_49033,N_48362);
nand UO_4765 (O_4765,N_49979,N_49141);
or UO_4766 (O_4766,N_48010,N_48313);
nand UO_4767 (O_4767,N_49527,N_48843);
nand UO_4768 (O_4768,N_49228,N_49126);
nor UO_4769 (O_4769,N_49244,N_49563);
xnor UO_4770 (O_4770,N_48169,N_49354);
and UO_4771 (O_4771,N_49382,N_49939);
or UO_4772 (O_4772,N_48098,N_48581);
and UO_4773 (O_4773,N_48559,N_48172);
xnor UO_4774 (O_4774,N_49399,N_48222);
nor UO_4775 (O_4775,N_49629,N_48890);
or UO_4776 (O_4776,N_48648,N_48216);
or UO_4777 (O_4777,N_48376,N_48635);
and UO_4778 (O_4778,N_48236,N_49731);
xor UO_4779 (O_4779,N_48732,N_48873);
xnor UO_4780 (O_4780,N_48498,N_48355);
or UO_4781 (O_4781,N_48684,N_49628);
nand UO_4782 (O_4782,N_49779,N_49459);
nor UO_4783 (O_4783,N_48026,N_49786);
xnor UO_4784 (O_4784,N_49235,N_49999);
nor UO_4785 (O_4785,N_48493,N_48426);
nor UO_4786 (O_4786,N_49713,N_49755);
xor UO_4787 (O_4787,N_48701,N_48510);
xnor UO_4788 (O_4788,N_48908,N_48526);
and UO_4789 (O_4789,N_48454,N_49634);
and UO_4790 (O_4790,N_49698,N_49627);
nor UO_4791 (O_4791,N_48892,N_48009);
nand UO_4792 (O_4792,N_48006,N_48925);
nand UO_4793 (O_4793,N_49958,N_49525);
nor UO_4794 (O_4794,N_48152,N_48182);
nor UO_4795 (O_4795,N_48522,N_48054);
or UO_4796 (O_4796,N_48982,N_48816);
nor UO_4797 (O_4797,N_48154,N_48379);
and UO_4798 (O_4798,N_48092,N_48648);
nand UO_4799 (O_4799,N_48585,N_48951);
nor UO_4800 (O_4800,N_49982,N_48781);
xor UO_4801 (O_4801,N_48495,N_48646);
and UO_4802 (O_4802,N_48692,N_49053);
xor UO_4803 (O_4803,N_48512,N_49609);
xnor UO_4804 (O_4804,N_49711,N_49191);
xor UO_4805 (O_4805,N_48139,N_48433);
nor UO_4806 (O_4806,N_48614,N_49319);
and UO_4807 (O_4807,N_48698,N_49470);
xor UO_4808 (O_4808,N_49295,N_49714);
or UO_4809 (O_4809,N_48692,N_49522);
or UO_4810 (O_4810,N_49754,N_49718);
nand UO_4811 (O_4811,N_49809,N_48911);
and UO_4812 (O_4812,N_49271,N_49552);
or UO_4813 (O_4813,N_48834,N_48048);
and UO_4814 (O_4814,N_49288,N_48797);
xnor UO_4815 (O_4815,N_48167,N_49465);
nand UO_4816 (O_4816,N_48662,N_48530);
xnor UO_4817 (O_4817,N_48056,N_49431);
nor UO_4818 (O_4818,N_48258,N_49058);
xnor UO_4819 (O_4819,N_49261,N_49172);
nor UO_4820 (O_4820,N_49333,N_49360);
xnor UO_4821 (O_4821,N_48324,N_48176);
xor UO_4822 (O_4822,N_49973,N_49074);
and UO_4823 (O_4823,N_49013,N_48923);
xor UO_4824 (O_4824,N_49004,N_48958);
and UO_4825 (O_4825,N_49995,N_49080);
nand UO_4826 (O_4826,N_49007,N_48588);
nor UO_4827 (O_4827,N_49358,N_49657);
nor UO_4828 (O_4828,N_48339,N_48704);
nand UO_4829 (O_4829,N_49307,N_49187);
nor UO_4830 (O_4830,N_48359,N_48682);
and UO_4831 (O_4831,N_49782,N_49232);
nand UO_4832 (O_4832,N_48474,N_49953);
or UO_4833 (O_4833,N_48993,N_49958);
xor UO_4834 (O_4834,N_49733,N_49380);
and UO_4835 (O_4835,N_48123,N_49544);
nand UO_4836 (O_4836,N_49394,N_49660);
and UO_4837 (O_4837,N_48368,N_48294);
xor UO_4838 (O_4838,N_49017,N_49895);
or UO_4839 (O_4839,N_49237,N_49759);
nor UO_4840 (O_4840,N_49638,N_49954);
xnor UO_4841 (O_4841,N_49416,N_48504);
nor UO_4842 (O_4842,N_49451,N_48428);
and UO_4843 (O_4843,N_49811,N_48710);
nand UO_4844 (O_4844,N_48899,N_49761);
nand UO_4845 (O_4845,N_49803,N_49488);
nand UO_4846 (O_4846,N_48615,N_49069);
nor UO_4847 (O_4847,N_49774,N_49518);
nor UO_4848 (O_4848,N_49389,N_48208);
xnor UO_4849 (O_4849,N_49898,N_48055);
nand UO_4850 (O_4850,N_48934,N_49824);
or UO_4851 (O_4851,N_49082,N_49391);
xor UO_4852 (O_4852,N_48220,N_49121);
nand UO_4853 (O_4853,N_48977,N_49930);
or UO_4854 (O_4854,N_48359,N_48823);
xnor UO_4855 (O_4855,N_48435,N_48058);
nand UO_4856 (O_4856,N_48809,N_48387);
nand UO_4857 (O_4857,N_49739,N_48257);
nand UO_4858 (O_4858,N_49099,N_48132);
nand UO_4859 (O_4859,N_49582,N_48081);
xnor UO_4860 (O_4860,N_48109,N_49539);
xnor UO_4861 (O_4861,N_48865,N_48054);
xor UO_4862 (O_4862,N_48813,N_49905);
and UO_4863 (O_4863,N_48097,N_48325);
and UO_4864 (O_4864,N_49395,N_48034);
and UO_4865 (O_4865,N_48081,N_49390);
or UO_4866 (O_4866,N_48331,N_49921);
and UO_4867 (O_4867,N_48504,N_48717);
nand UO_4868 (O_4868,N_48230,N_49344);
xnor UO_4869 (O_4869,N_48040,N_49368);
nand UO_4870 (O_4870,N_48613,N_49166);
or UO_4871 (O_4871,N_49794,N_49029);
xor UO_4872 (O_4872,N_49906,N_48824);
nand UO_4873 (O_4873,N_49435,N_48387);
or UO_4874 (O_4874,N_48787,N_48233);
nor UO_4875 (O_4875,N_49719,N_49027);
nand UO_4876 (O_4876,N_49499,N_49956);
and UO_4877 (O_4877,N_49734,N_49035);
nand UO_4878 (O_4878,N_49733,N_49531);
xor UO_4879 (O_4879,N_49523,N_48574);
nor UO_4880 (O_4880,N_48335,N_49897);
or UO_4881 (O_4881,N_49270,N_48116);
nor UO_4882 (O_4882,N_48210,N_49634);
or UO_4883 (O_4883,N_49750,N_49213);
or UO_4884 (O_4884,N_48106,N_48911);
and UO_4885 (O_4885,N_49165,N_48238);
nor UO_4886 (O_4886,N_48909,N_49242);
or UO_4887 (O_4887,N_48222,N_49126);
xnor UO_4888 (O_4888,N_48278,N_49914);
nand UO_4889 (O_4889,N_48130,N_48320);
xor UO_4890 (O_4890,N_48491,N_48486);
xor UO_4891 (O_4891,N_49710,N_49805);
or UO_4892 (O_4892,N_48626,N_49034);
or UO_4893 (O_4893,N_49274,N_48927);
or UO_4894 (O_4894,N_48500,N_49992);
or UO_4895 (O_4895,N_48637,N_48265);
nand UO_4896 (O_4896,N_49235,N_48835);
nor UO_4897 (O_4897,N_49865,N_48323);
and UO_4898 (O_4898,N_49406,N_49895);
or UO_4899 (O_4899,N_48150,N_48815);
xor UO_4900 (O_4900,N_48136,N_49914);
nor UO_4901 (O_4901,N_48674,N_49576);
or UO_4902 (O_4902,N_49226,N_49585);
nor UO_4903 (O_4903,N_49099,N_48754);
nor UO_4904 (O_4904,N_49567,N_48384);
xnor UO_4905 (O_4905,N_49041,N_49033);
nor UO_4906 (O_4906,N_49758,N_48236);
nand UO_4907 (O_4907,N_48940,N_49296);
or UO_4908 (O_4908,N_48259,N_48121);
or UO_4909 (O_4909,N_48589,N_49465);
xnor UO_4910 (O_4910,N_49860,N_49011);
xnor UO_4911 (O_4911,N_48920,N_49310);
or UO_4912 (O_4912,N_49534,N_49355);
xnor UO_4913 (O_4913,N_48269,N_49069);
and UO_4914 (O_4914,N_48790,N_49809);
nor UO_4915 (O_4915,N_48998,N_49728);
xnor UO_4916 (O_4916,N_48457,N_48638);
or UO_4917 (O_4917,N_49116,N_48849);
or UO_4918 (O_4918,N_49130,N_49194);
or UO_4919 (O_4919,N_48460,N_49404);
xnor UO_4920 (O_4920,N_48666,N_48735);
xor UO_4921 (O_4921,N_49086,N_48922);
nor UO_4922 (O_4922,N_48336,N_49463);
xnor UO_4923 (O_4923,N_48799,N_48783);
and UO_4924 (O_4924,N_48855,N_49003);
xnor UO_4925 (O_4925,N_49373,N_49832);
and UO_4926 (O_4926,N_49537,N_48592);
or UO_4927 (O_4927,N_48449,N_48863);
and UO_4928 (O_4928,N_48455,N_49597);
and UO_4929 (O_4929,N_49099,N_49148);
nand UO_4930 (O_4930,N_48173,N_49889);
and UO_4931 (O_4931,N_49669,N_49155);
nand UO_4932 (O_4932,N_48739,N_49071);
nand UO_4933 (O_4933,N_49803,N_49653);
or UO_4934 (O_4934,N_49265,N_48603);
or UO_4935 (O_4935,N_48526,N_49285);
nand UO_4936 (O_4936,N_48515,N_48786);
and UO_4937 (O_4937,N_48333,N_49223);
and UO_4938 (O_4938,N_48960,N_48198);
and UO_4939 (O_4939,N_49335,N_49187);
or UO_4940 (O_4940,N_49082,N_49937);
nand UO_4941 (O_4941,N_49842,N_48967);
xor UO_4942 (O_4942,N_49340,N_48833);
or UO_4943 (O_4943,N_48607,N_48749);
nor UO_4944 (O_4944,N_49848,N_49887);
and UO_4945 (O_4945,N_49820,N_49025);
nand UO_4946 (O_4946,N_48618,N_49905);
nand UO_4947 (O_4947,N_49744,N_49712);
and UO_4948 (O_4948,N_48843,N_49270);
or UO_4949 (O_4949,N_49949,N_48679);
or UO_4950 (O_4950,N_48902,N_48897);
xor UO_4951 (O_4951,N_48361,N_49498);
nand UO_4952 (O_4952,N_48963,N_48025);
nor UO_4953 (O_4953,N_49957,N_48164);
and UO_4954 (O_4954,N_48782,N_48883);
nand UO_4955 (O_4955,N_48398,N_49785);
nand UO_4956 (O_4956,N_49886,N_48250);
and UO_4957 (O_4957,N_48766,N_48612);
nor UO_4958 (O_4958,N_48693,N_49576);
nor UO_4959 (O_4959,N_48195,N_48955);
nand UO_4960 (O_4960,N_49201,N_49083);
nand UO_4961 (O_4961,N_49588,N_49797);
and UO_4962 (O_4962,N_49556,N_49439);
or UO_4963 (O_4963,N_48448,N_49857);
and UO_4964 (O_4964,N_49199,N_49446);
nor UO_4965 (O_4965,N_49225,N_48013);
xnor UO_4966 (O_4966,N_48143,N_48117);
xnor UO_4967 (O_4967,N_49078,N_49414);
or UO_4968 (O_4968,N_48061,N_49703);
and UO_4969 (O_4969,N_48459,N_49620);
and UO_4970 (O_4970,N_49555,N_49270);
nand UO_4971 (O_4971,N_48664,N_49223);
nor UO_4972 (O_4972,N_49424,N_49822);
nand UO_4973 (O_4973,N_49277,N_48504);
nand UO_4974 (O_4974,N_49534,N_49850);
xor UO_4975 (O_4975,N_48284,N_49231);
nand UO_4976 (O_4976,N_49099,N_48239);
and UO_4977 (O_4977,N_48000,N_49699);
or UO_4978 (O_4978,N_49596,N_49545);
xor UO_4979 (O_4979,N_49694,N_48431);
nand UO_4980 (O_4980,N_49212,N_48436);
xnor UO_4981 (O_4981,N_48003,N_48367);
and UO_4982 (O_4982,N_48993,N_48090);
and UO_4983 (O_4983,N_48977,N_48795);
nand UO_4984 (O_4984,N_48545,N_48293);
or UO_4985 (O_4985,N_49394,N_49283);
xor UO_4986 (O_4986,N_49929,N_49723);
xnor UO_4987 (O_4987,N_48144,N_49644);
or UO_4988 (O_4988,N_49490,N_49665);
nand UO_4989 (O_4989,N_48792,N_49269);
nand UO_4990 (O_4990,N_48996,N_48267);
and UO_4991 (O_4991,N_49135,N_48533);
and UO_4992 (O_4992,N_49694,N_48463);
xnor UO_4993 (O_4993,N_49989,N_48706);
nor UO_4994 (O_4994,N_49733,N_48902);
xnor UO_4995 (O_4995,N_49040,N_49053);
nand UO_4996 (O_4996,N_49854,N_49604);
nand UO_4997 (O_4997,N_48610,N_49263);
xnor UO_4998 (O_4998,N_48158,N_48011);
nand UO_4999 (O_4999,N_49032,N_49866);
endmodule