module basic_500_3000_500_4_levels_1xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_184,In_42);
and U1 (N_1,In_110,In_328);
nor U2 (N_2,In_457,In_209);
or U3 (N_3,In_473,In_34);
nand U4 (N_4,In_98,In_253);
nand U5 (N_5,In_409,In_484);
and U6 (N_6,In_237,In_337);
nand U7 (N_7,In_300,In_60);
or U8 (N_8,In_3,In_428);
or U9 (N_9,In_367,In_47);
or U10 (N_10,In_234,In_320);
and U11 (N_11,In_412,In_395);
nor U12 (N_12,In_171,In_496);
and U13 (N_13,In_69,In_493);
and U14 (N_14,In_138,In_68);
or U15 (N_15,In_108,In_434);
nor U16 (N_16,In_255,In_393);
nor U17 (N_17,In_453,In_202);
nand U18 (N_18,In_360,In_452);
nand U19 (N_19,In_423,In_93);
and U20 (N_20,In_181,In_21);
nor U21 (N_21,In_100,In_236);
nor U22 (N_22,In_246,In_262);
nor U23 (N_23,In_397,In_9);
and U24 (N_24,In_218,In_230);
nor U25 (N_25,In_4,In_358);
and U26 (N_26,In_144,In_391);
or U27 (N_27,In_425,In_469);
and U28 (N_28,In_329,In_418);
nor U29 (N_29,In_136,In_478);
and U30 (N_30,In_350,In_447);
nor U31 (N_31,In_23,In_207);
or U32 (N_32,In_338,In_497);
nor U33 (N_33,In_30,In_370);
or U34 (N_34,In_201,In_79);
or U35 (N_35,In_390,In_260);
nor U36 (N_36,In_431,In_235);
xnor U37 (N_37,In_58,In_489);
nor U38 (N_38,In_495,In_1);
nand U39 (N_39,In_116,In_420);
nand U40 (N_40,In_129,In_359);
and U41 (N_41,In_17,In_61);
or U42 (N_42,In_128,In_161);
nor U43 (N_43,In_74,In_53);
nor U44 (N_44,In_471,In_429);
nand U45 (N_45,In_339,In_466);
or U46 (N_46,In_52,In_373);
and U47 (N_47,In_156,In_215);
nand U48 (N_48,In_139,In_313);
nor U49 (N_49,In_266,In_118);
nand U50 (N_50,In_309,In_224);
nor U51 (N_51,In_8,In_333);
and U52 (N_52,In_55,In_400);
nor U53 (N_53,In_143,In_430);
nand U54 (N_54,In_459,In_155);
or U55 (N_55,In_342,In_212);
and U56 (N_56,In_112,In_99);
and U57 (N_57,In_270,In_238);
or U58 (N_58,In_46,In_316);
nor U59 (N_59,In_87,In_308);
nor U60 (N_60,In_199,In_140);
or U61 (N_61,In_82,In_56);
nand U62 (N_62,In_221,In_304);
nand U63 (N_63,In_63,In_267);
xnor U64 (N_64,In_323,In_286);
nand U65 (N_65,In_335,In_135);
nor U66 (N_66,In_91,In_51);
or U67 (N_67,In_384,In_205);
and U68 (N_68,In_382,In_402);
and U69 (N_69,In_427,In_18);
or U70 (N_70,In_377,In_88);
nand U71 (N_71,In_330,In_340);
and U72 (N_72,In_276,In_482);
nand U73 (N_73,In_59,In_96);
nor U74 (N_74,In_289,In_164);
nand U75 (N_75,In_374,In_186);
and U76 (N_76,In_232,In_89);
and U77 (N_77,In_449,In_64);
or U78 (N_78,In_33,In_10);
nand U79 (N_79,In_214,In_251);
or U80 (N_80,In_220,In_386);
and U81 (N_81,In_477,In_424);
xnor U82 (N_82,In_470,In_211);
nand U83 (N_83,In_203,In_448);
nor U84 (N_84,In_296,In_239);
nor U85 (N_85,In_62,In_222);
or U86 (N_86,In_70,In_7);
nor U87 (N_87,In_312,In_346);
nor U88 (N_88,In_241,In_403);
nor U89 (N_89,In_258,In_283);
or U90 (N_90,In_273,In_376);
nor U91 (N_91,In_381,In_204);
nand U92 (N_92,In_16,In_41);
nor U93 (N_93,In_76,In_254);
nor U94 (N_94,In_265,In_433);
nand U95 (N_95,In_40,In_455);
nand U96 (N_96,In_122,In_404);
or U97 (N_97,In_364,In_49);
and U98 (N_98,In_375,In_145);
nand U99 (N_99,In_476,In_168);
nand U100 (N_100,In_317,In_446);
nor U101 (N_101,In_292,In_450);
nand U102 (N_102,In_95,In_101);
or U103 (N_103,In_297,In_271);
and U104 (N_104,In_182,In_102);
nand U105 (N_105,In_356,In_278);
and U106 (N_106,In_387,In_32);
or U107 (N_107,In_307,In_27);
and U108 (N_108,In_252,In_28);
and U109 (N_109,In_491,In_78);
nand U110 (N_110,In_75,In_295);
and U111 (N_111,In_405,In_12);
nor U112 (N_112,In_198,In_303);
and U113 (N_113,In_369,In_2);
and U114 (N_114,In_306,In_104);
nor U115 (N_115,In_6,In_5);
nor U116 (N_116,In_465,In_245);
and U117 (N_117,In_157,In_106);
nand U118 (N_118,In_159,In_125);
nand U119 (N_119,In_107,In_322);
nand U120 (N_120,In_352,In_127);
nand U121 (N_121,In_410,In_72);
or U122 (N_122,In_413,In_318);
nand U123 (N_123,In_290,In_77);
or U124 (N_124,In_445,In_229);
nand U125 (N_125,In_490,In_406);
nand U126 (N_126,In_351,In_137);
and U127 (N_127,In_274,In_432);
or U128 (N_128,In_92,In_475);
nor U129 (N_129,In_151,In_26);
or U130 (N_130,In_65,In_353);
or U131 (N_131,In_302,In_389);
and U132 (N_132,In_460,In_486);
or U133 (N_133,In_311,In_472);
and U134 (N_134,In_365,In_256);
or U135 (N_135,In_13,In_268);
and U136 (N_136,In_111,In_385);
nand U137 (N_137,In_275,In_285);
and U138 (N_138,In_379,In_172);
and U139 (N_139,In_105,In_228);
or U140 (N_140,In_325,In_257);
nand U141 (N_141,In_35,In_123);
nand U142 (N_142,In_148,In_399);
nor U143 (N_143,In_345,In_279);
nor U144 (N_144,In_142,In_421);
and U145 (N_145,In_487,In_114);
nand U146 (N_146,In_227,In_174);
or U147 (N_147,In_280,In_305);
nor U148 (N_148,In_250,In_206);
and U149 (N_149,In_354,In_291);
and U150 (N_150,In_210,In_259);
xnor U151 (N_151,In_310,In_187);
nor U152 (N_152,In_494,In_334);
nand U153 (N_153,In_54,In_173);
and U154 (N_154,In_464,In_299);
nor U155 (N_155,In_247,In_176);
nor U156 (N_156,In_463,In_166);
or U157 (N_157,In_492,In_195);
or U158 (N_158,In_371,In_197);
or U159 (N_159,In_192,In_131);
or U160 (N_160,In_348,In_396);
nand U161 (N_161,In_226,In_378);
and U162 (N_162,In_39,In_388);
and U163 (N_163,In_38,In_438);
and U164 (N_164,In_152,In_153);
or U165 (N_165,In_48,In_115);
nand U166 (N_166,In_113,In_163);
nand U167 (N_167,In_217,In_357);
nor U168 (N_168,In_134,In_66);
nor U169 (N_169,In_0,In_499);
and U170 (N_170,In_158,In_474);
and U171 (N_171,In_165,In_347);
nor U172 (N_172,In_480,In_467);
nand U173 (N_173,In_435,In_193);
or U174 (N_174,In_269,In_277);
or U175 (N_175,In_319,In_343);
or U176 (N_176,In_213,In_314);
and U177 (N_177,In_461,In_240);
or U178 (N_178,In_479,In_185);
nor U179 (N_179,In_175,In_194);
or U180 (N_180,In_20,In_31);
nor U181 (N_181,In_415,In_331);
or U182 (N_182,In_398,In_439);
nand U183 (N_183,In_44,In_170);
nand U184 (N_184,In_344,In_14);
nand U185 (N_185,In_109,In_284);
nor U186 (N_186,In_321,In_298);
and U187 (N_187,In_244,In_24);
and U188 (N_188,In_456,In_454);
and U189 (N_189,In_149,In_368);
xnor U190 (N_190,In_301,In_481);
nor U191 (N_191,In_383,In_85);
and U192 (N_192,In_208,In_15);
nor U193 (N_193,In_444,In_200);
nor U194 (N_194,In_401,In_121);
nor U195 (N_195,In_81,In_261);
nor U196 (N_196,In_183,In_191);
nor U197 (N_197,In_332,In_485);
nand U198 (N_198,In_154,In_349);
and U199 (N_199,In_97,In_488);
and U200 (N_200,In_225,In_179);
nand U201 (N_201,In_117,In_130);
nor U202 (N_202,In_160,In_84);
nand U203 (N_203,In_50,In_80);
nor U204 (N_204,In_326,In_242);
nor U205 (N_205,In_189,In_294);
nor U206 (N_206,In_147,In_498);
and U207 (N_207,In_282,In_188);
nand U208 (N_208,In_37,In_223);
or U209 (N_209,In_327,In_19);
nand U210 (N_210,In_141,In_426);
or U211 (N_211,In_462,In_25);
and U212 (N_212,In_441,In_248);
nor U213 (N_213,In_180,In_288);
nand U214 (N_214,In_293,In_440);
nor U215 (N_215,In_436,In_362);
or U216 (N_216,In_380,In_86);
or U217 (N_217,In_249,In_83);
and U218 (N_218,In_90,In_22);
and U219 (N_219,In_57,In_315);
nand U220 (N_220,In_243,In_263);
nor U221 (N_221,In_133,In_196);
nor U222 (N_222,In_407,In_231);
nor U223 (N_223,In_169,In_437);
nand U224 (N_224,In_73,In_272);
and U225 (N_225,In_419,In_411);
or U226 (N_226,In_36,In_150);
nand U227 (N_227,In_119,In_468);
and U228 (N_228,In_408,In_126);
or U229 (N_229,In_363,In_94);
and U230 (N_230,In_71,In_372);
nand U231 (N_231,In_443,In_132);
and U232 (N_232,In_219,In_190);
nor U233 (N_233,In_177,In_287);
nand U234 (N_234,In_103,In_146);
or U235 (N_235,In_120,In_442);
nor U236 (N_236,In_392,In_483);
or U237 (N_237,In_341,In_178);
and U238 (N_238,In_11,In_216);
and U239 (N_239,In_394,In_451);
or U240 (N_240,In_324,In_233);
or U241 (N_241,In_281,In_162);
nor U242 (N_242,In_43,In_414);
or U243 (N_243,In_29,In_417);
or U244 (N_244,In_366,In_355);
and U245 (N_245,In_167,In_45);
and U246 (N_246,In_336,In_458);
nand U247 (N_247,In_416,In_124);
nor U248 (N_248,In_264,In_422);
nor U249 (N_249,In_67,In_361);
or U250 (N_250,In_173,In_482);
or U251 (N_251,In_468,In_138);
xor U252 (N_252,In_122,In_400);
nor U253 (N_253,In_95,In_384);
nor U254 (N_254,In_22,In_391);
nand U255 (N_255,In_81,In_118);
nor U256 (N_256,In_13,In_163);
nand U257 (N_257,In_129,In_231);
nand U258 (N_258,In_30,In_22);
nor U259 (N_259,In_45,In_192);
and U260 (N_260,In_377,In_400);
nor U261 (N_261,In_490,In_475);
nand U262 (N_262,In_223,In_149);
nand U263 (N_263,In_438,In_276);
nand U264 (N_264,In_254,In_154);
nor U265 (N_265,In_16,In_444);
nand U266 (N_266,In_245,In_97);
or U267 (N_267,In_280,In_375);
or U268 (N_268,In_492,In_417);
nor U269 (N_269,In_8,In_319);
or U270 (N_270,In_182,In_81);
nand U271 (N_271,In_148,In_159);
nor U272 (N_272,In_334,In_63);
nand U273 (N_273,In_25,In_110);
and U274 (N_274,In_463,In_344);
nor U275 (N_275,In_449,In_316);
or U276 (N_276,In_309,In_422);
nand U277 (N_277,In_285,In_118);
nor U278 (N_278,In_106,In_499);
and U279 (N_279,In_29,In_129);
or U280 (N_280,In_87,In_68);
nor U281 (N_281,In_284,In_337);
or U282 (N_282,In_359,In_72);
nand U283 (N_283,In_282,In_110);
and U284 (N_284,In_103,In_170);
nand U285 (N_285,In_234,In_417);
nor U286 (N_286,In_43,In_137);
and U287 (N_287,In_354,In_131);
nor U288 (N_288,In_139,In_86);
nand U289 (N_289,In_395,In_19);
and U290 (N_290,In_1,In_169);
nor U291 (N_291,In_402,In_407);
or U292 (N_292,In_488,In_291);
nand U293 (N_293,In_53,In_31);
nor U294 (N_294,In_176,In_350);
nor U295 (N_295,In_289,In_377);
and U296 (N_296,In_211,In_408);
or U297 (N_297,In_247,In_101);
and U298 (N_298,In_64,In_409);
and U299 (N_299,In_320,In_376);
or U300 (N_300,In_284,In_148);
or U301 (N_301,In_143,In_276);
nand U302 (N_302,In_224,In_39);
nand U303 (N_303,In_158,In_251);
nor U304 (N_304,In_58,In_233);
nor U305 (N_305,In_18,In_166);
nor U306 (N_306,In_338,In_484);
and U307 (N_307,In_371,In_169);
or U308 (N_308,In_190,In_384);
nor U309 (N_309,In_224,In_419);
nand U310 (N_310,In_394,In_164);
nand U311 (N_311,In_17,In_151);
nor U312 (N_312,In_31,In_60);
nor U313 (N_313,In_408,In_80);
nor U314 (N_314,In_489,In_311);
nor U315 (N_315,In_223,In_480);
and U316 (N_316,In_134,In_110);
and U317 (N_317,In_272,In_330);
or U318 (N_318,In_409,In_177);
and U319 (N_319,In_457,In_228);
xnor U320 (N_320,In_495,In_42);
nand U321 (N_321,In_313,In_470);
and U322 (N_322,In_385,In_196);
nand U323 (N_323,In_54,In_407);
nand U324 (N_324,In_442,In_225);
nor U325 (N_325,In_25,In_176);
nand U326 (N_326,In_175,In_152);
or U327 (N_327,In_497,In_457);
nor U328 (N_328,In_129,In_393);
nand U329 (N_329,In_344,In_77);
and U330 (N_330,In_359,In_332);
nor U331 (N_331,In_398,In_164);
and U332 (N_332,In_449,In_409);
nor U333 (N_333,In_329,In_70);
and U334 (N_334,In_133,In_257);
or U335 (N_335,In_254,In_183);
and U336 (N_336,In_404,In_217);
nor U337 (N_337,In_156,In_31);
nor U338 (N_338,In_248,In_91);
nand U339 (N_339,In_443,In_304);
nand U340 (N_340,In_444,In_397);
nor U341 (N_341,In_236,In_223);
or U342 (N_342,In_478,In_169);
nand U343 (N_343,In_302,In_292);
nor U344 (N_344,In_422,In_303);
and U345 (N_345,In_141,In_484);
and U346 (N_346,In_218,In_489);
and U347 (N_347,In_140,In_381);
nand U348 (N_348,In_353,In_428);
or U349 (N_349,In_235,In_305);
nor U350 (N_350,In_150,In_126);
nor U351 (N_351,In_312,In_54);
or U352 (N_352,In_285,In_24);
or U353 (N_353,In_466,In_51);
nand U354 (N_354,In_108,In_202);
or U355 (N_355,In_310,In_113);
nor U356 (N_356,In_436,In_56);
and U357 (N_357,In_357,In_272);
nand U358 (N_358,In_177,In_69);
and U359 (N_359,In_460,In_90);
nand U360 (N_360,In_455,In_114);
or U361 (N_361,In_234,In_206);
or U362 (N_362,In_51,In_110);
nor U363 (N_363,In_178,In_66);
and U364 (N_364,In_240,In_125);
and U365 (N_365,In_5,In_54);
and U366 (N_366,In_128,In_92);
and U367 (N_367,In_78,In_323);
nor U368 (N_368,In_403,In_81);
nor U369 (N_369,In_44,In_255);
nand U370 (N_370,In_227,In_476);
and U371 (N_371,In_84,In_64);
and U372 (N_372,In_203,In_388);
or U373 (N_373,In_394,In_358);
nor U374 (N_374,In_286,In_149);
and U375 (N_375,In_125,In_166);
or U376 (N_376,In_80,In_462);
or U377 (N_377,In_325,In_479);
or U378 (N_378,In_256,In_214);
nand U379 (N_379,In_278,In_165);
or U380 (N_380,In_483,In_151);
nand U381 (N_381,In_289,In_21);
xor U382 (N_382,In_233,In_231);
nor U383 (N_383,In_493,In_68);
or U384 (N_384,In_330,In_34);
and U385 (N_385,In_163,In_141);
nor U386 (N_386,In_301,In_87);
nor U387 (N_387,In_367,In_317);
nor U388 (N_388,In_75,In_42);
nand U389 (N_389,In_156,In_20);
or U390 (N_390,In_470,In_145);
and U391 (N_391,In_312,In_498);
or U392 (N_392,In_310,In_452);
and U393 (N_393,In_190,In_445);
nand U394 (N_394,In_304,In_336);
nor U395 (N_395,In_141,In_55);
nand U396 (N_396,In_20,In_455);
and U397 (N_397,In_196,In_12);
nor U398 (N_398,In_183,In_409);
nor U399 (N_399,In_111,In_181);
nand U400 (N_400,In_83,In_287);
nor U401 (N_401,In_0,In_202);
nor U402 (N_402,In_219,In_316);
or U403 (N_403,In_30,In_82);
nand U404 (N_404,In_312,In_301);
nand U405 (N_405,In_423,In_478);
and U406 (N_406,In_11,In_256);
and U407 (N_407,In_111,In_141);
nand U408 (N_408,In_128,In_495);
and U409 (N_409,In_228,In_153);
or U410 (N_410,In_130,In_472);
nand U411 (N_411,In_300,In_55);
or U412 (N_412,In_178,In_339);
nand U413 (N_413,In_371,In_411);
or U414 (N_414,In_221,In_248);
and U415 (N_415,In_455,In_89);
nand U416 (N_416,In_366,In_114);
and U417 (N_417,In_107,In_418);
nor U418 (N_418,In_227,In_90);
nand U419 (N_419,In_149,In_9);
nor U420 (N_420,In_283,In_477);
and U421 (N_421,In_86,In_426);
and U422 (N_422,In_316,In_84);
or U423 (N_423,In_260,In_143);
or U424 (N_424,In_128,In_365);
or U425 (N_425,In_234,In_394);
nand U426 (N_426,In_44,In_204);
nor U427 (N_427,In_306,In_65);
or U428 (N_428,In_412,In_279);
nand U429 (N_429,In_20,In_72);
or U430 (N_430,In_498,In_267);
nand U431 (N_431,In_335,In_482);
nand U432 (N_432,In_34,In_243);
and U433 (N_433,In_195,In_233);
or U434 (N_434,In_348,In_214);
nor U435 (N_435,In_222,In_265);
and U436 (N_436,In_115,In_312);
nor U437 (N_437,In_447,In_324);
nand U438 (N_438,In_35,In_380);
nor U439 (N_439,In_304,In_402);
and U440 (N_440,In_155,In_449);
nand U441 (N_441,In_395,In_411);
and U442 (N_442,In_52,In_228);
xnor U443 (N_443,In_272,In_159);
and U444 (N_444,In_202,In_326);
or U445 (N_445,In_313,In_360);
or U446 (N_446,In_185,In_480);
nand U447 (N_447,In_470,In_358);
nand U448 (N_448,In_15,In_391);
and U449 (N_449,In_383,In_232);
nor U450 (N_450,In_157,In_150);
and U451 (N_451,In_1,In_82);
nor U452 (N_452,In_73,In_454);
nor U453 (N_453,In_382,In_460);
or U454 (N_454,In_266,In_328);
and U455 (N_455,In_102,In_227);
and U456 (N_456,In_382,In_233);
nand U457 (N_457,In_79,In_135);
nand U458 (N_458,In_160,In_240);
nand U459 (N_459,In_71,In_150);
or U460 (N_460,In_394,In_113);
nor U461 (N_461,In_377,In_285);
and U462 (N_462,In_369,In_365);
nor U463 (N_463,In_153,In_315);
or U464 (N_464,In_446,In_171);
or U465 (N_465,In_243,In_213);
nand U466 (N_466,In_407,In_427);
nor U467 (N_467,In_100,In_222);
nor U468 (N_468,In_233,In_133);
nand U469 (N_469,In_85,In_342);
or U470 (N_470,In_337,In_21);
nand U471 (N_471,In_436,In_8);
nand U472 (N_472,In_478,In_1);
nor U473 (N_473,In_252,In_355);
and U474 (N_474,In_403,In_355);
or U475 (N_475,In_246,In_22);
nor U476 (N_476,In_161,In_52);
nand U477 (N_477,In_481,In_9);
nand U478 (N_478,In_429,In_491);
nand U479 (N_479,In_29,In_356);
nand U480 (N_480,In_320,In_329);
and U481 (N_481,In_456,In_307);
or U482 (N_482,In_465,In_87);
and U483 (N_483,In_208,In_44);
and U484 (N_484,In_234,In_26);
or U485 (N_485,In_200,In_389);
and U486 (N_486,In_152,In_42);
nor U487 (N_487,In_202,In_107);
or U488 (N_488,In_418,In_259);
nand U489 (N_489,In_73,In_143);
and U490 (N_490,In_287,In_10);
and U491 (N_491,In_491,In_444);
nor U492 (N_492,In_486,In_173);
nand U493 (N_493,In_7,In_375);
nor U494 (N_494,In_335,In_27);
and U495 (N_495,In_212,In_75);
nand U496 (N_496,In_263,In_382);
or U497 (N_497,In_380,In_139);
or U498 (N_498,In_160,In_59);
nor U499 (N_499,In_371,In_405);
or U500 (N_500,In_270,In_315);
nand U501 (N_501,In_361,In_282);
nand U502 (N_502,In_155,In_317);
nor U503 (N_503,In_451,In_323);
or U504 (N_504,In_268,In_443);
and U505 (N_505,In_105,In_109);
and U506 (N_506,In_22,In_441);
nor U507 (N_507,In_19,In_134);
xnor U508 (N_508,In_218,In_332);
nand U509 (N_509,In_139,In_208);
nor U510 (N_510,In_136,In_4);
or U511 (N_511,In_477,In_131);
or U512 (N_512,In_151,In_249);
nand U513 (N_513,In_341,In_139);
and U514 (N_514,In_338,In_262);
and U515 (N_515,In_138,In_33);
nor U516 (N_516,In_354,In_372);
nand U517 (N_517,In_81,In_444);
nand U518 (N_518,In_4,In_285);
and U519 (N_519,In_38,In_408);
nor U520 (N_520,In_462,In_325);
nand U521 (N_521,In_471,In_176);
nor U522 (N_522,In_232,In_171);
and U523 (N_523,In_324,In_323);
and U524 (N_524,In_296,In_149);
nor U525 (N_525,In_243,In_424);
and U526 (N_526,In_476,In_370);
nand U527 (N_527,In_346,In_276);
or U528 (N_528,In_153,In_318);
or U529 (N_529,In_317,In_351);
and U530 (N_530,In_249,In_174);
and U531 (N_531,In_63,In_129);
and U532 (N_532,In_331,In_194);
or U533 (N_533,In_240,In_420);
and U534 (N_534,In_61,In_330);
nor U535 (N_535,In_270,In_40);
or U536 (N_536,In_480,In_443);
or U537 (N_537,In_163,In_463);
nand U538 (N_538,In_296,In_242);
or U539 (N_539,In_128,In_416);
or U540 (N_540,In_83,In_283);
nand U541 (N_541,In_122,In_300);
nor U542 (N_542,In_53,In_202);
or U543 (N_543,In_115,In_128);
or U544 (N_544,In_496,In_72);
nor U545 (N_545,In_464,In_207);
or U546 (N_546,In_93,In_124);
or U547 (N_547,In_58,In_406);
or U548 (N_548,In_294,In_85);
nand U549 (N_549,In_146,In_60);
or U550 (N_550,In_471,In_424);
and U551 (N_551,In_209,In_322);
and U552 (N_552,In_4,In_207);
nand U553 (N_553,In_243,In_482);
nor U554 (N_554,In_461,In_85);
or U555 (N_555,In_198,In_201);
nor U556 (N_556,In_297,In_187);
nor U557 (N_557,In_450,In_397);
nand U558 (N_558,In_328,In_238);
nand U559 (N_559,In_286,In_266);
nor U560 (N_560,In_122,In_407);
and U561 (N_561,In_14,In_392);
or U562 (N_562,In_231,In_92);
nor U563 (N_563,In_460,In_333);
nand U564 (N_564,In_120,In_98);
and U565 (N_565,In_60,In_169);
or U566 (N_566,In_53,In_359);
nand U567 (N_567,In_95,In_135);
or U568 (N_568,In_194,In_308);
or U569 (N_569,In_478,In_134);
nand U570 (N_570,In_222,In_359);
or U571 (N_571,In_10,In_55);
or U572 (N_572,In_491,In_303);
and U573 (N_573,In_227,In_365);
or U574 (N_574,In_92,In_165);
nor U575 (N_575,In_133,In_340);
and U576 (N_576,In_456,In_332);
or U577 (N_577,In_391,In_123);
nor U578 (N_578,In_437,In_265);
nor U579 (N_579,In_242,In_51);
nor U580 (N_580,In_404,In_341);
or U581 (N_581,In_345,In_92);
and U582 (N_582,In_87,In_131);
nand U583 (N_583,In_412,In_78);
nor U584 (N_584,In_244,In_100);
and U585 (N_585,In_83,In_407);
and U586 (N_586,In_101,In_39);
nand U587 (N_587,In_73,In_252);
nand U588 (N_588,In_280,In_322);
and U589 (N_589,In_274,In_141);
nor U590 (N_590,In_209,In_363);
and U591 (N_591,In_282,In_494);
and U592 (N_592,In_492,In_34);
or U593 (N_593,In_394,In_285);
nand U594 (N_594,In_491,In_439);
nor U595 (N_595,In_194,In_312);
and U596 (N_596,In_368,In_118);
or U597 (N_597,In_270,In_24);
nor U598 (N_598,In_269,In_384);
or U599 (N_599,In_66,In_382);
nand U600 (N_600,In_494,In_495);
and U601 (N_601,In_108,In_211);
nor U602 (N_602,In_407,In_91);
nor U603 (N_603,In_87,In_88);
nand U604 (N_604,In_175,In_5);
or U605 (N_605,In_409,In_95);
nor U606 (N_606,In_90,In_459);
nand U607 (N_607,In_255,In_337);
and U608 (N_608,In_485,In_127);
nand U609 (N_609,In_79,In_189);
nand U610 (N_610,In_81,In_104);
nand U611 (N_611,In_318,In_128);
and U612 (N_612,In_381,In_42);
nand U613 (N_613,In_135,In_129);
and U614 (N_614,In_158,In_234);
or U615 (N_615,In_411,In_150);
or U616 (N_616,In_225,In_385);
nor U617 (N_617,In_243,In_150);
or U618 (N_618,In_203,In_400);
nand U619 (N_619,In_348,In_10);
nor U620 (N_620,In_408,In_425);
nand U621 (N_621,In_369,In_115);
nor U622 (N_622,In_148,In_301);
nor U623 (N_623,In_308,In_124);
and U624 (N_624,In_423,In_77);
or U625 (N_625,In_216,In_116);
or U626 (N_626,In_462,In_269);
or U627 (N_627,In_450,In_460);
nor U628 (N_628,In_240,In_93);
nand U629 (N_629,In_424,In_183);
nor U630 (N_630,In_380,In_392);
or U631 (N_631,In_400,In_485);
and U632 (N_632,In_106,In_472);
nor U633 (N_633,In_453,In_334);
and U634 (N_634,In_261,In_431);
or U635 (N_635,In_178,In_89);
nand U636 (N_636,In_80,In_34);
or U637 (N_637,In_32,In_209);
nor U638 (N_638,In_448,In_222);
or U639 (N_639,In_472,In_217);
nand U640 (N_640,In_120,In_395);
nor U641 (N_641,In_447,In_352);
nor U642 (N_642,In_48,In_246);
nor U643 (N_643,In_127,In_268);
nor U644 (N_644,In_49,In_299);
and U645 (N_645,In_183,In_496);
nand U646 (N_646,In_194,In_37);
and U647 (N_647,In_226,In_390);
nand U648 (N_648,In_167,In_328);
or U649 (N_649,In_52,In_213);
or U650 (N_650,In_170,In_429);
nor U651 (N_651,In_229,In_112);
and U652 (N_652,In_499,In_232);
nor U653 (N_653,In_193,In_39);
and U654 (N_654,In_270,In_495);
nor U655 (N_655,In_280,In_453);
or U656 (N_656,In_7,In_469);
nand U657 (N_657,In_278,In_36);
and U658 (N_658,In_121,In_102);
nand U659 (N_659,In_285,In_95);
nand U660 (N_660,In_180,In_34);
and U661 (N_661,In_307,In_236);
and U662 (N_662,In_167,In_221);
nand U663 (N_663,In_200,In_376);
nor U664 (N_664,In_408,In_267);
nand U665 (N_665,In_286,In_473);
and U666 (N_666,In_292,In_154);
nor U667 (N_667,In_468,In_170);
nand U668 (N_668,In_182,In_499);
or U669 (N_669,In_392,In_195);
nand U670 (N_670,In_114,In_207);
or U671 (N_671,In_215,In_10);
nor U672 (N_672,In_205,In_116);
nand U673 (N_673,In_319,In_382);
or U674 (N_674,In_446,In_13);
or U675 (N_675,In_116,In_394);
nand U676 (N_676,In_268,In_331);
and U677 (N_677,In_81,In_245);
or U678 (N_678,In_74,In_68);
or U679 (N_679,In_428,In_134);
nand U680 (N_680,In_336,In_383);
and U681 (N_681,In_494,In_486);
nor U682 (N_682,In_192,In_436);
nand U683 (N_683,In_321,In_404);
nor U684 (N_684,In_385,In_156);
and U685 (N_685,In_461,In_43);
and U686 (N_686,In_238,In_268);
and U687 (N_687,In_420,In_353);
nor U688 (N_688,In_240,In_76);
and U689 (N_689,In_58,In_317);
nand U690 (N_690,In_484,In_82);
nand U691 (N_691,In_415,In_316);
nor U692 (N_692,In_465,In_444);
and U693 (N_693,In_28,In_469);
nand U694 (N_694,In_8,In_180);
and U695 (N_695,In_100,In_246);
and U696 (N_696,In_38,In_274);
nand U697 (N_697,In_497,In_20);
nor U698 (N_698,In_333,In_89);
or U699 (N_699,In_197,In_117);
nand U700 (N_700,In_120,In_67);
or U701 (N_701,In_461,In_40);
nor U702 (N_702,In_85,In_238);
nand U703 (N_703,In_51,In_109);
nand U704 (N_704,In_462,In_72);
nor U705 (N_705,In_192,In_308);
and U706 (N_706,In_26,In_266);
or U707 (N_707,In_466,In_190);
nand U708 (N_708,In_396,In_452);
nor U709 (N_709,In_394,In_48);
nand U710 (N_710,In_477,In_197);
nand U711 (N_711,In_56,In_235);
nand U712 (N_712,In_59,In_182);
or U713 (N_713,In_339,In_480);
nor U714 (N_714,In_378,In_5);
nor U715 (N_715,In_148,In_493);
nand U716 (N_716,In_305,In_317);
nand U717 (N_717,In_287,In_434);
nand U718 (N_718,In_130,In_233);
nor U719 (N_719,In_25,In_113);
or U720 (N_720,In_468,In_213);
and U721 (N_721,In_467,In_298);
and U722 (N_722,In_442,In_492);
or U723 (N_723,In_286,In_253);
nor U724 (N_724,In_244,In_276);
nor U725 (N_725,In_354,In_424);
and U726 (N_726,In_263,In_104);
and U727 (N_727,In_156,In_431);
and U728 (N_728,In_301,In_176);
and U729 (N_729,In_417,In_433);
and U730 (N_730,In_492,In_477);
and U731 (N_731,In_123,In_167);
nand U732 (N_732,In_305,In_166);
nand U733 (N_733,In_398,In_246);
nor U734 (N_734,In_230,In_65);
or U735 (N_735,In_275,In_178);
nand U736 (N_736,In_45,In_297);
and U737 (N_737,In_497,In_464);
or U738 (N_738,In_284,In_488);
nand U739 (N_739,In_368,In_259);
nor U740 (N_740,In_427,In_99);
nand U741 (N_741,In_299,In_325);
or U742 (N_742,In_377,In_246);
nand U743 (N_743,In_422,In_409);
nand U744 (N_744,In_214,In_70);
nor U745 (N_745,In_36,In_280);
nand U746 (N_746,In_314,In_397);
nor U747 (N_747,In_310,In_334);
nand U748 (N_748,In_42,In_424);
nand U749 (N_749,In_74,In_109);
nor U750 (N_750,N_739,N_736);
nor U751 (N_751,N_330,N_737);
or U752 (N_752,N_6,N_68);
nand U753 (N_753,N_199,N_706);
or U754 (N_754,N_2,N_118);
or U755 (N_755,N_48,N_448);
or U756 (N_756,N_749,N_502);
and U757 (N_757,N_597,N_27);
nand U758 (N_758,N_434,N_120);
or U759 (N_759,N_315,N_506);
nand U760 (N_760,N_373,N_523);
or U761 (N_761,N_296,N_300);
or U762 (N_762,N_656,N_267);
nand U763 (N_763,N_198,N_620);
nor U764 (N_764,N_741,N_472);
or U765 (N_765,N_224,N_624);
or U766 (N_766,N_457,N_388);
nand U767 (N_767,N_39,N_318);
or U768 (N_768,N_596,N_602);
and U769 (N_769,N_274,N_676);
nand U770 (N_770,N_15,N_397);
nor U771 (N_771,N_137,N_7);
nor U772 (N_772,N_566,N_567);
or U773 (N_773,N_69,N_44);
and U774 (N_774,N_347,N_240);
nand U775 (N_775,N_356,N_541);
and U776 (N_776,N_495,N_108);
and U777 (N_777,N_217,N_212);
or U778 (N_778,N_192,N_278);
nor U779 (N_779,N_17,N_526);
and U780 (N_780,N_282,N_687);
nor U781 (N_781,N_555,N_497);
or U782 (N_782,N_579,N_134);
or U783 (N_783,N_586,N_420);
or U784 (N_784,N_3,N_115);
nor U785 (N_785,N_360,N_312);
nor U786 (N_786,N_548,N_626);
nand U787 (N_787,N_462,N_600);
nand U788 (N_788,N_400,N_326);
nor U789 (N_789,N_38,N_234);
nand U790 (N_790,N_691,N_371);
nor U791 (N_791,N_437,N_179);
and U792 (N_792,N_631,N_726);
or U793 (N_793,N_511,N_237);
and U794 (N_794,N_636,N_501);
nor U795 (N_795,N_452,N_94);
or U796 (N_796,N_510,N_389);
nor U797 (N_797,N_30,N_475);
and U798 (N_798,N_712,N_677);
or U799 (N_799,N_396,N_77);
and U800 (N_800,N_374,N_359);
or U801 (N_801,N_430,N_67);
nor U802 (N_802,N_305,N_669);
nor U803 (N_803,N_554,N_393);
nand U804 (N_804,N_365,N_191);
nand U805 (N_805,N_223,N_262);
nand U806 (N_806,N_288,N_163);
nor U807 (N_807,N_625,N_58);
or U808 (N_808,N_114,N_0);
nand U809 (N_809,N_246,N_28);
nor U810 (N_810,N_429,N_717);
or U811 (N_811,N_498,N_244);
nand U812 (N_812,N_560,N_439);
nand U813 (N_813,N_524,N_387);
and U814 (N_814,N_5,N_682);
and U815 (N_815,N_230,N_194);
and U816 (N_816,N_401,N_195);
or U817 (N_817,N_641,N_556);
nand U818 (N_818,N_723,N_404);
and U819 (N_819,N_173,N_500);
and U820 (N_820,N_285,N_344);
nand U821 (N_821,N_153,N_31);
and U822 (N_822,N_93,N_536);
nand U823 (N_823,N_508,N_61);
or U824 (N_824,N_86,N_418);
or U825 (N_825,N_352,N_152);
nor U826 (N_826,N_346,N_241);
nor U827 (N_827,N_692,N_612);
and U828 (N_828,N_126,N_391);
and U829 (N_829,N_689,N_422);
or U830 (N_830,N_369,N_84);
or U831 (N_831,N_317,N_445);
or U832 (N_832,N_202,N_379);
nand U833 (N_833,N_257,N_189);
nor U834 (N_834,N_181,N_154);
and U835 (N_835,N_129,N_14);
or U836 (N_836,N_187,N_663);
nand U837 (N_837,N_482,N_34);
nor U838 (N_838,N_539,N_29);
or U839 (N_839,N_99,N_286);
and U840 (N_840,N_405,N_688);
or U841 (N_841,N_458,N_245);
nand U842 (N_842,N_722,N_719);
nor U843 (N_843,N_307,N_518);
and U844 (N_844,N_178,N_188);
nand U845 (N_845,N_732,N_563);
or U846 (N_846,N_182,N_208);
nand U847 (N_847,N_639,N_43);
nand U848 (N_848,N_313,N_728);
and U849 (N_849,N_538,N_491);
or U850 (N_850,N_644,N_440);
or U851 (N_851,N_331,N_680);
or U852 (N_852,N_664,N_570);
nand U853 (N_853,N_564,N_604);
nand U854 (N_854,N_243,N_522);
nand U855 (N_855,N_339,N_714);
or U856 (N_856,N_258,N_247);
or U857 (N_857,N_529,N_213);
or U858 (N_858,N_415,N_532);
xor U859 (N_859,N_253,N_47);
and U860 (N_860,N_551,N_444);
and U861 (N_861,N_40,N_255);
nor U862 (N_862,N_725,N_711);
nor U863 (N_863,N_474,N_207);
or U864 (N_864,N_531,N_436);
or U865 (N_865,N_337,N_470);
nor U866 (N_866,N_228,N_362);
nor U867 (N_867,N_321,N_49);
nand U868 (N_868,N_112,N_643);
nor U869 (N_869,N_411,N_589);
nor U870 (N_870,N_568,N_138);
or U871 (N_871,N_746,N_708);
nor U872 (N_872,N_464,N_384);
and U873 (N_873,N_649,N_157);
and U874 (N_874,N_629,N_608);
nor U875 (N_875,N_351,N_176);
nand U876 (N_876,N_606,N_594);
or U877 (N_877,N_599,N_252);
or U878 (N_878,N_345,N_578);
nand U879 (N_879,N_562,N_239);
nor U880 (N_880,N_55,N_242);
nor U881 (N_881,N_268,N_698);
and U882 (N_882,N_561,N_638);
and U883 (N_883,N_250,N_75);
nand U884 (N_884,N_26,N_103);
nor U885 (N_885,N_336,N_302);
and U886 (N_886,N_665,N_184);
or U887 (N_887,N_130,N_168);
nor U888 (N_888,N_13,N_299);
nor U889 (N_889,N_316,N_21);
or U890 (N_890,N_20,N_503);
nor U891 (N_891,N_180,N_450);
or U892 (N_892,N_530,N_701);
or U893 (N_893,N_304,N_477);
nor U894 (N_894,N_117,N_324);
nor U895 (N_895,N_715,N_100);
nand U896 (N_896,N_167,N_459);
nand U897 (N_897,N_19,N_583);
nor U898 (N_898,N_341,N_332);
nand U899 (N_899,N_696,N_489);
and U900 (N_900,N_185,N_280);
or U901 (N_901,N_361,N_709);
nand U902 (N_902,N_54,N_71);
nand U903 (N_903,N_627,N_421);
or U904 (N_904,N_158,N_205);
and U905 (N_905,N_73,N_232);
and U906 (N_906,N_367,N_327);
nor U907 (N_907,N_291,N_544);
nand U908 (N_908,N_509,N_16);
nand U909 (N_909,N_517,N_174);
nand U910 (N_910,N_618,N_322);
xnor U911 (N_911,N_534,N_140);
nand U912 (N_912,N_710,N_479);
and U913 (N_913,N_628,N_478);
nor U914 (N_914,N_273,N_150);
nand U915 (N_915,N_289,N_201);
nor U916 (N_916,N_171,N_357);
nor U917 (N_917,N_309,N_319);
nor U918 (N_918,N_281,N_520);
and U919 (N_919,N_219,N_528);
nor U920 (N_920,N_424,N_146);
or U921 (N_921,N_175,N_582);
or U922 (N_922,N_702,N_220);
nor U923 (N_923,N_549,N_122);
and U924 (N_924,N_206,N_496);
xor U925 (N_925,N_661,N_662);
or U926 (N_926,N_674,N_64);
or U927 (N_927,N_413,N_558);
and U928 (N_928,N_571,N_377);
and U929 (N_929,N_169,N_637);
nor U930 (N_930,N_233,N_235);
and U931 (N_931,N_634,N_366);
nand U932 (N_932,N_729,N_90);
or U933 (N_933,N_8,N_101);
and U934 (N_934,N_260,N_368);
and U935 (N_935,N_587,N_92);
xnor U936 (N_936,N_325,N_514);
nor U937 (N_937,N_720,N_264);
and U938 (N_938,N_652,N_666);
nor U939 (N_939,N_190,N_142);
or U940 (N_940,N_236,N_121);
or U941 (N_941,N_53,N_623);
and U942 (N_942,N_699,N_298);
or U943 (N_943,N_588,N_395);
nor U944 (N_944,N_516,N_686);
or U945 (N_945,N_455,N_46);
nor U946 (N_946,N_416,N_406);
or U947 (N_947,N_461,N_227);
nand U948 (N_948,N_540,N_569);
or U949 (N_949,N_573,N_585);
and U950 (N_950,N_675,N_734);
or U951 (N_951,N_106,N_743);
nand U952 (N_952,N_667,N_287);
nand U953 (N_953,N_82,N_590);
nor U954 (N_954,N_1,N_438);
nor U955 (N_955,N_25,N_673);
nor U956 (N_956,N_527,N_276);
or U957 (N_957,N_139,N_22);
or U958 (N_958,N_601,N_607);
and U959 (N_959,N_671,N_290);
and U960 (N_960,N_441,N_454);
nand U961 (N_961,N_269,N_37);
nor U962 (N_962,N_159,N_172);
nand U963 (N_963,N_12,N_333);
and U964 (N_964,N_403,N_149);
and U965 (N_965,N_50,N_745);
nand U966 (N_966,N_226,N_132);
or U967 (N_967,N_216,N_125);
and U968 (N_968,N_731,N_694);
nand U969 (N_969,N_595,N_493);
nand U970 (N_970,N_363,N_613);
or U971 (N_971,N_266,N_135);
or U972 (N_972,N_412,N_229);
nor U973 (N_973,N_480,N_66);
or U974 (N_974,N_128,N_88);
or U975 (N_975,N_303,N_72);
nor U976 (N_976,N_147,N_721);
nand U977 (N_977,N_133,N_593);
nand U978 (N_978,N_577,N_654);
nor U979 (N_979,N_463,N_402);
nor U980 (N_980,N_695,N_151);
or U981 (N_981,N_398,N_297);
nand U982 (N_982,N_512,N_107);
nor U983 (N_983,N_301,N_645);
and U984 (N_984,N_89,N_483);
and U985 (N_985,N_204,N_700);
nand U986 (N_986,N_385,N_542);
or U987 (N_987,N_515,N_633);
nand U988 (N_988,N_308,N_200);
nor U989 (N_989,N_225,N_60);
or U990 (N_990,N_724,N_85);
or U991 (N_991,N_622,N_408);
nor U992 (N_992,N_113,N_553);
or U993 (N_993,N_443,N_131);
nand U994 (N_994,N_707,N_328);
and U995 (N_995,N_96,N_490);
nor U996 (N_996,N_610,N_136);
nor U997 (N_997,N_41,N_148);
nand U998 (N_998,N_78,N_653);
or U999 (N_999,N_466,N_611);
nor U1000 (N_1000,N_432,N_292);
and U1001 (N_1001,N_414,N_730);
or U1002 (N_1002,N_81,N_59);
or U1003 (N_1003,N_460,N_575);
nand U1004 (N_1004,N_314,N_294);
nand U1005 (N_1005,N_533,N_630);
nand U1006 (N_1006,N_42,N_592);
or U1007 (N_1007,N_660,N_183);
and U1008 (N_1008,N_433,N_487);
or U1009 (N_1009,N_355,N_162);
or U1010 (N_1010,N_380,N_231);
and U1011 (N_1011,N_295,N_119);
or U1012 (N_1012,N_218,N_358);
or U1013 (N_1013,N_565,N_476);
or U1014 (N_1014,N_605,N_581);
nor U1015 (N_1015,N_143,N_427);
or U1016 (N_1016,N_350,N_488);
nor U1017 (N_1017,N_650,N_431);
or U1018 (N_1018,N_453,N_335);
nand U1019 (N_1019,N_259,N_716);
nor U1020 (N_1020,N_256,N_283);
nor U1021 (N_1021,N_394,N_632);
or U1022 (N_1022,N_354,N_284);
nand U1023 (N_1023,N_83,N_616);
or U1024 (N_1024,N_580,N_382);
nor U1025 (N_1025,N_697,N_272);
nor U1026 (N_1026,N_423,N_197);
nand U1027 (N_1027,N_545,N_576);
or U1028 (N_1028,N_505,N_95);
nor U1029 (N_1029,N_123,N_51);
and U1030 (N_1030,N_145,N_619);
and U1031 (N_1031,N_672,N_504);
nor U1032 (N_1032,N_648,N_494);
and U1033 (N_1033,N_141,N_33);
and U1034 (N_1034,N_353,N_467);
and U1035 (N_1035,N_447,N_468);
and U1036 (N_1036,N_690,N_409);
and U1037 (N_1037,N_484,N_747);
and U1038 (N_1038,N_98,N_546);
or U1039 (N_1039,N_693,N_383);
nor U1040 (N_1040,N_407,N_486);
nand U1041 (N_1041,N_24,N_342);
nor U1042 (N_1042,N_559,N_340);
nor U1043 (N_1043,N_111,N_647);
nor U1044 (N_1044,N_547,N_70);
and U1045 (N_1045,N_214,N_525);
nand U1046 (N_1046,N_733,N_727);
and U1047 (N_1047,N_519,N_584);
and U1048 (N_1048,N_23,N_456);
nand U1049 (N_1049,N_63,N_215);
or U1050 (N_1050,N_557,N_210);
or U1051 (N_1051,N_9,N_10);
or U1052 (N_1052,N_364,N_473);
xor U1053 (N_1053,N_271,N_97);
nor U1054 (N_1054,N_62,N_221);
or U1055 (N_1055,N_165,N_376);
and U1056 (N_1056,N_18,N_196);
and U1057 (N_1057,N_381,N_704);
or U1058 (N_1058,N_343,N_646);
or U1059 (N_1059,N_57,N_426);
xor U1060 (N_1060,N_4,N_678);
nand U1061 (N_1061,N_572,N_32);
or U1062 (N_1062,N_378,N_742);
and U1063 (N_1063,N_386,N_670);
nand U1064 (N_1064,N_499,N_471);
nor U1065 (N_1065,N_744,N_249);
or U1066 (N_1066,N_311,N_375);
nor U1067 (N_1067,N_211,N_160);
and U1068 (N_1068,N_684,N_79);
nor U1069 (N_1069,N_451,N_659);
nand U1070 (N_1070,N_655,N_261);
and U1071 (N_1071,N_177,N_203);
or U1072 (N_1072,N_338,N_76);
or U1073 (N_1073,N_615,N_598);
nand U1074 (N_1074,N_507,N_668);
and U1075 (N_1075,N_435,N_657);
or U1076 (N_1076,N_640,N_102);
nand U1077 (N_1077,N_293,N_683);
xnor U1078 (N_1078,N_251,N_469);
nor U1079 (N_1079,N_537,N_552);
and U1080 (N_1080,N_428,N_87);
nand U1081 (N_1081,N_574,N_535);
or U1082 (N_1082,N_193,N_718);
nor U1083 (N_1083,N_161,N_617);
or U1084 (N_1084,N_110,N_446);
and U1085 (N_1085,N_170,N_277);
and U1086 (N_1086,N_209,N_442);
or U1087 (N_1087,N_609,N_91);
nand U1088 (N_1088,N_155,N_329);
or U1089 (N_1089,N_306,N_323);
and U1090 (N_1090,N_614,N_425);
and U1091 (N_1091,N_74,N_166);
and U1092 (N_1092,N_703,N_45);
nand U1093 (N_1093,N_348,N_679);
nor U1094 (N_1094,N_449,N_104);
nor U1095 (N_1095,N_513,N_658);
nor U1096 (N_1096,N_635,N_65);
nor U1097 (N_1097,N_399,N_334);
and U1098 (N_1098,N_521,N_238);
nand U1099 (N_1099,N_705,N_35);
and U1100 (N_1100,N_410,N_310);
nand U1101 (N_1101,N_320,N_279);
or U1102 (N_1102,N_127,N_349);
and U1103 (N_1103,N_265,N_685);
nor U1104 (N_1104,N_56,N_481);
or U1105 (N_1105,N_738,N_492);
nor U1106 (N_1106,N_124,N_417);
or U1107 (N_1107,N_222,N_144);
nor U1108 (N_1108,N_36,N_11);
or U1109 (N_1109,N_80,N_651);
nand U1110 (N_1110,N_392,N_186);
nand U1111 (N_1111,N_390,N_270);
and U1112 (N_1112,N_164,N_254);
nand U1113 (N_1113,N_105,N_275);
nand U1114 (N_1114,N_681,N_485);
or U1115 (N_1115,N_465,N_603);
or U1116 (N_1116,N_156,N_109);
or U1117 (N_1117,N_543,N_419);
nand U1118 (N_1118,N_642,N_735);
and U1119 (N_1119,N_591,N_248);
or U1120 (N_1120,N_263,N_748);
nand U1121 (N_1121,N_116,N_621);
and U1122 (N_1122,N_740,N_713);
and U1123 (N_1123,N_52,N_550);
nor U1124 (N_1124,N_372,N_370);
nor U1125 (N_1125,N_62,N_369);
nor U1126 (N_1126,N_494,N_426);
or U1127 (N_1127,N_566,N_726);
nor U1128 (N_1128,N_713,N_684);
and U1129 (N_1129,N_486,N_747);
or U1130 (N_1130,N_712,N_0);
nand U1131 (N_1131,N_109,N_192);
and U1132 (N_1132,N_72,N_497);
and U1133 (N_1133,N_606,N_249);
nor U1134 (N_1134,N_697,N_185);
or U1135 (N_1135,N_505,N_85);
and U1136 (N_1136,N_658,N_550);
or U1137 (N_1137,N_309,N_111);
nand U1138 (N_1138,N_524,N_243);
and U1139 (N_1139,N_260,N_571);
nand U1140 (N_1140,N_266,N_248);
or U1141 (N_1141,N_199,N_735);
nor U1142 (N_1142,N_193,N_467);
or U1143 (N_1143,N_283,N_721);
or U1144 (N_1144,N_160,N_545);
and U1145 (N_1145,N_620,N_172);
nand U1146 (N_1146,N_479,N_157);
nand U1147 (N_1147,N_629,N_287);
or U1148 (N_1148,N_296,N_255);
nand U1149 (N_1149,N_579,N_741);
nand U1150 (N_1150,N_179,N_682);
or U1151 (N_1151,N_236,N_601);
nor U1152 (N_1152,N_628,N_646);
nor U1153 (N_1153,N_54,N_322);
or U1154 (N_1154,N_28,N_649);
nand U1155 (N_1155,N_388,N_517);
or U1156 (N_1156,N_713,N_668);
and U1157 (N_1157,N_360,N_666);
or U1158 (N_1158,N_113,N_291);
and U1159 (N_1159,N_725,N_400);
nor U1160 (N_1160,N_546,N_122);
nand U1161 (N_1161,N_318,N_32);
and U1162 (N_1162,N_424,N_608);
nand U1163 (N_1163,N_95,N_527);
nand U1164 (N_1164,N_304,N_381);
nor U1165 (N_1165,N_691,N_620);
or U1166 (N_1166,N_356,N_341);
and U1167 (N_1167,N_689,N_381);
and U1168 (N_1168,N_236,N_424);
or U1169 (N_1169,N_208,N_682);
or U1170 (N_1170,N_85,N_54);
or U1171 (N_1171,N_512,N_446);
or U1172 (N_1172,N_98,N_291);
nand U1173 (N_1173,N_150,N_444);
nand U1174 (N_1174,N_492,N_441);
or U1175 (N_1175,N_40,N_737);
and U1176 (N_1176,N_342,N_57);
nor U1177 (N_1177,N_174,N_555);
and U1178 (N_1178,N_108,N_201);
nand U1179 (N_1179,N_240,N_107);
nand U1180 (N_1180,N_582,N_362);
or U1181 (N_1181,N_75,N_50);
nand U1182 (N_1182,N_558,N_442);
and U1183 (N_1183,N_436,N_270);
nand U1184 (N_1184,N_225,N_699);
nor U1185 (N_1185,N_568,N_595);
nand U1186 (N_1186,N_77,N_13);
xor U1187 (N_1187,N_192,N_290);
nor U1188 (N_1188,N_701,N_105);
nor U1189 (N_1189,N_44,N_335);
nor U1190 (N_1190,N_496,N_392);
or U1191 (N_1191,N_92,N_95);
and U1192 (N_1192,N_319,N_184);
or U1193 (N_1193,N_215,N_303);
and U1194 (N_1194,N_68,N_408);
and U1195 (N_1195,N_439,N_73);
or U1196 (N_1196,N_235,N_131);
nand U1197 (N_1197,N_727,N_524);
and U1198 (N_1198,N_167,N_22);
nand U1199 (N_1199,N_636,N_54);
or U1200 (N_1200,N_386,N_220);
and U1201 (N_1201,N_51,N_514);
nand U1202 (N_1202,N_80,N_632);
or U1203 (N_1203,N_644,N_103);
and U1204 (N_1204,N_207,N_314);
or U1205 (N_1205,N_180,N_108);
xnor U1206 (N_1206,N_418,N_561);
nor U1207 (N_1207,N_473,N_62);
or U1208 (N_1208,N_676,N_639);
nand U1209 (N_1209,N_376,N_19);
and U1210 (N_1210,N_207,N_686);
nand U1211 (N_1211,N_425,N_107);
nand U1212 (N_1212,N_560,N_410);
and U1213 (N_1213,N_650,N_460);
nor U1214 (N_1214,N_735,N_207);
nor U1215 (N_1215,N_210,N_351);
nand U1216 (N_1216,N_106,N_451);
or U1217 (N_1217,N_141,N_683);
nor U1218 (N_1218,N_90,N_614);
or U1219 (N_1219,N_555,N_240);
and U1220 (N_1220,N_428,N_465);
or U1221 (N_1221,N_499,N_653);
or U1222 (N_1222,N_629,N_9);
nor U1223 (N_1223,N_319,N_282);
and U1224 (N_1224,N_626,N_310);
or U1225 (N_1225,N_550,N_352);
nor U1226 (N_1226,N_378,N_160);
and U1227 (N_1227,N_652,N_450);
nor U1228 (N_1228,N_421,N_707);
nand U1229 (N_1229,N_737,N_742);
nand U1230 (N_1230,N_316,N_443);
nand U1231 (N_1231,N_153,N_38);
nor U1232 (N_1232,N_616,N_313);
or U1233 (N_1233,N_577,N_504);
or U1234 (N_1234,N_304,N_517);
nand U1235 (N_1235,N_253,N_472);
and U1236 (N_1236,N_529,N_118);
or U1237 (N_1237,N_46,N_445);
or U1238 (N_1238,N_662,N_596);
and U1239 (N_1239,N_158,N_423);
and U1240 (N_1240,N_138,N_722);
or U1241 (N_1241,N_509,N_328);
nor U1242 (N_1242,N_18,N_327);
or U1243 (N_1243,N_738,N_739);
or U1244 (N_1244,N_514,N_677);
or U1245 (N_1245,N_255,N_295);
and U1246 (N_1246,N_694,N_647);
and U1247 (N_1247,N_317,N_174);
and U1248 (N_1248,N_684,N_152);
or U1249 (N_1249,N_51,N_15);
or U1250 (N_1250,N_6,N_277);
or U1251 (N_1251,N_105,N_351);
or U1252 (N_1252,N_619,N_584);
nand U1253 (N_1253,N_76,N_95);
or U1254 (N_1254,N_521,N_13);
and U1255 (N_1255,N_112,N_216);
and U1256 (N_1256,N_581,N_441);
nand U1257 (N_1257,N_186,N_116);
and U1258 (N_1258,N_63,N_661);
and U1259 (N_1259,N_420,N_652);
nor U1260 (N_1260,N_355,N_373);
or U1261 (N_1261,N_307,N_699);
or U1262 (N_1262,N_235,N_8);
nor U1263 (N_1263,N_504,N_314);
xnor U1264 (N_1264,N_615,N_165);
nor U1265 (N_1265,N_631,N_563);
nor U1266 (N_1266,N_683,N_450);
nor U1267 (N_1267,N_523,N_599);
nor U1268 (N_1268,N_236,N_651);
and U1269 (N_1269,N_433,N_86);
or U1270 (N_1270,N_551,N_576);
nor U1271 (N_1271,N_287,N_628);
nor U1272 (N_1272,N_696,N_207);
nand U1273 (N_1273,N_614,N_234);
or U1274 (N_1274,N_659,N_97);
nand U1275 (N_1275,N_261,N_497);
nor U1276 (N_1276,N_386,N_705);
nor U1277 (N_1277,N_294,N_268);
or U1278 (N_1278,N_666,N_493);
or U1279 (N_1279,N_546,N_148);
nor U1280 (N_1280,N_403,N_12);
nor U1281 (N_1281,N_643,N_731);
nand U1282 (N_1282,N_260,N_589);
and U1283 (N_1283,N_441,N_734);
nor U1284 (N_1284,N_285,N_114);
and U1285 (N_1285,N_657,N_556);
nand U1286 (N_1286,N_702,N_205);
and U1287 (N_1287,N_63,N_568);
xnor U1288 (N_1288,N_557,N_297);
and U1289 (N_1289,N_258,N_542);
and U1290 (N_1290,N_282,N_12);
nand U1291 (N_1291,N_281,N_145);
or U1292 (N_1292,N_504,N_246);
or U1293 (N_1293,N_385,N_741);
nand U1294 (N_1294,N_482,N_748);
or U1295 (N_1295,N_648,N_510);
or U1296 (N_1296,N_212,N_159);
nand U1297 (N_1297,N_131,N_475);
nor U1298 (N_1298,N_689,N_286);
and U1299 (N_1299,N_117,N_493);
and U1300 (N_1300,N_727,N_448);
or U1301 (N_1301,N_174,N_28);
or U1302 (N_1302,N_182,N_40);
nor U1303 (N_1303,N_608,N_93);
nand U1304 (N_1304,N_203,N_679);
nor U1305 (N_1305,N_483,N_435);
nor U1306 (N_1306,N_738,N_203);
nand U1307 (N_1307,N_298,N_118);
and U1308 (N_1308,N_147,N_63);
nor U1309 (N_1309,N_720,N_259);
nand U1310 (N_1310,N_284,N_599);
and U1311 (N_1311,N_150,N_182);
nand U1312 (N_1312,N_176,N_649);
and U1313 (N_1313,N_70,N_669);
nor U1314 (N_1314,N_85,N_2);
nor U1315 (N_1315,N_539,N_463);
and U1316 (N_1316,N_286,N_192);
or U1317 (N_1317,N_11,N_80);
nor U1318 (N_1318,N_492,N_708);
or U1319 (N_1319,N_83,N_273);
or U1320 (N_1320,N_204,N_161);
nand U1321 (N_1321,N_420,N_493);
and U1322 (N_1322,N_286,N_295);
nand U1323 (N_1323,N_367,N_289);
or U1324 (N_1324,N_649,N_31);
nor U1325 (N_1325,N_435,N_129);
and U1326 (N_1326,N_92,N_337);
and U1327 (N_1327,N_472,N_124);
nor U1328 (N_1328,N_475,N_673);
and U1329 (N_1329,N_479,N_349);
nor U1330 (N_1330,N_746,N_377);
nor U1331 (N_1331,N_431,N_334);
nor U1332 (N_1332,N_721,N_107);
and U1333 (N_1333,N_606,N_67);
or U1334 (N_1334,N_366,N_103);
nand U1335 (N_1335,N_680,N_633);
or U1336 (N_1336,N_182,N_149);
and U1337 (N_1337,N_87,N_188);
and U1338 (N_1338,N_645,N_295);
and U1339 (N_1339,N_201,N_34);
or U1340 (N_1340,N_341,N_679);
nor U1341 (N_1341,N_340,N_441);
nand U1342 (N_1342,N_713,N_344);
or U1343 (N_1343,N_357,N_445);
and U1344 (N_1344,N_692,N_72);
or U1345 (N_1345,N_209,N_421);
nor U1346 (N_1346,N_338,N_14);
nor U1347 (N_1347,N_380,N_81);
or U1348 (N_1348,N_456,N_134);
and U1349 (N_1349,N_96,N_747);
nand U1350 (N_1350,N_81,N_603);
or U1351 (N_1351,N_310,N_494);
and U1352 (N_1352,N_121,N_532);
nor U1353 (N_1353,N_578,N_303);
and U1354 (N_1354,N_303,N_235);
or U1355 (N_1355,N_266,N_183);
or U1356 (N_1356,N_230,N_545);
and U1357 (N_1357,N_112,N_44);
nand U1358 (N_1358,N_465,N_739);
or U1359 (N_1359,N_83,N_132);
and U1360 (N_1360,N_84,N_748);
nand U1361 (N_1361,N_554,N_4);
or U1362 (N_1362,N_37,N_110);
or U1363 (N_1363,N_29,N_403);
nor U1364 (N_1364,N_282,N_250);
and U1365 (N_1365,N_666,N_59);
nor U1366 (N_1366,N_28,N_636);
nor U1367 (N_1367,N_404,N_22);
and U1368 (N_1368,N_63,N_261);
nand U1369 (N_1369,N_633,N_151);
nand U1370 (N_1370,N_486,N_65);
and U1371 (N_1371,N_283,N_682);
nor U1372 (N_1372,N_579,N_716);
nand U1373 (N_1373,N_159,N_104);
nand U1374 (N_1374,N_287,N_314);
nor U1375 (N_1375,N_476,N_287);
and U1376 (N_1376,N_215,N_163);
or U1377 (N_1377,N_638,N_159);
or U1378 (N_1378,N_587,N_397);
nand U1379 (N_1379,N_311,N_517);
nand U1380 (N_1380,N_721,N_397);
and U1381 (N_1381,N_552,N_688);
and U1382 (N_1382,N_599,N_173);
or U1383 (N_1383,N_560,N_199);
nor U1384 (N_1384,N_400,N_660);
nor U1385 (N_1385,N_628,N_501);
or U1386 (N_1386,N_532,N_232);
nor U1387 (N_1387,N_28,N_100);
nand U1388 (N_1388,N_569,N_469);
nand U1389 (N_1389,N_171,N_424);
nor U1390 (N_1390,N_536,N_382);
nor U1391 (N_1391,N_94,N_677);
and U1392 (N_1392,N_305,N_58);
nor U1393 (N_1393,N_37,N_439);
or U1394 (N_1394,N_139,N_274);
nor U1395 (N_1395,N_336,N_315);
or U1396 (N_1396,N_345,N_584);
nor U1397 (N_1397,N_37,N_521);
or U1398 (N_1398,N_406,N_439);
or U1399 (N_1399,N_478,N_533);
or U1400 (N_1400,N_274,N_401);
or U1401 (N_1401,N_183,N_734);
xnor U1402 (N_1402,N_242,N_717);
xor U1403 (N_1403,N_611,N_616);
nand U1404 (N_1404,N_645,N_560);
nor U1405 (N_1405,N_601,N_79);
or U1406 (N_1406,N_280,N_660);
nand U1407 (N_1407,N_739,N_512);
or U1408 (N_1408,N_449,N_203);
or U1409 (N_1409,N_337,N_720);
nand U1410 (N_1410,N_326,N_406);
and U1411 (N_1411,N_705,N_353);
and U1412 (N_1412,N_300,N_514);
nor U1413 (N_1413,N_613,N_265);
nor U1414 (N_1414,N_37,N_675);
nor U1415 (N_1415,N_377,N_292);
nand U1416 (N_1416,N_363,N_656);
nand U1417 (N_1417,N_651,N_229);
nand U1418 (N_1418,N_606,N_178);
nor U1419 (N_1419,N_733,N_666);
or U1420 (N_1420,N_707,N_505);
nor U1421 (N_1421,N_627,N_591);
nand U1422 (N_1422,N_362,N_52);
and U1423 (N_1423,N_28,N_348);
and U1424 (N_1424,N_21,N_282);
nand U1425 (N_1425,N_433,N_558);
nor U1426 (N_1426,N_673,N_222);
or U1427 (N_1427,N_356,N_672);
nor U1428 (N_1428,N_578,N_458);
and U1429 (N_1429,N_104,N_398);
nand U1430 (N_1430,N_226,N_111);
nor U1431 (N_1431,N_712,N_741);
or U1432 (N_1432,N_279,N_694);
nand U1433 (N_1433,N_658,N_249);
nor U1434 (N_1434,N_613,N_479);
nor U1435 (N_1435,N_134,N_216);
or U1436 (N_1436,N_712,N_261);
or U1437 (N_1437,N_398,N_127);
or U1438 (N_1438,N_26,N_537);
and U1439 (N_1439,N_203,N_126);
and U1440 (N_1440,N_516,N_124);
or U1441 (N_1441,N_524,N_707);
and U1442 (N_1442,N_209,N_355);
nor U1443 (N_1443,N_477,N_624);
and U1444 (N_1444,N_516,N_74);
or U1445 (N_1445,N_249,N_165);
or U1446 (N_1446,N_503,N_77);
and U1447 (N_1447,N_393,N_458);
nand U1448 (N_1448,N_701,N_689);
and U1449 (N_1449,N_267,N_595);
and U1450 (N_1450,N_287,N_326);
and U1451 (N_1451,N_223,N_642);
nor U1452 (N_1452,N_510,N_158);
and U1453 (N_1453,N_209,N_9);
nand U1454 (N_1454,N_220,N_675);
and U1455 (N_1455,N_132,N_554);
or U1456 (N_1456,N_616,N_326);
and U1457 (N_1457,N_540,N_117);
nor U1458 (N_1458,N_391,N_436);
or U1459 (N_1459,N_484,N_289);
or U1460 (N_1460,N_1,N_20);
or U1461 (N_1461,N_328,N_601);
nor U1462 (N_1462,N_196,N_675);
nand U1463 (N_1463,N_328,N_130);
nor U1464 (N_1464,N_518,N_689);
and U1465 (N_1465,N_289,N_175);
and U1466 (N_1466,N_445,N_590);
and U1467 (N_1467,N_520,N_114);
nand U1468 (N_1468,N_475,N_41);
and U1469 (N_1469,N_553,N_489);
or U1470 (N_1470,N_722,N_422);
nand U1471 (N_1471,N_64,N_489);
nand U1472 (N_1472,N_704,N_76);
nand U1473 (N_1473,N_749,N_539);
or U1474 (N_1474,N_609,N_183);
and U1475 (N_1475,N_598,N_272);
or U1476 (N_1476,N_147,N_567);
nor U1477 (N_1477,N_56,N_20);
and U1478 (N_1478,N_438,N_103);
and U1479 (N_1479,N_435,N_136);
and U1480 (N_1480,N_683,N_21);
xnor U1481 (N_1481,N_536,N_94);
or U1482 (N_1482,N_77,N_477);
or U1483 (N_1483,N_541,N_682);
nand U1484 (N_1484,N_559,N_656);
nand U1485 (N_1485,N_619,N_193);
nand U1486 (N_1486,N_666,N_90);
or U1487 (N_1487,N_397,N_633);
nor U1488 (N_1488,N_569,N_136);
and U1489 (N_1489,N_615,N_614);
xor U1490 (N_1490,N_133,N_482);
or U1491 (N_1491,N_86,N_341);
xor U1492 (N_1492,N_739,N_378);
nand U1493 (N_1493,N_493,N_86);
nand U1494 (N_1494,N_278,N_65);
xor U1495 (N_1495,N_477,N_625);
or U1496 (N_1496,N_81,N_341);
nor U1497 (N_1497,N_255,N_337);
or U1498 (N_1498,N_368,N_61);
nor U1499 (N_1499,N_284,N_203);
nor U1500 (N_1500,N_1423,N_844);
and U1501 (N_1501,N_923,N_850);
or U1502 (N_1502,N_1041,N_1203);
and U1503 (N_1503,N_1285,N_1164);
nor U1504 (N_1504,N_1351,N_901);
or U1505 (N_1505,N_1079,N_1362);
or U1506 (N_1506,N_1361,N_1274);
or U1507 (N_1507,N_1412,N_1102);
nand U1508 (N_1508,N_898,N_1488);
nand U1509 (N_1509,N_1359,N_945);
or U1510 (N_1510,N_940,N_1230);
nand U1511 (N_1511,N_1004,N_820);
nand U1512 (N_1512,N_1306,N_1127);
nor U1513 (N_1513,N_978,N_1204);
nor U1514 (N_1514,N_1290,N_1471);
nand U1515 (N_1515,N_963,N_888);
or U1516 (N_1516,N_902,N_1410);
and U1517 (N_1517,N_750,N_1128);
or U1518 (N_1518,N_753,N_1416);
or U1519 (N_1519,N_1263,N_860);
and U1520 (N_1520,N_1266,N_1155);
nand U1521 (N_1521,N_1427,N_979);
or U1522 (N_1522,N_1140,N_1473);
and U1523 (N_1523,N_786,N_755);
nand U1524 (N_1524,N_1382,N_774);
and U1525 (N_1525,N_976,N_1460);
nand U1526 (N_1526,N_1019,N_843);
and U1527 (N_1527,N_1322,N_920);
nand U1528 (N_1528,N_1420,N_1367);
and U1529 (N_1529,N_1307,N_832);
nand U1530 (N_1530,N_1134,N_1355);
and U1531 (N_1531,N_1078,N_758);
and U1532 (N_1532,N_1052,N_1441);
nor U1533 (N_1533,N_1113,N_1388);
and U1534 (N_1534,N_1235,N_1180);
and U1535 (N_1535,N_830,N_810);
nor U1536 (N_1536,N_964,N_1209);
or U1537 (N_1537,N_1479,N_1207);
nand U1538 (N_1538,N_1324,N_1063);
and U1539 (N_1539,N_781,N_1446);
nand U1540 (N_1540,N_854,N_1286);
or U1541 (N_1541,N_837,N_1492);
nor U1542 (N_1542,N_1454,N_1484);
or U1543 (N_1543,N_1316,N_1470);
xnor U1544 (N_1544,N_891,N_1458);
and U1545 (N_1545,N_927,N_1438);
nor U1546 (N_1546,N_947,N_1269);
nand U1547 (N_1547,N_1039,N_1025);
or U1548 (N_1548,N_1330,N_804);
nor U1549 (N_1549,N_1040,N_1291);
nand U1550 (N_1550,N_1225,N_1348);
nand U1551 (N_1551,N_790,N_1186);
nand U1552 (N_1552,N_909,N_809);
and U1553 (N_1553,N_1369,N_912);
nor U1554 (N_1554,N_879,N_778);
nor U1555 (N_1555,N_1073,N_1212);
or U1556 (N_1556,N_1157,N_1168);
or U1557 (N_1557,N_1270,N_1008);
nor U1558 (N_1558,N_1233,N_1001);
nor U1559 (N_1559,N_1401,N_1035);
nand U1560 (N_1560,N_1183,N_1424);
and U1561 (N_1561,N_1024,N_896);
and U1562 (N_1562,N_1245,N_1447);
nand U1563 (N_1563,N_1434,N_1363);
nor U1564 (N_1564,N_1053,N_868);
xnor U1565 (N_1565,N_1229,N_1453);
nor U1566 (N_1566,N_1328,N_1469);
and U1567 (N_1567,N_1103,N_1169);
or U1568 (N_1568,N_763,N_1301);
nor U1569 (N_1569,N_1390,N_766);
nor U1570 (N_1570,N_1399,N_792);
or U1571 (N_1571,N_1220,N_931);
and U1572 (N_1572,N_872,N_1248);
nand U1573 (N_1573,N_1122,N_1069);
and U1574 (N_1574,N_1459,N_1387);
and U1575 (N_1575,N_962,N_1413);
and U1576 (N_1576,N_1028,N_886);
and U1577 (N_1577,N_1014,N_1202);
and U1578 (N_1578,N_798,N_870);
and U1579 (N_1579,N_1214,N_955);
or U1580 (N_1580,N_1156,N_1298);
nand U1581 (N_1581,N_1100,N_1349);
nand U1582 (N_1582,N_1077,N_1497);
nand U1583 (N_1583,N_806,N_1027);
nor U1584 (N_1584,N_1241,N_797);
and U1585 (N_1585,N_1105,N_1275);
nand U1586 (N_1586,N_1036,N_1368);
and U1587 (N_1587,N_859,N_1189);
nand U1588 (N_1588,N_796,N_1007);
nand U1589 (N_1589,N_1231,N_835);
nor U1590 (N_1590,N_1430,N_1256);
xnor U1591 (N_1591,N_1477,N_1147);
nand U1592 (N_1592,N_1417,N_1345);
nor U1593 (N_1593,N_1236,N_1440);
nor U1594 (N_1594,N_895,N_1483);
or U1595 (N_1595,N_1129,N_760);
and U1596 (N_1596,N_1120,N_1197);
and U1597 (N_1597,N_1192,N_954);
nand U1598 (N_1598,N_1058,N_1003);
nand U1599 (N_1599,N_1398,N_929);
nor U1600 (N_1600,N_861,N_817);
and U1601 (N_1601,N_1373,N_941);
nor U1602 (N_1602,N_1211,N_1247);
nand U1603 (N_1603,N_1261,N_768);
nor U1604 (N_1604,N_932,N_1386);
nand U1605 (N_1605,N_939,N_918);
nor U1606 (N_1606,N_1449,N_1026);
nor U1607 (N_1607,N_1185,N_1087);
and U1608 (N_1608,N_974,N_1032);
nor U1609 (N_1609,N_771,N_1259);
nand U1610 (N_1610,N_1119,N_1173);
nand U1611 (N_1611,N_1246,N_1135);
and U1612 (N_1612,N_823,N_910);
or U1613 (N_1613,N_814,N_1486);
nand U1614 (N_1614,N_769,N_958);
nor U1615 (N_1615,N_1402,N_1415);
or U1616 (N_1616,N_871,N_1054);
nor U1617 (N_1617,N_1067,N_1457);
and U1618 (N_1618,N_1293,N_1494);
or U1619 (N_1619,N_1234,N_887);
nand U1620 (N_1620,N_1406,N_1123);
nor U1621 (N_1621,N_1048,N_1037);
and U1622 (N_1622,N_1170,N_876);
and U1623 (N_1623,N_928,N_1315);
xnor U1624 (N_1624,N_1276,N_1217);
nor U1625 (N_1625,N_1252,N_972);
and U1626 (N_1626,N_1174,N_1057);
and U1627 (N_1627,N_890,N_803);
nor U1628 (N_1628,N_1182,N_1300);
nor U1629 (N_1629,N_1319,N_825);
or U1630 (N_1630,N_1418,N_759);
and U1631 (N_1631,N_1033,N_1378);
or U1632 (N_1632,N_1422,N_1093);
xor U1633 (N_1633,N_1110,N_1193);
or U1634 (N_1634,N_829,N_867);
nand U1635 (N_1635,N_1085,N_1370);
nand U1636 (N_1636,N_1358,N_1137);
and U1637 (N_1637,N_1126,N_752);
or U1638 (N_1638,N_1200,N_767);
or U1639 (N_1639,N_1074,N_943);
and U1640 (N_1640,N_1199,N_987);
or U1641 (N_1641,N_805,N_1222);
nand U1642 (N_1642,N_1313,N_1442);
nand U1643 (N_1643,N_1435,N_1336);
nor U1644 (N_1644,N_1018,N_761);
nand U1645 (N_1645,N_1227,N_921);
or U1646 (N_1646,N_1012,N_926);
nand U1647 (N_1647,N_1172,N_1331);
and U1648 (N_1648,N_1021,N_1264);
nand U1649 (N_1649,N_840,N_1436);
nor U1650 (N_1650,N_773,N_828);
nor U1651 (N_1651,N_776,N_1303);
nor U1652 (N_1652,N_907,N_1339);
xor U1653 (N_1653,N_1108,N_1318);
nand U1654 (N_1654,N_1124,N_1044);
and U1655 (N_1655,N_1090,N_851);
and U1656 (N_1656,N_1254,N_1010);
or U1657 (N_1657,N_757,N_952);
nor U1658 (N_1658,N_908,N_1094);
or U1659 (N_1659,N_1342,N_1095);
and U1660 (N_1660,N_1480,N_869);
nor U1661 (N_1661,N_1112,N_1350);
nor U1662 (N_1662,N_933,N_1092);
and U1663 (N_1663,N_1042,N_1242);
or U1664 (N_1664,N_1190,N_1304);
and U1665 (N_1665,N_1467,N_1224);
nand U1666 (N_1666,N_973,N_970);
or U1667 (N_1667,N_1179,N_904);
nand U1668 (N_1668,N_756,N_1237);
or U1669 (N_1669,N_1076,N_1294);
nand U1670 (N_1670,N_802,N_1114);
or U1671 (N_1671,N_930,N_1226);
or U1672 (N_1672,N_1392,N_813);
nor U1673 (N_1673,N_1020,N_1064);
nor U1674 (N_1674,N_1148,N_905);
or U1675 (N_1675,N_1221,N_981);
nand U1676 (N_1676,N_866,N_1496);
nor U1677 (N_1677,N_882,N_1238);
nor U1678 (N_1678,N_807,N_1419);
or U1679 (N_1679,N_983,N_1279);
and U1680 (N_1680,N_922,N_925);
nor U1681 (N_1681,N_1409,N_1243);
and U1682 (N_1682,N_784,N_1111);
nor U1683 (N_1683,N_1393,N_1049);
or U1684 (N_1684,N_1091,N_821);
or U1685 (N_1685,N_1191,N_849);
and U1686 (N_1686,N_1347,N_1070);
and U1687 (N_1687,N_1136,N_960);
nor U1688 (N_1688,N_885,N_1353);
nand U1689 (N_1689,N_1059,N_999);
nor U1690 (N_1690,N_765,N_1320);
nand U1691 (N_1691,N_965,N_1489);
and U1692 (N_1692,N_1109,N_1375);
xnor U1693 (N_1693,N_1311,N_1096);
and U1694 (N_1694,N_975,N_1312);
nand U1695 (N_1695,N_864,N_1030);
or U1696 (N_1696,N_1163,N_1280);
and U1697 (N_1697,N_1196,N_889);
and U1698 (N_1698,N_1405,N_878);
and U1699 (N_1699,N_1142,N_1240);
or U1700 (N_1700,N_1364,N_906);
nand U1701 (N_1701,N_754,N_1407);
or U1702 (N_1702,N_841,N_1194);
nand U1703 (N_1703,N_1031,N_1062);
and U1704 (N_1704,N_1232,N_1421);
or U1705 (N_1705,N_811,N_996);
nand U1706 (N_1706,N_1490,N_1374);
and U1707 (N_1707,N_1425,N_1481);
nand U1708 (N_1708,N_998,N_1433);
or U1709 (N_1709,N_1167,N_1250);
or U1710 (N_1710,N_858,N_919);
and U1711 (N_1711,N_957,N_1450);
or U1712 (N_1712,N_1152,N_995);
or U1713 (N_1713,N_961,N_788);
nand U1714 (N_1714,N_1084,N_897);
or U1715 (N_1715,N_1268,N_1376);
or U1716 (N_1716,N_1205,N_934);
nor U1717 (N_1717,N_799,N_1029);
xor U1718 (N_1718,N_990,N_984);
and U1719 (N_1719,N_1060,N_1139);
or U1720 (N_1720,N_831,N_948);
nor U1721 (N_1721,N_779,N_953);
nand U1722 (N_1722,N_1287,N_1255);
or U1723 (N_1723,N_1452,N_1097);
and U1724 (N_1724,N_1144,N_827);
or U1725 (N_1725,N_772,N_847);
or U1726 (N_1726,N_1299,N_1456);
nor U1727 (N_1727,N_1160,N_1385);
nor U1728 (N_1728,N_1153,N_1166);
xor U1729 (N_1729,N_1218,N_1176);
nand U1730 (N_1730,N_1198,N_994);
nand U1731 (N_1731,N_1408,N_783);
nor U1732 (N_1732,N_1493,N_1475);
nand U1733 (N_1733,N_856,N_865);
and U1734 (N_1734,N_775,N_1448);
nand U1735 (N_1735,N_936,N_764);
nor U1736 (N_1736,N_1465,N_1283);
or U1737 (N_1737,N_992,N_1377);
and U1738 (N_1738,N_1338,N_1371);
nand U1739 (N_1739,N_1379,N_1472);
nand U1740 (N_1740,N_852,N_1143);
nor U1741 (N_1741,N_1265,N_1317);
or U1742 (N_1742,N_794,N_1133);
or U1743 (N_1743,N_1065,N_1171);
nand U1744 (N_1744,N_1432,N_1107);
or U1745 (N_1745,N_1281,N_1391);
or U1746 (N_1746,N_1272,N_1006);
nand U1747 (N_1747,N_1015,N_993);
nor U1748 (N_1748,N_1081,N_980);
nand U1749 (N_1749,N_977,N_1201);
and U1750 (N_1750,N_1016,N_1034);
or U1751 (N_1751,N_795,N_1075);
nand U1752 (N_1752,N_845,N_1474);
nand U1753 (N_1753,N_1098,N_1414);
nand U1754 (N_1754,N_1083,N_875);
nor U1755 (N_1755,N_1253,N_848);
and U1756 (N_1756,N_1005,N_1162);
and U1757 (N_1757,N_836,N_1175);
or U1758 (N_1758,N_880,N_1045);
and U1759 (N_1759,N_1444,N_1333);
or U1760 (N_1760,N_971,N_935);
nor U1761 (N_1761,N_881,N_1086);
nand U1762 (N_1762,N_1213,N_1013);
nor U1763 (N_1763,N_942,N_1258);
nand U1764 (N_1764,N_863,N_1101);
nor U1765 (N_1765,N_812,N_1149);
or U1766 (N_1766,N_877,N_1485);
nand U1767 (N_1767,N_1384,N_1437);
nand U1768 (N_1768,N_1321,N_1323);
nand U1769 (N_1769,N_853,N_1462);
nor U1770 (N_1770,N_1389,N_1468);
nand U1771 (N_1771,N_893,N_1099);
nor U1772 (N_1772,N_1177,N_1022);
or U1773 (N_1773,N_892,N_988);
nand U1774 (N_1774,N_751,N_1106);
nand U1775 (N_1775,N_1121,N_1343);
or U1776 (N_1776,N_1002,N_1260);
or U1777 (N_1777,N_1403,N_900);
or U1778 (N_1778,N_1145,N_1158);
nand U1779 (N_1779,N_1188,N_1118);
or U1780 (N_1780,N_1154,N_1340);
and U1781 (N_1781,N_1335,N_1326);
nand U1782 (N_1782,N_857,N_1404);
nand U1783 (N_1783,N_1043,N_1310);
nor U1784 (N_1784,N_1284,N_1066);
and U1785 (N_1785,N_1206,N_1038);
xor U1786 (N_1786,N_1394,N_1208);
nor U1787 (N_1787,N_873,N_969);
and U1788 (N_1788,N_913,N_1381);
nor U1789 (N_1789,N_924,N_789);
or U1790 (N_1790,N_1068,N_1277);
nand U1791 (N_1791,N_1327,N_1146);
nor U1792 (N_1792,N_1451,N_915);
and U1793 (N_1793,N_1165,N_1159);
nor U1794 (N_1794,N_1332,N_966);
nor U1795 (N_1795,N_834,N_1396);
or U1796 (N_1796,N_989,N_1082);
nand U1797 (N_1797,N_1297,N_1428);
or U1798 (N_1798,N_956,N_1249);
nand U1799 (N_1799,N_1228,N_1138);
or U1800 (N_1800,N_959,N_800);
or U1801 (N_1801,N_1499,N_1061);
nand U1802 (N_1802,N_1443,N_1491);
or U1803 (N_1803,N_982,N_985);
and U1804 (N_1804,N_1050,N_826);
nor U1805 (N_1805,N_1397,N_1150);
nor U1806 (N_1806,N_1047,N_1071);
nor U1807 (N_1807,N_1115,N_1278);
and U1808 (N_1808,N_808,N_1365);
and U1809 (N_1809,N_1354,N_862);
or U1810 (N_1810,N_1017,N_1411);
nor U1811 (N_1811,N_1051,N_1178);
and U1812 (N_1812,N_1439,N_1325);
nand U1813 (N_1813,N_1210,N_1055);
or U1814 (N_1814,N_1341,N_1187);
nor U1815 (N_1815,N_1466,N_1271);
nor U1816 (N_1816,N_1289,N_1292);
and U1817 (N_1817,N_946,N_1251);
and U1818 (N_1818,N_1498,N_1244);
nor U1819 (N_1819,N_1476,N_815);
nand U1820 (N_1820,N_1445,N_1056);
and U1821 (N_1821,N_1195,N_950);
and U1822 (N_1822,N_917,N_1366);
nor U1823 (N_1823,N_1495,N_838);
or U1824 (N_1824,N_1295,N_819);
and U1825 (N_1825,N_1239,N_1011);
and U1826 (N_1826,N_855,N_1357);
or U1827 (N_1827,N_1463,N_1181);
nand U1828 (N_1828,N_997,N_1273);
and U1829 (N_1829,N_818,N_822);
or U1830 (N_1830,N_1072,N_903);
and U1831 (N_1831,N_1132,N_787);
nor U1832 (N_1832,N_824,N_1464);
nor U1833 (N_1833,N_1426,N_1482);
nand U1834 (N_1834,N_968,N_1296);
and U1835 (N_1835,N_1352,N_967);
nor U1836 (N_1836,N_1334,N_833);
nor U1837 (N_1837,N_1308,N_1125);
nand U1838 (N_1838,N_1461,N_1429);
or U1839 (N_1839,N_916,N_991);
nor U1840 (N_1840,N_801,N_1288);
nor U1841 (N_1841,N_938,N_1257);
nor U1842 (N_1842,N_1223,N_780);
and U1843 (N_1843,N_1395,N_1329);
xor U1844 (N_1844,N_937,N_1360);
xor U1845 (N_1845,N_1455,N_1262);
nor U1846 (N_1846,N_874,N_1089);
nand U1847 (N_1847,N_785,N_1023);
nand U1848 (N_1848,N_1104,N_1383);
or U1849 (N_1849,N_1356,N_1305);
and U1850 (N_1850,N_1009,N_1219);
or U1851 (N_1851,N_899,N_1215);
and U1852 (N_1852,N_883,N_1372);
nand U1853 (N_1853,N_951,N_1478);
nand U1854 (N_1854,N_1141,N_816);
nand U1855 (N_1855,N_914,N_1117);
nor U1856 (N_1856,N_1314,N_1000);
nor U1857 (N_1857,N_1487,N_1130);
or U1858 (N_1858,N_894,N_1380);
and U1859 (N_1859,N_1184,N_1116);
or U1860 (N_1860,N_1344,N_782);
nor U1861 (N_1861,N_793,N_846);
and U1862 (N_1862,N_1267,N_949);
nand U1863 (N_1863,N_884,N_770);
nor U1864 (N_1864,N_1088,N_1431);
xnor U1865 (N_1865,N_839,N_1131);
or U1866 (N_1866,N_842,N_1400);
nand U1867 (N_1867,N_791,N_1337);
or U1868 (N_1868,N_1151,N_1216);
and U1869 (N_1869,N_762,N_777);
and U1870 (N_1870,N_1282,N_944);
nand U1871 (N_1871,N_1309,N_1046);
or U1872 (N_1872,N_1302,N_1161);
and U1873 (N_1873,N_911,N_1080);
and U1874 (N_1874,N_1346,N_986);
nor U1875 (N_1875,N_790,N_796);
and U1876 (N_1876,N_1299,N_948);
or U1877 (N_1877,N_1074,N_1159);
nand U1878 (N_1878,N_977,N_1159);
and U1879 (N_1879,N_864,N_1112);
nand U1880 (N_1880,N_994,N_834);
and U1881 (N_1881,N_1055,N_1125);
nor U1882 (N_1882,N_1336,N_1134);
xnor U1883 (N_1883,N_1177,N_1106);
nand U1884 (N_1884,N_1377,N_954);
nor U1885 (N_1885,N_1169,N_1305);
nand U1886 (N_1886,N_1050,N_1373);
or U1887 (N_1887,N_865,N_1210);
and U1888 (N_1888,N_1130,N_902);
nor U1889 (N_1889,N_1126,N_1112);
nor U1890 (N_1890,N_994,N_1415);
nand U1891 (N_1891,N_1143,N_831);
nor U1892 (N_1892,N_1242,N_990);
nor U1893 (N_1893,N_894,N_1068);
or U1894 (N_1894,N_1055,N_1349);
and U1895 (N_1895,N_1479,N_1180);
nand U1896 (N_1896,N_1006,N_1339);
xnor U1897 (N_1897,N_1403,N_1489);
nor U1898 (N_1898,N_1414,N_1121);
and U1899 (N_1899,N_861,N_1283);
nor U1900 (N_1900,N_1222,N_1258);
or U1901 (N_1901,N_1084,N_1149);
and U1902 (N_1902,N_1182,N_1079);
or U1903 (N_1903,N_1198,N_1262);
and U1904 (N_1904,N_1177,N_874);
and U1905 (N_1905,N_1203,N_1019);
or U1906 (N_1906,N_902,N_1402);
nand U1907 (N_1907,N_902,N_1349);
nand U1908 (N_1908,N_1108,N_1105);
nand U1909 (N_1909,N_953,N_1367);
nor U1910 (N_1910,N_1480,N_802);
nor U1911 (N_1911,N_1012,N_994);
xor U1912 (N_1912,N_1049,N_1452);
nand U1913 (N_1913,N_1126,N_1459);
and U1914 (N_1914,N_921,N_1353);
nor U1915 (N_1915,N_1283,N_1269);
or U1916 (N_1916,N_1036,N_1137);
nor U1917 (N_1917,N_872,N_837);
and U1918 (N_1918,N_1414,N_1341);
nor U1919 (N_1919,N_946,N_1450);
and U1920 (N_1920,N_1118,N_1019);
nand U1921 (N_1921,N_962,N_1283);
nor U1922 (N_1922,N_834,N_1057);
or U1923 (N_1923,N_1331,N_1269);
nor U1924 (N_1924,N_810,N_1290);
and U1925 (N_1925,N_997,N_1066);
nand U1926 (N_1926,N_874,N_757);
nand U1927 (N_1927,N_983,N_1213);
or U1928 (N_1928,N_828,N_1266);
or U1929 (N_1929,N_1081,N_1375);
nor U1930 (N_1930,N_863,N_1063);
and U1931 (N_1931,N_851,N_1229);
and U1932 (N_1932,N_1424,N_798);
nand U1933 (N_1933,N_1344,N_1126);
nand U1934 (N_1934,N_813,N_1099);
or U1935 (N_1935,N_881,N_965);
nand U1936 (N_1936,N_1199,N_1160);
nor U1937 (N_1937,N_1319,N_995);
or U1938 (N_1938,N_762,N_1013);
and U1939 (N_1939,N_1288,N_839);
nor U1940 (N_1940,N_1116,N_1243);
nor U1941 (N_1941,N_1073,N_970);
and U1942 (N_1942,N_949,N_770);
nor U1943 (N_1943,N_1123,N_1331);
and U1944 (N_1944,N_1271,N_1157);
and U1945 (N_1945,N_928,N_1090);
or U1946 (N_1946,N_1070,N_1378);
or U1947 (N_1947,N_1180,N_1338);
and U1948 (N_1948,N_1478,N_998);
and U1949 (N_1949,N_968,N_907);
or U1950 (N_1950,N_1431,N_767);
and U1951 (N_1951,N_1027,N_1107);
nor U1952 (N_1952,N_1277,N_1443);
nand U1953 (N_1953,N_1138,N_961);
nand U1954 (N_1954,N_1245,N_984);
or U1955 (N_1955,N_1219,N_1205);
and U1956 (N_1956,N_1186,N_1209);
or U1957 (N_1957,N_764,N_846);
or U1958 (N_1958,N_1270,N_975);
nand U1959 (N_1959,N_1168,N_1319);
nor U1960 (N_1960,N_1011,N_832);
and U1961 (N_1961,N_1430,N_1005);
nor U1962 (N_1962,N_1211,N_1085);
or U1963 (N_1963,N_987,N_1014);
nand U1964 (N_1964,N_1322,N_825);
nand U1965 (N_1965,N_973,N_1463);
and U1966 (N_1966,N_1278,N_947);
and U1967 (N_1967,N_1173,N_761);
and U1968 (N_1968,N_1478,N_1367);
nor U1969 (N_1969,N_1252,N_1439);
and U1970 (N_1970,N_1276,N_885);
nand U1971 (N_1971,N_1050,N_757);
and U1972 (N_1972,N_831,N_1468);
nor U1973 (N_1973,N_1355,N_1381);
nor U1974 (N_1974,N_1261,N_1477);
or U1975 (N_1975,N_1183,N_1145);
and U1976 (N_1976,N_786,N_1377);
or U1977 (N_1977,N_757,N_892);
nor U1978 (N_1978,N_779,N_1130);
nor U1979 (N_1979,N_1081,N_1195);
and U1980 (N_1980,N_891,N_1045);
or U1981 (N_1981,N_1095,N_1241);
or U1982 (N_1982,N_751,N_1081);
nor U1983 (N_1983,N_1084,N_966);
nor U1984 (N_1984,N_1377,N_1279);
or U1985 (N_1985,N_1323,N_907);
and U1986 (N_1986,N_1238,N_900);
and U1987 (N_1987,N_1010,N_1446);
xor U1988 (N_1988,N_1408,N_1375);
and U1989 (N_1989,N_815,N_1319);
and U1990 (N_1990,N_1204,N_1141);
nand U1991 (N_1991,N_1114,N_827);
or U1992 (N_1992,N_1237,N_863);
or U1993 (N_1993,N_1182,N_1417);
nand U1994 (N_1994,N_885,N_1008);
nor U1995 (N_1995,N_1463,N_1455);
or U1996 (N_1996,N_1279,N_1222);
or U1997 (N_1997,N_951,N_982);
nor U1998 (N_1998,N_1241,N_919);
nand U1999 (N_1999,N_1015,N_1075);
nand U2000 (N_2000,N_1002,N_1370);
or U2001 (N_2001,N_1418,N_1338);
and U2002 (N_2002,N_1200,N_1312);
nand U2003 (N_2003,N_1230,N_1444);
nor U2004 (N_2004,N_931,N_864);
and U2005 (N_2005,N_1003,N_878);
and U2006 (N_2006,N_1458,N_1042);
nand U2007 (N_2007,N_1322,N_959);
nor U2008 (N_2008,N_1296,N_1421);
nand U2009 (N_2009,N_1468,N_1432);
and U2010 (N_2010,N_1427,N_795);
nand U2011 (N_2011,N_1190,N_1430);
or U2012 (N_2012,N_855,N_1182);
nor U2013 (N_2013,N_1276,N_1016);
or U2014 (N_2014,N_1309,N_1483);
nor U2015 (N_2015,N_1332,N_1010);
and U2016 (N_2016,N_1005,N_857);
or U2017 (N_2017,N_1461,N_1218);
nand U2018 (N_2018,N_1041,N_809);
and U2019 (N_2019,N_1182,N_873);
or U2020 (N_2020,N_874,N_1139);
or U2021 (N_2021,N_848,N_1407);
nor U2022 (N_2022,N_932,N_1481);
or U2023 (N_2023,N_1327,N_931);
or U2024 (N_2024,N_957,N_1412);
nand U2025 (N_2025,N_1266,N_1454);
and U2026 (N_2026,N_1310,N_1207);
nand U2027 (N_2027,N_1474,N_1072);
or U2028 (N_2028,N_1176,N_1223);
or U2029 (N_2029,N_1338,N_1208);
nor U2030 (N_2030,N_1142,N_1033);
or U2031 (N_2031,N_968,N_1182);
or U2032 (N_2032,N_1199,N_1410);
nor U2033 (N_2033,N_1142,N_1189);
and U2034 (N_2034,N_1208,N_1334);
nor U2035 (N_2035,N_1473,N_896);
nor U2036 (N_2036,N_851,N_1424);
or U2037 (N_2037,N_1235,N_830);
or U2038 (N_2038,N_1131,N_1381);
nor U2039 (N_2039,N_1413,N_1182);
nor U2040 (N_2040,N_913,N_1114);
or U2041 (N_2041,N_1497,N_1486);
and U2042 (N_2042,N_871,N_1095);
or U2043 (N_2043,N_1339,N_1163);
nor U2044 (N_2044,N_1280,N_803);
or U2045 (N_2045,N_922,N_858);
or U2046 (N_2046,N_772,N_1396);
nand U2047 (N_2047,N_1467,N_831);
and U2048 (N_2048,N_785,N_1464);
nand U2049 (N_2049,N_1259,N_1124);
or U2050 (N_2050,N_1136,N_874);
or U2051 (N_2051,N_1454,N_969);
or U2052 (N_2052,N_1136,N_940);
or U2053 (N_2053,N_792,N_1035);
and U2054 (N_2054,N_1259,N_1474);
nand U2055 (N_2055,N_904,N_1480);
or U2056 (N_2056,N_1319,N_770);
nand U2057 (N_2057,N_1072,N_978);
and U2058 (N_2058,N_1223,N_754);
or U2059 (N_2059,N_935,N_1012);
and U2060 (N_2060,N_1117,N_1107);
nor U2061 (N_2061,N_1293,N_1143);
and U2062 (N_2062,N_949,N_803);
or U2063 (N_2063,N_1249,N_1138);
or U2064 (N_2064,N_929,N_1480);
nand U2065 (N_2065,N_1413,N_1149);
or U2066 (N_2066,N_1058,N_976);
nor U2067 (N_2067,N_1173,N_1290);
or U2068 (N_2068,N_787,N_1452);
nand U2069 (N_2069,N_1018,N_1171);
nor U2070 (N_2070,N_1088,N_1194);
or U2071 (N_2071,N_1201,N_1131);
or U2072 (N_2072,N_1436,N_814);
and U2073 (N_2073,N_1316,N_845);
nor U2074 (N_2074,N_1135,N_960);
or U2075 (N_2075,N_1164,N_1225);
or U2076 (N_2076,N_819,N_1117);
and U2077 (N_2077,N_1277,N_1215);
or U2078 (N_2078,N_1187,N_799);
nand U2079 (N_2079,N_1451,N_1462);
or U2080 (N_2080,N_1074,N_751);
or U2081 (N_2081,N_1324,N_1289);
nor U2082 (N_2082,N_879,N_958);
nor U2083 (N_2083,N_1180,N_1471);
and U2084 (N_2084,N_962,N_873);
nor U2085 (N_2085,N_880,N_1357);
nor U2086 (N_2086,N_773,N_901);
nand U2087 (N_2087,N_888,N_769);
nand U2088 (N_2088,N_1141,N_1363);
and U2089 (N_2089,N_1024,N_1277);
or U2090 (N_2090,N_939,N_1355);
or U2091 (N_2091,N_878,N_1429);
nor U2092 (N_2092,N_1231,N_1386);
or U2093 (N_2093,N_865,N_1143);
nand U2094 (N_2094,N_1267,N_1211);
or U2095 (N_2095,N_1171,N_1470);
and U2096 (N_2096,N_1403,N_760);
and U2097 (N_2097,N_1343,N_1265);
or U2098 (N_2098,N_1013,N_1319);
nor U2099 (N_2099,N_1131,N_1128);
nor U2100 (N_2100,N_1044,N_787);
and U2101 (N_2101,N_987,N_1034);
and U2102 (N_2102,N_1124,N_1069);
or U2103 (N_2103,N_1449,N_793);
and U2104 (N_2104,N_921,N_1032);
nand U2105 (N_2105,N_1223,N_784);
nand U2106 (N_2106,N_1112,N_1273);
and U2107 (N_2107,N_1011,N_939);
nor U2108 (N_2108,N_1271,N_984);
or U2109 (N_2109,N_977,N_1490);
nor U2110 (N_2110,N_1192,N_777);
or U2111 (N_2111,N_1297,N_1266);
and U2112 (N_2112,N_977,N_1145);
nand U2113 (N_2113,N_1250,N_1074);
and U2114 (N_2114,N_1099,N_999);
nand U2115 (N_2115,N_1238,N_871);
nand U2116 (N_2116,N_933,N_899);
or U2117 (N_2117,N_783,N_951);
nand U2118 (N_2118,N_1499,N_825);
or U2119 (N_2119,N_1229,N_1374);
and U2120 (N_2120,N_854,N_998);
nor U2121 (N_2121,N_1329,N_930);
nand U2122 (N_2122,N_1047,N_1106);
nor U2123 (N_2123,N_1063,N_1176);
or U2124 (N_2124,N_1049,N_864);
nand U2125 (N_2125,N_1266,N_1439);
or U2126 (N_2126,N_1344,N_1304);
nor U2127 (N_2127,N_1153,N_1095);
or U2128 (N_2128,N_1179,N_1441);
nand U2129 (N_2129,N_931,N_1104);
nand U2130 (N_2130,N_1098,N_903);
nor U2131 (N_2131,N_1477,N_1284);
or U2132 (N_2132,N_1378,N_1347);
nand U2133 (N_2133,N_782,N_843);
and U2134 (N_2134,N_861,N_1219);
xnor U2135 (N_2135,N_773,N_1401);
nand U2136 (N_2136,N_813,N_1351);
nor U2137 (N_2137,N_1325,N_1096);
nor U2138 (N_2138,N_994,N_1331);
xor U2139 (N_2139,N_1272,N_1443);
nor U2140 (N_2140,N_1418,N_1152);
and U2141 (N_2141,N_1029,N_1229);
nor U2142 (N_2142,N_908,N_986);
or U2143 (N_2143,N_982,N_1437);
nor U2144 (N_2144,N_1120,N_1110);
nor U2145 (N_2145,N_1209,N_1077);
nand U2146 (N_2146,N_1275,N_1080);
and U2147 (N_2147,N_1212,N_1282);
and U2148 (N_2148,N_1456,N_799);
nand U2149 (N_2149,N_1376,N_1136);
and U2150 (N_2150,N_1176,N_1466);
or U2151 (N_2151,N_865,N_1399);
nand U2152 (N_2152,N_1336,N_1361);
and U2153 (N_2153,N_767,N_1211);
nand U2154 (N_2154,N_1135,N_1312);
and U2155 (N_2155,N_1298,N_1347);
or U2156 (N_2156,N_984,N_963);
nand U2157 (N_2157,N_855,N_1448);
nor U2158 (N_2158,N_1084,N_1385);
and U2159 (N_2159,N_1305,N_1337);
nand U2160 (N_2160,N_1449,N_981);
nand U2161 (N_2161,N_1039,N_1173);
nor U2162 (N_2162,N_1355,N_1218);
or U2163 (N_2163,N_1037,N_927);
and U2164 (N_2164,N_938,N_1362);
nand U2165 (N_2165,N_810,N_874);
nand U2166 (N_2166,N_1359,N_1167);
nor U2167 (N_2167,N_910,N_1373);
or U2168 (N_2168,N_1251,N_1271);
or U2169 (N_2169,N_1134,N_1051);
nor U2170 (N_2170,N_1450,N_1115);
nand U2171 (N_2171,N_1349,N_1422);
nand U2172 (N_2172,N_1371,N_893);
and U2173 (N_2173,N_1381,N_765);
nor U2174 (N_2174,N_1063,N_1055);
or U2175 (N_2175,N_1264,N_1422);
or U2176 (N_2176,N_844,N_1120);
or U2177 (N_2177,N_941,N_1343);
nor U2178 (N_2178,N_952,N_1413);
nor U2179 (N_2179,N_1493,N_1118);
and U2180 (N_2180,N_1227,N_1291);
nor U2181 (N_2181,N_1138,N_989);
and U2182 (N_2182,N_1384,N_1087);
nor U2183 (N_2183,N_1007,N_963);
and U2184 (N_2184,N_1229,N_1494);
and U2185 (N_2185,N_1128,N_1468);
nand U2186 (N_2186,N_1363,N_934);
nand U2187 (N_2187,N_1472,N_1397);
and U2188 (N_2188,N_1334,N_908);
nand U2189 (N_2189,N_1369,N_870);
nor U2190 (N_2190,N_753,N_1334);
or U2191 (N_2191,N_1472,N_1367);
nand U2192 (N_2192,N_1138,N_1226);
or U2193 (N_2193,N_1332,N_832);
nand U2194 (N_2194,N_1286,N_1014);
nand U2195 (N_2195,N_798,N_1220);
or U2196 (N_2196,N_1157,N_774);
nand U2197 (N_2197,N_917,N_813);
nand U2198 (N_2198,N_930,N_1067);
and U2199 (N_2199,N_812,N_980);
or U2200 (N_2200,N_819,N_1433);
and U2201 (N_2201,N_1462,N_972);
or U2202 (N_2202,N_1385,N_1238);
nor U2203 (N_2203,N_1325,N_1378);
or U2204 (N_2204,N_1437,N_867);
nor U2205 (N_2205,N_778,N_1483);
or U2206 (N_2206,N_1206,N_1323);
nor U2207 (N_2207,N_1395,N_1015);
nand U2208 (N_2208,N_1227,N_1276);
nand U2209 (N_2209,N_758,N_1151);
or U2210 (N_2210,N_1368,N_1205);
nor U2211 (N_2211,N_1251,N_1003);
or U2212 (N_2212,N_1213,N_772);
and U2213 (N_2213,N_763,N_932);
or U2214 (N_2214,N_973,N_1288);
and U2215 (N_2215,N_1371,N_1101);
nor U2216 (N_2216,N_866,N_895);
and U2217 (N_2217,N_767,N_1283);
nand U2218 (N_2218,N_1046,N_1225);
or U2219 (N_2219,N_897,N_1486);
nand U2220 (N_2220,N_1104,N_1439);
nand U2221 (N_2221,N_1395,N_1299);
or U2222 (N_2222,N_1361,N_1286);
nand U2223 (N_2223,N_1062,N_1185);
and U2224 (N_2224,N_1312,N_1102);
or U2225 (N_2225,N_1130,N_1132);
nor U2226 (N_2226,N_939,N_1083);
and U2227 (N_2227,N_978,N_1467);
nor U2228 (N_2228,N_815,N_1161);
nor U2229 (N_2229,N_805,N_828);
nor U2230 (N_2230,N_838,N_845);
and U2231 (N_2231,N_1459,N_1076);
nand U2232 (N_2232,N_1113,N_1014);
and U2233 (N_2233,N_1258,N_758);
or U2234 (N_2234,N_1369,N_806);
nor U2235 (N_2235,N_858,N_1211);
or U2236 (N_2236,N_1250,N_1437);
and U2237 (N_2237,N_1356,N_985);
nand U2238 (N_2238,N_1462,N_870);
or U2239 (N_2239,N_926,N_1065);
nor U2240 (N_2240,N_788,N_962);
nand U2241 (N_2241,N_799,N_1373);
and U2242 (N_2242,N_782,N_825);
xnor U2243 (N_2243,N_1472,N_945);
and U2244 (N_2244,N_1226,N_782);
and U2245 (N_2245,N_1021,N_1170);
and U2246 (N_2246,N_876,N_972);
nor U2247 (N_2247,N_990,N_823);
and U2248 (N_2248,N_938,N_793);
xor U2249 (N_2249,N_884,N_1357);
nand U2250 (N_2250,N_1768,N_1934);
nand U2251 (N_2251,N_2227,N_1727);
or U2252 (N_2252,N_1619,N_2002);
and U2253 (N_2253,N_1938,N_1696);
and U2254 (N_2254,N_2130,N_1943);
nand U2255 (N_2255,N_1910,N_1530);
nand U2256 (N_2256,N_1911,N_1881);
nor U2257 (N_2257,N_1549,N_1793);
nand U2258 (N_2258,N_1571,N_1543);
nand U2259 (N_2259,N_1959,N_2137);
and U2260 (N_2260,N_2244,N_1994);
nor U2261 (N_2261,N_2077,N_1761);
nand U2262 (N_2262,N_2123,N_2019);
or U2263 (N_2263,N_2084,N_2201);
nor U2264 (N_2264,N_2057,N_1838);
nor U2265 (N_2265,N_2075,N_1947);
and U2266 (N_2266,N_1979,N_1770);
and U2267 (N_2267,N_1627,N_2173);
and U2268 (N_2268,N_1939,N_1975);
xnor U2269 (N_2269,N_1713,N_1992);
or U2270 (N_2270,N_1950,N_1836);
or U2271 (N_2271,N_2204,N_1822);
nor U2272 (N_2272,N_1623,N_1781);
nor U2273 (N_2273,N_1830,N_2016);
or U2274 (N_2274,N_2004,N_1574);
or U2275 (N_2275,N_2103,N_2199);
and U2276 (N_2276,N_1841,N_1964);
and U2277 (N_2277,N_1922,N_2117);
nor U2278 (N_2278,N_2000,N_1717);
xnor U2279 (N_2279,N_1692,N_2226);
and U2280 (N_2280,N_2025,N_2194);
and U2281 (N_2281,N_1594,N_2022);
and U2282 (N_2282,N_2098,N_2131);
and U2283 (N_2283,N_1519,N_1755);
or U2284 (N_2284,N_1779,N_2072);
and U2285 (N_2285,N_1652,N_2190);
or U2286 (N_2286,N_1883,N_1885);
nor U2287 (N_2287,N_2206,N_1699);
nand U2288 (N_2288,N_1752,N_1832);
nand U2289 (N_2289,N_1977,N_2221);
nor U2290 (N_2290,N_1579,N_1909);
or U2291 (N_2291,N_1914,N_1746);
nor U2292 (N_2292,N_2110,N_1509);
and U2293 (N_2293,N_2064,N_2030);
and U2294 (N_2294,N_1595,N_2026);
or U2295 (N_2295,N_1735,N_1680);
and U2296 (N_2296,N_1502,N_1695);
nand U2297 (N_2297,N_1917,N_2198);
and U2298 (N_2298,N_1672,N_1645);
or U2299 (N_2299,N_1702,N_1892);
or U2300 (N_2300,N_2050,N_2053);
nand U2301 (N_2301,N_1960,N_2178);
nor U2302 (N_2302,N_1511,N_2200);
nor U2303 (N_2303,N_1902,N_1870);
nor U2304 (N_2304,N_1775,N_1691);
nor U2305 (N_2305,N_1551,N_2031);
and U2306 (N_2306,N_1846,N_2008);
nor U2307 (N_2307,N_2018,N_1864);
nor U2308 (N_2308,N_1908,N_1617);
nor U2309 (N_2309,N_1585,N_1811);
or U2310 (N_2310,N_1515,N_1679);
nand U2311 (N_2311,N_1721,N_2024);
nand U2312 (N_2312,N_1807,N_2146);
or U2313 (N_2313,N_2055,N_1854);
or U2314 (N_2314,N_1527,N_1921);
or U2315 (N_2315,N_2073,N_1641);
nand U2316 (N_2316,N_2186,N_2080);
or U2317 (N_2317,N_2115,N_1657);
nor U2318 (N_2318,N_1941,N_2248);
and U2319 (N_2319,N_2195,N_1850);
nor U2320 (N_2320,N_2164,N_1654);
nand U2321 (N_2321,N_1969,N_1655);
nand U2322 (N_2322,N_2187,N_1971);
or U2323 (N_2323,N_1905,N_1681);
nand U2324 (N_2324,N_1820,N_1806);
nand U2325 (N_2325,N_2021,N_2143);
or U2326 (N_2326,N_1760,N_1804);
and U2327 (N_2327,N_1884,N_1895);
nand U2328 (N_2328,N_1833,N_1690);
nand U2329 (N_2329,N_1631,N_1757);
nor U2330 (N_2330,N_1732,N_2219);
and U2331 (N_2331,N_2136,N_1993);
or U2332 (N_2332,N_1665,N_1698);
nand U2333 (N_2333,N_2176,N_1687);
nor U2334 (N_2334,N_1714,N_2013);
nand U2335 (N_2335,N_1739,N_1728);
xnor U2336 (N_2336,N_2069,N_1888);
and U2337 (N_2337,N_1925,N_1569);
and U2338 (N_2338,N_1565,N_1988);
nand U2339 (N_2339,N_2135,N_1852);
nor U2340 (N_2340,N_1512,N_1664);
nor U2341 (N_2341,N_1622,N_1896);
and U2342 (N_2342,N_1916,N_1995);
nor U2343 (N_2343,N_1923,N_1765);
and U2344 (N_2344,N_1961,N_1991);
nor U2345 (N_2345,N_1869,N_1843);
nor U2346 (N_2346,N_2154,N_2092);
nand U2347 (N_2347,N_2066,N_1842);
and U2348 (N_2348,N_1951,N_1706);
and U2349 (N_2349,N_1650,N_2197);
nor U2350 (N_2350,N_2249,N_1879);
and U2351 (N_2351,N_1694,N_1827);
and U2352 (N_2352,N_1747,N_1928);
or U2353 (N_2353,N_2011,N_1797);
and U2354 (N_2354,N_1748,N_2202);
or U2355 (N_2355,N_1777,N_2116);
and U2356 (N_2356,N_2017,N_2168);
nor U2357 (N_2357,N_1766,N_1889);
or U2358 (N_2358,N_2047,N_1987);
nor U2359 (N_2359,N_1611,N_1535);
nor U2360 (N_2360,N_1981,N_1886);
or U2361 (N_2361,N_2074,N_2104);
or U2362 (N_2362,N_2045,N_1558);
and U2363 (N_2363,N_1956,N_1500);
nor U2364 (N_2364,N_2010,N_1897);
nor U2365 (N_2365,N_1999,N_1718);
or U2366 (N_2366,N_1805,N_1857);
or U2367 (N_2367,N_1784,N_2222);
nor U2368 (N_2368,N_2231,N_1828);
and U2369 (N_2369,N_1659,N_1904);
and U2370 (N_2370,N_1685,N_1529);
or U2371 (N_2371,N_2238,N_1965);
nand U2372 (N_2372,N_2211,N_1568);
nand U2373 (N_2373,N_2078,N_2079);
nor U2374 (N_2374,N_2169,N_1986);
and U2375 (N_2375,N_1704,N_1601);
nand U2376 (N_2376,N_1546,N_1609);
and U2377 (N_2377,N_1588,N_1762);
or U2378 (N_2378,N_1693,N_1505);
nand U2379 (N_2379,N_1637,N_1821);
or U2380 (N_2380,N_1788,N_1602);
and U2381 (N_2381,N_1867,N_2127);
nor U2382 (N_2382,N_1554,N_1572);
and U2383 (N_2383,N_1974,N_1773);
nor U2384 (N_2384,N_2145,N_1686);
and U2385 (N_2385,N_1658,N_2189);
nand U2386 (N_2386,N_2237,N_1935);
nand U2387 (N_2387,N_1570,N_1963);
and U2388 (N_2388,N_1890,N_2241);
nand U2389 (N_2389,N_1847,N_1639);
or U2390 (N_2390,N_1872,N_1859);
nand U2391 (N_2391,N_1591,N_1719);
or U2392 (N_2392,N_1855,N_1948);
or U2393 (N_2393,N_1849,N_1978);
nand U2394 (N_2394,N_1756,N_1697);
nand U2395 (N_2395,N_2183,N_2093);
nor U2396 (N_2396,N_1801,N_1526);
and U2397 (N_2397,N_2081,N_1845);
or U2398 (N_2398,N_1782,N_2128);
or U2399 (N_2399,N_1815,N_1944);
nor U2400 (N_2400,N_1638,N_1933);
or U2401 (N_2401,N_1539,N_1576);
nor U2402 (N_2402,N_2179,N_1656);
nand U2403 (N_2403,N_1523,N_2003);
or U2404 (N_2404,N_1513,N_1644);
and U2405 (N_2405,N_1898,N_1731);
nand U2406 (N_2406,N_1837,N_2082);
or U2407 (N_2407,N_1990,N_1774);
or U2408 (N_2408,N_1624,N_1940);
and U2409 (N_2409,N_1703,N_1592);
and U2410 (N_2410,N_1982,N_2102);
nand U2411 (N_2411,N_2174,N_2140);
or U2412 (N_2412,N_1678,N_1682);
or U2413 (N_2413,N_1649,N_1751);
nand U2414 (N_2414,N_1534,N_1817);
and U2415 (N_2415,N_2124,N_2165);
nand U2416 (N_2416,N_1802,N_1651);
or U2417 (N_2417,N_2193,N_2027);
or U2418 (N_2418,N_1813,N_2063);
or U2419 (N_2419,N_1531,N_1796);
nor U2420 (N_2420,N_1737,N_2015);
nand U2421 (N_2421,N_2091,N_1553);
or U2422 (N_2422,N_1967,N_2245);
nand U2423 (N_2423,N_1522,N_1630);
or U2424 (N_2424,N_2240,N_2109);
and U2425 (N_2425,N_1603,N_1520);
nor U2426 (N_2426,N_1606,N_1640);
nand U2427 (N_2427,N_1789,N_2218);
or U2428 (N_2428,N_1901,N_1771);
nor U2429 (N_2429,N_2039,N_1607);
and U2430 (N_2430,N_1557,N_1734);
nand U2431 (N_2431,N_2217,N_1671);
nor U2432 (N_2432,N_1517,N_1545);
and U2433 (N_2433,N_2108,N_1725);
nand U2434 (N_2434,N_2067,N_2223);
nor U2435 (N_2435,N_2121,N_2106);
and U2436 (N_2436,N_1736,N_2007);
and U2437 (N_2437,N_1575,N_2185);
or U2438 (N_2438,N_1794,N_1873);
and U2439 (N_2439,N_2134,N_2032);
or U2440 (N_2440,N_2161,N_2196);
or U2441 (N_2441,N_1581,N_2094);
nand U2442 (N_2442,N_1868,N_1810);
or U2443 (N_2443,N_1894,N_2099);
or U2444 (N_2444,N_1912,N_2001);
nor U2445 (N_2445,N_1878,N_1730);
nand U2446 (N_2446,N_2167,N_2139);
or U2447 (N_2447,N_2118,N_1976);
and U2448 (N_2448,N_2236,N_1809);
nand U2449 (N_2449,N_1937,N_1663);
or U2450 (N_2450,N_2155,N_1560);
nand U2451 (N_2451,N_2048,N_1738);
nor U2452 (N_2452,N_1626,N_1839);
and U2453 (N_2453,N_1688,N_1767);
nor U2454 (N_2454,N_1753,N_1660);
nand U2455 (N_2455,N_2180,N_1548);
xnor U2456 (N_2456,N_1858,N_2229);
and U2457 (N_2457,N_1628,N_1791);
nand U2458 (N_2458,N_1880,N_1701);
or U2459 (N_2459,N_1899,N_1700);
or U2460 (N_2460,N_1945,N_1620);
nor U2461 (N_2461,N_2162,N_2028);
or U2462 (N_2462,N_2060,N_1547);
nor U2463 (N_2463,N_2156,N_1599);
nor U2464 (N_2464,N_2051,N_2083);
nor U2465 (N_2465,N_1983,N_1742);
nand U2466 (N_2466,N_2037,N_1642);
nor U2467 (N_2467,N_1516,N_1772);
or U2468 (N_2468,N_2038,N_2170);
and U2469 (N_2469,N_1882,N_1653);
nor U2470 (N_2470,N_1799,N_2184);
and U2471 (N_2471,N_1920,N_2150);
nor U2472 (N_2472,N_1521,N_1893);
nor U2473 (N_2473,N_2023,N_1612);
nand U2474 (N_2474,N_1844,N_1705);
and U2475 (N_2475,N_2171,N_1544);
and U2476 (N_2476,N_1863,N_2006);
nor U2477 (N_2477,N_1524,N_1862);
or U2478 (N_2478,N_2177,N_1812);
nor U2479 (N_2479,N_1600,N_2182);
or U2480 (N_2480,N_1887,N_2228);
or U2481 (N_2481,N_2141,N_1724);
and U2482 (N_2482,N_2166,N_1851);
nand U2483 (N_2483,N_2086,N_1831);
nor U2484 (N_2484,N_1754,N_2076);
and U2485 (N_2485,N_2046,N_1996);
nand U2486 (N_2486,N_1953,N_2142);
nor U2487 (N_2487,N_1763,N_1783);
and U2488 (N_2488,N_2157,N_2230);
or U2489 (N_2489,N_1528,N_2090);
and U2490 (N_2490,N_1997,N_1795);
nand U2491 (N_2491,N_1798,N_2163);
or U2492 (N_2492,N_1615,N_1877);
nand U2493 (N_2493,N_2052,N_1677);
nand U2494 (N_2494,N_2040,N_1552);
and U2495 (N_2495,N_1675,N_1764);
nand U2496 (N_2496,N_2192,N_1954);
nand U2497 (N_2497,N_1936,N_1533);
or U2498 (N_2498,N_2159,N_1741);
nor U2499 (N_2499,N_2041,N_1707);
and U2500 (N_2500,N_1584,N_1712);
nor U2501 (N_2501,N_2151,N_1913);
and U2502 (N_2502,N_2208,N_1930);
nor U2503 (N_2503,N_1587,N_1668);
and U2504 (N_2504,N_2087,N_1740);
or U2505 (N_2505,N_2056,N_2020);
or U2506 (N_2506,N_1559,N_1929);
or U2507 (N_2507,N_1643,N_1563);
and U2508 (N_2508,N_1818,N_1708);
or U2509 (N_2509,N_1776,N_1932);
or U2510 (N_2510,N_2036,N_1667);
or U2511 (N_2511,N_1745,N_1583);
nand U2512 (N_2512,N_1790,N_1669);
xnor U2513 (N_2513,N_2224,N_1876);
or U2514 (N_2514,N_1952,N_1673);
nor U2515 (N_2515,N_2029,N_1564);
nand U2516 (N_2516,N_1662,N_2235);
nand U2517 (N_2517,N_1787,N_2209);
or U2518 (N_2518,N_2233,N_1968);
nor U2519 (N_2519,N_2133,N_1871);
and U2520 (N_2520,N_1891,N_1972);
or U2521 (N_2521,N_2068,N_2203);
nor U2522 (N_2522,N_2112,N_1834);
or U2523 (N_2523,N_1927,N_2070);
and U2524 (N_2524,N_2111,N_1984);
or U2525 (N_2525,N_2096,N_1621);
nand U2526 (N_2526,N_2239,N_1989);
and U2527 (N_2527,N_2188,N_2243);
nor U2528 (N_2528,N_1556,N_1723);
nand U2529 (N_2529,N_2005,N_1538);
and U2530 (N_2530,N_1785,N_1573);
nor U2531 (N_2531,N_2062,N_1618);
and U2532 (N_2532,N_2153,N_1726);
and U2533 (N_2533,N_2126,N_1501);
and U2534 (N_2534,N_2119,N_1605);
nor U2535 (N_2535,N_1826,N_1924);
nand U2536 (N_2536,N_2172,N_1633);
and U2537 (N_2537,N_2246,N_1759);
and U2538 (N_2538,N_1962,N_1590);
or U2539 (N_2539,N_1792,N_1980);
or U2540 (N_2540,N_2210,N_1875);
or U2541 (N_2541,N_2129,N_1958);
and U2542 (N_2542,N_1729,N_1758);
and U2543 (N_2543,N_2242,N_1710);
nand U2544 (N_2544,N_2215,N_2042);
and U2545 (N_2545,N_2100,N_2232);
or U2546 (N_2546,N_2138,N_2059);
nor U2547 (N_2547,N_1973,N_1503);
nand U2548 (N_2548,N_1865,N_1586);
and U2549 (N_2549,N_1541,N_1848);
nand U2550 (N_2550,N_1814,N_1646);
and U2551 (N_2551,N_1536,N_2049);
nor U2552 (N_2552,N_2144,N_1949);
and U2553 (N_2553,N_1780,N_1998);
or U2554 (N_2554,N_1715,N_1537);
nor U2555 (N_2555,N_1593,N_1825);
and U2556 (N_2556,N_1610,N_2088);
nor U2557 (N_2557,N_2101,N_1808);
nand U2558 (N_2558,N_2212,N_2191);
nand U2559 (N_2559,N_1733,N_1900);
or U2560 (N_2560,N_2234,N_1540);
or U2561 (N_2561,N_2085,N_1684);
or U2562 (N_2562,N_1578,N_1824);
or U2563 (N_2563,N_2181,N_2225);
nand U2564 (N_2564,N_2095,N_1518);
or U2565 (N_2565,N_2089,N_2132);
and U2566 (N_2566,N_2152,N_2058);
nand U2567 (N_2567,N_2216,N_1504);
or U2568 (N_2568,N_1566,N_1907);
nor U2569 (N_2569,N_1510,N_2097);
nand U2570 (N_2570,N_1647,N_1634);
and U2571 (N_2571,N_1743,N_1625);
or U2572 (N_2572,N_2175,N_1955);
or U2573 (N_2573,N_2033,N_1931);
nand U2574 (N_2574,N_1596,N_2113);
or U2575 (N_2575,N_1648,N_2034);
and U2576 (N_2576,N_1632,N_1856);
or U2577 (N_2577,N_1819,N_1966);
and U2578 (N_2578,N_2205,N_1716);
and U2579 (N_2579,N_2120,N_1970);
or U2580 (N_2580,N_1903,N_2214);
nand U2581 (N_2581,N_1555,N_2158);
or U2582 (N_2582,N_1514,N_1722);
and U2583 (N_2583,N_1750,N_1749);
nand U2584 (N_2584,N_1709,N_1598);
nand U2585 (N_2585,N_1582,N_1635);
nor U2586 (N_2586,N_1918,N_2054);
nand U2587 (N_2587,N_2149,N_1507);
nand U2588 (N_2588,N_1711,N_2107);
nand U2589 (N_2589,N_1720,N_1915);
xor U2590 (N_2590,N_1769,N_2207);
nand U2591 (N_2591,N_2071,N_1957);
nand U2592 (N_2592,N_1542,N_2065);
nand U2593 (N_2593,N_1942,N_2012);
nor U2594 (N_2594,N_1604,N_2125);
or U2595 (N_2595,N_2213,N_2114);
and U2596 (N_2596,N_2044,N_2014);
nor U2597 (N_2597,N_1874,N_1589);
or U2598 (N_2598,N_2105,N_1866);
or U2599 (N_2599,N_1985,N_1778);
and U2600 (N_2600,N_1636,N_1616);
xor U2601 (N_2601,N_1580,N_1674);
or U2602 (N_2602,N_1840,N_1613);
nor U2603 (N_2603,N_1786,N_1689);
nand U2604 (N_2604,N_2148,N_2147);
nand U2605 (N_2605,N_1861,N_1661);
or U2606 (N_2606,N_1676,N_1835);
or U2607 (N_2607,N_1550,N_2061);
nand U2608 (N_2608,N_2122,N_2247);
nor U2609 (N_2609,N_2220,N_1577);
and U2610 (N_2610,N_1803,N_1562);
nand U2611 (N_2611,N_1506,N_2009);
and U2612 (N_2612,N_1597,N_1683);
nand U2613 (N_2613,N_1860,N_2035);
or U2614 (N_2614,N_1816,N_1926);
or U2615 (N_2615,N_1823,N_1561);
and U2616 (N_2616,N_1919,N_1567);
and U2617 (N_2617,N_1508,N_1629);
nand U2618 (N_2618,N_1532,N_1614);
and U2619 (N_2619,N_2160,N_1608);
nand U2620 (N_2620,N_1670,N_1800);
nand U2621 (N_2621,N_1525,N_1906);
or U2622 (N_2622,N_1666,N_1744);
and U2623 (N_2623,N_1829,N_1853);
nor U2624 (N_2624,N_1946,N_2043);
and U2625 (N_2625,N_1902,N_1840);
and U2626 (N_2626,N_1569,N_2159);
nor U2627 (N_2627,N_2226,N_1636);
nand U2628 (N_2628,N_1869,N_1555);
and U2629 (N_2629,N_2046,N_1525);
nand U2630 (N_2630,N_1825,N_2230);
nor U2631 (N_2631,N_2148,N_2211);
or U2632 (N_2632,N_2051,N_1831);
nor U2633 (N_2633,N_1524,N_1977);
or U2634 (N_2634,N_2199,N_1844);
nand U2635 (N_2635,N_1972,N_1706);
nand U2636 (N_2636,N_1544,N_1506);
and U2637 (N_2637,N_1690,N_1546);
nand U2638 (N_2638,N_2123,N_2033);
and U2639 (N_2639,N_1630,N_1692);
nand U2640 (N_2640,N_1994,N_1987);
nor U2641 (N_2641,N_1543,N_1800);
nand U2642 (N_2642,N_2245,N_1867);
nand U2643 (N_2643,N_1515,N_1583);
or U2644 (N_2644,N_1803,N_2017);
nand U2645 (N_2645,N_2143,N_2245);
or U2646 (N_2646,N_1767,N_2011);
and U2647 (N_2647,N_2195,N_1992);
nor U2648 (N_2648,N_2223,N_1795);
nand U2649 (N_2649,N_2143,N_2069);
or U2650 (N_2650,N_1958,N_1652);
nand U2651 (N_2651,N_2096,N_1671);
and U2652 (N_2652,N_1551,N_1666);
or U2653 (N_2653,N_1886,N_1901);
nand U2654 (N_2654,N_1977,N_1792);
nand U2655 (N_2655,N_2022,N_2057);
and U2656 (N_2656,N_1720,N_1800);
nor U2657 (N_2657,N_2198,N_1690);
or U2658 (N_2658,N_1870,N_1895);
nor U2659 (N_2659,N_1535,N_1872);
or U2660 (N_2660,N_1649,N_1753);
and U2661 (N_2661,N_1815,N_1747);
and U2662 (N_2662,N_2121,N_1993);
xnor U2663 (N_2663,N_1555,N_2192);
or U2664 (N_2664,N_1906,N_1734);
nor U2665 (N_2665,N_1818,N_2058);
nor U2666 (N_2666,N_2052,N_1703);
nor U2667 (N_2667,N_1570,N_2205);
nor U2668 (N_2668,N_2179,N_1828);
nor U2669 (N_2669,N_2051,N_2054);
nand U2670 (N_2670,N_1870,N_2122);
nand U2671 (N_2671,N_2191,N_2201);
nor U2672 (N_2672,N_1683,N_2020);
nor U2673 (N_2673,N_1568,N_2226);
nor U2674 (N_2674,N_1915,N_2229);
and U2675 (N_2675,N_2081,N_2228);
or U2676 (N_2676,N_1537,N_1993);
and U2677 (N_2677,N_1867,N_1920);
or U2678 (N_2678,N_1595,N_2013);
xor U2679 (N_2679,N_1983,N_1784);
nand U2680 (N_2680,N_1566,N_2016);
or U2681 (N_2681,N_2100,N_2035);
nor U2682 (N_2682,N_1527,N_2001);
and U2683 (N_2683,N_2245,N_1922);
or U2684 (N_2684,N_1645,N_2154);
nand U2685 (N_2685,N_1676,N_1504);
nor U2686 (N_2686,N_2090,N_2009);
nand U2687 (N_2687,N_1546,N_1911);
nor U2688 (N_2688,N_1930,N_1970);
and U2689 (N_2689,N_1634,N_1948);
or U2690 (N_2690,N_1814,N_1868);
or U2691 (N_2691,N_2201,N_1825);
nand U2692 (N_2692,N_1695,N_1840);
nor U2693 (N_2693,N_1818,N_2019);
and U2694 (N_2694,N_1741,N_1574);
nor U2695 (N_2695,N_1546,N_1583);
and U2696 (N_2696,N_1830,N_1503);
nor U2697 (N_2697,N_1807,N_2048);
or U2698 (N_2698,N_1697,N_1946);
and U2699 (N_2699,N_1800,N_1983);
and U2700 (N_2700,N_1519,N_1677);
and U2701 (N_2701,N_1660,N_2076);
nor U2702 (N_2702,N_1595,N_2014);
nor U2703 (N_2703,N_1896,N_1702);
and U2704 (N_2704,N_2215,N_1807);
and U2705 (N_2705,N_2105,N_1564);
and U2706 (N_2706,N_1585,N_2215);
and U2707 (N_2707,N_1809,N_1739);
nand U2708 (N_2708,N_2007,N_1765);
or U2709 (N_2709,N_1546,N_2148);
or U2710 (N_2710,N_1823,N_1623);
and U2711 (N_2711,N_1543,N_1630);
and U2712 (N_2712,N_1887,N_1978);
nor U2713 (N_2713,N_1754,N_1706);
nor U2714 (N_2714,N_1681,N_1501);
and U2715 (N_2715,N_1980,N_2014);
nand U2716 (N_2716,N_2092,N_1775);
nor U2717 (N_2717,N_1957,N_1678);
and U2718 (N_2718,N_1587,N_1612);
or U2719 (N_2719,N_1585,N_2246);
nand U2720 (N_2720,N_2007,N_1813);
and U2721 (N_2721,N_2135,N_1715);
and U2722 (N_2722,N_1850,N_1576);
nor U2723 (N_2723,N_1689,N_2217);
nand U2724 (N_2724,N_2021,N_2212);
or U2725 (N_2725,N_2092,N_1533);
and U2726 (N_2726,N_1513,N_2164);
nand U2727 (N_2727,N_1908,N_2047);
and U2728 (N_2728,N_2205,N_1894);
nor U2729 (N_2729,N_2064,N_1605);
and U2730 (N_2730,N_1918,N_1902);
nor U2731 (N_2731,N_1597,N_2000);
nor U2732 (N_2732,N_2104,N_1768);
or U2733 (N_2733,N_1660,N_1984);
and U2734 (N_2734,N_2032,N_1851);
or U2735 (N_2735,N_1506,N_2190);
nand U2736 (N_2736,N_1607,N_1903);
nor U2737 (N_2737,N_1731,N_1976);
nand U2738 (N_2738,N_1517,N_2042);
xnor U2739 (N_2739,N_1530,N_1807);
or U2740 (N_2740,N_1618,N_1742);
nor U2741 (N_2741,N_1797,N_2118);
and U2742 (N_2742,N_2021,N_1539);
and U2743 (N_2743,N_2167,N_2018);
and U2744 (N_2744,N_1989,N_1988);
and U2745 (N_2745,N_1923,N_2188);
or U2746 (N_2746,N_1637,N_2080);
and U2747 (N_2747,N_2170,N_1707);
nand U2748 (N_2748,N_1857,N_1599);
and U2749 (N_2749,N_1575,N_1977);
or U2750 (N_2750,N_2151,N_1540);
or U2751 (N_2751,N_2078,N_1542);
nand U2752 (N_2752,N_1557,N_1859);
nand U2753 (N_2753,N_1645,N_2169);
and U2754 (N_2754,N_2011,N_2048);
nor U2755 (N_2755,N_2019,N_2221);
or U2756 (N_2756,N_2201,N_1627);
or U2757 (N_2757,N_1671,N_1820);
nand U2758 (N_2758,N_1686,N_1795);
or U2759 (N_2759,N_1810,N_2014);
and U2760 (N_2760,N_1527,N_2149);
nand U2761 (N_2761,N_1505,N_1549);
or U2762 (N_2762,N_2121,N_2167);
or U2763 (N_2763,N_1927,N_1569);
nor U2764 (N_2764,N_1526,N_1628);
or U2765 (N_2765,N_1913,N_2182);
nor U2766 (N_2766,N_1536,N_2027);
nand U2767 (N_2767,N_1689,N_1896);
nand U2768 (N_2768,N_2048,N_1778);
nor U2769 (N_2769,N_1632,N_2078);
nor U2770 (N_2770,N_2199,N_1957);
nand U2771 (N_2771,N_2057,N_1517);
nand U2772 (N_2772,N_2077,N_2106);
nand U2773 (N_2773,N_1989,N_2195);
nor U2774 (N_2774,N_1757,N_2248);
and U2775 (N_2775,N_1595,N_1715);
nor U2776 (N_2776,N_1539,N_1820);
and U2777 (N_2777,N_1950,N_2197);
nor U2778 (N_2778,N_1602,N_1817);
nand U2779 (N_2779,N_1871,N_2045);
or U2780 (N_2780,N_1945,N_1564);
nor U2781 (N_2781,N_1841,N_2183);
and U2782 (N_2782,N_2211,N_1679);
nor U2783 (N_2783,N_2108,N_1962);
nor U2784 (N_2784,N_1791,N_2027);
nand U2785 (N_2785,N_1651,N_2104);
nor U2786 (N_2786,N_1688,N_1618);
nor U2787 (N_2787,N_2233,N_1639);
or U2788 (N_2788,N_1599,N_1891);
or U2789 (N_2789,N_2235,N_2170);
and U2790 (N_2790,N_1513,N_2106);
nor U2791 (N_2791,N_1705,N_1867);
nand U2792 (N_2792,N_2111,N_2188);
nand U2793 (N_2793,N_2101,N_1538);
or U2794 (N_2794,N_1904,N_1800);
nor U2795 (N_2795,N_1822,N_1656);
or U2796 (N_2796,N_1761,N_2080);
or U2797 (N_2797,N_1759,N_2032);
nand U2798 (N_2798,N_1661,N_2171);
nand U2799 (N_2799,N_1996,N_1998);
and U2800 (N_2800,N_1930,N_1601);
or U2801 (N_2801,N_1983,N_2204);
or U2802 (N_2802,N_2238,N_2220);
nand U2803 (N_2803,N_1864,N_1728);
nand U2804 (N_2804,N_2177,N_1996);
or U2805 (N_2805,N_2231,N_1709);
nor U2806 (N_2806,N_2094,N_1672);
or U2807 (N_2807,N_1513,N_2101);
nor U2808 (N_2808,N_1682,N_1805);
nand U2809 (N_2809,N_1858,N_2084);
nor U2810 (N_2810,N_2051,N_1579);
and U2811 (N_2811,N_1895,N_1768);
nor U2812 (N_2812,N_1868,N_1938);
nor U2813 (N_2813,N_1521,N_1860);
or U2814 (N_2814,N_2191,N_1834);
nand U2815 (N_2815,N_1577,N_2190);
or U2816 (N_2816,N_2244,N_1893);
nor U2817 (N_2817,N_2089,N_2005);
and U2818 (N_2818,N_1981,N_1820);
nor U2819 (N_2819,N_1989,N_1880);
and U2820 (N_2820,N_1796,N_1979);
and U2821 (N_2821,N_1851,N_1565);
nand U2822 (N_2822,N_1548,N_1949);
or U2823 (N_2823,N_2135,N_1864);
and U2824 (N_2824,N_1630,N_1900);
or U2825 (N_2825,N_1825,N_1583);
nand U2826 (N_2826,N_1852,N_1833);
or U2827 (N_2827,N_2230,N_1777);
nand U2828 (N_2828,N_1941,N_2127);
or U2829 (N_2829,N_1700,N_1632);
and U2830 (N_2830,N_1939,N_1972);
or U2831 (N_2831,N_1519,N_2134);
nand U2832 (N_2832,N_1684,N_1555);
and U2833 (N_2833,N_1910,N_1648);
and U2834 (N_2834,N_1985,N_1961);
and U2835 (N_2835,N_1509,N_1854);
or U2836 (N_2836,N_1648,N_1866);
nand U2837 (N_2837,N_1611,N_2137);
nor U2838 (N_2838,N_1818,N_1817);
xor U2839 (N_2839,N_1570,N_2179);
nand U2840 (N_2840,N_1590,N_2079);
nor U2841 (N_2841,N_1883,N_1945);
nor U2842 (N_2842,N_2223,N_1604);
xor U2843 (N_2843,N_2178,N_1634);
and U2844 (N_2844,N_2180,N_2079);
nand U2845 (N_2845,N_2016,N_1625);
nand U2846 (N_2846,N_2054,N_1500);
nand U2847 (N_2847,N_1842,N_2121);
or U2848 (N_2848,N_1984,N_1635);
nand U2849 (N_2849,N_1832,N_2192);
nand U2850 (N_2850,N_2096,N_1543);
nand U2851 (N_2851,N_2136,N_1636);
nor U2852 (N_2852,N_1738,N_2120);
xnor U2853 (N_2853,N_1527,N_1933);
nor U2854 (N_2854,N_1730,N_2208);
nand U2855 (N_2855,N_1728,N_1784);
and U2856 (N_2856,N_1945,N_1654);
or U2857 (N_2857,N_2025,N_1704);
nor U2858 (N_2858,N_2235,N_1524);
or U2859 (N_2859,N_1548,N_2020);
and U2860 (N_2860,N_1839,N_1784);
or U2861 (N_2861,N_1886,N_1527);
nor U2862 (N_2862,N_2082,N_2054);
nand U2863 (N_2863,N_1522,N_1528);
and U2864 (N_2864,N_1993,N_1741);
nand U2865 (N_2865,N_2232,N_2193);
nand U2866 (N_2866,N_1656,N_1525);
nor U2867 (N_2867,N_2177,N_2172);
nor U2868 (N_2868,N_1767,N_2004);
nand U2869 (N_2869,N_1801,N_1836);
and U2870 (N_2870,N_1953,N_2125);
nor U2871 (N_2871,N_1988,N_2052);
nor U2872 (N_2872,N_1670,N_1568);
nor U2873 (N_2873,N_1920,N_1998);
or U2874 (N_2874,N_1645,N_1600);
nand U2875 (N_2875,N_1745,N_2058);
or U2876 (N_2876,N_1613,N_1780);
and U2877 (N_2877,N_1544,N_2041);
nand U2878 (N_2878,N_2204,N_1613);
nor U2879 (N_2879,N_1723,N_2204);
and U2880 (N_2880,N_1718,N_1972);
and U2881 (N_2881,N_1970,N_2191);
nor U2882 (N_2882,N_1971,N_2210);
nor U2883 (N_2883,N_2242,N_2082);
or U2884 (N_2884,N_2243,N_1703);
nand U2885 (N_2885,N_2163,N_1513);
or U2886 (N_2886,N_2148,N_1821);
or U2887 (N_2887,N_1881,N_2043);
and U2888 (N_2888,N_2050,N_1652);
nand U2889 (N_2889,N_1637,N_1556);
nand U2890 (N_2890,N_2036,N_1797);
nand U2891 (N_2891,N_1538,N_1624);
nand U2892 (N_2892,N_1554,N_2130);
or U2893 (N_2893,N_1549,N_2120);
nor U2894 (N_2894,N_1758,N_1712);
nand U2895 (N_2895,N_1891,N_1751);
or U2896 (N_2896,N_2108,N_1677);
and U2897 (N_2897,N_1672,N_2231);
and U2898 (N_2898,N_1833,N_1696);
nand U2899 (N_2899,N_2082,N_2237);
or U2900 (N_2900,N_1814,N_2244);
nor U2901 (N_2901,N_2182,N_2189);
nor U2902 (N_2902,N_1685,N_2151);
or U2903 (N_2903,N_1549,N_1880);
nor U2904 (N_2904,N_2211,N_1575);
or U2905 (N_2905,N_1508,N_1533);
nor U2906 (N_2906,N_1917,N_1895);
or U2907 (N_2907,N_1692,N_1615);
nand U2908 (N_2908,N_2202,N_1654);
nor U2909 (N_2909,N_2072,N_1554);
and U2910 (N_2910,N_2152,N_1588);
or U2911 (N_2911,N_2199,N_1904);
nor U2912 (N_2912,N_1798,N_1665);
and U2913 (N_2913,N_2148,N_1745);
and U2914 (N_2914,N_2026,N_1678);
nor U2915 (N_2915,N_1890,N_2186);
or U2916 (N_2916,N_1887,N_1977);
nor U2917 (N_2917,N_1843,N_2225);
nand U2918 (N_2918,N_1804,N_1598);
nor U2919 (N_2919,N_1601,N_2139);
nor U2920 (N_2920,N_1680,N_1816);
or U2921 (N_2921,N_1717,N_1899);
nand U2922 (N_2922,N_1848,N_2050);
or U2923 (N_2923,N_1660,N_2054);
or U2924 (N_2924,N_1703,N_1534);
nor U2925 (N_2925,N_1916,N_2239);
nor U2926 (N_2926,N_2157,N_1621);
and U2927 (N_2927,N_1545,N_1662);
and U2928 (N_2928,N_1825,N_1795);
nor U2929 (N_2929,N_1845,N_2193);
nor U2930 (N_2930,N_1579,N_2139);
and U2931 (N_2931,N_1516,N_2241);
and U2932 (N_2932,N_1821,N_1658);
and U2933 (N_2933,N_1596,N_1621);
or U2934 (N_2934,N_2062,N_1862);
nor U2935 (N_2935,N_1680,N_1518);
or U2936 (N_2936,N_1943,N_1913);
or U2937 (N_2937,N_1569,N_2027);
nand U2938 (N_2938,N_1870,N_1848);
or U2939 (N_2939,N_1675,N_1932);
and U2940 (N_2940,N_1847,N_1596);
nand U2941 (N_2941,N_1696,N_1780);
nand U2942 (N_2942,N_1808,N_2221);
nor U2943 (N_2943,N_2177,N_1781);
or U2944 (N_2944,N_1662,N_1756);
or U2945 (N_2945,N_1967,N_2014);
and U2946 (N_2946,N_1529,N_1950);
nor U2947 (N_2947,N_1736,N_1794);
or U2948 (N_2948,N_2014,N_2048);
or U2949 (N_2949,N_1975,N_1927);
xnor U2950 (N_2950,N_1927,N_1773);
nand U2951 (N_2951,N_1896,N_1670);
nor U2952 (N_2952,N_1625,N_1706);
xor U2953 (N_2953,N_1704,N_1502);
nor U2954 (N_2954,N_1993,N_1688);
nand U2955 (N_2955,N_1599,N_1678);
nor U2956 (N_2956,N_1554,N_2241);
nand U2957 (N_2957,N_1930,N_1889);
nor U2958 (N_2958,N_1741,N_1503);
and U2959 (N_2959,N_1624,N_1865);
nand U2960 (N_2960,N_2056,N_1508);
nor U2961 (N_2961,N_1712,N_2029);
nand U2962 (N_2962,N_1825,N_1678);
nor U2963 (N_2963,N_2012,N_1555);
or U2964 (N_2964,N_1629,N_1704);
and U2965 (N_2965,N_1502,N_1692);
and U2966 (N_2966,N_1571,N_2149);
and U2967 (N_2967,N_2203,N_1726);
and U2968 (N_2968,N_1785,N_1911);
nor U2969 (N_2969,N_1727,N_2124);
nor U2970 (N_2970,N_1889,N_1616);
or U2971 (N_2971,N_1967,N_2127);
or U2972 (N_2972,N_1768,N_2175);
nand U2973 (N_2973,N_1975,N_1589);
nand U2974 (N_2974,N_1937,N_2078);
or U2975 (N_2975,N_1583,N_1726);
or U2976 (N_2976,N_1826,N_1626);
or U2977 (N_2977,N_1770,N_1722);
and U2978 (N_2978,N_2167,N_2075);
nor U2979 (N_2979,N_2036,N_1639);
and U2980 (N_2980,N_1638,N_2028);
or U2981 (N_2981,N_1791,N_1619);
and U2982 (N_2982,N_2116,N_2241);
or U2983 (N_2983,N_2239,N_1948);
nor U2984 (N_2984,N_1991,N_1581);
and U2985 (N_2985,N_1690,N_2026);
or U2986 (N_2986,N_1672,N_1522);
nand U2987 (N_2987,N_1734,N_1941);
and U2988 (N_2988,N_1700,N_2110);
nand U2989 (N_2989,N_1536,N_1995);
nor U2990 (N_2990,N_2077,N_1813);
nor U2991 (N_2991,N_2240,N_1750);
and U2992 (N_2992,N_1923,N_1983);
or U2993 (N_2993,N_1874,N_2085);
and U2994 (N_2994,N_2133,N_1575);
nand U2995 (N_2995,N_2149,N_2238);
nor U2996 (N_2996,N_1726,N_1957);
and U2997 (N_2997,N_2150,N_1700);
nand U2998 (N_2998,N_1745,N_1652);
and U2999 (N_2999,N_1760,N_1837);
nand UO_0 (O_0,N_2577,N_2771);
nor UO_1 (O_1,N_2510,N_2744);
or UO_2 (O_2,N_2746,N_2343);
and UO_3 (O_3,N_2733,N_2415);
and UO_4 (O_4,N_2785,N_2992);
nand UO_5 (O_5,N_2742,N_2501);
nor UO_6 (O_6,N_2544,N_2970);
nand UO_7 (O_7,N_2298,N_2838);
and UO_8 (O_8,N_2592,N_2553);
nand UO_9 (O_9,N_2874,N_2349);
xor UO_10 (O_10,N_2885,N_2630);
nand UO_11 (O_11,N_2969,N_2810);
or UO_12 (O_12,N_2814,N_2853);
nor UO_13 (O_13,N_2937,N_2831);
nor UO_14 (O_14,N_2319,N_2791);
or UO_15 (O_15,N_2845,N_2911);
and UO_16 (O_16,N_2364,N_2328);
nor UO_17 (O_17,N_2753,N_2805);
and UO_18 (O_18,N_2432,N_2763);
nand UO_19 (O_19,N_2420,N_2910);
nand UO_20 (O_20,N_2569,N_2350);
nand UO_21 (O_21,N_2401,N_2703);
or UO_22 (O_22,N_2363,N_2826);
and UO_23 (O_23,N_2954,N_2545);
or UO_24 (O_24,N_2323,N_2884);
or UO_25 (O_25,N_2800,N_2387);
and UO_26 (O_26,N_2898,N_2311);
nand UO_27 (O_27,N_2927,N_2270);
or UO_28 (O_28,N_2920,N_2715);
and UO_29 (O_29,N_2416,N_2508);
nand UO_30 (O_30,N_2414,N_2440);
nand UO_31 (O_31,N_2978,N_2935);
and UO_32 (O_32,N_2903,N_2533);
or UO_33 (O_33,N_2317,N_2716);
and UO_34 (O_34,N_2655,N_2605);
nor UO_35 (O_35,N_2465,N_2535);
nand UO_36 (O_36,N_2264,N_2852);
nor UO_37 (O_37,N_2642,N_2691);
and UO_38 (O_38,N_2579,N_2489);
and UO_39 (O_39,N_2601,N_2855);
nor UO_40 (O_40,N_2513,N_2483);
nand UO_41 (O_41,N_2581,N_2811);
nor UO_42 (O_42,N_2770,N_2891);
or UO_43 (O_43,N_2447,N_2548);
or UO_44 (O_44,N_2677,N_2478);
nand UO_45 (O_45,N_2833,N_2723);
nand UO_46 (O_46,N_2308,N_2375);
and UO_47 (O_47,N_2384,N_2665);
or UO_48 (O_48,N_2976,N_2463);
and UO_49 (O_49,N_2768,N_2769);
nand UO_50 (O_50,N_2933,N_2547);
nor UO_51 (O_51,N_2580,N_2276);
nand UO_52 (O_52,N_2616,N_2895);
or UO_53 (O_53,N_2406,N_2296);
nand UO_54 (O_54,N_2473,N_2450);
xnor UO_55 (O_55,N_2321,N_2916);
and UO_56 (O_56,N_2486,N_2542);
nand UO_57 (O_57,N_2585,N_2452);
or UO_58 (O_58,N_2290,N_2528);
nor UO_59 (O_59,N_2449,N_2958);
nand UO_60 (O_60,N_2748,N_2731);
and UO_61 (O_61,N_2823,N_2552);
nand UO_62 (O_62,N_2775,N_2436);
nand UO_63 (O_63,N_2285,N_2736);
or UO_64 (O_64,N_2975,N_2640);
nor UO_65 (O_65,N_2869,N_2890);
and UO_66 (O_66,N_2951,N_2383);
and UO_67 (O_67,N_2946,N_2610);
nand UO_68 (O_68,N_2558,N_2626);
nand UO_69 (O_69,N_2362,N_2372);
or UO_70 (O_70,N_2477,N_2602);
nand UO_71 (O_71,N_2310,N_2507);
or UO_72 (O_72,N_2258,N_2688);
xor UO_73 (O_73,N_2638,N_2687);
nand UO_74 (O_74,N_2690,N_2980);
nand UO_75 (O_75,N_2609,N_2386);
nand UO_76 (O_76,N_2502,N_2983);
nor UO_77 (O_77,N_2998,N_2947);
or UO_78 (O_78,N_2278,N_2720);
and UO_79 (O_79,N_2265,N_2431);
nor UO_80 (O_80,N_2861,N_2423);
or UO_81 (O_81,N_2661,N_2701);
nor UO_82 (O_82,N_2700,N_2713);
nand UO_83 (O_83,N_2391,N_2302);
and UO_84 (O_84,N_2675,N_2588);
nor UO_85 (O_85,N_2491,N_2318);
and UO_86 (O_86,N_2427,N_2471);
and UO_87 (O_87,N_2400,N_2624);
or UO_88 (O_88,N_2422,N_2520);
nand UO_89 (O_89,N_2287,N_2667);
and UO_90 (O_90,N_2411,N_2370);
nand UO_91 (O_91,N_2267,N_2777);
and UO_92 (O_92,N_2525,N_2815);
and UO_93 (O_93,N_2405,N_2901);
nand UO_94 (O_94,N_2989,N_2348);
nor UO_95 (O_95,N_2851,N_2803);
nand UO_96 (O_96,N_2864,N_2281);
nand UO_97 (O_97,N_2797,N_2841);
nand UO_98 (O_98,N_2353,N_2576);
nor UO_99 (O_99,N_2309,N_2495);
or UO_100 (O_100,N_2698,N_2977);
nor UO_101 (O_101,N_2346,N_2556);
or UO_102 (O_102,N_2973,N_2286);
nand UO_103 (O_103,N_2407,N_2606);
and UO_104 (O_104,N_2627,N_2257);
and UO_105 (O_105,N_2398,N_2537);
and UO_106 (O_106,N_2480,N_2284);
and UO_107 (O_107,N_2360,N_2430);
nor UO_108 (O_108,N_2892,N_2275);
or UO_109 (O_109,N_2737,N_2526);
and UO_110 (O_110,N_2629,N_2435);
and UO_111 (O_111,N_2336,N_2439);
nor UO_112 (O_112,N_2648,N_2789);
nor UO_113 (O_113,N_2717,N_2283);
and UO_114 (O_114,N_2550,N_2358);
nand UO_115 (O_115,N_2949,N_2484);
nor UO_116 (O_116,N_2359,N_2918);
or UO_117 (O_117,N_2830,N_2551);
nor UO_118 (O_118,N_2497,N_2679);
and UO_119 (O_119,N_2458,N_2297);
or UO_120 (O_120,N_2279,N_2390);
nor UO_121 (O_121,N_2936,N_2639);
nand UO_122 (O_122,N_2333,N_2881);
nand UO_123 (O_123,N_2517,N_2725);
or UO_124 (O_124,N_2646,N_2836);
and UO_125 (O_125,N_2344,N_2664);
nand UO_126 (O_126,N_2574,N_2437);
nor UO_127 (O_127,N_2514,N_2554);
or UO_128 (O_128,N_2566,N_2924);
nor UO_129 (O_129,N_2320,N_2837);
nor UO_130 (O_130,N_2559,N_2740);
nor UO_131 (O_131,N_2905,N_2603);
or UO_132 (O_132,N_2809,N_2865);
nor UO_133 (O_133,N_2518,N_2650);
or UO_134 (O_134,N_2985,N_2995);
or UO_135 (O_135,N_2598,N_2674);
or UO_136 (O_136,N_2780,N_2338);
nor UO_137 (O_137,N_2636,N_2381);
and UO_138 (O_138,N_2291,N_2329);
nor UO_139 (O_139,N_2813,N_2324);
nor UO_140 (O_140,N_2994,N_2693);
or UO_141 (O_141,N_2676,N_2850);
nor UO_142 (O_142,N_2956,N_2568);
nand UO_143 (O_143,N_2354,N_2705);
nor UO_144 (O_144,N_2967,N_2858);
and UO_145 (O_145,N_2428,N_2482);
and UO_146 (O_146,N_2261,N_2498);
nor UO_147 (O_147,N_2256,N_2645);
nor UO_148 (O_148,N_2668,N_2825);
nand UO_149 (O_149,N_2560,N_2929);
nor UO_150 (O_150,N_2322,N_2678);
nand UO_151 (O_151,N_2351,N_2896);
nand UO_152 (O_152,N_2382,N_2527);
nor UO_153 (O_153,N_2945,N_2392);
and UO_154 (O_154,N_2345,N_2751);
nor UO_155 (O_155,N_2883,N_2848);
or UO_156 (O_156,N_2255,N_2806);
nand UO_157 (O_157,N_2888,N_2326);
nor UO_158 (O_158,N_2368,N_2681);
and UO_159 (O_159,N_2567,N_2963);
and UO_160 (O_160,N_2824,N_2570);
xor UO_161 (O_161,N_2614,N_2355);
and UO_162 (O_162,N_2893,N_2413);
or UO_163 (O_163,N_2369,N_2472);
nand UO_164 (O_164,N_2294,N_2718);
nor UO_165 (O_165,N_2334,N_2419);
or UO_166 (O_166,N_2378,N_2799);
or UO_167 (O_167,N_2794,N_2860);
nand UO_168 (O_168,N_2448,N_2738);
nor UO_169 (O_169,N_2882,N_2410);
nor UO_170 (O_170,N_2672,N_2897);
or UO_171 (O_171,N_2583,N_2979);
and UO_172 (O_172,N_2961,N_2925);
nor UO_173 (O_173,N_2695,N_2599);
nor UO_174 (O_174,N_2573,N_2663);
nor UO_175 (O_175,N_2408,N_2889);
and UO_176 (O_176,N_2727,N_2300);
nor UO_177 (O_177,N_2702,N_2371);
nand UO_178 (O_178,N_2494,N_2361);
and UO_179 (O_179,N_2704,N_2503);
or UO_180 (O_180,N_2524,N_2952);
xor UO_181 (O_181,N_2656,N_2443);
nand UO_182 (O_182,N_2834,N_2451);
or UO_183 (O_183,N_2259,N_2812);
nor UO_184 (O_184,N_2619,N_2591);
and UO_185 (O_185,N_2453,N_2615);
nand UO_186 (O_186,N_2397,N_2254);
or UO_187 (O_187,N_2557,N_2536);
nand UO_188 (O_188,N_2948,N_2766);
nand UO_189 (O_189,N_2714,N_2572);
or UO_190 (O_190,N_2467,N_2900);
and UO_191 (O_191,N_2671,N_2404);
nor UO_192 (O_192,N_2752,N_2697);
and UO_193 (O_193,N_2662,N_2365);
nand UO_194 (O_194,N_2442,N_2993);
and UO_195 (O_195,N_2446,N_2863);
nor UO_196 (O_196,N_2335,N_2367);
or UO_197 (O_197,N_2425,N_2521);
and UO_198 (O_198,N_2692,N_2496);
and UO_199 (O_199,N_2263,N_2641);
and UO_200 (O_200,N_2456,N_2561);
and UO_201 (O_201,N_2643,N_2538);
or UO_202 (O_202,N_2313,N_2539);
nand UO_203 (O_203,N_2868,N_2277);
nand UO_204 (O_204,N_2280,N_2402);
and UO_205 (O_205,N_2866,N_2352);
nand UO_206 (O_206,N_2906,N_2801);
or UO_207 (O_207,N_2586,N_2699);
nand UO_208 (O_208,N_2908,N_2827);
or UO_209 (O_209,N_2620,N_2464);
nand UO_210 (O_210,N_2342,N_2325);
nand UO_211 (O_211,N_2578,N_2926);
nand UO_212 (O_212,N_2461,N_2613);
or UO_213 (O_213,N_2760,N_2493);
or UO_214 (O_214,N_2475,N_2628);
and UO_215 (O_215,N_2622,N_2781);
nor UO_216 (O_216,N_2694,N_2870);
and UO_217 (O_217,N_2783,N_2563);
or UO_218 (O_218,N_2974,N_2798);
or UO_219 (O_219,N_2385,N_2840);
or UO_220 (O_220,N_2735,N_2996);
or UO_221 (O_221,N_2519,N_2393);
nor UO_222 (O_222,N_2757,N_2767);
or UO_223 (O_223,N_2680,N_2459);
or UO_224 (O_224,N_2859,N_2597);
or UO_225 (O_225,N_2894,N_2304);
nor UO_226 (O_226,N_2730,N_2575);
or UO_227 (O_227,N_2922,N_2394);
nand UO_228 (O_228,N_2492,N_2873);
and UO_229 (O_229,N_2634,N_2939);
and UO_230 (O_230,N_2773,N_2932);
and UO_231 (O_231,N_2269,N_2990);
nand UO_232 (O_232,N_2779,N_2741);
nand UO_233 (O_233,N_2772,N_2919);
nand UO_234 (O_234,N_2709,N_2843);
nand UO_235 (O_235,N_2724,N_2658);
nor UO_236 (O_236,N_2608,N_2747);
nor UO_237 (O_237,N_2584,N_2631);
nor UO_238 (O_238,N_2540,N_2942);
and UO_239 (O_239,N_2856,N_2657);
and UO_240 (O_240,N_2669,N_2988);
nor UO_241 (O_241,N_2871,N_2555);
nor UO_242 (O_242,N_2712,N_2562);
or UO_243 (O_243,N_2637,N_2396);
or UO_244 (O_244,N_2531,N_2706);
nand UO_245 (O_245,N_2880,N_2957);
and UO_246 (O_246,N_2293,N_2377);
and UO_247 (O_247,N_2541,N_2262);
or UO_248 (O_248,N_2822,N_2917);
or UO_249 (O_249,N_2653,N_2506);
nor UO_250 (O_250,N_2315,N_2647);
and UO_251 (O_251,N_2987,N_2786);
nor UO_252 (O_252,N_2522,N_2388);
or UO_253 (O_253,N_2959,N_2485);
nand UO_254 (O_254,N_2962,N_2749);
nor UO_255 (O_255,N_2707,N_2499);
nand UO_256 (O_256,N_2964,N_2689);
nand UO_257 (O_257,N_2250,N_2632);
and UO_258 (O_258,N_2955,N_2644);
nor UO_259 (O_259,N_2389,N_2332);
or UO_260 (O_260,N_2808,N_2844);
nor UO_261 (O_261,N_2412,N_2739);
nor UO_262 (O_262,N_2593,N_2943);
or UO_263 (O_263,N_2380,N_2792);
or UO_264 (O_264,N_2316,N_2950);
and UO_265 (O_265,N_2804,N_2305);
or UO_266 (O_266,N_2921,N_2877);
or UO_267 (O_267,N_2726,N_2515);
nand UO_268 (O_268,N_2403,N_2457);
nor UO_269 (O_269,N_2571,N_2816);
or UO_270 (O_270,N_2710,N_2312);
or UO_271 (O_271,N_2968,N_2612);
or UO_272 (O_272,N_2682,N_2374);
and UO_273 (O_273,N_2337,N_2913);
and UO_274 (O_274,N_2604,N_2886);
nor UO_275 (O_275,N_2842,N_2625);
nor UO_276 (O_276,N_2887,N_2429);
or UO_277 (O_277,N_2595,N_2282);
nor UO_278 (O_278,N_2529,N_2821);
or UO_279 (O_279,N_2788,N_2854);
nand UO_280 (O_280,N_2732,N_2589);
nand UO_281 (O_281,N_2366,N_2914);
nand UO_282 (O_282,N_2711,N_2418);
nand UO_283 (O_283,N_2399,N_2373);
nand UO_284 (O_284,N_2481,N_2288);
nand UO_285 (O_285,N_2633,N_2594);
or UO_286 (O_286,N_2982,N_2462);
nor UO_287 (O_287,N_2899,N_2981);
nor UO_288 (O_288,N_2764,N_2934);
nand UO_289 (O_289,N_2596,N_2849);
or UO_290 (O_290,N_2424,N_2847);
nand UO_291 (O_291,N_2379,N_2445);
nor UO_292 (O_292,N_2796,N_2649);
or UO_293 (O_293,N_2356,N_2938);
or UO_294 (O_294,N_2971,N_2829);
nand UO_295 (O_295,N_2879,N_2722);
nand UO_296 (O_296,N_2728,N_2607);
or UO_297 (O_297,N_2546,N_2516);
nor UO_298 (O_298,N_2512,N_2765);
and UO_299 (O_299,N_2953,N_2395);
nand UO_300 (O_300,N_2966,N_2817);
or UO_301 (O_301,N_2260,N_2330);
or UO_302 (O_302,N_2582,N_2509);
nor UO_303 (O_303,N_2673,N_2434);
nor UO_304 (O_304,N_2268,N_2292);
and UO_305 (O_305,N_2454,N_2876);
nor UO_306 (O_306,N_2778,N_2654);
or UO_307 (O_307,N_2339,N_2565);
and UO_308 (O_308,N_2729,N_2754);
nor UO_309 (O_309,N_2835,N_2683);
or UO_310 (O_310,N_2600,N_2867);
or UO_311 (O_311,N_2818,N_2266);
and UO_312 (O_312,N_2306,N_2659);
or UO_313 (O_313,N_2944,N_2660);
or UO_314 (O_314,N_2357,N_2758);
nor UO_315 (O_315,N_2273,N_2904);
or UO_316 (O_316,N_2734,N_2543);
and UO_317 (O_317,N_2928,N_2252);
or UO_318 (O_318,N_2564,N_2251);
nand UO_319 (O_319,N_2819,N_2666);
nor UO_320 (O_320,N_2468,N_2490);
nand UO_321 (O_321,N_2802,N_2902);
nand UO_322 (O_322,N_2417,N_2618);
or UO_323 (O_323,N_2761,N_2523);
or UO_324 (O_324,N_2303,N_2719);
nor UO_325 (O_325,N_2685,N_2421);
or UO_326 (O_326,N_2590,N_2931);
or UO_327 (O_327,N_2505,N_2530);
and UO_328 (O_328,N_2875,N_2941);
and UO_329 (O_329,N_2455,N_2479);
or UO_330 (O_330,N_2708,N_2376);
and UO_331 (O_331,N_2487,N_2960);
or UO_332 (O_332,N_2915,N_2623);
and UO_333 (O_333,N_2272,N_2474);
and UO_334 (O_334,N_2271,N_2828);
nor UO_335 (O_335,N_2549,N_2907);
nor UO_336 (O_336,N_2433,N_2846);
xnor UO_337 (O_337,N_2635,N_2488);
nor UO_338 (O_338,N_2444,N_2972);
or UO_339 (O_339,N_2438,N_2532);
nand UO_340 (O_340,N_2469,N_2984);
and UO_341 (O_341,N_2756,N_2940);
nor UO_342 (O_342,N_2466,N_2331);
and UO_343 (O_343,N_2787,N_2999);
and UO_344 (O_344,N_2930,N_2651);
nor UO_345 (O_345,N_2909,N_2670);
and UO_346 (O_346,N_2686,N_2289);
and UO_347 (O_347,N_2986,N_2500);
nor UO_348 (O_348,N_2274,N_2782);
and UO_349 (O_349,N_2460,N_2684);
and UO_350 (O_350,N_2743,N_2820);
nand UO_351 (O_351,N_2426,N_2878);
and UO_352 (O_352,N_2511,N_2750);
or UO_353 (O_353,N_2872,N_2587);
nor UO_354 (O_354,N_2441,N_2295);
or UO_355 (O_355,N_2759,N_2652);
nand UO_356 (O_356,N_2862,N_2307);
or UO_357 (O_357,N_2832,N_2340);
or UO_358 (O_358,N_2696,N_2253);
nand UO_359 (O_359,N_2795,N_2476);
and UO_360 (O_360,N_2347,N_2470);
nand UO_361 (O_361,N_2301,N_2621);
nor UO_362 (O_362,N_2504,N_2762);
nor UO_363 (O_363,N_2721,N_2807);
or UO_364 (O_364,N_2965,N_2774);
nand UO_365 (O_365,N_2991,N_2409);
and UO_366 (O_366,N_2617,N_2790);
or UO_367 (O_367,N_2784,N_2776);
or UO_368 (O_368,N_2299,N_2857);
and UO_369 (O_369,N_2912,N_2327);
nor UO_370 (O_370,N_2755,N_2997);
or UO_371 (O_371,N_2839,N_2341);
or UO_372 (O_372,N_2314,N_2745);
nor UO_373 (O_373,N_2793,N_2923);
nand UO_374 (O_374,N_2611,N_2534);
nor UO_375 (O_375,N_2382,N_2625);
and UO_376 (O_376,N_2797,N_2441);
and UO_377 (O_377,N_2692,N_2495);
nand UO_378 (O_378,N_2326,N_2517);
nor UO_379 (O_379,N_2383,N_2632);
or UO_380 (O_380,N_2804,N_2847);
and UO_381 (O_381,N_2565,N_2690);
or UO_382 (O_382,N_2424,N_2679);
and UO_383 (O_383,N_2299,N_2608);
or UO_384 (O_384,N_2741,N_2725);
nor UO_385 (O_385,N_2321,N_2283);
nor UO_386 (O_386,N_2847,N_2869);
nor UO_387 (O_387,N_2780,N_2731);
or UO_388 (O_388,N_2879,N_2306);
and UO_389 (O_389,N_2290,N_2355);
or UO_390 (O_390,N_2377,N_2889);
and UO_391 (O_391,N_2972,N_2279);
nand UO_392 (O_392,N_2319,N_2494);
nand UO_393 (O_393,N_2981,N_2813);
nor UO_394 (O_394,N_2633,N_2913);
or UO_395 (O_395,N_2834,N_2297);
or UO_396 (O_396,N_2836,N_2471);
nand UO_397 (O_397,N_2493,N_2388);
and UO_398 (O_398,N_2699,N_2290);
nand UO_399 (O_399,N_2842,N_2470);
or UO_400 (O_400,N_2535,N_2358);
or UO_401 (O_401,N_2349,N_2512);
and UO_402 (O_402,N_2445,N_2267);
or UO_403 (O_403,N_2462,N_2594);
nor UO_404 (O_404,N_2912,N_2442);
or UO_405 (O_405,N_2264,N_2509);
and UO_406 (O_406,N_2408,N_2811);
or UO_407 (O_407,N_2588,N_2658);
nor UO_408 (O_408,N_2280,N_2722);
nor UO_409 (O_409,N_2974,N_2559);
or UO_410 (O_410,N_2980,N_2917);
or UO_411 (O_411,N_2990,N_2933);
or UO_412 (O_412,N_2510,N_2546);
nor UO_413 (O_413,N_2574,N_2568);
nor UO_414 (O_414,N_2933,N_2342);
and UO_415 (O_415,N_2673,N_2265);
and UO_416 (O_416,N_2280,N_2567);
nand UO_417 (O_417,N_2993,N_2374);
and UO_418 (O_418,N_2261,N_2251);
nand UO_419 (O_419,N_2918,N_2632);
and UO_420 (O_420,N_2627,N_2633);
and UO_421 (O_421,N_2690,N_2879);
or UO_422 (O_422,N_2596,N_2985);
or UO_423 (O_423,N_2348,N_2868);
nor UO_424 (O_424,N_2549,N_2288);
nand UO_425 (O_425,N_2445,N_2303);
nor UO_426 (O_426,N_2542,N_2942);
nor UO_427 (O_427,N_2993,N_2437);
nor UO_428 (O_428,N_2398,N_2419);
nor UO_429 (O_429,N_2645,N_2672);
nand UO_430 (O_430,N_2489,N_2283);
nor UO_431 (O_431,N_2944,N_2409);
nor UO_432 (O_432,N_2347,N_2676);
and UO_433 (O_433,N_2687,N_2904);
and UO_434 (O_434,N_2386,N_2987);
nor UO_435 (O_435,N_2679,N_2454);
and UO_436 (O_436,N_2746,N_2325);
and UO_437 (O_437,N_2443,N_2469);
or UO_438 (O_438,N_2335,N_2253);
nor UO_439 (O_439,N_2618,N_2341);
or UO_440 (O_440,N_2381,N_2449);
and UO_441 (O_441,N_2459,N_2266);
and UO_442 (O_442,N_2825,N_2457);
or UO_443 (O_443,N_2473,N_2992);
and UO_444 (O_444,N_2927,N_2550);
or UO_445 (O_445,N_2534,N_2257);
nor UO_446 (O_446,N_2964,N_2893);
and UO_447 (O_447,N_2568,N_2299);
nor UO_448 (O_448,N_2576,N_2421);
or UO_449 (O_449,N_2304,N_2755);
nand UO_450 (O_450,N_2468,N_2519);
nor UO_451 (O_451,N_2947,N_2446);
and UO_452 (O_452,N_2642,N_2707);
or UO_453 (O_453,N_2557,N_2508);
or UO_454 (O_454,N_2583,N_2878);
nor UO_455 (O_455,N_2418,N_2835);
nand UO_456 (O_456,N_2905,N_2813);
nand UO_457 (O_457,N_2526,N_2596);
nand UO_458 (O_458,N_2310,N_2716);
or UO_459 (O_459,N_2973,N_2487);
nand UO_460 (O_460,N_2823,N_2541);
nand UO_461 (O_461,N_2387,N_2875);
and UO_462 (O_462,N_2510,N_2826);
nand UO_463 (O_463,N_2928,N_2711);
nor UO_464 (O_464,N_2629,N_2990);
and UO_465 (O_465,N_2657,N_2859);
and UO_466 (O_466,N_2353,N_2776);
nor UO_467 (O_467,N_2587,N_2312);
nand UO_468 (O_468,N_2463,N_2427);
or UO_469 (O_469,N_2669,N_2283);
nor UO_470 (O_470,N_2808,N_2609);
nand UO_471 (O_471,N_2604,N_2483);
nand UO_472 (O_472,N_2856,N_2470);
nor UO_473 (O_473,N_2888,N_2663);
nand UO_474 (O_474,N_2817,N_2880);
and UO_475 (O_475,N_2308,N_2962);
or UO_476 (O_476,N_2675,N_2799);
nor UO_477 (O_477,N_2995,N_2548);
nor UO_478 (O_478,N_2806,N_2418);
and UO_479 (O_479,N_2597,N_2255);
or UO_480 (O_480,N_2589,N_2502);
nand UO_481 (O_481,N_2458,N_2442);
nand UO_482 (O_482,N_2465,N_2905);
nor UO_483 (O_483,N_2408,N_2887);
nand UO_484 (O_484,N_2739,N_2974);
or UO_485 (O_485,N_2906,N_2259);
or UO_486 (O_486,N_2924,N_2542);
nand UO_487 (O_487,N_2517,N_2308);
nor UO_488 (O_488,N_2332,N_2998);
or UO_489 (O_489,N_2966,N_2969);
nand UO_490 (O_490,N_2663,N_2850);
nor UO_491 (O_491,N_2260,N_2455);
nor UO_492 (O_492,N_2435,N_2446);
and UO_493 (O_493,N_2398,N_2895);
or UO_494 (O_494,N_2466,N_2341);
nor UO_495 (O_495,N_2452,N_2450);
or UO_496 (O_496,N_2721,N_2327);
and UO_497 (O_497,N_2870,N_2613);
nor UO_498 (O_498,N_2911,N_2616);
or UO_499 (O_499,N_2260,N_2498);
endmodule