module basic_500_3000_500_3_levels_1xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nor U0 (N_0,In_142,In_99);
nor U1 (N_1,In_170,In_250);
and U2 (N_2,In_471,In_267);
nand U3 (N_3,In_102,In_1);
nor U4 (N_4,In_421,In_101);
nand U5 (N_5,In_371,In_254);
or U6 (N_6,In_374,In_401);
nor U7 (N_7,In_482,In_382);
nor U8 (N_8,In_78,In_350);
or U9 (N_9,In_289,In_18);
nand U10 (N_10,In_474,In_329);
nor U11 (N_11,In_36,In_288);
xor U12 (N_12,In_227,In_182);
nor U13 (N_13,In_187,In_37);
and U14 (N_14,In_148,In_2);
and U15 (N_15,In_320,In_273);
nor U16 (N_16,In_195,In_15);
or U17 (N_17,In_342,In_104);
nand U18 (N_18,In_33,In_292);
nand U19 (N_19,In_287,In_498);
nand U20 (N_20,In_476,In_439);
or U21 (N_21,In_262,In_236);
and U22 (N_22,In_135,In_461);
and U23 (N_23,In_144,In_352);
or U24 (N_24,In_149,In_68);
xnor U25 (N_25,In_456,In_167);
nor U26 (N_26,In_402,In_319);
nand U27 (N_27,In_107,In_245);
nor U28 (N_28,In_226,In_470);
nor U29 (N_29,In_260,In_274);
nand U30 (N_30,In_72,In_223);
or U31 (N_31,In_432,In_87);
nor U32 (N_32,In_466,In_190);
and U33 (N_33,In_120,In_263);
or U34 (N_34,In_185,In_345);
or U35 (N_35,In_290,In_192);
nor U36 (N_36,In_191,In_30);
nand U37 (N_37,In_307,In_283);
and U38 (N_38,In_302,In_141);
and U39 (N_39,In_242,In_451);
or U40 (N_40,In_11,In_477);
or U41 (N_41,In_340,In_113);
nor U42 (N_42,In_272,In_309);
nor U43 (N_43,In_394,In_325);
or U44 (N_44,In_48,In_128);
or U45 (N_45,In_480,In_330);
or U46 (N_46,In_259,In_431);
and U47 (N_47,In_24,In_317);
nor U48 (N_48,In_489,In_308);
nand U49 (N_49,In_447,In_479);
nand U50 (N_50,In_95,In_21);
or U51 (N_51,In_275,In_4);
or U52 (N_52,In_80,In_140);
and U53 (N_53,In_487,In_207);
nand U54 (N_54,In_218,In_429);
nand U55 (N_55,In_314,In_70);
nand U56 (N_56,In_433,In_111);
or U57 (N_57,In_246,In_184);
and U58 (N_58,In_279,In_249);
nor U59 (N_59,In_494,In_115);
nand U60 (N_60,In_328,In_383);
and U61 (N_61,In_305,In_150);
nand U62 (N_62,In_79,In_270);
nor U63 (N_63,In_388,In_166);
nand U64 (N_64,In_372,In_280);
and U65 (N_65,In_261,In_343);
nand U66 (N_66,In_493,In_415);
nor U67 (N_67,In_327,In_34);
nand U68 (N_68,In_248,In_392);
nand U69 (N_69,In_209,In_14);
or U70 (N_70,In_16,In_252);
and U71 (N_71,In_357,In_335);
nor U72 (N_72,In_136,In_106);
or U73 (N_73,In_51,In_119);
or U74 (N_74,In_285,In_12);
and U75 (N_75,In_497,In_444);
nand U76 (N_76,In_247,In_442);
or U77 (N_77,In_495,In_363);
or U78 (N_78,In_31,In_423);
nand U79 (N_79,In_88,In_424);
or U80 (N_80,In_397,In_331);
or U81 (N_81,In_194,In_169);
nand U82 (N_82,In_74,In_198);
or U83 (N_83,In_349,In_295);
nor U84 (N_84,In_436,In_411);
nand U85 (N_85,In_9,In_180);
nor U86 (N_86,In_323,In_449);
or U87 (N_87,In_417,In_450);
nor U88 (N_88,In_97,In_348);
or U89 (N_89,In_244,In_90);
or U90 (N_90,In_219,In_117);
nand U91 (N_91,In_174,In_59);
and U92 (N_92,In_19,In_364);
nor U93 (N_93,In_469,In_346);
nor U94 (N_94,In_324,In_358);
nand U95 (N_95,In_351,In_265);
and U96 (N_96,In_412,In_475);
and U97 (N_97,In_86,In_269);
or U98 (N_98,In_105,In_176);
nand U99 (N_99,In_64,In_304);
nand U100 (N_100,In_306,In_56);
nor U101 (N_101,In_293,In_10);
or U102 (N_102,In_386,In_77);
nand U103 (N_103,In_134,In_300);
nor U104 (N_104,In_229,In_213);
nor U105 (N_105,In_332,In_116);
and U106 (N_106,In_385,In_297);
or U107 (N_107,In_478,In_443);
nor U108 (N_108,In_264,In_152);
nand U109 (N_109,In_301,In_376);
nor U110 (N_110,In_132,In_276);
nor U111 (N_111,In_445,In_281);
nor U112 (N_112,In_256,In_438);
and U113 (N_113,In_109,In_422);
nand U114 (N_114,In_410,In_112);
nor U115 (N_115,In_98,In_139);
and U116 (N_116,In_404,In_370);
nor U117 (N_117,In_100,In_294);
nand U118 (N_118,In_123,In_403);
and U119 (N_119,In_7,In_131);
or U120 (N_120,In_147,In_125);
nand U121 (N_121,In_156,In_181);
and U122 (N_122,In_454,In_379);
nand U123 (N_123,In_233,In_409);
nand U124 (N_124,In_228,In_171);
and U125 (N_125,In_235,In_153);
nor U126 (N_126,In_464,In_318);
nor U127 (N_127,In_414,In_124);
or U128 (N_128,In_76,In_239);
and U129 (N_129,In_183,In_310);
or U130 (N_130,In_230,In_71);
or U131 (N_131,In_237,In_165);
or U132 (N_132,In_393,In_365);
nand U133 (N_133,In_362,In_481);
nor U134 (N_134,In_47,In_108);
nand U135 (N_135,In_130,In_483);
nor U136 (N_136,In_408,In_55);
nand U137 (N_137,In_419,In_61);
nand U138 (N_138,In_238,In_367);
and U139 (N_139,In_338,In_425);
and U140 (N_140,In_485,In_57);
nand U141 (N_141,In_40,In_222);
and U142 (N_142,In_395,In_368);
or U143 (N_143,In_315,In_8);
nor U144 (N_144,In_463,In_66);
nand U145 (N_145,In_126,In_496);
nand U146 (N_146,In_339,In_472);
nor U147 (N_147,In_312,In_303);
nand U148 (N_148,In_60,In_143);
nor U149 (N_149,In_396,In_284);
and U150 (N_150,In_29,In_197);
and U151 (N_151,In_175,In_225);
and U152 (N_152,In_65,In_93);
nand U153 (N_153,In_32,In_155);
nand U154 (N_154,In_154,In_62);
nor U155 (N_155,In_89,In_369);
nor U156 (N_156,In_234,In_178);
nor U157 (N_157,In_313,In_221);
or U158 (N_158,In_216,In_266);
or U159 (N_159,In_398,In_435);
nand U160 (N_160,In_428,In_486);
and U161 (N_161,In_85,In_202);
or U162 (N_162,In_5,In_291);
and U163 (N_163,In_361,In_241);
nand U164 (N_164,In_427,In_286);
nand U165 (N_165,In_311,In_458);
and U166 (N_166,In_441,In_416);
nor U167 (N_167,In_224,In_46);
and U168 (N_168,In_214,In_53);
and U169 (N_169,In_26,In_118);
nor U170 (N_170,In_211,In_437);
or U171 (N_171,In_138,In_163);
and U172 (N_172,In_54,In_296);
and U173 (N_173,In_366,In_44);
nor U174 (N_174,In_91,In_67);
and U175 (N_175,In_200,In_232);
nand U176 (N_176,In_258,In_137);
and U177 (N_177,In_282,In_321);
nand U178 (N_178,In_49,In_298);
or U179 (N_179,In_173,In_354);
and U180 (N_180,In_52,In_28);
nor U181 (N_181,In_359,In_206);
nor U182 (N_182,In_159,In_499);
or U183 (N_183,In_434,In_179);
nand U184 (N_184,In_189,In_83);
nand U185 (N_185,In_94,In_161);
nor U186 (N_186,In_199,In_491);
or U187 (N_187,In_448,In_217);
nor U188 (N_188,In_378,In_42);
nand U189 (N_189,In_243,In_459);
nand U190 (N_190,In_387,In_23);
nand U191 (N_191,In_344,In_84);
or U192 (N_192,In_460,In_271);
nor U193 (N_193,In_407,In_240);
and U194 (N_194,In_122,In_400);
nor U195 (N_195,In_103,In_333);
nand U196 (N_196,In_220,In_377);
and U197 (N_197,In_251,In_133);
or U198 (N_198,In_129,In_356);
nand U199 (N_199,In_114,In_334);
nor U200 (N_200,In_467,In_164);
and U201 (N_201,In_452,In_188);
nor U202 (N_202,In_418,In_492);
and U203 (N_203,In_462,In_446);
nor U204 (N_204,In_186,In_473);
nand U205 (N_205,In_210,In_203);
nor U206 (N_206,In_110,In_27);
or U207 (N_207,In_277,In_299);
and U208 (N_208,In_151,In_316);
nand U209 (N_209,In_158,In_58);
and U210 (N_210,In_390,In_121);
or U211 (N_211,In_146,In_405);
or U212 (N_212,In_0,In_389);
and U213 (N_213,In_75,In_453);
or U214 (N_214,In_127,In_212);
and U215 (N_215,In_347,In_196);
or U216 (N_216,In_255,In_25);
and U217 (N_217,In_13,In_157);
nand U218 (N_218,In_177,In_208);
or U219 (N_219,In_426,In_38);
or U220 (N_220,In_17,In_490);
and U221 (N_221,In_373,In_193);
or U222 (N_222,In_420,In_336);
nor U223 (N_223,In_205,In_50);
nand U224 (N_224,In_268,In_380);
nor U225 (N_225,In_440,In_341);
nand U226 (N_226,In_231,In_257);
and U227 (N_227,In_35,In_375);
nand U228 (N_228,In_465,In_69);
nor U229 (N_229,In_6,In_63);
or U230 (N_230,In_278,In_73);
or U231 (N_231,In_488,In_468);
and U232 (N_232,In_253,In_406);
nor U233 (N_233,In_96,In_20);
nand U234 (N_234,In_204,In_484);
nor U235 (N_235,In_22,In_92);
nand U236 (N_236,In_3,In_399);
or U237 (N_237,In_168,In_215);
and U238 (N_238,In_322,In_360);
or U239 (N_239,In_81,In_160);
nor U240 (N_240,In_82,In_162);
nor U241 (N_241,In_45,In_145);
and U242 (N_242,In_201,In_43);
nor U243 (N_243,In_430,In_384);
or U244 (N_244,In_413,In_355);
nand U245 (N_245,In_353,In_337);
or U246 (N_246,In_39,In_391);
nand U247 (N_247,In_457,In_455);
nor U248 (N_248,In_41,In_381);
nor U249 (N_249,In_326,In_172);
nand U250 (N_250,In_31,In_452);
nand U251 (N_251,In_240,In_272);
nor U252 (N_252,In_338,In_330);
or U253 (N_253,In_23,In_92);
and U254 (N_254,In_434,In_111);
xnor U255 (N_255,In_172,In_271);
nand U256 (N_256,In_430,In_203);
nor U257 (N_257,In_329,In_8);
and U258 (N_258,In_188,In_44);
nor U259 (N_259,In_274,In_96);
and U260 (N_260,In_447,In_57);
or U261 (N_261,In_305,In_257);
nand U262 (N_262,In_437,In_312);
or U263 (N_263,In_341,In_342);
nor U264 (N_264,In_250,In_186);
or U265 (N_265,In_77,In_267);
and U266 (N_266,In_320,In_292);
or U267 (N_267,In_229,In_202);
or U268 (N_268,In_315,In_232);
or U269 (N_269,In_376,In_69);
and U270 (N_270,In_402,In_438);
nor U271 (N_271,In_49,In_128);
nor U272 (N_272,In_289,In_445);
nor U273 (N_273,In_37,In_283);
nand U274 (N_274,In_468,In_203);
nor U275 (N_275,In_355,In_27);
and U276 (N_276,In_105,In_378);
nor U277 (N_277,In_62,In_140);
and U278 (N_278,In_12,In_204);
nand U279 (N_279,In_366,In_242);
xnor U280 (N_280,In_144,In_447);
nand U281 (N_281,In_8,In_67);
nand U282 (N_282,In_329,In_100);
or U283 (N_283,In_54,In_142);
nor U284 (N_284,In_291,In_210);
nor U285 (N_285,In_240,In_146);
or U286 (N_286,In_210,In_312);
nor U287 (N_287,In_366,In_271);
nor U288 (N_288,In_241,In_431);
nand U289 (N_289,In_312,In_85);
nor U290 (N_290,In_177,In_427);
and U291 (N_291,In_369,In_384);
nand U292 (N_292,In_160,In_104);
nor U293 (N_293,In_403,In_132);
or U294 (N_294,In_313,In_295);
and U295 (N_295,In_475,In_405);
or U296 (N_296,In_150,In_363);
nor U297 (N_297,In_412,In_67);
nor U298 (N_298,In_34,In_376);
nand U299 (N_299,In_365,In_295);
or U300 (N_300,In_109,In_24);
or U301 (N_301,In_208,In_294);
and U302 (N_302,In_282,In_336);
and U303 (N_303,In_373,In_266);
or U304 (N_304,In_136,In_188);
nor U305 (N_305,In_464,In_406);
and U306 (N_306,In_468,In_450);
nor U307 (N_307,In_167,In_290);
or U308 (N_308,In_5,In_309);
and U309 (N_309,In_131,In_491);
and U310 (N_310,In_210,In_148);
or U311 (N_311,In_478,In_62);
xor U312 (N_312,In_315,In_362);
nor U313 (N_313,In_268,In_178);
nor U314 (N_314,In_63,In_47);
nor U315 (N_315,In_449,In_201);
nor U316 (N_316,In_239,In_144);
or U317 (N_317,In_472,In_41);
or U318 (N_318,In_106,In_319);
nor U319 (N_319,In_400,In_148);
nand U320 (N_320,In_223,In_282);
or U321 (N_321,In_327,In_79);
nor U322 (N_322,In_218,In_146);
nand U323 (N_323,In_437,In_464);
nor U324 (N_324,In_68,In_224);
nand U325 (N_325,In_417,In_64);
or U326 (N_326,In_495,In_339);
and U327 (N_327,In_435,In_133);
nor U328 (N_328,In_262,In_398);
or U329 (N_329,In_276,In_373);
nand U330 (N_330,In_372,In_446);
nand U331 (N_331,In_186,In_244);
or U332 (N_332,In_32,In_101);
nand U333 (N_333,In_331,In_356);
nor U334 (N_334,In_412,In_381);
and U335 (N_335,In_176,In_59);
nor U336 (N_336,In_241,In_136);
nor U337 (N_337,In_240,In_139);
nand U338 (N_338,In_126,In_29);
and U339 (N_339,In_187,In_479);
and U340 (N_340,In_136,In_261);
and U341 (N_341,In_422,In_417);
nor U342 (N_342,In_127,In_328);
nor U343 (N_343,In_183,In_28);
nor U344 (N_344,In_454,In_399);
or U345 (N_345,In_457,In_109);
nand U346 (N_346,In_396,In_428);
nor U347 (N_347,In_209,In_307);
or U348 (N_348,In_8,In_111);
nor U349 (N_349,In_374,In_152);
nand U350 (N_350,In_312,In_136);
nand U351 (N_351,In_134,In_215);
and U352 (N_352,In_311,In_296);
nand U353 (N_353,In_288,In_435);
nor U354 (N_354,In_372,In_250);
or U355 (N_355,In_158,In_281);
and U356 (N_356,In_75,In_466);
or U357 (N_357,In_495,In_26);
xor U358 (N_358,In_49,In_132);
nor U359 (N_359,In_438,In_300);
nor U360 (N_360,In_69,In_200);
nand U361 (N_361,In_90,In_266);
or U362 (N_362,In_186,In_209);
nand U363 (N_363,In_129,In_238);
or U364 (N_364,In_394,In_66);
and U365 (N_365,In_454,In_455);
nor U366 (N_366,In_180,In_195);
nor U367 (N_367,In_490,In_179);
nand U368 (N_368,In_169,In_2);
nand U369 (N_369,In_201,In_256);
or U370 (N_370,In_11,In_281);
or U371 (N_371,In_365,In_89);
or U372 (N_372,In_191,In_40);
and U373 (N_373,In_419,In_195);
or U374 (N_374,In_73,In_279);
nand U375 (N_375,In_413,In_374);
nand U376 (N_376,In_81,In_209);
xor U377 (N_377,In_425,In_380);
and U378 (N_378,In_324,In_38);
nor U379 (N_379,In_263,In_361);
and U380 (N_380,In_119,In_416);
and U381 (N_381,In_251,In_418);
nor U382 (N_382,In_63,In_151);
nor U383 (N_383,In_417,In_463);
or U384 (N_384,In_125,In_491);
and U385 (N_385,In_5,In_438);
nand U386 (N_386,In_108,In_403);
or U387 (N_387,In_104,In_411);
nor U388 (N_388,In_267,In_469);
and U389 (N_389,In_389,In_266);
nor U390 (N_390,In_182,In_216);
nor U391 (N_391,In_46,In_396);
and U392 (N_392,In_203,In_372);
nand U393 (N_393,In_210,In_445);
and U394 (N_394,In_477,In_79);
nand U395 (N_395,In_279,In_52);
nor U396 (N_396,In_205,In_211);
nor U397 (N_397,In_15,In_400);
nor U398 (N_398,In_188,In_487);
nor U399 (N_399,In_14,In_345);
and U400 (N_400,In_238,In_457);
and U401 (N_401,In_339,In_117);
nor U402 (N_402,In_383,In_30);
nor U403 (N_403,In_323,In_268);
nor U404 (N_404,In_120,In_176);
or U405 (N_405,In_338,In_496);
nand U406 (N_406,In_166,In_224);
nand U407 (N_407,In_76,In_251);
nor U408 (N_408,In_160,In_135);
and U409 (N_409,In_265,In_250);
nor U410 (N_410,In_314,In_278);
and U411 (N_411,In_224,In_83);
or U412 (N_412,In_296,In_126);
or U413 (N_413,In_251,In_342);
and U414 (N_414,In_301,In_283);
nand U415 (N_415,In_8,In_240);
and U416 (N_416,In_227,In_143);
nand U417 (N_417,In_149,In_23);
nor U418 (N_418,In_151,In_296);
or U419 (N_419,In_219,In_351);
nor U420 (N_420,In_109,In_463);
or U421 (N_421,In_400,In_383);
nand U422 (N_422,In_219,In_154);
or U423 (N_423,In_290,In_22);
nor U424 (N_424,In_46,In_108);
nand U425 (N_425,In_185,In_489);
nand U426 (N_426,In_458,In_218);
and U427 (N_427,In_452,In_392);
nand U428 (N_428,In_339,In_240);
and U429 (N_429,In_155,In_375);
nor U430 (N_430,In_29,In_381);
or U431 (N_431,In_420,In_210);
or U432 (N_432,In_402,In_18);
nor U433 (N_433,In_382,In_208);
nand U434 (N_434,In_291,In_425);
or U435 (N_435,In_408,In_159);
or U436 (N_436,In_249,In_221);
or U437 (N_437,In_458,In_307);
or U438 (N_438,In_32,In_217);
nand U439 (N_439,In_113,In_351);
and U440 (N_440,In_159,In_399);
nand U441 (N_441,In_424,In_157);
nand U442 (N_442,In_419,In_54);
nor U443 (N_443,In_257,In_384);
nor U444 (N_444,In_154,In_164);
nor U445 (N_445,In_170,In_361);
and U446 (N_446,In_77,In_370);
nor U447 (N_447,In_7,In_439);
or U448 (N_448,In_485,In_231);
or U449 (N_449,In_148,In_59);
or U450 (N_450,In_39,In_218);
or U451 (N_451,In_397,In_335);
or U452 (N_452,In_431,In_177);
nor U453 (N_453,In_242,In_397);
or U454 (N_454,In_67,In_328);
and U455 (N_455,In_147,In_413);
and U456 (N_456,In_351,In_235);
nor U457 (N_457,In_231,In_307);
and U458 (N_458,In_440,In_444);
nor U459 (N_459,In_392,In_129);
nand U460 (N_460,In_194,In_490);
and U461 (N_461,In_26,In_316);
and U462 (N_462,In_115,In_246);
or U463 (N_463,In_81,In_465);
or U464 (N_464,In_5,In_6);
nand U465 (N_465,In_463,In_497);
and U466 (N_466,In_259,In_485);
and U467 (N_467,In_145,In_280);
nor U468 (N_468,In_355,In_28);
and U469 (N_469,In_322,In_91);
or U470 (N_470,In_470,In_101);
nand U471 (N_471,In_296,In_218);
nor U472 (N_472,In_42,In_395);
nand U473 (N_473,In_38,In_375);
and U474 (N_474,In_411,In_216);
or U475 (N_475,In_279,In_317);
and U476 (N_476,In_256,In_258);
or U477 (N_477,In_284,In_491);
and U478 (N_478,In_231,In_494);
nor U479 (N_479,In_58,In_349);
nand U480 (N_480,In_406,In_203);
or U481 (N_481,In_26,In_373);
or U482 (N_482,In_169,In_152);
nor U483 (N_483,In_104,In_481);
nand U484 (N_484,In_416,In_281);
or U485 (N_485,In_314,In_222);
and U486 (N_486,In_75,In_27);
nor U487 (N_487,In_258,In_350);
and U488 (N_488,In_407,In_159);
nor U489 (N_489,In_424,In_242);
or U490 (N_490,In_279,In_67);
and U491 (N_491,In_442,In_256);
nand U492 (N_492,In_309,In_19);
and U493 (N_493,In_0,In_447);
nor U494 (N_494,In_410,In_194);
xor U495 (N_495,In_172,In_414);
and U496 (N_496,In_416,In_39);
and U497 (N_497,In_112,In_239);
nand U498 (N_498,In_472,In_125);
nor U499 (N_499,In_262,In_316);
and U500 (N_500,In_496,In_463);
xor U501 (N_501,In_479,In_145);
nor U502 (N_502,In_411,In_210);
nor U503 (N_503,In_141,In_499);
nand U504 (N_504,In_89,In_398);
or U505 (N_505,In_437,In_75);
or U506 (N_506,In_273,In_245);
nand U507 (N_507,In_87,In_156);
nor U508 (N_508,In_300,In_148);
nor U509 (N_509,In_384,In_372);
or U510 (N_510,In_305,In_306);
nand U511 (N_511,In_420,In_166);
or U512 (N_512,In_192,In_172);
and U513 (N_513,In_383,In_24);
nor U514 (N_514,In_186,In_309);
and U515 (N_515,In_383,In_373);
and U516 (N_516,In_24,In_128);
and U517 (N_517,In_422,In_431);
or U518 (N_518,In_269,In_68);
nand U519 (N_519,In_73,In_13);
xnor U520 (N_520,In_248,In_315);
or U521 (N_521,In_407,In_13);
nor U522 (N_522,In_4,In_497);
and U523 (N_523,In_167,In_188);
or U524 (N_524,In_178,In_351);
or U525 (N_525,In_137,In_246);
or U526 (N_526,In_308,In_145);
nand U527 (N_527,In_87,In_376);
nand U528 (N_528,In_271,In_478);
nor U529 (N_529,In_53,In_64);
or U530 (N_530,In_131,In_372);
or U531 (N_531,In_84,In_468);
or U532 (N_532,In_186,In_73);
or U533 (N_533,In_186,In_417);
nand U534 (N_534,In_361,In_167);
and U535 (N_535,In_434,In_128);
or U536 (N_536,In_438,In_166);
nand U537 (N_537,In_449,In_118);
and U538 (N_538,In_490,In_446);
nor U539 (N_539,In_138,In_271);
nor U540 (N_540,In_52,In_68);
and U541 (N_541,In_255,In_335);
or U542 (N_542,In_49,In_395);
or U543 (N_543,In_302,In_357);
or U544 (N_544,In_71,In_480);
nor U545 (N_545,In_119,In_397);
nand U546 (N_546,In_341,In_408);
nand U547 (N_547,In_169,In_464);
xor U548 (N_548,In_237,In_242);
and U549 (N_549,In_210,In_403);
nor U550 (N_550,In_424,In_165);
nor U551 (N_551,In_471,In_181);
and U552 (N_552,In_70,In_356);
or U553 (N_553,In_445,In_303);
or U554 (N_554,In_197,In_40);
and U555 (N_555,In_320,In_172);
nand U556 (N_556,In_434,In_242);
or U557 (N_557,In_96,In_77);
xor U558 (N_558,In_199,In_222);
or U559 (N_559,In_372,In_284);
nor U560 (N_560,In_266,In_489);
and U561 (N_561,In_291,In_104);
nand U562 (N_562,In_70,In_297);
nand U563 (N_563,In_29,In_85);
nor U564 (N_564,In_155,In_488);
nand U565 (N_565,In_386,In_102);
nor U566 (N_566,In_261,In_375);
and U567 (N_567,In_134,In_109);
and U568 (N_568,In_10,In_370);
nand U569 (N_569,In_367,In_319);
nand U570 (N_570,In_4,In_149);
and U571 (N_571,In_365,In_96);
nor U572 (N_572,In_497,In_362);
nor U573 (N_573,In_300,In_351);
and U574 (N_574,In_332,In_20);
nor U575 (N_575,In_205,In_306);
nor U576 (N_576,In_414,In_143);
and U577 (N_577,In_160,In_230);
xor U578 (N_578,In_112,In_341);
or U579 (N_579,In_322,In_236);
nand U580 (N_580,In_64,In_422);
nor U581 (N_581,In_364,In_157);
and U582 (N_582,In_46,In_168);
xnor U583 (N_583,In_162,In_313);
or U584 (N_584,In_417,In_444);
nand U585 (N_585,In_40,In_390);
nand U586 (N_586,In_330,In_473);
nand U587 (N_587,In_270,In_112);
nand U588 (N_588,In_331,In_277);
or U589 (N_589,In_496,In_383);
or U590 (N_590,In_121,In_252);
and U591 (N_591,In_168,In_326);
nor U592 (N_592,In_317,In_313);
and U593 (N_593,In_242,In_179);
nand U594 (N_594,In_499,In_113);
or U595 (N_595,In_420,In_262);
nand U596 (N_596,In_442,In_155);
and U597 (N_597,In_295,In_235);
or U598 (N_598,In_139,In_156);
nand U599 (N_599,In_406,In_432);
and U600 (N_600,In_324,In_254);
and U601 (N_601,In_197,In_150);
nand U602 (N_602,In_92,In_394);
nor U603 (N_603,In_86,In_279);
nand U604 (N_604,In_77,In_53);
nor U605 (N_605,In_99,In_68);
or U606 (N_606,In_487,In_422);
and U607 (N_607,In_61,In_478);
and U608 (N_608,In_349,In_286);
nand U609 (N_609,In_369,In_166);
nor U610 (N_610,In_475,In_96);
and U611 (N_611,In_358,In_181);
and U612 (N_612,In_380,In_318);
and U613 (N_613,In_113,In_72);
and U614 (N_614,In_454,In_103);
and U615 (N_615,In_239,In_17);
nor U616 (N_616,In_120,In_164);
and U617 (N_617,In_453,In_209);
nand U618 (N_618,In_351,In_216);
nand U619 (N_619,In_311,In_115);
nor U620 (N_620,In_10,In_368);
nor U621 (N_621,In_58,In_368);
nand U622 (N_622,In_43,In_182);
nor U623 (N_623,In_460,In_165);
or U624 (N_624,In_222,In_184);
and U625 (N_625,In_326,In_207);
or U626 (N_626,In_287,In_234);
and U627 (N_627,In_101,In_180);
or U628 (N_628,In_469,In_200);
and U629 (N_629,In_206,In_224);
or U630 (N_630,In_372,In_32);
nor U631 (N_631,In_138,In_416);
or U632 (N_632,In_70,In_294);
and U633 (N_633,In_483,In_180);
nand U634 (N_634,In_98,In_138);
nand U635 (N_635,In_240,In_37);
nand U636 (N_636,In_31,In_129);
nand U637 (N_637,In_444,In_170);
or U638 (N_638,In_391,In_302);
nand U639 (N_639,In_158,In_333);
or U640 (N_640,In_172,In_128);
and U641 (N_641,In_298,In_354);
nor U642 (N_642,In_408,In_253);
nand U643 (N_643,In_232,In_287);
nor U644 (N_644,In_10,In_189);
nand U645 (N_645,In_378,In_219);
and U646 (N_646,In_389,In_429);
or U647 (N_647,In_3,In_151);
or U648 (N_648,In_315,In_247);
nor U649 (N_649,In_366,In_364);
nor U650 (N_650,In_73,In_121);
xor U651 (N_651,In_297,In_52);
nor U652 (N_652,In_140,In_201);
and U653 (N_653,In_453,In_374);
nor U654 (N_654,In_56,In_110);
or U655 (N_655,In_212,In_405);
nor U656 (N_656,In_266,In_208);
nor U657 (N_657,In_405,In_233);
nand U658 (N_658,In_231,In_354);
nand U659 (N_659,In_178,In_441);
nor U660 (N_660,In_117,In_384);
nand U661 (N_661,In_171,In_304);
nor U662 (N_662,In_294,In_202);
or U663 (N_663,In_398,In_91);
and U664 (N_664,In_440,In_25);
nand U665 (N_665,In_366,In_395);
and U666 (N_666,In_442,In_16);
or U667 (N_667,In_460,In_309);
and U668 (N_668,In_291,In_142);
and U669 (N_669,In_378,In_395);
or U670 (N_670,In_210,In_101);
nor U671 (N_671,In_326,In_399);
and U672 (N_672,In_34,In_115);
and U673 (N_673,In_273,In_379);
and U674 (N_674,In_204,In_393);
or U675 (N_675,In_470,In_194);
and U676 (N_676,In_128,In_237);
and U677 (N_677,In_222,In_477);
or U678 (N_678,In_195,In_375);
nand U679 (N_679,In_387,In_215);
nor U680 (N_680,In_460,In_384);
or U681 (N_681,In_184,In_77);
or U682 (N_682,In_181,In_478);
or U683 (N_683,In_55,In_108);
or U684 (N_684,In_30,In_116);
nor U685 (N_685,In_265,In_257);
nand U686 (N_686,In_472,In_213);
nand U687 (N_687,In_410,In_258);
or U688 (N_688,In_186,In_138);
and U689 (N_689,In_415,In_183);
nand U690 (N_690,In_109,In_110);
or U691 (N_691,In_432,In_33);
nor U692 (N_692,In_334,In_0);
or U693 (N_693,In_113,In_237);
xor U694 (N_694,In_482,In_187);
nand U695 (N_695,In_225,In_291);
nor U696 (N_696,In_302,In_472);
nor U697 (N_697,In_334,In_472);
or U698 (N_698,In_46,In_423);
nand U699 (N_699,In_426,In_260);
nor U700 (N_700,In_385,In_424);
or U701 (N_701,In_426,In_242);
and U702 (N_702,In_13,In_456);
or U703 (N_703,In_38,In_441);
and U704 (N_704,In_459,In_132);
and U705 (N_705,In_122,In_284);
or U706 (N_706,In_126,In_219);
or U707 (N_707,In_3,In_449);
nand U708 (N_708,In_394,In_204);
nor U709 (N_709,In_206,In_127);
and U710 (N_710,In_189,In_154);
and U711 (N_711,In_327,In_75);
or U712 (N_712,In_154,In_32);
nand U713 (N_713,In_180,In_346);
and U714 (N_714,In_375,In_451);
nand U715 (N_715,In_370,In_352);
or U716 (N_716,In_237,In_68);
nor U717 (N_717,In_229,In_105);
and U718 (N_718,In_73,In_432);
nor U719 (N_719,In_60,In_116);
and U720 (N_720,In_296,In_445);
nand U721 (N_721,In_297,In_271);
nand U722 (N_722,In_468,In_366);
nor U723 (N_723,In_479,In_14);
and U724 (N_724,In_249,In_33);
nor U725 (N_725,In_112,In_471);
or U726 (N_726,In_42,In_75);
and U727 (N_727,In_312,In_257);
nor U728 (N_728,In_328,In_345);
and U729 (N_729,In_285,In_266);
nor U730 (N_730,In_2,In_85);
and U731 (N_731,In_209,In_221);
nor U732 (N_732,In_314,In_308);
and U733 (N_733,In_178,In_235);
nand U734 (N_734,In_162,In_475);
and U735 (N_735,In_128,In_272);
and U736 (N_736,In_492,In_24);
and U737 (N_737,In_408,In_484);
nor U738 (N_738,In_20,In_356);
nand U739 (N_739,In_25,In_364);
or U740 (N_740,In_369,In_179);
or U741 (N_741,In_456,In_124);
and U742 (N_742,In_319,In_90);
and U743 (N_743,In_77,In_133);
nor U744 (N_744,In_263,In_271);
nand U745 (N_745,In_271,In_481);
nand U746 (N_746,In_221,In_72);
or U747 (N_747,In_350,In_245);
nor U748 (N_748,In_250,In_160);
nor U749 (N_749,In_304,In_197);
and U750 (N_750,In_202,In_262);
nand U751 (N_751,In_434,In_267);
nand U752 (N_752,In_45,In_449);
or U753 (N_753,In_219,In_411);
or U754 (N_754,In_152,In_332);
nand U755 (N_755,In_153,In_318);
nand U756 (N_756,In_79,In_95);
nand U757 (N_757,In_280,In_478);
nor U758 (N_758,In_415,In_35);
or U759 (N_759,In_450,In_104);
nand U760 (N_760,In_324,In_71);
and U761 (N_761,In_269,In_57);
nor U762 (N_762,In_350,In_131);
nor U763 (N_763,In_487,In_183);
nor U764 (N_764,In_439,In_374);
nand U765 (N_765,In_210,In_302);
or U766 (N_766,In_324,In_128);
nor U767 (N_767,In_481,In_34);
and U768 (N_768,In_21,In_44);
and U769 (N_769,In_464,In_271);
or U770 (N_770,In_218,In_385);
nor U771 (N_771,In_215,In_425);
and U772 (N_772,In_15,In_96);
nand U773 (N_773,In_40,In_169);
nand U774 (N_774,In_375,In_207);
nand U775 (N_775,In_379,In_258);
or U776 (N_776,In_408,In_322);
and U777 (N_777,In_493,In_451);
and U778 (N_778,In_44,In_432);
nand U779 (N_779,In_48,In_393);
nand U780 (N_780,In_358,In_247);
and U781 (N_781,In_0,In_331);
nor U782 (N_782,In_117,In_52);
nand U783 (N_783,In_464,In_102);
and U784 (N_784,In_134,In_262);
and U785 (N_785,In_390,In_99);
or U786 (N_786,In_386,In_401);
nor U787 (N_787,In_17,In_488);
nor U788 (N_788,In_214,In_138);
or U789 (N_789,In_332,In_340);
nor U790 (N_790,In_89,In_351);
nor U791 (N_791,In_253,In_63);
and U792 (N_792,In_340,In_474);
or U793 (N_793,In_224,In_310);
xnor U794 (N_794,In_360,In_345);
or U795 (N_795,In_309,In_149);
or U796 (N_796,In_489,In_412);
or U797 (N_797,In_481,In_147);
and U798 (N_798,In_340,In_191);
nor U799 (N_799,In_374,In_91);
and U800 (N_800,In_447,In_102);
nor U801 (N_801,In_60,In_317);
and U802 (N_802,In_91,In_243);
nand U803 (N_803,In_96,In_331);
nor U804 (N_804,In_293,In_470);
nor U805 (N_805,In_191,In_389);
nor U806 (N_806,In_311,In_335);
and U807 (N_807,In_222,In_382);
and U808 (N_808,In_393,In_412);
or U809 (N_809,In_376,In_131);
or U810 (N_810,In_306,In_369);
nor U811 (N_811,In_220,In_462);
and U812 (N_812,In_232,In_372);
nor U813 (N_813,In_288,In_75);
and U814 (N_814,In_457,In_153);
and U815 (N_815,In_73,In_434);
nand U816 (N_816,In_288,In_67);
nand U817 (N_817,In_177,In_87);
and U818 (N_818,In_371,In_85);
xnor U819 (N_819,In_367,In_376);
or U820 (N_820,In_350,In_358);
nor U821 (N_821,In_106,In_389);
and U822 (N_822,In_193,In_335);
and U823 (N_823,In_266,In_252);
xnor U824 (N_824,In_56,In_191);
nor U825 (N_825,In_426,In_57);
and U826 (N_826,In_458,In_347);
or U827 (N_827,In_429,In_297);
nor U828 (N_828,In_109,In_73);
or U829 (N_829,In_116,In_356);
or U830 (N_830,In_235,In_377);
nor U831 (N_831,In_458,In_280);
and U832 (N_832,In_174,In_262);
nor U833 (N_833,In_94,In_151);
and U834 (N_834,In_430,In_489);
nor U835 (N_835,In_234,In_32);
or U836 (N_836,In_122,In_265);
and U837 (N_837,In_150,In_382);
nor U838 (N_838,In_256,In_380);
or U839 (N_839,In_53,In_271);
or U840 (N_840,In_7,In_277);
or U841 (N_841,In_367,In_446);
or U842 (N_842,In_135,In_76);
nor U843 (N_843,In_295,In_246);
nor U844 (N_844,In_96,In_445);
and U845 (N_845,In_395,In_361);
and U846 (N_846,In_150,In_146);
or U847 (N_847,In_332,In_47);
nor U848 (N_848,In_195,In_425);
and U849 (N_849,In_225,In_236);
nand U850 (N_850,In_65,In_55);
and U851 (N_851,In_144,In_21);
nor U852 (N_852,In_325,In_395);
and U853 (N_853,In_56,In_292);
nor U854 (N_854,In_167,In_129);
or U855 (N_855,In_191,In_184);
nor U856 (N_856,In_320,In_79);
nor U857 (N_857,In_375,In_445);
and U858 (N_858,In_179,In_455);
or U859 (N_859,In_14,In_397);
and U860 (N_860,In_8,In_207);
and U861 (N_861,In_85,In_237);
or U862 (N_862,In_41,In_353);
and U863 (N_863,In_115,In_465);
and U864 (N_864,In_494,In_123);
and U865 (N_865,In_350,In_209);
nor U866 (N_866,In_377,In_487);
nand U867 (N_867,In_289,In_396);
and U868 (N_868,In_325,In_48);
and U869 (N_869,In_153,In_194);
nand U870 (N_870,In_390,In_241);
nand U871 (N_871,In_270,In_442);
nor U872 (N_872,In_37,In_282);
and U873 (N_873,In_249,In_202);
nand U874 (N_874,In_307,In_24);
and U875 (N_875,In_26,In_388);
nor U876 (N_876,In_393,In_137);
nand U877 (N_877,In_77,In_334);
nand U878 (N_878,In_178,In_107);
and U879 (N_879,In_254,In_196);
or U880 (N_880,In_147,In_38);
nand U881 (N_881,In_377,In_27);
nor U882 (N_882,In_394,In_198);
or U883 (N_883,In_365,In_389);
and U884 (N_884,In_451,In_446);
nand U885 (N_885,In_272,In_298);
and U886 (N_886,In_133,In_397);
and U887 (N_887,In_100,In_349);
nor U888 (N_888,In_141,In_219);
nor U889 (N_889,In_112,In_61);
nand U890 (N_890,In_68,In_110);
nand U891 (N_891,In_253,In_459);
nand U892 (N_892,In_193,In_11);
nor U893 (N_893,In_277,In_160);
nand U894 (N_894,In_62,In_330);
or U895 (N_895,In_234,In_136);
nand U896 (N_896,In_282,In_4);
and U897 (N_897,In_308,In_270);
and U898 (N_898,In_107,In_426);
and U899 (N_899,In_281,In_349);
or U900 (N_900,In_11,In_43);
and U901 (N_901,In_394,In_337);
and U902 (N_902,In_142,In_470);
nand U903 (N_903,In_45,In_34);
and U904 (N_904,In_201,In_462);
nor U905 (N_905,In_28,In_127);
or U906 (N_906,In_145,In_289);
nor U907 (N_907,In_239,In_15);
or U908 (N_908,In_470,In_300);
or U909 (N_909,In_235,In_328);
and U910 (N_910,In_205,In_110);
and U911 (N_911,In_289,In_183);
or U912 (N_912,In_239,In_72);
and U913 (N_913,In_484,In_4);
nor U914 (N_914,In_74,In_240);
nand U915 (N_915,In_273,In_26);
nand U916 (N_916,In_499,In_28);
or U917 (N_917,In_47,In_413);
and U918 (N_918,In_259,In_421);
nand U919 (N_919,In_62,In_318);
and U920 (N_920,In_194,In_74);
nor U921 (N_921,In_156,In_499);
nand U922 (N_922,In_107,In_419);
or U923 (N_923,In_447,In_46);
and U924 (N_924,In_302,In_355);
or U925 (N_925,In_280,In_344);
and U926 (N_926,In_241,In_247);
nor U927 (N_927,In_333,In_116);
or U928 (N_928,In_120,In_448);
or U929 (N_929,In_327,In_46);
nor U930 (N_930,In_430,In_143);
nand U931 (N_931,In_118,In_399);
or U932 (N_932,In_422,In_359);
nor U933 (N_933,In_289,In_405);
or U934 (N_934,In_397,In_240);
nor U935 (N_935,In_63,In_130);
and U936 (N_936,In_300,In_281);
nor U937 (N_937,In_417,In_282);
nor U938 (N_938,In_419,In_332);
and U939 (N_939,In_68,In_279);
or U940 (N_940,In_71,In_60);
nor U941 (N_941,In_480,In_456);
nand U942 (N_942,In_227,In_254);
nor U943 (N_943,In_84,In_78);
and U944 (N_944,In_246,In_207);
xnor U945 (N_945,In_265,In_21);
and U946 (N_946,In_227,In_104);
nand U947 (N_947,In_326,In_251);
nand U948 (N_948,In_311,In_236);
nand U949 (N_949,In_216,In_358);
nand U950 (N_950,In_287,In_92);
and U951 (N_951,In_251,In_383);
nor U952 (N_952,In_289,In_466);
and U953 (N_953,In_297,In_299);
and U954 (N_954,In_275,In_416);
nand U955 (N_955,In_416,In_270);
and U956 (N_956,In_168,In_157);
or U957 (N_957,In_137,In_157);
nor U958 (N_958,In_347,In_149);
and U959 (N_959,In_184,In_466);
or U960 (N_960,In_60,In_454);
nor U961 (N_961,In_302,In_256);
or U962 (N_962,In_95,In_223);
nand U963 (N_963,In_99,In_498);
or U964 (N_964,In_449,In_210);
or U965 (N_965,In_293,In_192);
or U966 (N_966,In_96,In_498);
or U967 (N_967,In_99,In_23);
nand U968 (N_968,In_79,In_87);
nor U969 (N_969,In_492,In_17);
nand U970 (N_970,In_88,In_382);
nand U971 (N_971,In_176,In_7);
and U972 (N_972,In_322,In_272);
nor U973 (N_973,In_180,In_349);
nor U974 (N_974,In_289,In_304);
and U975 (N_975,In_315,In_203);
nor U976 (N_976,In_64,In_356);
or U977 (N_977,In_68,In_307);
xor U978 (N_978,In_396,In_51);
nor U979 (N_979,In_383,In_294);
or U980 (N_980,In_230,In_37);
nor U981 (N_981,In_252,In_378);
and U982 (N_982,In_83,In_423);
and U983 (N_983,In_220,In_456);
nor U984 (N_984,In_409,In_414);
nor U985 (N_985,In_301,In_92);
nand U986 (N_986,In_256,In_464);
nor U987 (N_987,In_186,In_421);
nand U988 (N_988,In_323,In_330);
and U989 (N_989,In_205,In_472);
and U990 (N_990,In_349,In_193);
nand U991 (N_991,In_260,In_332);
xnor U992 (N_992,In_245,In_94);
and U993 (N_993,In_86,In_371);
or U994 (N_994,In_401,In_429);
or U995 (N_995,In_77,In_270);
and U996 (N_996,In_258,In_204);
nand U997 (N_997,In_55,In_427);
nand U998 (N_998,In_184,In_330);
and U999 (N_999,In_179,In_38);
nor U1000 (N_1000,N_869,N_440);
and U1001 (N_1001,N_933,N_258);
and U1002 (N_1002,N_732,N_542);
and U1003 (N_1003,N_294,N_118);
or U1004 (N_1004,N_25,N_361);
and U1005 (N_1005,N_901,N_721);
nand U1006 (N_1006,N_739,N_94);
or U1007 (N_1007,N_283,N_375);
nor U1008 (N_1008,N_62,N_301);
and U1009 (N_1009,N_667,N_726);
nor U1010 (N_1010,N_180,N_686);
and U1011 (N_1011,N_167,N_782);
nand U1012 (N_1012,N_146,N_663);
or U1013 (N_1013,N_989,N_97);
nand U1014 (N_1014,N_14,N_508);
and U1015 (N_1015,N_829,N_854);
or U1016 (N_1016,N_221,N_904);
nand U1017 (N_1017,N_80,N_572);
nand U1018 (N_1018,N_99,N_831);
nor U1019 (N_1019,N_130,N_10);
or U1020 (N_1020,N_597,N_677);
and U1021 (N_1021,N_599,N_308);
or U1022 (N_1022,N_557,N_928);
nand U1023 (N_1023,N_90,N_287);
nor U1024 (N_1024,N_817,N_973);
and U1025 (N_1025,N_816,N_656);
nand U1026 (N_1026,N_551,N_967);
nand U1027 (N_1027,N_596,N_332);
nor U1028 (N_1028,N_73,N_290);
nor U1029 (N_1029,N_704,N_864);
and U1030 (N_1030,N_101,N_281);
or U1031 (N_1031,N_250,N_859);
and U1032 (N_1032,N_780,N_911);
nand U1033 (N_1033,N_405,N_601);
or U1034 (N_1034,N_564,N_809);
nor U1035 (N_1035,N_365,N_211);
nand U1036 (N_1036,N_842,N_333);
and U1037 (N_1037,N_735,N_451);
xor U1038 (N_1038,N_231,N_875);
nor U1039 (N_1039,N_756,N_335);
nor U1040 (N_1040,N_835,N_494);
and U1041 (N_1041,N_45,N_456);
nor U1042 (N_1042,N_255,N_822);
and U1043 (N_1043,N_515,N_662);
or U1044 (N_1044,N_34,N_555);
nand U1045 (N_1045,N_806,N_749);
or U1046 (N_1046,N_549,N_593);
or U1047 (N_1047,N_522,N_181);
nor U1048 (N_1048,N_468,N_434);
or U1049 (N_1049,N_107,N_958);
nor U1050 (N_1050,N_903,N_188);
nor U1051 (N_1051,N_190,N_879);
or U1052 (N_1052,N_32,N_988);
or U1053 (N_1053,N_364,N_998);
and U1054 (N_1054,N_942,N_923);
and U1055 (N_1055,N_486,N_356);
nand U1056 (N_1056,N_999,N_675);
and U1057 (N_1057,N_846,N_166);
and U1058 (N_1058,N_337,N_743);
or U1059 (N_1059,N_128,N_204);
nor U1060 (N_1060,N_591,N_27);
nor U1061 (N_1061,N_446,N_125);
nand U1062 (N_1062,N_470,N_814);
nor U1063 (N_1063,N_793,N_908);
and U1064 (N_1064,N_303,N_262);
nand U1065 (N_1065,N_855,N_905);
and U1066 (N_1066,N_55,N_254);
and U1067 (N_1067,N_733,N_100);
nor U1068 (N_1068,N_552,N_981);
or U1069 (N_1069,N_21,N_789);
nand U1070 (N_1070,N_305,N_659);
or U1071 (N_1071,N_219,N_61);
and U1072 (N_1072,N_98,N_42);
or U1073 (N_1073,N_285,N_89);
nor U1074 (N_1074,N_917,N_629);
nand U1075 (N_1075,N_883,N_347);
nor U1076 (N_1076,N_171,N_397);
nand U1077 (N_1077,N_723,N_443);
or U1078 (N_1078,N_380,N_968);
or U1079 (N_1079,N_853,N_319);
or U1080 (N_1080,N_409,N_830);
or U1081 (N_1081,N_577,N_536);
and U1082 (N_1082,N_872,N_530);
or U1083 (N_1083,N_896,N_401);
and U1084 (N_1084,N_37,N_202);
and U1085 (N_1085,N_623,N_529);
and U1086 (N_1086,N_613,N_289);
or U1087 (N_1087,N_873,N_275);
or U1088 (N_1088,N_438,N_709);
or U1089 (N_1089,N_787,N_189);
and U1090 (N_1090,N_436,N_40);
nand U1091 (N_1091,N_897,N_509);
and U1092 (N_1092,N_479,N_769);
nor U1093 (N_1093,N_783,N_102);
and U1094 (N_1094,N_352,N_791);
or U1095 (N_1095,N_444,N_105);
nand U1096 (N_1096,N_495,N_909);
or U1097 (N_1097,N_164,N_785);
and U1098 (N_1098,N_428,N_306);
nor U1099 (N_1099,N_516,N_573);
nor U1100 (N_1100,N_241,N_149);
and U1101 (N_1101,N_651,N_417);
or U1102 (N_1102,N_671,N_960);
or U1103 (N_1103,N_758,N_60);
or U1104 (N_1104,N_912,N_626);
nand U1105 (N_1105,N_565,N_433);
or U1106 (N_1106,N_278,N_950);
and U1107 (N_1107,N_658,N_886);
nand U1108 (N_1108,N_194,N_8);
and U1109 (N_1109,N_569,N_488);
nand U1110 (N_1110,N_583,N_839);
or U1111 (N_1111,N_725,N_578);
nor U1112 (N_1112,N_236,N_199);
nor U1113 (N_1113,N_799,N_646);
or U1114 (N_1114,N_946,N_453);
and U1115 (N_1115,N_710,N_505);
or U1116 (N_1116,N_172,N_74);
or U1117 (N_1117,N_96,N_421);
nor U1118 (N_1118,N_330,N_874);
and U1119 (N_1119,N_884,N_888);
nor U1120 (N_1120,N_110,N_638);
nor U1121 (N_1121,N_771,N_235);
and U1122 (N_1122,N_770,N_684);
or U1123 (N_1123,N_695,N_19);
or U1124 (N_1124,N_630,N_768);
and U1125 (N_1125,N_863,N_373);
and U1126 (N_1126,N_997,N_270);
and U1127 (N_1127,N_512,N_339);
and U1128 (N_1128,N_13,N_681);
and U1129 (N_1129,N_574,N_68);
nand U1130 (N_1130,N_594,N_585);
nand U1131 (N_1131,N_891,N_28);
nand U1132 (N_1132,N_95,N_767);
and U1133 (N_1133,N_992,N_366);
or U1134 (N_1134,N_72,N_866);
or U1135 (N_1135,N_498,N_159);
or U1136 (N_1136,N_900,N_419);
xor U1137 (N_1137,N_325,N_331);
nand U1138 (N_1138,N_393,N_198);
or U1139 (N_1139,N_852,N_466);
nand U1140 (N_1140,N_711,N_913);
or U1141 (N_1141,N_930,N_961);
nand U1142 (N_1142,N_56,N_895);
nand U1143 (N_1143,N_396,N_476);
nor U1144 (N_1144,N_122,N_416);
nor U1145 (N_1145,N_947,N_408);
nand U1146 (N_1146,N_642,N_535);
or U1147 (N_1147,N_309,N_83);
nand U1148 (N_1148,N_272,N_265);
or U1149 (N_1149,N_877,N_261);
nand U1150 (N_1150,N_819,N_918);
nand U1151 (N_1151,N_131,N_773);
nor U1152 (N_1152,N_567,N_894);
or U1153 (N_1153,N_970,N_385);
nor U1154 (N_1154,N_291,N_459);
nor U1155 (N_1155,N_774,N_959);
nor U1156 (N_1156,N_136,N_398);
nor U1157 (N_1157,N_78,N_951);
nor U1158 (N_1158,N_197,N_279);
nand U1159 (N_1159,N_581,N_632);
nor U1160 (N_1160,N_423,N_251);
or U1161 (N_1161,N_841,N_374);
and U1162 (N_1162,N_457,N_161);
and U1163 (N_1163,N_445,N_966);
nand U1164 (N_1164,N_203,N_617);
nor U1165 (N_1165,N_639,N_314);
xnor U1166 (N_1166,N_145,N_943);
nor U1167 (N_1167,N_742,N_304);
and U1168 (N_1168,N_969,N_519);
and U1169 (N_1169,N_588,N_134);
and U1170 (N_1170,N_354,N_82);
or U1171 (N_1171,N_195,N_391);
nor U1172 (N_1172,N_160,N_79);
nor U1173 (N_1173,N_697,N_592);
and U1174 (N_1174,N_600,N_266);
nand U1175 (N_1175,N_316,N_182);
or U1176 (N_1176,N_232,N_112);
nor U1177 (N_1177,N_399,N_129);
or U1178 (N_1178,N_679,N_367);
nor U1179 (N_1179,N_158,N_851);
or U1180 (N_1180,N_482,N_926);
nor U1181 (N_1181,N_276,N_245);
nor U1182 (N_1182,N_964,N_868);
or U1183 (N_1183,N_400,N_76);
or U1184 (N_1184,N_702,N_485);
nor U1185 (N_1185,N_802,N_746);
nor U1186 (N_1186,N_755,N_560);
nand U1187 (N_1187,N_18,N_718);
and U1188 (N_1188,N_307,N_507);
or U1189 (N_1189,N_982,N_383);
and U1190 (N_1190,N_532,N_827);
and U1191 (N_1191,N_528,N_193);
and U1192 (N_1192,N_323,N_680);
or U1193 (N_1193,N_857,N_716);
nand U1194 (N_1194,N_389,N_558);
and U1195 (N_1195,N_329,N_708);
nor U1196 (N_1196,N_431,N_929);
or U1197 (N_1197,N_889,N_86);
and U1198 (N_1198,N_526,N_700);
or U1199 (N_1199,N_493,N_545);
and U1200 (N_1200,N_22,N_907);
nand U1201 (N_1201,N_664,N_922);
nand U1202 (N_1202,N_993,N_411);
and U1203 (N_1203,N_985,N_313);
or U1204 (N_1204,N_388,N_355);
and U1205 (N_1205,N_893,N_412);
nor U1206 (N_1206,N_510,N_682);
or U1207 (N_1207,N_832,N_673);
nand U1208 (N_1208,N_111,N_442);
and U1209 (N_1209,N_514,N_604);
or U1210 (N_1210,N_44,N_243);
or U1211 (N_1211,N_688,N_991);
and U1212 (N_1212,N_404,N_848);
nand U1213 (N_1213,N_284,N_990);
nand U1214 (N_1214,N_685,N_847);
and U1215 (N_1215,N_731,N_127);
nor U1216 (N_1216,N_792,N_69);
or U1217 (N_1217,N_467,N_690);
nand U1218 (N_1218,N_437,N_226);
or U1219 (N_1219,N_489,N_286);
nor U1220 (N_1220,N_384,N_887);
nand U1221 (N_1221,N_3,N_871);
nand U1222 (N_1222,N_582,N_17);
and U1223 (N_1223,N_106,N_694);
or U1224 (N_1224,N_33,N_778);
nand U1225 (N_1225,N_51,N_715);
nand U1226 (N_1226,N_899,N_501);
nand U1227 (N_1227,N_174,N_425);
nand U1228 (N_1228,N_840,N_363);
nor U1229 (N_1229,N_815,N_260);
or U1230 (N_1230,N_475,N_296);
nor U1231 (N_1231,N_312,N_935);
nand U1232 (N_1232,N_187,N_531);
and U1233 (N_1233,N_201,N_561);
and U1234 (N_1234,N_644,N_916);
and U1235 (N_1235,N_687,N_775);
and U1236 (N_1236,N_183,N_571);
xor U1237 (N_1237,N_280,N_580);
nor U1238 (N_1238,N_579,N_327);
and U1239 (N_1239,N_402,N_665);
nor U1240 (N_1240,N_661,N_120);
and U1241 (N_1241,N_953,N_302);
or U1242 (N_1242,N_293,N_297);
or U1243 (N_1243,N_734,N_714);
and U1244 (N_1244,N_372,N_234);
nor U1245 (N_1245,N_628,N_184);
nand U1246 (N_1246,N_669,N_794);
nand U1247 (N_1247,N_359,N_455);
or U1248 (N_1248,N_70,N_30);
nand U1249 (N_1249,N_547,N_945);
or U1250 (N_1250,N_796,N_504);
nor U1251 (N_1251,N_965,N_995);
and U1252 (N_1252,N_225,N_539);
nand U1253 (N_1253,N_621,N_382);
or U1254 (N_1254,N_826,N_392);
nand U1255 (N_1255,N_103,N_503);
nor U1256 (N_1256,N_150,N_138);
or U1257 (N_1257,N_473,N_538);
and U1258 (N_1258,N_633,N_244);
nand U1259 (N_1259,N_533,N_776);
or U1260 (N_1260,N_518,N_341);
and U1261 (N_1261,N_208,N_540);
nand U1262 (N_1262,N_26,N_834);
and U1263 (N_1263,N_439,N_606);
nand U1264 (N_1264,N_91,N_744);
nor U1265 (N_1265,N_932,N_2);
or U1266 (N_1266,N_403,N_747);
or U1267 (N_1267,N_546,N_925);
or U1268 (N_1268,N_169,N_67);
and U1269 (N_1269,N_213,N_605);
nand U1270 (N_1270,N_570,N_607);
nor U1271 (N_1271,N_880,N_524);
and U1272 (N_1272,N_484,N_240);
or U1273 (N_1273,N_104,N_952);
or U1274 (N_1274,N_590,N_919);
nor U1275 (N_1275,N_821,N_348);
or U1276 (N_1276,N_870,N_616);
nor U1277 (N_1277,N_0,N_228);
and U1278 (N_1278,N_192,N_766);
or U1279 (N_1279,N_556,N_119);
nand U1280 (N_1280,N_781,N_420);
or U1281 (N_1281,N_608,N_263);
or U1282 (N_1282,N_59,N_563);
or U1283 (N_1283,N_653,N_618);
and U1284 (N_1284,N_788,N_523);
nand U1285 (N_1285,N_462,N_748);
and U1286 (N_1286,N_71,N_483);
or U1287 (N_1287,N_620,N_757);
or U1288 (N_1288,N_689,N_975);
or U1289 (N_1289,N_506,N_954);
nor U1290 (N_1290,N_386,N_343);
nor U1291 (N_1291,N_155,N_387);
and U1292 (N_1292,N_427,N_311);
or U1293 (N_1293,N_862,N_490);
xor U1294 (N_1294,N_649,N_962);
nand U1295 (N_1295,N_902,N_414);
or U1296 (N_1296,N_619,N_804);
nor U1297 (N_1297,N_141,N_625);
nand U1298 (N_1298,N_41,N_740);
nand U1299 (N_1299,N_610,N_299);
nand U1300 (N_1300,N_940,N_974);
nor U1301 (N_1301,N_39,N_713);
nand U1302 (N_1302,N_274,N_843);
nor U1303 (N_1303,N_537,N_336);
nand U1304 (N_1304,N_239,N_116);
or U1305 (N_1305,N_481,N_142);
or U1306 (N_1306,N_683,N_924);
and U1307 (N_1307,N_360,N_471);
nor U1308 (N_1308,N_906,N_492);
nand U1309 (N_1309,N_148,N_818);
or U1310 (N_1310,N_828,N_252);
and U1311 (N_1311,N_666,N_271);
nand U1312 (N_1312,N_185,N_268);
nand U1313 (N_1313,N_795,N_371);
and U1314 (N_1314,N_595,N_223);
and U1315 (N_1315,N_139,N_117);
and U1316 (N_1316,N_315,N_282);
nor U1317 (N_1317,N_342,N_29);
or U1318 (N_1318,N_892,N_121);
or U1319 (N_1319,N_318,N_267);
or U1320 (N_1320,N_249,N_153);
nor U1321 (N_1321,N_43,N_75);
and U1322 (N_1322,N_728,N_586);
nor U1323 (N_1323,N_738,N_670);
and U1324 (N_1324,N_469,N_986);
nor U1325 (N_1325,N_353,N_979);
nor U1326 (N_1326,N_338,N_132);
nand U1327 (N_1327,N_752,N_701);
nand U1328 (N_1328,N_452,N_256);
nand U1329 (N_1329,N_491,N_465);
nand U1330 (N_1330,N_890,N_340);
nand U1331 (N_1331,N_635,N_177);
and U1332 (N_1332,N_277,N_322);
and U1333 (N_1333,N_429,N_641);
and U1334 (N_1334,N_449,N_57);
or U1335 (N_1335,N_810,N_422);
nor U1336 (N_1336,N_779,N_882);
and U1337 (N_1337,N_165,N_430);
nor U1338 (N_1338,N_636,N_797);
nand U1339 (N_1339,N_936,N_114);
or U1340 (N_1340,N_205,N_948);
nor U1341 (N_1341,N_938,N_762);
or U1342 (N_1342,N_584,N_645);
nor U1343 (N_1343,N_937,N_634);
and U1344 (N_1344,N_233,N_66);
or U1345 (N_1345,N_5,N_461);
or U1346 (N_1346,N_273,N_115);
nand U1347 (N_1347,N_759,N_980);
nor U1348 (N_1348,N_648,N_175);
nand U1349 (N_1349,N_212,N_589);
nor U1350 (N_1350,N_963,N_217);
and U1351 (N_1351,N_643,N_248);
and U1352 (N_1352,N_63,N_381);
nand U1353 (N_1353,N_813,N_300);
and U1354 (N_1354,N_124,N_820);
and U1355 (N_1355,N_178,N_377);
and U1356 (N_1356,N_84,N_844);
nand U1357 (N_1357,N_849,N_587);
nor U1358 (N_1358,N_707,N_502);
xor U1359 (N_1359,N_257,N_370);
or U1360 (N_1360,N_154,N_612);
or U1361 (N_1361,N_737,N_224);
or U1362 (N_1362,N_576,N_151);
and U1363 (N_1363,N_562,N_237);
and U1364 (N_1364,N_511,N_113);
and U1365 (N_1365,N_603,N_441);
nor U1366 (N_1366,N_144,N_133);
nor U1367 (N_1367,N_956,N_173);
and U1368 (N_1368,N_46,N_741);
or U1369 (N_1369,N_460,N_777);
nor U1370 (N_1370,N_362,N_939);
and U1371 (N_1371,N_58,N_477);
nor U1372 (N_1372,N_949,N_824);
nor U1373 (N_1373,N_369,N_676);
or U1374 (N_1374,N_298,N_93);
or U1375 (N_1375,N_344,N_81);
nand U1376 (N_1376,N_525,N_140);
or U1377 (N_1377,N_147,N_521);
or U1378 (N_1378,N_227,N_931);
nand U1379 (N_1379,N_760,N_432);
and U1380 (N_1380,N_602,N_152);
nor U1381 (N_1381,N_914,N_668);
nor U1382 (N_1382,N_126,N_881);
and U1383 (N_1383,N_915,N_31);
and U1384 (N_1384,N_786,N_196);
and U1385 (N_1385,N_898,N_168);
and U1386 (N_1386,N_487,N_143);
and U1387 (N_1387,N_259,N_837);
or U1388 (N_1388,N_611,N_876);
nor U1389 (N_1389,N_800,N_54);
and U1390 (N_1390,N_207,N_418);
nor U1391 (N_1391,N_88,N_415);
and U1392 (N_1392,N_253,N_288);
nor U1393 (N_1393,N_246,N_699);
nand U1394 (N_1394,N_861,N_660);
or U1395 (N_1395,N_358,N_238);
nand U1396 (N_1396,N_705,N_614);
or U1397 (N_1397,N_350,N_520);
nand U1398 (N_1398,N_957,N_672);
or U1399 (N_1399,N_978,N_87);
nor U1400 (N_1400,N_765,N_229);
nand U1401 (N_1401,N_627,N_654);
or U1402 (N_1402,N_230,N_410);
nor U1403 (N_1403,N_550,N_772);
and U1404 (N_1404,N_368,N_696);
nand U1405 (N_1405,N_801,N_320);
nor U1406 (N_1406,N_860,N_424);
or U1407 (N_1407,N_135,N_764);
nor U1408 (N_1408,N_983,N_376);
nand U1409 (N_1409,N_480,N_811);
or U1410 (N_1410,N_220,N_264);
nor U1411 (N_1411,N_210,N_326);
nand U1412 (N_1412,N_47,N_463);
and U1413 (N_1413,N_631,N_163);
and U1414 (N_1414,N_109,N_971);
nor U1415 (N_1415,N_9,N_807);
and U1416 (N_1416,N_703,N_295);
or U1417 (N_1417,N_534,N_652);
nand U1418 (N_1418,N_609,N_729);
or U1419 (N_1419,N_994,N_678);
and U1420 (N_1420,N_38,N_598);
nor U1421 (N_1421,N_214,N_750);
nor U1422 (N_1422,N_16,N_317);
or U1423 (N_1423,N_186,N_176);
or U1424 (N_1424,N_833,N_500);
nand U1425 (N_1425,N_987,N_996);
and U1426 (N_1426,N_458,N_35);
nand U1427 (N_1427,N_170,N_191);
nand U1428 (N_1428,N_77,N_858);
or U1429 (N_1429,N_379,N_247);
nand U1430 (N_1430,N_885,N_691);
or U1431 (N_1431,N_790,N_559);
and U1432 (N_1432,N_717,N_349);
or U1433 (N_1433,N_637,N_753);
nand U1434 (N_1434,N_413,N_910);
or U1435 (N_1435,N_655,N_334);
or U1436 (N_1436,N_693,N_209);
nand U1437 (N_1437,N_798,N_23);
nor U1438 (N_1438,N_447,N_215);
and U1439 (N_1439,N_543,N_20);
nor U1440 (N_1440,N_823,N_328);
or U1441 (N_1441,N_692,N_108);
nand U1442 (N_1442,N_568,N_216);
nor U1443 (N_1443,N_838,N_137);
nor U1444 (N_1444,N_53,N_977);
nand U1445 (N_1445,N_944,N_49);
nor U1446 (N_1446,N_156,N_941);
and U1447 (N_1447,N_865,N_984);
and U1448 (N_1448,N_497,N_724);
nand U1449 (N_1449,N_162,N_269);
nor U1450 (N_1450,N_921,N_706);
and U1451 (N_1451,N_657,N_7);
and U1452 (N_1452,N_394,N_730);
and U1453 (N_1453,N_722,N_395);
nor U1454 (N_1454,N_200,N_650);
nand U1455 (N_1455,N_242,N_218);
nor U1456 (N_1456,N_407,N_496);
nand U1457 (N_1457,N_499,N_123);
and U1458 (N_1458,N_513,N_464);
and U1459 (N_1459,N_761,N_48);
nor U1460 (N_1460,N_927,N_24);
or U1461 (N_1461,N_292,N_553);
and U1462 (N_1462,N_622,N_1);
and U1463 (N_1463,N_351,N_920);
or U1464 (N_1464,N_36,N_745);
and U1465 (N_1465,N_544,N_541);
nand U1466 (N_1466,N_450,N_754);
or U1467 (N_1467,N_719,N_972);
nand U1468 (N_1468,N_517,N_751);
nor U1469 (N_1469,N_92,N_4);
or U1470 (N_1470,N_640,N_812);
and U1471 (N_1471,N_478,N_934);
nor U1472 (N_1472,N_845,N_736);
and U1473 (N_1473,N_346,N_378);
and U1474 (N_1474,N_65,N_527);
and U1475 (N_1475,N_850,N_52);
and U1476 (N_1476,N_803,N_406);
and U1477 (N_1477,N_805,N_615);
nand U1478 (N_1478,N_390,N_878);
nor U1479 (N_1479,N_345,N_647);
and U1480 (N_1480,N_825,N_976);
and U1481 (N_1481,N_674,N_206);
and U1482 (N_1482,N_426,N_179);
or U1483 (N_1483,N_856,N_698);
nand U1484 (N_1484,N_472,N_554);
and U1485 (N_1485,N_867,N_566);
and U1486 (N_1486,N_727,N_784);
or U1487 (N_1487,N_157,N_808);
nand U1488 (N_1488,N_624,N_64);
or U1489 (N_1489,N_763,N_435);
or U1490 (N_1490,N_15,N_836);
nand U1491 (N_1491,N_6,N_474);
and U1492 (N_1492,N_222,N_720);
and U1493 (N_1493,N_955,N_357);
or U1494 (N_1494,N_454,N_575);
nor U1495 (N_1495,N_712,N_321);
and U1496 (N_1496,N_324,N_548);
and U1497 (N_1497,N_50,N_11);
and U1498 (N_1498,N_85,N_12);
nor U1499 (N_1499,N_310,N_448);
and U1500 (N_1500,N_177,N_731);
nor U1501 (N_1501,N_655,N_443);
nor U1502 (N_1502,N_504,N_615);
nand U1503 (N_1503,N_971,N_430);
or U1504 (N_1504,N_130,N_654);
or U1505 (N_1505,N_363,N_892);
nor U1506 (N_1506,N_393,N_545);
or U1507 (N_1507,N_196,N_448);
nor U1508 (N_1508,N_638,N_39);
and U1509 (N_1509,N_192,N_657);
nor U1510 (N_1510,N_949,N_317);
nand U1511 (N_1511,N_124,N_808);
nand U1512 (N_1512,N_582,N_5);
or U1513 (N_1513,N_318,N_268);
and U1514 (N_1514,N_798,N_380);
nor U1515 (N_1515,N_642,N_293);
and U1516 (N_1516,N_540,N_266);
nand U1517 (N_1517,N_479,N_0);
or U1518 (N_1518,N_413,N_566);
and U1519 (N_1519,N_209,N_180);
nand U1520 (N_1520,N_597,N_707);
or U1521 (N_1521,N_855,N_512);
nand U1522 (N_1522,N_395,N_820);
and U1523 (N_1523,N_326,N_967);
nand U1524 (N_1524,N_56,N_587);
and U1525 (N_1525,N_871,N_337);
and U1526 (N_1526,N_496,N_3);
nand U1527 (N_1527,N_975,N_206);
or U1528 (N_1528,N_524,N_267);
or U1529 (N_1529,N_957,N_864);
nand U1530 (N_1530,N_426,N_400);
nor U1531 (N_1531,N_509,N_226);
or U1532 (N_1532,N_202,N_772);
nor U1533 (N_1533,N_528,N_625);
nand U1534 (N_1534,N_245,N_80);
and U1535 (N_1535,N_514,N_731);
nand U1536 (N_1536,N_168,N_284);
nor U1537 (N_1537,N_135,N_326);
nor U1538 (N_1538,N_410,N_397);
nor U1539 (N_1539,N_50,N_209);
or U1540 (N_1540,N_239,N_441);
and U1541 (N_1541,N_695,N_594);
nand U1542 (N_1542,N_424,N_383);
and U1543 (N_1543,N_286,N_684);
nor U1544 (N_1544,N_75,N_821);
nand U1545 (N_1545,N_1,N_175);
or U1546 (N_1546,N_843,N_874);
nand U1547 (N_1547,N_648,N_210);
and U1548 (N_1548,N_165,N_985);
nor U1549 (N_1549,N_604,N_998);
nand U1550 (N_1550,N_563,N_812);
nand U1551 (N_1551,N_208,N_955);
nor U1552 (N_1552,N_48,N_873);
nor U1553 (N_1553,N_784,N_815);
and U1554 (N_1554,N_127,N_965);
or U1555 (N_1555,N_71,N_552);
nand U1556 (N_1556,N_835,N_889);
nand U1557 (N_1557,N_873,N_182);
nor U1558 (N_1558,N_0,N_641);
nor U1559 (N_1559,N_775,N_493);
and U1560 (N_1560,N_622,N_865);
and U1561 (N_1561,N_784,N_127);
nor U1562 (N_1562,N_258,N_211);
and U1563 (N_1563,N_89,N_192);
nor U1564 (N_1564,N_525,N_126);
nand U1565 (N_1565,N_780,N_262);
or U1566 (N_1566,N_290,N_864);
or U1567 (N_1567,N_245,N_576);
and U1568 (N_1568,N_182,N_231);
nor U1569 (N_1569,N_317,N_72);
nor U1570 (N_1570,N_386,N_468);
or U1571 (N_1571,N_134,N_350);
nand U1572 (N_1572,N_282,N_942);
or U1573 (N_1573,N_39,N_172);
nor U1574 (N_1574,N_816,N_422);
or U1575 (N_1575,N_390,N_686);
or U1576 (N_1576,N_719,N_15);
nor U1577 (N_1577,N_173,N_336);
nand U1578 (N_1578,N_976,N_238);
or U1579 (N_1579,N_611,N_741);
nand U1580 (N_1580,N_924,N_872);
and U1581 (N_1581,N_927,N_405);
and U1582 (N_1582,N_422,N_659);
or U1583 (N_1583,N_996,N_972);
or U1584 (N_1584,N_784,N_497);
nand U1585 (N_1585,N_181,N_938);
xnor U1586 (N_1586,N_576,N_244);
or U1587 (N_1587,N_573,N_320);
nor U1588 (N_1588,N_56,N_825);
and U1589 (N_1589,N_556,N_621);
nor U1590 (N_1590,N_58,N_688);
and U1591 (N_1591,N_365,N_100);
nor U1592 (N_1592,N_531,N_647);
nand U1593 (N_1593,N_290,N_939);
nor U1594 (N_1594,N_656,N_471);
nand U1595 (N_1595,N_121,N_65);
or U1596 (N_1596,N_262,N_679);
and U1597 (N_1597,N_512,N_626);
or U1598 (N_1598,N_363,N_743);
nor U1599 (N_1599,N_413,N_572);
and U1600 (N_1600,N_34,N_80);
nor U1601 (N_1601,N_603,N_894);
and U1602 (N_1602,N_202,N_380);
nand U1603 (N_1603,N_256,N_301);
or U1604 (N_1604,N_914,N_910);
nor U1605 (N_1605,N_430,N_667);
nand U1606 (N_1606,N_46,N_393);
nor U1607 (N_1607,N_287,N_79);
nand U1608 (N_1608,N_868,N_172);
nand U1609 (N_1609,N_630,N_9);
and U1610 (N_1610,N_558,N_73);
or U1611 (N_1611,N_350,N_235);
nand U1612 (N_1612,N_538,N_345);
xor U1613 (N_1613,N_215,N_866);
or U1614 (N_1614,N_415,N_4);
and U1615 (N_1615,N_255,N_966);
or U1616 (N_1616,N_940,N_337);
xnor U1617 (N_1617,N_524,N_713);
nor U1618 (N_1618,N_772,N_549);
and U1619 (N_1619,N_51,N_968);
nand U1620 (N_1620,N_218,N_631);
or U1621 (N_1621,N_713,N_228);
nor U1622 (N_1622,N_196,N_860);
and U1623 (N_1623,N_83,N_490);
and U1624 (N_1624,N_363,N_134);
nand U1625 (N_1625,N_243,N_17);
nor U1626 (N_1626,N_495,N_103);
or U1627 (N_1627,N_145,N_367);
and U1628 (N_1628,N_880,N_694);
and U1629 (N_1629,N_67,N_580);
nor U1630 (N_1630,N_589,N_778);
or U1631 (N_1631,N_706,N_397);
and U1632 (N_1632,N_771,N_230);
nor U1633 (N_1633,N_113,N_526);
nor U1634 (N_1634,N_89,N_182);
nor U1635 (N_1635,N_432,N_972);
or U1636 (N_1636,N_73,N_710);
nor U1637 (N_1637,N_818,N_537);
and U1638 (N_1638,N_362,N_438);
nand U1639 (N_1639,N_438,N_575);
nand U1640 (N_1640,N_673,N_367);
and U1641 (N_1641,N_847,N_608);
nor U1642 (N_1642,N_231,N_781);
or U1643 (N_1643,N_139,N_924);
nor U1644 (N_1644,N_228,N_184);
and U1645 (N_1645,N_883,N_279);
xnor U1646 (N_1646,N_759,N_446);
nor U1647 (N_1647,N_868,N_921);
and U1648 (N_1648,N_140,N_574);
or U1649 (N_1649,N_341,N_326);
and U1650 (N_1650,N_158,N_29);
or U1651 (N_1651,N_591,N_443);
nand U1652 (N_1652,N_805,N_785);
nor U1653 (N_1653,N_849,N_244);
and U1654 (N_1654,N_115,N_375);
and U1655 (N_1655,N_791,N_907);
or U1656 (N_1656,N_387,N_582);
nand U1657 (N_1657,N_725,N_737);
and U1658 (N_1658,N_770,N_929);
or U1659 (N_1659,N_428,N_94);
nor U1660 (N_1660,N_416,N_227);
and U1661 (N_1661,N_754,N_674);
or U1662 (N_1662,N_104,N_337);
nand U1663 (N_1663,N_871,N_403);
and U1664 (N_1664,N_449,N_829);
nand U1665 (N_1665,N_197,N_61);
or U1666 (N_1666,N_437,N_537);
or U1667 (N_1667,N_852,N_433);
nor U1668 (N_1668,N_301,N_375);
nor U1669 (N_1669,N_385,N_880);
nor U1670 (N_1670,N_580,N_363);
nand U1671 (N_1671,N_765,N_272);
and U1672 (N_1672,N_324,N_831);
or U1673 (N_1673,N_254,N_654);
nor U1674 (N_1674,N_151,N_267);
and U1675 (N_1675,N_862,N_956);
nand U1676 (N_1676,N_161,N_288);
or U1677 (N_1677,N_370,N_187);
or U1678 (N_1678,N_292,N_787);
nand U1679 (N_1679,N_362,N_599);
nor U1680 (N_1680,N_602,N_935);
nand U1681 (N_1681,N_355,N_384);
nand U1682 (N_1682,N_827,N_466);
nor U1683 (N_1683,N_616,N_895);
nor U1684 (N_1684,N_33,N_558);
and U1685 (N_1685,N_149,N_611);
and U1686 (N_1686,N_126,N_55);
nor U1687 (N_1687,N_116,N_758);
or U1688 (N_1688,N_70,N_88);
nor U1689 (N_1689,N_451,N_702);
nand U1690 (N_1690,N_4,N_407);
nand U1691 (N_1691,N_717,N_557);
or U1692 (N_1692,N_980,N_138);
nand U1693 (N_1693,N_241,N_862);
nor U1694 (N_1694,N_929,N_651);
nor U1695 (N_1695,N_678,N_542);
nor U1696 (N_1696,N_726,N_262);
nor U1697 (N_1697,N_250,N_72);
nor U1698 (N_1698,N_899,N_268);
and U1699 (N_1699,N_360,N_489);
or U1700 (N_1700,N_603,N_11);
and U1701 (N_1701,N_58,N_502);
or U1702 (N_1702,N_400,N_450);
or U1703 (N_1703,N_491,N_518);
nor U1704 (N_1704,N_624,N_353);
or U1705 (N_1705,N_972,N_43);
nand U1706 (N_1706,N_283,N_719);
nand U1707 (N_1707,N_875,N_419);
or U1708 (N_1708,N_809,N_429);
nand U1709 (N_1709,N_395,N_657);
or U1710 (N_1710,N_957,N_654);
nand U1711 (N_1711,N_939,N_504);
or U1712 (N_1712,N_155,N_545);
and U1713 (N_1713,N_703,N_942);
nor U1714 (N_1714,N_838,N_407);
and U1715 (N_1715,N_792,N_433);
nor U1716 (N_1716,N_657,N_685);
nor U1717 (N_1717,N_37,N_857);
nor U1718 (N_1718,N_0,N_991);
or U1719 (N_1719,N_622,N_129);
nor U1720 (N_1720,N_37,N_996);
nor U1721 (N_1721,N_719,N_999);
nand U1722 (N_1722,N_387,N_912);
nor U1723 (N_1723,N_406,N_151);
and U1724 (N_1724,N_150,N_395);
and U1725 (N_1725,N_530,N_395);
nor U1726 (N_1726,N_988,N_607);
and U1727 (N_1727,N_377,N_456);
or U1728 (N_1728,N_869,N_244);
nor U1729 (N_1729,N_844,N_443);
nand U1730 (N_1730,N_52,N_363);
nor U1731 (N_1731,N_251,N_228);
nand U1732 (N_1732,N_884,N_400);
nand U1733 (N_1733,N_965,N_889);
nor U1734 (N_1734,N_790,N_425);
or U1735 (N_1735,N_458,N_774);
and U1736 (N_1736,N_353,N_145);
nor U1737 (N_1737,N_979,N_12);
nor U1738 (N_1738,N_472,N_948);
or U1739 (N_1739,N_298,N_900);
nor U1740 (N_1740,N_428,N_833);
or U1741 (N_1741,N_470,N_899);
or U1742 (N_1742,N_640,N_53);
nand U1743 (N_1743,N_136,N_472);
nand U1744 (N_1744,N_501,N_486);
nand U1745 (N_1745,N_778,N_375);
nand U1746 (N_1746,N_456,N_996);
nand U1747 (N_1747,N_403,N_358);
nor U1748 (N_1748,N_962,N_419);
and U1749 (N_1749,N_395,N_582);
and U1750 (N_1750,N_792,N_699);
nand U1751 (N_1751,N_445,N_353);
nand U1752 (N_1752,N_24,N_164);
nor U1753 (N_1753,N_232,N_931);
nand U1754 (N_1754,N_471,N_452);
nor U1755 (N_1755,N_381,N_899);
or U1756 (N_1756,N_110,N_810);
or U1757 (N_1757,N_437,N_617);
nor U1758 (N_1758,N_642,N_540);
nor U1759 (N_1759,N_342,N_332);
nand U1760 (N_1760,N_789,N_551);
or U1761 (N_1761,N_669,N_601);
and U1762 (N_1762,N_58,N_797);
nor U1763 (N_1763,N_387,N_663);
nor U1764 (N_1764,N_661,N_719);
nand U1765 (N_1765,N_811,N_334);
nand U1766 (N_1766,N_606,N_13);
nand U1767 (N_1767,N_973,N_257);
nor U1768 (N_1768,N_872,N_711);
nor U1769 (N_1769,N_311,N_468);
xor U1770 (N_1770,N_186,N_414);
or U1771 (N_1771,N_9,N_85);
nor U1772 (N_1772,N_80,N_938);
or U1773 (N_1773,N_404,N_512);
nand U1774 (N_1774,N_864,N_333);
nand U1775 (N_1775,N_532,N_420);
or U1776 (N_1776,N_928,N_480);
or U1777 (N_1777,N_391,N_261);
nor U1778 (N_1778,N_230,N_691);
nand U1779 (N_1779,N_621,N_337);
and U1780 (N_1780,N_86,N_382);
or U1781 (N_1781,N_772,N_764);
or U1782 (N_1782,N_184,N_224);
nor U1783 (N_1783,N_439,N_455);
or U1784 (N_1784,N_621,N_684);
nor U1785 (N_1785,N_316,N_305);
and U1786 (N_1786,N_996,N_888);
and U1787 (N_1787,N_5,N_377);
and U1788 (N_1788,N_690,N_520);
or U1789 (N_1789,N_527,N_208);
and U1790 (N_1790,N_819,N_931);
or U1791 (N_1791,N_653,N_146);
or U1792 (N_1792,N_55,N_841);
nand U1793 (N_1793,N_759,N_423);
nand U1794 (N_1794,N_849,N_270);
or U1795 (N_1795,N_457,N_218);
nor U1796 (N_1796,N_609,N_911);
or U1797 (N_1797,N_968,N_397);
or U1798 (N_1798,N_390,N_527);
nand U1799 (N_1799,N_512,N_679);
nor U1800 (N_1800,N_524,N_83);
and U1801 (N_1801,N_965,N_818);
or U1802 (N_1802,N_515,N_927);
or U1803 (N_1803,N_63,N_9);
or U1804 (N_1804,N_771,N_958);
and U1805 (N_1805,N_294,N_430);
nor U1806 (N_1806,N_90,N_624);
nand U1807 (N_1807,N_471,N_344);
nor U1808 (N_1808,N_634,N_442);
or U1809 (N_1809,N_20,N_283);
and U1810 (N_1810,N_783,N_129);
nand U1811 (N_1811,N_936,N_207);
and U1812 (N_1812,N_492,N_755);
nor U1813 (N_1813,N_941,N_856);
and U1814 (N_1814,N_211,N_592);
nor U1815 (N_1815,N_847,N_784);
or U1816 (N_1816,N_873,N_568);
and U1817 (N_1817,N_359,N_40);
nand U1818 (N_1818,N_935,N_628);
nor U1819 (N_1819,N_648,N_73);
or U1820 (N_1820,N_698,N_828);
nand U1821 (N_1821,N_153,N_44);
and U1822 (N_1822,N_762,N_650);
or U1823 (N_1823,N_617,N_821);
nand U1824 (N_1824,N_724,N_977);
nand U1825 (N_1825,N_413,N_550);
or U1826 (N_1826,N_717,N_549);
nor U1827 (N_1827,N_863,N_321);
nor U1828 (N_1828,N_463,N_904);
or U1829 (N_1829,N_349,N_555);
nand U1830 (N_1830,N_982,N_203);
nor U1831 (N_1831,N_13,N_567);
or U1832 (N_1832,N_496,N_951);
nand U1833 (N_1833,N_452,N_654);
or U1834 (N_1834,N_337,N_440);
and U1835 (N_1835,N_591,N_282);
xnor U1836 (N_1836,N_831,N_466);
or U1837 (N_1837,N_310,N_523);
nand U1838 (N_1838,N_418,N_908);
and U1839 (N_1839,N_795,N_728);
and U1840 (N_1840,N_641,N_417);
or U1841 (N_1841,N_652,N_191);
nor U1842 (N_1842,N_466,N_498);
nand U1843 (N_1843,N_849,N_718);
nand U1844 (N_1844,N_12,N_420);
and U1845 (N_1845,N_218,N_19);
nor U1846 (N_1846,N_597,N_172);
nand U1847 (N_1847,N_891,N_441);
or U1848 (N_1848,N_662,N_440);
nor U1849 (N_1849,N_986,N_700);
or U1850 (N_1850,N_623,N_285);
or U1851 (N_1851,N_882,N_325);
nor U1852 (N_1852,N_752,N_142);
nand U1853 (N_1853,N_432,N_983);
nand U1854 (N_1854,N_883,N_854);
or U1855 (N_1855,N_872,N_211);
nor U1856 (N_1856,N_310,N_227);
nand U1857 (N_1857,N_885,N_664);
nor U1858 (N_1858,N_322,N_232);
nand U1859 (N_1859,N_638,N_9);
or U1860 (N_1860,N_617,N_606);
or U1861 (N_1861,N_965,N_492);
and U1862 (N_1862,N_342,N_441);
and U1863 (N_1863,N_538,N_574);
nor U1864 (N_1864,N_651,N_777);
or U1865 (N_1865,N_491,N_515);
nor U1866 (N_1866,N_501,N_966);
and U1867 (N_1867,N_500,N_233);
and U1868 (N_1868,N_313,N_426);
nor U1869 (N_1869,N_512,N_746);
nor U1870 (N_1870,N_815,N_18);
xor U1871 (N_1871,N_952,N_117);
or U1872 (N_1872,N_997,N_88);
nand U1873 (N_1873,N_889,N_460);
nand U1874 (N_1874,N_638,N_647);
nand U1875 (N_1875,N_163,N_465);
or U1876 (N_1876,N_92,N_488);
nor U1877 (N_1877,N_455,N_839);
nand U1878 (N_1878,N_333,N_826);
and U1879 (N_1879,N_345,N_266);
nand U1880 (N_1880,N_92,N_17);
xnor U1881 (N_1881,N_596,N_726);
nand U1882 (N_1882,N_198,N_684);
or U1883 (N_1883,N_965,N_942);
nand U1884 (N_1884,N_156,N_947);
nand U1885 (N_1885,N_317,N_426);
nor U1886 (N_1886,N_586,N_74);
and U1887 (N_1887,N_286,N_493);
or U1888 (N_1888,N_833,N_246);
nor U1889 (N_1889,N_575,N_608);
and U1890 (N_1890,N_850,N_37);
nand U1891 (N_1891,N_723,N_156);
nor U1892 (N_1892,N_504,N_143);
or U1893 (N_1893,N_878,N_421);
or U1894 (N_1894,N_77,N_116);
and U1895 (N_1895,N_528,N_810);
or U1896 (N_1896,N_730,N_836);
and U1897 (N_1897,N_88,N_720);
xnor U1898 (N_1898,N_769,N_365);
nor U1899 (N_1899,N_153,N_453);
and U1900 (N_1900,N_65,N_473);
or U1901 (N_1901,N_797,N_953);
or U1902 (N_1902,N_448,N_702);
and U1903 (N_1903,N_722,N_243);
or U1904 (N_1904,N_565,N_84);
or U1905 (N_1905,N_785,N_276);
and U1906 (N_1906,N_796,N_294);
and U1907 (N_1907,N_990,N_94);
and U1908 (N_1908,N_227,N_661);
and U1909 (N_1909,N_233,N_862);
and U1910 (N_1910,N_350,N_682);
or U1911 (N_1911,N_925,N_991);
nand U1912 (N_1912,N_348,N_25);
nor U1913 (N_1913,N_335,N_679);
nor U1914 (N_1914,N_247,N_252);
or U1915 (N_1915,N_694,N_865);
nand U1916 (N_1916,N_188,N_33);
nand U1917 (N_1917,N_772,N_259);
nand U1918 (N_1918,N_329,N_459);
nand U1919 (N_1919,N_311,N_792);
or U1920 (N_1920,N_331,N_702);
and U1921 (N_1921,N_409,N_137);
nand U1922 (N_1922,N_813,N_685);
and U1923 (N_1923,N_249,N_844);
and U1924 (N_1924,N_284,N_497);
and U1925 (N_1925,N_357,N_690);
and U1926 (N_1926,N_84,N_809);
xor U1927 (N_1927,N_450,N_777);
nor U1928 (N_1928,N_801,N_150);
and U1929 (N_1929,N_166,N_580);
or U1930 (N_1930,N_378,N_324);
nand U1931 (N_1931,N_7,N_772);
and U1932 (N_1932,N_384,N_181);
nand U1933 (N_1933,N_300,N_861);
or U1934 (N_1934,N_936,N_939);
and U1935 (N_1935,N_190,N_474);
nor U1936 (N_1936,N_760,N_391);
nor U1937 (N_1937,N_566,N_379);
or U1938 (N_1938,N_684,N_791);
or U1939 (N_1939,N_896,N_645);
or U1940 (N_1940,N_846,N_307);
nand U1941 (N_1941,N_349,N_426);
nor U1942 (N_1942,N_283,N_239);
nand U1943 (N_1943,N_775,N_544);
or U1944 (N_1944,N_798,N_15);
and U1945 (N_1945,N_516,N_868);
and U1946 (N_1946,N_851,N_283);
and U1947 (N_1947,N_200,N_20);
nor U1948 (N_1948,N_197,N_811);
and U1949 (N_1949,N_136,N_830);
or U1950 (N_1950,N_516,N_568);
or U1951 (N_1951,N_374,N_599);
and U1952 (N_1952,N_218,N_71);
nor U1953 (N_1953,N_654,N_61);
or U1954 (N_1954,N_175,N_910);
nand U1955 (N_1955,N_686,N_370);
or U1956 (N_1956,N_975,N_773);
nor U1957 (N_1957,N_837,N_26);
nor U1958 (N_1958,N_269,N_856);
nand U1959 (N_1959,N_958,N_133);
and U1960 (N_1960,N_214,N_953);
and U1961 (N_1961,N_640,N_276);
nor U1962 (N_1962,N_581,N_855);
nor U1963 (N_1963,N_234,N_982);
nand U1964 (N_1964,N_517,N_663);
nand U1965 (N_1965,N_321,N_507);
nand U1966 (N_1966,N_393,N_489);
or U1967 (N_1967,N_217,N_763);
nor U1968 (N_1968,N_194,N_714);
nor U1969 (N_1969,N_648,N_145);
and U1970 (N_1970,N_744,N_413);
and U1971 (N_1971,N_409,N_740);
or U1972 (N_1972,N_640,N_572);
and U1973 (N_1973,N_296,N_192);
nand U1974 (N_1974,N_986,N_298);
and U1975 (N_1975,N_111,N_79);
nand U1976 (N_1976,N_115,N_25);
and U1977 (N_1977,N_634,N_628);
nand U1978 (N_1978,N_425,N_933);
xor U1979 (N_1979,N_577,N_255);
or U1980 (N_1980,N_274,N_22);
or U1981 (N_1981,N_807,N_537);
or U1982 (N_1982,N_738,N_875);
or U1983 (N_1983,N_10,N_258);
and U1984 (N_1984,N_904,N_317);
nand U1985 (N_1985,N_52,N_610);
nand U1986 (N_1986,N_528,N_218);
nor U1987 (N_1987,N_335,N_801);
nor U1988 (N_1988,N_666,N_166);
nand U1989 (N_1989,N_218,N_103);
and U1990 (N_1990,N_749,N_211);
nor U1991 (N_1991,N_973,N_818);
or U1992 (N_1992,N_807,N_449);
nand U1993 (N_1993,N_494,N_896);
and U1994 (N_1994,N_491,N_37);
nor U1995 (N_1995,N_219,N_25);
and U1996 (N_1996,N_651,N_375);
and U1997 (N_1997,N_490,N_942);
and U1998 (N_1998,N_649,N_730);
xor U1999 (N_1999,N_630,N_212);
and U2000 (N_2000,N_1036,N_1661);
and U2001 (N_2001,N_1308,N_1443);
or U2002 (N_2002,N_1237,N_1226);
and U2003 (N_2003,N_1204,N_1949);
nor U2004 (N_2004,N_1960,N_1235);
or U2005 (N_2005,N_1494,N_1143);
or U2006 (N_2006,N_1145,N_1472);
or U2007 (N_2007,N_1331,N_1532);
nand U2008 (N_2008,N_1455,N_1219);
nand U2009 (N_2009,N_1172,N_1840);
nand U2010 (N_2010,N_1280,N_1883);
nand U2011 (N_2011,N_1712,N_1084);
xnor U2012 (N_2012,N_1918,N_1801);
or U2013 (N_2013,N_1464,N_1909);
nand U2014 (N_2014,N_1778,N_1647);
nand U2015 (N_2015,N_1651,N_1310);
nor U2016 (N_2016,N_1147,N_1123);
or U2017 (N_2017,N_1350,N_1183);
and U2018 (N_2018,N_1868,N_1886);
nand U2019 (N_2019,N_1378,N_1466);
nor U2020 (N_2020,N_1176,N_1862);
nor U2021 (N_2021,N_1784,N_1866);
or U2022 (N_2022,N_1521,N_1323);
or U2023 (N_2023,N_1516,N_1765);
and U2024 (N_2024,N_1577,N_1001);
nand U2025 (N_2025,N_1045,N_1556);
nor U2026 (N_2026,N_1880,N_1985);
nand U2027 (N_2027,N_1065,N_1966);
and U2028 (N_2028,N_1191,N_1769);
nor U2029 (N_2029,N_1368,N_1870);
nand U2030 (N_2030,N_1160,N_1122);
and U2031 (N_2031,N_1022,N_1201);
nor U2032 (N_2032,N_1469,N_1248);
nor U2033 (N_2033,N_1621,N_1630);
nor U2034 (N_2034,N_1477,N_1366);
or U2035 (N_2035,N_1081,N_1389);
or U2036 (N_2036,N_1570,N_1066);
and U2037 (N_2037,N_1602,N_1761);
nand U2038 (N_2038,N_1328,N_1326);
and U2039 (N_2039,N_1457,N_1316);
nand U2040 (N_2040,N_1322,N_1168);
nor U2041 (N_2041,N_1076,N_1385);
nor U2042 (N_2042,N_1083,N_1749);
nand U2043 (N_2043,N_1265,N_1159);
or U2044 (N_2044,N_1380,N_1559);
or U2045 (N_2045,N_1044,N_1460);
nor U2046 (N_2046,N_1085,N_1211);
and U2047 (N_2047,N_1290,N_1436);
nand U2048 (N_2048,N_1991,N_1864);
or U2049 (N_2049,N_1161,N_1674);
nor U2050 (N_2050,N_1422,N_1774);
or U2051 (N_2051,N_1994,N_1781);
and U2052 (N_2052,N_1585,N_1246);
nor U2053 (N_2053,N_1666,N_1349);
nor U2054 (N_2054,N_1397,N_1509);
or U2055 (N_2055,N_1105,N_1024);
nand U2056 (N_2056,N_1853,N_1069);
nor U2057 (N_2057,N_1415,N_1503);
nor U2058 (N_2058,N_1701,N_1470);
or U2059 (N_2059,N_1135,N_1982);
or U2060 (N_2060,N_1106,N_1640);
nor U2061 (N_2061,N_1236,N_1110);
and U2062 (N_2062,N_1279,N_1873);
nor U2063 (N_2063,N_1905,N_1806);
nand U2064 (N_2064,N_1791,N_1244);
nand U2065 (N_2065,N_1462,N_1927);
and U2066 (N_2066,N_1283,N_1010);
or U2067 (N_2067,N_1206,N_1500);
nand U2068 (N_2068,N_1089,N_1673);
nor U2069 (N_2069,N_1860,N_1569);
nor U2070 (N_2070,N_1555,N_1216);
nor U2071 (N_2071,N_1164,N_1075);
nor U2072 (N_2072,N_1212,N_1723);
or U2073 (N_2073,N_1591,N_1009);
or U2074 (N_2074,N_1408,N_1273);
nor U2075 (N_2075,N_1895,N_1770);
nor U2076 (N_2076,N_1102,N_1600);
nor U2077 (N_2077,N_1433,N_1298);
nor U2078 (N_2078,N_1692,N_1360);
nand U2079 (N_2079,N_1534,N_1357);
and U2080 (N_2080,N_1192,N_1340);
and U2081 (N_2081,N_1245,N_1482);
nand U2082 (N_2082,N_1847,N_1973);
nor U2083 (N_2083,N_1259,N_1261);
and U2084 (N_2084,N_1867,N_1240);
or U2085 (N_2085,N_1751,N_1590);
and U2086 (N_2086,N_1238,N_1669);
and U2087 (N_2087,N_1394,N_1842);
nor U2088 (N_2088,N_1239,N_1064);
or U2089 (N_2089,N_1221,N_1314);
nor U2090 (N_2090,N_1151,N_1040);
and U2091 (N_2091,N_1764,N_1515);
nor U2092 (N_2092,N_1440,N_1499);
nor U2093 (N_2093,N_1307,N_1182);
nor U2094 (N_2094,N_1033,N_1805);
and U2095 (N_2095,N_1813,N_1554);
nor U2096 (N_2096,N_1100,N_1353);
or U2097 (N_2097,N_1605,N_1538);
nor U2098 (N_2098,N_1485,N_1525);
nor U2099 (N_2099,N_1746,N_1548);
nand U2100 (N_2100,N_1432,N_1714);
xnor U2101 (N_2101,N_1155,N_1043);
or U2102 (N_2102,N_1888,N_1984);
nor U2103 (N_2103,N_1533,N_1344);
nand U2104 (N_2104,N_1288,N_1969);
or U2105 (N_2105,N_1333,N_1233);
or U2106 (N_2106,N_1507,N_1463);
or U2107 (N_2107,N_1289,N_1291);
and U2108 (N_2108,N_1171,N_1592);
nand U2109 (N_2109,N_1018,N_1465);
nand U2110 (N_2110,N_1094,N_1384);
or U2111 (N_2111,N_1109,N_1926);
or U2112 (N_2112,N_1120,N_1752);
nor U2113 (N_2113,N_1179,N_1073);
nor U2114 (N_2114,N_1149,N_1890);
and U2115 (N_2115,N_1272,N_1718);
or U2116 (N_2116,N_1613,N_1413);
or U2117 (N_2117,N_1940,N_1048);
and U2118 (N_2118,N_1373,N_1406);
and U2119 (N_2119,N_1262,N_1971);
and U2120 (N_2120,N_1919,N_1101);
or U2121 (N_2121,N_1028,N_1923);
nand U2122 (N_2122,N_1524,N_1996);
nand U2123 (N_2123,N_1039,N_1404);
nand U2124 (N_2124,N_1762,N_1691);
or U2125 (N_2125,N_1557,N_1875);
nor U2126 (N_2126,N_1623,N_1364);
nor U2127 (N_2127,N_1027,N_1187);
nand U2128 (N_2128,N_1127,N_1839);
or U2129 (N_2129,N_1136,N_1471);
nand U2130 (N_2130,N_1553,N_1427);
and U2131 (N_2131,N_1650,N_1197);
nor U2132 (N_2132,N_1810,N_1777);
or U2133 (N_2133,N_1584,N_1872);
nor U2134 (N_2134,N_1059,N_1648);
nand U2135 (N_2135,N_1811,N_1278);
nand U2136 (N_2136,N_1739,N_1572);
and U2137 (N_2137,N_1632,N_1410);
and U2138 (N_2138,N_1831,N_1479);
and U2139 (N_2139,N_1727,N_1906);
nand U2140 (N_2140,N_1792,N_1571);
nor U2141 (N_2141,N_1067,N_1337);
nor U2142 (N_2142,N_1374,N_1999);
and U2143 (N_2143,N_1270,N_1948);
and U2144 (N_2144,N_1946,N_1299);
nand U2145 (N_2145,N_1797,N_1203);
or U2146 (N_2146,N_1823,N_1678);
nor U2147 (N_2147,N_1351,N_1476);
nand U2148 (N_2148,N_1858,N_1582);
nor U2149 (N_2149,N_1051,N_1997);
and U2150 (N_2150,N_1950,N_1473);
and U2151 (N_2151,N_1829,N_1565);
nor U2152 (N_2152,N_1983,N_1871);
or U2153 (N_2153,N_1167,N_1011);
nand U2154 (N_2154,N_1733,N_1990);
nor U2155 (N_2155,N_1795,N_1091);
and U2156 (N_2156,N_1504,N_1398);
and U2157 (N_2157,N_1779,N_1185);
or U2158 (N_2158,N_1581,N_1690);
nor U2159 (N_2159,N_1421,N_1268);
or U2160 (N_2160,N_1070,N_1250);
or U2161 (N_2161,N_1638,N_1367);
nor U2162 (N_2162,N_1717,N_1814);
nor U2163 (N_2163,N_1744,N_1552);
and U2164 (N_2164,N_1841,N_1058);
nand U2165 (N_2165,N_1859,N_1227);
nand U2166 (N_2166,N_1134,N_1937);
or U2167 (N_2167,N_1052,N_1330);
nor U2168 (N_2168,N_1411,N_1908);
nand U2169 (N_2169,N_1843,N_1992);
nand U2170 (N_2170,N_1738,N_1610);
and U2171 (N_2171,N_1720,N_1498);
or U2172 (N_2172,N_1945,N_1297);
and U2173 (N_2173,N_1785,N_1451);
nand U2174 (N_2174,N_1523,N_1327);
nor U2175 (N_2175,N_1150,N_1713);
or U2176 (N_2176,N_1885,N_1579);
or U2177 (N_2177,N_1153,N_1832);
or U2178 (N_2178,N_1818,N_1856);
or U2179 (N_2179,N_1562,N_1920);
or U2180 (N_2180,N_1266,N_1865);
or U2181 (N_2181,N_1511,N_1144);
and U2182 (N_2182,N_1311,N_1074);
nor U2183 (N_2183,N_1332,N_1205);
and U2184 (N_2184,N_1978,N_1108);
nor U2185 (N_2185,N_1126,N_1583);
and U2186 (N_2186,N_1693,N_1726);
nand U2187 (N_2187,N_1295,N_1077);
and U2188 (N_2188,N_1348,N_1133);
and U2189 (N_2189,N_1838,N_1060);
nor U2190 (N_2190,N_1376,N_1213);
or U2191 (N_2191,N_1611,N_1169);
nor U2192 (N_2192,N_1200,N_1459);
and U2193 (N_2193,N_1104,N_1467);
or U2194 (N_2194,N_1345,N_1399);
and U2195 (N_2195,N_1484,N_1597);
and U2196 (N_2196,N_1038,N_1241);
and U2197 (N_2197,N_1644,N_1125);
nor U2198 (N_2198,N_1697,N_1852);
or U2199 (N_2199,N_1708,N_1363);
and U2200 (N_2200,N_1252,N_1755);
nor U2201 (N_2201,N_1961,N_1229);
nor U2202 (N_2202,N_1452,N_1596);
nand U2203 (N_2203,N_1857,N_1281);
or U2204 (N_2204,N_1882,N_1822);
and U2205 (N_2205,N_1341,N_1177);
nor U2206 (N_2206,N_1401,N_1963);
nand U2207 (N_2207,N_1189,N_1114);
nor U2208 (N_2208,N_1220,N_1707);
nand U2209 (N_2209,N_1913,N_1416);
nor U2210 (N_2210,N_1218,N_1124);
and U2211 (N_2211,N_1531,N_1851);
nor U2212 (N_2212,N_1371,N_1400);
or U2213 (N_2213,N_1137,N_1113);
or U2214 (N_2214,N_1014,N_1446);
nand U2215 (N_2215,N_1274,N_1276);
nand U2216 (N_2216,N_1492,N_1506);
and U2217 (N_2217,N_1293,N_1305);
nand U2218 (N_2218,N_1403,N_1501);
nor U2219 (N_2219,N_1257,N_1685);
or U2220 (N_2220,N_1512,N_1668);
and U2221 (N_2221,N_1624,N_1362);
nor U2222 (N_2222,N_1407,N_1098);
or U2223 (N_2223,N_1988,N_1780);
and U2224 (N_2224,N_1753,N_1931);
nor U2225 (N_2225,N_1437,N_1116);
nand U2226 (N_2226,N_1645,N_1893);
nand U2227 (N_2227,N_1119,N_1315);
and U2228 (N_2228,N_1008,N_1628);
nand U2229 (N_2229,N_1223,N_1099);
nor U2230 (N_2230,N_1794,N_1951);
nor U2231 (N_2231,N_1646,N_1256);
nand U2232 (N_2232,N_1772,N_1210);
and U2233 (N_2233,N_1734,N_1952);
nor U2234 (N_2234,N_1339,N_1031);
nor U2235 (N_2235,N_1750,N_1546);
nor U2236 (N_2236,N_1877,N_1545);
nor U2237 (N_2237,N_1998,N_1202);
and U2238 (N_2238,N_1230,N_1529);
and U2239 (N_2239,N_1514,N_1361);
or U2240 (N_2240,N_1728,N_1030);
nor U2241 (N_2241,N_1224,N_1194);
and U2242 (N_2242,N_1543,N_1830);
nor U2243 (N_2243,N_1193,N_1391);
and U2244 (N_2244,N_1370,N_1497);
or U2245 (N_2245,N_1510,N_1542);
nor U2246 (N_2246,N_1037,N_1286);
or U2247 (N_2247,N_1309,N_1652);
nand U2248 (N_2248,N_1802,N_1003);
xnor U2249 (N_2249,N_1130,N_1625);
or U2250 (N_2250,N_1879,N_1547);
nor U2251 (N_2251,N_1993,N_1115);
and U2252 (N_2252,N_1891,N_1000);
nor U2253 (N_2253,N_1863,N_1696);
and U2254 (N_2254,N_1488,N_1771);
nor U2255 (N_2255,N_1522,N_1705);
nand U2256 (N_2256,N_1812,N_1747);
or U2257 (N_2257,N_1026,N_1836);
nand U2258 (N_2258,N_1884,N_1251);
nand U2259 (N_2259,N_1953,N_1317);
nand U2260 (N_2260,N_1354,N_1664);
and U2261 (N_2261,N_1986,N_1178);
nor U2262 (N_2262,N_1980,N_1844);
or U2263 (N_2263,N_1916,N_1017);
nor U2264 (N_2264,N_1020,N_1783);
or U2265 (N_2265,N_1215,N_1915);
and U2266 (N_2266,N_1209,N_1263);
and U2267 (N_2267,N_1958,N_1336);
nor U2268 (N_2268,N_1053,N_1063);
and U2269 (N_2269,N_1242,N_1379);
nor U2270 (N_2270,N_1910,N_1535);
or U2271 (N_2271,N_1558,N_1775);
nor U2272 (N_2272,N_1152,N_1604);
and U2273 (N_2273,N_1047,N_1972);
or U2274 (N_2274,N_1835,N_1264);
nor U2275 (N_2275,N_1505,N_1869);
nand U2276 (N_2276,N_1850,N_1313);
nand U2277 (N_2277,N_1899,N_1711);
or U2278 (N_2278,N_1166,N_1878);
nand U2279 (N_2279,N_1682,N_1679);
and U2280 (N_2280,N_1414,N_1025);
and U2281 (N_2281,N_1759,N_1392);
or U2282 (N_2282,N_1184,N_1658);
nor U2283 (N_2283,N_1903,N_1006);
or U2284 (N_2284,N_1402,N_1247);
nand U2285 (N_2285,N_1849,N_1825);
and U2286 (N_2286,N_1737,N_1382);
nand U2287 (N_2287,N_1249,N_1627);
nor U2288 (N_2288,N_1491,N_1444);
nor U2289 (N_2289,N_1355,N_1170);
nand U2290 (N_2290,N_1418,N_1208);
nand U2291 (N_2291,N_1243,N_1320);
or U2292 (N_2292,N_1222,N_1438);
or U2293 (N_2293,N_1260,N_1933);
xnor U2294 (N_2294,N_1082,N_1277);
nand U2295 (N_2295,N_1944,N_1925);
nand U2296 (N_2296,N_1942,N_1359);
nand U2297 (N_2297,N_1095,N_1618);
or U2298 (N_2298,N_1163,N_1269);
nor U2299 (N_2299,N_1448,N_1453);
and U2300 (N_2300,N_1921,N_1938);
nor U2301 (N_2301,N_1688,N_1267);
or U2302 (N_2302,N_1588,N_1072);
nor U2303 (N_2303,N_1670,N_1090);
and U2304 (N_2304,N_1458,N_1007);
nand U2305 (N_2305,N_1536,N_1544);
and U2306 (N_2306,N_1776,N_1729);
or U2307 (N_2307,N_1703,N_1757);
and U2308 (N_2308,N_1663,N_1741);
nor U2309 (N_2309,N_1481,N_1773);
or U2310 (N_2310,N_1325,N_1056);
nand U2311 (N_2311,N_1656,N_1405);
nor U2312 (N_2312,N_1660,N_1657);
nand U2313 (N_2313,N_1032,N_1725);
and U2314 (N_2314,N_1939,N_1549);
or U2315 (N_2315,N_1846,N_1156);
nand U2316 (N_2316,N_1616,N_1180);
and U2317 (N_2317,N_1107,N_1140);
nor U2318 (N_2318,N_1900,N_1306);
nor U2319 (N_2319,N_1981,N_1907);
and U2320 (N_2320,N_1480,N_1987);
or U2321 (N_2321,N_1055,N_1409);
or U2322 (N_2322,N_1287,N_1489);
or U2323 (N_2323,N_1977,N_1803);
and U2324 (N_2324,N_1381,N_1589);
nor U2325 (N_2325,N_1807,N_1282);
nor U2326 (N_2326,N_1898,N_1587);
nand U2327 (N_2327,N_1365,N_1275);
nor U2328 (N_2328,N_1386,N_1198);
and U2329 (N_2329,N_1347,N_1428);
nand U2330 (N_2330,N_1911,N_1786);
nor U2331 (N_2331,N_1112,N_1478);
and U2332 (N_2332,N_1930,N_1672);
nor U2333 (N_2333,N_1148,N_1121);
nor U2334 (N_2334,N_1196,N_1606);
or U2335 (N_2335,N_1580,N_1955);
nor U2336 (N_2336,N_1526,N_1425);
nand U2337 (N_2337,N_1303,N_1637);
and U2338 (N_2338,N_1800,N_1162);
nand U2339 (N_2339,N_1541,N_1093);
or U2340 (N_2340,N_1896,N_1019);
nor U2341 (N_2341,N_1012,N_1550);
nand U2342 (N_2342,N_1285,N_1833);
and U2343 (N_2343,N_1540,N_1808);
nand U2344 (N_2344,N_1894,N_1730);
and U2345 (N_2345,N_1924,N_1490);
nor U2346 (N_2346,N_1861,N_1612);
nand U2347 (N_2347,N_1486,N_1643);
nor U2348 (N_2348,N_1042,N_1848);
or U2349 (N_2349,N_1487,N_1854);
or U2350 (N_2350,N_1787,N_1461);
nor U2351 (N_2351,N_1573,N_1046);
or U2352 (N_2352,N_1254,N_1129);
and U2353 (N_2353,N_1342,N_1175);
nand U2354 (N_2354,N_1041,N_1225);
and U2355 (N_2355,N_1343,N_1702);
and U2356 (N_2356,N_1564,N_1518);
xor U2357 (N_2357,N_1493,N_1214);
nand U2358 (N_2358,N_1804,N_1423);
and U2359 (N_2359,N_1876,N_1447);
and U2360 (N_2360,N_1767,N_1396);
nor U2361 (N_2361,N_1968,N_1654);
or U2362 (N_2362,N_1527,N_1614);
and U2363 (N_2363,N_1642,N_1683);
and U2364 (N_2364,N_1721,N_1424);
or U2365 (N_2365,N_1659,N_1731);
or U2366 (N_2366,N_1329,N_1782);
or U2367 (N_2367,N_1092,N_1681);
and U2368 (N_2368,N_1594,N_1190);
or U2369 (N_2369,N_1595,N_1141);
or U2370 (N_2370,N_1956,N_1002);
nor U2371 (N_2371,N_1680,N_1551);
nand U2372 (N_2372,N_1566,N_1821);
nor U2373 (N_2373,N_1917,N_1560);
or U2374 (N_2374,N_1495,N_1417);
nor U2375 (N_2375,N_1947,N_1964);
nand U2376 (N_2376,N_1352,N_1071);
nor U2377 (N_2377,N_1724,N_1483);
xor U2378 (N_2378,N_1304,N_1902);
nor U2379 (N_2379,N_1431,N_1671);
nand U2380 (N_2380,N_1965,N_1517);
or U2381 (N_2381,N_1271,N_1537);
or U2382 (N_2382,N_1631,N_1128);
nor U2383 (N_2383,N_1686,N_1334);
or U2384 (N_2384,N_1034,N_1441);
nor U2385 (N_2385,N_1146,N_1928);
nand U2386 (N_2386,N_1016,N_1439);
nand U2387 (N_2387,N_1454,N_1513);
nand U2388 (N_2388,N_1619,N_1633);
nor U2389 (N_2389,N_1608,N_1819);
or U2390 (N_2390,N_1388,N_1302);
or U2391 (N_2391,N_1798,N_1706);
nand U2392 (N_2392,N_1475,N_1598);
and U2393 (N_2393,N_1111,N_1929);
nand U2394 (N_2394,N_1817,N_1607);
and U2395 (N_2395,N_1695,N_1601);
and U2396 (N_2396,N_1232,N_1837);
nand U2397 (N_2397,N_1228,N_1743);
or U2398 (N_2398,N_1957,N_1442);
or U2399 (N_2399,N_1173,N_1676);
or U2400 (N_2400,N_1599,N_1375);
nand U2401 (N_2401,N_1586,N_1827);
or U2402 (N_2402,N_1881,N_1062);
nor U2403 (N_2403,N_1207,N_1258);
and U2404 (N_2404,N_1335,N_1346);
nand U2405 (N_2405,N_1689,N_1117);
nand U2406 (N_2406,N_1138,N_1698);
nor U2407 (N_2407,N_1790,N_1296);
nor U2408 (N_2408,N_1449,N_1383);
nand U2409 (N_2409,N_1429,N_1975);
nand U2410 (N_2410,N_1634,N_1165);
or U2411 (N_2411,N_1292,N_1892);
and U2412 (N_2412,N_1004,N_1217);
or U2413 (N_2413,N_1426,N_1576);
nor U2414 (N_2414,N_1539,N_1815);
and U2415 (N_2415,N_1834,N_1393);
and U2416 (N_2416,N_1430,N_1434);
and U2417 (N_2417,N_1096,N_1321);
nor U2418 (N_2418,N_1530,N_1231);
or U2419 (N_2419,N_1620,N_1561);
and U2420 (N_2420,N_1061,N_1057);
nand U2421 (N_2421,N_1300,N_1356);
or U2422 (N_2422,N_1722,N_1029);
nor U2423 (N_2423,N_1284,N_1901);
or U2424 (N_2424,N_1760,N_1694);
nor U2425 (N_2425,N_1174,N_1845);
nand U2426 (N_2426,N_1474,N_1914);
or U2427 (N_2427,N_1758,N_1622);
nor U2428 (N_2428,N_1742,N_1740);
nand U2429 (N_2429,N_1828,N_1035);
nor U2430 (N_2430,N_1567,N_1704);
or U2431 (N_2431,N_1677,N_1142);
or U2432 (N_2432,N_1954,N_1528);
nand U2433 (N_2433,N_1390,N_1395);
and U2434 (N_2434,N_1502,N_1932);
nor U2435 (N_2435,N_1412,N_1979);
and U2436 (N_2436,N_1736,N_1234);
nand U2437 (N_2437,N_1756,N_1088);
nand U2438 (N_2438,N_1639,N_1897);
nand U2439 (N_2439,N_1763,N_1719);
nand U2440 (N_2440,N_1078,N_1626);
nand U2441 (N_2441,N_1976,N_1103);
or U2442 (N_2442,N_1824,N_1575);
or U2443 (N_2443,N_1735,N_1974);
nand U2444 (N_2444,N_1675,N_1609);
or U2445 (N_2445,N_1732,N_1387);
nand U2446 (N_2446,N_1377,N_1793);
nand U2447 (N_2447,N_1809,N_1989);
nand U2448 (N_2448,N_1338,N_1684);
and U2449 (N_2449,N_1603,N_1301);
or U2450 (N_2450,N_1080,N_1157);
and U2451 (N_2451,N_1635,N_1716);
nand U2452 (N_2452,N_1943,N_1520);
nor U2453 (N_2453,N_1420,N_1023);
nand U2454 (N_2454,N_1699,N_1139);
nand U2455 (N_2455,N_1874,N_1312);
and U2456 (N_2456,N_1687,N_1068);
nor U2457 (N_2457,N_1855,N_1959);
nand U2458 (N_2458,N_1049,N_1054);
nand U2459 (N_2459,N_1294,N_1912);
or U2460 (N_2460,N_1419,N_1629);
or U2461 (N_2461,N_1995,N_1131);
nand U2462 (N_2462,N_1941,N_1887);
nand U2463 (N_2463,N_1050,N_1253);
and U2464 (N_2464,N_1021,N_1715);
and U2465 (N_2465,N_1086,N_1496);
nand U2466 (N_2466,N_1636,N_1788);
nand U2467 (N_2467,N_1700,N_1641);
or U2468 (N_2468,N_1745,N_1934);
nand U2469 (N_2469,N_1186,N_1967);
nand U2470 (N_2470,N_1665,N_1662);
or U2471 (N_2471,N_1255,N_1369);
and U2472 (N_2472,N_1132,N_1319);
nor U2473 (N_2473,N_1936,N_1748);
nand U2474 (N_2474,N_1158,N_1005);
nor U2475 (N_2475,N_1796,N_1456);
nor U2476 (N_2476,N_1593,N_1962);
and U2477 (N_2477,N_1709,N_1154);
nor U2478 (N_2478,N_1655,N_1445);
and U2479 (N_2479,N_1617,N_1820);
and U2480 (N_2480,N_1816,N_1889);
and U2481 (N_2481,N_1789,N_1199);
nand U2482 (N_2482,N_1574,N_1097);
nand U2483 (N_2483,N_1766,N_1615);
and U2484 (N_2484,N_1450,N_1768);
or U2485 (N_2485,N_1318,N_1935);
or U2486 (N_2486,N_1435,N_1667);
nor U2487 (N_2487,N_1970,N_1324);
nor U2488 (N_2488,N_1649,N_1754);
and U2489 (N_2489,N_1508,N_1118);
and U2490 (N_2490,N_1013,N_1519);
nor U2491 (N_2491,N_1195,N_1710);
and U2492 (N_2492,N_1079,N_1826);
and U2493 (N_2493,N_1653,N_1922);
and U2494 (N_2494,N_1087,N_1563);
and U2495 (N_2495,N_1372,N_1904);
and U2496 (N_2496,N_1468,N_1568);
nand U2497 (N_2497,N_1015,N_1799);
nand U2498 (N_2498,N_1578,N_1181);
and U2499 (N_2499,N_1188,N_1358);
or U2500 (N_2500,N_1765,N_1281);
nand U2501 (N_2501,N_1689,N_1010);
and U2502 (N_2502,N_1118,N_1929);
nand U2503 (N_2503,N_1528,N_1413);
nand U2504 (N_2504,N_1614,N_1136);
nand U2505 (N_2505,N_1796,N_1289);
nor U2506 (N_2506,N_1040,N_1670);
or U2507 (N_2507,N_1413,N_1238);
nor U2508 (N_2508,N_1582,N_1093);
nor U2509 (N_2509,N_1797,N_1199);
nor U2510 (N_2510,N_1179,N_1257);
or U2511 (N_2511,N_1179,N_1850);
nor U2512 (N_2512,N_1017,N_1452);
nor U2513 (N_2513,N_1759,N_1599);
or U2514 (N_2514,N_1250,N_1429);
nor U2515 (N_2515,N_1282,N_1345);
nor U2516 (N_2516,N_1001,N_1293);
and U2517 (N_2517,N_1343,N_1362);
or U2518 (N_2518,N_1660,N_1840);
and U2519 (N_2519,N_1701,N_1584);
or U2520 (N_2520,N_1453,N_1520);
or U2521 (N_2521,N_1855,N_1719);
xnor U2522 (N_2522,N_1561,N_1137);
nand U2523 (N_2523,N_1717,N_1982);
nand U2524 (N_2524,N_1783,N_1421);
and U2525 (N_2525,N_1661,N_1334);
nand U2526 (N_2526,N_1880,N_1665);
nor U2527 (N_2527,N_1181,N_1426);
nor U2528 (N_2528,N_1668,N_1400);
nand U2529 (N_2529,N_1698,N_1057);
nor U2530 (N_2530,N_1169,N_1286);
and U2531 (N_2531,N_1664,N_1019);
nor U2532 (N_2532,N_1355,N_1944);
or U2533 (N_2533,N_1769,N_1500);
nand U2534 (N_2534,N_1715,N_1437);
nor U2535 (N_2535,N_1176,N_1595);
nand U2536 (N_2536,N_1027,N_1443);
nor U2537 (N_2537,N_1144,N_1362);
nand U2538 (N_2538,N_1126,N_1040);
or U2539 (N_2539,N_1492,N_1655);
or U2540 (N_2540,N_1080,N_1122);
nor U2541 (N_2541,N_1300,N_1427);
or U2542 (N_2542,N_1135,N_1539);
and U2543 (N_2543,N_1677,N_1716);
and U2544 (N_2544,N_1448,N_1911);
nor U2545 (N_2545,N_1882,N_1350);
nand U2546 (N_2546,N_1147,N_1342);
and U2547 (N_2547,N_1166,N_1091);
nor U2548 (N_2548,N_1289,N_1866);
nand U2549 (N_2549,N_1821,N_1207);
nor U2550 (N_2550,N_1373,N_1007);
nand U2551 (N_2551,N_1611,N_1999);
and U2552 (N_2552,N_1795,N_1586);
and U2553 (N_2553,N_1873,N_1754);
and U2554 (N_2554,N_1794,N_1087);
nand U2555 (N_2555,N_1657,N_1991);
or U2556 (N_2556,N_1902,N_1200);
or U2557 (N_2557,N_1649,N_1021);
or U2558 (N_2558,N_1417,N_1258);
and U2559 (N_2559,N_1399,N_1421);
and U2560 (N_2560,N_1106,N_1663);
nor U2561 (N_2561,N_1803,N_1141);
nor U2562 (N_2562,N_1896,N_1056);
or U2563 (N_2563,N_1430,N_1641);
nand U2564 (N_2564,N_1471,N_1947);
and U2565 (N_2565,N_1020,N_1814);
or U2566 (N_2566,N_1663,N_1041);
or U2567 (N_2567,N_1241,N_1755);
and U2568 (N_2568,N_1488,N_1870);
nand U2569 (N_2569,N_1396,N_1281);
nor U2570 (N_2570,N_1637,N_1214);
or U2571 (N_2571,N_1312,N_1290);
and U2572 (N_2572,N_1386,N_1393);
nand U2573 (N_2573,N_1502,N_1606);
nand U2574 (N_2574,N_1239,N_1160);
nor U2575 (N_2575,N_1093,N_1367);
or U2576 (N_2576,N_1333,N_1525);
and U2577 (N_2577,N_1442,N_1785);
or U2578 (N_2578,N_1509,N_1666);
and U2579 (N_2579,N_1757,N_1001);
nor U2580 (N_2580,N_1862,N_1675);
nand U2581 (N_2581,N_1632,N_1926);
nor U2582 (N_2582,N_1829,N_1642);
and U2583 (N_2583,N_1387,N_1737);
nor U2584 (N_2584,N_1063,N_1466);
nor U2585 (N_2585,N_1494,N_1964);
or U2586 (N_2586,N_1032,N_1432);
nand U2587 (N_2587,N_1028,N_1976);
nor U2588 (N_2588,N_1544,N_1200);
and U2589 (N_2589,N_1244,N_1718);
nand U2590 (N_2590,N_1496,N_1850);
or U2591 (N_2591,N_1692,N_1684);
nand U2592 (N_2592,N_1705,N_1397);
and U2593 (N_2593,N_1032,N_1813);
nor U2594 (N_2594,N_1853,N_1309);
nor U2595 (N_2595,N_1111,N_1073);
nor U2596 (N_2596,N_1686,N_1594);
or U2597 (N_2597,N_1312,N_1079);
nor U2598 (N_2598,N_1112,N_1095);
or U2599 (N_2599,N_1804,N_1845);
nor U2600 (N_2600,N_1789,N_1810);
nor U2601 (N_2601,N_1435,N_1887);
or U2602 (N_2602,N_1682,N_1530);
and U2603 (N_2603,N_1577,N_1120);
nor U2604 (N_2604,N_1769,N_1768);
nor U2605 (N_2605,N_1037,N_1474);
and U2606 (N_2606,N_1309,N_1570);
nand U2607 (N_2607,N_1666,N_1459);
or U2608 (N_2608,N_1484,N_1757);
nand U2609 (N_2609,N_1272,N_1894);
nor U2610 (N_2610,N_1335,N_1299);
or U2611 (N_2611,N_1892,N_1987);
or U2612 (N_2612,N_1323,N_1336);
nor U2613 (N_2613,N_1557,N_1892);
nand U2614 (N_2614,N_1145,N_1021);
nand U2615 (N_2615,N_1202,N_1016);
nand U2616 (N_2616,N_1671,N_1563);
or U2617 (N_2617,N_1737,N_1448);
and U2618 (N_2618,N_1787,N_1388);
nand U2619 (N_2619,N_1265,N_1094);
or U2620 (N_2620,N_1302,N_1983);
and U2621 (N_2621,N_1896,N_1988);
or U2622 (N_2622,N_1441,N_1657);
nor U2623 (N_2623,N_1022,N_1662);
or U2624 (N_2624,N_1230,N_1628);
nand U2625 (N_2625,N_1232,N_1403);
or U2626 (N_2626,N_1763,N_1493);
nand U2627 (N_2627,N_1090,N_1717);
nand U2628 (N_2628,N_1825,N_1999);
and U2629 (N_2629,N_1464,N_1375);
and U2630 (N_2630,N_1082,N_1102);
nor U2631 (N_2631,N_1100,N_1258);
and U2632 (N_2632,N_1337,N_1849);
or U2633 (N_2633,N_1890,N_1620);
nor U2634 (N_2634,N_1302,N_1104);
nand U2635 (N_2635,N_1351,N_1234);
or U2636 (N_2636,N_1399,N_1450);
nand U2637 (N_2637,N_1185,N_1875);
nand U2638 (N_2638,N_1326,N_1664);
and U2639 (N_2639,N_1625,N_1740);
or U2640 (N_2640,N_1814,N_1408);
nor U2641 (N_2641,N_1080,N_1752);
xnor U2642 (N_2642,N_1269,N_1838);
nor U2643 (N_2643,N_1159,N_1854);
nand U2644 (N_2644,N_1622,N_1899);
nand U2645 (N_2645,N_1811,N_1623);
or U2646 (N_2646,N_1804,N_1780);
nor U2647 (N_2647,N_1814,N_1003);
and U2648 (N_2648,N_1516,N_1823);
and U2649 (N_2649,N_1160,N_1191);
nand U2650 (N_2650,N_1027,N_1534);
nand U2651 (N_2651,N_1306,N_1018);
nand U2652 (N_2652,N_1515,N_1876);
and U2653 (N_2653,N_1840,N_1200);
xor U2654 (N_2654,N_1798,N_1352);
nand U2655 (N_2655,N_1589,N_1435);
nor U2656 (N_2656,N_1783,N_1077);
or U2657 (N_2657,N_1666,N_1684);
nand U2658 (N_2658,N_1977,N_1639);
nand U2659 (N_2659,N_1069,N_1044);
or U2660 (N_2660,N_1333,N_1813);
nor U2661 (N_2661,N_1434,N_1232);
or U2662 (N_2662,N_1982,N_1686);
and U2663 (N_2663,N_1349,N_1080);
nand U2664 (N_2664,N_1573,N_1636);
or U2665 (N_2665,N_1437,N_1289);
or U2666 (N_2666,N_1149,N_1357);
nor U2667 (N_2667,N_1940,N_1613);
nor U2668 (N_2668,N_1104,N_1927);
or U2669 (N_2669,N_1731,N_1764);
and U2670 (N_2670,N_1067,N_1061);
nand U2671 (N_2671,N_1572,N_1025);
nor U2672 (N_2672,N_1945,N_1923);
or U2673 (N_2673,N_1156,N_1449);
nand U2674 (N_2674,N_1165,N_1532);
nor U2675 (N_2675,N_1387,N_1099);
and U2676 (N_2676,N_1029,N_1226);
nor U2677 (N_2677,N_1681,N_1432);
nor U2678 (N_2678,N_1787,N_1118);
nand U2679 (N_2679,N_1675,N_1638);
nor U2680 (N_2680,N_1916,N_1966);
and U2681 (N_2681,N_1883,N_1192);
and U2682 (N_2682,N_1631,N_1902);
or U2683 (N_2683,N_1066,N_1948);
nor U2684 (N_2684,N_1839,N_1283);
nand U2685 (N_2685,N_1787,N_1823);
or U2686 (N_2686,N_1469,N_1029);
and U2687 (N_2687,N_1387,N_1070);
or U2688 (N_2688,N_1310,N_1144);
nand U2689 (N_2689,N_1248,N_1495);
or U2690 (N_2690,N_1067,N_1924);
nor U2691 (N_2691,N_1249,N_1797);
and U2692 (N_2692,N_1214,N_1170);
nand U2693 (N_2693,N_1694,N_1848);
or U2694 (N_2694,N_1995,N_1198);
and U2695 (N_2695,N_1478,N_1957);
and U2696 (N_2696,N_1743,N_1206);
nand U2697 (N_2697,N_1468,N_1195);
nand U2698 (N_2698,N_1451,N_1255);
or U2699 (N_2699,N_1323,N_1957);
and U2700 (N_2700,N_1497,N_1160);
nand U2701 (N_2701,N_1845,N_1512);
and U2702 (N_2702,N_1096,N_1329);
or U2703 (N_2703,N_1865,N_1592);
nand U2704 (N_2704,N_1334,N_1994);
or U2705 (N_2705,N_1003,N_1066);
or U2706 (N_2706,N_1788,N_1786);
and U2707 (N_2707,N_1208,N_1357);
and U2708 (N_2708,N_1395,N_1314);
and U2709 (N_2709,N_1191,N_1860);
and U2710 (N_2710,N_1615,N_1788);
or U2711 (N_2711,N_1414,N_1457);
or U2712 (N_2712,N_1874,N_1061);
xnor U2713 (N_2713,N_1616,N_1097);
nand U2714 (N_2714,N_1284,N_1559);
nor U2715 (N_2715,N_1530,N_1087);
or U2716 (N_2716,N_1335,N_1772);
or U2717 (N_2717,N_1895,N_1261);
nor U2718 (N_2718,N_1442,N_1010);
xor U2719 (N_2719,N_1577,N_1223);
nand U2720 (N_2720,N_1129,N_1209);
or U2721 (N_2721,N_1263,N_1549);
or U2722 (N_2722,N_1563,N_1050);
or U2723 (N_2723,N_1145,N_1047);
or U2724 (N_2724,N_1604,N_1682);
or U2725 (N_2725,N_1738,N_1162);
xnor U2726 (N_2726,N_1596,N_1429);
nand U2727 (N_2727,N_1539,N_1247);
or U2728 (N_2728,N_1789,N_1699);
nor U2729 (N_2729,N_1559,N_1293);
nand U2730 (N_2730,N_1351,N_1029);
nor U2731 (N_2731,N_1877,N_1503);
and U2732 (N_2732,N_1693,N_1581);
nor U2733 (N_2733,N_1493,N_1428);
nand U2734 (N_2734,N_1729,N_1506);
nand U2735 (N_2735,N_1251,N_1344);
nand U2736 (N_2736,N_1476,N_1469);
nor U2737 (N_2737,N_1373,N_1741);
nor U2738 (N_2738,N_1347,N_1264);
and U2739 (N_2739,N_1333,N_1048);
and U2740 (N_2740,N_1224,N_1262);
and U2741 (N_2741,N_1991,N_1520);
nor U2742 (N_2742,N_1017,N_1396);
or U2743 (N_2743,N_1894,N_1632);
nor U2744 (N_2744,N_1802,N_1856);
and U2745 (N_2745,N_1768,N_1551);
nand U2746 (N_2746,N_1846,N_1700);
or U2747 (N_2747,N_1962,N_1575);
nor U2748 (N_2748,N_1383,N_1441);
nand U2749 (N_2749,N_1293,N_1643);
and U2750 (N_2750,N_1198,N_1875);
or U2751 (N_2751,N_1841,N_1332);
xnor U2752 (N_2752,N_1494,N_1799);
nand U2753 (N_2753,N_1335,N_1814);
and U2754 (N_2754,N_1840,N_1400);
nand U2755 (N_2755,N_1616,N_1956);
xnor U2756 (N_2756,N_1024,N_1591);
nand U2757 (N_2757,N_1710,N_1867);
nand U2758 (N_2758,N_1408,N_1219);
and U2759 (N_2759,N_1662,N_1729);
nor U2760 (N_2760,N_1879,N_1909);
and U2761 (N_2761,N_1364,N_1978);
or U2762 (N_2762,N_1143,N_1168);
nand U2763 (N_2763,N_1163,N_1766);
or U2764 (N_2764,N_1725,N_1210);
nor U2765 (N_2765,N_1079,N_1538);
nand U2766 (N_2766,N_1846,N_1999);
nor U2767 (N_2767,N_1189,N_1127);
and U2768 (N_2768,N_1213,N_1804);
nand U2769 (N_2769,N_1500,N_1633);
nand U2770 (N_2770,N_1640,N_1042);
nand U2771 (N_2771,N_1353,N_1654);
nand U2772 (N_2772,N_1978,N_1104);
and U2773 (N_2773,N_1215,N_1684);
and U2774 (N_2774,N_1622,N_1962);
nor U2775 (N_2775,N_1948,N_1025);
and U2776 (N_2776,N_1396,N_1666);
nand U2777 (N_2777,N_1731,N_1484);
nand U2778 (N_2778,N_1150,N_1241);
nand U2779 (N_2779,N_1950,N_1413);
or U2780 (N_2780,N_1773,N_1568);
and U2781 (N_2781,N_1659,N_1619);
and U2782 (N_2782,N_1156,N_1428);
or U2783 (N_2783,N_1482,N_1019);
nand U2784 (N_2784,N_1365,N_1724);
and U2785 (N_2785,N_1120,N_1405);
nor U2786 (N_2786,N_1744,N_1789);
nand U2787 (N_2787,N_1459,N_1327);
and U2788 (N_2788,N_1069,N_1687);
or U2789 (N_2789,N_1461,N_1853);
nand U2790 (N_2790,N_1079,N_1760);
or U2791 (N_2791,N_1167,N_1182);
or U2792 (N_2792,N_1235,N_1028);
or U2793 (N_2793,N_1280,N_1920);
nand U2794 (N_2794,N_1910,N_1696);
nor U2795 (N_2795,N_1129,N_1292);
nand U2796 (N_2796,N_1659,N_1942);
or U2797 (N_2797,N_1190,N_1545);
and U2798 (N_2798,N_1432,N_1404);
nor U2799 (N_2799,N_1495,N_1615);
and U2800 (N_2800,N_1903,N_1081);
or U2801 (N_2801,N_1022,N_1166);
or U2802 (N_2802,N_1052,N_1808);
nor U2803 (N_2803,N_1146,N_1491);
nor U2804 (N_2804,N_1649,N_1480);
or U2805 (N_2805,N_1497,N_1855);
or U2806 (N_2806,N_1975,N_1219);
nand U2807 (N_2807,N_1990,N_1153);
nand U2808 (N_2808,N_1119,N_1256);
or U2809 (N_2809,N_1561,N_1993);
nor U2810 (N_2810,N_1834,N_1967);
or U2811 (N_2811,N_1796,N_1116);
and U2812 (N_2812,N_1417,N_1161);
nor U2813 (N_2813,N_1168,N_1137);
nor U2814 (N_2814,N_1669,N_1061);
xor U2815 (N_2815,N_1203,N_1015);
or U2816 (N_2816,N_1752,N_1575);
nor U2817 (N_2817,N_1968,N_1228);
and U2818 (N_2818,N_1695,N_1911);
or U2819 (N_2819,N_1275,N_1576);
nand U2820 (N_2820,N_1193,N_1580);
nor U2821 (N_2821,N_1741,N_1788);
and U2822 (N_2822,N_1842,N_1262);
and U2823 (N_2823,N_1074,N_1312);
or U2824 (N_2824,N_1465,N_1988);
nand U2825 (N_2825,N_1280,N_1179);
nor U2826 (N_2826,N_1412,N_1942);
or U2827 (N_2827,N_1098,N_1794);
or U2828 (N_2828,N_1147,N_1569);
or U2829 (N_2829,N_1599,N_1501);
and U2830 (N_2830,N_1618,N_1404);
nor U2831 (N_2831,N_1600,N_1419);
or U2832 (N_2832,N_1381,N_1438);
nand U2833 (N_2833,N_1250,N_1910);
and U2834 (N_2834,N_1619,N_1547);
nor U2835 (N_2835,N_1814,N_1758);
or U2836 (N_2836,N_1753,N_1284);
nand U2837 (N_2837,N_1888,N_1060);
and U2838 (N_2838,N_1183,N_1431);
and U2839 (N_2839,N_1048,N_1794);
nor U2840 (N_2840,N_1514,N_1794);
or U2841 (N_2841,N_1480,N_1021);
nor U2842 (N_2842,N_1071,N_1664);
nand U2843 (N_2843,N_1467,N_1609);
nand U2844 (N_2844,N_1371,N_1332);
nor U2845 (N_2845,N_1579,N_1722);
and U2846 (N_2846,N_1604,N_1383);
nand U2847 (N_2847,N_1993,N_1991);
nor U2848 (N_2848,N_1768,N_1270);
and U2849 (N_2849,N_1385,N_1532);
nand U2850 (N_2850,N_1712,N_1061);
nor U2851 (N_2851,N_1979,N_1396);
and U2852 (N_2852,N_1553,N_1636);
nor U2853 (N_2853,N_1582,N_1238);
and U2854 (N_2854,N_1236,N_1121);
and U2855 (N_2855,N_1409,N_1893);
nor U2856 (N_2856,N_1891,N_1178);
nand U2857 (N_2857,N_1230,N_1972);
and U2858 (N_2858,N_1131,N_1010);
and U2859 (N_2859,N_1279,N_1190);
and U2860 (N_2860,N_1107,N_1963);
or U2861 (N_2861,N_1429,N_1821);
and U2862 (N_2862,N_1039,N_1234);
and U2863 (N_2863,N_1605,N_1617);
nor U2864 (N_2864,N_1703,N_1969);
or U2865 (N_2865,N_1821,N_1707);
nand U2866 (N_2866,N_1136,N_1399);
nor U2867 (N_2867,N_1190,N_1707);
nand U2868 (N_2868,N_1936,N_1266);
and U2869 (N_2869,N_1076,N_1424);
nor U2870 (N_2870,N_1488,N_1863);
nor U2871 (N_2871,N_1463,N_1414);
nand U2872 (N_2872,N_1024,N_1658);
or U2873 (N_2873,N_1114,N_1142);
nor U2874 (N_2874,N_1963,N_1561);
nand U2875 (N_2875,N_1131,N_1841);
and U2876 (N_2876,N_1364,N_1936);
or U2877 (N_2877,N_1514,N_1641);
and U2878 (N_2878,N_1880,N_1653);
and U2879 (N_2879,N_1755,N_1378);
nor U2880 (N_2880,N_1296,N_1517);
and U2881 (N_2881,N_1002,N_1257);
nand U2882 (N_2882,N_1855,N_1100);
nand U2883 (N_2883,N_1569,N_1205);
and U2884 (N_2884,N_1036,N_1810);
and U2885 (N_2885,N_1037,N_1957);
or U2886 (N_2886,N_1413,N_1615);
and U2887 (N_2887,N_1794,N_1268);
or U2888 (N_2888,N_1001,N_1194);
and U2889 (N_2889,N_1195,N_1795);
nand U2890 (N_2890,N_1230,N_1404);
and U2891 (N_2891,N_1616,N_1126);
nor U2892 (N_2892,N_1594,N_1803);
nand U2893 (N_2893,N_1848,N_1720);
and U2894 (N_2894,N_1597,N_1963);
nand U2895 (N_2895,N_1537,N_1815);
and U2896 (N_2896,N_1579,N_1732);
nor U2897 (N_2897,N_1595,N_1994);
and U2898 (N_2898,N_1156,N_1990);
and U2899 (N_2899,N_1111,N_1383);
nand U2900 (N_2900,N_1506,N_1612);
or U2901 (N_2901,N_1022,N_1497);
nand U2902 (N_2902,N_1982,N_1654);
nand U2903 (N_2903,N_1211,N_1993);
or U2904 (N_2904,N_1969,N_1256);
nor U2905 (N_2905,N_1700,N_1674);
and U2906 (N_2906,N_1174,N_1817);
or U2907 (N_2907,N_1534,N_1111);
or U2908 (N_2908,N_1142,N_1297);
nor U2909 (N_2909,N_1876,N_1400);
nor U2910 (N_2910,N_1567,N_1484);
or U2911 (N_2911,N_1320,N_1253);
or U2912 (N_2912,N_1196,N_1251);
or U2913 (N_2913,N_1630,N_1590);
nor U2914 (N_2914,N_1003,N_1812);
and U2915 (N_2915,N_1088,N_1102);
nand U2916 (N_2916,N_1644,N_1887);
or U2917 (N_2917,N_1400,N_1398);
or U2918 (N_2918,N_1452,N_1287);
and U2919 (N_2919,N_1517,N_1254);
nor U2920 (N_2920,N_1402,N_1337);
or U2921 (N_2921,N_1191,N_1641);
and U2922 (N_2922,N_1494,N_1974);
and U2923 (N_2923,N_1078,N_1028);
or U2924 (N_2924,N_1129,N_1778);
or U2925 (N_2925,N_1850,N_1084);
or U2926 (N_2926,N_1576,N_1931);
and U2927 (N_2927,N_1984,N_1478);
nand U2928 (N_2928,N_1428,N_1877);
or U2929 (N_2929,N_1556,N_1479);
and U2930 (N_2930,N_1672,N_1733);
or U2931 (N_2931,N_1796,N_1495);
and U2932 (N_2932,N_1598,N_1223);
and U2933 (N_2933,N_1605,N_1578);
nor U2934 (N_2934,N_1055,N_1139);
nand U2935 (N_2935,N_1503,N_1051);
nand U2936 (N_2936,N_1684,N_1397);
nor U2937 (N_2937,N_1243,N_1730);
and U2938 (N_2938,N_1209,N_1170);
nor U2939 (N_2939,N_1355,N_1826);
or U2940 (N_2940,N_1696,N_1150);
and U2941 (N_2941,N_1369,N_1629);
nand U2942 (N_2942,N_1083,N_1563);
nand U2943 (N_2943,N_1571,N_1050);
nor U2944 (N_2944,N_1906,N_1180);
and U2945 (N_2945,N_1181,N_1711);
nor U2946 (N_2946,N_1731,N_1587);
and U2947 (N_2947,N_1290,N_1594);
and U2948 (N_2948,N_1292,N_1483);
and U2949 (N_2949,N_1952,N_1402);
nand U2950 (N_2950,N_1134,N_1907);
nand U2951 (N_2951,N_1906,N_1372);
nor U2952 (N_2952,N_1009,N_1048);
and U2953 (N_2953,N_1591,N_1968);
nor U2954 (N_2954,N_1662,N_1092);
nand U2955 (N_2955,N_1802,N_1118);
nand U2956 (N_2956,N_1804,N_1706);
or U2957 (N_2957,N_1196,N_1619);
or U2958 (N_2958,N_1974,N_1342);
nand U2959 (N_2959,N_1744,N_1855);
and U2960 (N_2960,N_1320,N_1514);
or U2961 (N_2961,N_1521,N_1310);
or U2962 (N_2962,N_1925,N_1752);
nor U2963 (N_2963,N_1209,N_1441);
nand U2964 (N_2964,N_1333,N_1202);
nor U2965 (N_2965,N_1182,N_1975);
or U2966 (N_2966,N_1265,N_1076);
nand U2967 (N_2967,N_1093,N_1995);
nor U2968 (N_2968,N_1124,N_1294);
or U2969 (N_2969,N_1052,N_1352);
and U2970 (N_2970,N_1649,N_1550);
nand U2971 (N_2971,N_1311,N_1362);
or U2972 (N_2972,N_1481,N_1114);
nand U2973 (N_2973,N_1106,N_1039);
nand U2974 (N_2974,N_1494,N_1441);
nand U2975 (N_2975,N_1130,N_1658);
or U2976 (N_2976,N_1195,N_1260);
nand U2977 (N_2977,N_1180,N_1101);
nand U2978 (N_2978,N_1098,N_1644);
and U2979 (N_2979,N_1691,N_1204);
nand U2980 (N_2980,N_1152,N_1338);
nand U2981 (N_2981,N_1172,N_1054);
or U2982 (N_2982,N_1499,N_1158);
or U2983 (N_2983,N_1736,N_1979);
or U2984 (N_2984,N_1945,N_1453);
or U2985 (N_2985,N_1073,N_1953);
nand U2986 (N_2986,N_1068,N_1769);
nor U2987 (N_2987,N_1409,N_1730);
or U2988 (N_2988,N_1048,N_1375);
or U2989 (N_2989,N_1647,N_1277);
and U2990 (N_2990,N_1576,N_1668);
and U2991 (N_2991,N_1654,N_1404);
and U2992 (N_2992,N_1960,N_1409);
nand U2993 (N_2993,N_1679,N_1953);
and U2994 (N_2994,N_1850,N_1718);
or U2995 (N_2995,N_1366,N_1283);
nand U2996 (N_2996,N_1284,N_1720);
nor U2997 (N_2997,N_1823,N_1301);
nor U2998 (N_2998,N_1072,N_1686);
or U2999 (N_2999,N_1333,N_1475);
and UO_0 (O_0,N_2475,N_2987);
nand UO_1 (O_1,N_2691,N_2986);
nor UO_2 (O_2,N_2410,N_2737);
nor UO_3 (O_3,N_2403,N_2396);
and UO_4 (O_4,N_2721,N_2659);
nand UO_5 (O_5,N_2941,N_2505);
and UO_6 (O_6,N_2338,N_2142);
and UO_7 (O_7,N_2347,N_2872);
nand UO_8 (O_8,N_2368,N_2062);
or UO_9 (O_9,N_2975,N_2816);
and UO_10 (O_10,N_2759,N_2565);
or UO_11 (O_11,N_2594,N_2307);
or UO_12 (O_12,N_2133,N_2749);
nor UO_13 (O_13,N_2481,N_2956);
and UO_14 (O_14,N_2595,N_2453);
nand UO_15 (O_15,N_2220,N_2025);
and UO_16 (O_16,N_2778,N_2241);
nor UO_17 (O_17,N_2576,N_2797);
nor UO_18 (O_18,N_2512,N_2988);
nor UO_19 (O_19,N_2443,N_2240);
or UO_20 (O_20,N_2803,N_2262);
or UO_21 (O_21,N_2924,N_2501);
or UO_22 (O_22,N_2442,N_2112);
and UO_23 (O_23,N_2199,N_2952);
or UO_24 (O_24,N_2040,N_2104);
nor UO_25 (O_25,N_2331,N_2369);
and UO_26 (O_26,N_2490,N_2680);
or UO_27 (O_27,N_2276,N_2179);
nor UO_28 (O_28,N_2796,N_2111);
or UO_29 (O_29,N_2608,N_2309);
and UO_30 (O_30,N_2878,N_2838);
and UO_31 (O_31,N_2468,N_2929);
and UO_32 (O_32,N_2406,N_2108);
nor UO_33 (O_33,N_2429,N_2556);
and UO_34 (O_34,N_2761,N_2200);
nand UO_35 (O_35,N_2944,N_2847);
or UO_36 (O_36,N_2817,N_2123);
or UO_37 (O_37,N_2160,N_2055);
or UO_38 (O_38,N_2416,N_2516);
and UO_39 (O_39,N_2744,N_2425);
and UO_40 (O_40,N_2640,N_2903);
nand UO_41 (O_41,N_2122,N_2943);
and UO_42 (O_42,N_2794,N_2017);
or UO_43 (O_43,N_2626,N_2320);
nand UO_44 (O_44,N_2867,N_2694);
and UO_45 (O_45,N_2426,N_2610);
nand UO_46 (O_46,N_2682,N_2086);
nor UO_47 (O_47,N_2243,N_2820);
nor UO_48 (O_48,N_2402,N_2921);
nor UO_49 (O_49,N_2272,N_2973);
xor UO_50 (O_50,N_2035,N_2885);
and UO_51 (O_51,N_2394,N_2689);
nor UO_52 (O_52,N_2837,N_2587);
nand UO_53 (O_53,N_2831,N_2101);
nor UO_54 (O_54,N_2934,N_2568);
and UO_55 (O_55,N_2553,N_2033);
nand UO_56 (O_56,N_2018,N_2213);
and UO_57 (O_57,N_2738,N_2939);
nand UO_58 (O_58,N_2823,N_2539);
or UO_59 (O_59,N_2182,N_2912);
nand UO_60 (O_60,N_2683,N_2642);
nand UO_61 (O_61,N_2011,N_2418);
nand UO_62 (O_62,N_2190,N_2487);
nor UO_63 (O_63,N_2357,N_2137);
and UO_64 (O_64,N_2319,N_2084);
nor UO_65 (O_65,N_2494,N_2644);
and UO_66 (O_66,N_2703,N_2981);
nor UO_67 (O_67,N_2162,N_2128);
nand UO_68 (O_68,N_2381,N_2269);
or UO_69 (O_69,N_2109,N_2541);
nand UO_70 (O_70,N_2016,N_2284);
nor UO_71 (O_71,N_2664,N_2253);
and UO_72 (O_72,N_2238,N_2379);
and UO_73 (O_73,N_2853,N_2917);
and UO_74 (O_74,N_2449,N_2730);
and UO_75 (O_75,N_2012,N_2953);
nand UO_76 (O_76,N_2722,N_2521);
and UO_77 (O_77,N_2047,N_2962);
or UO_78 (O_78,N_2914,N_2554);
and UO_79 (O_79,N_2584,N_2651);
and UO_80 (O_80,N_2242,N_2827);
nor UO_81 (O_81,N_2996,N_2804);
and UO_82 (O_82,N_2311,N_2138);
nand UO_83 (O_83,N_2513,N_2520);
and UO_84 (O_84,N_2997,N_2968);
nor UO_85 (O_85,N_2909,N_2447);
nor UO_86 (O_86,N_2881,N_2714);
nand UO_87 (O_87,N_2883,N_2264);
and UO_88 (O_88,N_2724,N_2150);
nor UO_89 (O_89,N_2788,N_2223);
or UO_90 (O_90,N_2469,N_2672);
nor UO_91 (O_91,N_2898,N_2419);
or UO_92 (O_92,N_2464,N_2155);
nand UO_93 (O_93,N_2908,N_2544);
xnor UO_94 (O_94,N_2135,N_2792);
or UO_95 (O_95,N_2052,N_2774);
nand UO_96 (O_96,N_2857,N_2600);
or UO_97 (O_97,N_2573,N_2446);
nor UO_98 (O_98,N_2221,N_2994);
nor UO_99 (O_99,N_2334,N_2198);
nor UO_100 (O_100,N_2583,N_2391);
and UO_101 (O_101,N_2614,N_2329);
and UO_102 (O_102,N_2219,N_2550);
nand UO_103 (O_103,N_2799,N_2725);
nor UO_104 (O_104,N_2913,N_2234);
nand UO_105 (O_105,N_2631,N_2578);
or UO_106 (O_106,N_2060,N_2299);
nand UO_107 (O_107,N_2189,N_2826);
or UO_108 (O_108,N_2059,N_2606);
nand UO_109 (O_109,N_2280,N_2237);
and UO_110 (O_110,N_2212,N_2326);
or UO_111 (O_111,N_2066,N_2302);
nand UO_112 (O_112,N_2582,N_2581);
nand UO_113 (O_113,N_2008,N_2648);
and UO_114 (O_114,N_2586,N_2151);
or UO_115 (O_115,N_2099,N_2641);
and UO_116 (O_116,N_2423,N_2174);
or UO_117 (O_117,N_2531,N_2841);
and UO_118 (O_118,N_2897,N_2688);
nand UO_119 (O_119,N_2285,N_2766);
nor UO_120 (O_120,N_2843,N_2315);
xor UO_121 (O_121,N_2668,N_2627);
and UO_122 (O_122,N_2291,N_2471);
nand UO_123 (O_123,N_2348,N_2764);
or UO_124 (O_124,N_2455,N_2239);
and UO_125 (O_125,N_2144,N_2933);
or UO_126 (O_126,N_2364,N_2875);
and UO_127 (O_127,N_2547,N_2965);
nand UO_128 (O_128,N_2014,N_2925);
nand UO_129 (O_129,N_2617,N_2798);
nand UO_130 (O_130,N_2963,N_2545);
nand UO_131 (O_131,N_2624,N_2720);
and UO_132 (O_132,N_2166,N_2528);
or UO_133 (O_133,N_2218,N_2769);
nor UO_134 (O_134,N_2157,N_2283);
nand UO_135 (O_135,N_2785,N_2222);
nand UO_136 (O_136,N_2492,N_2932);
or UO_137 (O_137,N_2655,N_2890);
or UO_138 (O_138,N_2902,N_2639);
or UO_139 (O_139,N_2267,N_2716);
or UO_140 (O_140,N_2718,N_2032);
nand UO_141 (O_141,N_2662,N_2966);
or UO_142 (O_142,N_2409,N_2509);
or UO_143 (O_143,N_2957,N_2844);
nand UO_144 (O_144,N_2984,N_2169);
or UO_145 (O_145,N_2630,N_2927);
and UO_146 (O_146,N_2660,N_2700);
and UO_147 (O_147,N_2643,N_2559);
nor UO_148 (O_148,N_2846,N_2667);
and UO_149 (O_149,N_2736,N_2652);
and UO_150 (O_150,N_2090,N_2072);
or UO_151 (O_151,N_2413,N_2039);
nor UO_152 (O_152,N_2435,N_2275);
nor UO_153 (O_153,N_2712,N_2762);
nand UO_154 (O_154,N_2760,N_2673);
nor UO_155 (O_155,N_2589,N_2611);
nor UO_156 (O_156,N_2258,N_2585);
nand UO_157 (O_157,N_2830,N_2260);
or UO_158 (O_158,N_2923,N_2955);
nand UO_159 (O_159,N_2729,N_2503);
nand UO_160 (O_160,N_2197,N_2196);
nor UO_161 (O_161,N_2607,N_2980);
nor UO_162 (O_162,N_2085,N_2812);
and UO_163 (O_163,N_2244,N_2916);
and UO_164 (O_164,N_2438,N_2650);
nor UO_165 (O_165,N_2753,N_2656);
and UO_166 (O_166,N_2739,N_2633);
nor UO_167 (O_167,N_2010,N_2612);
and UO_168 (O_168,N_2873,N_2282);
nand UO_169 (O_169,N_2960,N_2312);
nand UO_170 (O_170,N_2510,N_2719);
nor UO_171 (O_171,N_2967,N_2888);
and UO_172 (O_172,N_2236,N_2819);
or UO_173 (O_173,N_2593,N_2972);
nand UO_174 (O_174,N_2715,N_2995);
nand UO_175 (O_175,N_2246,N_2519);
and UO_176 (O_176,N_2003,N_2482);
or UO_177 (O_177,N_2188,N_2681);
nor UO_178 (O_178,N_2530,N_2910);
nor UO_179 (O_179,N_2874,N_2733);
nor UO_180 (O_180,N_2027,N_2065);
nor UO_181 (O_181,N_2982,N_2839);
xor UO_182 (O_182,N_2470,N_2036);
nand UO_183 (O_183,N_2942,N_2177);
or UO_184 (O_184,N_2918,N_2105);
or UO_185 (O_185,N_2328,N_2495);
nor UO_186 (O_186,N_2524,N_2444);
and UO_187 (O_187,N_2178,N_2723);
nand UO_188 (O_188,N_2063,N_2193);
nand UO_189 (O_189,N_2287,N_2459);
or UO_190 (O_190,N_2095,N_2231);
nand UO_191 (O_191,N_2552,N_2863);
nor UO_192 (O_192,N_2344,N_2833);
nor UO_193 (O_193,N_2677,N_2743);
and UO_194 (O_194,N_2534,N_2895);
and UO_195 (O_195,N_2834,N_2889);
and UO_196 (O_196,N_2810,N_2332);
or UO_197 (O_197,N_2336,N_2690);
nand UO_198 (O_198,N_2054,N_2658);
nand UO_199 (O_199,N_2367,N_2207);
and UO_200 (O_200,N_2590,N_2570);
nand UO_201 (O_201,N_2339,N_2560);
nand UO_202 (O_202,N_2731,N_2257);
nor UO_203 (O_203,N_2814,N_2388);
nor UO_204 (O_204,N_2674,N_2372);
or UO_205 (O_205,N_2615,N_2015);
or UO_206 (O_206,N_2949,N_2161);
nand UO_207 (O_207,N_2907,N_2609);
nand UO_208 (O_208,N_2170,N_2389);
nor UO_209 (O_209,N_2599,N_2130);
nor UO_210 (O_210,N_2784,N_2051);
nor UO_211 (O_211,N_2536,N_2928);
and UO_212 (O_212,N_2143,N_2758);
and UO_213 (O_213,N_2954,N_2415);
nor UO_214 (O_214,N_2024,N_2210);
and UO_215 (O_215,N_2430,N_2303);
or UO_216 (O_216,N_2686,N_2555);
nand UO_217 (O_217,N_2567,N_2097);
or UO_218 (O_218,N_2373,N_2868);
and UO_219 (O_219,N_2383,N_2786);
and UO_220 (O_220,N_2164,N_2399);
or UO_221 (O_221,N_2670,N_2374);
xor UO_222 (O_222,N_2249,N_2103);
and UO_223 (O_223,N_2575,N_2605);
nor UO_224 (O_224,N_2647,N_2855);
or UO_225 (O_225,N_2261,N_2476);
nand UO_226 (O_226,N_2361,N_2864);
nand UO_227 (O_227,N_2851,N_2542);
and UO_228 (O_228,N_2489,N_2022);
or UO_229 (O_229,N_2124,N_2358);
and UO_230 (O_230,N_2472,N_2202);
nand UO_231 (O_231,N_2629,N_2692);
and UO_232 (O_232,N_2397,N_2288);
nor UO_233 (O_233,N_2323,N_2789);
nand UO_234 (O_234,N_2896,N_2945);
nand UO_235 (O_235,N_2300,N_2549);
and UO_236 (O_236,N_2071,N_2286);
and UO_237 (O_237,N_2499,N_2382);
nor UO_238 (O_238,N_2380,N_2049);
nor UO_239 (O_239,N_2698,N_2079);
and UO_240 (O_240,N_2488,N_2508);
nor UO_241 (O_241,N_2707,N_2871);
and UO_242 (O_242,N_2622,N_2526);
or UO_243 (O_243,N_2001,N_2392);
nand UO_244 (O_244,N_2543,N_2989);
and UO_245 (O_245,N_2330,N_2214);
or UO_246 (O_246,N_2901,N_2821);
nor UO_247 (O_247,N_2306,N_2290);
nand UO_248 (O_248,N_2384,N_2046);
nand UO_249 (O_249,N_2842,N_2529);
nand UO_250 (O_250,N_2407,N_2776);
nand UO_251 (O_251,N_2119,N_2882);
and UO_252 (O_252,N_2637,N_2517);
nor UO_253 (O_253,N_2461,N_2129);
and UO_254 (O_254,N_2087,N_2825);
nor UO_255 (O_255,N_2279,N_2006);
nand UO_256 (O_256,N_2704,N_2400);
nor UO_257 (O_257,N_2616,N_2184);
nand UO_258 (O_258,N_2665,N_2195);
nand UO_259 (O_259,N_2106,N_2362);
nand UO_260 (O_260,N_2533,N_2645);
nand UO_261 (O_261,N_2993,N_2678);
nand UO_262 (O_262,N_2978,N_2057);
xor UO_263 (O_263,N_2206,N_2225);
and UO_264 (O_264,N_2779,N_2434);
nor UO_265 (O_265,N_2327,N_2000);
nand UO_266 (O_266,N_2661,N_2301);
nand UO_267 (O_267,N_2156,N_2603);
or UO_268 (O_268,N_2412,N_2795);
or UO_269 (O_269,N_2800,N_2205);
nor UO_270 (O_270,N_2822,N_2037);
nand UO_271 (O_271,N_2706,N_2393);
or UO_272 (O_272,N_2848,N_2741);
nor UO_273 (O_273,N_2181,N_2551);
nand UO_274 (O_274,N_2859,N_2904);
nor UO_275 (O_275,N_2346,N_2209);
nand UO_276 (O_276,N_2964,N_2163);
nor UO_277 (O_277,N_2751,N_2992);
nand UO_278 (O_278,N_2740,N_2755);
nor UO_279 (O_279,N_2783,N_2961);
nor UO_280 (O_280,N_2563,N_2313);
and UO_281 (O_281,N_2906,N_2805);
and UO_282 (O_282,N_2491,N_2201);
nor UO_283 (O_283,N_2118,N_2548);
nor UO_284 (O_284,N_2891,N_2705);
or UO_285 (O_285,N_2745,N_2951);
or UO_286 (O_286,N_2292,N_2748);
or UO_287 (O_287,N_2793,N_2376);
nand UO_288 (O_288,N_2165,N_2638);
or UO_289 (O_289,N_2815,N_2935);
or UO_290 (O_290,N_2363,N_2452);
and UO_291 (O_291,N_2773,N_2696);
nor UO_292 (O_292,N_2370,N_2985);
nand UO_293 (O_293,N_2849,N_2592);
nor UO_294 (O_294,N_2147,N_2088);
or UO_295 (O_295,N_2734,N_2070);
nand UO_296 (O_296,N_2131,N_2480);
nor UO_297 (O_297,N_2116,N_2096);
nand UO_298 (O_298,N_2132,N_2056);
nor UO_299 (O_299,N_2171,N_2628);
nor UO_300 (O_300,N_2440,N_2148);
or UO_301 (O_301,N_2938,N_2417);
and UO_302 (O_302,N_2523,N_2601);
and UO_303 (O_303,N_2149,N_2958);
nand UO_304 (O_304,N_2337,N_2224);
and UO_305 (O_305,N_2437,N_2884);
and UO_306 (O_306,N_2034,N_2504);
nand UO_307 (O_307,N_2002,N_2294);
or UO_308 (O_308,N_2588,N_2619);
nor UO_309 (O_309,N_2304,N_2340);
and UO_310 (O_310,N_2771,N_2031);
and UO_311 (O_311,N_2298,N_2044);
nand UO_312 (O_312,N_2634,N_2742);
or UO_313 (O_313,N_2126,N_2893);
and UO_314 (O_314,N_2950,N_2140);
nand UO_315 (O_315,N_2041,N_2926);
and UO_316 (O_316,N_2089,N_2646);
or UO_317 (O_317,N_2345,N_2693);
nor UO_318 (O_318,N_2676,N_2977);
and UO_319 (O_319,N_2602,N_2421);
nand UO_320 (O_320,N_2094,N_2146);
or UO_321 (O_321,N_2876,N_2377);
and UO_322 (O_322,N_2445,N_2232);
and UO_323 (O_323,N_2450,N_2710);
nand UO_324 (O_324,N_2020,N_2562);
or UO_325 (O_325,N_2657,N_2728);
or UO_326 (O_326,N_2082,N_2102);
nand UO_327 (O_327,N_2990,N_2502);
nand UO_328 (O_328,N_2577,N_2801);
nor UO_329 (O_329,N_2463,N_2525);
or UO_330 (O_330,N_2900,N_2078);
and UO_331 (O_331,N_2411,N_2152);
nand UO_332 (O_332,N_2937,N_2620);
and UO_333 (O_333,N_2043,N_2974);
nand UO_334 (O_334,N_2333,N_2217);
and UO_335 (O_335,N_2053,N_2321);
nor UO_336 (O_336,N_2979,N_2457);
nor UO_337 (O_337,N_2699,N_2113);
or UO_338 (O_338,N_2271,N_2216);
nand UO_339 (O_339,N_2750,N_2009);
and UO_340 (O_340,N_2959,N_2813);
nor UO_341 (O_341,N_2424,N_2013);
nand UO_342 (O_342,N_2856,N_2064);
nor UO_343 (O_343,N_2832,N_2768);
nor UO_344 (O_344,N_2727,N_2076);
or UO_345 (O_345,N_2467,N_2654);
and UO_346 (O_346,N_2756,N_2192);
or UO_347 (O_347,N_2247,N_2100);
nand UO_348 (O_348,N_2946,N_2752);
nor UO_349 (O_349,N_2173,N_2564);
nor UO_350 (O_350,N_2121,N_2653);
or UO_351 (O_351,N_2506,N_2865);
and UO_352 (O_352,N_2887,N_2120);
nor UO_353 (O_353,N_2777,N_2763);
and UO_354 (O_354,N_2145,N_2404);
nor UO_355 (O_355,N_2360,N_2414);
nor UO_356 (O_356,N_2685,N_2840);
or UO_357 (O_357,N_2515,N_2806);
nand UO_358 (O_358,N_2366,N_2324);
nor UO_359 (O_359,N_2824,N_2277);
and UO_360 (O_360,N_2462,N_2527);
nand UO_361 (O_361,N_2432,N_2858);
nand UO_362 (O_362,N_2483,N_2073);
or UO_363 (O_363,N_2067,N_2852);
nor UO_364 (O_364,N_2540,N_2317);
and UO_365 (O_365,N_2458,N_2836);
nor UO_366 (O_366,N_2354,N_2021);
and UO_367 (O_367,N_2316,N_2068);
or UO_368 (O_368,N_2127,N_2879);
nor UO_369 (O_369,N_2473,N_2061);
or UO_370 (O_370,N_2649,N_2746);
nand UO_371 (O_371,N_2405,N_2375);
nor UO_372 (O_372,N_2711,N_2083);
and UO_373 (O_373,N_2183,N_2259);
or UO_374 (O_374,N_2613,N_2572);
or UO_375 (O_375,N_2598,N_2134);
nor UO_376 (O_376,N_2350,N_2931);
or UO_377 (O_377,N_2922,N_2862);
nor UO_378 (O_378,N_2256,N_2180);
nor UO_379 (O_379,N_2341,N_2532);
xor UO_380 (O_380,N_2511,N_2781);
nor UO_381 (O_381,N_2114,N_2349);
nand UO_382 (O_382,N_2477,N_2186);
or UO_383 (O_383,N_2514,N_2310);
and UO_384 (O_384,N_2308,N_2870);
and UO_385 (O_385,N_2451,N_2398);
nand UO_386 (O_386,N_2618,N_2747);
nand UO_387 (O_387,N_2666,N_2365);
nor UO_388 (O_388,N_2561,N_2093);
or UO_389 (O_389,N_2167,N_2669);
and UO_390 (O_390,N_2172,N_2296);
or UO_391 (O_391,N_2940,N_2695);
nand UO_392 (O_392,N_2325,N_2697);
and UO_393 (O_393,N_2970,N_2636);
and UO_394 (O_394,N_2030,N_2625);
nor UO_395 (O_395,N_2204,N_2175);
and UO_396 (O_396,N_2886,N_2081);
nand UO_397 (O_397,N_2765,N_2230);
and UO_398 (O_398,N_2050,N_2702);
nor UO_399 (O_399,N_2187,N_2281);
nand UO_400 (O_400,N_2305,N_2735);
or UO_401 (O_401,N_2537,N_2635);
nand UO_402 (O_402,N_2623,N_2775);
nand UO_403 (O_403,N_2770,N_2215);
nor UO_404 (O_404,N_2808,N_2936);
nand UO_405 (O_405,N_2250,N_2058);
nand UO_406 (O_406,N_2265,N_2486);
and UO_407 (O_407,N_2289,N_2454);
or UO_408 (O_408,N_2228,N_2971);
or UO_409 (O_409,N_2546,N_2969);
and UO_410 (O_410,N_2478,N_2091);
nor UO_411 (O_411,N_2322,N_2048);
nor UO_412 (O_412,N_2159,N_2535);
and UO_413 (O_413,N_2191,N_2948);
or UO_414 (O_414,N_2436,N_2107);
or UO_415 (O_415,N_2732,N_2019);
nor UO_416 (O_416,N_2754,N_2401);
or UO_417 (O_417,N_2386,N_2075);
or UO_418 (O_418,N_2597,N_2905);
or UO_419 (O_419,N_2790,N_2497);
nor UO_420 (O_420,N_2371,N_2098);
nor UO_421 (O_421,N_2782,N_2356);
nand UO_422 (O_422,N_2420,N_2915);
or UO_423 (O_423,N_2355,N_2663);
or UO_424 (O_424,N_2077,N_2117);
and UO_425 (O_425,N_2042,N_2894);
nand UO_426 (O_426,N_2484,N_2390);
nor UO_427 (O_427,N_2465,N_2251);
and UO_428 (O_428,N_2866,N_2791);
and UO_429 (O_429,N_2342,N_2235);
or UO_430 (O_430,N_2580,N_2999);
nor UO_431 (O_431,N_2828,N_2226);
or UO_432 (O_432,N_2558,N_2496);
or UO_433 (O_433,N_2168,N_2136);
nor UO_434 (O_434,N_2538,N_2139);
and UO_435 (O_435,N_2485,N_2991);
nand UO_436 (O_436,N_2899,N_2203);
nor UO_437 (O_437,N_2353,N_2185);
or UO_438 (O_438,N_2807,N_2930);
nand UO_439 (O_439,N_2154,N_2479);
or UO_440 (O_440,N_2211,N_2273);
and UO_441 (O_441,N_2684,N_2518);
or UO_442 (O_442,N_2522,N_2233);
nand UO_443 (O_443,N_2023,N_2274);
or UO_444 (O_444,N_2671,N_2767);
and UO_445 (O_445,N_2708,N_2818);
nor UO_446 (O_446,N_2566,N_2431);
and UO_447 (O_447,N_2701,N_2428);
nor UO_448 (O_448,N_2433,N_2352);
or UO_449 (O_449,N_2632,N_2408);
nor UO_450 (O_450,N_2141,N_2687);
nand UO_451 (O_451,N_2787,N_2026);
and UO_452 (O_452,N_2110,N_2498);
nand UO_453 (O_453,N_2208,N_2675);
nor UO_454 (O_454,N_2318,N_2474);
nand UO_455 (O_455,N_2176,N_2713);
and UO_456 (O_456,N_2293,N_2297);
and UO_457 (O_457,N_2571,N_2880);
or UO_458 (O_458,N_2252,N_2314);
or UO_459 (O_459,N_2877,N_2278);
nor UO_460 (O_460,N_2245,N_2074);
nor UO_461 (O_461,N_2829,N_2850);
nor UO_462 (O_462,N_2569,N_2709);
nor UO_463 (O_463,N_2579,N_2809);
xnor UO_464 (O_464,N_2359,N_2493);
nand UO_465 (O_465,N_2780,N_2835);
and UO_466 (O_466,N_2466,N_2069);
or UO_467 (O_467,N_2460,N_2947);
nor UO_468 (O_468,N_2621,N_2004);
nor UO_469 (O_469,N_2919,N_2757);
nor UO_470 (O_470,N_2385,N_2263);
nor UO_471 (O_471,N_2920,N_2255);
nor UO_472 (O_472,N_2295,N_2115);
nand UO_473 (O_473,N_2422,N_2854);
nand UO_474 (O_474,N_2227,N_2194);
nor UO_475 (O_475,N_2158,N_2845);
and UO_476 (O_476,N_2351,N_2507);
nor UO_477 (O_477,N_2726,N_2395);
and UO_478 (O_478,N_2229,N_2335);
nor UO_479 (O_479,N_2268,N_2911);
nand UO_480 (O_480,N_2456,N_2427);
or UO_481 (O_481,N_2596,N_2892);
nor UO_482 (O_482,N_2254,N_2387);
and UO_483 (O_483,N_2574,N_2441);
nand UO_484 (O_484,N_2270,N_2976);
nand UO_485 (O_485,N_2448,N_2679);
nor UO_486 (O_486,N_2591,N_2007);
nor UO_487 (O_487,N_2998,N_2869);
and UO_488 (O_488,N_2860,N_2811);
nor UO_489 (O_489,N_2802,N_2500);
nand UO_490 (O_490,N_2029,N_2028);
nor UO_491 (O_491,N_2861,N_2983);
or UO_492 (O_492,N_2378,N_2080);
xnor UO_493 (O_493,N_2772,N_2125);
and UO_494 (O_494,N_2439,N_2266);
or UO_495 (O_495,N_2005,N_2038);
nand UO_496 (O_496,N_2604,N_2343);
and UO_497 (O_497,N_2248,N_2045);
and UO_498 (O_498,N_2557,N_2717);
or UO_499 (O_499,N_2092,N_2153);
endmodule