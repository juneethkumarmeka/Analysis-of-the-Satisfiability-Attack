module basic_750_5000_1000_10_levels_1xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
or U0 (N_0,In_418,In_708);
and U1 (N_1,In_365,In_293);
and U2 (N_2,In_172,In_717);
nor U3 (N_3,In_521,In_308);
nor U4 (N_4,In_360,In_488);
or U5 (N_5,In_292,In_223);
or U6 (N_6,In_90,In_562);
nand U7 (N_7,In_167,In_355);
nor U8 (N_8,In_291,In_736);
nand U9 (N_9,In_24,In_102);
or U10 (N_10,In_120,In_249);
and U11 (N_11,In_195,In_647);
nor U12 (N_12,In_83,In_53);
nand U13 (N_13,In_105,In_613);
or U14 (N_14,In_454,In_440);
or U15 (N_15,In_396,In_162);
or U16 (N_16,In_523,In_146);
and U17 (N_17,In_629,In_70);
or U18 (N_18,In_47,In_101);
nor U19 (N_19,In_286,In_408);
and U20 (N_20,In_151,In_137);
nor U21 (N_21,In_208,In_669);
nand U22 (N_22,In_502,In_362);
nor U23 (N_23,In_742,In_489);
or U24 (N_24,In_327,In_287);
and U25 (N_25,In_199,In_226);
and U26 (N_26,In_580,In_182);
nand U27 (N_27,In_354,In_675);
and U28 (N_28,In_649,In_439);
nor U29 (N_29,In_343,In_247);
and U30 (N_30,In_155,In_159);
nor U31 (N_31,In_433,In_670);
and U32 (N_32,In_325,In_201);
or U33 (N_33,In_683,In_635);
and U34 (N_34,In_381,In_737);
nor U35 (N_35,In_676,In_642);
nor U36 (N_36,In_278,In_480);
and U37 (N_37,In_495,In_432);
or U38 (N_38,In_700,In_460);
and U39 (N_39,In_300,In_48);
or U40 (N_40,In_733,In_34);
and U41 (N_41,In_621,In_482);
and U42 (N_42,In_58,In_338);
nand U43 (N_43,In_250,In_674);
xnor U44 (N_44,In_281,In_748);
nand U45 (N_45,In_662,In_387);
and U46 (N_46,In_461,In_479);
nand U47 (N_47,In_380,In_22);
nor U48 (N_48,In_391,In_261);
or U49 (N_49,In_14,In_546);
and U50 (N_50,In_156,In_552);
nor U51 (N_51,In_583,In_739);
nor U52 (N_52,In_745,In_361);
nor U53 (N_53,In_470,In_628);
or U54 (N_54,In_69,In_288);
nor U55 (N_55,In_253,In_61);
nor U56 (N_56,In_503,In_125);
nor U57 (N_57,In_135,In_657);
nand U58 (N_58,In_453,In_118);
and U59 (N_59,In_274,In_695);
or U60 (N_60,In_477,In_272);
nand U61 (N_61,In_124,In_255);
or U62 (N_62,In_612,In_595);
nand U63 (N_63,In_55,In_18);
or U64 (N_64,In_339,In_499);
nand U65 (N_65,In_483,In_533);
or U66 (N_66,In_224,In_424);
nand U67 (N_67,In_264,In_409);
or U68 (N_68,In_590,In_506);
and U69 (N_69,In_410,In_248);
nand U70 (N_70,In_42,In_652);
and U71 (N_71,In_333,In_75);
nand U72 (N_72,In_260,In_358);
nor U73 (N_73,In_237,In_62);
and U74 (N_74,In_245,In_569);
nor U75 (N_75,In_66,In_522);
nor U76 (N_76,In_659,In_721);
or U77 (N_77,In_566,In_89);
nand U78 (N_78,In_103,In_712);
nand U79 (N_79,In_400,In_307);
nor U80 (N_80,In_517,In_238);
or U81 (N_81,In_266,In_498);
or U82 (N_82,In_405,In_451);
nand U83 (N_83,In_283,In_254);
nor U84 (N_84,In_267,In_464);
and U85 (N_85,In_234,In_618);
or U86 (N_86,In_666,In_184);
nor U87 (N_87,In_21,In_140);
and U88 (N_88,In_486,In_602);
nor U89 (N_89,In_23,In_169);
nand U90 (N_90,In_743,In_382);
or U91 (N_91,In_427,In_529);
nand U92 (N_92,In_49,In_205);
and U93 (N_93,In_701,In_271);
nor U94 (N_94,In_352,In_530);
nor U95 (N_95,In_112,In_218);
nand U96 (N_96,In_122,In_269);
or U97 (N_97,In_384,In_92);
nor U98 (N_98,In_228,In_604);
and U99 (N_99,In_10,In_420);
and U100 (N_100,In_678,In_141);
and U101 (N_101,In_322,In_235);
nor U102 (N_102,In_445,In_476);
or U103 (N_103,In_746,In_715);
nor U104 (N_104,In_344,In_672);
nor U105 (N_105,In_532,In_484);
and U106 (N_106,In_637,In_709);
nor U107 (N_107,In_154,In_45);
nor U108 (N_108,In_12,In_527);
nand U109 (N_109,In_513,In_421);
or U110 (N_110,In_656,In_364);
or U111 (N_111,In_611,In_321);
nand U112 (N_112,In_658,In_719);
or U113 (N_113,In_456,In_598);
or U114 (N_114,In_393,In_126);
and U115 (N_115,In_607,In_707);
nor U116 (N_116,In_578,In_720);
and U117 (N_117,In_681,In_641);
nand U118 (N_118,In_620,In_221);
nor U119 (N_119,In_181,In_402);
nor U120 (N_120,In_526,In_655);
and U121 (N_121,In_213,In_104);
and U122 (N_122,In_277,In_316);
and U123 (N_123,In_749,In_109);
nor U124 (N_124,In_175,In_207);
and U125 (N_125,In_349,In_106);
nor U126 (N_126,In_383,In_588);
nand U127 (N_127,In_56,In_206);
and U128 (N_128,In_121,In_183);
or U129 (N_129,In_727,In_113);
or U130 (N_130,In_403,In_587);
nor U131 (N_131,In_331,In_559);
or U132 (N_132,In_44,In_230);
and U133 (N_133,In_487,In_689);
or U134 (N_134,In_597,In_95);
and U135 (N_135,In_17,In_713);
nand U136 (N_136,In_728,In_345);
or U137 (N_137,In_448,In_653);
and U138 (N_138,In_372,In_747);
nor U139 (N_139,In_741,In_216);
nand U140 (N_140,In_340,In_504);
and U141 (N_141,In_665,In_663);
nor U142 (N_142,In_632,In_481);
nor U143 (N_143,In_220,In_654);
or U144 (N_144,In_397,In_192);
and U145 (N_145,In_176,In_469);
and U146 (N_146,In_493,In_80);
and U147 (N_147,In_680,In_514);
nand U148 (N_148,In_548,In_568);
and U149 (N_149,In_510,In_646);
and U150 (N_150,In_699,In_204);
nor U151 (N_151,In_236,In_645);
nand U152 (N_152,In_687,In_542);
nand U153 (N_153,In_317,In_537);
nand U154 (N_154,In_471,In_553);
nor U155 (N_155,In_593,In_614);
or U156 (N_156,In_373,In_289);
nor U157 (N_157,In_139,In_730);
nor U158 (N_158,In_462,In_459);
or U159 (N_159,In_217,In_38);
and U160 (N_160,In_442,In_341);
nor U161 (N_161,In_188,In_97);
and U162 (N_162,In_594,In_246);
nor U163 (N_163,In_390,In_688);
and U164 (N_164,In_225,In_544);
nand U165 (N_165,In_33,In_6);
or U166 (N_166,In_518,In_450);
nand U167 (N_167,In_19,In_512);
nand U168 (N_168,In_4,In_153);
xor U169 (N_169,In_294,In_65);
nor U170 (N_170,In_78,In_134);
nor U171 (N_171,In_564,In_584);
or U172 (N_172,In_475,In_634);
and U173 (N_173,In_609,In_738);
nand U174 (N_174,In_303,In_368);
or U175 (N_175,In_241,In_437);
or U176 (N_176,In_714,In_263);
or U177 (N_177,In_229,In_3);
or U178 (N_178,In_356,In_435);
nor U179 (N_179,In_744,In_543);
or U180 (N_180,In_540,In_474);
nand U181 (N_181,In_74,In_531);
nor U182 (N_182,In_516,In_166);
nand U183 (N_183,In_631,In_585);
and U184 (N_184,In_366,In_686);
and U185 (N_185,In_376,In_127);
and U186 (N_186,In_581,In_35);
and U187 (N_187,In_414,In_262);
nand U188 (N_188,In_473,In_36);
nand U189 (N_189,In_571,In_379);
nand U190 (N_190,In_693,In_640);
nand U191 (N_191,In_404,In_697);
nor U192 (N_192,In_93,In_444);
nor U193 (N_193,In_491,In_457);
and U194 (N_194,In_296,In_501);
nor U195 (N_195,In_615,In_187);
xor U196 (N_196,In_11,In_1);
nand U197 (N_197,In_485,In_72);
nor U198 (N_198,In_579,In_59);
and U199 (N_199,In_734,In_596);
nor U200 (N_200,In_79,In_399);
nand U201 (N_201,In_633,In_240);
nor U202 (N_202,In_244,In_377);
nand U203 (N_203,In_41,In_452);
nor U204 (N_204,In_575,In_32);
nand U205 (N_205,In_458,In_200);
and U206 (N_206,In_123,In_7);
nand U207 (N_207,In_179,In_73);
or U208 (N_208,In_203,In_592);
and U209 (N_209,In_441,In_648);
nand U210 (N_210,In_682,In_71);
or U211 (N_211,In_627,In_15);
and U212 (N_212,In_731,In_82);
and U213 (N_213,In_87,In_696);
or U214 (N_214,In_429,In_375);
nand U215 (N_215,In_64,In_115);
nor U216 (N_216,In_145,In_50);
nor U217 (N_217,In_367,In_117);
nand U218 (N_218,In_301,In_636);
nor U219 (N_219,In_305,In_419);
or U220 (N_220,In_233,In_554);
or U221 (N_221,In_555,In_116);
or U222 (N_222,In_25,In_425);
nand U223 (N_223,In_130,In_668);
or U224 (N_224,In_174,In_13);
nand U225 (N_225,In_430,In_60);
nor U226 (N_226,In_625,In_497);
and U227 (N_227,In_723,In_639);
nor U228 (N_228,In_243,In_535);
and U229 (N_229,In_500,In_463);
nor U230 (N_230,In_574,In_299);
and U231 (N_231,In_417,In_407);
and U232 (N_232,In_524,In_694);
and U233 (N_233,In_144,In_210);
and U234 (N_234,In_591,In_99);
and U235 (N_235,In_212,In_326);
and U236 (N_236,In_332,In_431);
and U237 (N_237,In_624,In_622);
and U238 (N_238,In_84,In_667);
or U239 (N_239,In_704,In_209);
and U240 (N_240,In_570,In_285);
or U241 (N_241,In_88,In_147);
nor U242 (N_242,In_194,In_550);
nor U243 (N_243,In_57,In_610);
nand U244 (N_244,In_690,In_100);
or U245 (N_245,In_398,In_679);
nand U246 (N_246,In_436,In_388);
and U247 (N_247,In_280,In_31);
or U248 (N_248,In_163,In_161);
or U249 (N_249,In_661,In_528);
nor U250 (N_250,In_198,In_323);
and U251 (N_251,In_313,In_386);
nor U252 (N_252,In_348,In_107);
nor U253 (N_253,In_547,In_511);
or U254 (N_254,In_576,In_443);
and U255 (N_255,In_494,In_385);
and U256 (N_256,In_302,In_310);
xor U257 (N_257,In_258,In_98);
nor U258 (N_258,In_315,In_465);
nand U259 (N_259,In_557,In_446);
nor U260 (N_260,In_111,In_702);
and U261 (N_261,In_219,In_197);
and U262 (N_262,In_351,In_691);
or U263 (N_263,In_318,In_705);
or U264 (N_264,In_509,In_626);
or U265 (N_265,In_328,In_297);
or U266 (N_266,In_692,In_282);
nor U267 (N_267,In_392,In_395);
and U268 (N_268,In_671,In_214);
and U269 (N_269,In_85,In_211);
nand U270 (N_270,In_157,In_582);
nor U271 (N_271,In_374,In_558);
and U272 (N_272,In_706,In_724);
or U273 (N_273,In_77,In_170);
nand U274 (N_274,In_729,In_586);
or U275 (N_275,In_573,In_68);
or U276 (N_276,In_20,In_478);
nand U277 (N_277,In_335,In_46);
or U278 (N_278,In_560,In_599);
or U279 (N_279,In_468,In_505);
nand U280 (N_280,In_94,In_9);
nor U281 (N_281,In_684,In_319);
nor U282 (N_282,In_490,In_39);
nor U283 (N_283,In_132,In_467);
or U284 (N_284,In_256,In_28);
or U285 (N_285,In_150,In_617);
or U286 (N_286,In_314,In_371);
and U287 (N_287,In_539,In_133);
nand U288 (N_288,In_359,In_515);
nor U289 (N_289,In_202,In_298);
and U290 (N_290,In_508,In_173);
and U291 (N_291,In_40,In_311);
and U292 (N_292,In_608,In_342);
and U293 (N_293,In_143,In_295);
and U294 (N_294,In_416,In_158);
or U295 (N_295,In_411,In_54);
or U296 (N_296,In_589,In_196);
and U297 (N_297,In_273,In_227);
or U298 (N_298,In_346,In_718);
nand U299 (N_299,In_616,In_378);
nand U300 (N_300,In_401,In_177);
nor U301 (N_301,In_447,In_136);
and U302 (N_302,In_434,In_148);
and U303 (N_303,In_191,In_52);
nor U304 (N_304,In_525,In_231);
nor U305 (N_305,In_171,In_673);
nor U306 (N_306,In_239,In_270);
or U307 (N_307,In_698,In_334);
nor U308 (N_308,In_725,In_370);
and U309 (N_309,In_545,In_551);
nand U310 (N_310,In_189,In_8);
nand U311 (N_311,In_128,In_119);
nor U312 (N_312,In_413,In_556);
or U313 (N_313,In_638,In_81);
or U314 (N_314,In_186,In_309);
and U315 (N_315,In_538,In_76);
nand U316 (N_316,In_129,In_330);
or U317 (N_317,In_449,In_353);
or U318 (N_318,In_350,In_519);
or U319 (N_319,In_347,In_265);
or U320 (N_320,In_369,In_222);
nor U321 (N_321,In_567,In_185);
or U322 (N_322,In_630,In_541);
nand U323 (N_323,In_290,In_428);
nand U324 (N_324,In_232,In_43);
or U325 (N_325,In_252,In_30);
or U326 (N_326,In_735,In_160);
or U327 (N_327,In_394,In_131);
nand U328 (N_328,In_561,In_96);
xnor U329 (N_329,In_406,In_242);
nor U330 (N_330,In_577,In_619);
or U331 (N_331,In_63,In_5);
and U332 (N_332,In_438,In_651);
nand U333 (N_333,In_664,In_455);
nor U334 (N_334,In_110,In_26);
nand U335 (N_335,In_320,In_312);
nor U336 (N_336,In_644,In_152);
or U337 (N_337,In_534,In_466);
or U338 (N_338,In_732,In_276);
or U339 (N_339,In_304,In_650);
or U340 (N_340,In_86,In_643);
nand U341 (N_341,In_492,In_108);
and U342 (N_342,In_726,In_138);
nand U343 (N_343,In_275,In_685);
nor U344 (N_344,In_114,In_572);
nand U345 (N_345,In_415,In_193);
and U346 (N_346,In_180,In_279);
nor U347 (N_347,In_605,In_496);
nand U348 (N_348,In_27,In_215);
and U349 (N_349,In_2,In_422);
nor U350 (N_350,In_565,In_507);
nor U351 (N_351,In_51,In_740);
nor U352 (N_352,In_67,In_549);
nor U353 (N_353,In_716,In_306);
nor U354 (N_354,In_412,In_16);
nor U355 (N_355,In_91,In_284);
nor U356 (N_356,In_329,In_606);
nor U357 (N_357,In_426,In_165);
xnor U358 (N_358,In_37,In_268);
or U359 (N_359,In_29,In_149);
nand U360 (N_360,In_603,In_363);
nor U361 (N_361,In_337,In_677);
or U362 (N_362,In_722,In_251);
nor U363 (N_363,In_142,In_660);
and U364 (N_364,In_389,In_600);
or U365 (N_365,In_472,In_336);
or U366 (N_366,In_623,In_563);
and U367 (N_367,In_190,In_164);
and U368 (N_368,In_259,In_601);
or U369 (N_369,In_257,In_536);
nand U370 (N_370,In_168,In_357);
or U371 (N_371,In_711,In_423);
nand U372 (N_372,In_0,In_710);
nand U373 (N_373,In_520,In_703);
nor U374 (N_374,In_324,In_178);
or U375 (N_375,In_129,In_557);
or U376 (N_376,In_327,In_229);
nor U377 (N_377,In_320,In_50);
nand U378 (N_378,In_409,In_328);
nand U379 (N_379,In_32,In_67);
nand U380 (N_380,In_660,In_110);
or U381 (N_381,In_233,In_4);
and U382 (N_382,In_695,In_229);
and U383 (N_383,In_675,In_99);
nor U384 (N_384,In_305,In_319);
nor U385 (N_385,In_739,In_277);
or U386 (N_386,In_71,In_207);
or U387 (N_387,In_424,In_609);
nor U388 (N_388,In_620,In_193);
nand U389 (N_389,In_277,In_692);
and U390 (N_390,In_223,In_339);
or U391 (N_391,In_453,In_345);
nor U392 (N_392,In_305,In_577);
or U393 (N_393,In_157,In_595);
nor U394 (N_394,In_379,In_422);
nand U395 (N_395,In_459,In_61);
nand U396 (N_396,In_518,In_662);
nand U397 (N_397,In_401,In_104);
and U398 (N_398,In_680,In_299);
or U399 (N_399,In_531,In_657);
and U400 (N_400,In_568,In_745);
and U401 (N_401,In_368,In_684);
or U402 (N_402,In_729,In_435);
nor U403 (N_403,In_205,In_354);
nand U404 (N_404,In_366,In_165);
or U405 (N_405,In_98,In_575);
nor U406 (N_406,In_88,In_302);
nor U407 (N_407,In_644,In_158);
nor U408 (N_408,In_218,In_554);
nand U409 (N_409,In_725,In_708);
and U410 (N_410,In_566,In_578);
or U411 (N_411,In_224,In_270);
nor U412 (N_412,In_174,In_517);
nand U413 (N_413,In_616,In_531);
and U414 (N_414,In_56,In_435);
nor U415 (N_415,In_542,In_214);
and U416 (N_416,In_610,In_744);
nor U417 (N_417,In_713,In_396);
and U418 (N_418,In_439,In_157);
nor U419 (N_419,In_554,In_418);
nand U420 (N_420,In_6,In_727);
nor U421 (N_421,In_610,In_651);
nand U422 (N_422,In_193,In_25);
nand U423 (N_423,In_216,In_562);
nor U424 (N_424,In_451,In_165);
or U425 (N_425,In_253,In_146);
nand U426 (N_426,In_246,In_359);
nand U427 (N_427,In_178,In_685);
or U428 (N_428,In_574,In_607);
nand U429 (N_429,In_601,In_674);
and U430 (N_430,In_732,In_52);
or U431 (N_431,In_365,In_141);
and U432 (N_432,In_60,In_593);
or U433 (N_433,In_219,In_86);
nand U434 (N_434,In_493,In_407);
or U435 (N_435,In_732,In_194);
or U436 (N_436,In_748,In_539);
nor U437 (N_437,In_725,In_335);
nand U438 (N_438,In_227,In_635);
nand U439 (N_439,In_460,In_485);
nor U440 (N_440,In_270,In_147);
and U441 (N_441,In_412,In_410);
or U442 (N_442,In_468,In_225);
nand U443 (N_443,In_111,In_193);
nand U444 (N_444,In_8,In_164);
nor U445 (N_445,In_523,In_540);
or U446 (N_446,In_374,In_604);
and U447 (N_447,In_96,In_338);
or U448 (N_448,In_245,In_496);
or U449 (N_449,In_220,In_65);
nand U450 (N_450,In_546,In_167);
and U451 (N_451,In_673,In_603);
or U452 (N_452,In_151,In_265);
or U453 (N_453,In_384,In_459);
nand U454 (N_454,In_96,In_466);
or U455 (N_455,In_307,In_258);
and U456 (N_456,In_256,In_600);
and U457 (N_457,In_112,In_193);
or U458 (N_458,In_188,In_254);
nand U459 (N_459,In_80,In_32);
nand U460 (N_460,In_49,In_712);
or U461 (N_461,In_467,In_455);
nor U462 (N_462,In_729,In_714);
nor U463 (N_463,In_96,In_365);
and U464 (N_464,In_378,In_623);
and U465 (N_465,In_330,In_613);
nor U466 (N_466,In_26,In_314);
nand U467 (N_467,In_50,In_121);
nor U468 (N_468,In_510,In_38);
nor U469 (N_469,In_160,In_213);
or U470 (N_470,In_117,In_198);
or U471 (N_471,In_423,In_249);
nor U472 (N_472,In_208,In_9);
nand U473 (N_473,In_114,In_299);
and U474 (N_474,In_682,In_331);
or U475 (N_475,In_446,In_352);
or U476 (N_476,In_20,In_589);
or U477 (N_477,In_357,In_331);
and U478 (N_478,In_204,In_746);
nand U479 (N_479,In_674,In_648);
or U480 (N_480,In_547,In_98);
nor U481 (N_481,In_7,In_380);
nor U482 (N_482,In_673,In_279);
nor U483 (N_483,In_107,In_316);
or U484 (N_484,In_496,In_285);
xnor U485 (N_485,In_358,In_550);
and U486 (N_486,In_577,In_636);
and U487 (N_487,In_117,In_186);
and U488 (N_488,In_68,In_445);
or U489 (N_489,In_498,In_651);
and U490 (N_490,In_563,In_402);
nand U491 (N_491,In_167,In_261);
nor U492 (N_492,In_447,In_39);
nor U493 (N_493,In_199,In_331);
or U494 (N_494,In_299,In_204);
and U495 (N_495,In_353,In_242);
nor U496 (N_496,In_388,In_331);
nor U497 (N_497,In_525,In_425);
or U498 (N_498,In_312,In_12);
and U499 (N_499,In_547,In_352);
and U500 (N_500,N_487,N_304);
and U501 (N_501,N_65,N_414);
nand U502 (N_502,N_183,N_457);
and U503 (N_503,N_30,N_403);
or U504 (N_504,N_300,N_164);
nor U505 (N_505,N_150,N_413);
or U506 (N_506,N_353,N_165);
nand U507 (N_507,N_21,N_205);
nor U508 (N_508,N_73,N_134);
or U509 (N_509,N_110,N_285);
nand U510 (N_510,N_376,N_105);
and U511 (N_511,N_286,N_323);
nor U512 (N_512,N_405,N_60);
or U513 (N_513,N_120,N_404);
and U514 (N_514,N_426,N_228);
nand U515 (N_515,N_423,N_31);
nand U516 (N_516,N_495,N_425);
and U517 (N_517,N_123,N_187);
or U518 (N_518,N_95,N_329);
nor U519 (N_519,N_80,N_239);
nand U520 (N_520,N_58,N_320);
and U521 (N_521,N_339,N_305);
nand U522 (N_522,N_484,N_282);
nor U523 (N_523,N_59,N_342);
nand U524 (N_524,N_326,N_447);
and U525 (N_525,N_335,N_365);
or U526 (N_526,N_398,N_399);
nor U527 (N_527,N_433,N_108);
or U528 (N_528,N_200,N_49);
or U529 (N_529,N_464,N_406);
or U530 (N_530,N_453,N_470);
and U531 (N_531,N_211,N_126);
or U532 (N_532,N_374,N_369);
or U533 (N_533,N_332,N_462);
or U534 (N_534,N_328,N_161);
nand U535 (N_535,N_131,N_477);
and U536 (N_536,N_74,N_273);
nand U537 (N_537,N_391,N_140);
nor U538 (N_538,N_142,N_288);
nor U539 (N_539,N_209,N_368);
and U540 (N_540,N_124,N_195);
nor U541 (N_541,N_159,N_54);
nor U542 (N_542,N_136,N_192);
and U543 (N_543,N_361,N_51);
and U544 (N_544,N_83,N_264);
and U545 (N_545,N_352,N_307);
and U546 (N_546,N_38,N_390);
or U547 (N_547,N_483,N_363);
nor U548 (N_548,N_162,N_325);
nor U549 (N_549,N_291,N_217);
nand U550 (N_550,N_212,N_292);
and U551 (N_551,N_468,N_154);
or U552 (N_552,N_249,N_415);
nand U553 (N_553,N_71,N_82);
nor U554 (N_554,N_461,N_4);
or U555 (N_555,N_170,N_394);
nand U556 (N_556,N_392,N_400);
or U557 (N_557,N_283,N_254);
or U558 (N_558,N_15,N_189);
nand U559 (N_559,N_272,N_245);
and U560 (N_560,N_367,N_432);
nand U561 (N_561,N_451,N_106);
and U562 (N_562,N_77,N_175);
nor U563 (N_563,N_160,N_107);
nor U564 (N_564,N_303,N_445);
nor U565 (N_565,N_206,N_301);
nand U566 (N_566,N_338,N_50);
xor U567 (N_567,N_166,N_492);
nand U568 (N_568,N_144,N_346);
nor U569 (N_569,N_318,N_455);
xor U570 (N_570,N_100,N_355);
or U571 (N_571,N_449,N_78);
or U572 (N_572,N_459,N_358);
nor U573 (N_573,N_137,N_472);
or U574 (N_574,N_316,N_475);
or U575 (N_575,N_8,N_479);
or U576 (N_576,N_176,N_424);
and U577 (N_577,N_310,N_357);
or U578 (N_578,N_334,N_17);
nand U579 (N_579,N_446,N_379);
and U580 (N_580,N_155,N_204);
or U581 (N_581,N_135,N_256);
or U582 (N_582,N_488,N_220);
nor U583 (N_583,N_79,N_247);
or U584 (N_584,N_42,N_218);
and U585 (N_585,N_222,N_86);
or U586 (N_586,N_485,N_437);
nor U587 (N_587,N_333,N_314);
and U588 (N_588,N_321,N_349);
or U589 (N_589,N_362,N_72);
nor U590 (N_590,N_194,N_360);
or U591 (N_591,N_93,N_274);
or U592 (N_592,N_198,N_2);
nand U593 (N_593,N_97,N_319);
or U594 (N_594,N_240,N_260);
nor U595 (N_595,N_372,N_177);
nand U596 (N_596,N_439,N_47);
or U597 (N_597,N_13,N_190);
and U598 (N_598,N_19,N_486);
or U599 (N_599,N_337,N_104);
or U600 (N_600,N_243,N_389);
xnor U601 (N_601,N_10,N_48);
and U602 (N_602,N_213,N_186);
or U603 (N_603,N_490,N_45);
nand U604 (N_604,N_474,N_378);
or U605 (N_605,N_241,N_179);
nor U606 (N_606,N_441,N_172);
or U607 (N_607,N_132,N_43);
nand U608 (N_608,N_387,N_364);
and U609 (N_609,N_356,N_436);
or U610 (N_610,N_122,N_253);
and U611 (N_611,N_109,N_227);
and U612 (N_612,N_296,N_75);
nor U613 (N_613,N_295,N_147);
or U614 (N_614,N_157,N_489);
nor U615 (N_615,N_22,N_202);
nand U616 (N_616,N_450,N_336);
nor U617 (N_617,N_199,N_235);
xor U618 (N_618,N_149,N_129);
or U619 (N_619,N_299,N_70);
nand U620 (N_620,N_112,N_163);
or U621 (N_621,N_309,N_422);
nand U622 (N_622,N_234,N_182);
or U623 (N_623,N_481,N_252);
nand U624 (N_624,N_215,N_366);
and U625 (N_625,N_61,N_324);
nand U626 (N_626,N_69,N_139);
nor U627 (N_627,N_36,N_354);
nand U628 (N_628,N_0,N_258);
or U629 (N_629,N_87,N_133);
nor U630 (N_630,N_128,N_44);
or U631 (N_631,N_259,N_40);
nand U632 (N_632,N_238,N_233);
and U633 (N_633,N_277,N_178);
or U634 (N_634,N_152,N_67);
nor U635 (N_635,N_236,N_345);
or U636 (N_636,N_409,N_418);
or U637 (N_637,N_6,N_298);
and U638 (N_638,N_55,N_18);
or U639 (N_639,N_435,N_293);
nor U640 (N_640,N_203,N_452);
and U641 (N_641,N_223,N_262);
and U642 (N_642,N_121,N_471);
and U643 (N_643,N_276,N_116);
xor U644 (N_644,N_383,N_440);
nor U645 (N_645,N_429,N_28);
nand U646 (N_646,N_76,N_208);
and U647 (N_647,N_89,N_99);
nand U648 (N_648,N_279,N_41);
and U649 (N_649,N_322,N_494);
nand U650 (N_650,N_499,N_32);
nand U651 (N_651,N_221,N_347);
nand U652 (N_652,N_327,N_119);
or U653 (N_653,N_251,N_113);
or U654 (N_654,N_226,N_380);
nor U655 (N_655,N_350,N_115);
and U656 (N_656,N_313,N_156);
and U657 (N_657,N_52,N_85);
or U658 (N_658,N_180,N_396);
and U659 (N_659,N_225,N_145);
or U660 (N_660,N_456,N_171);
and U661 (N_661,N_306,N_88);
nor U662 (N_662,N_1,N_386);
xor U663 (N_663,N_434,N_444);
or U664 (N_664,N_498,N_12);
and U665 (N_665,N_14,N_469);
nor U666 (N_666,N_497,N_5);
and U667 (N_667,N_66,N_269);
nand U668 (N_668,N_385,N_261);
and U669 (N_669,N_402,N_458);
nor U670 (N_670,N_33,N_188);
or U671 (N_671,N_242,N_57);
xor U672 (N_672,N_141,N_416);
or U673 (N_673,N_63,N_377);
nor U674 (N_674,N_181,N_270);
nand U675 (N_675,N_427,N_463);
nand U676 (N_676,N_25,N_267);
nand U677 (N_677,N_493,N_90);
xor U678 (N_678,N_118,N_53);
and U679 (N_679,N_169,N_397);
or U680 (N_680,N_248,N_173);
or U681 (N_681,N_407,N_35);
nand U682 (N_682,N_401,N_257);
or U683 (N_683,N_294,N_230);
nor U684 (N_684,N_168,N_11);
or U685 (N_685,N_417,N_265);
or U686 (N_686,N_7,N_284);
or U687 (N_687,N_20,N_193);
or U688 (N_688,N_56,N_410);
nor U689 (N_689,N_370,N_34);
nand U690 (N_690,N_197,N_102);
nand U691 (N_691,N_411,N_68);
xnor U692 (N_692,N_81,N_117);
or U693 (N_693,N_454,N_64);
or U694 (N_694,N_185,N_315);
nand U695 (N_695,N_37,N_311);
nand U696 (N_696,N_229,N_207);
nand U697 (N_697,N_281,N_3);
nor U698 (N_698,N_382,N_84);
nor U699 (N_699,N_148,N_359);
or U700 (N_700,N_196,N_375);
nor U701 (N_701,N_393,N_174);
and U702 (N_702,N_146,N_101);
nor U703 (N_703,N_419,N_289);
or U704 (N_704,N_16,N_430);
or U705 (N_705,N_224,N_341);
nor U706 (N_706,N_98,N_351);
nor U707 (N_707,N_478,N_278);
and U708 (N_708,N_94,N_467);
or U709 (N_709,N_143,N_91);
nor U710 (N_710,N_473,N_24);
and U711 (N_711,N_214,N_448);
nor U712 (N_712,N_330,N_125);
nor U713 (N_713,N_395,N_158);
nand U714 (N_714,N_312,N_280);
nand U715 (N_715,N_219,N_412);
nor U716 (N_716,N_482,N_237);
nor U717 (N_717,N_428,N_191);
nor U718 (N_718,N_331,N_476);
nand U719 (N_719,N_62,N_96);
or U720 (N_720,N_271,N_343);
nor U721 (N_721,N_348,N_460);
and U722 (N_722,N_268,N_167);
or U723 (N_723,N_431,N_151);
or U724 (N_724,N_421,N_340);
or U725 (N_725,N_153,N_302);
and U726 (N_726,N_111,N_266);
nand U727 (N_727,N_92,N_438);
or U728 (N_728,N_184,N_275);
and U729 (N_729,N_114,N_216);
nand U730 (N_730,N_420,N_138);
nand U731 (N_731,N_384,N_381);
nand U732 (N_732,N_491,N_231);
nand U733 (N_733,N_297,N_210);
nor U734 (N_734,N_290,N_496);
nor U735 (N_735,N_103,N_443);
or U736 (N_736,N_466,N_373);
nor U737 (N_737,N_127,N_371);
and U738 (N_738,N_26,N_344);
and U739 (N_739,N_308,N_263);
nor U740 (N_740,N_480,N_27);
nor U741 (N_741,N_46,N_29);
nand U742 (N_742,N_232,N_201);
and U743 (N_743,N_39,N_246);
nor U744 (N_744,N_388,N_317);
nand U745 (N_745,N_9,N_287);
and U746 (N_746,N_244,N_255);
and U747 (N_747,N_130,N_442);
nand U748 (N_748,N_408,N_250);
nand U749 (N_749,N_23,N_465);
and U750 (N_750,N_316,N_335);
nand U751 (N_751,N_234,N_72);
nor U752 (N_752,N_495,N_179);
or U753 (N_753,N_399,N_236);
or U754 (N_754,N_403,N_32);
or U755 (N_755,N_27,N_424);
or U756 (N_756,N_352,N_347);
and U757 (N_757,N_277,N_397);
nand U758 (N_758,N_41,N_412);
nand U759 (N_759,N_277,N_268);
or U760 (N_760,N_41,N_221);
nand U761 (N_761,N_233,N_0);
nor U762 (N_762,N_156,N_97);
nor U763 (N_763,N_479,N_260);
nor U764 (N_764,N_132,N_153);
nor U765 (N_765,N_58,N_221);
and U766 (N_766,N_394,N_96);
or U767 (N_767,N_69,N_342);
nand U768 (N_768,N_32,N_345);
nor U769 (N_769,N_470,N_142);
or U770 (N_770,N_411,N_230);
and U771 (N_771,N_330,N_458);
and U772 (N_772,N_236,N_431);
and U773 (N_773,N_270,N_437);
or U774 (N_774,N_362,N_335);
and U775 (N_775,N_156,N_461);
and U776 (N_776,N_461,N_309);
and U777 (N_777,N_355,N_416);
or U778 (N_778,N_76,N_132);
xor U779 (N_779,N_45,N_453);
and U780 (N_780,N_55,N_41);
and U781 (N_781,N_470,N_250);
and U782 (N_782,N_85,N_11);
nor U783 (N_783,N_453,N_391);
nand U784 (N_784,N_105,N_284);
nand U785 (N_785,N_350,N_149);
nand U786 (N_786,N_454,N_170);
or U787 (N_787,N_244,N_475);
nand U788 (N_788,N_188,N_179);
or U789 (N_789,N_53,N_389);
and U790 (N_790,N_106,N_170);
and U791 (N_791,N_469,N_290);
or U792 (N_792,N_352,N_103);
nor U793 (N_793,N_454,N_32);
nand U794 (N_794,N_267,N_313);
or U795 (N_795,N_290,N_168);
nor U796 (N_796,N_419,N_267);
or U797 (N_797,N_249,N_426);
and U798 (N_798,N_372,N_496);
nor U799 (N_799,N_26,N_27);
and U800 (N_800,N_342,N_359);
or U801 (N_801,N_482,N_360);
nor U802 (N_802,N_158,N_201);
nand U803 (N_803,N_434,N_375);
xor U804 (N_804,N_345,N_163);
nor U805 (N_805,N_63,N_68);
and U806 (N_806,N_102,N_294);
and U807 (N_807,N_364,N_422);
nand U808 (N_808,N_170,N_248);
nand U809 (N_809,N_190,N_302);
and U810 (N_810,N_284,N_431);
or U811 (N_811,N_172,N_247);
nand U812 (N_812,N_192,N_316);
nor U813 (N_813,N_363,N_361);
nor U814 (N_814,N_153,N_241);
nor U815 (N_815,N_493,N_4);
nand U816 (N_816,N_431,N_115);
nand U817 (N_817,N_192,N_378);
nor U818 (N_818,N_66,N_43);
nand U819 (N_819,N_382,N_378);
or U820 (N_820,N_350,N_171);
or U821 (N_821,N_220,N_149);
and U822 (N_822,N_244,N_320);
or U823 (N_823,N_89,N_358);
or U824 (N_824,N_308,N_387);
or U825 (N_825,N_222,N_2);
nand U826 (N_826,N_78,N_238);
nand U827 (N_827,N_434,N_376);
or U828 (N_828,N_151,N_489);
and U829 (N_829,N_312,N_190);
and U830 (N_830,N_202,N_31);
and U831 (N_831,N_457,N_199);
and U832 (N_832,N_406,N_238);
and U833 (N_833,N_316,N_180);
nand U834 (N_834,N_358,N_91);
nand U835 (N_835,N_233,N_96);
nand U836 (N_836,N_456,N_289);
nand U837 (N_837,N_379,N_309);
nor U838 (N_838,N_331,N_233);
and U839 (N_839,N_446,N_293);
or U840 (N_840,N_65,N_495);
nor U841 (N_841,N_461,N_315);
or U842 (N_842,N_272,N_459);
and U843 (N_843,N_432,N_134);
nor U844 (N_844,N_286,N_85);
or U845 (N_845,N_377,N_253);
or U846 (N_846,N_301,N_27);
nor U847 (N_847,N_418,N_106);
and U848 (N_848,N_387,N_298);
nor U849 (N_849,N_156,N_358);
and U850 (N_850,N_310,N_331);
and U851 (N_851,N_152,N_445);
and U852 (N_852,N_335,N_60);
or U853 (N_853,N_220,N_340);
and U854 (N_854,N_404,N_30);
or U855 (N_855,N_251,N_84);
nand U856 (N_856,N_12,N_151);
and U857 (N_857,N_297,N_396);
nor U858 (N_858,N_441,N_109);
nor U859 (N_859,N_485,N_338);
and U860 (N_860,N_397,N_481);
and U861 (N_861,N_74,N_240);
or U862 (N_862,N_387,N_254);
nor U863 (N_863,N_60,N_339);
nand U864 (N_864,N_167,N_484);
nand U865 (N_865,N_254,N_39);
nand U866 (N_866,N_428,N_36);
and U867 (N_867,N_77,N_72);
and U868 (N_868,N_370,N_42);
or U869 (N_869,N_169,N_487);
nand U870 (N_870,N_337,N_199);
and U871 (N_871,N_388,N_411);
nor U872 (N_872,N_76,N_128);
nand U873 (N_873,N_309,N_426);
and U874 (N_874,N_103,N_458);
nor U875 (N_875,N_297,N_427);
and U876 (N_876,N_438,N_159);
nand U877 (N_877,N_470,N_80);
or U878 (N_878,N_102,N_321);
or U879 (N_879,N_449,N_198);
or U880 (N_880,N_131,N_319);
nor U881 (N_881,N_170,N_480);
nor U882 (N_882,N_321,N_10);
nor U883 (N_883,N_475,N_499);
and U884 (N_884,N_225,N_369);
nor U885 (N_885,N_239,N_18);
nand U886 (N_886,N_389,N_32);
nor U887 (N_887,N_232,N_51);
and U888 (N_888,N_293,N_258);
nand U889 (N_889,N_376,N_397);
or U890 (N_890,N_68,N_30);
or U891 (N_891,N_176,N_34);
and U892 (N_892,N_492,N_363);
nor U893 (N_893,N_259,N_401);
and U894 (N_894,N_245,N_465);
nand U895 (N_895,N_147,N_33);
or U896 (N_896,N_279,N_166);
and U897 (N_897,N_190,N_10);
and U898 (N_898,N_337,N_437);
nand U899 (N_899,N_21,N_457);
nor U900 (N_900,N_280,N_175);
or U901 (N_901,N_306,N_350);
or U902 (N_902,N_270,N_245);
nor U903 (N_903,N_191,N_194);
nand U904 (N_904,N_414,N_146);
nor U905 (N_905,N_162,N_461);
or U906 (N_906,N_63,N_462);
nor U907 (N_907,N_68,N_256);
or U908 (N_908,N_355,N_59);
or U909 (N_909,N_483,N_370);
or U910 (N_910,N_447,N_371);
or U911 (N_911,N_194,N_253);
nor U912 (N_912,N_89,N_253);
nand U913 (N_913,N_115,N_226);
nor U914 (N_914,N_177,N_323);
nand U915 (N_915,N_261,N_73);
or U916 (N_916,N_61,N_28);
and U917 (N_917,N_331,N_159);
and U918 (N_918,N_21,N_204);
nor U919 (N_919,N_293,N_248);
nor U920 (N_920,N_201,N_27);
nor U921 (N_921,N_25,N_234);
or U922 (N_922,N_108,N_486);
or U923 (N_923,N_9,N_278);
nand U924 (N_924,N_225,N_490);
nand U925 (N_925,N_385,N_32);
or U926 (N_926,N_102,N_415);
or U927 (N_927,N_230,N_129);
nor U928 (N_928,N_100,N_146);
nor U929 (N_929,N_50,N_75);
or U930 (N_930,N_397,N_93);
or U931 (N_931,N_499,N_217);
or U932 (N_932,N_93,N_49);
or U933 (N_933,N_80,N_391);
nand U934 (N_934,N_328,N_416);
nor U935 (N_935,N_352,N_164);
and U936 (N_936,N_132,N_350);
nand U937 (N_937,N_141,N_386);
nor U938 (N_938,N_221,N_497);
nor U939 (N_939,N_151,N_212);
nand U940 (N_940,N_445,N_221);
and U941 (N_941,N_183,N_415);
nor U942 (N_942,N_33,N_356);
or U943 (N_943,N_260,N_78);
and U944 (N_944,N_414,N_351);
or U945 (N_945,N_452,N_82);
or U946 (N_946,N_168,N_432);
nand U947 (N_947,N_416,N_491);
and U948 (N_948,N_286,N_187);
nor U949 (N_949,N_88,N_141);
or U950 (N_950,N_163,N_494);
or U951 (N_951,N_53,N_444);
and U952 (N_952,N_213,N_336);
nor U953 (N_953,N_490,N_221);
or U954 (N_954,N_126,N_242);
nand U955 (N_955,N_228,N_266);
or U956 (N_956,N_121,N_455);
nor U957 (N_957,N_406,N_283);
nor U958 (N_958,N_367,N_349);
and U959 (N_959,N_188,N_118);
nand U960 (N_960,N_148,N_480);
nand U961 (N_961,N_442,N_89);
nand U962 (N_962,N_385,N_34);
or U963 (N_963,N_304,N_209);
nor U964 (N_964,N_467,N_359);
and U965 (N_965,N_308,N_413);
or U966 (N_966,N_34,N_50);
xor U967 (N_967,N_419,N_126);
nand U968 (N_968,N_354,N_62);
and U969 (N_969,N_238,N_288);
and U970 (N_970,N_418,N_42);
nor U971 (N_971,N_421,N_406);
and U972 (N_972,N_316,N_387);
nor U973 (N_973,N_172,N_298);
and U974 (N_974,N_464,N_222);
and U975 (N_975,N_383,N_69);
nand U976 (N_976,N_316,N_67);
and U977 (N_977,N_86,N_366);
nand U978 (N_978,N_337,N_194);
nor U979 (N_979,N_349,N_486);
nand U980 (N_980,N_28,N_38);
nor U981 (N_981,N_138,N_152);
nand U982 (N_982,N_397,N_49);
nor U983 (N_983,N_26,N_64);
and U984 (N_984,N_390,N_253);
or U985 (N_985,N_480,N_442);
or U986 (N_986,N_335,N_313);
nand U987 (N_987,N_281,N_78);
and U988 (N_988,N_64,N_338);
and U989 (N_989,N_34,N_183);
nand U990 (N_990,N_441,N_150);
nand U991 (N_991,N_140,N_102);
and U992 (N_992,N_114,N_471);
nor U993 (N_993,N_403,N_466);
or U994 (N_994,N_225,N_231);
or U995 (N_995,N_450,N_301);
or U996 (N_996,N_430,N_415);
or U997 (N_997,N_70,N_262);
or U998 (N_998,N_454,N_414);
or U999 (N_999,N_153,N_433);
nor U1000 (N_1000,N_904,N_762);
nand U1001 (N_1001,N_502,N_874);
nor U1002 (N_1002,N_801,N_960);
or U1003 (N_1003,N_720,N_846);
nand U1004 (N_1004,N_728,N_527);
nor U1005 (N_1005,N_973,N_648);
nand U1006 (N_1006,N_741,N_954);
nor U1007 (N_1007,N_659,N_767);
nand U1008 (N_1008,N_630,N_522);
nor U1009 (N_1009,N_573,N_740);
nand U1010 (N_1010,N_884,N_508);
and U1011 (N_1011,N_634,N_805);
nor U1012 (N_1012,N_707,N_618);
nor U1013 (N_1013,N_706,N_709);
nor U1014 (N_1014,N_865,N_557);
or U1015 (N_1015,N_896,N_887);
nand U1016 (N_1016,N_732,N_932);
and U1017 (N_1017,N_673,N_772);
or U1018 (N_1018,N_743,N_918);
nand U1019 (N_1019,N_638,N_962);
or U1020 (N_1020,N_753,N_696);
or U1021 (N_1021,N_705,N_770);
nand U1022 (N_1022,N_951,N_632);
and U1023 (N_1023,N_543,N_604);
nor U1024 (N_1024,N_524,N_730);
nand U1025 (N_1025,N_978,N_941);
or U1026 (N_1026,N_729,N_867);
nor U1027 (N_1027,N_711,N_553);
xnor U1028 (N_1028,N_796,N_652);
or U1029 (N_1029,N_975,N_986);
nor U1030 (N_1030,N_777,N_945);
nand U1031 (N_1031,N_763,N_776);
or U1032 (N_1032,N_703,N_654);
nor U1033 (N_1033,N_828,N_566);
nand U1034 (N_1034,N_784,N_526);
nand U1035 (N_1035,N_597,N_506);
or U1036 (N_1036,N_864,N_658);
nor U1037 (N_1037,N_518,N_641);
nand U1038 (N_1038,N_688,N_861);
nand U1039 (N_1039,N_797,N_644);
or U1040 (N_1040,N_523,N_882);
or U1041 (N_1041,N_555,N_546);
nor U1042 (N_1042,N_934,N_745);
nand U1043 (N_1043,N_656,N_579);
nand U1044 (N_1044,N_869,N_625);
or U1045 (N_1045,N_627,N_739);
nor U1046 (N_1046,N_970,N_662);
or U1047 (N_1047,N_542,N_930);
and U1048 (N_1048,N_999,N_534);
nand U1049 (N_1049,N_830,N_544);
or U1050 (N_1050,N_742,N_853);
and U1051 (N_1051,N_812,N_750);
and U1052 (N_1052,N_606,N_842);
or U1053 (N_1053,N_645,N_775);
nand U1054 (N_1054,N_898,N_953);
and U1055 (N_1055,N_541,N_552);
nand U1056 (N_1056,N_833,N_909);
nor U1057 (N_1057,N_794,N_948);
or U1058 (N_1058,N_836,N_871);
nor U1059 (N_1059,N_961,N_571);
and U1060 (N_1060,N_577,N_787);
or U1061 (N_1061,N_890,N_969);
nor U1062 (N_1062,N_949,N_708);
nand U1063 (N_1063,N_854,N_609);
nand U1064 (N_1064,N_879,N_968);
and U1065 (N_1065,N_799,N_614);
nor U1066 (N_1066,N_868,N_572);
or U1067 (N_1067,N_907,N_878);
nor U1068 (N_1068,N_860,N_576);
nand U1069 (N_1069,N_859,N_674);
and U1070 (N_1070,N_806,N_780);
or U1071 (N_1071,N_605,N_990);
nand U1072 (N_1072,N_870,N_501);
nand U1073 (N_1073,N_533,N_849);
or U1074 (N_1074,N_624,N_623);
and U1075 (N_1075,N_760,N_781);
and U1076 (N_1076,N_798,N_845);
and U1077 (N_1077,N_839,N_565);
and U1078 (N_1078,N_642,N_992);
nand U1079 (N_1079,N_827,N_923);
nand U1080 (N_1080,N_795,N_966);
and U1081 (N_1081,N_681,N_710);
and U1082 (N_1082,N_704,N_835);
nor U1083 (N_1083,N_880,N_578);
nand U1084 (N_1084,N_899,N_788);
nand U1085 (N_1085,N_718,N_831);
nor U1086 (N_1086,N_944,N_569);
nand U1087 (N_1087,N_723,N_619);
or U1088 (N_1088,N_976,N_995);
and U1089 (N_1089,N_936,N_749);
xnor U1090 (N_1090,N_758,N_851);
and U1091 (N_1091,N_620,N_615);
nand U1092 (N_1092,N_549,N_537);
or U1093 (N_1093,N_816,N_922);
nor U1094 (N_1094,N_939,N_668);
or U1095 (N_1095,N_545,N_778);
nor U1096 (N_1096,N_792,N_785);
and U1097 (N_1097,N_691,N_687);
nor U1098 (N_1098,N_856,N_626);
and U1099 (N_1099,N_832,N_616);
nand U1100 (N_1100,N_829,N_719);
nor U1101 (N_1101,N_988,N_809);
nor U1102 (N_1102,N_554,N_751);
or U1103 (N_1103,N_893,N_540);
nor U1104 (N_1104,N_724,N_580);
and U1105 (N_1105,N_629,N_950);
and U1106 (N_1106,N_981,N_804);
and U1107 (N_1107,N_929,N_538);
nand U1108 (N_1108,N_693,N_803);
and U1109 (N_1109,N_591,N_581);
or U1110 (N_1110,N_905,N_808);
or U1111 (N_1111,N_562,N_759);
and U1112 (N_1112,N_505,N_737);
or U1113 (N_1113,N_983,N_752);
or U1114 (N_1114,N_985,N_998);
or U1115 (N_1115,N_660,N_727);
nor U1116 (N_1116,N_952,N_684);
or U1117 (N_1117,N_601,N_955);
or U1118 (N_1118,N_570,N_586);
and U1119 (N_1119,N_611,N_957);
nor U1120 (N_1120,N_560,N_735);
or U1121 (N_1121,N_593,N_789);
nor U1122 (N_1122,N_574,N_612);
or U1123 (N_1123,N_974,N_682);
nor U1124 (N_1124,N_825,N_940);
nand U1125 (N_1125,N_590,N_771);
and U1126 (N_1126,N_663,N_819);
nor U1127 (N_1127,N_664,N_779);
nand U1128 (N_1128,N_547,N_669);
nor U1129 (N_1129,N_643,N_513);
and U1130 (N_1130,N_733,N_714);
or U1131 (N_1131,N_702,N_734);
nand U1132 (N_1132,N_509,N_933);
or U1133 (N_1133,N_588,N_889);
and U1134 (N_1134,N_598,N_550);
and U1135 (N_1135,N_584,N_912);
nor U1136 (N_1136,N_989,N_903);
and U1137 (N_1137,N_919,N_608);
nor U1138 (N_1138,N_843,N_655);
and U1139 (N_1139,N_726,N_971);
nor U1140 (N_1140,N_521,N_906);
nor U1141 (N_1141,N_877,N_525);
nor U1142 (N_1142,N_997,N_722);
nand U1143 (N_1143,N_633,N_820);
xnor U1144 (N_1144,N_921,N_814);
nand U1145 (N_1145,N_866,N_564);
or U1146 (N_1146,N_510,N_563);
and U1147 (N_1147,N_972,N_786);
nor U1148 (N_1148,N_858,N_535);
nand U1149 (N_1149,N_585,N_716);
and U1150 (N_1150,N_862,N_942);
or U1151 (N_1151,N_979,N_617);
nor U1152 (N_1152,N_755,N_665);
and U1153 (N_1153,N_667,N_567);
and U1154 (N_1154,N_791,N_528);
nand U1155 (N_1155,N_937,N_685);
and U1156 (N_1156,N_511,N_602);
and U1157 (N_1157,N_982,N_900);
and U1158 (N_1158,N_556,N_531);
and U1159 (N_1159,N_977,N_765);
or U1160 (N_1160,N_913,N_712);
nand U1161 (N_1161,N_818,N_875);
or U1162 (N_1162,N_947,N_639);
and U1163 (N_1163,N_744,N_500);
nand U1164 (N_1164,N_914,N_679);
nand U1165 (N_1165,N_507,N_517);
nand U1166 (N_1166,N_911,N_915);
and U1167 (N_1167,N_583,N_902);
nor U1168 (N_1168,N_761,N_873);
nand U1169 (N_1169,N_698,N_686);
nor U1170 (N_1170,N_603,N_876);
and U1171 (N_1171,N_766,N_844);
or U1172 (N_1172,N_613,N_807);
nand U1173 (N_1173,N_910,N_764);
or U1174 (N_1174,N_647,N_916);
nor U1175 (N_1175,N_888,N_840);
and U1176 (N_1176,N_512,N_848);
or U1177 (N_1177,N_993,N_946);
and U1178 (N_1178,N_748,N_607);
nor U1179 (N_1179,N_895,N_599);
nor U1180 (N_1180,N_754,N_721);
nor U1181 (N_1181,N_938,N_782);
and U1182 (N_1182,N_595,N_813);
nand U1183 (N_1183,N_589,N_823);
nor U1184 (N_1184,N_925,N_943);
or U1185 (N_1185,N_725,N_697);
and U1186 (N_1186,N_891,N_640);
nor U1187 (N_1187,N_649,N_596);
nand U1188 (N_1188,N_855,N_678);
and U1189 (N_1189,N_756,N_575);
nand U1190 (N_1190,N_610,N_559);
nor U1191 (N_1191,N_582,N_987);
nand U1192 (N_1192,N_935,N_920);
nand U1193 (N_1193,N_991,N_815);
or U1194 (N_1194,N_959,N_551);
nand U1195 (N_1195,N_783,N_967);
and U1196 (N_1196,N_746,N_558);
nand U1197 (N_1197,N_671,N_773);
nand U1198 (N_1198,N_532,N_863);
nor U1199 (N_1199,N_637,N_817);
nor U1200 (N_1200,N_837,N_631);
nand U1201 (N_1201,N_927,N_885);
and U1202 (N_1202,N_768,N_680);
or U1203 (N_1203,N_715,N_568);
nor U1204 (N_1204,N_515,N_731);
or U1205 (N_1205,N_519,N_872);
xor U1206 (N_1206,N_826,N_653);
or U1207 (N_1207,N_802,N_651);
and U1208 (N_1208,N_931,N_892);
nor U1209 (N_1209,N_881,N_713);
and U1210 (N_1210,N_736,N_822);
and U1211 (N_1211,N_883,N_901);
or U1212 (N_1212,N_897,N_963);
nand U1213 (N_1213,N_657,N_757);
nor U1214 (N_1214,N_592,N_850);
or U1215 (N_1215,N_980,N_841);
nand U1216 (N_1216,N_958,N_548);
or U1217 (N_1217,N_650,N_600);
or U1218 (N_1218,N_699,N_800);
nor U1219 (N_1219,N_838,N_690);
and U1220 (N_1220,N_692,N_790);
or U1221 (N_1221,N_503,N_646);
and U1222 (N_1222,N_536,N_956);
nor U1223 (N_1223,N_994,N_774);
nand U1224 (N_1224,N_676,N_847);
and U1225 (N_1225,N_824,N_834);
nand U1226 (N_1226,N_635,N_717);
nand U1227 (N_1227,N_928,N_514);
nand U1228 (N_1228,N_666,N_670);
and U1229 (N_1229,N_857,N_675);
nor U1230 (N_1230,N_683,N_821);
nand U1231 (N_1231,N_908,N_628);
or U1232 (N_1232,N_964,N_701);
or U1233 (N_1233,N_661,N_886);
nand U1234 (N_1234,N_924,N_689);
or U1235 (N_1235,N_695,N_516);
or U1236 (N_1236,N_700,N_672);
and U1237 (N_1237,N_917,N_530);
and U1238 (N_1238,N_793,N_677);
or U1239 (N_1239,N_852,N_539);
nand U1240 (N_1240,N_810,N_769);
and U1241 (N_1241,N_561,N_694);
nor U1242 (N_1242,N_587,N_520);
nor U1243 (N_1243,N_984,N_894);
and U1244 (N_1244,N_926,N_747);
and U1245 (N_1245,N_636,N_811);
or U1246 (N_1246,N_529,N_594);
or U1247 (N_1247,N_504,N_621);
and U1248 (N_1248,N_965,N_622);
nand U1249 (N_1249,N_996,N_738);
nor U1250 (N_1250,N_998,N_548);
nor U1251 (N_1251,N_710,N_782);
nor U1252 (N_1252,N_831,N_939);
nor U1253 (N_1253,N_905,N_919);
or U1254 (N_1254,N_679,N_743);
nor U1255 (N_1255,N_808,N_562);
and U1256 (N_1256,N_508,N_715);
or U1257 (N_1257,N_657,N_551);
nand U1258 (N_1258,N_826,N_903);
or U1259 (N_1259,N_782,N_961);
and U1260 (N_1260,N_591,N_553);
nand U1261 (N_1261,N_594,N_551);
nand U1262 (N_1262,N_757,N_531);
or U1263 (N_1263,N_516,N_739);
xnor U1264 (N_1264,N_741,N_763);
and U1265 (N_1265,N_579,N_852);
or U1266 (N_1266,N_623,N_630);
and U1267 (N_1267,N_966,N_722);
nor U1268 (N_1268,N_791,N_693);
nand U1269 (N_1269,N_732,N_901);
nand U1270 (N_1270,N_943,N_708);
and U1271 (N_1271,N_641,N_919);
nor U1272 (N_1272,N_942,N_697);
nand U1273 (N_1273,N_542,N_894);
or U1274 (N_1274,N_690,N_627);
and U1275 (N_1275,N_570,N_850);
xor U1276 (N_1276,N_958,N_979);
or U1277 (N_1277,N_729,N_851);
and U1278 (N_1278,N_716,N_805);
or U1279 (N_1279,N_605,N_733);
or U1280 (N_1280,N_582,N_713);
and U1281 (N_1281,N_812,N_950);
nand U1282 (N_1282,N_980,N_581);
nor U1283 (N_1283,N_752,N_863);
and U1284 (N_1284,N_770,N_772);
nor U1285 (N_1285,N_836,N_999);
and U1286 (N_1286,N_565,N_780);
xor U1287 (N_1287,N_761,N_551);
or U1288 (N_1288,N_619,N_610);
or U1289 (N_1289,N_852,N_966);
nand U1290 (N_1290,N_598,N_687);
and U1291 (N_1291,N_565,N_555);
and U1292 (N_1292,N_583,N_893);
nand U1293 (N_1293,N_916,N_913);
and U1294 (N_1294,N_751,N_567);
and U1295 (N_1295,N_906,N_666);
nand U1296 (N_1296,N_709,N_654);
nor U1297 (N_1297,N_724,N_575);
nor U1298 (N_1298,N_860,N_670);
or U1299 (N_1299,N_882,N_781);
and U1300 (N_1300,N_632,N_874);
and U1301 (N_1301,N_665,N_539);
and U1302 (N_1302,N_655,N_502);
or U1303 (N_1303,N_604,N_613);
nor U1304 (N_1304,N_885,N_687);
nor U1305 (N_1305,N_818,N_585);
or U1306 (N_1306,N_615,N_965);
nand U1307 (N_1307,N_515,N_811);
and U1308 (N_1308,N_969,N_836);
and U1309 (N_1309,N_781,N_777);
or U1310 (N_1310,N_516,N_663);
nand U1311 (N_1311,N_775,N_539);
nand U1312 (N_1312,N_595,N_880);
nor U1313 (N_1313,N_824,N_930);
nor U1314 (N_1314,N_854,N_546);
or U1315 (N_1315,N_814,N_882);
nand U1316 (N_1316,N_503,N_938);
and U1317 (N_1317,N_680,N_805);
nor U1318 (N_1318,N_612,N_932);
nand U1319 (N_1319,N_822,N_790);
nor U1320 (N_1320,N_679,N_627);
nor U1321 (N_1321,N_533,N_840);
nor U1322 (N_1322,N_521,N_933);
nor U1323 (N_1323,N_827,N_592);
or U1324 (N_1324,N_740,N_691);
nand U1325 (N_1325,N_776,N_730);
nor U1326 (N_1326,N_689,N_603);
and U1327 (N_1327,N_967,N_625);
and U1328 (N_1328,N_566,N_895);
nand U1329 (N_1329,N_589,N_888);
or U1330 (N_1330,N_878,N_777);
nor U1331 (N_1331,N_513,N_566);
nor U1332 (N_1332,N_586,N_659);
nor U1333 (N_1333,N_785,N_967);
or U1334 (N_1334,N_849,N_732);
or U1335 (N_1335,N_856,N_796);
nor U1336 (N_1336,N_923,N_743);
nor U1337 (N_1337,N_863,N_762);
or U1338 (N_1338,N_614,N_735);
or U1339 (N_1339,N_978,N_546);
or U1340 (N_1340,N_720,N_821);
nand U1341 (N_1341,N_529,N_968);
and U1342 (N_1342,N_625,N_859);
and U1343 (N_1343,N_795,N_749);
and U1344 (N_1344,N_821,N_916);
or U1345 (N_1345,N_619,N_843);
and U1346 (N_1346,N_886,N_807);
nand U1347 (N_1347,N_646,N_580);
and U1348 (N_1348,N_827,N_514);
and U1349 (N_1349,N_704,N_849);
nor U1350 (N_1350,N_579,N_819);
and U1351 (N_1351,N_639,N_702);
and U1352 (N_1352,N_631,N_859);
or U1353 (N_1353,N_624,N_977);
nor U1354 (N_1354,N_636,N_711);
nand U1355 (N_1355,N_857,N_866);
nand U1356 (N_1356,N_877,N_507);
nor U1357 (N_1357,N_736,N_731);
and U1358 (N_1358,N_658,N_745);
nor U1359 (N_1359,N_746,N_842);
nor U1360 (N_1360,N_939,N_830);
or U1361 (N_1361,N_950,N_556);
or U1362 (N_1362,N_641,N_950);
or U1363 (N_1363,N_777,N_948);
nand U1364 (N_1364,N_769,N_871);
nor U1365 (N_1365,N_910,N_946);
or U1366 (N_1366,N_688,N_756);
and U1367 (N_1367,N_761,N_784);
nand U1368 (N_1368,N_759,N_864);
xor U1369 (N_1369,N_610,N_849);
or U1370 (N_1370,N_656,N_502);
or U1371 (N_1371,N_829,N_532);
and U1372 (N_1372,N_743,N_719);
nand U1373 (N_1373,N_764,N_991);
or U1374 (N_1374,N_602,N_822);
nand U1375 (N_1375,N_778,N_745);
nor U1376 (N_1376,N_862,N_508);
or U1377 (N_1377,N_881,N_514);
nand U1378 (N_1378,N_663,N_610);
nand U1379 (N_1379,N_909,N_503);
and U1380 (N_1380,N_720,N_816);
or U1381 (N_1381,N_914,N_807);
and U1382 (N_1382,N_632,N_977);
nor U1383 (N_1383,N_540,N_742);
or U1384 (N_1384,N_892,N_501);
nand U1385 (N_1385,N_870,N_959);
or U1386 (N_1386,N_510,N_741);
or U1387 (N_1387,N_764,N_707);
nor U1388 (N_1388,N_798,N_998);
nor U1389 (N_1389,N_696,N_954);
nor U1390 (N_1390,N_900,N_787);
and U1391 (N_1391,N_553,N_592);
and U1392 (N_1392,N_939,N_760);
and U1393 (N_1393,N_830,N_940);
nand U1394 (N_1394,N_513,N_674);
and U1395 (N_1395,N_950,N_768);
or U1396 (N_1396,N_691,N_818);
nand U1397 (N_1397,N_582,N_985);
nor U1398 (N_1398,N_709,N_728);
or U1399 (N_1399,N_834,N_637);
nor U1400 (N_1400,N_504,N_850);
xnor U1401 (N_1401,N_885,N_963);
or U1402 (N_1402,N_966,N_738);
nand U1403 (N_1403,N_610,N_701);
nor U1404 (N_1404,N_688,N_528);
nor U1405 (N_1405,N_871,N_970);
or U1406 (N_1406,N_830,N_829);
nand U1407 (N_1407,N_972,N_737);
or U1408 (N_1408,N_998,N_696);
and U1409 (N_1409,N_912,N_694);
or U1410 (N_1410,N_717,N_841);
nor U1411 (N_1411,N_894,N_522);
nand U1412 (N_1412,N_546,N_612);
nor U1413 (N_1413,N_694,N_678);
and U1414 (N_1414,N_917,N_978);
nand U1415 (N_1415,N_747,N_959);
and U1416 (N_1416,N_692,N_711);
nor U1417 (N_1417,N_502,N_930);
nand U1418 (N_1418,N_986,N_525);
nand U1419 (N_1419,N_838,N_592);
nand U1420 (N_1420,N_546,N_668);
nand U1421 (N_1421,N_911,N_852);
nand U1422 (N_1422,N_501,N_822);
or U1423 (N_1423,N_518,N_818);
or U1424 (N_1424,N_596,N_630);
or U1425 (N_1425,N_823,N_850);
nand U1426 (N_1426,N_755,N_778);
nand U1427 (N_1427,N_626,N_527);
and U1428 (N_1428,N_731,N_868);
nor U1429 (N_1429,N_677,N_956);
or U1430 (N_1430,N_998,N_675);
nor U1431 (N_1431,N_917,N_886);
or U1432 (N_1432,N_705,N_583);
nor U1433 (N_1433,N_838,N_824);
and U1434 (N_1434,N_888,N_837);
nand U1435 (N_1435,N_619,N_800);
nor U1436 (N_1436,N_581,N_774);
nor U1437 (N_1437,N_645,N_936);
nor U1438 (N_1438,N_763,N_978);
or U1439 (N_1439,N_882,N_502);
and U1440 (N_1440,N_964,N_793);
nand U1441 (N_1441,N_980,N_700);
nand U1442 (N_1442,N_570,N_938);
nand U1443 (N_1443,N_564,N_682);
or U1444 (N_1444,N_530,N_861);
nor U1445 (N_1445,N_833,N_923);
or U1446 (N_1446,N_732,N_916);
nor U1447 (N_1447,N_902,N_688);
or U1448 (N_1448,N_816,N_694);
or U1449 (N_1449,N_798,N_973);
or U1450 (N_1450,N_951,N_569);
or U1451 (N_1451,N_580,N_816);
and U1452 (N_1452,N_534,N_551);
and U1453 (N_1453,N_659,N_517);
nand U1454 (N_1454,N_947,N_682);
or U1455 (N_1455,N_595,N_584);
nand U1456 (N_1456,N_997,N_677);
or U1457 (N_1457,N_604,N_843);
or U1458 (N_1458,N_746,N_598);
nand U1459 (N_1459,N_635,N_832);
or U1460 (N_1460,N_880,N_518);
and U1461 (N_1461,N_753,N_936);
or U1462 (N_1462,N_640,N_892);
or U1463 (N_1463,N_805,N_765);
or U1464 (N_1464,N_519,N_693);
and U1465 (N_1465,N_890,N_678);
or U1466 (N_1466,N_791,N_961);
and U1467 (N_1467,N_501,N_835);
nand U1468 (N_1468,N_963,N_862);
and U1469 (N_1469,N_927,N_721);
nor U1470 (N_1470,N_915,N_631);
and U1471 (N_1471,N_870,N_532);
nand U1472 (N_1472,N_548,N_735);
nand U1473 (N_1473,N_825,N_631);
and U1474 (N_1474,N_688,N_727);
nor U1475 (N_1475,N_996,N_532);
nor U1476 (N_1476,N_550,N_876);
nor U1477 (N_1477,N_898,N_546);
or U1478 (N_1478,N_922,N_720);
or U1479 (N_1479,N_586,N_826);
xor U1480 (N_1480,N_743,N_740);
or U1481 (N_1481,N_627,N_947);
or U1482 (N_1482,N_536,N_757);
or U1483 (N_1483,N_664,N_680);
nand U1484 (N_1484,N_893,N_890);
nor U1485 (N_1485,N_581,N_665);
or U1486 (N_1486,N_627,N_845);
or U1487 (N_1487,N_567,N_647);
or U1488 (N_1488,N_871,N_727);
nor U1489 (N_1489,N_663,N_981);
nand U1490 (N_1490,N_877,N_881);
nor U1491 (N_1491,N_936,N_767);
nor U1492 (N_1492,N_557,N_563);
nand U1493 (N_1493,N_780,N_805);
nand U1494 (N_1494,N_845,N_765);
nor U1495 (N_1495,N_861,N_949);
and U1496 (N_1496,N_501,N_790);
nand U1497 (N_1497,N_773,N_935);
and U1498 (N_1498,N_778,N_741);
and U1499 (N_1499,N_815,N_564);
nor U1500 (N_1500,N_1255,N_1224);
or U1501 (N_1501,N_1284,N_1377);
nand U1502 (N_1502,N_1287,N_1374);
nor U1503 (N_1503,N_1273,N_1106);
nand U1504 (N_1504,N_1188,N_1469);
nand U1505 (N_1505,N_1295,N_1068);
nor U1506 (N_1506,N_1193,N_1135);
nor U1507 (N_1507,N_1153,N_1014);
and U1508 (N_1508,N_1015,N_1343);
and U1509 (N_1509,N_1242,N_1052);
nor U1510 (N_1510,N_1365,N_1380);
and U1511 (N_1511,N_1372,N_1436);
nor U1512 (N_1512,N_1311,N_1084);
nand U1513 (N_1513,N_1168,N_1375);
nor U1514 (N_1514,N_1041,N_1249);
nand U1515 (N_1515,N_1075,N_1254);
nor U1516 (N_1516,N_1386,N_1216);
and U1517 (N_1517,N_1376,N_1165);
or U1518 (N_1518,N_1102,N_1160);
and U1519 (N_1519,N_1349,N_1332);
and U1520 (N_1520,N_1393,N_1400);
and U1521 (N_1521,N_1241,N_1336);
and U1522 (N_1522,N_1435,N_1370);
nor U1523 (N_1523,N_1159,N_1077);
and U1524 (N_1524,N_1317,N_1211);
nand U1525 (N_1525,N_1210,N_1272);
or U1526 (N_1526,N_1341,N_1267);
nand U1527 (N_1527,N_1225,N_1302);
nor U1528 (N_1528,N_1209,N_1117);
or U1529 (N_1529,N_1268,N_1474);
or U1530 (N_1530,N_1213,N_1038);
nor U1531 (N_1531,N_1059,N_1490);
or U1532 (N_1532,N_1244,N_1115);
and U1533 (N_1533,N_1230,N_1166);
and U1534 (N_1534,N_1199,N_1324);
nor U1535 (N_1535,N_1437,N_1013);
nor U1536 (N_1536,N_1422,N_1124);
nor U1537 (N_1537,N_1489,N_1017);
nor U1538 (N_1538,N_1382,N_1360);
nand U1539 (N_1539,N_1089,N_1095);
nand U1540 (N_1540,N_1090,N_1478);
or U1541 (N_1541,N_1133,N_1246);
nor U1542 (N_1542,N_1368,N_1183);
and U1543 (N_1543,N_1439,N_1288);
nand U1544 (N_1544,N_1196,N_1062);
nand U1545 (N_1545,N_1050,N_1040);
and U1546 (N_1546,N_1446,N_1137);
and U1547 (N_1547,N_1410,N_1261);
nor U1548 (N_1548,N_1345,N_1082);
or U1549 (N_1549,N_1163,N_1329);
or U1550 (N_1550,N_1339,N_1367);
nand U1551 (N_1551,N_1328,N_1071);
nand U1552 (N_1552,N_1308,N_1304);
or U1553 (N_1553,N_1202,N_1477);
and U1554 (N_1554,N_1141,N_1310);
and U1555 (N_1555,N_1229,N_1378);
nand U1556 (N_1556,N_1011,N_1479);
and U1557 (N_1557,N_1259,N_1399);
or U1558 (N_1558,N_1187,N_1155);
nor U1559 (N_1559,N_1274,N_1081);
or U1560 (N_1560,N_1282,N_1006);
nor U1561 (N_1561,N_1042,N_1428);
and U1562 (N_1562,N_1420,N_1495);
or U1563 (N_1563,N_1045,N_1313);
or U1564 (N_1564,N_1114,N_1108);
and U1565 (N_1565,N_1214,N_1444);
or U1566 (N_1566,N_1096,N_1481);
nor U1567 (N_1567,N_1233,N_1236);
and U1568 (N_1568,N_1491,N_1001);
nor U1569 (N_1569,N_1192,N_1238);
or U1570 (N_1570,N_1113,N_1174);
and U1571 (N_1571,N_1130,N_1316);
and U1572 (N_1572,N_1167,N_1072);
or U1573 (N_1573,N_1322,N_1407);
and U1574 (N_1574,N_1004,N_1172);
nor U1575 (N_1575,N_1227,N_1154);
or U1576 (N_1576,N_1381,N_1087);
and U1577 (N_1577,N_1487,N_1335);
nand U1578 (N_1578,N_1197,N_1066);
nor U1579 (N_1579,N_1025,N_1306);
nor U1580 (N_1580,N_1093,N_1118);
and U1581 (N_1581,N_1440,N_1352);
or U1582 (N_1582,N_1007,N_1148);
or U1583 (N_1583,N_1391,N_1046);
nand U1584 (N_1584,N_1403,N_1411);
or U1585 (N_1585,N_1499,N_1270);
xor U1586 (N_1586,N_1262,N_1021);
nand U1587 (N_1587,N_1049,N_1362);
nor U1588 (N_1588,N_1026,N_1150);
nand U1589 (N_1589,N_1398,N_1286);
or U1590 (N_1590,N_1454,N_1088);
and U1591 (N_1591,N_1323,N_1098);
nor U1592 (N_1592,N_1024,N_1239);
or U1593 (N_1593,N_1047,N_1488);
nor U1594 (N_1594,N_1320,N_1285);
or U1595 (N_1595,N_1147,N_1484);
or U1596 (N_1596,N_1494,N_1279);
or U1597 (N_1597,N_1109,N_1458);
and U1598 (N_1598,N_1461,N_1441);
nor U1599 (N_1599,N_1460,N_1340);
and U1600 (N_1600,N_1053,N_1426);
or U1601 (N_1601,N_1182,N_1373);
or U1602 (N_1602,N_1292,N_1347);
and U1603 (N_1603,N_1146,N_1390);
or U1604 (N_1604,N_1305,N_1003);
nand U1605 (N_1605,N_1486,N_1111);
and U1606 (N_1606,N_1010,N_1116);
or U1607 (N_1607,N_1100,N_1122);
or U1608 (N_1608,N_1212,N_1475);
nor U1609 (N_1609,N_1140,N_1097);
or U1610 (N_1610,N_1278,N_1438);
nor U1611 (N_1611,N_1421,N_1019);
and U1612 (N_1612,N_1034,N_1151);
nand U1613 (N_1613,N_1152,N_1351);
or U1614 (N_1614,N_1215,N_1307);
and U1615 (N_1615,N_1303,N_1016);
or U1616 (N_1616,N_1466,N_1432);
or U1617 (N_1617,N_1318,N_1472);
or U1618 (N_1618,N_1492,N_1326);
nand U1619 (N_1619,N_1157,N_1482);
or U1620 (N_1620,N_1131,N_1094);
and U1621 (N_1621,N_1371,N_1260);
and U1622 (N_1622,N_1190,N_1346);
and U1623 (N_1623,N_1344,N_1033);
and U1624 (N_1624,N_1110,N_1257);
and U1625 (N_1625,N_1423,N_1069);
or U1626 (N_1626,N_1051,N_1379);
nand U1627 (N_1627,N_1175,N_1226);
nand U1628 (N_1628,N_1496,N_1277);
or U1629 (N_1629,N_1291,N_1470);
and U1630 (N_1630,N_1433,N_1392);
nor U1631 (N_1631,N_1498,N_1309);
and U1632 (N_1632,N_1086,N_1235);
or U1633 (N_1633,N_1383,N_1067);
nor U1634 (N_1634,N_1080,N_1385);
and U1635 (N_1635,N_1493,N_1315);
nand U1636 (N_1636,N_1266,N_1121);
or U1637 (N_1637,N_1330,N_1389);
and U1638 (N_1638,N_1120,N_1397);
nor U1639 (N_1639,N_1416,N_1206);
and U1640 (N_1640,N_1388,N_1497);
and U1641 (N_1641,N_1463,N_1350);
and U1642 (N_1642,N_1301,N_1105);
nor U1643 (N_1643,N_1417,N_1099);
nor U1644 (N_1644,N_1280,N_1162);
or U1645 (N_1645,N_1186,N_1468);
xor U1646 (N_1646,N_1419,N_1180);
or U1647 (N_1647,N_1178,N_1065);
nor U1648 (N_1648,N_1465,N_1312);
or U1649 (N_1649,N_1445,N_1325);
nand U1650 (N_1650,N_1144,N_1048);
and U1651 (N_1651,N_1177,N_1237);
or U1652 (N_1652,N_1198,N_1402);
or U1653 (N_1653,N_1338,N_1476);
xor U1654 (N_1654,N_1200,N_1447);
nand U1655 (N_1655,N_1023,N_1408);
nor U1656 (N_1656,N_1248,N_1195);
nand U1657 (N_1657,N_1185,N_1353);
nand U1658 (N_1658,N_1161,N_1064);
and U1659 (N_1659,N_1451,N_1387);
nand U1660 (N_1660,N_1107,N_1358);
nor U1661 (N_1661,N_1364,N_1404);
or U1662 (N_1662,N_1143,N_1028);
or U1663 (N_1663,N_1058,N_1314);
nand U1664 (N_1664,N_1369,N_1223);
nand U1665 (N_1665,N_1258,N_1030);
and U1666 (N_1666,N_1092,N_1263);
or U1667 (N_1667,N_1355,N_1061);
or U1668 (N_1668,N_1427,N_1164);
nor U1669 (N_1669,N_1036,N_1022);
nand U1670 (N_1670,N_1189,N_1057);
nand U1671 (N_1671,N_1290,N_1128);
nand U1672 (N_1672,N_1129,N_1348);
nand U1673 (N_1673,N_1060,N_1289);
or U1674 (N_1674,N_1243,N_1055);
nor U1675 (N_1675,N_1431,N_1138);
or U1676 (N_1676,N_1173,N_1449);
nand U1677 (N_1677,N_1293,N_1405);
or U1678 (N_1678,N_1222,N_1276);
and U1679 (N_1679,N_1296,N_1018);
or U1680 (N_1680,N_1139,N_1044);
and U1681 (N_1681,N_1253,N_1076);
or U1682 (N_1682,N_1181,N_1204);
nand U1683 (N_1683,N_1363,N_1169);
or U1684 (N_1684,N_1356,N_1418);
or U1685 (N_1685,N_1250,N_1337);
or U1686 (N_1686,N_1158,N_1299);
or U1687 (N_1687,N_1119,N_1415);
and U1688 (N_1688,N_1112,N_1251);
nand U1689 (N_1689,N_1170,N_1231);
and U1690 (N_1690,N_1283,N_1078);
and U1691 (N_1691,N_1430,N_1009);
or U1692 (N_1692,N_1264,N_1459);
and U1693 (N_1693,N_1271,N_1194);
nor U1694 (N_1694,N_1256,N_1035);
or U1695 (N_1695,N_1275,N_1083);
nor U1696 (N_1696,N_1039,N_1450);
xnor U1697 (N_1697,N_1027,N_1101);
nand U1698 (N_1698,N_1218,N_1240);
or U1699 (N_1699,N_1091,N_1395);
nor U1700 (N_1700,N_1245,N_1073);
or U1701 (N_1701,N_1205,N_1191);
or U1702 (N_1702,N_1471,N_1104);
nor U1703 (N_1703,N_1462,N_1145);
and U1704 (N_1704,N_1480,N_1396);
or U1705 (N_1705,N_1000,N_1043);
nand U1706 (N_1706,N_1125,N_1134);
and U1707 (N_1707,N_1149,N_1414);
and U1708 (N_1708,N_1228,N_1232);
or U1709 (N_1709,N_1448,N_1333);
or U1710 (N_1710,N_1220,N_1269);
or U1711 (N_1711,N_1409,N_1054);
or U1712 (N_1712,N_1334,N_1176);
or U1713 (N_1713,N_1142,N_1354);
and U1714 (N_1714,N_1300,N_1203);
nand U1715 (N_1715,N_1031,N_1074);
nand U1716 (N_1716,N_1452,N_1455);
nand U1717 (N_1717,N_1359,N_1171);
nor U1718 (N_1718,N_1126,N_1361);
nor U1719 (N_1719,N_1221,N_1056);
nand U1720 (N_1720,N_1457,N_1037);
nand U1721 (N_1721,N_1029,N_1252);
nor U1722 (N_1722,N_1384,N_1485);
nand U1723 (N_1723,N_1008,N_1467);
xnor U1724 (N_1724,N_1413,N_1085);
nor U1725 (N_1725,N_1429,N_1297);
nand U1726 (N_1726,N_1394,N_1219);
nor U1727 (N_1727,N_1366,N_1201);
or U1728 (N_1728,N_1217,N_1434);
and U1729 (N_1729,N_1103,N_1342);
nand U1730 (N_1730,N_1247,N_1184);
nor U1731 (N_1731,N_1005,N_1207);
or U1732 (N_1732,N_1424,N_1132);
nor U1733 (N_1733,N_1464,N_1294);
or U1734 (N_1734,N_1357,N_1063);
and U1735 (N_1735,N_1453,N_1473);
or U1736 (N_1736,N_1406,N_1208);
and U1737 (N_1737,N_1234,N_1331);
or U1738 (N_1738,N_1442,N_1265);
nand U1739 (N_1739,N_1327,N_1136);
nand U1740 (N_1740,N_1156,N_1456);
nand U1741 (N_1741,N_1443,N_1070);
or U1742 (N_1742,N_1401,N_1127);
and U1743 (N_1743,N_1298,N_1321);
or U1744 (N_1744,N_1319,N_1412);
or U1745 (N_1745,N_1483,N_1179);
nand U1746 (N_1746,N_1079,N_1123);
and U1747 (N_1747,N_1020,N_1281);
and U1748 (N_1748,N_1032,N_1012);
nor U1749 (N_1749,N_1425,N_1002);
nor U1750 (N_1750,N_1196,N_1031);
nand U1751 (N_1751,N_1096,N_1235);
nor U1752 (N_1752,N_1464,N_1378);
or U1753 (N_1753,N_1463,N_1335);
nand U1754 (N_1754,N_1055,N_1189);
and U1755 (N_1755,N_1369,N_1175);
and U1756 (N_1756,N_1245,N_1438);
nand U1757 (N_1757,N_1137,N_1284);
nor U1758 (N_1758,N_1105,N_1414);
nand U1759 (N_1759,N_1484,N_1474);
nor U1760 (N_1760,N_1356,N_1100);
or U1761 (N_1761,N_1090,N_1034);
nand U1762 (N_1762,N_1092,N_1066);
or U1763 (N_1763,N_1396,N_1308);
nand U1764 (N_1764,N_1264,N_1187);
or U1765 (N_1765,N_1297,N_1338);
xor U1766 (N_1766,N_1001,N_1414);
and U1767 (N_1767,N_1289,N_1019);
nor U1768 (N_1768,N_1216,N_1086);
nand U1769 (N_1769,N_1101,N_1395);
and U1770 (N_1770,N_1199,N_1492);
and U1771 (N_1771,N_1333,N_1057);
nor U1772 (N_1772,N_1024,N_1232);
nand U1773 (N_1773,N_1094,N_1231);
nand U1774 (N_1774,N_1041,N_1094);
nand U1775 (N_1775,N_1335,N_1377);
nand U1776 (N_1776,N_1217,N_1334);
nand U1777 (N_1777,N_1262,N_1165);
or U1778 (N_1778,N_1043,N_1287);
and U1779 (N_1779,N_1120,N_1496);
nor U1780 (N_1780,N_1035,N_1308);
nand U1781 (N_1781,N_1006,N_1050);
nand U1782 (N_1782,N_1458,N_1043);
nor U1783 (N_1783,N_1283,N_1433);
nor U1784 (N_1784,N_1116,N_1190);
nor U1785 (N_1785,N_1027,N_1177);
nor U1786 (N_1786,N_1159,N_1466);
and U1787 (N_1787,N_1256,N_1193);
nand U1788 (N_1788,N_1222,N_1075);
nand U1789 (N_1789,N_1406,N_1006);
and U1790 (N_1790,N_1184,N_1317);
nor U1791 (N_1791,N_1276,N_1271);
nor U1792 (N_1792,N_1007,N_1279);
nor U1793 (N_1793,N_1141,N_1484);
or U1794 (N_1794,N_1217,N_1416);
or U1795 (N_1795,N_1217,N_1108);
or U1796 (N_1796,N_1461,N_1294);
nand U1797 (N_1797,N_1393,N_1249);
nor U1798 (N_1798,N_1449,N_1122);
or U1799 (N_1799,N_1034,N_1075);
or U1800 (N_1800,N_1234,N_1347);
nand U1801 (N_1801,N_1135,N_1014);
nand U1802 (N_1802,N_1369,N_1108);
or U1803 (N_1803,N_1495,N_1406);
or U1804 (N_1804,N_1401,N_1476);
and U1805 (N_1805,N_1424,N_1400);
nor U1806 (N_1806,N_1050,N_1312);
and U1807 (N_1807,N_1023,N_1493);
xnor U1808 (N_1808,N_1165,N_1496);
or U1809 (N_1809,N_1312,N_1371);
or U1810 (N_1810,N_1478,N_1425);
or U1811 (N_1811,N_1263,N_1003);
nor U1812 (N_1812,N_1422,N_1226);
nand U1813 (N_1813,N_1256,N_1391);
or U1814 (N_1814,N_1109,N_1371);
nor U1815 (N_1815,N_1178,N_1346);
nor U1816 (N_1816,N_1470,N_1390);
nor U1817 (N_1817,N_1260,N_1277);
or U1818 (N_1818,N_1243,N_1061);
nor U1819 (N_1819,N_1290,N_1151);
or U1820 (N_1820,N_1272,N_1189);
or U1821 (N_1821,N_1012,N_1454);
and U1822 (N_1822,N_1394,N_1476);
nand U1823 (N_1823,N_1132,N_1494);
or U1824 (N_1824,N_1484,N_1019);
or U1825 (N_1825,N_1476,N_1048);
or U1826 (N_1826,N_1321,N_1494);
and U1827 (N_1827,N_1324,N_1063);
and U1828 (N_1828,N_1252,N_1309);
and U1829 (N_1829,N_1091,N_1255);
nor U1830 (N_1830,N_1218,N_1236);
or U1831 (N_1831,N_1382,N_1312);
nor U1832 (N_1832,N_1099,N_1143);
and U1833 (N_1833,N_1293,N_1072);
nor U1834 (N_1834,N_1209,N_1069);
xnor U1835 (N_1835,N_1285,N_1476);
and U1836 (N_1836,N_1262,N_1195);
or U1837 (N_1837,N_1463,N_1457);
nand U1838 (N_1838,N_1279,N_1120);
and U1839 (N_1839,N_1010,N_1419);
nor U1840 (N_1840,N_1498,N_1169);
nor U1841 (N_1841,N_1183,N_1424);
nor U1842 (N_1842,N_1136,N_1474);
nand U1843 (N_1843,N_1107,N_1051);
or U1844 (N_1844,N_1117,N_1379);
or U1845 (N_1845,N_1411,N_1123);
and U1846 (N_1846,N_1137,N_1007);
or U1847 (N_1847,N_1451,N_1012);
nand U1848 (N_1848,N_1012,N_1148);
nand U1849 (N_1849,N_1347,N_1293);
nand U1850 (N_1850,N_1395,N_1043);
or U1851 (N_1851,N_1106,N_1360);
nor U1852 (N_1852,N_1408,N_1435);
nor U1853 (N_1853,N_1323,N_1327);
xnor U1854 (N_1854,N_1294,N_1312);
nand U1855 (N_1855,N_1214,N_1139);
nand U1856 (N_1856,N_1323,N_1029);
nand U1857 (N_1857,N_1132,N_1229);
nor U1858 (N_1858,N_1398,N_1275);
and U1859 (N_1859,N_1275,N_1042);
or U1860 (N_1860,N_1374,N_1038);
or U1861 (N_1861,N_1182,N_1170);
nor U1862 (N_1862,N_1035,N_1407);
nand U1863 (N_1863,N_1347,N_1459);
and U1864 (N_1864,N_1144,N_1435);
nand U1865 (N_1865,N_1465,N_1212);
and U1866 (N_1866,N_1055,N_1120);
and U1867 (N_1867,N_1001,N_1224);
nand U1868 (N_1868,N_1183,N_1406);
or U1869 (N_1869,N_1306,N_1411);
or U1870 (N_1870,N_1002,N_1107);
and U1871 (N_1871,N_1350,N_1313);
or U1872 (N_1872,N_1059,N_1425);
and U1873 (N_1873,N_1408,N_1442);
nand U1874 (N_1874,N_1285,N_1271);
nand U1875 (N_1875,N_1427,N_1333);
nor U1876 (N_1876,N_1409,N_1343);
nor U1877 (N_1877,N_1162,N_1062);
nand U1878 (N_1878,N_1245,N_1087);
nand U1879 (N_1879,N_1474,N_1038);
or U1880 (N_1880,N_1203,N_1378);
nand U1881 (N_1881,N_1290,N_1392);
and U1882 (N_1882,N_1243,N_1266);
nand U1883 (N_1883,N_1138,N_1452);
nand U1884 (N_1884,N_1478,N_1318);
nand U1885 (N_1885,N_1256,N_1374);
nor U1886 (N_1886,N_1172,N_1269);
or U1887 (N_1887,N_1380,N_1219);
and U1888 (N_1888,N_1216,N_1384);
nand U1889 (N_1889,N_1440,N_1318);
or U1890 (N_1890,N_1190,N_1252);
and U1891 (N_1891,N_1335,N_1133);
or U1892 (N_1892,N_1045,N_1439);
nand U1893 (N_1893,N_1420,N_1398);
and U1894 (N_1894,N_1481,N_1071);
nor U1895 (N_1895,N_1080,N_1375);
nor U1896 (N_1896,N_1438,N_1218);
or U1897 (N_1897,N_1383,N_1320);
or U1898 (N_1898,N_1023,N_1196);
or U1899 (N_1899,N_1274,N_1253);
nor U1900 (N_1900,N_1035,N_1459);
nor U1901 (N_1901,N_1049,N_1353);
nand U1902 (N_1902,N_1391,N_1475);
nor U1903 (N_1903,N_1443,N_1366);
and U1904 (N_1904,N_1429,N_1462);
and U1905 (N_1905,N_1262,N_1337);
or U1906 (N_1906,N_1064,N_1270);
or U1907 (N_1907,N_1159,N_1422);
and U1908 (N_1908,N_1020,N_1200);
nor U1909 (N_1909,N_1031,N_1261);
nor U1910 (N_1910,N_1474,N_1173);
and U1911 (N_1911,N_1094,N_1487);
or U1912 (N_1912,N_1320,N_1420);
nand U1913 (N_1913,N_1223,N_1328);
nor U1914 (N_1914,N_1294,N_1497);
and U1915 (N_1915,N_1155,N_1053);
or U1916 (N_1916,N_1473,N_1489);
and U1917 (N_1917,N_1027,N_1342);
or U1918 (N_1918,N_1483,N_1434);
nor U1919 (N_1919,N_1121,N_1022);
nor U1920 (N_1920,N_1087,N_1324);
nor U1921 (N_1921,N_1168,N_1208);
and U1922 (N_1922,N_1250,N_1089);
or U1923 (N_1923,N_1226,N_1126);
and U1924 (N_1924,N_1450,N_1334);
or U1925 (N_1925,N_1271,N_1416);
nor U1926 (N_1926,N_1491,N_1328);
and U1927 (N_1927,N_1233,N_1446);
and U1928 (N_1928,N_1391,N_1487);
and U1929 (N_1929,N_1254,N_1200);
or U1930 (N_1930,N_1059,N_1075);
nand U1931 (N_1931,N_1279,N_1131);
nor U1932 (N_1932,N_1367,N_1402);
nor U1933 (N_1933,N_1422,N_1033);
nor U1934 (N_1934,N_1459,N_1186);
nor U1935 (N_1935,N_1306,N_1212);
nand U1936 (N_1936,N_1140,N_1494);
nor U1937 (N_1937,N_1220,N_1361);
and U1938 (N_1938,N_1382,N_1379);
nor U1939 (N_1939,N_1334,N_1278);
nor U1940 (N_1940,N_1262,N_1146);
and U1941 (N_1941,N_1272,N_1494);
or U1942 (N_1942,N_1060,N_1428);
nand U1943 (N_1943,N_1492,N_1491);
nor U1944 (N_1944,N_1466,N_1072);
or U1945 (N_1945,N_1420,N_1437);
and U1946 (N_1946,N_1344,N_1284);
nand U1947 (N_1947,N_1042,N_1036);
or U1948 (N_1948,N_1029,N_1166);
nand U1949 (N_1949,N_1252,N_1371);
and U1950 (N_1950,N_1414,N_1310);
nand U1951 (N_1951,N_1006,N_1418);
or U1952 (N_1952,N_1066,N_1154);
and U1953 (N_1953,N_1474,N_1374);
or U1954 (N_1954,N_1061,N_1053);
nand U1955 (N_1955,N_1094,N_1481);
or U1956 (N_1956,N_1205,N_1473);
or U1957 (N_1957,N_1089,N_1439);
or U1958 (N_1958,N_1424,N_1347);
nor U1959 (N_1959,N_1293,N_1244);
nor U1960 (N_1960,N_1402,N_1365);
or U1961 (N_1961,N_1205,N_1480);
or U1962 (N_1962,N_1416,N_1188);
and U1963 (N_1963,N_1295,N_1456);
or U1964 (N_1964,N_1342,N_1497);
and U1965 (N_1965,N_1284,N_1341);
and U1966 (N_1966,N_1260,N_1247);
nand U1967 (N_1967,N_1192,N_1039);
nor U1968 (N_1968,N_1171,N_1177);
or U1969 (N_1969,N_1207,N_1088);
nor U1970 (N_1970,N_1133,N_1177);
nor U1971 (N_1971,N_1307,N_1205);
nand U1972 (N_1972,N_1084,N_1288);
nand U1973 (N_1973,N_1211,N_1167);
and U1974 (N_1974,N_1121,N_1188);
nand U1975 (N_1975,N_1351,N_1376);
and U1976 (N_1976,N_1253,N_1309);
nand U1977 (N_1977,N_1291,N_1392);
or U1978 (N_1978,N_1200,N_1071);
nand U1979 (N_1979,N_1141,N_1313);
nand U1980 (N_1980,N_1339,N_1238);
nand U1981 (N_1981,N_1426,N_1185);
or U1982 (N_1982,N_1131,N_1107);
or U1983 (N_1983,N_1398,N_1468);
nor U1984 (N_1984,N_1284,N_1296);
and U1985 (N_1985,N_1304,N_1126);
or U1986 (N_1986,N_1273,N_1363);
or U1987 (N_1987,N_1204,N_1055);
nor U1988 (N_1988,N_1293,N_1420);
nand U1989 (N_1989,N_1314,N_1175);
nor U1990 (N_1990,N_1064,N_1469);
nand U1991 (N_1991,N_1199,N_1378);
and U1992 (N_1992,N_1394,N_1082);
and U1993 (N_1993,N_1346,N_1071);
nand U1994 (N_1994,N_1016,N_1341);
or U1995 (N_1995,N_1082,N_1014);
or U1996 (N_1996,N_1369,N_1435);
and U1997 (N_1997,N_1170,N_1480);
nor U1998 (N_1998,N_1197,N_1417);
or U1999 (N_1999,N_1454,N_1400);
and U2000 (N_2000,N_1878,N_1686);
nor U2001 (N_2001,N_1659,N_1892);
and U2002 (N_2002,N_1998,N_1724);
or U2003 (N_2003,N_1553,N_1531);
or U2004 (N_2004,N_1916,N_1954);
nand U2005 (N_2005,N_1559,N_1695);
nand U2006 (N_2006,N_1544,N_1680);
nor U2007 (N_2007,N_1898,N_1860);
or U2008 (N_2008,N_1574,N_1921);
nor U2009 (N_2009,N_1525,N_1834);
and U2010 (N_2010,N_1712,N_1554);
or U2011 (N_2011,N_1508,N_1633);
or U2012 (N_2012,N_1551,N_1550);
or U2013 (N_2013,N_1883,N_1764);
or U2014 (N_2014,N_1858,N_1759);
or U2015 (N_2015,N_1933,N_1762);
or U2016 (N_2016,N_1943,N_1993);
or U2017 (N_2017,N_1516,N_1884);
or U2018 (N_2018,N_1619,N_1994);
and U2019 (N_2019,N_1861,N_1895);
or U2020 (N_2020,N_1957,N_1698);
nand U2021 (N_2021,N_1997,N_1945);
nand U2022 (N_2022,N_1747,N_1709);
and U2023 (N_2023,N_1571,N_1576);
and U2024 (N_2024,N_1730,N_1922);
nor U2025 (N_2025,N_1879,N_1951);
nand U2026 (N_2026,N_1671,N_1914);
and U2027 (N_2027,N_1563,N_1928);
and U2028 (N_2028,N_1609,N_1811);
nand U2029 (N_2029,N_1944,N_1580);
and U2030 (N_2030,N_1751,N_1765);
nand U2031 (N_2031,N_1814,N_1542);
or U2032 (N_2032,N_1539,N_1979);
and U2033 (N_2033,N_1556,N_1649);
nor U2034 (N_2034,N_1932,N_1645);
nor U2035 (N_2035,N_1777,N_1564);
and U2036 (N_2036,N_1547,N_1502);
nand U2037 (N_2037,N_1742,N_1596);
or U2038 (N_2038,N_1591,N_1526);
or U2039 (N_2039,N_1833,N_1911);
nand U2040 (N_2040,N_1940,N_1830);
and U2041 (N_2041,N_1968,N_1784);
nand U2042 (N_2042,N_1674,N_1782);
nand U2043 (N_2043,N_1831,N_1687);
and U2044 (N_2044,N_1915,N_1842);
nor U2045 (N_2045,N_1637,N_1909);
and U2046 (N_2046,N_1902,N_1501);
or U2047 (N_2047,N_1618,N_1634);
nor U2048 (N_2048,N_1780,N_1942);
and U2049 (N_2049,N_1668,N_1702);
and U2050 (N_2050,N_1887,N_1991);
and U2051 (N_2051,N_1797,N_1621);
nand U2052 (N_2052,N_1681,N_1738);
nor U2053 (N_2053,N_1512,N_1820);
nor U2054 (N_2054,N_1983,N_1607);
and U2055 (N_2055,N_1611,N_1992);
and U2056 (N_2056,N_1632,N_1774);
and U2057 (N_2057,N_1602,N_1673);
nand U2058 (N_2058,N_1952,N_1927);
nand U2059 (N_2059,N_1567,N_1807);
nand U2060 (N_2060,N_1958,N_1701);
and U2061 (N_2061,N_1984,N_1785);
nor U2062 (N_2062,N_1877,N_1623);
and U2063 (N_2063,N_1740,N_1737);
nor U2064 (N_2064,N_1899,N_1826);
and U2065 (N_2065,N_1725,N_1566);
nand U2066 (N_2066,N_1857,N_1813);
nand U2067 (N_2067,N_1662,N_1949);
nand U2068 (N_2068,N_1758,N_1848);
nor U2069 (N_2069,N_1770,N_1518);
nand U2070 (N_2070,N_1707,N_1626);
and U2071 (N_2071,N_1799,N_1912);
nor U2072 (N_2072,N_1638,N_1635);
nor U2073 (N_2073,N_1560,N_1715);
or U2074 (N_2074,N_1608,N_1966);
nand U2075 (N_2075,N_1776,N_1655);
nor U2076 (N_2076,N_1903,N_1658);
xor U2077 (N_2077,N_1669,N_1908);
nand U2078 (N_2078,N_1772,N_1515);
nand U2079 (N_2079,N_1821,N_1804);
and U2080 (N_2080,N_1622,N_1852);
or U2081 (N_2081,N_1552,N_1523);
and U2082 (N_2082,N_1521,N_1736);
nand U2083 (N_2083,N_1555,N_1844);
and U2084 (N_2084,N_1627,N_1534);
nand U2085 (N_2085,N_1793,N_1855);
nand U2086 (N_2086,N_1536,N_1947);
or U2087 (N_2087,N_1885,N_1750);
and U2088 (N_2088,N_1636,N_1642);
nor U2089 (N_2089,N_1605,N_1876);
nand U2090 (N_2090,N_1988,N_1739);
xnor U2091 (N_2091,N_1973,N_1976);
and U2092 (N_2092,N_1809,N_1620);
nand U2093 (N_2093,N_1828,N_1822);
nand U2094 (N_2094,N_1504,N_1529);
and U2095 (N_2095,N_1846,N_1546);
and U2096 (N_2096,N_1693,N_1744);
nor U2097 (N_2097,N_1977,N_1528);
nor U2098 (N_2098,N_1881,N_1906);
or U2099 (N_2099,N_1520,N_1696);
or U2100 (N_2100,N_1705,N_1616);
or U2101 (N_2101,N_1829,N_1593);
nand U2102 (N_2102,N_1880,N_1741);
nand U2103 (N_2103,N_1630,N_1716);
or U2104 (N_2104,N_1972,N_1766);
nand U2105 (N_2105,N_1896,N_1549);
or U2106 (N_2106,N_1786,N_1548);
or U2107 (N_2107,N_1961,N_1955);
or U2108 (N_2108,N_1692,N_1723);
and U2109 (N_2109,N_1981,N_1919);
nor U2110 (N_2110,N_1708,N_1936);
or U2111 (N_2111,N_1850,N_1875);
or U2112 (N_2112,N_1893,N_1978);
nand U2113 (N_2113,N_1870,N_1953);
or U2114 (N_2114,N_1950,N_1853);
nand U2115 (N_2115,N_1868,N_1891);
and U2116 (N_2116,N_1652,N_1578);
or U2117 (N_2117,N_1982,N_1790);
and U2118 (N_2118,N_1889,N_1996);
and U2119 (N_2119,N_1507,N_1631);
nand U2120 (N_2120,N_1558,N_1963);
and U2121 (N_2121,N_1532,N_1610);
nor U2122 (N_2122,N_1513,N_1648);
and U2123 (N_2123,N_1806,N_1923);
nor U2124 (N_2124,N_1872,N_1859);
or U2125 (N_2125,N_1678,N_1812);
or U2126 (N_2126,N_1689,N_1823);
nor U2127 (N_2127,N_1753,N_1752);
nand U2128 (N_2128,N_1711,N_1644);
nor U2129 (N_2129,N_1871,N_1665);
nor U2130 (N_2130,N_1836,N_1519);
or U2131 (N_2131,N_1768,N_1841);
nand U2132 (N_2132,N_1557,N_1901);
nand U2133 (N_2133,N_1779,N_1545);
or U2134 (N_2134,N_1615,N_1714);
and U2135 (N_2135,N_1676,N_1946);
nand U2136 (N_2136,N_1628,N_1694);
nor U2137 (N_2137,N_1543,N_1967);
nor U2138 (N_2138,N_1613,N_1587);
or U2139 (N_2139,N_1767,N_1733);
and U2140 (N_2140,N_1755,N_1960);
and U2141 (N_2141,N_1843,N_1731);
and U2142 (N_2142,N_1690,N_1761);
or U2143 (N_2143,N_1783,N_1939);
nor U2144 (N_2144,N_1805,N_1987);
nand U2145 (N_2145,N_1594,N_1540);
and U2146 (N_2146,N_1827,N_1787);
or U2147 (N_2147,N_1964,N_1980);
nor U2148 (N_2148,N_1825,N_1541);
and U2149 (N_2149,N_1651,N_1684);
and U2150 (N_2150,N_1788,N_1538);
and U2151 (N_2151,N_1920,N_1910);
nand U2152 (N_2152,N_1710,N_1735);
or U2153 (N_2153,N_1660,N_1970);
or U2154 (N_2154,N_1754,N_1604);
nand U2155 (N_2155,N_1904,N_1929);
nor U2156 (N_2156,N_1930,N_1986);
or U2157 (N_2157,N_1838,N_1917);
nor U2158 (N_2158,N_1832,N_1606);
and U2159 (N_2159,N_1926,N_1990);
and U2160 (N_2160,N_1583,N_1663);
nor U2161 (N_2161,N_1794,N_1962);
and U2162 (N_2162,N_1713,N_1948);
nor U2163 (N_2163,N_1718,N_1503);
and U2164 (N_2164,N_1646,N_1688);
nor U2165 (N_2165,N_1845,N_1700);
nor U2166 (N_2166,N_1575,N_1819);
or U2167 (N_2167,N_1522,N_1565);
and U2168 (N_2168,N_1938,N_1802);
or U2169 (N_2169,N_1506,N_1975);
or U2170 (N_2170,N_1641,N_1913);
nor U2171 (N_2171,N_1756,N_1728);
and U2172 (N_2172,N_1847,N_1769);
nand U2173 (N_2173,N_1989,N_1569);
and U2174 (N_2174,N_1959,N_1937);
or U2175 (N_2175,N_1699,N_1882);
nor U2176 (N_2176,N_1771,N_1612);
nor U2177 (N_2177,N_1837,N_1601);
and U2178 (N_2178,N_1661,N_1629);
nand U2179 (N_2179,N_1685,N_1840);
nor U2180 (N_2180,N_1995,N_1999);
and U2181 (N_2181,N_1598,N_1818);
or U2182 (N_2182,N_1517,N_1816);
nor U2183 (N_2183,N_1726,N_1734);
nand U2184 (N_2184,N_1561,N_1934);
or U2185 (N_2185,N_1677,N_1568);
or U2186 (N_2186,N_1500,N_1749);
or U2187 (N_2187,N_1640,N_1869);
nand U2188 (N_2188,N_1624,N_1666);
nor U2189 (N_2189,N_1595,N_1717);
nand U2190 (N_2190,N_1572,N_1727);
or U2191 (N_2191,N_1527,N_1675);
and U2192 (N_2192,N_1743,N_1808);
or U2193 (N_2193,N_1697,N_1654);
nor U2194 (N_2194,N_1815,N_1886);
nor U2195 (N_2195,N_1511,N_1907);
nand U2196 (N_2196,N_1746,N_1935);
nor U2197 (N_2197,N_1918,N_1789);
nand U2198 (N_2198,N_1897,N_1530);
or U2199 (N_2199,N_1656,N_1905);
nor U2200 (N_2200,N_1582,N_1650);
and U2201 (N_2201,N_1900,N_1537);
nand U2202 (N_2202,N_1760,N_1803);
and U2203 (N_2203,N_1510,N_1894);
or U2204 (N_2204,N_1763,N_1703);
nor U2205 (N_2205,N_1577,N_1625);
xnor U2206 (N_2206,N_1657,N_1672);
and U2207 (N_2207,N_1617,N_1849);
or U2208 (N_2208,N_1720,N_1956);
xnor U2209 (N_2209,N_1865,N_1985);
or U2210 (N_2210,N_1924,N_1796);
nand U2211 (N_2211,N_1683,N_1667);
nand U2212 (N_2212,N_1839,N_1679);
nor U2213 (N_2213,N_1863,N_1757);
nand U2214 (N_2214,N_1719,N_1603);
and U2215 (N_2215,N_1931,N_1570);
and U2216 (N_2216,N_1969,N_1748);
xnor U2217 (N_2217,N_1589,N_1597);
nor U2218 (N_2218,N_1773,N_1775);
nor U2219 (N_2219,N_1835,N_1890);
nand U2220 (N_2220,N_1965,N_1524);
or U2221 (N_2221,N_1682,N_1801);
nor U2222 (N_2222,N_1810,N_1745);
nand U2223 (N_2223,N_1817,N_1579);
nor U2224 (N_2224,N_1864,N_1691);
nor U2225 (N_2225,N_1509,N_1704);
or U2226 (N_2226,N_1653,N_1664);
nand U2227 (N_2227,N_1590,N_1824);
or U2228 (N_2228,N_1791,N_1873);
nand U2229 (N_2229,N_1614,N_1925);
nor U2230 (N_2230,N_1722,N_1599);
nand U2231 (N_2231,N_1792,N_1581);
nor U2232 (N_2232,N_1535,N_1505);
nor U2233 (N_2233,N_1862,N_1643);
or U2234 (N_2234,N_1562,N_1874);
and U2235 (N_2235,N_1798,N_1533);
nand U2236 (N_2236,N_1866,N_1778);
nand U2237 (N_2237,N_1573,N_1585);
or U2238 (N_2238,N_1851,N_1729);
nand U2239 (N_2239,N_1721,N_1888);
and U2240 (N_2240,N_1586,N_1971);
and U2241 (N_2241,N_1592,N_1639);
nand U2242 (N_2242,N_1670,N_1867);
nor U2243 (N_2243,N_1974,N_1795);
nand U2244 (N_2244,N_1647,N_1941);
nor U2245 (N_2245,N_1800,N_1732);
and U2246 (N_2246,N_1584,N_1588);
nor U2247 (N_2247,N_1706,N_1600);
nand U2248 (N_2248,N_1514,N_1781);
nor U2249 (N_2249,N_1856,N_1854);
nand U2250 (N_2250,N_1819,N_1673);
or U2251 (N_2251,N_1741,N_1839);
nand U2252 (N_2252,N_1818,N_1568);
nor U2253 (N_2253,N_1622,N_1915);
xor U2254 (N_2254,N_1811,N_1749);
or U2255 (N_2255,N_1588,N_1861);
and U2256 (N_2256,N_1831,N_1506);
nor U2257 (N_2257,N_1719,N_1989);
or U2258 (N_2258,N_1741,N_1677);
nor U2259 (N_2259,N_1939,N_1904);
nor U2260 (N_2260,N_1788,N_1626);
nand U2261 (N_2261,N_1989,N_1819);
nor U2262 (N_2262,N_1850,N_1686);
and U2263 (N_2263,N_1770,N_1879);
or U2264 (N_2264,N_1609,N_1558);
and U2265 (N_2265,N_1522,N_1908);
or U2266 (N_2266,N_1545,N_1838);
nand U2267 (N_2267,N_1872,N_1905);
nand U2268 (N_2268,N_1936,N_1535);
and U2269 (N_2269,N_1613,N_1934);
and U2270 (N_2270,N_1538,N_1532);
and U2271 (N_2271,N_1716,N_1881);
or U2272 (N_2272,N_1676,N_1710);
and U2273 (N_2273,N_1909,N_1652);
nor U2274 (N_2274,N_1900,N_1551);
or U2275 (N_2275,N_1568,N_1617);
nor U2276 (N_2276,N_1553,N_1656);
nor U2277 (N_2277,N_1945,N_1898);
nand U2278 (N_2278,N_1654,N_1743);
and U2279 (N_2279,N_1553,N_1511);
or U2280 (N_2280,N_1876,N_1838);
or U2281 (N_2281,N_1891,N_1862);
or U2282 (N_2282,N_1619,N_1659);
nand U2283 (N_2283,N_1646,N_1683);
xor U2284 (N_2284,N_1975,N_1961);
and U2285 (N_2285,N_1671,N_1786);
and U2286 (N_2286,N_1884,N_1626);
or U2287 (N_2287,N_1680,N_1602);
and U2288 (N_2288,N_1847,N_1580);
nor U2289 (N_2289,N_1548,N_1631);
nor U2290 (N_2290,N_1719,N_1899);
nor U2291 (N_2291,N_1619,N_1800);
nand U2292 (N_2292,N_1538,N_1946);
and U2293 (N_2293,N_1644,N_1796);
nor U2294 (N_2294,N_1997,N_1602);
nor U2295 (N_2295,N_1760,N_1878);
or U2296 (N_2296,N_1548,N_1551);
nor U2297 (N_2297,N_1593,N_1652);
or U2298 (N_2298,N_1573,N_1676);
nor U2299 (N_2299,N_1638,N_1886);
nor U2300 (N_2300,N_1644,N_1767);
nor U2301 (N_2301,N_1629,N_1605);
or U2302 (N_2302,N_1555,N_1506);
and U2303 (N_2303,N_1800,N_1968);
and U2304 (N_2304,N_1807,N_1548);
or U2305 (N_2305,N_1518,N_1826);
nor U2306 (N_2306,N_1906,N_1547);
and U2307 (N_2307,N_1687,N_1691);
nand U2308 (N_2308,N_1597,N_1643);
and U2309 (N_2309,N_1531,N_1901);
nand U2310 (N_2310,N_1821,N_1904);
and U2311 (N_2311,N_1907,N_1577);
nor U2312 (N_2312,N_1990,N_1924);
or U2313 (N_2313,N_1569,N_1954);
nor U2314 (N_2314,N_1979,N_1904);
nor U2315 (N_2315,N_1841,N_1750);
nor U2316 (N_2316,N_1981,N_1577);
nor U2317 (N_2317,N_1562,N_1945);
nor U2318 (N_2318,N_1815,N_1722);
and U2319 (N_2319,N_1642,N_1797);
nor U2320 (N_2320,N_1580,N_1911);
nand U2321 (N_2321,N_1881,N_1516);
and U2322 (N_2322,N_1722,N_1813);
nand U2323 (N_2323,N_1870,N_1812);
nand U2324 (N_2324,N_1626,N_1924);
nor U2325 (N_2325,N_1558,N_1752);
nor U2326 (N_2326,N_1651,N_1712);
nor U2327 (N_2327,N_1649,N_1789);
and U2328 (N_2328,N_1677,N_1777);
xnor U2329 (N_2329,N_1625,N_1512);
nor U2330 (N_2330,N_1587,N_1869);
nand U2331 (N_2331,N_1850,N_1914);
and U2332 (N_2332,N_1921,N_1999);
and U2333 (N_2333,N_1721,N_1517);
nor U2334 (N_2334,N_1758,N_1590);
nand U2335 (N_2335,N_1606,N_1660);
nor U2336 (N_2336,N_1655,N_1568);
nand U2337 (N_2337,N_1552,N_1710);
and U2338 (N_2338,N_1647,N_1913);
and U2339 (N_2339,N_1574,N_1828);
nand U2340 (N_2340,N_1673,N_1766);
nand U2341 (N_2341,N_1626,N_1618);
nand U2342 (N_2342,N_1568,N_1741);
and U2343 (N_2343,N_1667,N_1648);
and U2344 (N_2344,N_1678,N_1803);
or U2345 (N_2345,N_1951,N_1595);
and U2346 (N_2346,N_1567,N_1512);
or U2347 (N_2347,N_1685,N_1636);
or U2348 (N_2348,N_1680,N_1706);
or U2349 (N_2349,N_1505,N_1735);
nor U2350 (N_2350,N_1907,N_1500);
and U2351 (N_2351,N_1676,N_1910);
xnor U2352 (N_2352,N_1665,N_1755);
and U2353 (N_2353,N_1621,N_1751);
nor U2354 (N_2354,N_1710,N_1875);
nor U2355 (N_2355,N_1607,N_1972);
or U2356 (N_2356,N_1861,N_1712);
and U2357 (N_2357,N_1636,N_1617);
nor U2358 (N_2358,N_1854,N_1573);
nand U2359 (N_2359,N_1601,N_1980);
nor U2360 (N_2360,N_1993,N_1722);
nand U2361 (N_2361,N_1822,N_1727);
nor U2362 (N_2362,N_1892,N_1823);
nor U2363 (N_2363,N_1580,N_1894);
nor U2364 (N_2364,N_1690,N_1676);
and U2365 (N_2365,N_1519,N_1554);
nand U2366 (N_2366,N_1954,N_1656);
and U2367 (N_2367,N_1702,N_1829);
nor U2368 (N_2368,N_1787,N_1791);
nand U2369 (N_2369,N_1511,N_1969);
nor U2370 (N_2370,N_1514,N_1855);
and U2371 (N_2371,N_1613,N_1618);
nor U2372 (N_2372,N_1808,N_1654);
or U2373 (N_2373,N_1941,N_1973);
and U2374 (N_2374,N_1741,N_1868);
or U2375 (N_2375,N_1866,N_1799);
nor U2376 (N_2376,N_1804,N_1560);
nor U2377 (N_2377,N_1843,N_1975);
nand U2378 (N_2378,N_1660,N_1535);
or U2379 (N_2379,N_1588,N_1919);
or U2380 (N_2380,N_1676,N_1601);
nor U2381 (N_2381,N_1865,N_1779);
and U2382 (N_2382,N_1794,N_1747);
and U2383 (N_2383,N_1876,N_1790);
nor U2384 (N_2384,N_1994,N_1849);
and U2385 (N_2385,N_1940,N_1568);
nand U2386 (N_2386,N_1660,N_1865);
or U2387 (N_2387,N_1948,N_1954);
and U2388 (N_2388,N_1630,N_1684);
or U2389 (N_2389,N_1775,N_1782);
nor U2390 (N_2390,N_1701,N_1734);
xor U2391 (N_2391,N_1736,N_1760);
nor U2392 (N_2392,N_1773,N_1519);
nand U2393 (N_2393,N_1718,N_1940);
or U2394 (N_2394,N_1700,N_1555);
nor U2395 (N_2395,N_1936,N_1525);
and U2396 (N_2396,N_1629,N_1794);
or U2397 (N_2397,N_1756,N_1708);
nor U2398 (N_2398,N_1832,N_1646);
nor U2399 (N_2399,N_1727,N_1978);
nand U2400 (N_2400,N_1575,N_1926);
nor U2401 (N_2401,N_1750,N_1927);
nand U2402 (N_2402,N_1772,N_1706);
nand U2403 (N_2403,N_1516,N_1808);
nor U2404 (N_2404,N_1603,N_1636);
nand U2405 (N_2405,N_1526,N_1841);
and U2406 (N_2406,N_1905,N_1776);
nand U2407 (N_2407,N_1672,N_1707);
nand U2408 (N_2408,N_1742,N_1819);
or U2409 (N_2409,N_1720,N_1902);
nor U2410 (N_2410,N_1838,N_1720);
nor U2411 (N_2411,N_1970,N_1678);
and U2412 (N_2412,N_1913,N_1826);
nand U2413 (N_2413,N_1909,N_1694);
nor U2414 (N_2414,N_1987,N_1699);
nand U2415 (N_2415,N_1764,N_1910);
nor U2416 (N_2416,N_1798,N_1512);
and U2417 (N_2417,N_1809,N_1793);
and U2418 (N_2418,N_1972,N_1653);
or U2419 (N_2419,N_1971,N_1615);
and U2420 (N_2420,N_1924,N_1844);
or U2421 (N_2421,N_1779,N_1831);
or U2422 (N_2422,N_1899,N_1910);
and U2423 (N_2423,N_1749,N_1740);
or U2424 (N_2424,N_1509,N_1826);
nor U2425 (N_2425,N_1678,N_1532);
and U2426 (N_2426,N_1801,N_1541);
nand U2427 (N_2427,N_1525,N_1886);
nor U2428 (N_2428,N_1995,N_1601);
and U2429 (N_2429,N_1681,N_1634);
nand U2430 (N_2430,N_1561,N_1585);
or U2431 (N_2431,N_1832,N_1785);
nor U2432 (N_2432,N_1542,N_1537);
nor U2433 (N_2433,N_1949,N_1774);
and U2434 (N_2434,N_1849,N_1550);
nand U2435 (N_2435,N_1853,N_1517);
or U2436 (N_2436,N_1599,N_1990);
nor U2437 (N_2437,N_1847,N_1867);
and U2438 (N_2438,N_1757,N_1540);
nand U2439 (N_2439,N_1748,N_1764);
or U2440 (N_2440,N_1654,N_1818);
nand U2441 (N_2441,N_1654,N_1578);
nand U2442 (N_2442,N_1995,N_1849);
and U2443 (N_2443,N_1517,N_1980);
nand U2444 (N_2444,N_1768,N_1935);
nor U2445 (N_2445,N_1929,N_1999);
or U2446 (N_2446,N_1882,N_1810);
nor U2447 (N_2447,N_1805,N_1777);
or U2448 (N_2448,N_1828,N_1596);
and U2449 (N_2449,N_1940,N_1906);
or U2450 (N_2450,N_1896,N_1801);
nor U2451 (N_2451,N_1937,N_1704);
xnor U2452 (N_2452,N_1842,N_1732);
nor U2453 (N_2453,N_1520,N_1647);
nand U2454 (N_2454,N_1541,N_1588);
nor U2455 (N_2455,N_1738,N_1894);
or U2456 (N_2456,N_1508,N_1511);
nor U2457 (N_2457,N_1535,N_1542);
and U2458 (N_2458,N_1687,N_1536);
or U2459 (N_2459,N_1571,N_1777);
nor U2460 (N_2460,N_1898,N_1748);
nand U2461 (N_2461,N_1827,N_1605);
nand U2462 (N_2462,N_1766,N_1968);
and U2463 (N_2463,N_1809,N_1762);
or U2464 (N_2464,N_1954,N_1600);
nand U2465 (N_2465,N_1779,N_1951);
nor U2466 (N_2466,N_1514,N_1646);
nand U2467 (N_2467,N_1588,N_1614);
or U2468 (N_2468,N_1943,N_1868);
nand U2469 (N_2469,N_1728,N_1863);
and U2470 (N_2470,N_1658,N_1705);
or U2471 (N_2471,N_1766,N_1723);
nor U2472 (N_2472,N_1978,N_1975);
nor U2473 (N_2473,N_1697,N_1784);
or U2474 (N_2474,N_1937,N_1898);
nor U2475 (N_2475,N_1604,N_1768);
nand U2476 (N_2476,N_1626,N_1524);
and U2477 (N_2477,N_1972,N_1774);
or U2478 (N_2478,N_1878,N_1981);
nand U2479 (N_2479,N_1512,N_1748);
or U2480 (N_2480,N_1701,N_1902);
and U2481 (N_2481,N_1771,N_1853);
nor U2482 (N_2482,N_1723,N_1870);
nand U2483 (N_2483,N_1844,N_1560);
and U2484 (N_2484,N_1841,N_1534);
and U2485 (N_2485,N_1628,N_1636);
and U2486 (N_2486,N_1578,N_1630);
or U2487 (N_2487,N_1890,N_1675);
or U2488 (N_2488,N_1908,N_1799);
nand U2489 (N_2489,N_1576,N_1728);
or U2490 (N_2490,N_1725,N_1826);
and U2491 (N_2491,N_1757,N_1659);
nor U2492 (N_2492,N_1856,N_1791);
nor U2493 (N_2493,N_1752,N_1913);
or U2494 (N_2494,N_1750,N_1871);
and U2495 (N_2495,N_1660,N_1802);
or U2496 (N_2496,N_1819,N_1636);
nor U2497 (N_2497,N_1528,N_1895);
nor U2498 (N_2498,N_1802,N_1957);
nor U2499 (N_2499,N_1886,N_1657);
and U2500 (N_2500,N_2151,N_2109);
or U2501 (N_2501,N_2396,N_2329);
and U2502 (N_2502,N_2223,N_2257);
or U2503 (N_2503,N_2243,N_2429);
nor U2504 (N_2504,N_2069,N_2014);
or U2505 (N_2505,N_2205,N_2310);
nor U2506 (N_2506,N_2141,N_2334);
or U2507 (N_2507,N_2318,N_2388);
and U2508 (N_2508,N_2174,N_2186);
and U2509 (N_2509,N_2082,N_2092);
and U2510 (N_2510,N_2458,N_2013);
and U2511 (N_2511,N_2282,N_2441);
nor U2512 (N_2512,N_2316,N_2049);
or U2513 (N_2513,N_2083,N_2454);
nor U2514 (N_2514,N_2315,N_2161);
or U2515 (N_2515,N_2036,N_2279);
nand U2516 (N_2516,N_2299,N_2154);
or U2517 (N_2517,N_2107,N_2380);
or U2518 (N_2518,N_2032,N_2152);
nor U2519 (N_2519,N_2215,N_2081);
nand U2520 (N_2520,N_2187,N_2037);
or U2521 (N_2521,N_2123,N_2115);
nor U2522 (N_2522,N_2440,N_2355);
nor U2523 (N_2523,N_2136,N_2012);
nor U2524 (N_2524,N_2073,N_2264);
and U2525 (N_2525,N_2090,N_2241);
nor U2526 (N_2526,N_2006,N_2095);
nand U2527 (N_2527,N_2072,N_2457);
nor U2528 (N_2528,N_2419,N_2056);
nor U2529 (N_2529,N_2498,N_2084);
and U2530 (N_2530,N_2167,N_2459);
nand U2531 (N_2531,N_2331,N_2010);
and U2532 (N_2532,N_2265,N_2430);
nand U2533 (N_2533,N_2249,N_2127);
nand U2534 (N_2534,N_2426,N_2170);
nor U2535 (N_2535,N_2022,N_2319);
and U2536 (N_2536,N_2119,N_2134);
nand U2537 (N_2537,N_2475,N_2280);
nor U2538 (N_2538,N_2252,N_2066);
or U2539 (N_2539,N_2325,N_2444);
and U2540 (N_2540,N_2307,N_2484);
or U2541 (N_2541,N_2412,N_2131);
or U2542 (N_2542,N_2428,N_2333);
or U2543 (N_2543,N_2464,N_2338);
nor U2544 (N_2544,N_2213,N_2352);
or U2545 (N_2545,N_2108,N_2422);
nor U2546 (N_2546,N_2079,N_2350);
nor U2547 (N_2547,N_2204,N_2099);
nor U2548 (N_2548,N_2258,N_2229);
and U2549 (N_2549,N_2017,N_2046);
or U2550 (N_2550,N_2261,N_2237);
nor U2551 (N_2551,N_2025,N_2034);
nor U2552 (N_2552,N_2283,N_2358);
nor U2553 (N_2553,N_2030,N_2183);
and U2554 (N_2554,N_2011,N_2337);
and U2555 (N_2555,N_2271,N_2449);
nor U2556 (N_2556,N_2489,N_2044);
nand U2557 (N_2557,N_2005,N_2179);
and U2558 (N_2558,N_2364,N_2004);
nor U2559 (N_2559,N_2041,N_2497);
and U2560 (N_2560,N_2365,N_2322);
xnor U2561 (N_2561,N_2147,N_2112);
nand U2562 (N_2562,N_2086,N_2348);
or U2563 (N_2563,N_2102,N_2418);
or U2564 (N_2564,N_2201,N_2436);
or U2565 (N_2565,N_2461,N_2155);
or U2566 (N_2566,N_2050,N_2111);
nor U2567 (N_2567,N_2055,N_2381);
or U2568 (N_2568,N_2376,N_2217);
nor U2569 (N_2569,N_2284,N_2297);
nand U2570 (N_2570,N_2002,N_2210);
or U2571 (N_2571,N_2130,N_2052);
or U2572 (N_2572,N_2270,N_2339);
nor U2573 (N_2573,N_2374,N_2024);
or U2574 (N_2574,N_2373,N_2114);
nor U2575 (N_2575,N_2239,N_2197);
or U2576 (N_2576,N_2476,N_2230);
or U2577 (N_2577,N_2026,N_2477);
and U2578 (N_2578,N_2240,N_2203);
and U2579 (N_2579,N_2278,N_2324);
nor U2580 (N_2580,N_2456,N_2409);
nand U2581 (N_2581,N_2450,N_2043);
nor U2582 (N_2582,N_2251,N_2490);
and U2583 (N_2583,N_2145,N_2173);
nand U2584 (N_2584,N_2312,N_2100);
nand U2585 (N_2585,N_2238,N_2447);
and U2586 (N_2586,N_2360,N_2070);
and U2587 (N_2587,N_2298,N_2367);
nand U2588 (N_2588,N_2274,N_2277);
nand U2589 (N_2589,N_2033,N_2295);
nor U2590 (N_2590,N_2078,N_2227);
or U2591 (N_2591,N_2347,N_2425);
and U2592 (N_2592,N_2077,N_2200);
nor U2593 (N_2593,N_2138,N_2062);
nand U2594 (N_2594,N_2420,N_2465);
nor U2595 (N_2595,N_2047,N_2424);
or U2596 (N_2596,N_2341,N_2309);
xor U2597 (N_2597,N_2494,N_2051);
nand U2598 (N_2598,N_2357,N_2402);
nor U2599 (N_2599,N_2300,N_2222);
and U2600 (N_2600,N_2122,N_2394);
nand U2601 (N_2601,N_2260,N_2427);
or U2602 (N_2602,N_2410,N_2031);
nor U2603 (N_2603,N_2413,N_2445);
and U2604 (N_2604,N_2080,N_2281);
nor U2605 (N_2605,N_2291,N_2190);
nor U2606 (N_2606,N_2142,N_2220);
and U2607 (N_2607,N_2434,N_2481);
or U2608 (N_2608,N_2496,N_2221);
nor U2609 (N_2609,N_2391,N_2015);
or U2610 (N_2610,N_2242,N_2219);
nand U2611 (N_2611,N_2343,N_2178);
nand U2612 (N_2612,N_2415,N_2185);
nor U2613 (N_2613,N_2029,N_2231);
or U2614 (N_2614,N_2269,N_2305);
nor U2615 (N_2615,N_2294,N_2483);
nand U2616 (N_2616,N_2275,N_2349);
and U2617 (N_2617,N_2035,N_2354);
and U2618 (N_2618,N_2168,N_2495);
or U2619 (N_2619,N_2019,N_2214);
and U2620 (N_2620,N_2194,N_2383);
and U2621 (N_2621,N_2110,N_2491);
nor U2622 (N_2622,N_2172,N_2106);
nand U2623 (N_2623,N_2267,N_2384);
or U2624 (N_2624,N_2370,N_2443);
or U2625 (N_2625,N_2001,N_2328);
or U2626 (N_2626,N_2135,N_2228);
nand U2627 (N_2627,N_2074,N_2336);
nor U2628 (N_2628,N_2385,N_2163);
and U2629 (N_2629,N_2361,N_2027);
nor U2630 (N_2630,N_2306,N_2262);
or U2631 (N_2631,N_2156,N_2304);
nor U2632 (N_2632,N_2403,N_2254);
nand U2633 (N_2633,N_2202,N_2301);
nand U2634 (N_2634,N_2438,N_2144);
or U2635 (N_2635,N_2149,N_2075);
or U2636 (N_2636,N_2302,N_2129);
or U2637 (N_2637,N_2089,N_2366);
nor U2638 (N_2638,N_2256,N_2382);
and U2639 (N_2639,N_2473,N_2063);
and U2640 (N_2640,N_2093,N_2191);
nand U2641 (N_2641,N_2068,N_2390);
xor U2642 (N_2642,N_2276,N_2054);
or U2643 (N_2643,N_2346,N_2375);
nand U2644 (N_2644,N_2368,N_2113);
nor U2645 (N_2645,N_2235,N_2345);
or U2646 (N_2646,N_2259,N_2059);
nand U2647 (N_2647,N_2393,N_2314);
nor U2648 (N_2648,N_2218,N_2404);
and U2649 (N_2649,N_2146,N_2018);
nand U2650 (N_2650,N_2485,N_2362);
nor U2651 (N_2651,N_2016,N_2407);
and U2652 (N_2652,N_2266,N_2323);
or U2653 (N_2653,N_2389,N_2303);
nand U2654 (N_2654,N_2285,N_2332);
and U2655 (N_2655,N_2293,N_2363);
or U2656 (N_2656,N_2175,N_2245);
or U2657 (N_2657,N_2166,N_2096);
nor U2658 (N_2658,N_2273,N_2248);
or U2659 (N_2659,N_2246,N_2133);
or U2660 (N_2660,N_2263,N_2128);
and U2661 (N_2661,N_2207,N_2148);
nor U2662 (N_2662,N_2028,N_2061);
nor U2663 (N_2663,N_2023,N_2158);
nor U2664 (N_2664,N_2125,N_2164);
nor U2665 (N_2665,N_2225,N_2209);
or U2666 (N_2666,N_2021,N_2091);
nor U2667 (N_2667,N_2467,N_2493);
nor U2668 (N_2668,N_2103,N_2272);
and U2669 (N_2669,N_2097,N_2342);
and U2670 (N_2670,N_2372,N_2208);
or U2671 (N_2671,N_2188,N_2399);
and U2672 (N_2672,N_2058,N_2432);
and U2673 (N_2673,N_2488,N_2401);
nor U2674 (N_2674,N_2326,N_2460);
nor U2675 (N_2675,N_2369,N_2289);
nand U2676 (N_2676,N_2233,N_2153);
and U2677 (N_2677,N_2181,N_2417);
nand U2678 (N_2678,N_2048,N_2397);
nor U2679 (N_2679,N_2060,N_2292);
nand U2680 (N_2680,N_2020,N_2439);
or U2681 (N_2681,N_2453,N_2437);
nand U2682 (N_2682,N_2150,N_2196);
nor U2683 (N_2683,N_2340,N_2189);
nor U2684 (N_2684,N_2255,N_2126);
and U2685 (N_2685,N_2253,N_2165);
or U2686 (N_2686,N_2492,N_2479);
and U2687 (N_2687,N_2250,N_2226);
nand U2688 (N_2688,N_2000,N_2038);
nand U2689 (N_2689,N_2120,N_2177);
or U2690 (N_2690,N_2040,N_2320);
nand U2691 (N_2691,N_2169,N_2311);
or U2692 (N_2692,N_2198,N_2317);
nor U2693 (N_2693,N_2212,N_2121);
xor U2694 (N_2694,N_2486,N_2104);
nand U2695 (N_2695,N_2124,N_2139);
nor U2696 (N_2696,N_2101,N_2431);
and U2697 (N_2697,N_2435,N_2007);
or U2698 (N_2698,N_2414,N_2421);
nor U2699 (N_2699,N_2232,N_2351);
and U2700 (N_2700,N_2065,N_2499);
nor U2701 (N_2701,N_2480,N_2094);
or U2702 (N_2702,N_2448,N_2433);
nor U2703 (N_2703,N_2057,N_2474);
or U2704 (N_2704,N_2268,N_2359);
nor U2705 (N_2705,N_2184,N_2160);
or U2706 (N_2706,N_2117,N_2171);
nor U2707 (N_2707,N_2137,N_2442);
or U2708 (N_2708,N_2470,N_2408);
or U2709 (N_2709,N_2088,N_2159);
or U2710 (N_2710,N_2193,N_2462);
nand U2711 (N_2711,N_2405,N_2353);
nor U2712 (N_2712,N_2321,N_2118);
nor U2713 (N_2713,N_2344,N_2206);
and U2714 (N_2714,N_2471,N_2045);
nand U2715 (N_2715,N_2287,N_2236);
and U2716 (N_2716,N_2286,N_2335);
nand U2717 (N_2717,N_2466,N_2216);
nor U2718 (N_2718,N_2482,N_2469);
or U2719 (N_2719,N_2463,N_2039);
nor U2720 (N_2720,N_2009,N_2371);
and U2721 (N_2721,N_2451,N_2085);
or U2722 (N_2722,N_2327,N_2157);
or U2723 (N_2723,N_2290,N_2395);
and U2724 (N_2724,N_2105,N_2067);
and U2725 (N_2725,N_2392,N_2162);
nor U2726 (N_2726,N_2455,N_2377);
or U2727 (N_2727,N_2042,N_2132);
or U2728 (N_2728,N_2180,N_2313);
nor U2729 (N_2729,N_2386,N_2296);
nand U2730 (N_2730,N_2356,N_2176);
nand U2731 (N_2731,N_2288,N_2143);
nand U2732 (N_2732,N_2098,N_2199);
nor U2733 (N_2733,N_2195,N_2446);
or U2734 (N_2734,N_2398,N_2478);
and U2735 (N_2735,N_2487,N_2247);
and U2736 (N_2736,N_2411,N_2387);
or U2737 (N_2737,N_2472,N_2140);
nor U2738 (N_2738,N_2224,N_2003);
nor U2739 (N_2739,N_2406,N_2244);
nand U2740 (N_2740,N_2071,N_2211);
and U2741 (N_2741,N_2308,N_2182);
nor U2742 (N_2742,N_2076,N_2234);
or U2743 (N_2743,N_2116,N_2416);
nor U2744 (N_2744,N_2087,N_2330);
and U2745 (N_2745,N_2378,N_2468);
nor U2746 (N_2746,N_2192,N_2452);
xnor U2747 (N_2747,N_2423,N_2379);
and U2748 (N_2748,N_2053,N_2008);
nand U2749 (N_2749,N_2064,N_2400);
or U2750 (N_2750,N_2396,N_2355);
and U2751 (N_2751,N_2148,N_2054);
nand U2752 (N_2752,N_2047,N_2179);
nor U2753 (N_2753,N_2435,N_2492);
nor U2754 (N_2754,N_2435,N_2473);
or U2755 (N_2755,N_2314,N_2499);
nor U2756 (N_2756,N_2066,N_2013);
nand U2757 (N_2757,N_2360,N_2246);
nand U2758 (N_2758,N_2388,N_2442);
xor U2759 (N_2759,N_2043,N_2306);
nand U2760 (N_2760,N_2241,N_2151);
and U2761 (N_2761,N_2485,N_2300);
and U2762 (N_2762,N_2213,N_2132);
nand U2763 (N_2763,N_2042,N_2399);
or U2764 (N_2764,N_2398,N_2401);
nand U2765 (N_2765,N_2493,N_2341);
nor U2766 (N_2766,N_2098,N_2130);
nand U2767 (N_2767,N_2402,N_2093);
nand U2768 (N_2768,N_2439,N_2125);
nor U2769 (N_2769,N_2171,N_2144);
nor U2770 (N_2770,N_2095,N_2056);
and U2771 (N_2771,N_2211,N_2120);
nand U2772 (N_2772,N_2321,N_2158);
nand U2773 (N_2773,N_2479,N_2009);
or U2774 (N_2774,N_2441,N_2036);
nand U2775 (N_2775,N_2421,N_2196);
and U2776 (N_2776,N_2106,N_2251);
nand U2777 (N_2777,N_2080,N_2054);
nand U2778 (N_2778,N_2114,N_2388);
and U2779 (N_2779,N_2075,N_2002);
nor U2780 (N_2780,N_2015,N_2014);
nand U2781 (N_2781,N_2472,N_2236);
or U2782 (N_2782,N_2091,N_2374);
and U2783 (N_2783,N_2093,N_2225);
and U2784 (N_2784,N_2386,N_2464);
xnor U2785 (N_2785,N_2321,N_2257);
nand U2786 (N_2786,N_2161,N_2263);
nand U2787 (N_2787,N_2437,N_2141);
nor U2788 (N_2788,N_2436,N_2243);
or U2789 (N_2789,N_2314,N_2129);
nand U2790 (N_2790,N_2292,N_2255);
nand U2791 (N_2791,N_2105,N_2085);
nand U2792 (N_2792,N_2336,N_2008);
nor U2793 (N_2793,N_2069,N_2079);
xnor U2794 (N_2794,N_2450,N_2253);
and U2795 (N_2795,N_2499,N_2083);
and U2796 (N_2796,N_2285,N_2094);
or U2797 (N_2797,N_2284,N_2438);
and U2798 (N_2798,N_2257,N_2133);
or U2799 (N_2799,N_2040,N_2115);
nand U2800 (N_2800,N_2244,N_2387);
nand U2801 (N_2801,N_2469,N_2465);
nor U2802 (N_2802,N_2278,N_2429);
nand U2803 (N_2803,N_2154,N_2159);
and U2804 (N_2804,N_2084,N_2246);
nand U2805 (N_2805,N_2395,N_2068);
or U2806 (N_2806,N_2488,N_2133);
nand U2807 (N_2807,N_2169,N_2401);
and U2808 (N_2808,N_2454,N_2270);
and U2809 (N_2809,N_2253,N_2478);
nor U2810 (N_2810,N_2476,N_2220);
and U2811 (N_2811,N_2236,N_2155);
nor U2812 (N_2812,N_2322,N_2496);
and U2813 (N_2813,N_2456,N_2436);
nor U2814 (N_2814,N_2095,N_2378);
nand U2815 (N_2815,N_2342,N_2300);
nand U2816 (N_2816,N_2004,N_2473);
or U2817 (N_2817,N_2257,N_2091);
and U2818 (N_2818,N_2163,N_2128);
or U2819 (N_2819,N_2132,N_2253);
nand U2820 (N_2820,N_2216,N_2326);
and U2821 (N_2821,N_2057,N_2273);
nor U2822 (N_2822,N_2030,N_2203);
and U2823 (N_2823,N_2195,N_2016);
or U2824 (N_2824,N_2080,N_2115);
nor U2825 (N_2825,N_2466,N_2023);
nand U2826 (N_2826,N_2320,N_2134);
or U2827 (N_2827,N_2293,N_2085);
and U2828 (N_2828,N_2323,N_2493);
nand U2829 (N_2829,N_2292,N_2278);
nor U2830 (N_2830,N_2403,N_2341);
and U2831 (N_2831,N_2467,N_2290);
nand U2832 (N_2832,N_2200,N_2154);
and U2833 (N_2833,N_2144,N_2404);
nand U2834 (N_2834,N_2306,N_2199);
or U2835 (N_2835,N_2253,N_2491);
or U2836 (N_2836,N_2110,N_2215);
and U2837 (N_2837,N_2405,N_2499);
and U2838 (N_2838,N_2401,N_2076);
nand U2839 (N_2839,N_2079,N_2134);
nand U2840 (N_2840,N_2361,N_2164);
and U2841 (N_2841,N_2050,N_2467);
nand U2842 (N_2842,N_2405,N_2471);
and U2843 (N_2843,N_2467,N_2355);
or U2844 (N_2844,N_2432,N_2401);
nand U2845 (N_2845,N_2312,N_2244);
or U2846 (N_2846,N_2425,N_2292);
or U2847 (N_2847,N_2379,N_2033);
xor U2848 (N_2848,N_2369,N_2036);
nor U2849 (N_2849,N_2361,N_2386);
nand U2850 (N_2850,N_2065,N_2271);
or U2851 (N_2851,N_2326,N_2323);
and U2852 (N_2852,N_2257,N_2194);
or U2853 (N_2853,N_2305,N_2281);
nor U2854 (N_2854,N_2065,N_2243);
and U2855 (N_2855,N_2104,N_2063);
nand U2856 (N_2856,N_2417,N_2415);
or U2857 (N_2857,N_2360,N_2149);
nand U2858 (N_2858,N_2249,N_2351);
nand U2859 (N_2859,N_2292,N_2224);
nand U2860 (N_2860,N_2058,N_2226);
and U2861 (N_2861,N_2032,N_2024);
or U2862 (N_2862,N_2171,N_2421);
nand U2863 (N_2863,N_2482,N_2378);
and U2864 (N_2864,N_2104,N_2482);
nand U2865 (N_2865,N_2398,N_2314);
or U2866 (N_2866,N_2081,N_2451);
or U2867 (N_2867,N_2378,N_2194);
nand U2868 (N_2868,N_2421,N_2116);
nor U2869 (N_2869,N_2215,N_2360);
and U2870 (N_2870,N_2000,N_2082);
nor U2871 (N_2871,N_2376,N_2191);
and U2872 (N_2872,N_2479,N_2000);
or U2873 (N_2873,N_2224,N_2157);
or U2874 (N_2874,N_2043,N_2217);
nand U2875 (N_2875,N_2451,N_2426);
nand U2876 (N_2876,N_2426,N_2307);
and U2877 (N_2877,N_2259,N_2394);
and U2878 (N_2878,N_2363,N_2474);
or U2879 (N_2879,N_2237,N_2081);
or U2880 (N_2880,N_2140,N_2134);
nand U2881 (N_2881,N_2453,N_2305);
nor U2882 (N_2882,N_2352,N_2115);
nand U2883 (N_2883,N_2192,N_2205);
nand U2884 (N_2884,N_2093,N_2452);
and U2885 (N_2885,N_2277,N_2380);
or U2886 (N_2886,N_2408,N_2047);
nand U2887 (N_2887,N_2039,N_2454);
nor U2888 (N_2888,N_2174,N_2026);
and U2889 (N_2889,N_2082,N_2403);
nor U2890 (N_2890,N_2234,N_2295);
or U2891 (N_2891,N_2394,N_2476);
or U2892 (N_2892,N_2324,N_2185);
or U2893 (N_2893,N_2212,N_2456);
or U2894 (N_2894,N_2161,N_2304);
nor U2895 (N_2895,N_2414,N_2357);
nand U2896 (N_2896,N_2002,N_2304);
nor U2897 (N_2897,N_2106,N_2412);
and U2898 (N_2898,N_2213,N_2244);
nand U2899 (N_2899,N_2174,N_2499);
nand U2900 (N_2900,N_2315,N_2437);
nand U2901 (N_2901,N_2467,N_2049);
nor U2902 (N_2902,N_2464,N_2080);
or U2903 (N_2903,N_2105,N_2414);
and U2904 (N_2904,N_2234,N_2112);
or U2905 (N_2905,N_2197,N_2305);
xor U2906 (N_2906,N_2011,N_2407);
nand U2907 (N_2907,N_2333,N_2129);
nor U2908 (N_2908,N_2218,N_2477);
xor U2909 (N_2909,N_2342,N_2069);
nand U2910 (N_2910,N_2232,N_2436);
or U2911 (N_2911,N_2309,N_2290);
or U2912 (N_2912,N_2246,N_2401);
or U2913 (N_2913,N_2455,N_2357);
and U2914 (N_2914,N_2192,N_2480);
nand U2915 (N_2915,N_2248,N_2276);
nor U2916 (N_2916,N_2211,N_2268);
and U2917 (N_2917,N_2092,N_2116);
and U2918 (N_2918,N_2430,N_2088);
or U2919 (N_2919,N_2126,N_2124);
nor U2920 (N_2920,N_2242,N_2189);
nor U2921 (N_2921,N_2216,N_2360);
or U2922 (N_2922,N_2181,N_2036);
nor U2923 (N_2923,N_2218,N_2438);
nand U2924 (N_2924,N_2467,N_2169);
and U2925 (N_2925,N_2464,N_2405);
nor U2926 (N_2926,N_2360,N_2295);
and U2927 (N_2927,N_2156,N_2100);
nand U2928 (N_2928,N_2380,N_2086);
nor U2929 (N_2929,N_2373,N_2400);
or U2930 (N_2930,N_2453,N_2329);
or U2931 (N_2931,N_2115,N_2326);
nor U2932 (N_2932,N_2277,N_2302);
and U2933 (N_2933,N_2065,N_2070);
nor U2934 (N_2934,N_2306,N_2085);
nand U2935 (N_2935,N_2353,N_2282);
or U2936 (N_2936,N_2437,N_2061);
nand U2937 (N_2937,N_2296,N_2377);
and U2938 (N_2938,N_2394,N_2091);
and U2939 (N_2939,N_2450,N_2031);
or U2940 (N_2940,N_2101,N_2336);
nor U2941 (N_2941,N_2288,N_2168);
or U2942 (N_2942,N_2480,N_2295);
nor U2943 (N_2943,N_2477,N_2429);
nand U2944 (N_2944,N_2358,N_2012);
nand U2945 (N_2945,N_2133,N_2128);
nand U2946 (N_2946,N_2052,N_2442);
nor U2947 (N_2947,N_2141,N_2206);
or U2948 (N_2948,N_2145,N_2304);
or U2949 (N_2949,N_2104,N_2406);
nor U2950 (N_2950,N_2378,N_2383);
nand U2951 (N_2951,N_2058,N_2031);
nand U2952 (N_2952,N_2490,N_2336);
or U2953 (N_2953,N_2043,N_2346);
or U2954 (N_2954,N_2390,N_2005);
nand U2955 (N_2955,N_2153,N_2229);
or U2956 (N_2956,N_2459,N_2303);
nand U2957 (N_2957,N_2186,N_2006);
nand U2958 (N_2958,N_2259,N_2237);
nand U2959 (N_2959,N_2138,N_2348);
nand U2960 (N_2960,N_2147,N_2203);
and U2961 (N_2961,N_2371,N_2269);
or U2962 (N_2962,N_2088,N_2330);
nor U2963 (N_2963,N_2209,N_2145);
and U2964 (N_2964,N_2180,N_2145);
and U2965 (N_2965,N_2258,N_2212);
or U2966 (N_2966,N_2181,N_2391);
and U2967 (N_2967,N_2328,N_2190);
nand U2968 (N_2968,N_2018,N_2312);
or U2969 (N_2969,N_2220,N_2291);
nand U2970 (N_2970,N_2296,N_2215);
and U2971 (N_2971,N_2477,N_2057);
nand U2972 (N_2972,N_2235,N_2412);
nor U2973 (N_2973,N_2064,N_2288);
nor U2974 (N_2974,N_2387,N_2168);
nor U2975 (N_2975,N_2036,N_2341);
nand U2976 (N_2976,N_2189,N_2001);
nand U2977 (N_2977,N_2116,N_2040);
nor U2978 (N_2978,N_2407,N_2390);
and U2979 (N_2979,N_2434,N_2452);
or U2980 (N_2980,N_2136,N_2159);
nand U2981 (N_2981,N_2319,N_2355);
and U2982 (N_2982,N_2319,N_2393);
and U2983 (N_2983,N_2067,N_2109);
nor U2984 (N_2984,N_2165,N_2217);
nand U2985 (N_2985,N_2279,N_2122);
nand U2986 (N_2986,N_2428,N_2113);
nor U2987 (N_2987,N_2211,N_2112);
nor U2988 (N_2988,N_2145,N_2364);
or U2989 (N_2989,N_2174,N_2450);
or U2990 (N_2990,N_2089,N_2256);
or U2991 (N_2991,N_2381,N_2385);
nor U2992 (N_2992,N_2200,N_2471);
nor U2993 (N_2993,N_2114,N_2418);
or U2994 (N_2994,N_2139,N_2350);
or U2995 (N_2995,N_2267,N_2297);
nor U2996 (N_2996,N_2386,N_2195);
or U2997 (N_2997,N_2230,N_2444);
nor U2998 (N_2998,N_2362,N_2250);
nor U2999 (N_2999,N_2286,N_2155);
or U3000 (N_3000,N_2759,N_2543);
or U3001 (N_3001,N_2605,N_2980);
nor U3002 (N_3002,N_2767,N_2779);
nand U3003 (N_3003,N_2549,N_2925);
or U3004 (N_3004,N_2742,N_2915);
nand U3005 (N_3005,N_2973,N_2793);
nand U3006 (N_3006,N_2653,N_2849);
nor U3007 (N_3007,N_2539,N_2700);
nand U3008 (N_3008,N_2546,N_2967);
nor U3009 (N_3009,N_2703,N_2950);
nor U3010 (N_3010,N_2500,N_2707);
nand U3011 (N_3011,N_2981,N_2978);
or U3012 (N_3012,N_2773,N_2595);
or U3013 (N_3013,N_2762,N_2880);
nor U3014 (N_3014,N_2988,N_2725);
and U3015 (N_3015,N_2658,N_2809);
and U3016 (N_3016,N_2801,N_2839);
and U3017 (N_3017,N_2853,N_2506);
nor U3018 (N_3018,N_2600,N_2995);
nand U3019 (N_3019,N_2984,N_2528);
or U3020 (N_3020,N_2518,N_2642);
and U3021 (N_3021,N_2679,N_2895);
and U3022 (N_3022,N_2567,N_2774);
nand U3023 (N_3023,N_2515,N_2982);
nand U3024 (N_3024,N_2558,N_2743);
nand U3025 (N_3025,N_2667,N_2881);
and U3026 (N_3026,N_2805,N_2845);
or U3027 (N_3027,N_2798,N_2990);
or U3028 (N_3028,N_2908,N_2714);
nand U3029 (N_3029,N_2891,N_2766);
nand U3030 (N_3030,N_2717,N_2636);
or U3031 (N_3031,N_2641,N_2815);
nand U3032 (N_3032,N_2632,N_2581);
nor U3033 (N_3033,N_2735,N_2781);
nor U3034 (N_3034,N_2593,N_2624);
or U3035 (N_3035,N_2623,N_2724);
nand U3036 (N_3036,N_2813,N_2806);
and U3037 (N_3037,N_2587,N_2618);
nand U3038 (N_3038,N_2777,N_2789);
nand U3039 (N_3039,N_2873,N_2772);
nand U3040 (N_3040,N_2736,N_2657);
or U3041 (N_3041,N_2907,N_2927);
nand U3042 (N_3042,N_2812,N_2857);
and U3043 (N_3043,N_2942,N_2937);
nor U3044 (N_3044,N_2933,N_2918);
nand U3045 (N_3045,N_2723,N_2616);
nor U3046 (N_3046,N_2606,N_2770);
or U3047 (N_3047,N_2564,N_2843);
nand U3048 (N_3048,N_2877,N_2673);
nand U3049 (N_3049,N_2591,N_2934);
nand U3050 (N_3050,N_2956,N_2987);
and U3051 (N_3051,N_2569,N_2989);
or U3052 (N_3052,N_2530,N_2875);
nor U3053 (N_3053,N_2503,N_2921);
nor U3054 (N_3054,N_2741,N_2999);
nor U3055 (N_3055,N_2751,N_2599);
nor U3056 (N_3056,N_2696,N_2792);
or U3057 (N_3057,N_2512,N_2551);
or U3058 (N_3058,N_2951,N_2803);
or U3059 (N_3059,N_2722,N_2565);
nand U3060 (N_3060,N_2846,N_2834);
and U3061 (N_3061,N_2681,N_2754);
nand U3062 (N_3062,N_2851,N_2504);
nand U3063 (N_3063,N_2731,N_2669);
and U3064 (N_3064,N_2886,N_2711);
nor U3065 (N_3065,N_2685,N_2882);
or U3066 (N_3066,N_2583,N_2524);
and U3067 (N_3067,N_2602,N_2998);
nor U3068 (N_3068,N_2749,N_2825);
nand U3069 (N_3069,N_2910,N_2906);
and U3070 (N_3070,N_2662,N_2935);
nor U3071 (N_3071,N_2620,N_2784);
or U3072 (N_3072,N_2720,N_2960);
nor U3073 (N_3073,N_2847,N_2860);
nand U3074 (N_3074,N_2598,N_2656);
nor U3075 (N_3075,N_2975,N_2579);
nor U3076 (N_3076,N_2629,N_2695);
nor U3077 (N_3077,N_2688,N_2889);
or U3078 (N_3078,N_2661,N_2566);
or U3079 (N_3079,N_2892,N_2710);
or U3080 (N_3080,N_2525,N_2807);
nor U3081 (N_3081,N_2713,N_2943);
nor U3082 (N_3082,N_2702,N_2890);
nor U3083 (N_3083,N_2811,N_2699);
nand U3084 (N_3084,N_2655,N_2986);
nor U3085 (N_3085,N_2705,N_2876);
nand U3086 (N_3086,N_2726,N_2554);
nor U3087 (N_3087,N_2867,N_2948);
nor U3088 (N_3088,N_2919,N_2586);
or U3089 (N_3089,N_2517,N_2733);
and U3090 (N_3090,N_2622,N_2625);
nand U3091 (N_3091,N_2976,N_2870);
nand U3092 (N_3092,N_2550,N_2757);
and U3093 (N_3093,N_2966,N_2831);
and U3094 (N_3094,N_2974,N_2536);
nor U3095 (N_3095,N_2756,N_2824);
nand U3096 (N_3096,N_2574,N_2621);
or U3097 (N_3097,N_2559,N_2628);
nor U3098 (N_3098,N_2938,N_2944);
and U3099 (N_3099,N_2947,N_2985);
and U3100 (N_3100,N_2597,N_2992);
or U3101 (N_3101,N_2728,N_2727);
or U3102 (N_3102,N_2844,N_2835);
nor U3103 (N_3103,N_2848,N_2959);
nand U3104 (N_3104,N_2674,N_2610);
and U3105 (N_3105,N_2592,N_2708);
nor U3106 (N_3106,N_2562,N_2855);
nor U3107 (N_3107,N_2765,N_2603);
and U3108 (N_3108,N_2573,N_2648);
nor U3109 (N_3109,N_2893,N_2612);
nand U3110 (N_3110,N_2904,N_2866);
nor U3111 (N_3111,N_2862,N_2568);
or U3112 (N_3112,N_2836,N_2531);
nand U3113 (N_3113,N_2903,N_2972);
nand U3114 (N_3114,N_2913,N_2686);
or U3115 (N_3115,N_2917,N_2869);
and U3116 (N_3116,N_2521,N_2544);
nor U3117 (N_3117,N_2795,N_2532);
nor U3118 (N_3118,N_2678,N_2683);
and U3119 (N_3119,N_2734,N_2914);
or U3120 (N_3120,N_2874,N_2507);
nand U3121 (N_3121,N_2896,N_2671);
or U3122 (N_3122,N_2775,N_2953);
nor U3123 (N_3123,N_2526,N_2930);
nand U3124 (N_3124,N_2589,N_2508);
nand U3125 (N_3125,N_2520,N_2899);
or U3126 (N_3126,N_2883,N_2548);
nor U3127 (N_3127,N_2842,N_2799);
nor U3128 (N_3128,N_2868,N_2808);
nor U3129 (N_3129,N_2794,N_2965);
nand U3130 (N_3130,N_2514,N_2850);
nor U3131 (N_3131,N_2952,N_2778);
nor U3132 (N_3132,N_2962,N_2630);
nor U3133 (N_3133,N_2646,N_2509);
nor U3134 (N_3134,N_2822,N_2823);
nand U3135 (N_3135,N_2534,N_2796);
and U3136 (N_3136,N_2828,N_2588);
or U3137 (N_3137,N_2936,N_2582);
and U3138 (N_3138,N_2900,N_2994);
nand U3139 (N_3139,N_2764,N_2827);
or U3140 (N_3140,N_2615,N_2820);
xnor U3141 (N_3141,N_2563,N_2692);
and U3142 (N_3142,N_2701,N_2676);
nand U3143 (N_3143,N_2833,N_2929);
nand U3144 (N_3144,N_2542,N_2739);
nor U3145 (N_3145,N_2644,N_2580);
nand U3146 (N_3146,N_2555,N_2819);
nor U3147 (N_3147,N_2797,N_2601);
or U3148 (N_3148,N_2771,N_2553);
nand U3149 (N_3149,N_2716,N_2758);
and U3150 (N_3150,N_2516,N_2859);
nand U3151 (N_3151,N_2670,N_2584);
nand U3152 (N_3152,N_2991,N_2761);
nor U3153 (N_3153,N_2510,N_2638);
and U3154 (N_3154,N_2885,N_2852);
and U3155 (N_3155,N_2923,N_2746);
or U3156 (N_3156,N_2665,N_2790);
and U3157 (N_3157,N_2556,N_2755);
nand U3158 (N_3158,N_2704,N_2926);
and U3159 (N_3159,N_2712,N_2753);
and U3160 (N_3160,N_2861,N_2887);
nor U3161 (N_3161,N_2802,N_2816);
nand U3162 (N_3162,N_2637,N_2993);
nor U3163 (N_3163,N_2968,N_2715);
or U3164 (N_3164,N_2690,N_2800);
nor U3165 (N_3165,N_2768,N_2578);
and U3166 (N_3166,N_2769,N_2590);
nand U3167 (N_3167,N_2830,N_2545);
nor U3168 (N_3168,N_2838,N_2745);
or U3169 (N_3169,N_2617,N_2954);
nor U3170 (N_3170,N_2577,N_2939);
or U3171 (N_3171,N_2924,N_2570);
nand U3172 (N_3172,N_2730,N_2786);
and U3173 (N_3173,N_2604,N_2791);
or U3174 (N_3174,N_2804,N_2872);
nand U3175 (N_3175,N_2752,N_2654);
nor U3176 (N_3176,N_2680,N_2912);
and U3177 (N_3177,N_2560,N_2501);
and U3178 (N_3178,N_2787,N_2821);
or U3179 (N_3179,N_2996,N_2763);
nand U3180 (N_3180,N_2652,N_2729);
nand U3181 (N_3181,N_2522,N_2502);
nor U3182 (N_3182,N_2829,N_2718);
and U3183 (N_3183,N_2619,N_2633);
and U3184 (N_3184,N_2689,N_2709);
nor U3185 (N_3185,N_2535,N_2898);
or U3186 (N_3186,N_2832,N_2783);
and U3187 (N_3187,N_2613,N_2858);
nor U3188 (N_3188,N_2922,N_2888);
nor U3189 (N_3189,N_2905,N_2884);
nor U3190 (N_3190,N_2660,N_2901);
or U3191 (N_3191,N_2571,N_2826);
and U3192 (N_3192,N_2523,N_2666);
nand U3193 (N_3193,N_2647,N_2958);
or U3194 (N_3194,N_2609,N_2650);
and U3195 (N_3195,N_2776,N_2608);
and U3196 (N_3196,N_2782,N_2780);
nand U3197 (N_3197,N_2511,N_2817);
nand U3198 (N_3198,N_2540,N_2684);
or U3199 (N_3199,N_2691,N_2505);
xnor U3200 (N_3200,N_2611,N_2607);
nor U3201 (N_3201,N_2932,N_2977);
or U3202 (N_3202,N_2663,N_2909);
nor U3203 (N_3203,N_2879,N_2631);
nor U3204 (N_3204,N_2694,N_2547);
nand U3205 (N_3205,N_2940,N_2785);
and U3206 (N_3206,N_2561,N_2856);
nand U3207 (N_3207,N_2810,N_2970);
nor U3208 (N_3208,N_2675,N_2668);
nand U3209 (N_3209,N_2957,N_2732);
or U3210 (N_3210,N_2649,N_2738);
nor U3211 (N_3211,N_2818,N_2635);
or U3212 (N_3212,N_2854,N_2719);
nand U3213 (N_3213,N_2865,N_2814);
nor U3214 (N_3214,N_2537,N_2788);
or U3215 (N_3215,N_2575,N_2697);
nand U3216 (N_3216,N_2645,N_2594);
nand U3217 (N_3217,N_2533,N_2627);
nor U3218 (N_3218,N_2651,N_2750);
nor U3219 (N_3219,N_2949,N_2760);
nand U3220 (N_3220,N_2894,N_2961);
nand U3221 (N_3221,N_2682,N_2529);
or U3222 (N_3222,N_2634,N_2596);
nor U3223 (N_3223,N_2971,N_2664);
and U3224 (N_3224,N_2837,N_2840);
nand U3225 (N_3225,N_2916,N_2721);
nand U3226 (N_3226,N_2576,N_2541);
nand U3227 (N_3227,N_2693,N_2538);
nand U3228 (N_3228,N_2677,N_2955);
or U3229 (N_3229,N_2643,N_2969);
or U3230 (N_3230,N_2687,N_2864);
and U3231 (N_3231,N_2659,N_2744);
nor U3232 (N_3232,N_2963,N_2519);
and U3233 (N_3233,N_2747,N_2740);
nor U3234 (N_3234,N_2878,N_2552);
nor U3235 (N_3235,N_2841,N_2920);
nand U3236 (N_3236,N_2640,N_2572);
or U3237 (N_3237,N_2614,N_2527);
nand U3238 (N_3238,N_2946,N_2737);
nand U3239 (N_3239,N_2672,N_2557);
and U3240 (N_3240,N_2639,N_2945);
or U3241 (N_3241,N_2871,N_2698);
nand U3242 (N_3242,N_2513,N_2997);
and U3243 (N_3243,N_2964,N_2863);
and U3244 (N_3244,N_2585,N_2902);
and U3245 (N_3245,N_2979,N_2626);
and U3246 (N_3246,N_2931,N_2983);
nor U3247 (N_3247,N_2941,N_2928);
nor U3248 (N_3248,N_2748,N_2706);
and U3249 (N_3249,N_2911,N_2897);
and U3250 (N_3250,N_2843,N_2504);
nor U3251 (N_3251,N_2876,N_2958);
nand U3252 (N_3252,N_2845,N_2886);
or U3253 (N_3253,N_2609,N_2542);
nor U3254 (N_3254,N_2719,N_2532);
and U3255 (N_3255,N_2513,N_2634);
nor U3256 (N_3256,N_2546,N_2910);
nor U3257 (N_3257,N_2552,N_2834);
and U3258 (N_3258,N_2779,N_2789);
nand U3259 (N_3259,N_2859,N_2993);
xnor U3260 (N_3260,N_2524,N_2718);
and U3261 (N_3261,N_2509,N_2839);
or U3262 (N_3262,N_2661,N_2739);
or U3263 (N_3263,N_2526,N_2680);
nor U3264 (N_3264,N_2500,N_2771);
nand U3265 (N_3265,N_2975,N_2956);
nor U3266 (N_3266,N_2723,N_2558);
nand U3267 (N_3267,N_2643,N_2673);
or U3268 (N_3268,N_2919,N_2708);
or U3269 (N_3269,N_2697,N_2905);
nor U3270 (N_3270,N_2659,N_2818);
nor U3271 (N_3271,N_2710,N_2970);
and U3272 (N_3272,N_2811,N_2760);
nand U3273 (N_3273,N_2806,N_2975);
nor U3274 (N_3274,N_2902,N_2816);
and U3275 (N_3275,N_2850,N_2810);
nand U3276 (N_3276,N_2810,N_2701);
or U3277 (N_3277,N_2750,N_2830);
nor U3278 (N_3278,N_2914,N_2731);
nand U3279 (N_3279,N_2631,N_2934);
nand U3280 (N_3280,N_2652,N_2539);
nand U3281 (N_3281,N_2677,N_2556);
nor U3282 (N_3282,N_2770,N_2695);
or U3283 (N_3283,N_2854,N_2844);
and U3284 (N_3284,N_2871,N_2790);
and U3285 (N_3285,N_2862,N_2587);
or U3286 (N_3286,N_2923,N_2879);
nor U3287 (N_3287,N_2840,N_2666);
nand U3288 (N_3288,N_2697,N_2929);
or U3289 (N_3289,N_2735,N_2551);
nor U3290 (N_3290,N_2776,N_2793);
nand U3291 (N_3291,N_2869,N_2719);
and U3292 (N_3292,N_2763,N_2927);
or U3293 (N_3293,N_2622,N_2736);
and U3294 (N_3294,N_2885,N_2778);
nand U3295 (N_3295,N_2621,N_2888);
nor U3296 (N_3296,N_2798,N_2841);
nand U3297 (N_3297,N_2734,N_2547);
and U3298 (N_3298,N_2673,N_2692);
nor U3299 (N_3299,N_2859,N_2550);
and U3300 (N_3300,N_2916,N_2637);
or U3301 (N_3301,N_2711,N_2945);
and U3302 (N_3302,N_2986,N_2522);
nand U3303 (N_3303,N_2541,N_2619);
nor U3304 (N_3304,N_2597,N_2583);
and U3305 (N_3305,N_2644,N_2754);
xor U3306 (N_3306,N_2869,N_2563);
and U3307 (N_3307,N_2557,N_2902);
nor U3308 (N_3308,N_2627,N_2820);
nand U3309 (N_3309,N_2569,N_2906);
and U3310 (N_3310,N_2624,N_2741);
and U3311 (N_3311,N_2790,N_2632);
nand U3312 (N_3312,N_2558,N_2535);
and U3313 (N_3313,N_2883,N_2788);
and U3314 (N_3314,N_2918,N_2692);
or U3315 (N_3315,N_2704,N_2539);
nor U3316 (N_3316,N_2803,N_2942);
and U3317 (N_3317,N_2912,N_2941);
nor U3318 (N_3318,N_2526,N_2802);
nor U3319 (N_3319,N_2644,N_2708);
nand U3320 (N_3320,N_2920,N_2759);
nand U3321 (N_3321,N_2507,N_2960);
or U3322 (N_3322,N_2915,N_2789);
nand U3323 (N_3323,N_2602,N_2973);
or U3324 (N_3324,N_2551,N_2874);
xor U3325 (N_3325,N_2864,N_2921);
or U3326 (N_3326,N_2700,N_2776);
nor U3327 (N_3327,N_2505,N_2650);
nand U3328 (N_3328,N_2650,N_2923);
nor U3329 (N_3329,N_2902,N_2653);
nand U3330 (N_3330,N_2531,N_2737);
or U3331 (N_3331,N_2721,N_2963);
nand U3332 (N_3332,N_2529,N_2873);
or U3333 (N_3333,N_2683,N_2583);
or U3334 (N_3334,N_2791,N_2833);
and U3335 (N_3335,N_2605,N_2896);
xnor U3336 (N_3336,N_2852,N_2997);
and U3337 (N_3337,N_2962,N_2755);
nor U3338 (N_3338,N_2712,N_2574);
nand U3339 (N_3339,N_2970,N_2697);
nand U3340 (N_3340,N_2865,N_2821);
nor U3341 (N_3341,N_2545,N_2778);
nand U3342 (N_3342,N_2870,N_2589);
or U3343 (N_3343,N_2978,N_2626);
nand U3344 (N_3344,N_2532,N_2605);
nor U3345 (N_3345,N_2784,N_2762);
and U3346 (N_3346,N_2886,N_2597);
nand U3347 (N_3347,N_2937,N_2521);
nor U3348 (N_3348,N_2858,N_2893);
or U3349 (N_3349,N_2768,N_2749);
nor U3350 (N_3350,N_2750,N_2650);
or U3351 (N_3351,N_2944,N_2530);
and U3352 (N_3352,N_2538,N_2999);
and U3353 (N_3353,N_2623,N_2869);
nand U3354 (N_3354,N_2838,N_2916);
nand U3355 (N_3355,N_2534,N_2639);
nor U3356 (N_3356,N_2598,N_2801);
nand U3357 (N_3357,N_2745,N_2974);
nand U3358 (N_3358,N_2677,N_2702);
and U3359 (N_3359,N_2716,N_2936);
nor U3360 (N_3360,N_2505,N_2525);
nand U3361 (N_3361,N_2926,N_2728);
nand U3362 (N_3362,N_2791,N_2709);
nand U3363 (N_3363,N_2748,N_2941);
or U3364 (N_3364,N_2892,N_2689);
nor U3365 (N_3365,N_2990,N_2584);
and U3366 (N_3366,N_2959,N_2987);
and U3367 (N_3367,N_2963,N_2930);
and U3368 (N_3368,N_2753,N_2863);
and U3369 (N_3369,N_2802,N_2984);
nand U3370 (N_3370,N_2992,N_2658);
nor U3371 (N_3371,N_2559,N_2720);
nand U3372 (N_3372,N_2532,N_2791);
and U3373 (N_3373,N_2831,N_2708);
nor U3374 (N_3374,N_2571,N_2650);
nor U3375 (N_3375,N_2665,N_2956);
and U3376 (N_3376,N_2838,N_2728);
and U3377 (N_3377,N_2586,N_2811);
nor U3378 (N_3378,N_2656,N_2906);
and U3379 (N_3379,N_2567,N_2781);
or U3380 (N_3380,N_2529,N_2616);
xnor U3381 (N_3381,N_2537,N_2833);
nor U3382 (N_3382,N_2946,N_2928);
nor U3383 (N_3383,N_2585,N_2921);
nor U3384 (N_3384,N_2790,N_2751);
xor U3385 (N_3385,N_2861,N_2754);
and U3386 (N_3386,N_2520,N_2815);
nand U3387 (N_3387,N_2602,N_2864);
and U3388 (N_3388,N_2813,N_2576);
nand U3389 (N_3389,N_2981,N_2550);
or U3390 (N_3390,N_2888,N_2826);
or U3391 (N_3391,N_2990,N_2917);
nor U3392 (N_3392,N_2969,N_2537);
and U3393 (N_3393,N_2524,N_2622);
nor U3394 (N_3394,N_2763,N_2938);
nor U3395 (N_3395,N_2822,N_2573);
or U3396 (N_3396,N_2541,N_2819);
nor U3397 (N_3397,N_2553,N_2852);
or U3398 (N_3398,N_2660,N_2526);
nand U3399 (N_3399,N_2660,N_2930);
nor U3400 (N_3400,N_2641,N_2919);
nor U3401 (N_3401,N_2880,N_2951);
or U3402 (N_3402,N_2915,N_2701);
nand U3403 (N_3403,N_2906,N_2592);
nor U3404 (N_3404,N_2740,N_2505);
or U3405 (N_3405,N_2861,N_2725);
nor U3406 (N_3406,N_2768,N_2914);
nor U3407 (N_3407,N_2928,N_2959);
nor U3408 (N_3408,N_2711,N_2547);
or U3409 (N_3409,N_2792,N_2515);
or U3410 (N_3410,N_2844,N_2895);
or U3411 (N_3411,N_2814,N_2640);
or U3412 (N_3412,N_2681,N_2596);
or U3413 (N_3413,N_2979,N_2840);
or U3414 (N_3414,N_2829,N_2623);
nand U3415 (N_3415,N_2523,N_2887);
or U3416 (N_3416,N_2969,N_2928);
nor U3417 (N_3417,N_2810,N_2988);
or U3418 (N_3418,N_2836,N_2890);
or U3419 (N_3419,N_2500,N_2813);
nand U3420 (N_3420,N_2670,N_2774);
or U3421 (N_3421,N_2651,N_2834);
nor U3422 (N_3422,N_2632,N_2566);
nand U3423 (N_3423,N_2606,N_2916);
and U3424 (N_3424,N_2597,N_2767);
and U3425 (N_3425,N_2835,N_2841);
nor U3426 (N_3426,N_2609,N_2820);
and U3427 (N_3427,N_2947,N_2829);
or U3428 (N_3428,N_2662,N_2789);
nor U3429 (N_3429,N_2882,N_2872);
or U3430 (N_3430,N_2917,N_2691);
and U3431 (N_3431,N_2827,N_2619);
and U3432 (N_3432,N_2501,N_2847);
nand U3433 (N_3433,N_2553,N_2528);
and U3434 (N_3434,N_2722,N_2501);
or U3435 (N_3435,N_2951,N_2822);
nor U3436 (N_3436,N_2739,N_2818);
nor U3437 (N_3437,N_2730,N_2691);
nor U3438 (N_3438,N_2989,N_2761);
nor U3439 (N_3439,N_2845,N_2566);
nand U3440 (N_3440,N_2810,N_2962);
and U3441 (N_3441,N_2769,N_2616);
and U3442 (N_3442,N_2788,N_2735);
nor U3443 (N_3443,N_2764,N_2728);
nand U3444 (N_3444,N_2863,N_2736);
nor U3445 (N_3445,N_2675,N_2795);
nor U3446 (N_3446,N_2984,N_2711);
or U3447 (N_3447,N_2903,N_2728);
and U3448 (N_3448,N_2630,N_2610);
nand U3449 (N_3449,N_2812,N_2511);
and U3450 (N_3450,N_2974,N_2659);
or U3451 (N_3451,N_2579,N_2878);
nor U3452 (N_3452,N_2726,N_2638);
and U3453 (N_3453,N_2558,N_2510);
or U3454 (N_3454,N_2501,N_2574);
or U3455 (N_3455,N_2959,N_2811);
nand U3456 (N_3456,N_2799,N_2722);
nand U3457 (N_3457,N_2791,N_2522);
and U3458 (N_3458,N_2838,N_2507);
and U3459 (N_3459,N_2773,N_2568);
nand U3460 (N_3460,N_2629,N_2836);
nor U3461 (N_3461,N_2531,N_2948);
nor U3462 (N_3462,N_2647,N_2577);
nor U3463 (N_3463,N_2885,N_2569);
xnor U3464 (N_3464,N_2950,N_2658);
or U3465 (N_3465,N_2881,N_2950);
or U3466 (N_3466,N_2914,N_2520);
and U3467 (N_3467,N_2503,N_2781);
and U3468 (N_3468,N_2780,N_2924);
nor U3469 (N_3469,N_2568,N_2671);
and U3470 (N_3470,N_2925,N_2586);
nor U3471 (N_3471,N_2859,N_2621);
nand U3472 (N_3472,N_2859,N_2737);
or U3473 (N_3473,N_2957,N_2986);
nor U3474 (N_3474,N_2951,N_2744);
or U3475 (N_3475,N_2937,N_2684);
and U3476 (N_3476,N_2514,N_2565);
nor U3477 (N_3477,N_2777,N_2848);
or U3478 (N_3478,N_2786,N_2679);
nor U3479 (N_3479,N_2588,N_2652);
nor U3480 (N_3480,N_2892,N_2772);
nor U3481 (N_3481,N_2745,N_2687);
and U3482 (N_3482,N_2925,N_2829);
nor U3483 (N_3483,N_2832,N_2556);
nor U3484 (N_3484,N_2691,N_2668);
and U3485 (N_3485,N_2890,N_2804);
nor U3486 (N_3486,N_2563,N_2688);
nor U3487 (N_3487,N_2843,N_2933);
nand U3488 (N_3488,N_2981,N_2582);
and U3489 (N_3489,N_2766,N_2919);
nor U3490 (N_3490,N_2634,N_2784);
nor U3491 (N_3491,N_2583,N_2908);
nand U3492 (N_3492,N_2667,N_2731);
or U3493 (N_3493,N_2990,N_2513);
nor U3494 (N_3494,N_2558,N_2934);
or U3495 (N_3495,N_2606,N_2805);
nand U3496 (N_3496,N_2819,N_2691);
and U3497 (N_3497,N_2830,N_2564);
and U3498 (N_3498,N_2511,N_2663);
nor U3499 (N_3499,N_2541,N_2639);
nand U3500 (N_3500,N_3049,N_3270);
and U3501 (N_3501,N_3114,N_3120);
and U3502 (N_3502,N_3147,N_3258);
nor U3503 (N_3503,N_3362,N_3444);
nor U3504 (N_3504,N_3351,N_3212);
nor U3505 (N_3505,N_3411,N_3467);
and U3506 (N_3506,N_3405,N_3034);
nand U3507 (N_3507,N_3140,N_3245);
nor U3508 (N_3508,N_3051,N_3456);
nor U3509 (N_3509,N_3307,N_3356);
xnor U3510 (N_3510,N_3058,N_3075);
or U3511 (N_3511,N_3230,N_3018);
xnor U3512 (N_3512,N_3243,N_3095);
nor U3513 (N_3513,N_3195,N_3072);
or U3514 (N_3514,N_3478,N_3129);
nor U3515 (N_3515,N_3443,N_3479);
nand U3516 (N_3516,N_3215,N_3182);
nor U3517 (N_3517,N_3224,N_3176);
nand U3518 (N_3518,N_3241,N_3311);
or U3519 (N_3519,N_3400,N_3488);
nand U3520 (N_3520,N_3396,N_3015);
and U3521 (N_3521,N_3021,N_3343);
nor U3522 (N_3522,N_3056,N_3216);
and U3523 (N_3523,N_3206,N_3229);
nor U3524 (N_3524,N_3457,N_3030);
nor U3525 (N_3525,N_3221,N_3352);
and U3526 (N_3526,N_3069,N_3361);
or U3527 (N_3527,N_3165,N_3298);
nand U3528 (N_3528,N_3103,N_3225);
or U3529 (N_3529,N_3177,N_3117);
nand U3530 (N_3530,N_3432,N_3135);
nand U3531 (N_3531,N_3438,N_3346);
nand U3532 (N_3532,N_3272,N_3423);
nor U3533 (N_3533,N_3308,N_3223);
or U3534 (N_3534,N_3257,N_3242);
and U3535 (N_3535,N_3252,N_3286);
and U3536 (N_3536,N_3306,N_3294);
and U3537 (N_3537,N_3116,N_3374);
nor U3538 (N_3538,N_3439,N_3373);
and U3539 (N_3539,N_3131,N_3145);
nor U3540 (N_3540,N_3290,N_3202);
and U3541 (N_3541,N_3259,N_3050);
or U3542 (N_3542,N_3434,N_3435);
and U3543 (N_3543,N_3424,N_3480);
nand U3544 (N_3544,N_3265,N_3020);
nor U3545 (N_3545,N_3084,N_3204);
nor U3546 (N_3546,N_3172,N_3232);
and U3547 (N_3547,N_3275,N_3149);
and U3548 (N_3548,N_3261,N_3217);
nand U3549 (N_3549,N_3345,N_3474);
nand U3550 (N_3550,N_3440,N_3137);
nor U3551 (N_3551,N_3236,N_3445);
nor U3552 (N_3552,N_3318,N_3200);
and U3553 (N_3553,N_3295,N_3039);
and U3554 (N_3554,N_3074,N_3162);
or U3555 (N_3555,N_3151,N_3323);
nand U3556 (N_3556,N_3452,N_3004);
nand U3557 (N_3557,N_3128,N_3062);
nand U3558 (N_3558,N_3139,N_3080);
nand U3559 (N_3559,N_3322,N_3031);
or U3560 (N_3560,N_3477,N_3130);
or U3561 (N_3561,N_3449,N_3256);
and U3562 (N_3562,N_3010,N_3313);
or U3563 (N_3563,N_3088,N_3040);
and U3564 (N_3564,N_3150,N_3384);
or U3565 (N_3565,N_3025,N_3155);
nand U3566 (N_3566,N_3187,N_3238);
nor U3567 (N_3567,N_3097,N_3002);
and U3568 (N_3568,N_3099,N_3142);
or U3569 (N_3569,N_3170,N_3458);
nor U3570 (N_3570,N_3174,N_3027);
or U3571 (N_3571,N_3016,N_3262);
or U3572 (N_3572,N_3093,N_3017);
nand U3573 (N_3573,N_3285,N_3302);
nor U3574 (N_3574,N_3353,N_3124);
and U3575 (N_3575,N_3363,N_3032);
nand U3576 (N_3576,N_3317,N_3288);
or U3577 (N_3577,N_3268,N_3481);
and U3578 (N_3578,N_3381,N_3102);
nand U3579 (N_3579,N_3462,N_3240);
and U3580 (N_3580,N_3448,N_3047);
and U3581 (N_3581,N_3246,N_3420);
nand U3582 (N_3582,N_3186,N_3418);
nand U3583 (N_3583,N_3293,N_3070);
nor U3584 (N_3584,N_3184,N_3447);
nor U3585 (N_3585,N_3228,N_3159);
nand U3586 (N_3586,N_3278,N_3372);
and U3587 (N_3587,N_3086,N_3408);
or U3588 (N_3588,N_3210,N_3327);
nor U3589 (N_3589,N_3104,N_3334);
nor U3590 (N_3590,N_3158,N_3161);
and U3591 (N_3591,N_3416,N_3003);
and U3592 (N_3592,N_3152,N_3496);
and U3593 (N_3593,N_3013,N_3377);
nor U3594 (N_3594,N_3109,N_3183);
nor U3595 (N_3595,N_3297,N_3375);
nor U3596 (N_3596,N_3329,N_3348);
and U3597 (N_3597,N_3430,N_3365);
nand U3598 (N_3598,N_3284,N_3391);
or U3599 (N_3599,N_3341,N_3105);
or U3600 (N_3600,N_3055,N_3407);
and U3601 (N_3601,N_3271,N_3185);
nor U3602 (N_3602,N_3357,N_3154);
or U3603 (N_3603,N_3392,N_3083);
and U3604 (N_3604,N_3024,N_3390);
nand U3605 (N_3605,N_3226,N_3429);
nor U3606 (N_3606,N_3280,N_3468);
and U3607 (N_3607,N_3332,N_3368);
nor U3608 (N_3608,N_3376,N_3325);
or U3609 (N_3609,N_3469,N_3219);
xor U3610 (N_3610,N_3354,N_3442);
and U3611 (N_3611,N_3132,N_3495);
or U3612 (N_3612,N_3211,N_3493);
or U3613 (N_3613,N_3143,N_3157);
or U3614 (N_3614,N_3235,N_3399);
and U3615 (N_3615,N_3193,N_3299);
nor U3616 (N_3616,N_3309,N_3173);
nor U3617 (N_3617,N_3009,N_3492);
or U3618 (N_3618,N_3045,N_3199);
nand U3619 (N_3619,N_3388,N_3196);
and U3620 (N_3620,N_3037,N_3414);
and U3621 (N_3621,N_3061,N_3378);
or U3622 (N_3622,N_3036,N_3310);
xor U3623 (N_3623,N_3498,N_3483);
nand U3624 (N_3624,N_3119,N_3098);
or U3625 (N_3625,N_3121,N_3059);
nor U3626 (N_3626,N_3472,N_3427);
nor U3627 (N_3627,N_3274,N_3181);
and U3628 (N_3628,N_3428,N_3335);
and U3629 (N_3629,N_3136,N_3266);
nand U3630 (N_3630,N_3324,N_3071);
or U3631 (N_3631,N_3042,N_3019);
or U3632 (N_3632,N_3475,N_3291);
nand U3633 (N_3633,N_3389,N_3250);
nor U3634 (N_3634,N_3450,N_3222);
and U3635 (N_3635,N_3277,N_3383);
or U3636 (N_3636,N_3328,N_3404);
and U3637 (N_3637,N_3461,N_3022);
nand U3638 (N_3638,N_3422,N_3198);
nand U3639 (N_3639,N_3330,N_3459);
nand U3640 (N_3640,N_3041,N_3484);
and U3641 (N_3641,N_3100,N_3491);
nor U3642 (N_3642,N_3292,N_3369);
or U3643 (N_3643,N_3350,N_3436);
and U3644 (N_3644,N_3048,N_3397);
nor U3645 (N_3645,N_3126,N_3141);
or U3646 (N_3646,N_3453,N_3044);
and U3647 (N_3647,N_3065,N_3092);
and U3648 (N_3648,N_3296,N_3340);
and U3649 (N_3649,N_3090,N_3267);
nand U3650 (N_3650,N_3473,N_3276);
nor U3651 (N_3651,N_3494,N_3054);
and U3652 (N_3652,N_3251,N_3077);
nor U3653 (N_3653,N_3387,N_3007);
nand U3654 (N_3654,N_3209,N_3189);
or U3655 (N_3655,N_3180,N_3314);
or U3656 (N_3656,N_3413,N_3033);
and U3657 (N_3657,N_3487,N_3499);
or U3658 (N_3658,N_3273,N_3412);
and U3659 (N_3659,N_3426,N_3067);
or U3660 (N_3660,N_3066,N_3089);
nor U3661 (N_3661,N_3455,N_3106);
or U3662 (N_3662,N_3281,N_3260);
or U3663 (N_3663,N_3360,N_3153);
nand U3664 (N_3664,N_3289,N_3192);
nand U3665 (N_3665,N_3227,N_3344);
xor U3666 (N_3666,N_3207,N_3421);
nor U3667 (N_3667,N_3111,N_3085);
nor U3668 (N_3668,N_3108,N_3203);
or U3669 (N_3669,N_3094,N_3486);
nor U3670 (N_3670,N_3367,N_3433);
nor U3671 (N_3671,N_3029,N_3073);
and U3672 (N_3672,N_3415,N_3220);
and U3673 (N_3673,N_3167,N_3255);
and U3674 (N_3674,N_3485,N_3336);
nor U3675 (N_3675,N_3023,N_3213);
and U3676 (N_3676,N_3287,N_3454);
and U3677 (N_3677,N_3446,N_3038);
nand U3678 (N_3678,N_3078,N_3026);
nor U3679 (N_3679,N_3464,N_3279);
nor U3680 (N_3680,N_3057,N_3282);
or U3681 (N_3681,N_3338,N_3122);
and U3682 (N_3682,N_3382,N_3239);
nor U3683 (N_3683,N_3133,N_3466);
nand U3684 (N_3684,N_3028,N_3315);
nand U3685 (N_3685,N_3231,N_3123);
nor U3686 (N_3686,N_3410,N_3096);
or U3687 (N_3687,N_3403,N_3208);
and U3688 (N_3688,N_3014,N_3398);
nor U3689 (N_3689,N_3333,N_3321);
and U3690 (N_3690,N_3197,N_3248);
or U3691 (N_3691,N_3385,N_3342);
or U3692 (N_3692,N_3043,N_3355);
nand U3693 (N_3693,N_3076,N_3303);
or U3694 (N_3694,N_3006,N_3393);
and U3695 (N_3695,N_3247,N_3316);
or U3696 (N_3696,N_3087,N_3349);
and U3697 (N_3697,N_3409,N_3264);
nand U3698 (N_3698,N_3146,N_3451);
nand U3699 (N_3699,N_3359,N_3402);
or U3700 (N_3700,N_3001,N_3068);
and U3701 (N_3701,N_3079,N_3425);
nand U3702 (N_3702,N_3138,N_3441);
or U3703 (N_3703,N_3320,N_3134);
or U3704 (N_3704,N_3371,N_3331);
or U3705 (N_3705,N_3091,N_3263);
nand U3706 (N_3706,N_3107,N_3489);
nand U3707 (N_3707,N_3304,N_3237);
or U3708 (N_3708,N_3326,N_3300);
and U3709 (N_3709,N_3319,N_3156);
or U3710 (N_3710,N_3012,N_3190);
nand U3711 (N_3711,N_3188,N_3000);
or U3712 (N_3712,N_3253,N_3490);
and U3713 (N_3713,N_3301,N_3171);
nor U3714 (N_3714,N_3234,N_3118);
nor U3715 (N_3715,N_3347,N_3148);
nand U3716 (N_3716,N_3166,N_3005);
or U3717 (N_3717,N_3125,N_3179);
and U3718 (N_3718,N_3339,N_3312);
and U3719 (N_3719,N_3431,N_3366);
nand U3720 (N_3720,N_3110,N_3233);
or U3721 (N_3721,N_3364,N_3470);
or U3722 (N_3722,N_3194,N_3254);
nor U3723 (N_3723,N_3283,N_3115);
and U3724 (N_3724,N_3249,N_3380);
nor U3725 (N_3725,N_3163,N_3386);
nand U3726 (N_3726,N_3463,N_3417);
and U3727 (N_3727,N_3060,N_3437);
and U3728 (N_3728,N_3064,N_3218);
or U3729 (N_3729,N_3214,N_3305);
nor U3730 (N_3730,N_3337,N_3011);
or U3731 (N_3731,N_3160,N_3175);
or U3732 (N_3732,N_3112,N_3035);
and U3733 (N_3733,N_3113,N_3370);
xor U3734 (N_3734,N_3465,N_3379);
nand U3735 (N_3735,N_3191,N_3053);
nor U3736 (N_3736,N_3244,N_3205);
or U3737 (N_3737,N_3144,N_3497);
or U3738 (N_3738,N_3482,N_3052);
or U3739 (N_3739,N_3471,N_3101);
or U3740 (N_3740,N_3394,N_3081);
or U3741 (N_3741,N_3164,N_3476);
nand U3742 (N_3742,N_3201,N_3169);
and U3743 (N_3743,N_3082,N_3460);
nand U3744 (N_3744,N_3419,N_3008);
or U3745 (N_3745,N_3178,N_3046);
and U3746 (N_3746,N_3168,N_3269);
or U3747 (N_3747,N_3127,N_3401);
nand U3748 (N_3748,N_3358,N_3063);
or U3749 (N_3749,N_3406,N_3395);
nor U3750 (N_3750,N_3467,N_3348);
or U3751 (N_3751,N_3189,N_3434);
nand U3752 (N_3752,N_3253,N_3405);
and U3753 (N_3753,N_3152,N_3196);
nand U3754 (N_3754,N_3054,N_3106);
or U3755 (N_3755,N_3076,N_3185);
nor U3756 (N_3756,N_3058,N_3055);
nand U3757 (N_3757,N_3051,N_3383);
or U3758 (N_3758,N_3412,N_3310);
nand U3759 (N_3759,N_3329,N_3386);
nand U3760 (N_3760,N_3142,N_3202);
nand U3761 (N_3761,N_3013,N_3104);
nand U3762 (N_3762,N_3474,N_3333);
nand U3763 (N_3763,N_3095,N_3323);
nand U3764 (N_3764,N_3007,N_3050);
nor U3765 (N_3765,N_3208,N_3419);
nand U3766 (N_3766,N_3431,N_3343);
nand U3767 (N_3767,N_3255,N_3036);
nor U3768 (N_3768,N_3016,N_3142);
nor U3769 (N_3769,N_3050,N_3112);
or U3770 (N_3770,N_3442,N_3135);
or U3771 (N_3771,N_3392,N_3498);
nand U3772 (N_3772,N_3409,N_3460);
and U3773 (N_3773,N_3009,N_3233);
or U3774 (N_3774,N_3026,N_3050);
or U3775 (N_3775,N_3206,N_3126);
nand U3776 (N_3776,N_3025,N_3115);
nor U3777 (N_3777,N_3317,N_3083);
nand U3778 (N_3778,N_3467,N_3341);
nand U3779 (N_3779,N_3241,N_3039);
nor U3780 (N_3780,N_3125,N_3335);
or U3781 (N_3781,N_3069,N_3024);
nor U3782 (N_3782,N_3308,N_3325);
nor U3783 (N_3783,N_3053,N_3242);
nor U3784 (N_3784,N_3155,N_3014);
nand U3785 (N_3785,N_3430,N_3134);
nor U3786 (N_3786,N_3256,N_3216);
or U3787 (N_3787,N_3070,N_3296);
or U3788 (N_3788,N_3106,N_3434);
and U3789 (N_3789,N_3001,N_3373);
nand U3790 (N_3790,N_3445,N_3273);
nor U3791 (N_3791,N_3291,N_3223);
or U3792 (N_3792,N_3095,N_3322);
and U3793 (N_3793,N_3376,N_3193);
or U3794 (N_3794,N_3413,N_3153);
or U3795 (N_3795,N_3349,N_3146);
or U3796 (N_3796,N_3148,N_3054);
and U3797 (N_3797,N_3397,N_3092);
nor U3798 (N_3798,N_3252,N_3247);
nor U3799 (N_3799,N_3487,N_3174);
nand U3800 (N_3800,N_3029,N_3472);
and U3801 (N_3801,N_3199,N_3346);
or U3802 (N_3802,N_3132,N_3383);
nor U3803 (N_3803,N_3239,N_3437);
and U3804 (N_3804,N_3154,N_3352);
and U3805 (N_3805,N_3286,N_3308);
and U3806 (N_3806,N_3299,N_3321);
or U3807 (N_3807,N_3109,N_3259);
nor U3808 (N_3808,N_3080,N_3199);
and U3809 (N_3809,N_3317,N_3460);
and U3810 (N_3810,N_3349,N_3214);
and U3811 (N_3811,N_3210,N_3371);
and U3812 (N_3812,N_3445,N_3440);
or U3813 (N_3813,N_3210,N_3025);
and U3814 (N_3814,N_3081,N_3241);
and U3815 (N_3815,N_3350,N_3154);
or U3816 (N_3816,N_3220,N_3109);
and U3817 (N_3817,N_3395,N_3051);
nor U3818 (N_3818,N_3236,N_3402);
nand U3819 (N_3819,N_3067,N_3366);
nor U3820 (N_3820,N_3039,N_3037);
and U3821 (N_3821,N_3369,N_3035);
xor U3822 (N_3822,N_3174,N_3108);
or U3823 (N_3823,N_3095,N_3173);
or U3824 (N_3824,N_3174,N_3194);
and U3825 (N_3825,N_3332,N_3127);
or U3826 (N_3826,N_3060,N_3046);
and U3827 (N_3827,N_3381,N_3045);
or U3828 (N_3828,N_3067,N_3186);
and U3829 (N_3829,N_3214,N_3006);
or U3830 (N_3830,N_3107,N_3167);
nand U3831 (N_3831,N_3006,N_3364);
nand U3832 (N_3832,N_3053,N_3238);
nor U3833 (N_3833,N_3191,N_3483);
nand U3834 (N_3834,N_3332,N_3135);
and U3835 (N_3835,N_3449,N_3060);
nand U3836 (N_3836,N_3149,N_3182);
nor U3837 (N_3837,N_3221,N_3032);
and U3838 (N_3838,N_3356,N_3202);
nand U3839 (N_3839,N_3268,N_3429);
nand U3840 (N_3840,N_3405,N_3019);
or U3841 (N_3841,N_3181,N_3164);
nand U3842 (N_3842,N_3149,N_3018);
or U3843 (N_3843,N_3082,N_3011);
nand U3844 (N_3844,N_3225,N_3387);
or U3845 (N_3845,N_3153,N_3117);
or U3846 (N_3846,N_3174,N_3266);
nor U3847 (N_3847,N_3202,N_3383);
and U3848 (N_3848,N_3008,N_3262);
or U3849 (N_3849,N_3188,N_3022);
nand U3850 (N_3850,N_3252,N_3330);
nor U3851 (N_3851,N_3280,N_3021);
or U3852 (N_3852,N_3191,N_3095);
or U3853 (N_3853,N_3441,N_3167);
nor U3854 (N_3854,N_3399,N_3107);
nor U3855 (N_3855,N_3492,N_3053);
and U3856 (N_3856,N_3473,N_3235);
and U3857 (N_3857,N_3179,N_3361);
nand U3858 (N_3858,N_3480,N_3361);
nand U3859 (N_3859,N_3005,N_3135);
and U3860 (N_3860,N_3411,N_3196);
nor U3861 (N_3861,N_3441,N_3208);
and U3862 (N_3862,N_3306,N_3136);
or U3863 (N_3863,N_3126,N_3106);
or U3864 (N_3864,N_3087,N_3402);
nor U3865 (N_3865,N_3073,N_3288);
nand U3866 (N_3866,N_3323,N_3297);
nand U3867 (N_3867,N_3324,N_3040);
nor U3868 (N_3868,N_3049,N_3314);
and U3869 (N_3869,N_3406,N_3392);
nor U3870 (N_3870,N_3318,N_3467);
and U3871 (N_3871,N_3149,N_3185);
and U3872 (N_3872,N_3346,N_3404);
nand U3873 (N_3873,N_3017,N_3248);
and U3874 (N_3874,N_3308,N_3270);
or U3875 (N_3875,N_3276,N_3394);
and U3876 (N_3876,N_3097,N_3106);
nand U3877 (N_3877,N_3098,N_3006);
nor U3878 (N_3878,N_3341,N_3457);
or U3879 (N_3879,N_3207,N_3081);
and U3880 (N_3880,N_3317,N_3428);
and U3881 (N_3881,N_3298,N_3282);
nor U3882 (N_3882,N_3305,N_3464);
nand U3883 (N_3883,N_3415,N_3393);
nor U3884 (N_3884,N_3327,N_3154);
and U3885 (N_3885,N_3353,N_3369);
or U3886 (N_3886,N_3388,N_3099);
nor U3887 (N_3887,N_3178,N_3064);
and U3888 (N_3888,N_3024,N_3063);
or U3889 (N_3889,N_3466,N_3422);
nand U3890 (N_3890,N_3232,N_3057);
nand U3891 (N_3891,N_3376,N_3471);
and U3892 (N_3892,N_3199,N_3284);
and U3893 (N_3893,N_3147,N_3189);
and U3894 (N_3894,N_3040,N_3458);
and U3895 (N_3895,N_3449,N_3498);
and U3896 (N_3896,N_3008,N_3045);
or U3897 (N_3897,N_3424,N_3190);
xnor U3898 (N_3898,N_3192,N_3256);
and U3899 (N_3899,N_3435,N_3012);
or U3900 (N_3900,N_3447,N_3219);
or U3901 (N_3901,N_3245,N_3369);
nor U3902 (N_3902,N_3058,N_3354);
nand U3903 (N_3903,N_3192,N_3175);
or U3904 (N_3904,N_3074,N_3313);
or U3905 (N_3905,N_3283,N_3175);
or U3906 (N_3906,N_3075,N_3378);
and U3907 (N_3907,N_3437,N_3333);
or U3908 (N_3908,N_3437,N_3349);
nand U3909 (N_3909,N_3150,N_3373);
and U3910 (N_3910,N_3384,N_3062);
and U3911 (N_3911,N_3003,N_3045);
and U3912 (N_3912,N_3289,N_3087);
and U3913 (N_3913,N_3060,N_3460);
or U3914 (N_3914,N_3134,N_3331);
nand U3915 (N_3915,N_3021,N_3035);
and U3916 (N_3916,N_3326,N_3017);
nand U3917 (N_3917,N_3209,N_3139);
or U3918 (N_3918,N_3283,N_3011);
and U3919 (N_3919,N_3082,N_3239);
nor U3920 (N_3920,N_3287,N_3104);
nand U3921 (N_3921,N_3262,N_3005);
or U3922 (N_3922,N_3453,N_3380);
and U3923 (N_3923,N_3302,N_3338);
nor U3924 (N_3924,N_3440,N_3411);
nand U3925 (N_3925,N_3278,N_3102);
and U3926 (N_3926,N_3220,N_3443);
nor U3927 (N_3927,N_3021,N_3358);
nor U3928 (N_3928,N_3015,N_3482);
or U3929 (N_3929,N_3448,N_3063);
or U3930 (N_3930,N_3336,N_3121);
and U3931 (N_3931,N_3141,N_3434);
or U3932 (N_3932,N_3023,N_3323);
nand U3933 (N_3933,N_3202,N_3419);
and U3934 (N_3934,N_3133,N_3485);
nor U3935 (N_3935,N_3417,N_3420);
or U3936 (N_3936,N_3228,N_3145);
nor U3937 (N_3937,N_3077,N_3483);
nand U3938 (N_3938,N_3094,N_3205);
or U3939 (N_3939,N_3233,N_3190);
or U3940 (N_3940,N_3088,N_3010);
or U3941 (N_3941,N_3188,N_3068);
or U3942 (N_3942,N_3186,N_3041);
nor U3943 (N_3943,N_3446,N_3225);
nor U3944 (N_3944,N_3274,N_3328);
nand U3945 (N_3945,N_3356,N_3155);
and U3946 (N_3946,N_3475,N_3157);
or U3947 (N_3947,N_3132,N_3493);
and U3948 (N_3948,N_3457,N_3407);
nor U3949 (N_3949,N_3003,N_3303);
and U3950 (N_3950,N_3295,N_3495);
nor U3951 (N_3951,N_3286,N_3030);
and U3952 (N_3952,N_3235,N_3128);
or U3953 (N_3953,N_3467,N_3238);
nor U3954 (N_3954,N_3301,N_3291);
or U3955 (N_3955,N_3282,N_3268);
and U3956 (N_3956,N_3290,N_3378);
nand U3957 (N_3957,N_3103,N_3403);
nand U3958 (N_3958,N_3411,N_3248);
nor U3959 (N_3959,N_3255,N_3268);
and U3960 (N_3960,N_3258,N_3226);
nor U3961 (N_3961,N_3235,N_3136);
or U3962 (N_3962,N_3326,N_3185);
nor U3963 (N_3963,N_3431,N_3066);
nor U3964 (N_3964,N_3004,N_3231);
nor U3965 (N_3965,N_3436,N_3448);
nand U3966 (N_3966,N_3311,N_3163);
nand U3967 (N_3967,N_3373,N_3381);
nor U3968 (N_3968,N_3257,N_3483);
and U3969 (N_3969,N_3266,N_3190);
xnor U3970 (N_3970,N_3219,N_3124);
and U3971 (N_3971,N_3051,N_3364);
and U3972 (N_3972,N_3253,N_3227);
nor U3973 (N_3973,N_3140,N_3148);
and U3974 (N_3974,N_3039,N_3173);
or U3975 (N_3975,N_3060,N_3072);
or U3976 (N_3976,N_3191,N_3213);
nor U3977 (N_3977,N_3320,N_3214);
nor U3978 (N_3978,N_3397,N_3263);
or U3979 (N_3979,N_3386,N_3421);
nand U3980 (N_3980,N_3168,N_3239);
nand U3981 (N_3981,N_3222,N_3494);
or U3982 (N_3982,N_3444,N_3031);
nor U3983 (N_3983,N_3304,N_3287);
nand U3984 (N_3984,N_3393,N_3322);
or U3985 (N_3985,N_3396,N_3226);
or U3986 (N_3986,N_3272,N_3405);
or U3987 (N_3987,N_3038,N_3260);
and U3988 (N_3988,N_3134,N_3216);
nor U3989 (N_3989,N_3349,N_3444);
nor U3990 (N_3990,N_3093,N_3496);
nor U3991 (N_3991,N_3364,N_3421);
and U3992 (N_3992,N_3253,N_3155);
and U3993 (N_3993,N_3393,N_3039);
nor U3994 (N_3994,N_3294,N_3166);
or U3995 (N_3995,N_3117,N_3286);
and U3996 (N_3996,N_3420,N_3268);
and U3997 (N_3997,N_3293,N_3146);
nand U3998 (N_3998,N_3346,N_3448);
nor U3999 (N_3999,N_3468,N_3184);
nor U4000 (N_4000,N_3744,N_3611);
or U4001 (N_4001,N_3580,N_3655);
or U4002 (N_4002,N_3661,N_3576);
nor U4003 (N_4003,N_3685,N_3652);
nand U4004 (N_4004,N_3830,N_3686);
nor U4005 (N_4005,N_3837,N_3834);
nand U4006 (N_4006,N_3894,N_3940);
nand U4007 (N_4007,N_3500,N_3528);
nor U4008 (N_4008,N_3907,N_3753);
and U4009 (N_4009,N_3949,N_3647);
and U4010 (N_4010,N_3738,N_3663);
and U4011 (N_4011,N_3566,N_3970);
or U4012 (N_4012,N_3516,N_3570);
nand U4013 (N_4013,N_3918,N_3610);
and U4014 (N_4014,N_3881,N_3552);
nand U4015 (N_4015,N_3680,N_3897);
nand U4016 (N_4016,N_3936,N_3768);
nand U4017 (N_4017,N_3865,N_3653);
and U4018 (N_4018,N_3778,N_3850);
nor U4019 (N_4019,N_3715,N_3501);
or U4020 (N_4020,N_3641,N_3846);
and U4021 (N_4021,N_3793,N_3941);
or U4022 (N_4022,N_3542,N_3856);
and U4023 (N_4023,N_3898,N_3631);
or U4024 (N_4024,N_3607,N_3646);
nor U4025 (N_4025,N_3946,N_3529);
xor U4026 (N_4026,N_3947,N_3925);
nor U4027 (N_4027,N_3575,N_3562);
xor U4028 (N_4028,N_3887,N_3989);
and U4029 (N_4029,N_3687,N_3526);
nor U4030 (N_4030,N_3901,N_3809);
nand U4031 (N_4031,N_3730,N_3979);
nor U4032 (N_4032,N_3600,N_3513);
nand U4033 (N_4033,N_3863,N_3868);
and U4034 (N_4034,N_3882,N_3991);
nand U4035 (N_4035,N_3869,N_3756);
and U4036 (N_4036,N_3737,N_3975);
and U4037 (N_4037,N_3911,N_3832);
nor U4038 (N_4038,N_3779,N_3508);
nand U4039 (N_4039,N_3976,N_3914);
or U4040 (N_4040,N_3536,N_3801);
nor U4041 (N_4041,N_3594,N_3662);
or U4042 (N_4042,N_3681,N_3823);
nor U4043 (N_4043,N_3582,N_3533);
nand U4044 (N_4044,N_3884,N_3699);
or U4045 (N_4045,N_3598,N_3952);
and U4046 (N_4046,N_3588,N_3718);
xor U4047 (N_4047,N_3899,N_3571);
or U4048 (N_4048,N_3844,N_3617);
nand U4049 (N_4049,N_3568,N_3978);
or U4050 (N_4050,N_3831,N_3560);
and U4051 (N_4051,N_3710,N_3913);
and U4052 (N_4052,N_3980,N_3625);
nor U4053 (N_4053,N_3777,N_3740);
and U4054 (N_4054,N_3957,N_3602);
nor U4055 (N_4055,N_3593,N_3698);
or U4056 (N_4056,N_3822,N_3847);
or U4057 (N_4057,N_3569,N_3912);
nor U4058 (N_4058,N_3972,N_3992);
nor U4059 (N_4059,N_3728,N_3567);
nor U4060 (N_4060,N_3623,N_3998);
nand U4061 (N_4061,N_3919,N_3751);
nand U4062 (N_4062,N_3966,N_3731);
or U4063 (N_4063,N_3955,N_3961);
nand U4064 (N_4064,N_3608,N_3864);
and U4065 (N_4065,N_3609,N_3637);
nand U4066 (N_4066,N_3712,N_3807);
and U4067 (N_4067,N_3616,N_3761);
or U4068 (N_4068,N_3512,N_3942);
nor U4069 (N_4069,N_3620,N_3968);
nor U4070 (N_4070,N_3857,N_3732);
and U4071 (N_4071,N_3634,N_3999);
or U4072 (N_4072,N_3764,N_3904);
nand U4073 (N_4073,N_3951,N_3855);
and U4074 (N_4074,N_3648,N_3665);
nor U4075 (N_4075,N_3780,N_3725);
or U4076 (N_4076,N_3658,N_3595);
or U4077 (N_4077,N_3606,N_3987);
or U4078 (N_4078,N_3719,N_3675);
or U4079 (N_4079,N_3775,N_3826);
and U4080 (N_4080,N_3795,N_3910);
nand U4081 (N_4081,N_3541,N_3684);
nand U4082 (N_4082,N_3977,N_3592);
and U4083 (N_4083,N_3960,N_3814);
nor U4084 (N_4084,N_3532,N_3923);
or U4085 (N_4085,N_3633,N_3835);
nor U4086 (N_4086,N_3997,N_3547);
nor U4087 (N_4087,N_3693,N_3723);
and U4088 (N_4088,N_3587,N_3530);
nand U4089 (N_4089,N_3875,N_3804);
nor U4090 (N_4090,N_3510,N_3861);
or U4091 (N_4091,N_3578,N_3581);
nand U4092 (N_4092,N_3928,N_3971);
nor U4093 (N_4093,N_3591,N_3829);
nor U4094 (N_4094,N_3930,N_3599);
nor U4095 (N_4095,N_3691,N_3553);
nand U4096 (N_4096,N_3603,N_3983);
and U4097 (N_4097,N_3534,N_3762);
nand U4098 (N_4098,N_3852,N_3584);
nor U4099 (N_4099,N_3802,N_3618);
nand U4100 (N_4100,N_3917,N_3706);
nand U4101 (N_4101,N_3676,N_3805);
nand U4102 (N_4102,N_3745,N_3798);
nand U4103 (N_4103,N_3996,N_3563);
and U4104 (N_4104,N_3962,N_3511);
or U4105 (N_4105,N_3702,N_3916);
nor U4106 (N_4106,N_3994,N_3520);
nand U4107 (N_4107,N_3726,N_3736);
nand U4108 (N_4108,N_3927,N_3721);
nand U4109 (N_4109,N_3539,N_3810);
nand U4110 (N_4110,N_3935,N_3836);
and U4111 (N_4111,N_3514,N_3880);
nor U4112 (N_4112,N_3773,N_3729);
nand U4113 (N_4113,N_3550,N_3808);
and U4114 (N_4114,N_3853,N_3589);
nor U4115 (N_4115,N_3555,N_3890);
nor U4116 (N_4116,N_3540,N_3689);
nand U4117 (N_4117,N_3903,N_3796);
nand U4118 (N_4118,N_3614,N_3934);
and U4119 (N_4119,N_3985,N_3818);
or U4120 (N_4120,N_3671,N_3551);
and U4121 (N_4121,N_3733,N_3895);
and U4122 (N_4122,N_3554,N_3943);
nor U4123 (N_4123,N_3694,N_3544);
and U4124 (N_4124,N_3522,N_3921);
and U4125 (N_4125,N_3527,N_3817);
nand U4126 (N_4126,N_3537,N_3507);
nor U4127 (N_4127,N_3650,N_3848);
nand U4128 (N_4128,N_3774,N_3759);
nand U4129 (N_4129,N_3535,N_3871);
or U4130 (N_4130,N_3543,N_3549);
and U4131 (N_4131,N_3776,N_3678);
nand U4132 (N_4132,N_3883,N_3643);
nor U4133 (N_4133,N_3788,N_3765);
nor U4134 (N_4134,N_3644,N_3717);
nand U4135 (N_4135,N_3673,N_3659);
and U4136 (N_4136,N_3866,N_3929);
or U4137 (N_4137,N_3878,N_3629);
nor U4138 (N_4138,N_3859,N_3521);
nand U4139 (N_4139,N_3735,N_3749);
nor U4140 (N_4140,N_3626,N_3724);
nand U4141 (N_4141,N_3790,N_3757);
and U4142 (N_4142,N_3615,N_3954);
and U4143 (N_4143,N_3622,N_3639);
nand U4144 (N_4144,N_3619,N_3766);
nand U4145 (N_4145,N_3915,N_3771);
and U4146 (N_4146,N_3945,N_3789);
nand U4147 (N_4147,N_3502,N_3799);
nand U4148 (N_4148,N_3937,N_3654);
and U4149 (N_4149,N_3666,N_3565);
xor U4150 (N_4150,N_3677,N_3656);
nor U4151 (N_4151,N_3583,N_3548);
nand U4152 (N_4152,N_3703,N_3862);
nand U4153 (N_4153,N_3932,N_3843);
nor U4154 (N_4154,N_3969,N_3519);
nand U4155 (N_4155,N_3959,N_3574);
nand U4156 (N_4156,N_3948,N_3931);
nand U4157 (N_4157,N_3791,N_3748);
nor U4158 (N_4158,N_3752,N_3523);
nor U4159 (N_4159,N_3596,N_3638);
and U4160 (N_4160,N_3545,N_3953);
nand U4161 (N_4161,N_3640,N_3630);
or U4162 (N_4162,N_3700,N_3900);
or U4163 (N_4163,N_3995,N_3964);
or U4164 (N_4164,N_3585,N_3770);
nand U4165 (N_4165,N_3896,N_3908);
or U4166 (N_4166,N_3785,N_3632);
nor U4167 (N_4167,N_3559,N_3696);
nand U4168 (N_4168,N_3509,N_3842);
nand U4169 (N_4169,N_3709,N_3819);
nor U4170 (N_4170,N_3813,N_3950);
and U4171 (N_4171,N_3668,N_3982);
nor U4172 (N_4172,N_3743,N_3739);
and U4173 (N_4173,N_3538,N_3783);
and U4174 (N_4174,N_3993,N_3682);
or U4175 (N_4175,N_3926,N_3572);
nand U4176 (N_4176,N_3704,N_3613);
nor U4177 (N_4177,N_3605,N_3628);
or U4178 (N_4178,N_3839,N_3933);
nor U4179 (N_4179,N_3590,N_3672);
and U4180 (N_4180,N_3742,N_3909);
nor U4181 (N_4181,N_3722,N_3664);
nor U4182 (N_4182,N_3504,N_3838);
or U4183 (N_4183,N_3797,N_3956);
nor U4184 (N_4184,N_3787,N_3860);
or U4185 (N_4185,N_3651,N_3758);
nor U4186 (N_4186,N_3827,N_3924);
nor U4187 (N_4187,N_3760,N_3657);
and U4188 (N_4188,N_3558,N_3747);
and U4189 (N_4189,N_3573,N_3701);
and U4190 (N_4190,N_3825,N_3828);
nand U4191 (N_4191,N_3794,N_3531);
or U4192 (N_4192,N_3645,N_3517);
and U4193 (N_4193,N_3988,N_3800);
nand U4194 (N_4194,N_3984,N_3958);
nor U4195 (N_4195,N_3873,N_3889);
and U4196 (N_4196,N_3627,N_3683);
nand U4197 (N_4197,N_3525,N_3518);
nand U4198 (N_4198,N_3679,N_3811);
and U4199 (N_4199,N_3965,N_3967);
or U4200 (N_4200,N_3515,N_3944);
or U4201 (N_4201,N_3697,N_3816);
nand U4202 (N_4202,N_3750,N_3867);
nor U4203 (N_4203,N_3782,N_3746);
nand U4204 (N_4204,N_3755,N_3784);
and U4205 (N_4205,N_3561,N_3711);
or U4206 (N_4206,N_3688,N_3604);
and U4207 (N_4207,N_3635,N_3886);
or U4208 (N_4208,N_3874,N_3674);
or U4209 (N_4209,N_3769,N_3524);
and U4210 (N_4210,N_3872,N_3939);
nor U4211 (N_4211,N_3845,N_3705);
nand U4212 (N_4212,N_3564,N_3877);
or U4213 (N_4213,N_3597,N_3905);
and U4214 (N_4214,N_3891,N_3893);
or U4215 (N_4215,N_3660,N_3849);
nor U4216 (N_4216,N_3986,N_3754);
or U4217 (N_4217,N_3690,N_3556);
or U4218 (N_4218,N_3990,N_3579);
nand U4219 (N_4219,N_3727,N_3505);
and U4220 (N_4220,N_3557,N_3767);
nand U4221 (N_4221,N_3888,N_3920);
nand U4222 (N_4222,N_3708,N_3624);
nand U4223 (N_4223,N_3649,N_3546);
nand U4224 (N_4224,N_3612,N_3786);
nand U4225 (N_4225,N_3707,N_3636);
or U4226 (N_4226,N_3621,N_3841);
and U4227 (N_4227,N_3821,N_3840);
nor U4228 (N_4228,N_3669,N_3506);
nor U4229 (N_4229,N_3902,N_3851);
or U4230 (N_4230,N_3876,N_3885);
and U4231 (N_4231,N_3670,N_3734);
or U4232 (N_4232,N_3870,N_3781);
or U4233 (N_4233,N_3667,N_3858);
nand U4234 (N_4234,N_3906,N_3963);
nor U4235 (N_4235,N_3695,N_3763);
or U4236 (N_4236,N_3503,N_3974);
nand U4237 (N_4237,N_3973,N_3833);
nand U4238 (N_4238,N_3692,N_3981);
nand U4239 (N_4239,N_3922,N_3716);
nand U4240 (N_4240,N_3812,N_3642);
and U4241 (N_4241,N_3586,N_3601);
nor U4242 (N_4242,N_3803,N_3820);
nor U4243 (N_4243,N_3824,N_3879);
or U4244 (N_4244,N_3713,N_3806);
and U4245 (N_4245,N_3792,N_3772);
or U4246 (N_4246,N_3741,N_3938);
or U4247 (N_4247,N_3714,N_3577);
or U4248 (N_4248,N_3815,N_3854);
nand U4249 (N_4249,N_3892,N_3720);
nand U4250 (N_4250,N_3841,N_3556);
nand U4251 (N_4251,N_3602,N_3971);
nand U4252 (N_4252,N_3572,N_3723);
or U4253 (N_4253,N_3567,N_3630);
nor U4254 (N_4254,N_3592,N_3768);
nand U4255 (N_4255,N_3955,N_3732);
and U4256 (N_4256,N_3837,N_3700);
and U4257 (N_4257,N_3563,N_3810);
and U4258 (N_4258,N_3600,N_3641);
or U4259 (N_4259,N_3508,N_3808);
xnor U4260 (N_4260,N_3665,N_3586);
nand U4261 (N_4261,N_3844,N_3734);
and U4262 (N_4262,N_3642,N_3734);
nand U4263 (N_4263,N_3533,N_3517);
xor U4264 (N_4264,N_3649,N_3533);
and U4265 (N_4265,N_3854,N_3833);
nor U4266 (N_4266,N_3912,N_3919);
nor U4267 (N_4267,N_3587,N_3737);
and U4268 (N_4268,N_3850,N_3508);
and U4269 (N_4269,N_3684,N_3797);
nand U4270 (N_4270,N_3581,N_3689);
or U4271 (N_4271,N_3935,N_3657);
nand U4272 (N_4272,N_3832,N_3965);
and U4273 (N_4273,N_3711,N_3579);
and U4274 (N_4274,N_3543,N_3831);
nor U4275 (N_4275,N_3871,N_3807);
nand U4276 (N_4276,N_3851,N_3572);
nor U4277 (N_4277,N_3508,N_3623);
nand U4278 (N_4278,N_3674,N_3797);
and U4279 (N_4279,N_3630,N_3748);
or U4280 (N_4280,N_3572,N_3592);
or U4281 (N_4281,N_3723,N_3592);
or U4282 (N_4282,N_3640,N_3735);
nor U4283 (N_4283,N_3998,N_3656);
or U4284 (N_4284,N_3784,N_3745);
nand U4285 (N_4285,N_3965,N_3568);
or U4286 (N_4286,N_3821,N_3799);
and U4287 (N_4287,N_3880,N_3552);
and U4288 (N_4288,N_3603,N_3696);
or U4289 (N_4289,N_3814,N_3927);
and U4290 (N_4290,N_3997,N_3833);
or U4291 (N_4291,N_3849,N_3580);
nor U4292 (N_4292,N_3933,N_3528);
nor U4293 (N_4293,N_3889,N_3545);
nand U4294 (N_4294,N_3578,N_3617);
nand U4295 (N_4295,N_3535,N_3840);
and U4296 (N_4296,N_3981,N_3718);
nor U4297 (N_4297,N_3791,N_3933);
and U4298 (N_4298,N_3756,N_3710);
nor U4299 (N_4299,N_3536,N_3508);
nor U4300 (N_4300,N_3588,N_3920);
nor U4301 (N_4301,N_3532,N_3627);
nand U4302 (N_4302,N_3682,N_3743);
and U4303 (N_4303,N_3682,N_3630);
nor U4304 (N_4304,N_3838,N_3659);
nand U4305 (N_4305,N_3868,N_3691);
nor U4306 (N_4306,N_3559,N_3750);
or U4307 (N_4307,N_3835,N_3979);
or U4308 (N_4308,N_3619,N_3651);
nor U4309 (N_4309,N_3685,N_3960);
nor U4310 (N_4310,N_3711,N_3596);
nor U4311 (N_4311,N_3513,N_3679);
nand U4312 (N_4312,N_3637,N_3759);
nor U4313 (N_4313,N_3903,N_3829);
or U4314 (N_4314,N_3908,N_3544);
and U4315 (N_4315,N_3745,N_3642);
nor U4316 (N_4316,N_3912,N_3935);
nor U4317 (N_4317,N_3857,N_3975);
nor U4318 (N_4318,N_3978,N_3836);
nor U4319 (N_4319,N_3796,N_3753);
and U4320 (N_4320,N_3653,N_3550);
nor U4321 (N_4321,N_3750,N_3928);
nand U4322 (N_4322,N_3832,N_3816);
nand U4323 (N_4323,N_3620,N_3754);
or U4324 (N_4324,N_3732,N_3571);
nor U4325 (N_4325,N_3681,N_3897);
nor U4326 (N_4326,N_3507,N_3964);
or U4327 (N_4327,N_3507,N_3867);
nand U4328 (N_4328,N_3808,N_3598);
nand U4329 (N_4329,N_3993,N_3542);
and U4330 (N_4330,N_3532,N_3571);
nand U4331 (N_4331,N_3599,N_3740);
and U4332 (N_4332,N_3786,N_3510);
and U4333 (N_4333,N_3969,N_3795);
or U4334 (N_4334,N_3898,N_3948);
or U4335 (N_4335,N_3541,N_3812);
nand U4336 (N_4336,N_3518,N_3865);
nand U4337 (N_4337,N_3810,N_3742);
nand U4338 (N_4338,N_3842,N_3745);
or U4339 (N_4339,N_3536,N_3501);
or U4340 (N_4340,N_3564,N_3792);
nor U4341 (N_4341,N_3866,N_3921);
nand U4342 (N_4342,N_3987,N_3893);
nand U4343 (N_4343,N_3801,N_3628);
nand U4344 (N_4344,N_3960,N_3976);
and U4345 (N_4345,N_3750,N_3912);
nor U4346 (N_4346,N_3699,N_3890);
and U4347 (N_4347,N_3943,N_3957);
nor U4348 (N_4348,N_3616,N_3572);
or U4349 (N_4349,N_3599,N_3809);
or U4350 (N_4350,N_3887,N_3731);
nand U4351 (N_4351,N_3779,N_3557);
nand U4352 (N_4352,N_3841,N_3654);
and U4353 (N_4353,N_3685,N_3828);
nor U4354 (N_4354,N_3983,N_3535);
nor U4355 (N_4355,N_3565,N_3870);
or U4356 (N_4356,N_3533,N_3716);
nor U4357 (N_4357,N_3513,N_3580);
nand U4358 (N_4358,N_3681,N_3596);
nor U4359 (N_4359,N_3913,N_3785);
nor U4360 (N_4360,N_3662,N_3551);
or U4361 (N_4361,N_3964,N_3623);
and U4362 (N_4362,N_3789,N_3979);
and U4363 (N_4363,N_3926,N_3538);
and U4364 (N_4364,N_3630,N_3596);
nand U4365 (N_4365,N_3839,N_3511);
nor U4366 (N_4366,N_3699,N_3716);
nand U4367 (N_4367,N_3590,N_3513);
nor U4368 (N_4368,N_3687,N_3959);
and U4369 (N_4369,N_3902,N_3704);
and U4370 (N_4370,N_3791,N_3892);
or U4371 (N_4371,N_3974,N_3786);
and U4372 (N_4372,N_3789,N_3686);
nor U4373 (N_4373,N_3924,N_3549);
nor U4374 (N_4374,N_3609,N_3848);
nor U4375 (N_4375,N_3542,N_3701);
nor U4376 (N_4376,N_3686,N_3618);
nor U4377 (N_4377,N_3870,N_3690);
nand U4378 (N_4378,N_3533,N_3669);
or U4379 (N_4379,N_3565,N_3992);
nor U4380 (N_4380,N_3705,N_3602);
nand U4381 (N_4381,N_3705,N_3626);
nor U4382 (N_4382,N_3844,N_3555);
nor U4383 (N_4383,N_3618,N_3631);
and U4384 (N_4384,N_3659,N_3771);
and U4385 (N_4385,N_3792,N_3945);
nor U4386 (N_4386,N_3961,N_3654);
or U4387 (N_4387,N_3858,N_3749);
and U4388 (N_4388,N_3821,N_3837);
or U4389 (N_4389,N_3672,N_3804);
nor U4390 (N_4390,N_3677,N_3993);
nand U4391 (N_4391,N_3683,N_3635);
or U4392 (N_4392,N_3678,N_3995);
and U4393 (N_4393,N_3910,N_3842);
nor U4394 (N_4394,N_3718,N_3627);
and U4395 (N_4395,N_3514,N_3745);
nor U4396 (N_4396,N_3851,N_3696);
nand U4397 (N_4397,N_3591,N_3946);
or U4398 (N_4398,N_3981,N_3934);
and U4399 (N_4399,N_3959,N_3547);
or U4400 (N_4400,N_3681,N_3758);
or U4401 (N_4401,N_3618,N_3923);
nor U4402 (N_4402,N_3858,N_3645);
or U4403 (N_4403,N_3506,N_3639);
or U4404 (N_4404,N_3503,N_3519);
nand U4405 (N_4405,N_3809,N_3928);
nor U4406 (N_4406,N_3999,N_3879);
nor U4407 (N_4407,N_3684,N_3532);
nand U4408 (N_4408,N_3585,N_3908);
or U4409 (N_4409,N_3971,N_3519);
or U4410 (N_4410,N_3611,N_3570);
nand U4411 (N_4411,N_3687,N_3622);
nand U4412 (N_4412,N_3785,N_3728);
and U4413 (N_4413,N_3822,N_3583);
and U4414 (N_4414,N_3842,N_3594);
or U4415 (N_4415,N_3926,N_3517);
nand U4416 (N_4416,N_3548,N_3846);
nor U4417 (N_4417,N_3894,N_3779);
or U4418 (N_4418,N_3921,N_3847);
or U4419 (N_4419,N_3517,N_3754);
nor U4420 (N_4420,N_3979,N_3930);
and U4421 (N_4421,N_3652,N_3751);
nor U4422 (N_4422,N_3771,N_3920);
nand U4423 (N_4423,N_3871,N_3532);
or U4424 (N_4424,N_3727,N_3986);
or U4425 (N_4425,N_3587,N_3856);
and U4426 (N_4426,N_3804,N_3508);
and U4427 (N_4427,N_3888,N_3810);
or U4428 (N_4428,N_3830,N_3998);
nor U4429 (N_4429,N_3981,N_3829);
and U4430 (N_4430,N_3504,N_3825);
and U4431 (N_4431,N_3868,N_3748);
nor U4432 (N_4432,N_3630,N_3959);
or U4433 (N_4433,N_3697,N_3602);
and U4434 (N_4434,N_3736,N_3881);
nor U4435 (N_4435,N_3739,N_3853);
nand U4436 (N_4436,N_3895,N_3816);
xor U4437 (N_4437,N_3904,N_3583);
nor U4438 (N_4438,N_3966,N_3709);
nor U4439 (N_4439,N_3809,N_3780);
nand U4440 (N_4440,N_3785,N_3556);
or U4441 (N_4441,N_3762,N_3809);
or U4442 (N_4442,N_3563,N_3959);
or U4443 (N_4443,N_3740,N_3582);
and U4444 (N_4444,N_3945,N_3708);
nand U4445 (N_4445,N_3810,N_3775);
nor U4446 (N_4446,N_3934,N_3665);
or U4447 (N_4447,N_3809,N_3848);
or U4448 (N_4448,N_3501,N_3691);
nand U4449 (N_4449,N_3656,N_3858);
nand U4450 (N_4450,N_3792,N_3930);
or U4451 (N_4451,N_3814,N_3598);
nor U4452 (N_4452,N_3826,N_3572);
nand U4453 (N_4453,N_3505,N_3716);
and U4454 (N_4454,N_3779,N_3548);
nand U4455 (N_4455,N_3815,N_3694);
nor U4456 (N_4456,N_3723,N_3755);
or U4457 (N_4457,N_3788,N_3735);
or U4458 (N_4458,N_3578,N_3827);
nand U4459 (N_4459,N_3926,N_3504);
and U4460 (N_4460,N_3857,N_3897);
or U4461 (N_4461,N_3704,N_3677);
nand U4462 (N_4462,N_3753,N_3555);
nor U4463 (N_4463,N_3909,N_3775);
nand U4464 (N_4464,N_3778,N_3722);
nand U4465 (N_4465,N_3944,N_3558);
nor U4466 (N_4466,N_3616,N_3938);
nor U4467 (N_4467,N_3954,N_3608);
nand U4468 (N_4468,N_3735,N_3845);
and U4469 (N_4469,N_3670,N_3991);
or U4470 (N_4470,N_3728,N_3862);
nand U4471 (N_4471,N_3851,N_3561);
or U4472 (N_4472,N_3705,N_3564);
and U4473 (N_4473,N_3549,N_3738);
or U4474 (N_4474,N_3738,N_3629);
and U4475 (N_4475,N_3855,N_3996);
or U4476 (N_4476,N_3754,N_3963);
nand U4477 (N_4477,N_3615,N_3627);
nor U4478 (N_4478,N_3588,N_3886);
nor U4479 (N_4479,N_3693,N_3760);
or U4480 (N_4480,N_3775,N_3736);
or U4481 (N_4481,N_3571,N_3721);
nand U4482 (N_4482,N_3886,N_3959);
xnor U4483 (N_4483,N_3581,N_3810);
nand U4484 (N_4484,N_3602,N_3571);
nor U4485 (N_4485,N_3989,N_3855);
or U4486 (N_4486,N_3836,N_3616);
or U4487 (N_4487,N_3935,N_3568);
and U4488 (N_4488,N_3912,N_3754);
nor U4489 (N_4489,N_3678,N_3684);
nor U4490 (N_4490,N_3661,N_3553);
or U4491 (N_4491,N_3836,N_3628);
and U4492 (N_4492,N_3990,N_3558);
and U4493 (N_4493,N_3900,N_3533);
nand U4494 (N_4494,N_3810,N_3504);
and U4495 (N_4495,N_3813,N_3819);
and U4496 (N_4496,N_3902,N_3640);
nor U4497 (N_4497,N_3627,N_3775);
nor U4498 (N_4498,N_3761,N_3603);
nand U4499 (N_4499,N_3995,N_3967);
nand U4500 (N_4500,N_4060,N_4196);
and U4501 (N_4501,N_4365,N_4072);
and U4502 (N_4502,N_4013,N_4306);
nor U4503 (N_4503,N_4165,N_4046);
nand U4504 (N_4504,N_4349,N_4273);
nor U4505 (N_4505,N_4333,N_4201);
nand U4506 (N_4506,N_4498,N_4023);
or U4507 (N_4507,N_4081,N_4454);
and U4508 (N_4508,N_4112,N_4123);
and U4509 (N_4509,N_4445,N_4444);
nand U4510 (N_4510,N_4235,N_4172);
and U4511 (N_4511,N_4101,N_4193);
nand U4512 (N_4512,N_4077,N_4153);
or U4513 (N_4513,N_4238,N_4326);
nand U4514 (N_4514,N_4400,N_4405);
and U4515 (N_4515,N_4259,N_4140);
and U4516 (N_4516,N_4006,N_4265);
nand U4517 (N_4517,N_4499,N_4244);
nand U4518 (N_4518,N_4103,N_4262);
or U4519 (N_4519,N_4299,N_4289);
or U4520 (N_4520,N_4319,N_4404);
nand U4521 (N_4521,N_4494,N_4082);
nor U4522 (N_4522,N_4144,N_4460);
or U4523 (N_4523,N_4314,N_4278);
or U4524 (N_4524,N_4078,N_4045);
or U4525 (N_4525,N_4497,N_4455);
or U4526 (N_4526,N_4426,N_4474);
nor U4527 (N_4527,N_4283,N_4166);
nand U4528 (N_4528,N_4363,N_4391);
and U4529 (N_4529,N_4020,N_4067);
or U4530 (N_4530,N_4243,N_4209);
nor U4531 (N_4531,N_4245,N_4486);
nor U4532 (N_4532,N_4302,N_4431);
and U4533 (N_4533,N_4436,N_4441);
nand U4534 (N_4534,N_4121,N_4155);
and U4535 (N_4535,N_4128,N_4254);
nor U4536 (N_4536,N_4312,N_4104);
nand U4537 (N_4537,N_4269,N_4401);
xor U4538 (N_4538,N_4068,N_4053);
or U4539 (N_4539,N_4339,N_4105);
and U4540 (N_4540,N_4371,N_4040);
or U4541 (N_4541,N_4424,N_4331);
or U4542 (N_4542,N_4233,N_4458);
and U4543 (N_4543,N_4228,N_4096);
and U4544 (N_4544,N_4202,N_4145);
nand U4545 (N_4545,N_4329,N_4280);
and U4546 (N_4546,N_4465,N_4386);
or U4547 (N_4547,N_4217,N_4059);
nor U4548 (N_4548,N_4338,N_4159);
nor U4549 (N_4549,N_4242,N_4032);
or U4550 (N_4550,N_4161,N_4004);
nand U4551 (N_4551,N_4291,N_4396);
or U4552 (N_4552,N_4050,N_4357);
and U4553 (N_4553,N_4070,N_4197);
or U4554 (N_4554,N_4021,N_4073);
nand U4555 (N_4555,N_4352,N_4389);
nand U4556 (N_4556,N_4491,N_4071);
nand U4557 (N_4557,N_4025,N_4261);
nand U4558 (N_4558,N_4055,N_4337);
and U4559 (N_4559,N_4147,N_4394);
or U4560 (N_4560,N_4036,N_4198);
xnor U4561 (N_4561,N_4210,N_4415);
nor U4562 (N_4562,N_4037,N_4309);
and U4563 (N_4563,N_4100,N_4124);
and U4564 (N_4564,N_4179,N_4409);
or U4565 (N_4565,N_4336,N_4276);
or U4566 (N_4566,N_4324,N_4168);
xnor U4567 (N_4567,N_4018,N_4412);
or U4568 (N_4568,N_4419,N_4133);
nand U4569 (N_4569,N_4328,N_4093);
and U4570 (N_4570,N_4019,N_4051);
nor U4571 (N_4571,N_4322,N_4281);
and U4572 (N_4572,N_4111,N_4129);
or U4573 (N_4573,N_4471,N_4134);
nor U4574 (N_4574,N_4315,N_4251);
nor U4575 (N_4575,N_4479,N_4260);
and U4576 (N_4576,N_4402,N_4122);
xnor U4577 (N_4577,N_4493,N_4170);
and U4578 (N_4578,N_4447,N_4188);
nor U4579 (N_4579,N_4301,N_4407);
or U4580 (N_4580,N_4131,N_4249);
nand U4581 (N_4581,N_4485,N_4113);
nand U4582 (N_4582,N_4156,N_4207);
nor U4583 (N_4583,N_4219,N_4086);
and U4584 (N_4584,N_4057,N_4483);
nor U4585 (N_4585,N_4293,N_4359);
and U4586 (N_4586,N_4195,N_4489);
nor U4587 (N_4587,N_4488,N_4164);
or U4588 (N_4588,N_4038,N_4356);
and U4589 (N_4589,N_4468,N_4017);
or U4590 (N_4590,N_4169,N_4181);
and U4591 (N_4591,N_4298,N_4440);
nor U4592 (N_4592,N_4184,N_4061);
nand U4593 (N_4593,N_4204,N_4380);
nand U4594 (N_4594,N_4099,N_4428);
nor U4595 (N_4595,N_4208,N_4403);
and U4596 (N_4596,N_4158,N_4229);
nor U4597 (N_4597,N_4152,N_4002);
nor U4598 (N_4598,N_4031,N_4080);
or U4599 (N_4599,N_4011,N_4150);
and U4600 (N_4600,N_4342,N_4285);
and U4601 (N_4601,N_4360,N_4212);
nand U4602 (N_4602,N_4347,N_4425);
nand U4603 (N_4603,N_4343,N_4496);
nor U4604 (N_4604,N_4227,N_4463);
nand U4605 (N_4605,N_4149,N_4015);
nand U4606 (N_4606,N_4054,N_4484);
or U4607 (N_4607,N_4028,N_4058);
nor U4608 (N_4608,N_4317,N_4437);
or U4609 (N_4609,N_4139,N_4399);
nor U4610 (N_4610,N_4423,N_4182);
nor U4611 (N_4611,N_4237,N_4187);
nand U4612 (N_4612,N_4065,N_4146);
nand U4613 (N_4613,N_4287,N_4034);
and U4614 (N_4614,N_4030,N_4282);
or U4615 (N_4615,N_4473,N_4033);
or U4616 (N_4616,N_4115,N_4083);
and U4617 (N_4617,N_4213,N_4016);
nor U4618 (N_4618,N_4316,N_4064);
nand U4619 (N_4619,N_4481,N_4022);
nor U4620 (N_4620,N_4464,N_4413);
and U4621 (N_4621,N_4452,N_4069);
and U4622 (N_4622,N_4010,N_4087);
and U4623 (N_4623,N_4175,N_4305);
xor U4624 (N_4624,N_4221,N_4311);
or U4625 (N_4625,N_4374,N_4120);
or U4626 (N_4626,N_4255,N_4137);
nor U4627 (N_4627,N_4390,N_4239);
xor U4628 (N_4628,N_4325,N_4286);
or U4629 (N_4629,N_4194,N_4226);
and U4630 (N_4630,N_4205,N_4236);
or U4631 (N_4631,N_4014,N_4354);
nand U4632 (N_4632,N_4151,N_4108);
nand U4633 (N_4633,N_4272,N_4136);
nand U4634 (N_4634,N_4183,N_4477);
nor U4635 (N_4635,N_4167,N_4098);
nand U4636 (N_4636,N_4252,N_4148);
or U4637 (N_4637,N_4308,N_4005);
nand U4638 (N_4638,N_4117,N_4266);
nand U4639 (N_4639,N_4476,N_4443);
nand U4640 (N_4640,N_4327,N_4049);
nand U4641 (N_4641,N_4351,N_4384);
nor U4642 (N_4642,N_4085,N_4001);
nor U4643 (N_4643,N_4303,N_4421);
or U4644 (N_4644,N_4110,N_4430);
nor U4645 (N_4645,N_4387,N_4066);
nor U4646 (N_4646,N_4089,N_4224);
nor U4647 (N_4647,N_4388,N_4042);
or U4648 (N_4648,N_4230,N_4162);
or U4649 (N_4649,N_4130,N_4368);
nand U4650 (N_4650,N_4027,N_4275);
and U4651 (N_4651,N_4366,N_4459);
nor U4652 (N_4652,N_4264,N_4041);
nor U4653 (N_4653,N_4076,N_4433);
nor U4654 (N_4654,N_4457,N_4469);
and U4655 (N_4655,N_4330,N_4418);
xnor U4656 (N_4656,N_4092,N_4417);
or U4657 (N_4657,N_4383,N_4449);
and U4658 (N_4658,N_4190,N_4218);
or U4659 (N_4659,N_4408,N_4176);
nand U4660 (N_4660,N_4012,N_4127);
nand U4661 (N_4661,N_4332,N_4231);
nand U4662 (N_4662,N_4379,N_4478);
and U4663 (N_4663,N_4313,N_4398);
or U4664 (N_4664,N_4043,N_4392);
or U4665 (N_4665,N_4307,N_4373);
nand U4666 (N_4666,N_4106,N_4257);
xor U4667 (N_4667,N_4296,N_4340);
nand U4668 (N_4668,N_4186,N_4422);
or U4669 (N_4669,N_4321,N_4375);
nor U4670 (N_4670,N_4482,N_4263);
or U4671 (N_4671,N_4267,N_4125);
nand U4672 (N_4672,N_4427,N_4344);
and U4673 (N_4673,N_4116,N_4088);
and U4674 (N_4674,N_4126,N_4284);
nor U4675 (N_4675,N_4397,N_4461);
nand U4676 (N_4676,N_4029,N_4138);
or U4677 (N_4677,N_4318,N_4420);
nor U4678 (N_4678,N_4044,N_4353);
or U4679 (N_4679,N_4438,N_4240);
xor U4680 (N_4680,N_4174,N_4079);
or U4681 (N_4681,N_4300,N_4102);
nor U4682 (N_4682,N_4450,N_4211);
and U4683 (N_4683,N_4487,N_4268);
nand U4684 (N_4684,N_4395,N_4256);
and U4685 (N_4685,N_4185,N_4372);
nor U4686 (N_4686,N_4382,N_4406);
nand U4687 (N_4687,N_4432,N_4361);
nand U4688 (N_4688,N_4270,N_4090);
nor U4689 (N_4689,N_4097,N_4056);
or U4690 (N_4690,N_4157,N_4214);
nand U4691 (N_4691,N_4446,N_4295);
nand U4692 (N_4692,N_4203,N_4304);
nor U4693 (N_4693,N_4492,N_4414);
nand U4694 (N_4694,N_4323,N_4075);
and U4695 (N_4695,N_4035,N_4490);
and U4696 (N_4696,N_4191,N_4451);
nor U4697 (N_4697,N_4480,N_4223);
or U4698 (N_4698,N_4225,N_4345);
and U4699 (N_4699,N_4114,N_4290);
and U4700 (N_4700,N_4119,N_4495);
nand U4701 (N_4701,N_4132,N_4385);
nand U4702 (N_4702,N_4222,N_4220);
or U4703 (N_4703,N_4253,N_4074);
nor U4704 (N_4704,N_4376,N_4335);
or U4705 (N_4705,N_4355,N_4358);
nor U4706 (N_4706,N_4442,N_4448);
nand U4707 (N_4707,N_4393,N_4334);
and U4708 (N_4708,N_4274,N_4142);
nor U4709 (N_4709,N_4258,N_4362);
or U4710 (N_4710,N_4206,N_4277);
and U4711 (N_4711,N_4234,N_4416);
and U4712 (N_4712,N_4434,N_4466);
nand U4713 (N_4713,N_4118,N_4216);
nor U4714 (N_4714,N_4135,N_4310);
nor U4715 (N_4715,N_4154,N_4232);
or U4716 (N_4716,N_4297,N_4271);
and U4717 (N_4717,N_4288,N_4435);
and U4718 (N_4718,N_4364,N_4063);
and U4719 (N_4719,N_4009,N_4143);
or U4720 (N_4720,N_4160,N_4279);
or U4721 (N_4721,N_4350,N_4008);
or U4722 (N_4722,N_4370,N_4007);
and U4723 (N_4723,N_4200,N_4456);
nor U4724 (N_4724,N_4091,N_4346);
nand U4725 (N_4725,N_4367,N_4248);
nor U4726 (N_4726,N_4052,N_4178);
xor U4727 (N_4727,N_4163,N_4378);
nand U4728 (N_4728,N_4024,N_4247);
nor U4729 (N_4729,N_4062,N_4439);
nor U4730 (N_4730,N_4199,N_4003);
and U4731 (N_4731,N_4453,N_4189);
or U4732 (N_4732,N_4410,N_4246);
and U4733 (N_4733,N_4177,N_4381);
nor U4734 (N_4734,N_4348,N_4215);
or U4735 (N_4735,N_4369,N_4429);
or U4736 (N_4736,N_4320,N_4250);
and U4737 (N_4737,N_4173,N_4462);
or U4738 (N_4738,N_4475,N_4094);
nor U4739 (N_4739,N_4292,N_4411);
nand U4740 (N_4740,N_4047,N_4241);
or U4741 (N_4741,N_4048,N_4294);
or U4742 (N_4742,N_4039,N_4341);
nor U4743 (N_4743,N_4095,N_4107);
or U4744 (N_4744,N_4472,N_4467);
and U4745 (N_4745,N_4141,N_4171);
and U4746 (N_4746,N_4377,N_4026);
nand U4747 (N_4747,N_4109,N_4180);
nor U4748 (N_4748,N_4192,N_4000);
or U4749 (N_4749,N_4084,N_4470);
and U4750 (N_4750,N_4079,N_4287);
or U4751 (N_4751,N_4492,N_4335);
and U4752 (N_4752,N_4478,N_4056);
and U4753 (N_4753,N_4191,N_4460);
nor U4754 (N_4754,N_4165,N_4385);
nand U4755 (N_4755,N_4129,N_4265);
or U4756 (N_4756,N_4200,N_4289);
and U4757 (N_4757,N_4138,N_4122);
nand U4758 (N_4758,N_4233,N_4360);
and U4759 (N_4759,N_4145,N_4459);
and U4760 (N_4760,N_4070,N_4108);
and U4761 (N_4761,N_4435,N_4480);
or U4762 (N_4762,N_4130,N_4016);
and U4763 (N_4763,N_4498,N_4233);
nand U4764 (N_4764,N_4237,N_4260);
or U4765 (N_4765,N_4205,N_4312);
and U4766 (N_4766,N_4183,N_4385);
or U4767 (N_4767,N_4271,N_4371);
nor U4768 (N_4768,N_4300,N_4424);
or U4769 (N_4769,N_4166,N_4221);
or U4770 (N_4770,N_4065,N_4219);
or U4771 (N_4771,N_4428,N_4176);
nor U4772 (N_4772,N_4046,N_4293);
nor U4773 (N_4773,N_4348,N_4363);
and U4774 (N_4774,N_4263,N_4311);
and U4775 (N_4775,N_4080,N_4244);
nand U4776 (N_4776,N_4084,N_4417);
nor U4777 (N_4777,N_4208,N_4364);
nand U4778 (N_4778,N_4471,N_4414);
or U4779 (N_4779,N_4441,N_4409);
or U4780 (N_4780,N_4374,N_4305);
nor U4781 (N_4781,N_4489,N_4284);
nor U4782 (N_4782,N_4370,N_4473);
and U4783 (N_4783,N_4429,N_4380);
nand U4784 (N_4784,N_4092,N_4218);
nand U4785 (N_4785,N_4300,N_4171);
nor U4786 (N_4786,N_4248,N_4230);
or U4787 (N_4787,N_4209,N_4179);
or U4788 (N_4788,N_4048,N_4379);
nor U4789 (N_4789,N_4115,N_4005);
and U4790 (N_4790,N_4050,N_4030);
nor U4791 (N_4791,N_4091,N_4383);
nand U4792 (N_4792,N_4447,N_4054);
nor U4793 (N_4793,N_4147,N_4297);
or U4794 (N_4794,N_4014,N_4074);
nor U4795 (N_4795,N_4394,N_4230);
nor U4796 (N_4796,N_4493,N_4471);
nor U4797 (N_4797,N_4363,N_4309);
or U4798 (N_4798,N_4334,N_4112);
nand U4799 (N_4799,N_4317,N_4418);
nor U4800 (N_4800,N_4357,N_4018);
nor U4801 (N_4801,N_4372,N_4097);
and U4802 (N_4802,N_4292,N_4302);
nand U4803 (N_4803,N_4006,N_4065);
nand U4804 (N_4804,N_4196,N_4035);
nand U4805 (N_4805,N_4065,N_4025);
nand U4806 (N_4806,N_4087,N_4497);
or U4807 (N_4807,N_4015,N_4043);
or U4808 (N_4808,N_4306,N_4154);
or U4809 (N_4809,N_4294,N_4170);
and U4810 (N_4810,N_4435,N_4097);
nand U4811 (N_4811,N_4208,N_4370);
or U4812 (N_4812,N_4241,N_4016);
and U4813 (N_4813,N_4351,N_4221);
nand U4814 (N_4814,N_4399,N_4183);
and U4815 (N_4815,N_4014,N_4033);
and U4816 (N_4816,N_4227,N_4055);
and U4817 (N_4817,N_4069,N_4029);
nand U4818 (N_4818,N_4174,N_4081);
nand U4819 (N_4819,N_4198,N_4100);
nand U4820 (N_4820,N_4412,N_4210);
nand U4821 (N_4821,N_4364,N_4140);
nor U4822 (N_4822,N_4137,N_4077);
nand U4823 (N_4823,N_4254,N_4064);
or U4824 (N_4824,N_4468,N_4074);
and U4825 (N_4825,N_4337,N_4001);
nand U4826 (N_4826,N_4016,N_4166);
or U4827 (N_4827,N_4018,N_4297);
and U4828 (N_4828,N_4048,N_4164);
or U4829 (N_4829,N_4143,N_4070);
nor U4830 (N_4830,N_4339,N_4277);
nand U4831 (N_4831,N_4043,N_4136);
and U4832 (N_4832,N_4446,N_4006);
or U4833 (N_4833,N_4143,N_4442);
or U4834 (N_4834,N_4246,N_4321);
nand U4835 (N_4835,N_4373,N_4120);
and U4836 (N_4836,N_4249,N_4139);
nor U4837 (N_4837,N_4322,N_4125);
and U4838 (N_4838,N_4035,N_4170);
or U4839 (N_4839,N_4291,N_4267);
nor U4840 (N_4840,N_4457,N_4462);
xnor U4841 (N_4841,N_4425,N_4368);
nor U4842 (N_4842,N_4377,N_4046);
nor U4843 (N_4843,N_4265,N_4397);
and U4844 (N_4844,N_4283,N_4387);
or U4845 (N_4845,N_4486,N_4151);
and U4846 (N_4846,N_4490,N_4241);
nand U4847 (N_4847,N_4320,N_4051);
or U4848 (N_4848,N_4440,N_4175);
or U4849 (N_4849,N_4279,N_4402);
nand U4850 (N_4850,N_4223,N_4429);
and U4851 (N_4851,N_4364,N_4444);
nand U4852 (N_4852,N_4208,N_4036);
and U4853 (N_4853,N_4434,N_4380);
and U4854 (N_4854,N_4443,N_4013);
nand U4855 (N_4855,N_4077,N_4463);
and U4856 (N_4856,N_4301,N_4087);
nand U4857 (N_4857,N_4494,N_4486);
nand U4858 (N_4858,N_4148,N_4461);
nor U4859 (N_4859,N_4218,N_4284);
nor U4860 (N_4860,N_4356,N_4480);
or U4861 (N_4861,N_4443,N_4129);
nand U4862 (N_4862,N_4446,N_4494);
xor U4863 (N_4863,N_4308,N_4087);
or U4864 (N_4864,N_4450,N_4352);
nand U4865 (N_4865,N_4271,N_4153);
and U4866 (N_4866,N_4042,N_4341);
nand U4867 (N_4867,N_4456,N_4055);
or U4868 (N_4868,N_4217,N_4279);
and U4869 (N_4869,N_4200,N_4381);
nor U4870 (N_4870,N_4291,N_4229);
or U4871 (N_4871,N_4356,N_4464);
nor U4872 (N_4872,N_4319,N_4111);
and U4873 (N_4873,N_4153,N_4166);
and U4874 (N_4874,N_4284,N_4395);
and U4875 (N_4875,N_4444,N_4131);
and U4876 (N_4876,N_4143,N_4309);
nand U4877 (N_4877,N_4415,N_4197);
and U4878 (N_4878,N_4410,N_4155);
and U4879 (N_4879,N_4143,N_4490);
nor U4880 (N_4880,N_4012,N_4225);
and U4881 (N_4881,N_4381,N_4064);
nor U4882 (N_4882,N_4115,N_4158);
or U4883 (N_4883,N_4181,N_4246);
nand U4884 (N_4884,N_4363,N_4015);
nor U4885 (N_4885,N_4226,N_4156);
nor U4886 (N_4886,N_4382,N_4149);
nor U4887 (N_4887,N_4297,N_4359);
nand U4888 (N_4888,N_4030,N_4054);
or U4889 (N_4889,N_4384,N_4483);
or U4890 (N_4890,N_4466,N_4386);
and U4891 (N_4891,N_4063,N_4335);
nor U4892 (N_4892,N_4328,N_4145);
nor U4893 (N_4893,N_4473,N_4261);
nand U4894 (N_4894,N_4235,N_4385);
nor U4895 (N_4895,N_4382,N_4395);
and U4896 (N_4896,N_4215,N_4091);
nand U4897 (N_4897,N_4487,N_4089);
nand U4898 (N_4898,N_4407,N_4345);
nor U4899 (N_4899,N_4179,N_4287);
or U4900 (N_4900,N_4322,N_4317);
and U4901 (N_4901,N_4076,N_4123);
nor U4902 (N_4902,N_4174,N_4085);
or U4903 (N_4903,N_4137,N_4129);
and U4904 (N_4904,N_4329,N_4347);
nand U4905 (N_4905,N_4091,N_4251);
or U4906 (N_4906,N_4231,N_4434);
and U4907 (N_4907,N_4172,N_4198);
or U4908 (N_4908,N_4348,N_4337);
nand U4909 (N_4909,N_4297,N_4448);
and U4910 (N_4910,N_4355,N_4091);
xnor U4911 (N_4911,N_4228,N_4068);
or U4912 (N_4912,N_4346,N_4288);
and U4913 (N_4913,N_4265,N_4333);
nand U4914 (N_4914,N_4243,N_4361);
nor U4915 (N_4915,N_4413,N_4030);
nor U4916 (N_4916,N_4223,N_4002);
nand U4917 (N_4917,N_4230,N_4351);
and U4918 (N_4918,N_4196,N_4029);
or U4919 (N_4919,N_4190,N_4287);
or U4920 (N_4920,N_4405,N_4128);
or U4921 (N_4921,N_4219,N_4255);
or U4922 (N_4922,N_4010,N_4104);
and U4923 (N_4923,N_4092,N_4471);
or U4924 (N_4924,N_4446,N_4183);
and U4925 (N_4925,N_4108,N_4390);
and U4926 (N_4926,N_4297,N_4492);
and U4927 (N_4927,N_4321,N_4148);
or U4928 (N_4928,N_4101,N_4103);
nand U4929 (N_4929,N_4491,N_4233);
and U4930 (N_4930,N_4131,N_4432);
nor U4931 (N_4931,N_4168,N_4347);
and U4932 (N_4932,N_4317,N_4085);
nand U4933 (N_4933,N_4349,N_4435);
and U4934 (N_4934,N_4210,N_4308);
and U4935 (N_4935,N_4492,N_4091);
nor U4936 (N_4936,N_4041,N_4467);
nor U4937 (N_4937,N_4202,N_4117);
and U4938 (N_4938,N_4147,N_4381);
or U4939 (N_4939,N_4480,N_4333);
nor U4940 (N_4940,N_4272,N_4303);
nand U4941 (N_4941,N_4335,N_4278);
and U4942 (N_4942,N_4061,N_4079);
or U4943 (N_4943,N_4346,N_4336);
or U4944 (N_4944,N_4066,N_4271);
nor U4945 (N_4945,N_4326,N_4283);
or U4946 (N_4946,N_4251,N_4374);
and U4947 (N_4947,N_4223,N_4168);
nand U4948 (N_4948,N_4147,N_4102);
or U4949 (N_4949,N_4240,N_4435);
and U4950 (N_4950,N_4224,N_4163);
or U4951 (N_4951,N_4315,N_4318);
or U4952 (N_4952,N_4347,N_4013);
or U4953 (N_4953,N_4489,N_4454);
or U4954 (N_4954,N_4162,N_4175);
or U4955 (N_4955,N_4470,N_4015);
nor U4956 (N_4956,N_4224,N_4188);
or U4957 (N_4957,N_4272,N_4298);
or U4958 (N_4958,N_4250,N_4118);
nand U4959 (N_4959,N_4187,N_4420);
or U4960 (N_4960,N_4008,N_4386);
nand U4961 (N_4961,N_4489,N_4400);
nor U4962 (N_4962,N_4160,N_4197);
or U4963 (N_4963,N_4450,N_4347);
nand U4964 (N_4964,N_4383,N_4271);
and U4965 (N_4965,N_4225,N_4300);
and U4966 (N_4966,N_4256,N_4084);
nand U4967 (N_4967,N_4166,N_4323);
nor U4968 (N_4968,N_4303,N_4444);
nor U4969 (N_4969,N_4072,N_4444);
nor U4970 (N_4970,N_4271,N_4238);
nand U4971 (N_4971,N_4113,N_4122);
nor U4972 (N_4972,N_4074,N_4312);
or U4973 (N_4973,N_4405,N_4328);
nor U4974 (N_4974,N_4417,N_4317);
nor U4975 (N_4975,N_4099,N_4253);
or U4976 (N_4976,N_4012,N_4180);
or U4977 (N_4977,N_4138,N_4210);
nor U4978 (N_4978,N_4446,N_4122);
nor U4979 (N_4979,N_4240,N_4385);
or U4980 (N_4980,N_4422,N_4033);
and U4981 (N_4981,N_4122,N_4469);
nand U4982 (N_4982,N_4150,N_4389);
and U4983 (N_4983,N_4422,N_4162);
and U4984 (N_4984,N_4167,N_4273);
nand U4985 (N_4985,N_4250,N_4276);
nor U4986 (N_4986,N_4291,N_4099);
nor U4987 (N_4987,N_4461,N_4496);
nand U4988 (N_4988,N_4330,N_4447);
or U4989 (N_4989,N_4367,N_4409);
nor U4990 (N_4990,N_4330,N_4120);
nor U4991 (N_4991,N_4235,N_4204);
and U4992 (N_4992,N_4096,N_4347);
nand U4993 (N_4993,N_4383,N_4050);
or U4994 (N_4994,N_4051,N_4117);
or U4995 (N_4995,N_4137,N_4435);
or U4996 (N_4996,N_4014,N_4061);
nor U4997 (N_4997,N_4025,N_4151);
nor U4998 (N_4998,N_4032,N_4134);
nand U4999 (N_4999,N_4438,N_4295);
nand UO_0 (O_0,N_4545,N_4788);
nand UO_1 (O_1,N_4926,N_4694);
and UO_2 (O_2,N_4904,N_4618);
nand UO_3 (O_3,N_4560,N_4623);
nand UO_4 (O_4,N_4679,N_4999);
nand UO_5 (O_5,N_4707,N_4577);
nor UO_6 (O_6,N_4656,N_4833);
or UO_7 (O_7,N_4581,N_4948);
and UO_8 (O_8,N_4789,N_4663);
nand UO_9 (O_9,N_4959,N_4685);
nor UO_10 (O_10,N_4676,N_4972);
nand UO_11 (O_11,N_4559,N_4633);
and UO_12 (O_12,N_4555,N_4554);
or UO_13 (O_13,N_4681,N_4834);
and UO_14 (O_14,N_4553,N_4645);
and UO_15 (O_15,N_4544,N_4803);
and UO_16 (O_16,N_4539,N_4882);
xnor UO_17 (O_17,N_4701,N_4761);
or UO_18 (O_18,N_4818,N_4911);
or UO_19 (O_19,N_4835,N_4787);
nand UO_20 (O_20,N_4903,N_4712);
or UO_21 (O_21,N_4783,N_4689);
nand UO_22 (O_22,N_4604,N_4859);
nor UO_23 (O_23,N_4868,N_4775);
and UO_24 (O_24,N_4827,N_4897);
nand UO_25 (O_25,N_4507,N_4901);
nand UO_26 (O_26,N_4763,N_4664);
or UO_27 (O_27,N_4905,N_4612);
or UO_28 (O_28,N_4921,N_4639);
or UO_29 (O_29,N_4705,N_4816);
nand UO_30 (O_30,N_4751,N_4806);
and UO_31 (O_31,N_4776,N_4980);
and UO_32 (O_32,N_4831,N_4938);
nand UO_33 (O_33,N_4965,N_4923);
or UO_34 (O_34,N_4884,N_4703);
nor UO_35 (O_35,N_4536,N_4865);
nor UO_36 (O_36,N_4919,N_4608);
nand UO_37 (O_37,N_4771,N_4525);
nand UO_38 (O_38,N_4743,N_4971);
nor UO_39 (O_39,N_4616,N_4768);
nor UO_40 (O_40,N_4651,N_4994);
nor UO_41 (O_41,N_4993,N_4609);
or UO_42 (O_42,N_4836,N_4519);
nand UO_43 (O_43,N_4652,N_4711);
or UO_44 (O_44,N_4590,N_4879);
or UO_45 (O_45,N_4832,N_4774);
nand UO_46 (O_46,N_4632,N_4625);
and UO_47 (O_47,N_4706,N_4671);
nor UO_48 (O_48,N_4702,N_4697);
and UO_49 (O_49,N_4855,N_4801);
or UO_50 (O_50,N_4515,N_4637);
or UO_51 (O_51,N_4951,N_4532);
and UO_52 (O_52,N_4924,N_4682);
and UO_53 (O_53,N_4692,N_4683);
nand UO_54 (O_54,N_4798,N_4728);
or UO_55 (O_55,N_4543,N_4770);
nor UO_56 (O_56,N_4538,N_4819);
or UO_57 (O_57,N_4873,N_4867);
and UO_58 (O_58,N_4860,N_4778);
or UO_59 (O_59,N_4755,N_4760);
or UO_60 (O_60,N_4793,N_4517);
or UO_61 (O_61,N_4635,N_4918);
or UO_62 (O_62,N_4957,N_4826);
xnor UO_63 (O_63,N_4922,N_4857);
nor UO_64 (O_64,N_4622,N_4804);
nand UO_65 (O_65,N_4847,N_4624);
or UO_66 (O_66,N_4546,N_4717);
and UO_67 (O_67,N_4968,N_4841);
or UO_68 (O_68,N_4513,N_4962);
or UO_69 (O_69,N_4933,N_4643);
nor UO_70 (O_70,N_4942,N_4753);
or UO_71 (O_71,N_4662,N_4772);
and UO_72 (O_72,N_4805,N_4665);
nor UO_73 (O_73,N_4666,N_4534);
and UO_74 (O_74,N_4802,N_4878);
and UO_75 (O_75,N_4947,N_4747);
or UO_76 (O_76,N_4790,N_4812);
nand UO_77 (O_77,N_4893,N_4709);
nor UO_78 (O_78,N_4563,N_4907);
and UO_79 (O_79,N_4851,N_4686);
and UO_80 (O_80,N_4784,N_4731);
nor UO_81 (O_81,N_4687,N_4601);
and UO_82 (O_82,N_4529,N_4528);
or UO_83 (O_83,N_4823,N_4571);
nor UO_84 (O_84,N_4883,N_4648);
and UO_85 (O_85,N_4509,N_4605);
nor UO_86 (O_86,N_4750,N_4880);
or UO_87 (O_87,N_4562,N_4892);
nand UO_88 (O_88,N_4874,N_4650);
or UO_89 (O_89,N_4730,N_4973);
and UO_90 (O_90,N_4886,N_4655);
and UO_91 (O_91,N_4729,N_4822);
nor UO_92 (O_92,N_4510,N_4786);
nand UO_93 (O_93,N_4724,N_4738);
or UO_94 (O_94,N_4927,N_4955);
or UO_95 (O_95,N_4673,N_4698);
nor UO_96 (O_96,N_4762,N_4533);
or UO_97 (O_97,N_4896,N_4952);
or UO_98 (O_98,N_4548,N_4912);
nand UO_99 (O_99,N_4654,N_4675);
and UO_100 (O_100,N_4839,N_4591);
and UO_101 (O_101,N_4758,N_4714);
and UO_102 (O_102,N_4735,N_4589);
and UO_103 (O_103,N_4920,N_4766);
and UO_104 (O_104,N_4792,N_4906);
nor UO_105 (O_105,N_4570,N_4785);
nor UO_106 (O_106,N_4757,N_4582);
or UO_107 (O_107,N_4887,N_4986);
nor UO_108 (O_108,N_4902,N_4644);
nand UO_109 (O_109,N_4657,N_4863);
or UO_110 (O_110,N_4628,N_4630);
or UO_111 (O_111,N_4615,N_4889);
xor UO_112 (O_112,N_4592,N_4574);
or UO_113 (O_113,N_4820,N_4984);
nand UO_114 (O_114,N_4696,N_4930);
nand UO_115 (O_115,N_4742,N_4537);
nand UO_116 (O_116,N_4983,N_4815);
and UO_117 (O_117,N_4575,N_4849);
and UO_118 (O_118,N_4708,N_4810);
nand UO_119 (O_119,N_4503,N_4531);
or UO_120 (O_120,N_4749,N_4716);
and UO_121 (O_121,N_4607,N_4721);
or UO_122 (O_122,N_4580,N_4936);
and UO_123 (O_123,N_4521,N_4518);
and UO_124 (O_124,N_4794,N_4916);
nor UO_125 (O_125,N_4995,N_4606);
nand UO_126 (O_126,N_4670,N_4830);
nand UO_127 (O_127,N_4723,N_4547);
and UO_128 (O_128,N_4552,N_4585);
nor UO_129 (O_129,N_4568,N_4595);
or UO_130 (O_130,N_4773,N_4915);
nor UO_131 (O_131,N_4909,N_4726);
or UO_132 (O_132,N_4900,N_4733);
and UO_133 (O_133,N_4985,N_4791);
or UO_134 (O_134,N_4695,N_4727);
or UO_135 (O_135,N_4556,N_4913);
nor UO_136 (O_136,N_4894,N_4780);
or UO_137 (O_137,N_4877,N_4713);
and UO_138 (O_138,N_4501,N_4871);
and UO_139 (O_139,N_4739,N_4514);
nor UO_140 (O_140,N_4808,N_4704);
or UO_141 (O_141,N_4939,N_4576);
nand UO_142 (O_142,N_4541,N_4677);
nand UO_143 (O_143,N_4691,N_4566);
and UO_144 (O_144,N_4987,N_4744);
nor UO_145 (O_145,N_4524,N_4688);
nor UO_146 (O_146,N_4781,N_4958);
nor UO_147 (O_147,N_4549,N_4872);
nand UO_148 (O_148,N_4950,N_4626);
nand UO_149 (O_149,N_4858,N_4535);
and UO_150 (O_150,N_4526,N_4597);
xnor UO_151 (O_151,N_4672,N_4989);
nor UO_152 (O_152,N_4977,N_4557);
or UO_153 (O_153,N_4634,N_4898);
nor UO_154 (O_154,N_4578,N_4891);
or UO_155 (O_155,N_4807,N_4734);
and UO_156 (O_156,N_4573,N_4954);
nor UO_157 (O_157,N_4684,N_4795);
nor UO_158 (O_158,N_4917,N_4963);
nor UO_159 (O_159,N_4504,N_4500);
or UO_160 (O_160,N_4838,N_4602);
nand UO_161 (O_161,N_4854,N_4505);
or UO_162 (O_162,N_4748,N_4956);
or UO_163 (O_163,N_4551,N_4925);
or UO_164 (O_164,N_4719,N_4678);
nor UO_165 (O_165,N_4814,N_4975);
or UO_166 (O_166,N_4653,N_4640);
or UO_167 (O_167,N_4953,N_4611);
and UO_168 (O_168,N_4584,N_4850);
nor UO_169 (O_169,N_4759,N_4564);
or UO_170 (O_170,N_4964,N_4588);
and UO_171 (O_171,N_4991,N_4741);
nor UO_172 (O_172,N_4800,N_4813);
nor UO_173 (O_173,N_4988,N_4944);
nor UO_174 (O_174,N_4558,N_4869);
or UO_175 (O_175,N_4899,N_4565);
and UO_176 (O_176,N_4843,N_4946);
nor UO_177 (O_177,N_4527,N_4567);
or UO_178 (O_178,N_4967,N_4603);
and UO_179 (O_179,N_4797,N_4799);
and UO_180 (O_180,N_4767,N_4636);
or UO_181 (O_181,N_4680,N_4777);
or UO_182 (O_182,N_4572,N_4910);
nor UO_183 (O_183,N_4598,N_4668);
or UO_184 (O_184,N_4523,N_4885);
and UO_185 (O_185,N_4600,N_4979);
nand UO_186 (O_186,N_4508,N_4970);
nor UO_187 (O_187,N_4661,N_4502);
nor UO_188 (O_188,N_4620,N_4737);
and UO_189 (O_189,N_4614,N_4718);
nor UO_190 (O_190,N_4715,N_4875);
or UO_191 (O_191,N_4997,N_4593);
nand UO_192 (O_192,N_4845,N_4914);
nor UO_193 (O_193,N_4961,N_4647);
nor UO_194 (O_194,N_4722,N_4610);
nor UO_195 (O_195,N_4674,N_4736);
nor UO_196 (O_196,N_4725,N_4613);
nand UO_197 (O_197,N_4710,N_4631);
nor UO_198 (O_198,N_4881,N_4829);
nand UO_199 (O_199,N_4649,N_4669);
and UO_200 (O_200,N_4542,N_4745);
or UO_201 (O_201,N_4540,N_4935);
nor UO_202 (O_202,N_4996,N_4779);
nand UO_203 (O_203,N_4516,N_4599);
and UO_204 (O_204,N_4617,N_4929);
nor UO_205 (O_205,N_4828,N_4629);
nand UO_206 (O_206,N_4861,N_4928);
nand UO_207 (O_207,N_4522,N_4811);
and UO_208 (O_208,N_4658,N_4949);
and UO_209 (O_209,N_4732,N_4638);
nor UO_210 (O_210,N_4825,N_4908);
nand UO_211 (O_211,N_4583,N_4876);
nand UO_212 (O_212,N_4943,N_4842);
nor UO_213 (O_213,N_4693,N_4853);
xor UO_214 (O_214,N_4530,N_4866);
nand UO_215 (O_215,N_4756,N_4809);
or UO_216 (O_216,N_4844,N_4667);
nor UO_217 (O_217,N_4506,N_4769);
nor UO_218 (O_218,N_4932,N_4740);
or UO_219 (O_219,N_4945,N_4690);
or UO_220 (O_220,N_4940,N_4837);
nor UO_221 (O_221,N_4782,N_4596);
or UO_222 (O_222,N_4966,N_4550);
nor UO_223 (O_223,N_4990,N_4752);
nand UO_224 (O_224,N_4579,N_4992);
or UO_225 (O_225,N_4998,N_4594);
nor UO_226 (O_226,N_4862,N_4864);
nor UO_227 (O_227,N_4982,N_4659);
and UO_228 (O_228,N_4700,N_4642);
nor UO_229 (O_229,N_4974,N_4646);
and UO_230 (O_230,N_4978,N_4764);
and UO_231 (O_231,N_4621,N_4512);
nand UO_232 (O_232,N_4856,N_4699);
nand UO_233 (O_233,N_4754,N_4848);
and UO_234 (O_234,N_4821,N_4587);
nand UO_235 (O_235,N_4969,N_4890);
nand UO_236 (O_236,N_4569,N_4561);
nand UO_237 (O_237,N_4981,N_4941);
or UO_238 (O_238,N_4976,N_4840);
and UO_239 (O_239,N_4619,N_4586);
and UO_240 (O_240,N_4720,N_4960);
or UO_241 (O_241,N_4846,N_4660);
nor UO_242 (O_242,N_4641,N_4627);
nor UO_243 (O_243,N_4796,N_4937);
nor UO_244 (O_244,N_4765,N_4824);
xnor UO_245 (O_245,N_4934,N_4852);
nor UO_246 (O_246,N_4511,N_4817);
and UO_247 (O_247,N_4895,N_4746);
nor UO_248 (O_248,N_4520,N_4888);
and UO_249 (O_249,N_4931,N_4870);
or UO_250 (O_250,N_4851,N_4681);
nand UO_251 (O_251,N_4525,N_4501);
and UO_252 (O_252,N_4749,N_4506);
and UO_253 (O_253,N_4920,N_4965);
or UO_254 (O_254,N_4538,N_4547);
and UO_255 (O_255,N_4732,N_4949);
nand UO_256 (O_256,N_4841,N_4576);
nand UO_257 (O_257,N_4982,N_4957);
nand UO_258 (O_258,N_4943,N_4817);
nor UO_259 (O_259,N_4896,N_4743);
and UO_260 (O_260,N_4843,N_4608);
and UO_261 (O_261,N_4942,N_4603);
nand UO_262 (O_262,N_4885,N_4963);
or UO_263 (O_263,N_4518,N_4729);
nor UO_264 (O_264,N_4660,N_4723);
nand UO_265 (O_265,N_4604,N_4567);
and UO_266 (O_266,N_4876,N_4766);
nor UO_267 (O_267,N_4720,N_4628);
and UO_268 (O_268,N_4638,N_4628);
nand UO_269 (O_269,N_4766,N_4879);
nand UO_270 (O_270,N_4619,N_4684);
or UO_271 (O_271,N_4784,N_4774);
nor UO_272 (O_272,N_4853,N_4944);
and UO_273 (O_273,N_4879,N_4661);
nor UO_274 (O_274,N_4853,N_4615);
or UO_275 (O_275,N_4979,N_4772);
nand UO_276 (O_276,N_4645,N_4734);
and UO_277 (O_277,N_4899,N_4829);
or UO_278 (O_278,N_4505,N_4889);
nor UO_279 (O_279,N_4846,N_4944);
nand UO_280 (O_280,N_4695,N_4758);
nor UO_281 (O_281,N_4970,N_4539);
or UO_282 (O_282,N_4695,N_4702);
and UO_283 (O_283,N_4503,N_4580);
and UO_284 (O_284,N_4603,N_4779);
and UO_285 (O_285,N_4668,N_4558);
and UO_286 (O_286,N_4916,N_4533);
xor UO_287 (O_287,N_4874,N_4986);
nor UO_288 (O_288,N_4764,N_4722);
or UO_289 (O_289,N_4690,N_4988);
nand UO_290 (O_290,N_4934,N_4823);
or UO_291 (O_291,N_4886,N_4616);
and UO_292 (O_292,N_4611,N_4875);
nand UO_293 (O_293,N_4829,N_4787);
nor UO_294 (O_294,N_4965,N_4558);
and UO_295 (O_295,N_4616,N_4585);
nor UO_296 (O_296,N_4781,N_4695);
and UO_297 (O_297,N_4890,N_4713);
nand UO_298 (O_298,N_4867,N_4766);
nand UO_299 (O_299,N_4777,N_4943);
nor UO_300 (O_300,N_4742,N_4957);
nor UO_301 (O_301,N_4541,N_4706);
nand UO_302 (O_302,N_4619,N_4746);
or UO_303 (O_303,N_4769,N_4800);
and UO_304 (O_304,N_4668,N_4912);
and UO_305 (O_305,N_4579,N_4718);
and UO_306 (O_306,N_4517,N_4588);
nor UO_307 (O_307,N_4582,N_4680);
nor UO_308 (O_308,N_4822,N_4651);
and UO_309 (O_309,N_4850,N_4553);
or UO_310 (O_310,N_4858,N_4949);
or UO_311 (O_311,N_4864,N_4908);
nand UO_312 (O_312,N_4993,N_4566);
nand UO_313 (O_313,N_4779,N_4545);
nand UO_314 (O_314,N_4764,N_4703);
or UO_315 (O_315,N_4992,N_4706);
and UO_316 (O_316,N_4688,N_4638);
nor UO_317 (O_317,N_4557,N_4912);
nor UO_318 (O_318,N_4989,N_4990);
nor UO_319 (O_319,N_4993,N_4884);
nand UO_320 (O_320,N_4525,N_4825);
nand UO_321 (O_321,N_4994,N_4875);
or UO_322 (O_322,N_4545,N_4868);
or UO_323 (O_323,N_4750,N_4792);
and UO_324 (O_324,N_4670,N_4769);
or UO_325 (O_325,N_4510,N_4906);
and UO_326 (O_326,N_4898,N_4934);
or UO_327 (O_327,N_4821,N_4914);
nand UO_328 (O_328,N_4903,N_4937);
and UO_329 (O_329,N_4813,N_4614);
nand UO_330 (O_330,N_4970,N_4874);
and UO_331 (O_331,N_4813,N_4921);
xnor UO_332 (O_332,N_4545,N_4583);
or UO_333 (O_333,N_4835,N_4788);
nand UO_334 (O_334,N_4874,N_4717);
nor UO_335 (O_335,N_4911,N_4874);
or UO_336 (O_336,N_4820,N_4794);
and UO_337 (O_337,N_4607,N_4526);
nand UO_338 (O_338,N_4548,N_4538);
or UO_339 (O_339,N_4575,N_4821);
xnor UO_340 (O_340,N_4665,N_4986);
or UO_341 (O_341,N_4756,N_4798);
nand UO_342 (O_342,N_4988,N_4529);
nand UO_343 (O_343,N_4534,N_4629);
nor UO_344 (O_344,N_4626,N_4735);
and UO_345 (O_345,N_4511,N_4509);
nor UO_346 (O_346,N_4939,N_4861);
and UO_347 (O_347,N_4518,N_4760);
and UO_348 (O_348,N_4588,N_4682);
and UO_349 (O_349,N_4862,N_4663);
nand UO_350 (O_350,N_4751,N_4712);
nor UO_351 (O_351,N_4727,N_4842);
or UO_352 (O_352,N_4586,N_4732);
nor UO_353 (O_353,N_4604,N_4608);
nor UO_354 (O_354,N_4735,N_4728);
or UO_355 (O_355,N_4599,N_4517);
nor UO_356 (O_356,N_4543,N_4533);
nand UO_357 (O_357,N_4596,N_4683);
and UO_358 (O_358,N_4898,N_4907);
and UO_359 (O_359,N_4880,N_4983);
nand UO_360 (O_360,N_4954,N_4891);
or UO_361 (O_361,N_4895,N_4508);
and UO_362 (O_362,N_4587,N_4725);
nor UO_363 (O_363,N_4969,N_4780);
nand UO_364 (O_364,N_4885,N_4692);
nor UO_365 (O_365,N_4582,N_4953);
nor UO_366 (O_366,N_4652,N_4863);
or UO_367 (O_367,N_4653,N_4782);
and UO_368 (O_368,N_4795,N_4712);
or UO_369 (O_369,N_4639,N_4631);
nor UO_370 (O_370,N_4647,N_4889);
and UO_371 (O_371,N_4896,N_4616);
nor UO_372 (O_372,N_4511,N_4636);
nand UO_373 (O_373,N_4600,N_4847);
nand UO_374 (O_374,N_4847,N_4930);
nand UO_375 (O_375,N_4839,N_4580);
or UO_376 (O_376,N_4525,N_4864);
nor UO_377 (O_377,N_4738,N_4672);
xnor UO_378 (O_378,N_4841,N_4619);
nor UO_379 (O_379,N_4945,N_4521);
or UO_380 (O_380,N_4761,N_4506);
or UO_381 (O_381,N_4975,N_4766);
nand UO_382 (O_382,N_4669,N_4575);
or UO_383 (O_383,N_4862,N_4647);
nand UO_384 (O_384,N_4702,N_4710);
or UO_385 (O_385,N_4643,N_4904);
nand UO_386 (O_386,N_4858,N_4637);
nor UO_387 (O_387,N_4884,N_4637);
nand UO_388 (O_388,N_4732,N_4832);
nand UO_389 (O_389,N_4773,N_4595);
nand UO_390 (O_390,N_4722,N_4672);
xnor UO_391 (O_391,N_4789,N_4555);
and UO_392 (O_392,N_4626,N_4784);
nor UO_393 (O_393,N_4983,N_4852);
nor UO_394 (O_394,N_4883,N_4573);
or UO_395 (O_395,N_4892,N_4745);
nand UO_396 (O_396,N_4938,N_4960);
nand UO_397 (O_397,N_4846,N_4528);
nand UO_398 (O_398,N_4580,N_4690);
and UO_399 (O_399,N_4981,N_4926);
nor UO_400 (O_400,N_4638,N_4997);
or UO_401 (O_401,N_4627,N_4700);
and UO_402 (O_402,N_4934,N_4717);
and UO_403 (O_403,N_4811,N_4621);
nor UO_404 (O_404,N_4542,N_4834);
and UO_405 (O_405,N_4521,N_4587);
and UO_406 (O_406,N_4652,N_4671);
and UO_407 (O_407,N_4969,N_4829);
or UO_408 (O_408,N_4712,N_4610);
nand UO_409 (O_409,N_4920,N_4641);
or UO_410 (O_410,N_4827,N_4788);
nand UO_411 (O_411,N_4603,N_4637);
nand UO_412 (O_412,N_4582,N_4738);
nand UO_413 (O_413,N_4634,N_4754);
and UO_414 (O_414,N_4612,N_4932);
and UO_415 (O_415,N_4632,N_4876);
nand UO_416 (O_416,N_4785,N_4896);
or UO_417 (O_417,N_4528,N_4791);
nand UO_418 (O_418,N_4962,N_4607);
nor UO_419 (O_419,N_4897,N_4692);
nand UO_420 (O_420,N_4837,N_4831);
xor UO_421 (O_421,N_4502,N_4642);
nand UO_422 (O_422,N_4615,N_4521);
and UO_423 (O_423,N_4649,N_4500);
nor UO_424 (O_424,N_4521,N_4721);
and UO_425 (O_425,N_4881,N_4918);
nand UO_426 (O_426,N_4796,N_4874);
nand UO_427 (O_427,N_4795,N_4580);
nor UO_428 (O_428,N_4641,N_4553);
nand UO_429 (O_429,N_4897,N_4643);
nor UO_430 (O_430,N_4679,N_4639);
nand UO_431 (O_431,N_4899,N_4796);
nor UO_432 (O_432,N_4937,N_4815);
nand UO_433 (O_433,N_4990,N_4675);
nor UO_434 (O_434,N_4671,N_4828);
nand UO_435 (O_435,N_4774,N_4604);
and UO_436 (O_436,N_4692,N_4671);
nor UO_437 (O_437,N_4860,N_4622);
nand UO_438 (O_438,N_4641,N_4904);
nand UO_439 (O_439,N_4541,N_4857);
nor UO_440 (O_440,N_4634,N_4918);
nor UO_441 (O_441,N_4890,N_4758);
or UO_442 (O_442,N_4992,N_4912);
nor UO_443 (O_443,N_4933,N_4858);
nor UO_444 (O_444,N_4753,N_4565);
or UO_445 (O_445,N_4899,N_4925);
nand UO_446 (O_446,N_4771,N_4576);
or UO_447 (O_447,N_4739,N_4542);
and UO_448 (O_448,N_4773,N_4549);
nand UO_449 (O_449,N_4664,N_4945);
nand UO_450 (O_450,N_4537,N_4712);
and UO_451 (O_451,N_4528,N_4591);
or UO_452 (O_452,N_4799,N_4558);
nand UO_453 (O_453,N_4823,N_4727);
nand UO_454 (O_454,N_4606,N_4828);
nand UO_455 (O_455,N_4991,N_4940);
nor UO_456 (O_456,N_4963,N_4548);
nand UO_457 (O_457,N_4638,N_4955);
or UO_458 (O_458,N_4518,N_4771);
and UO_459 (O_459,N_4610,N_4632);
or UO_460 (O_460,N_4901,N_4823);
or UO_461 (O_461,N_4923,N_4599);
nand UO_462 (O_462,N_4883,N_4911);
xor UO_463 (O_463,N_4594,N_4827);
or UO_464 (O_464,N_4534,N_4718);
nand UO_465 (O_465,N_4719,N_4796);
nor UO_466 (O_466,N_4536,N_4528);
nand UO_467 (O_467,N_4916,N_4593);
nand UO_468 (O_468,N_4757,N_4967);
nand UO_469 (O_469,N_4809,N_4912);
nor UO_470 (O_470,N_4626,N_4863);
or UO_471 (O_471,N_4536,N_4818);
nand UO_472 (O_472,N_4520,N_4781);
or UO_473 (O_473,N_4730,N_4663);
nor UO_474 (O_474,N_4895,N_4683);
and UO_475 (O_475,N_4891,N_4598);
nor UO_476 (O_476,N_4944,N_4632);
nand UO_477 (O_477,N_4577,N_4639);
nand UO_478 (O_478,N_4803,N_4662);
nor UO_479 (O_479,N_4587,N_4731);
nand UO_480 (O_480,N_4868,N_4652);
nor UO_481 (O_481,N_4773,N_4632);
nor UO_482 (O_482,N_4523,N_4558);
or UO_483 (O_483,N_4801,N_4550);
nand UO_484 (O_484,N_4728,N_4918);
nand UO_485 (O_485,N_4869,N_4980);
nor UO_486 (O_486,N_4775,N_4671);
nor UO_487 (O_487,N_4922,N_4946);
nand UO_488 (O_488,N_4859,N_4827);
nand UO_489 (O_489,N_4761,N_4881);
and UO_490 (O_490,N_4838,N_4756);
nor UO_491 (O_491,N_4796,N_4970);
nor UO_492 (O_492,N_4907,N_4867);
nand UO_493 (O_493,N_4606,N_4633);
or UO_494 (O_494,N_4862,N_4767);
and UO_495 (O_495,N_4944,N_4935);
nor UO_496 (O_496,N_4874,N_4931);
or UO_497 (O_497,N_4556,N_4974);
nand UO_498 (O_498,N_4726,N_4648);
or UO_499 (O_499,N_4887,N_4634);
and UO_500 (O_500,N_4975,N_4926);
nor UO_501 (O_501,N_4579,N_4894);
nand UO_502 (O_502,N_4886,N_4570);
or UO_503 (O_503,N_4554,N_4773);
nand UO_504 (O_504,N_4955,N_4842);
and UO_505 (O_505,N_4727,N_4618);
and UO_506 (O_506,N_4976,N_4592);
nor UO_507 (O_507,N_4619,N_4871);
nand UO_508 (O_508,N_4719,N_4790);
or UO_509 (O_509,N_4801,N_4854);
nor UO_510 (O_510,N_4980,N_4778);
nor UO_511 (O_511,N_4572,N_4582);
nor UO_512 (O_512,N_4959,N_4662);
nor UO_513 (O_513,N_4579,N_4668);
or UO_514 (O_514,N_4917,N_4854);
and UO_515 (O_515,N_4748,N_4808);
or UO_516 (O_516,N_4592,N_4545);
nor UO_517 (O_517,N_4700,N_4503);
or UO_518 (O_518,N_4556,N_4672);
and UO_519 (O_519,N_4674,N_4864);
nor UO_520 (O_520,N_4779,N_4906);
or UO_521 (O_521,N_4909,N_4522);
or UO_522 (O_522,N_4600,N_4801);
and UO_523 (O_523,N_4837,N_4994);
or UO_524 (O_524,N_4646,N_4761);
nor UO_525 (O_525,N_4789,N_4635);
and UO_526 (O_526,N_4881,N_4906);
nor UO_527 (O_527,N_4907,N_4583);
and UO_528 (O_528,N_4658,N_4595);
or UO_529 (O_529,N_4669,N_4984);
nand UO_530 (O_530,N_4680,N_4866);
and UO_531 (O_531,N_4906,N_4841);
or UO_532 (O_532,N_4505,N_4744);
nor UO_533 (O_533,N_4594,N_4634);
and UO_534 (O_534,N_4547,N_4604);
and UO_535 (O_535,N_4984,N_4909);
nor UO_536 (O_536,N_4860,N_4983);
and UO_537 (O_537,N_4953,N_4858);
nand UO_538 (O_538,N_4687,N_4988);
nand UO_539 (O_539,N_4737,N_4962);
and UO_540 (O_540,N_4646,N_4855);
or UO_541 (O_541,N_4682,N_4902);
nand UO_542 (O_542,N_4989,N_4663);
or UO_543 (O_543,N_4767,N_4906);
and UO_544 (O_544,N_4946,N_4637);
and UO_545 (O_545,N_4756,N_4565);
or UO_546 (O_546,N_4508,N_4600);
and UO_547 (O_547,N_4921,N_4946);
nand UO_548 (O_548,N_4525,N_4571);
and UO_549 (O_549,N_4610,N_4612);
and UO_550 (O_550,N_4899,N_4948);
and UO_551 (O_551,N_4774,N_4933);
nor UO_552 (O_552,N_4797,N_4764);
nor UO_553 (O_553,N_4683,N_4703);
nand UO_554 (O_554,N_4552,N_4626);
nand UO_555 (O_555,N_4593,N_4553);
and UO_556 (O_556,N_4935,N_4714);
or UO_557 (O_557,N_4563,N_4610);
and UO_558 (O_558,N_4667,N_4599);
nand UO_559 (O_559,N_4800,N_4740);
xnor UO_560 (O_560,N_4908,N_4787);
and UO_561 (O_561,N_4604,N_4706);
nor UO_562 (O_562,N_4735,N_4609);
and UO_563 (O_563,N_4761,N_4513);
nand UO_564 (O_564,N_4904,N_4986);
nor UO_565 (O_565,N_4983,N_4947);
nor UO_566 (O_566,N_4897,N_4789);
nand UO_567 (O_567,N_4650,N_4602);
nor UO_568 (O_568,N_4693,N_4660);
nor UO_569 (O_569,N_4926,N_4955);
and UO_570 (O_570,N_4625,N_4662);
or UO_571 (O_571,N_4586,N_4596);
nand UO_572 (O_572,N_4889,N_4703);
nor UO_573 (O_573,N_4717,N_4889);
nand UO_574 (O_574,N_4685,N_4705);
nor UO_575 (O_575,N_4757,N_4953);
nor UO_576 (O_576,N_4997,N_4950);
and UO_577 (O_577,N_4503,N_4706);
nand UO_578 (O_578,N_4926,N_4635);
or UO_579 (O_579,N_4907,N_4689);
nand UO_580 (O_580,N_4896,N_4682);
or UO_581 (O_581,N_4805,N_4840);
nor UO_582 (O_582,N_4849,N_4937);
nand UO_583 (O_583,N_4537,N_4918);
or UO_584 (O_584,N_4928,N_4814);
nand UO_585 (O_585,N_4899,N_4955);
or UO_586 (O_586,N_4888,N_4649);
nor UO_587 (O_587,N_4994,N_4726);
nand UO_588 (O_588,N_4864,N_4721);
and UO_589 (O_589,N_4690,N_4636);
or UO_590 (O_590,N_4994,N_4722);
or UO_591 (O_591,N_4861,N_4812);
nor UO_592 (O_592,N_4549,N_4885);
nor UO_593 (O_593,N_4967,N_4764);
nand UO_594 (O_594,N_4885,N_4952);
nand UO_595 (O_595,N_4654,N_4988);
nand UO_596 (O_596,N_4718,N_4631);
nand UO_597 (O_597,N_4826,N_4597);
xor UO_598 (O_598,N_4930,N_4691);
nand UO_599 (O_599,N_4910,N_4538);
and UO_600 (O_600,N_4825,N_4927);
nand UO_601 (O_601,N_4876,N_4936);
nand UO_602 (O_602,N_4923,N_4676);
and UO_603 (O_603,N_4916,N_4946);
nand UO_604 (O_604,N_4772,N_4803);
nor UO_605 (O_605,N_4517,N_4918);
nand UO_606 (O_606,N_4538,N_4977);
nand UO_607 (O_607,N_4623,N_4818);
nand UO_608 (O_608,N_4978,N_4828);
xor UO_609 (O_609,N_4672,N_4688);
and UO_610 (O_610,N_4946,N_4821);
nor UO_611 (O_611,N_4915,N_4825);
nand UO_612 (O_612,N_4529,N_4673);
or UO_613 (O_613,N_4888,N_4983);
or UO_614 (O_614,N_4627,N_4816);
or UO_615 (O_615,N_4624,N_4896);
and UO_616 (O_616,N_4597,N_4562);
and UO_617 (O_617,N_4736,N_4706);
or UO_618 (O_618,N_4526,N_4652);
nor UO_619 (O_619,N_4964,N_4678);
and UO_620 (O_620,N_4666,N_4793);
nand UO_621 (O_621,N_4926,N_4999);
nand UO_622 (O_622,N_4703,N_4958);
or UO_623 (O_623,N_4777,N_4915);
nand UO_624 (O_624,N_4501,N_4629);
nand UO_625 (O_625,N_4934,N_4661);
xor UO_626 (O_626,N_4671,N_4864);
nor UO_627 (O_627,N_4803,N_4504);
or UO_628 (O_628,N_4568,N_4615);
nand UO_629 (O_629,N_4960,N_4940);
and UO_630 (O_630,N_4984,N_4730);
or UO_631 (O_631,N_4717,N_4854);
nand UO_632 (O_632,N_4754,N_4612);
nor UO_633 (O_633,N_4677,N_4996);
or UO_634 (O_634,N_4755,N_4947);
nor UO_635 (O_635,N_4795,N_4595);
nor UO_636 (O_636,N_4968,N_4906);
and UO_637 (O_637,N_4774,N_4821);
nand UO_638 (O_638,N_4996,N_4700);
or UO_639 (O_639,N_4576,N_4716);
and UO_640 (O_640,N_4631,N_4745);
nand UO_641 (O_641,N_4804,N_4737);
and UO_642 (O_642,N_4908,N_4518);
nor UO_643 (O_643,N_4632,N_4788);
nand UO_644 (O_644,N_4714,N_4981);
or UO_645 (O_645,N_4807,N_4822);
nor UO_646 (O_646,N_4513,N_4663);
nand UO_647 (O_647,N_4808,N_4503);
or UO_648 (O_648,N_4665,N_4897);
nand UO_649 (O_649,N_4852,N_4567);
nand UO_650 (O_650,N_4774,N_4801);
nor UO_651 (O_651,N_4716,N_4510);
xnor UO_652 (O_652,N_4968,N_4525);
or UO_653 (O_653,N_4788,N_4959);
nor UO_654 (O_654,N_4680,N_4992);
and UO_655 (O_655,N_4943,N_4980);
nor UO_656 (O_656,N_4896,N_4651);
nor UO_657 (O_657,N_4605,N_4765);
or UO_658 (O_658,N_4985,N_4989);
and UO_659 (O_659,N_4729,N_4883);
and UO_660 (O_660,N_4545,N_4889);
or UO_661 (O_661,N_4549,N_4709);
and UO_662 (O_662,N_4566,N_4660);
and UO_663 (O_663,N_4965,N_4544);
nand UO_664 (O_664,N_4746,N_4876);
nor UO_665 (O_665,N_4927,N_4939);
nand UO_666 (O_666,N_4699,N_4503);
nand UO_667 (O_667,N_4613,N_4994);
and UO_668 (O_668,N_4632,N_4721);
nand UO_669 (O_669,N_4722,N_4951);
nor UO_670 (O_670,N_4852,N_4864);
or UO_671 (O_671,N_4559,N_4861);
nand UO_672 (O_672,N_4528,N_4680);
nand UO_673 (O_673,N_4827,N_4940);
and UO_674 (O_674,N_4554,N_4941);
or UO_675 (O_675,N_4956,N_4996);
or UO_676 (O_676,N_4584,N_4980);
or UO_677 (O_677,N_4853,N_4974);
nand UO_678 (O_678,N_4627,N_4716);
or UO_679 (O_679,N_4633,N_4616);
nor UO_680 (O_680,N_4685,N_4669);
or UO_681 (O_681,N_4935,N_4979);
nor UO_682 (O_682,N_4703,N_4724);
nand UO_683 (O_683,N_4951,N_4906);
nor UO_684 (O_684,N_4583,N_4697);
and UO_685 (O_685,N_4948,N_4504);
and UO_686 (O_686,N_4531,N_4819);
or UO_687 (O_687,N_4744,N_4673);
and UO_688 (O_688,N_4841,N_4965);
and UO_689 (O_689,N_4826,N_4601);
and UO_690 (O_690,N_4884,N_4538);
nand UO_691 (O_691,N_4861,N_4751);
or UO_692 (O_692,N_4965,N_4884);
and UO_693 (O_693,N_4738,N_4737);
nand UO_694 (O_694,N_4680,N_4697);
and UO_695 (O_695,N_4773,N_4783);
nand UO_696 (O_696,N_4573,N_4866);
and UO_697 (O_697,N_4916,N_4650);
nor UO_698 (O_698,N_4609,N_4851);
nor UO_699 (O_699,N_4608,N_4861);
nor UO_700 (O_700,N_4605,N_4922);
nor UO_701 (O_701,N_4584,N_4852);
nor UO_702 (O_702,N_4573,N_4747);
and UO_703 (O_703,N_4730,N_4616);
nor UO_704 (O_704,N_4687,N_4564);
nand UO_705 (O_705,N_4990,N_4740);
nor UO_706 (O_706,N_4675,N_4515);
and UO_707 (O_707,N_4725,N_4843);
nand UO_708 (O_708,N_4649,N_4581);
nor UO_709 (O_709,N_4629,N_4746);
and UO_710 (O_710,N_4903,N_4651);
and UO_711 (O_711,N_4706,N_4921);
nor UO_712 (O_712,N_4784,N_4974);
and UO_713 (O_713,N_4795,N_4752);
or UO_714 (O_714,N_4687,N_4590);
nand UO_715 (O_715,N_4522,N_4623);
and UO_716 (O_716,N_4689,N_4754);
nand UO_717 (O_717,N_4538,N_4625);
and UO_718 (O_718,N_4685,N_4718);
or UO_719 (O_719,N_4744,N_4972);
nor UO_720 (O_720,N_4961,N_4859);
nor UO_721 (O_721,N_4864,N_4798);
and UO_722 (O_722,N_4772,N_4729);
or UO_723 (O_723,N_4715,N_4645);
and UO_724 (O_724,N_4684,N_4509);
and UO_725 (O_725,N_4967,N_4796);
and UO_726 (O_726,N_4646,N_4746);
or UO_727 (O_727,N_4529,N_4971);
nand UO_728 (O_728,N_4975,N_4532);
nand UO_729 (O_729,N_4655,N_4902);
nand UO_730 (O_730,N_4661,N_4573);
nand UO_731 (O_731,N_4835,N_4892);
and UO_732 (O_732,N_4869,N_4989);
nand UO_733 (O_733,N_4754,N_4780);
and UO_734 (O_734,N_4728,N_4994);
nor UO_735 (O_735,N_4552,N_4763);
or UO_736 (O_736,N_4924,N_4958);
and UO_737 (O_737,N_4961,N_4832);
nand UO_738 (O_738,N_4855,N_4753);
nor UO_739 (O_739,N_4729,N_4621);
or UO_740 (O_740,N_4819,N_4895);
and UO_741 (O_741,N_4991,N_4658);
nor UO_742 (O_742,N_4979,N_4863);
nand UO_743 (O_743,N_4521,N_4558);
or UO_744 (O_744,N_4745,N_4808);
or UO_745 (O_745,N_4934,N_4822);
and UO_746 (O_746,N_4996,N_4980);
nand UO_747 (O_747,N_4507,N_4847);
nand UO_748 (O_748,N_4975,N_4634);
and UO_749 (O_749,N_4721,N_4831);
nor UO_750 (O_750,N_4838,N_4640);
nor UO_751 (O_751,N_4595,N_4764);
nand UO_752 (O_752,N_4679,N_4772);
or UO_753 (O_753,N_4801,N_4844);
nand UO_754 (O_754,N_4750,N_4975);
nor UO_755 (O_755,N_4555,N_4540);
nand UO_756 (O_756,N_4843,N_4545);
nor UO_757 (O_757,N_4974,N_4791);
or UO_758 (O_758,N_4505,N_4798);
nor UO_759 (O_759,N_4916,N_4800);
or UO_760 (O_760,N_4877,N_4880);
and UO_761 (O_761,N_4638,N_4949);
or UO_762 (O_762,N_4995,N_4740);
nand UO_763 (O_763,N_4968,N_4797);
and UO_764 (O_764,N_4617,N_4775);
and UO_765 (O_765,N_4500,N_4651);
nand UO_766 (O_766,N_4939,N_4637);
or UO_767 (O_767,N_4793,N_4680);
or UO_768 (O_768,N_4527,N_4987);
or UO_769 (O_769,N_4590,N_4507);
nand UO_770 (O_770,N_4814,N_4878);
nor UO_771 (O_771,N_4583,N_4524);
and UO_772 (O_772,N_4568,N_4581);
nor UO_773 (O_773,N_4857,N_4724);
or UO_774 (O_774,N_4622,N_4923);
nand UO_775 (O_775,N_4511,N_4983);
nor UO_776 (O_776,N_4783,N_4997);
or UO_777 (O_777,N_4592,N_4511);
or UO_778 (O_778,N_4889,N_4746);
nand UO_779 (O_779,N_4591,N_4834);
or UO_780 (O_780,N_4989,N_4683);
or UO_781 (O_781,N_4919,N_4616);
nor UO_782 (O_782,N_4909,N_4615);
nor UO_783 (O_783,N_4790,N_4593);
and UO_784 (O_784,N_4791,N_4817);
nor UO_785 (O_785,N_4981,N_4879);
nand UO_786 (O_786,N_4623,N_4757);
nand UO_787 (O_787,N_4751,N_4645);
or UO_788 (O_788,N_4551,N_4955);
nand UO_789 (O_789,N_4561,N_4977);
or UO_790 (O_790,N_4719,N_4873);
and UO_791 (O_791,N_4873,N_4686);
and UO_792 (O_792,N_4978,N_4936);
or UO_793 (O_793,N_4987,N_4722);
nor UO_794 (O_794,N_4942,N_4654);
and UO_795 (O_795,N_4948,N_4789);
or UO_796 (O_796,N_4609,N_4513);
nand UO_797 (O_797,N_4761,N_4975);
or UO_798 (O_798,N_4512,N_4949);
nor UO_799 (O_799,N_4532,N_4833);
nand UO_800 (O_800,N_4789,N_4747);
and UO_801 (O_801,N_4781,N_4516);
nand UO_802 (O_802,N_4531,N_4594);
and UO_803 (O_803,N_4777,N_4999);
or UO_804 (O_804,N_4524,N_4968);
and UO_805 (O_805,N_4515,N_4987);
and UO_806 (O_806,N_4526,N_4746);
nor UO_807 (O_807,N_4680,N_4553);
nor UO_808 (O_808,N_4699,N_4974);
nor UO_809 (O_809,N_4921,N_4894);
nor UO_810 (O_810,N_4742,N_4574);
and UO_811 (O_811,N_4759,N_4663);
and UO_812 (O_812,N_4865,N_4545);
or UO_813 (O_813,N_4557,N_4994);
nor UO_814 (O_814,N_4662,N_4516);
nand UO_815 (O_815,N_4578,N_4870);
nand UO_816 (O_816,N_4742,N_4863);
nand UO_817 (O_817,N_4708,N_4978);
and UO_818 (O_818,N_4512,N_4685);
or UO_819 (O_819,N_4983,N_4735);
nor UO_820 (O_820,N_4933,N_4579);
nor UO_821 (O_821,N_4862,N_4795);
nand UO_822 (O_822,N_4745,N_4881);
nor UO_823 (O_823,N_4810,N_4508);
nor UO_824 (O_824,N_4786,N_4720);
or UO_825 (O_825,N_4744,N_4808);
and UO_826 (O_826,N_4749,N_4654);
nor UO_827 (O_827,N_4668,N_4500);
nand UO_828 (O_828,N_4768,N_4518);
or UO_829 (O_829,N_4911,N_4984);
or UO_830 (O_830,N_4681,N_4747);
or UO_831 (O_831,N_4784,N_4577);
nand UO_832 (O_832,N_4983,N_4949);
or UO_833 (O_833,N_4740,N_4885);
nor UO_834 (O_834,N_4998,N_4507);
or UO_835 (O_835,N_4819,N_4928);
nor UO_836 (O_836,N_4692,N_4922);
or UO_837 (O_837,N_4903,N_4661);
or UO_838 (O_838,N_4657,N_4792);
nor UO_839 (O_839,N_4791,N_4834);
nor UO_840 (O_840,N_4981,N_4794);
nand UO_841 (O_841,N_4977,N_4639);
nand UO_842 (O_842,N_4640,N_4836);
nor UO_843 (O_843,N_4768,N_4937);
nand UO_844 (O_844,N_4673,N_4767);
nor UO_845 (O_845,N_4733,N_4931);
nor UO_846 (O_846,N_4550,N_4542);
nand UO_847 (O_847,N_4671,N_4973);
and UO_848 (O_848,N_4838,N_4962);
and UO_849 (O_849,N_4906,N_4940);
or UO_850 (O_850,N_4640,N_4631);
or UO_851 (O_851,N_4502,N_4881);
nand UO_852 (O_852,N_4592,N_4869);
nand UO_853 (O_853,N_4635,N_4698);
and UO_854 (O_854,N_4896,N_4531);
and UO_855 (O_855,N_4911,N_4971);
or UO_856 (O_856,N_4531,N_4624);
or UO_857 (O_857,N_4749,N_4679);
and UO_858 (O_858,N_4663,N_4807);
or UO_859 (O_859,N_4722,N_4772);
nor UO_860 (O_860,N_4987,N_4697);
or UO_861 (O_861,N_4908,N_4971);
nor UO_862 (O_862,N_4934,N_4994);
and UO_863 (O_863,N_4655,N_4630);
nand UO_864 (O_864,N_4957,N_4867);
and UO_865 (O_865,N_4647,N_4643);
nand UO_866 (O_866,N_4793,N_4780);
nor UO_867 (O_867,N_4926,N_4695);
nor UO_868 (O_868,N_4771,N_4568);
or UO_869 (O_869,N_4915,N_4554);
and UO_870 (O_870,N_4919,N_4750);
nand UO_871 (O_871,N_4614,N_4565);
nand UO_872 (O_872,N_4763,N_4561);
or UO_873 (O_873,N_4962,N_4567);
or UO_874 (O_874,N_4811,N_4917);
nand UO_875 (O_875,N_4787,N_4664);
nand UO_876 (O_876,N_4715,N_4908);
nand UO_877 (O_877,N_4776,N_4791);
nand UO_878 (O_878,N_4853,N_4673);
nand UO_879 (O_879,N_4586,N_4708);
and UO_880 (O_880,N_4667,N_4526);
nor UO_881 (O_881,N_4509,N_4772);
and UO_882 (O_882,N_4550,N_4795);
nand UO_883 (O_883,N_4702,N_4892);
or UO_884 (O_884,N_4581,N_4645);
nor UO_885 (O_885,N_4884,N_4809);
nand UO_886 (O_886,N_4719,N_4895);
nor UO_887 (O_887,N_4910,N_4564);
or UO_888 (O_888,N_4985,N_4959);
and UO_889 (O_889,N_4740,N_4653);
nand UO_890 (O_890,N_4779,N_4803);
or UO_891 (O_891,N_4679,N_4838);
xor UO_892 (O_892,N_4941,N_4849);
nor UO_893 (O_893,N_4582,N_4514);
nand UO_894 (O_894,N_4794,N_4731);
nand UO_895 (O_895,N_4521,N_4841);
xnor UO_896 (O_896,N_4802,N_4788);
and UO_897 (O_897,N_4568,N_4540);
or UO_898 (O_898,N_4931,N_4916);
or UO_899 (O_899,N_4924,N_4788);
nand UO_900 (O_900,N_4692,N_4755);
nor UO_901 (O_901,N_4804,N_4878);
and UO_902 (O_902,N_4671,N_4704);
nor UO_903 (O_903,N_4596,N_4627);
nor UO_904 (O_904,N_4766,N_4629);
and UO_905 (O_905,N_4754,N_4755);
nor UO_906 (O_906,N_4868,N_4576);
or UO_907 (O_907,N_4667,N_4967);
or UO_908 (O_908,N_4927,N_4603);
nor UO_909 (O_909,N_4836,N_4931);
or UO_910 (O_910,N_4835,N_4674);
and UO_911 (O_911,N_4895,N_4860);
or UO_912 (O_912,N_4814,N_4953);
or UO_913 (O_913,N_4940,N_4521);
or UO_914 (O_914,N_4545,N_4748);
nor UO_915 (O_915,N_4669,N_4629);
xnor UO_916 (O_916,N_4509,N_4850);
nand UO_917 (O_917,N_4711,N_4606);
and UO_918 (O_918,N_4665,N_4648);
and UO_919 (O_919,N_4953,N_4939);
or UO_920 (O_920,N_4912,N_4812);
nor UO_921 (O_921,N_4510,N_4856);
or UO_922 (O_922,N_4500,N_4955);
and UO_923 (O_923,N_4517,N_4864);
and UO_924 (O_924,N_4729,N_4741);
nand UO_925 (O_925,N_4700,N_4570);
nand UO_926 (O_926,N_4887,N_4984);
nor UO_927 (O_927,N_4501,N_4755);
and UO_928 (O_928,N_4838,N_4798);
and UO_929 (O_929,N_4611,N_4844);
and UO_930 (O_930,N_4713,N_4981);
nand UO_931 (O_931,N_4917,N_4531);
nor UO_932 (O_932,N_4940,N_4691);
or UO_933 (O_933,N_4589,N_4928);
nor UO_934 (O_934,N_4932,N_4733);
nor UO_935 (O_935,N_4840,N_4510);
xnor UO_936 (O_936,N_4844,N_4843);
and UO_937 (O_937,N_4817,N_4728);
nand UO_938 (O_938,N_4895,N_4876);
and UO_939 (O_939,N_4533,N_4571);
and UO_940 (O_940,N_4996,N_4755);
nor UO_941 (O_941,N_4941,N_4922);
or UO_942 (O_942,N_4871,N_4940);
and UO_943 (O_943,N_4647,N_4916);
nor UO_944 (O_944,N_4764,N_4798);
and UO_945 (O_945,N_4746,N_4992);
nor UO_946 (O_946,N_4670,N_4726);
nor UO_947 (O_947,N_4629,N_4957);
and UO_948 (O_948,N_4563,N_4712);
nor UO_949 (O_949,N_4986,N_4556);
and UO_950 (O_950,N_4942,N_4762);
and UO_951 (O_951,N_4864,N_4810);
nor UO_952 (O_952,N_4632,N_4874);
and UO_953 (O_953,N_4961,N_4962);
nand UO_954 (O_954,N_4646,N_4573);
nand UO_955 (O_955,N_4961,N_4814);
or UO_956 (O_956,N_4818,N_4851);
nand UO_957 (O_957,N_4637,N_4739);
nand UO_958 (O_958,N_4552,N_4668);
and UO_959 (O_959,N_4726,N_4906);
or UO_960 (O_960,N_4517,N_4809);
or UO_961 (O_961,N_4887,N_4780);
nor UO_962 (O_962,N_4870,N_4672);
and UO_963 (O_963,N_4869,N_4730);
nor UO_964 (O_964,N_4591,N_4845);
xor UO_965 (O_965,N_4786,N_4544);
or UO_966 (O_966,N_4900,N_4626);
nand UO_967 (O_967,N_4808,N_4801);
nand UO_968 (O_968,N_4968,N_4582);
nor UO_969 (O_969,N_4655,N_4674);
or UO_970 (O_970,N_4615,N_4867);
nand UO_971 (O_971,N_4559,N_4596);
nor UO_972 (O_972,N_4595,N_4936);
or UO_973 (O_973,N_4991,N_4666);
nand UO_974 (O_974,N_4556,N_4825);
nand UO_975 (O_975,N_4555,N_4641);
or UO_976 (O_976,N_4762,N_4715);
nor UO_977 (O_977,N_4642,N_4553);
nor UO_978 (O_978,N_4837,N_4567);
nor UO_979 (O_979,N_4917,N_4736);
and UO_980 (O_980,N_4708,N_4686);
nand UO_981 (O_981,N_4623,N_4636);
nor UO_982 (O_982,N_4709,N_4723);
and UO_983 (O_983,N_4804,N_4707);
and UO_984 (O_984,N_4593,N_4830);
or UO_985 (O_985,N_4536,N_4731);
or UO_986 (O_986,N_4608,N_4675);
or UO_987 (O_987,N_4607,N_4890);
or UO_988 (O_988,N_4547,N_4797);
and UO_989 (O_989,N_4873,N_4882);
or UO_990 (O_990,N_4603,N_4502);
nor UO_991 (O_991,N_4683,N_4802);
and UO_992 (O_992,N_4646,N_4586);
and UO_993 (O_993,N_4596,N_4793);
and UO_994 (O_994,N_4832,N_4626);
nand UO_995 (O_995,N_4756,N_4672);
and UO_996 (O_996,N_4758,N_4816);
nor UO_997 (O_997,N_4733,N_4923);
nor UO_998 (O_998,N_4537,N_4722);
nor UO_999 (O_999,N_4604,N_4537);
endmodule