module basic_2000_20000_2500_4_levels_10xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
nand U0 (N_0,In_1582,In_921);
xor U1 (N_1,In_1143,In_1992);
nand U2 (N_2,In_631,In_427);
xor U3 (N_3,In_825,In_1394);
and U4 (N_4,In_1431,In_1270);
nand U5 (N_5,In_221,In_1997);
or U6 (N_6,In_562,In_176);
nand U7 (N_7,In_7,In_367);
nor U8 (N_8,In_891,In_1730);
or U9 (N_9,In_1037,In_775);
xnor U10 (N_10,In_502,In_1441);
and U11 (N_11,In_766,In_1468);
or U12 (N_12,In_1741,In_1744);
and U13 (N_13,In_513,In_71);
nor U14 (N_14,In_1624,In_191);
nand U15 (N_15,In_153,In_1971);
nand U16 (N_16,In_1746,In_226);
xnor U17 (N_17,In_1692,In_377);
or U18 (N_18,In_146,In_1599);
nand U19 (N_19,In_983,In_135);
nand U20 (N_20,In_1285,In_187);
nand U21 (N_21,In_339,In_333);
and U22 (N_22,In_1793,In_735);
or U23 (N_23,In_899,In_1488);
or U24 (N_24,In_1379,In_1178);
nor U25 (N_25,In_843,In_755);
xnor U26 (N_26,In_764,In_1225);
nand U27 (N_27,In_1045,In_1575);
or U28 (N_28,In_1515,In_1986);
xnor U29 (N_29,In_656,In_232);
nor U30 (N_30,In_204,In_1069);
nand U31 (N_31,In_138,In_760);
nand U32 (N_32,In_1372,In_1328);
or U33 (N_33,In_475,In_711);
or U34 (N_34,In_1234,In_72);
or U35 (N_35,In_1299,In_456);
nand U36 (N_36,In_1381,In_9);
xnor U37 (N_37,In_1214,In_1851);
xnor U38 (N_38,In_391,In_1338);
and U39 (N_39,In_621,In_602);
xnor U40 (N_40,In_452,In_1665);
xnor U41 (N_41,In_1137,In_590);
nor U42 (N_42,In_1048,In_43);
and U43 (N_43,In_8,In_1713);
nand U44 (N_44,In_1640,In_1836);
or U45 (N_45,In_811,In_1422);
and U46 (N_46,In_1718,In_985);
nor U47 (N_47,In_346,In_3);
or U48 (N_48,In_402,In_797);
and U49 (N_49,In_235,In_1322);
xor U50 (N_50,In_1082,In_512);
nand U51 (N_51,In_1922,In_231);
nor U52 (N_52,In_1462,In_575);
nor U53 (N_53,In_595,In_464);
and U54 (N_54,In_682,In_1238);
or U55 (N_55,In_1546,In_348);
and U56 (N_56,In_1768,In_253);
nand U57 (N_57,In_1346,In_1789);
or U58 (N_58,In_522,In_931);
and U59 (N_59,In_940,In_211);
nor U60 (N_60,In_1762,In_1170);
xnor U61 (N_61,In_571,In_1895);
nand U62 (N_62,In_696,In_67);
or U63 (N_63,In_1129,In_203);
nand U64 (N_64,In_27,In_1426);
nand U65 (N_65,In_1516,In_1551);
nor U66 (N_66,In_1091,In_1146);
nand U67 (N_67,In_1866,In_417);
or U68 (N_68,In_795,In_802);
xnor U69 (N_69,In_295,In_1024);
nand U70 (N_70,In_1926,In_468);
nor U71 (N_71,In_1152,In_220);
and U72 (N_72,In_1994,In_936);
xor U73 (N_73,In_1587,In_761);
and U74 (N_74,In_1106,In_1061);
or U75 (N_75,In_1919,In_1331);
or U76 (N_76,In_465,In_1827);
nand U77 (N_77,In_774,In_932);
nor U78 (N_78,In_360,In_1850);
or U79 (N_79,In_1983,In_1219);
and U80 (N_80,In_1969,In_1620);
xor U81 (N_81,In_544,In_1077);
nand U82 (N_82,In_256,In_1728);
nand U83 (N_83,In_205,In_779);
and U84 (N_84,In_1279,In_788);
or U85 (N_85,In_1401,In_167);
or U86 (N_86,In_325,In_83);
nor U87 (N_87,In_658,In_183);
and U88 (N_88,In_1709,In_920);
and U89 (N_89,In_1953,In_819);
nand U90 (N_90,In_925,In_816);
nand U91 (N_91,In_474,In_103);
nor U92 (N_92,In_1016,In_1612);
nand U93 (N_93,In_414,In_42);
or U94 (N_94,In_335,In_1852);
nor U95 (N_95,In_94,In_1068);
nor U96 (N_96,In_1255,In_286);
nand U97 (N_97,In_494,In_28);
nor U98 (N_98,In_127,In_1253);
nand U99 (N_99,In_1326,In_292);
nand U100 (N_100,In_1585,In_1662);
or U101 (N_101,In_479,In_147);
or U102 (N_102,In_1882,In_1151);
or U103 (N_103,In_177,In_115);
nor U104 (N_104,In_1165,In_1311);
and U105 (N_105,In_408,In_1708);
and U106 (N_106,In_61,In_1180);
or U107 (N_107,In_1561,In_619);
nor U108 (N_108,In_1650,In_1795);
and U109 (N_109,In_1248,In_1360);
nor U110 (N_110,In_1192,In_1549);
and U111 (N_111,In_87,In_1678);
nand U112 (N_112,In_1093,In_1456);
or U113 (N_113,In_1593,In_1875);
nand U114 (N_114,In_1140,In_706);
nor U115 (N_115,In_1352,In_959);
nand U116 (N_116,In_726,In_1382);
and U117 (N_117,In_813,In_1797);
nand U118 (N_118,In_809,In_1130);
xnor U119 (N_119,In_1450,In_283);
nand U120 (N_120,In_1675,In_481);
nand U121 (N_121,In_1935,In_879);
and U122 (N_122,In_1230,In_587);
and U123 (N_123,In_355,In_987);
xor U124 (N_124,In_1108,In_1763);
xor U125 (N_125,In_1489,In_1453);
or U126 (N_126,In_1358,In_285);
nor U127 (N_127,In_551,In_1415);
and U128 (N_128,In_1378,In_1803);
and U129 (N_129,In_1752,In_1622);
and U130 (N_130,In_910,In_160);
and U131 (N_131,In_1288,In_25);
and U132 (N_132,In_1890,In_884);
nand U133 (N_133,In_1723,In_1569);
nor U134 (N_134,In_1128,In_1492);
nand U135 (N_135,In_466,In_1505);
nand U136 (N_136,In_158,In_1679);
or U137 (N_137,In_54,In_1740);
or U138 (N_138,In_1161,In_1993);
nor U139 (N_139,In_933,In_405);
or U140 (N_140,In_1033,In_316);
or U141 (N_141,In_1122,In_413);
or U142 (N_142,In_269,In_944);
nand U143 (N_143,In_865,In_1780);
xor U144 (N_144,In_1863,In_381);
and U145 (N_145,In_792,In_287);
nand U146 (N_146,In_574,In_1461);
nand U147 (N_147,In_1788,In_1065);
xnor U148 (N_148,In_275,In_659);
xor U149 (N_149,In_1658,In_796);
and U150 (N_150,In_576,In_569);
xor U151 (N_151,In_1908,In_582);
nand U152 (N_152,In_496,In_839);
and U153 (N_153,In_652,In_608);
xor U154 (N_154,In_1790,In_1974);
and U155 (N_155,In_1501,In_1308);
nor U156 (N_156,In_165,In_1846);
xor U157 (N_157,In_1179,In_1548);
or U158 (N_158,In_1717,In_1055);
nand U159 (N_159,In_1446,In_1083);
xor U160 (N_160,In_1252,In_965);
and U161 (N_161,In_1282,In_803);
xnor U162 (N_162,In_1547,In_154);
xnor U163 (N_163,In_584,In_937);
or U164 (N_164,In_151,In_1517);
nand U165 (N_165,In_1949,In_1941);
nor U166 (N_166,In_1268,In_332);
or U167 (N_167,In_470,In_596);
xor U168 (N_168,In_1104,In_1811);
nand U169 (N_169,In_666,In_1646);
nor U170 (N_170,In_1909,In_1275);
xnor U171 (N_171,In_445,In_1476);
nand U172 (N_172,In_871,In_1274);
xnor U173 (N_173,In_1062,In_106);
xor U174 (N_174,In_1873,In_1059);
and U175 (N_175,In_943,In_1364);
or U176 (N_176,In_1472,In_1534);
nand U177 (N_177,In_780,In_493);
and U178 (N_178,In_1817,In_1353);
and U179 (N_179,In_923,In_1403);
xor U180 (N_180,In_639,In_527);
and U181 (N_181,In_1816,In_859);
and U182 (N_182,In_174,In_505);
nand U183 (N_183,In_1094,In_208);
or U184 (N_184,In_901,In_998);
nand U185 (N_185,In_1757,In_16);
nor U186 (N_186,In_1791,In_46);
xor U187 (N_187,In_1075,In_314);
nand U188 (N_188,In_31,In_585);
and U189 (N_189,In_353,In_1030);
nor U190 (N_190,In_1749,In_1089);
nor U191 (N_191,In_1959,In_261);
xnor U192 (N_192,In_1627,In_876);
and U193 (N_193,In_1000,In_1519);
or U194 (N_194,In_1204,In_961);
and U195 (N_195,In_84,In_1747);
xor U196 (N_196,In_553,In_842);
or U197 (N_197,In_438,In_1638);
xnor U198 (N_198,In_1283,In_44);
nor U199 (N_199,In_129,In_689);
or U200 (N_200,In_1583,In_69);
nand U201 (N_201,In_834,In_672);
or U202 (N_202,In_17,In_1444);
xnor U203 (N_203,In_412,In_1900);
and U204 (N_204,In_111,In_1023);
nor U205 (N_205,In_1742,In_1018);
and U206 (N_206,In_238,In_701);
nor U207 (N_207,In_592,In_559);
nor U208 (N_208,In_1296,In_1921);
nand U209 (N_209,In_53,In_1772);
and U210 (N_210,In_1525,In_756);
and U211 (N_211,In_896,In_1554);
nand U212 (N_212,In_1384,In_827);
xnor U213 (N_213,In_958,In_180);
and U214 (N_214,In_173,In_258);
or U215 (N_215,In_1177,In_38);
nor U216 (N_216,In_302,In_971);
nand U217 (N_217,In_172,In_1854);
or U218 (N_218,In_1370,In_1464);
nand U219 (N_219,In_1293,In_249);
xor U220 (N_220,In_1373,In_573);
nand U221 (N_221,In_1079,In_826);
or U222 (N_222,In_323,In_1071);
or U223 (N_223,In_199,In_447);
or U224 (N_224,In_312,In_1318);
and U225 (N_225,In_380,In_949);
and U226 (N_226,In_1920,In_1758);
xor U227 (N_227,In_1292,In_246);
xor U228 (N_228,In_815,In_1819);
nor U229 (N_229,In_928,In_1934);
and U230 (N_230,In_1957,In_887);
or U231 (N_231,In_1374,In_1375);
and U232 (N_232,In_984,In_968);
nand U233 (N_233,In_1300,In_1483);
nor U234 (N_234,In_432,In_732);
nor U235 (N_235,In_555,In_924);
or U236 (N_236,In_123,In_1266);
nand U237 (N_237,In_311,In_885);
nor U238 (N_238,In_1820,In_860);
nand U239 (N_239,In_1429,In_955);
nor U240 (N_240,In_1998,In_718);
nor U241 (N_241,In_651,In_1944);
nand U242 (N_242,In_620,In_1681);
nor U243 (N_243,In_422,In_1112);
and U244 (N_244,In_653,In_953);
nand U245 (N_245,In_1743,In_421);
nor U246 (N_246,In_516,In_583);
nor U247 (N_247,In_678,In_579);
nor U248 (N_248,In_1427,In_416);
nor U249 (N_249,In_533,In_1298);
and U250 (N_250,In_1197,In_1171);
xor U251 (N_251,In_547,In_124);
nor U252 (N_252,In_1015,In_446);
nor U253 (N_253,In_790,In_59);
nor U254 (N_254,In_349,In_1903);
and U255 (N_255,In_1859,In_1669);
nand U256 (N_256,In_473,In_1878);
xor U257 (N_257,In_1247,In_1990);
and U258 (N_258,In_1495,In_0);
xor U259 (N_259,In_476,In_1007);
or U260 (N_260,In_1436,In_260);
nor U261 (N_261,In_1078,In_1195);
nor U262 (N_262,In_560,In_1223);
and U263 (N_263,In_1212,In_964);
nand U264 (N_264,In_1262,In_1226);
and U265 (N_265,In_1034,In_1887);
nor U266 (N_266,In_1163,In_1088);
xor U267 (N_267,In_1616,In_47);
nand U268 (N_268,In_1063,In_1932);
nand U269 (N_269,In_1750,In_601);
nand U270 (N_270,In_169,In_1691);
xor U271 (N_271,In_744,In_60);
nand U272 (N_272,In_273,In_155);
and U273 (N_273,In_749,In_686);
nor U274 (N_274,In_771,In_681);
or U275 (N_275,In_93,In_1821);
or U276 (N_276,In_477,In_981);
and U277 (N_277,In_159,In_540);
nand U278 (N_278,In_120,In_1241);
nand U279 (N_279,In_2,In_1265);
nor U280 (N_280,In_948,In_463);
nand U281 (N_281,In_1754,In_1564);
and U282 (N_282,In_1142,In_21);
nand U283 (N_283,In_808,In_277);
nand U284 (N_284,In_1786,In_1207);
or U285 (N_285,In_498,In_1798);
and U286 (N_286,In_1003,In_1860);
or U287 (N_287,In_1240,In_472);
nand U288 (N_288,In_733,In_1397);
or U289 (N_289,In_442,In_846);
nor U290 (N_290,In_1208,In_1837);
or U291 (N_291,In_233,In_556);
nand U292 (N_292,In_912,In_529);
nand U293 (N_293,In_1702,In_716);
or U294 (N_294,In_404,In_1448);
and U295 (N_295,In_700,In_611);
nand U296 (N_296,In_57,In_327);
or U297 (N_297,In_1443,In_561);
and U298 (N_298,In_274,In_1064);
or U299 (N_299,In_1916,In_55);
or U300 (N_300,In_471,In_1139);
nor U301 (N_301,In_960,In_80);
nand U302 (N_302,In_1654,In_1251);
xor U303 (N_303,In_684,In_1630);
and U304 (N_304,In_952,In_444);
nand U305 (N_305,In_1565,In_1703);
or U306 (N_306,In_101,In_1726);
and U307 (N_307,In_1209,In_1343);
or U308 (N_308,In_1591,In_216);
and U309 (N_309,In_791,In_210);
nor U310 (N_310,In_1838,In_436);
or U311 (N_311,In_102,In_1345);
or U312 (N_312,In_1341,In_1416);
and U313 (N_313,In_1822,In_1216);
xor U314 (N_314,In_1008,In_492);
nand U315 (N_315,In_1473,In_137);
and U316 (N_316,In_1655,In_1438);
nand U317 (N_317,In_1670,In_117);
nor U318 (N_318,In_1315,In_19);
nand U319 (N_319,In_637,In_1608);
nand U320 (N_320,In_298,In_886);
nand U321 (N_321,In_874,In_130);
nor U322 (N_322,In_1787,In_1309);
nand U323 (N_323,In_1276,In_484);
or U324 (N_324,In_114,In_534);
and U325 (N_325,In_1533,In_623);
nand U326 (N_326,In_1522,In_890);
xor U327 (N_327,In_1399,In_1155);
xnor U328 (N_328,In_1267,In_1110);
or U329 (N_329,In_1169,In_36);
or U330 (N_330,In_1294,In_1904);
nor U331 (N_331,In_1391,In_1220);
or U332 (N_332,In_324,In_1644);
and U333 (N_333,In_1150,In_1651);
or U334 (N_334,In_1537,In_1503);
nand U335 (N_335,In_543,In_291);
nor U336 (N_336,In_134,In_1536);
nand U337 (N_337,In_1556,In_708);
nor U338 (N_338,In_1945,In_900);
and U339 (N_339,In_23,In_632);
xor U340 (N_340,In_1694,In_1383);
or U341 (N_341,In_748,In_1245);
nand U342 (N_342,In_1290,In_223);
or U343 (N_343,In_91,In_1720);
xnor U344 (N_344,In_1733,In_1645);
and U345 (N_345,In_1567,In_108);
and U346 (N_346,In_352,In_1305);
and U347 (N_347,In_593,In_613);
or U348 (N_348,In_1159,In_250);
nand U349 (N_349,In_1674,In_1526);
and U350 (N_350,In_357,In_1596);
nand U351 (N_351,In_804,In_143);
or U352 (N_352,In_81,In_1404);
and U353 (N_353,In_946,In_300);
and U354 (N_354,In_1938,In_1231);
or U355 (N_355,In_239,In_186);
nand U356 (N_356,In_424,In_1289);
nor U357 (N_357,In_703,In_96);
xnor U358 (N_358,In_838,In_1357);
xnor U359 (N_359,In_1261,In_941);
or U360 (N_360,In_104,In_752);
nor U361 (N_361,In_1423,In_1160);
or U362 (N_362,In_1518,In_977);
nor U363 (N_363,In_1125,In_1497);
and U364 (N_364,In_1010,In_1101);
nand U365 (N_365,In_1542,In_1400);
xor U366 (N_366,In_1676,In_1474);
and U367 (N_367,In_1452,In_926);
and U368 (N_368,In_1,In_1175);
and U369 (N_369,In_996,In_618);
and U370 (N_370,In_999,In_1395);
xnor U371 (N_371,In_1109,In_1297);
and U372 (N_372,In_1661,In_832);
xor U373 (N_373,In_854,In_290);
and U374 (N_374,In_1936,In_1040);
nor U375 (N_375,In_1043,In_100);
nand U376 (N_376,In_599,In_1482);
xor U377 (N_377,In_1025,In_64);
nor U378 (N_378,In_66,In_1144);
nand U379 (N_379,In_457,In_673);
or U380 (N_380,In_1221,In_1393);
or U381 (N_381,In_1893,In_904);
nor U382 (N_382,In_604,In_616);
nor U383 (N_383,In_1842,In_1340);
xor U384 (N_384,In_1258,In_409);
xnor U385 (N_385,In_164,In_1877);
xor U386 (N_386,In_32,In_1099);
and U387 (N_387,In_453,In_1347);
or U388 (N_388,In_1454,In_162);
xnor U389 (N_389,In_175,In_1136);
or U390 (N_390,In_1832,In_95);
nor U391 (N_391,In_1652,In_383);
nor U392 (N_392,In_699,In_730);
or U393 (N_393,In_594,In_1408);
nor U394 (N_394,In_6,In_259);
xor U395 (N_395,In_480,In_1779);
and U396 (N_396,In_709,In_746);
xor U397 (N_397,In_459,In_1633);
or U398 (N_398,In_688,In_423);
nor U399 (N_399,In_939,In_310);
nand U400 (N_400,In_79,In_1313);
nor U401 (N_401,In_818,In_554);
nor U402 (N_402,In_693,In_638);
or U403 (N_403,In_384,In_1269);
nor U404 (N_404,In_1637,In_5);
xnor U405 (N_405,In_1133,In_1685);
or U406 (N_406,In_369,In_801);
xnor U407 (N_407,In_301,In_857);
or U408 (N_408,In_970,In_1712);
nand U409 (N_409,In_1500,In_988);
nand U410 (N_410,In_705,In_1853);
or U411 (N_411,In_878,In_1046);
nor U412 (N_412,In_430,In_1405);
nand U413 (N_413,In_491,In_642);
nor U414 (N_414,In_1614,In_640);
and U415 (N_415,In_1491,In_1814);
nand U416 (N_416,In_1359,In_1433);
xor U417 (N_417,In_782,In_829);
and U418 (N_418,In_668,In_1553);
and U419 (N_419,In_1734,In_541);
and U420 (N_420,In_1958,In_1156);
and U421 (N_421,In_850,In_128);
nor U422 (N_422,In_338,In_548);
nor U423 (N_423,In_263,In_580);
or U424 (N_424,In_598,In_1930);
and U425 (N_425,In_1508,In_1312);
or U426 (N_426,In_257,In_1287);
nand U427 (N_427,In_467,In_462);
and U428 (N_428,In_136,In_1985);
nand U429 (N_429,In_893,In_1244);
nand U430 (N_430,In_724,In_1199);
xnor U431 (N_431,In_228,In_858);
and U432 (N_432,In_1799,In_1153);
and U433 (N_433,In_1070,In_282);
nor U434 (N_434,In_1232,In_1074);
nand U435 (N_435,In_1684,In_429);
nand U436 (N_436,In_1172,In_506);
nand U437 (N_437,In_644,In_1050);
nor U438 (N_438,In_76,In_1615);
or U439 (N_439,In_773,In_1092);
and U440 (N_440,In_515,In_1806);
xor U441 (N_441,In_1126,In_497);
and U442 (N_442,In_1700,In_992);
xnor U443 (N_443,In_1410,In_1613);
nor U444 (N_444,In_1200,In_51);
nor U445 (N_445,In_190,In_655);
nor U446 (N_446,In_168,In_1598);
xnor U447 (N_447,In_329,In_1164);
and U448 (N_448,In_1215,In_1603);
nand U449 (N_449,In_715,In_617);
nand U450 (N_450,In_1970,In_1978);
xor U451 (N_451,In_519,In_552);
nand U452 (N_452,In_1925,In_806);
nor U453 (N_453,In_1434,In_1227);
xnor U454 (N_454,In_1871,In_189);
and U455 (N_455,In_1579,In_646);
xor U456 (N_456,In_206,In_880);
xnor U457 (N_457,In_1738,In_1987);
nand U458 (N_458,In_1166,In_306);
nand U459 (N_459,In_1504,In_1705);
nand U460 (N_460,In_119,In_989);
and U461 (N_461,In_1531,In_279);
and U462 (N_462,In_193,In_605);
or U463 (N_463,In_271,In_1918);
nand U464 (N_464,In_823,In_1988);
or U465 (N_465,In_694,In_1629);
nand U466 (N_466,In_1335,In_1385);
or U467 (N_467,In_488,In_1727);
xnor U468 (N_468,In_1864,In_1514);
nor U469 (N_469,In_1590,In_1176);
nor U470 (N_470,In_1597,In_1604);
and U471 (N_471,In_37,In_793);
or U472 (N_472,In_1337,In_1568);
and U473 (N_473,In_1745,In_1571);
or U474 (N_474,In_411,In_909);
or U475 (N_475,In_240,In_237);
nand U476 (N_476,In_660,In_1507);
nor U477 (N_477,In_934,In_905);
or U478 (N_478,In_1584,In_1607);
and U479 (N_479,In_1719,In_550);
nand U480 (N_480,In_683,In_455);
or U481 (N_481,In_898,In_1001);
or U482 (N_482,In_1035,In_1872);
and U483 (N_483,In_99,In_1967);
xnor U484 (N_484,In_1813,In_528);
nor U485 (N_485,In_62,In_13);
nand U486 (N_486,In_535,In_1147);
xnor U487 (N_487,In_787,In_1609);
nand U488 (N_488,In_525,In_156);
nand U489 (N_489,In_577,In_647);
xnor U490 (N_490,In_754,In_1186);
xor U491 (N_491,In_1329,In_524);
or U492 (N_492,In_636,In_1148);
nor U493 (N_493,In_370,In_490);
or U494 (N_494,In_918,In_1032);
or U495 (N_495,In_1162,In_624);
or U496 (N_496,In_1342,In_313);
nor U497 (N_497,In_49,In_1884);
xnor U498 (N_498,In_1004,In_1102);
and U499 (N_499,In_1901,In_1915);
or U500 (N_500,In_1688,In_1021);
nor U501 (N_501,In_326,In_671);
and U502 (N_502,In_1770,In_821);
and U503 (N_503,In_1664,In_1229);
and U504 (N_504,In_566,In_869);
and U505 (N_505,In_1013,In_1354);
and U506 (N_506,In_1849,In_112);
or U507 (N_507,In_1984,In_1527);
and U508 (N_508,In_320,In_1611);
or U509 (N_509,In_1979,In_1595);
nand U510 (N_510,In_1281,In_1509);
xnor U511 (N_511,In_916,In_1862);
or U512 (N_512,In_304,In_628);
nor U513 (N_513,In_1103,In_1237);
nor U514 (N_514,In_1550,In_163);
and U515 (N_515,In_1559,In_35);
nor U516 (N_516,In_1931,In_1725);
xnor U517 (N_517,In_741,In_1044);
nor U518 (N_518,In_670,In_407);
and U519 (N_519,In_627,In_1320);
xor U520 (N_520,In_431,In_510);
or U521 (N_521,In_737,In_1291);
nor U522 (N_522,In_1181,In_1933);
or U523 (N_523,In_1100,In_1280);
nor U524 (N_524,In_1540,In_1927);
nor U525 (N_525,In_537,In_1996);
and U526 (N_526,In_1115,In_345);
nor U527 (N_527,In_954,In_676);
nor U528 (N_528,In_366,In_1699);
and U529 (N_529,In_1809,In_1572);
nand U530 (N_530,In_875,In_1766);
and U531 (N_531,In_1330,In_1490);
nand U532 (N_532,In_690,In_1022);
and U533 (N_533,In_68,In_1881);
or U534 (N_534,In_1457,In_1698);
xnor U535 (N_535,In_1060,In_990);
or U536 (N_536,In_1689,In_1277);
or U537 (N_537,In_74,In_1783);
or U538 (N_538,In_1191,In_906);
nor U539 (N_539,In_1390,In_1955);
and U540 (N_540,In_1116,In_105);
or U541 (N_541,In_1991,In_1049);
and U542 (N_542,In_1167,In_1419);
xnor U543 (N_543,In_1924,In_1885);
xnor U544 (N_544,In_685,In_1861);
or U545 (N_545,In_350,In_1962);
xnor U546 (N_546,In_212,In_382);
and U547 (N_547,In_663,In_243);
nor U548 (N_548,In_1697,In_245);
nand U549 (N_549,In_770,In_1217);
and U550 (N_550,In_213,In_845);
nor U551 (N_551,In_1543,In_1566);
or U552 (N_552,In_680,In_1336);
xnor U553 (N_553,In_1802,In_1532);
or U554 (N_554,In_1467,In_511);
nor U555 (N_555,In_1671,In_951);
and U556 (N_556,In_1442,In_1722);
nor U557 (N_557,In_1605,In_1301);
xnor U558 (N_558,In_1833,In_1947);
and U559 (N_559,In_1939,In_530);
nor U560 (N_560,In_1141,In_1867);
xnor U561 (N_561,In_1222,In_1012);
nor U562 (N_562,In_772,In_1892);
xor U563 (N_563,In_836,In_361);
or U564 (N_564,In_662,In_1203);
nand U565 (N_565,In_364,In_1090);
nand U566 (N_566,In_41,In_1963);
nand U567 (N_567,In_139,In_1677);
and U568 (N_568,In_1306,In_1610);
nor U569 (N_569,In_868,In_478);
nand U570 (N_570,In_778,In_626);
nor U571 (N_571,In_938,In_789);
or U572 (N_572,In_588,In_1544);
or U573 (N_573,In_200,In_739);
and U574 (N_574,In_1663,In_945);
nand U575 (N_575,In_398,In_166);
nor U576 (N_576,In_1190,In_641);
nand U577 (N_577,In_215,In_86);
nor U578 (N_578,In_1641,In_1765);
nor U579 (N_579,In_1848,In_1425);
nand U580 (N_580,In_1493,In_435);
or U581 (N_581,In_1316,In_386);
nand U582 (N_582,In_1812,In_1889);
nor U583 (N_583,In_643,In_1521);
nor U584 (N_584,In_1005,In_1858);
and U585 (N_585,In_131,In_1350);
nand U586 (N_586,In_374,In_33);
nor U587 (N_587,In_434,In_109);
and U588 (N_588,In_4,In_1981);
xnor U589 (N_589,In_1801,In_1756);
and U590 (N_590,In_39,In_634);
nand U591 (N_591,In_1825,In_1577);
or U592 (N_592,In_317,In_161);
nand U593 (N_593,In_1977,In_674);
or U594 (N_594,In_1246,In_942);
or U595 (N_595,In_675,In_753);
and U596 (N_596,In_1038,In_888);
and U597 (N_597,In_1946,In_1829);
xnor U598 (N_598,In_373,In_1445);
nand U599 (N_599,In_786,In_1185);
nor U600 (N_600,In_1520,In_976);
or U601 (N_601,In_1530,In_242);
nor U602 (N_602,In_974,In_557);
nand U603 (N_603,In_1942,In_1430);
xnor U604 (N_604,In_667,In_956);
xnor U605 (N_605,In_1656,In_1834);
nand U606 (N_606,In_336,In_307);
nand U607 (N_607,In_777,In_1760);
xnor U608 (N_608,In_1898,In_219);
or U609 (N_609,In_1307,In_305);
nor U610 (N_610,In_1249,In_1396);
or U611 (N_611,In_610,In_1417);
or U612 (N_612,In_820,In_1117);
and U613 (N_613,In_514,In_725);
nor U614 (N_614,In_657,In_1562);
and U615 (N_615,In_1810,In_448);
and U616 (N_616,In_1907,In_197);
xor U617 (N_617,In_88,In_633);
xor U618 (N_618,In_665,In_319);
and U619 (N_619,In_1107,In_1524);
xor U620 (N_620,In_1158,In_1498);
nand U621 (N_621,In_1905,In_1928);
nor U622 (N_622,In_1239,In_1051);
or U623 (N_623,In_840,In_736);
xnor U624 (N_624,In_600,In_687);
and U625 (N_625,In_1824,In_520);
nor U626 (N_626,In_218,In_692);
or U627 (N_627,In_1484,In_1475);
or U628 (N_628,In_1707,In_52);
and U629 (N_629,In_1420,In_280);
nand U630 (N_630,In_1377,In_581);
xnor U631 (N_631,In_1339,In_654);
or U632 (N_632,In_1672,In_1736);
and U633 (N_633,In_758,In_288);
nor U634 (N_634,In_1923,In_831);
nand U635 (N_635,In_281,In_1844);
nor U636 (N_636,In_1891,In_1714);
or U637 (N_637,In_1830,In_769);
xor U638 (N_638,In_1334,In_1224);
nand U639 (N_639,In_248,In_399);
nor U640 (N_640,In_195,In_1696);
and U641 (N_641,In_376,In_1729);
and U642 (N_642,In_727,In_864);
nand U643 (N_643,In_1632,In_482);
xor U644 (N_644,In_1960,In_720);
xnor U645 (N_645,In_1659,In_1113);
and U646 (N_646,In_1487,In_1643);
xnor U647 (N_647,In_1841,In_719);
nor U648 (N_648,In_1260,In_1459);
nor U649 (N_649,In_1600,In_1631);
xor U650 (N_650,In_1259,In_1471);
nand U651 (N_651,In_980,In_415);
nor U652 (N_652,In_1096,In_378);
nand U653 (N_653,In_1014,In_837);
and U654 (N_654,In_1796,In_244);
and U655 (N_655,In_400,In_118);
nor U656 (N_656,In_1201,In_927);
or U657 (N_657,In_1606,In_1870);
and U658 (N_658,In_1460,In_255);
nor U659 (N_659,In_814,In_1418);
and U660 (N_660,In_503,In_697);
nand U661 (N_661,In_145,In_1243);
or U662 (N_662,In_517,In_828);
or U663 (N_663,In_201,In_1193);
nor U664 (N_664,In_1794,In_1362);
xor U665 (N_665,In_63,In_612);
and U666 (N_666,In_1463,In_1072);
nand U667 (N_667,In_406,In_460);
nor U668 (N_668,In_1499,In_783);
nand U669 (N_669,In_1999,In_297);
nor U670 (N_670,In_184,In_499);
nor U671 (N_671,In_1325,In_1594);
nand U672 (N_672,In_1095,In_141);
nor U673 (N_673,In_48,In_1589);
nand U674 (N_674,In_568,In_897);
xnor U675 (N_675,In_1545,In_629);
or U676 (N_676,In_523,In_1168);
and U677 (N_677,In_747,In_1210);
xnor U678 (N_678,In_1800,In_1529);
and U679 (N_679,In_1759,In_1687);
or U680 (N_680,In_1512,In_1017);
nand U681 (N_681,In_1961,In_379);
nor U682 (N_682,In_1120,In_536);
nor U683 (N_683,In_1213,In_1052);
nor U684 (N_684,In_1271,In_892);
nor U685 (N_685,In_365,In_861);
nand U686 (N_686,In_1952,In_794);
and U687 (N_687,In_731,In_181);
nand U688 (N_688,In_1826,In_188);
and U689 (N_689,In_545,In_606);
xor U690 (N_690,In_1804,In_1428);
nor U691 (N_691,In_734,In_1363);
xnor U692 (N_692,In_1781,In_441);
nand U693 (N_693,In_1421,In_1538);
and U694 (N_694,In_1218,In_759);
nor U695 (N_695,In_351,In_501);
nand U696 (N_696,In_714,In_1782);
and U697 (N_697,In_371,In_1706);
or U698 (N_698,In_776,In_1211);
nand U699 (N_699,In_284,In_1173);
or U700 (N_700,In_1975,In_1154);
and U701 (N_701,In_1348,In_1560);
or U702 (N_702,In_526,In_170);
nor U703 (N_703,In_603,In_1535);
nand U704 (N_704,In_895,In_337);
nor U705 (N_705,In_798,In_867);
xnor U706 (N_706,In_1097,In_1174);
nand U707 (N_707,In_691,In_1323);
nor U708 (N_708,In_1807,In_1386);
nand U709 (N_709,In_328,In_194);
or U710 (N_710,In_65,In_1388);
or U711 (N_711,In_1286,In_648);
and U712 (N_712,In_1412,In_1695);
xor U713 (N_713,In_1496,In_1368);
and U714 (N_714,In_1948,In_1732);
xor U715 (N_715,In_1680,In_863);
xor U716 (N_716,In_847,In_133);
nand U717 (N_717,In_34,In_1389);
xnor U718 (N_718,In_558,In_372);
nand U719 (N_719,In_241,In_1494);
and U720 (N_720,In_150,In_922);
and U721 (N_721,In_1808,In_810);
or U722 (N_722,In_917,In_707);
or U723 (N_723,In_1704,In_293);
and U724 (N_724,In_1902,In_1578);
xor U725 (N_725,In_1361,In_375);
nand U726 (N_726,In_1576,In_171);
xnor U727 (N_727,In_1897,In_1968);
nor U728 (N_728,In_1701,In_1673);
or U729 (N_729,In_1073,In_833);
xor U730 (N_730,In_403,In_722);
nand U731 (N_731,In_132,In_1776);
nor U732 (N_732,In_1666,In_995);
xnor U733 (N_733,In_1124,In_542);
xnor U734 (N_734,In_1715,In_401);
nor U735 (N_735,In_1914,In_830);
nand U736 (N_736,In_704,In_1828);
xor U737 (N_737,In_1965,In_883);
and U738 (N_738,In_1573,In_433);
xnor U739 (N_739,In_1138,In_1202);
and U740 (N_740,In_1009,In_1721);
nand U741 (N_741,In_1036,In_784);
and U742 (N_742,In_1039,In_1601);
xnor U743 (N_743,In_1710,In_589);
or U744 (N_744,In_1189,In_1769);
xnor U745 (N_745,In_504,In_877);
xor U746 (N_746,In_1228,In_907);
nor U747 (N_747,In_267,In_207);
or U748 (N_748,In_679,In_1502);
nor U749 (N_749,In_1478,In_539);
nand U750 (N_750,In_1029,In_1626);
or U751 (N_751,In_1123,In_1635);
and U752 (N_752,In_1753,In_278);
and U753 (N_753,In_1319,In_388);
or U754 (N_754,In_538,In_1087);
nand U755 (N_755,In_967,In_1660);
or U756 (N_756,In_852,In_570);
and U757 (N_757,In_1523,In_1653);
nor U758 (N_758,In_224,In_1856);
nor U759 (N_759,In_1563,In_1634);
nand U760 (N_760,In_389,In_717);
nor U761 (N_761,In_1899,In_1042);
xnor U762 (N_762,In_70,In_1131);
nand U763 (N_763,In_763,In_1541);
nor U764 (N_764,In_113,In_966);
xnor U765 (N_765,In_1406,In_1026);
nand U766 (N_766,In_1080,In_410);
nor U767 (N_767,In_508,In_1648);
xor U768 (N_768,In_807,In_1731);
xor U769 (N_769,In_800,In_40);
or U770 (N_770,In_178,In_740);
or U771 (N_771,In_1182,In_609);
and U772 (N_772,In_712,In_1937);
and U773 (N_773,In_1387,In_1440);
nand U774 (N_774,In_1735,In_341);
nand U775 (N_775,In_518,In_1888);
xnor U776 (N_776,In_394,In_1011);
and U777 (N_777,In_1823,In_973);
and U778 (N_778,In_835,In_450);
or U779 (N_779,In_1847,In_919);
and U780 (N_780,In_1256,In_742);
and U781 (N_781,In_1076,In_1031);
and U782 (N_782,In_1906,In_855);
or U783 (N_783,In_483,In_1205);
or U784 (N_784,In_1435,In_994);
xor U785 (N_785,In_1552,In_1966);
xnor U786 (N_786,In_1815,In_1690);
and U787 (N_787,In_567,In_911);
nand U788 (N_788,In_1455,In_532);
xor U789 (N_789,In_1465,In_849);
or U790 (N_790,In_1951,In_1424);
xnor U791 (N_791,In_698,In_451);
xor U792 (N_792,In_1964,In_270);
or U793 (N_793,In_1628,In_330);
and U794 (N_794,In_1845,In_661);
or U795 (N_795,In_50,In_1657);
nand U796 (N_796,In_1510,In_254);
nand U797 (N_797,In_1686,In_225);
nor U798 (N_798,In_597,In_1912);
nand U799 (N_799,In_318,In_1580);
nor U800 (N_800,In_77,In_1145);
and U801 (N_801,In_751,In_29);
nor U802 (N_802,In_321,In_1047);
xnor U803 (N_803,In_1511,In_1865);
nor U804 (N_804,In_1623,In_738);
and U805 (N_805,In_1321,In_1081);
nand U806 (N_806,In_461,In_247);
or U807 (N_807,In_1777,In_85);
nor U808 (N_808,In_1874,In_1263);
or U809 (N_809,In_1084,In_824);
nand U810 (N_810,In_289,In_1184);
or U811 (N_811,In_1458,In_1855);
or U812 (N_812,In_507,In_1149);
nand U813 (N_813,In_1716,In_1402);
nand U814 (N_814,In_1206,In_363);
nor U815 (N_815,In_586,In_1785);
nor U816 (N_816,In_268,In_1913);
xnor U817 (N_817,In_309,In_1792);
xor U818 (N_818,In_294,In_625);
nor U819 (N_819,In_426,In_882);
xnor U820 (N_820,In_1840,In_1198);
or U821 (N_821,In_1910,In_664);
nor U822 (N_822,In_1592,In_1755);
nor U823 (N_823,In_30,In_1413);
and U824 (N_824,In_222,In_1943);
nand U825 (N_825,In_1896,In_142);
nand U826 (N_826,In_152,In_45);
and U827 (N_827,In_947,In_591);
and U828 (N_828,In_20,In_1355);
nand U829 (N_829,In_914,In_872);
or U830 (N_830,In_157,In_1917);
nand U831 (N_831,In_1767,In_993);
and U832 (N_832,In_368,In_1006);
nor U833 (N_833,In_702,In_58);
xnor U834 (N_834,In_1414,In_344);
or U835 (N_835,In_1639,In_1588);
nand U836 (N_836,In_930,In_767);
nand U837 (N_837,In_1118,In_1911);
or U838 (N_838,In_757,In_359);
xnor U839 (N_839,In_1477,In_486);
nor U840 (N_840,In_1773,In_1751);
and U841 (N_841,In_710,In_489);
nor U842 (N_842,In_851,In_340);
nor U843 (N_843,In_1570,In_1295);
xnor U844 (N_844,In_1365,In_1127);
nor U845 (N_845,In_458,In_1950);
and U846 (N_846,In_439,In_308);
or U847 (N_847,In_862,In_1683);
and U848 (N_848,In_848,In_1157);
nor U849 (N_849,In_428,In_649);
nor U850 (N_850,In_1085,In_1880);
nand U851 (N_851,In_500,In_397);
and U852 (N_852,In_179,In_1349);
and U853 (N_853,In_1183,In_669);
xor U854 (N_854,In_1392,In_509);
or U855 (N_855,In_1778,In_870);
or U856 (N_856,In_1513,In_229);
xor U857 (N_857,In_419,In_768);
or U858 (N_858,In_92,In_978);
xor U859 (N_859,In_564,In_750);
nand U860 (N_860,In_1278,In_1121);
and U861 (N_861,In_1086,In_10);
and U862 (N_862,In_844,In_82);
nor U863 (N_863,In_622,In_1973);
nand U864 (N_864,In_1027,In_1839);
and U865 (N_865,In_1879,In_495);
xnor U866 (N_866,In_1647,In_252);
and U867 (N_867,In_1114,In_192);
xor U868 (N_868,In_805,In_979);
nand U869 (N_869,In_1621,In_125);
or U870 (N_870,In_392,In_1098);
or U871 (N_871,In_73,In_1324);
nand U872 (N_872,In_1284,In_915);
or U873 (N_873,In_485,In_799);
nor U874 (N_874,In_531,In_1451);
nand U875 (N_875,In_1054,In_975);
nand U876 (N_876,In_230,In_1642);
or U877 (N_877,In_1105,In_1481);
nand U878 (N_878,In_1188,In_1649);
or U879 (N_879,In_1250,In_14);
xor U880 (N_880,In_1868,In_1470);
nand U881 (N_881,In_98,In_913);
and U882 (N_882,In_565,In_1761);
and U883 (N_883,In_1619,In_149);
and U884 (N_884,In_1775,In_122);
or U885 (N_885,In_356,In_1310);
nand U886 (N_886,In_615,In_1257);
nand U887 (N_887,In_1028,In_1954);
nand U888 (N_888,In_635,In_24);
and U889 (N_889,In_1976,In_343);
xor U890 (N_890,In_198,In_1366);
or U891 (N_891,In_90,In_866);
and U892 (N_892,In_1236,In_1667);
xor U893 (N_893,In_743,In_469);
nor U894 (N_894,In_1869,In_1376);
xor U895 (N_895,In_18,In_75);
nor U896 (N_896,In_713,In_1929);
nor U897 (N_897,In_695,In_22);
xor U898 (N_898,In_1407,In_645);
xor U899 (N_899,In_578,In_56);
nor U900 (N_900,In_1254,In_1327);
and U901 (N_901,In_1196,In_873);
xor U902 (N_902,In_331,In_1711);
and U903 (N_903,In_1739,In_1989);
nand U904 (N_904,In_1411,In_299);
nor U905 (N_905,In_1469,In_266);
nand U906 (N_906,In_1771,In_1135);
nand U907 (N_907,In_1302,In_549);
nor U908 (N_908,In_296,In_121);
nor U909 (N_909,In_817,In_1317);
nand U910 (N_910,In_929,In_202);
and U911 (N_911,In_196,In_563);
nor U912 (N_912,In_454,In_15);
nand U913 (N_913,In_962,In_1020);
or U914 (N_914,In_342,In_853);
and U915 (N_915,In_390,In_234);
nand U916 (N_916,In_986,In_841);
and U917 (N_917,In_972,In_322);
nand U918 (N_918,In_1774,In_1982);
and U919 (N_919,In_963,In_1618);
and U920 (N_920,In_902,In_107);
nand U921 (N_921,In_1480,In_1617);
and U922 (N_922,In_1805,In_1486);
xnor U923 (N_923,In_1439,In_1682);
and U924 (N_924,In_856,In_607);
or U925 (N_925,In_1539,In_1367);
or U926 (N_926,In_1272,In_358);
nand U927 (N_927,In_1233,In_991);
nor U928 (N_928,In_969,In_894);
xor U929 (N_929,In_982,In_276);
and U930 (N_930,In_1972,In_236);
or U931 (N_931,In_1058,In_1980);
or U932 (N_932,In_889,In_1041);
xnor U933 (N_933,In_1724,In_1737);
nand U934 (N_934,In_521,In_78);
nand U935 (N_935,In_1693,In_723);
nand U936 (N_936,In_1356,In_209);
or U937 (N_937,In_26,In_1764);
and U938 (N_938,In_1894,In_1784);
or U939 (N_939,In_126,In_1371);
nand U940 (N_940,In_1264,In_614);
nand U941 (N_941,In_1134,In_1194);
nor U942 (N_942,In_1835,In_144);
xnor U943 (N_943,In_251,In_1409);
and U944 (N_944,In_11,In_393);
nor U945 (N_945,In_1940,In_1581);
xor U946 (N_946,In_997,In_650);
or U947 (N_947,In_449,In_1956);
and U948 (N_948,In_950,In_334);
and U949 (N_949,In_1057,In_437);
and U950 (N_950,In_418,In_1019);
nand U951 (N_951,In_677,In_785);
xnor U952 (N_952,In_546,In_110);
nor U953 (N_953,In_89,In_1479);
nand U954 (N_954,In_1187,In_140);
and U955 (N_955,In_1586,In_395);
nand U956 (N_956,In_487,In_362);
and U957 (N_957,In_1528,In_148);
and U958 (N_958,In_272,In_1273);
xnor U959 (N_959,In_572,In_265);
nor U960 (N_960,In_425,In_1111);
and U961 (N_961,In_396,In_1831);
xor U962 (N_962,In_1235,In_1369);
nand U963 (N_963,In_1242,In_957);
and U964 (N_964,In_1332,In_1485);
nand U965 (N_965,In_227,In_1132);
and U966 (N_966,In_387,In_217);
or U967 (N_967,In_1602,In_1995);
nor U968 (N_968,In_728,In_354);
or U969 (N_969,In_116,In_1557);
and U970 (N_970,In_1625,In_1876);
or U971 (N_971,In_1056,In_1304);
xnor U972 (N_972,In_385,In_264);
or U973 (N_973,In_185,In_1067);
and U974 (N_974,In_1447,In_1857);
xnor U975 (N_975,In_97,In_1333);
or U976 (N_976,In_822,In_630);
and U977 (N_977,In_745,In_729);
xor U978 (N_978,In_1748,In_765);
or U979 (N_979,In_908,In_1555);
nor U980 (N_980,In_440,In_762);
and U981 (N_981,In_443,In_1398);
nand U982 (N_982,In_1574,In_781);
and U983 (N_983,In_721,In_1668);
or U984 (N_984,In_12,In_1843);
nor U985 (N_985,In_1432,In_420);
xnor U986 (N_986,In_1558,In_881);
nand U987 (N_987,In_1449,In_812);
nand U988 (N_988,In_1506,In_315);
xor U989 (N_989,In_1886,In_1119);
or U990 (N_990,In_347,In_1818);
or U991 (N_991,In_1351,In_262);
and U992 (N_992,In_1053,In_1437);
nor U993 (N_993,In_1303,In_214);
or U994 (N_994,In_1636,In_1314);
or U995 (N_995,In_1002,In_1344);
nor U996 (N_996,In_1066,In_1380);
nand U997 (N_997,In_903,In_303);
nor U998 (N_998,In_182,In_1883);
xor U999 (N_999,In_935,In_1466);
nor U1000 (N_1000,In_1586,In_660);
nor U1001 (N_1001,In_526,In_1647);
and U1002 (N_1002,In_1070,In_678);
and U1003 (N_1003,In_1,In_716);
nand U1004 (N_1004,In_1653,In_962);
or U1005 (N_1005,In_145,In_1868);
nand U1006 (N_1006,In_734,In_799);
xor U1007 (N_1007,In_1455,In_1809);
and U1008 (N_1008,In_1282,In_235);
and U1009 (N_1009,In_1628,In_1791);
nor U1010 (N_1010,In_1861,In_261);
xnor U1011 (N_1011,In_126,In_169);
or U1012 (N_1012,In_85,In_342);
or U1013 (N_1013,In_56,In_1918);
xnor U1014 (N_1014,In_912,In_1650);
nor U1015 (N_1015,In_1947,In_1175);
xnor U1016 (N_1016,In_728,In_1203);
or U1017 (N_1017,In_1131,In_606);
or U1018 (N_1018,In_48,In_1397);
nand U1019 (N_1019,In_1120,In_1820);
or U1020 (N_1020,In_1825,In_44);
xor U1021 (N_1021,In_1091,In_1099);
nor U1022 (N_1022,In_246,In_1805);
nor U1023 (N_1023,In_41,In_1402);
xnor U1024 (N_1024,In_1555,In_1730);
and U1025 (N_1025,In_112,In_627);
or U1026 (N_1026,In_744,In_192);
or U1027 (N_1027,In_1780,In_378);
xnor U1028 (N_1028,In_1267,In_170);
xnor U1029 (N_1029,In_1970,In_869);
nand U1030 (N_1030,In_1658,In_380);
and U1031 (N_1031,In_1880,In_1969);
xnor U1032 (N_1032,In_453,In_555);
or U1033 (N_1033,In_643,In_286);
nand U1034 (N_1034,In_348,In_817);
nor U1035 (N_1035,In_623,In_360);
nand U1036 (N_1036,In_443,In_792);
or U1037 (N_1037,In_1946,In_1469);
and U1038 (N_1038,In_1993,In_297);
and U1039 (N_1039,In_118,In_1233);
nand U1040 (N_1040,In_482,In_1833);
or U1041 (N_1041,In_775,In_1914);
nor U1042 (N_1042,In_1492,In_213);
nand U1043 (N_1043,In_175,In_1646);
nor U1044 (N_1044,In_166,In_439);
and U1045 (N_1045,In_1574,In_150);
xor U1046 (N_1046,In_473,In_1651);
xor U1047 (N_1047,In_420,In_220);
nand U1048 (N_1048,In_1831,In_1729);
or U1049 (N_1049,In_1486,In_622);
xnor U1050 (N_1050,In_1936,In_1971);
nor U1051 (N_1051,In_245,In_145);
nor U1052 (N_1052,In_257,In_717);
or U1053 (N_1053,In_1832,In_1988);
nand U1054 (N_1054,In_634,In_1532);
nor U1055 (N_1055,In_1509,In_800);
or U1056 (N_1056,In_970,In_1167);
xnor U1057 (N_1057,In_700,In_1779);
xor U1058 (N_1058,In_508,In_620);
nand U1059 (N_1059,In_1660,In_510);
nor U1060 (N_1060,In_458,In_63);
nand U1061 (N_1061,In_1486,In_155);
nor U1062 (N_1062,In_813,In_1982);
or U1063 (N_1063,In_450,In_1904);
or U1064 (N_1064,In_1184,In_1999);
or U1065 (N_1065,In_1598,In_1380);
or U1066 (N_1066,In_1891,In_359);
and U1067 (N_1067,In_1596,In_1584);
or U1068 (N_1068,In_1749,In_640);
nor U1069 (N_1069,In_868,In_699);
nor U1070 (N_1070,In_1971,In_456);
xor U1071 (N_1071,In_150,In_631);
xnor U1072 (N_1072,In_1270,In_1689);
and U1073 (N_1073,In_1202,In_441);
nand U1074 (N_1074,In_1237,In_1724);
nor U1075 (N_1075,In_976,In_619);
and U1076 (N_1076,In_1605,In_1409);
and U1077 (N_1077,In_278,In_1686);
nor U1078 (N_1078,In_1744,In_1713);
nor U1079 (N_1079,In_1002,In_398);
xnor U1080 (N_1080,In_233,In_882);
or U1081 (N_1081,In_245,In_533);
nor U1082 (N_1082,In_17,In_528);
nand U1083 (N_1083,In_1042,In_833);
nor U1084 (N_1084,In_1987,In_1305);
and U1085 (N_1085,In_135,In_1444);
and U1086 (N_1086,In_151,In_1627);
xnor U1087 (N_1087,In_1703,In_824);
and U1088 (N_1088,In_1632,In_497);
and U1089 (N_1089,In_1204,In_728);
and U1090 (N_1090,In_783,In_238);
nor U1091 (N_1091,In_191,In_1762);
and U1092 (N_1092,In_1215,In_1662);
and U1093 (N_1093,In_993,In_1745);
nand U1094 (N_1094,In_1645,In_220);
nor U1095 (N_1095,In_807,In_1139);
xor U1096 (N_1096,In_1778,In_1984);
nor U1097 (N_1097,In_1681,In_1215);
xnor U1098 (N_1098,In_1316,In_1177);
and U1099 (N_1099,In_1417,In_1902);
and U1100 (N_1100,In_1847,In_133);
and U1101 (N_1101,In_1837,In_1236);
nand U1102 (N_1102,In_338,In_1710);
nor U1103 (N_1103,In_1704,In_1375);
xor U1104 (N_1104,In_1153,In_488);
nor U1105 (N_1105,In_1928,In_897);
xor U1106 (N_1106,In_1519,In_1434);
and U1107 (N_1107,In_1009,In_1937);
or U1108 (N_1108,In_610,In_1544);
nand U1109 (N_1109,In_1866,In_26);
or U1110 (N_1110,In_1463,In_1428);
nand U1111 (N_1111,In_353,In_1771);
nand U1112 (N_1112,In_213,In_94);
nor U1113 (N_1113,In_444,In_978);
nor U1114 (N_1114,In_1065,In_1233);
and U1115 (N_1115,In_957,In_1022);
or U1116 (N_1116,In_1952,In_491);
nand U1117 (N_1117,In_1349,In_1203);
xor U1118 (N_1118,In_764,In_1817);
and U1119 (N_1119,In_410,In_834);
and U1120 (N_1120,In_1822,In_1267);
xnor U1121 (N_1121,In_1492,In_55);
and U1122 (N_1122,In_100,In_143);
or U1123 (N_1123,In_388,In_401);
or U1124 (N_1124,In_1558,In_1440);
nor U1125 (N_1125,In_524,In_1341);
or U1126 (N_1126,In_283,In_127);
nor U1127 (N_1127,In_1300,In_256);
xor U1128 (N_1128,In_909,In_1009);
nand U1129 (N_1129,In_359,In_183);
nor U1130 (N_1130,In_1279,In_132);
xor U1131 (N_1131,In_1532,In_1970);
or U1132 (N_1132,In_1738,In_959);
nand U1133 (N_1133,In_1922,In_1422);
xor U1134 (N_1134,In_737,In_62);
xor U1135 (N_1135,In_1842,In_1276);
xnor U1136 (N_1136,In_1780,In_597);
or U1137 (N_1137,In_1607,In_794);
nor U1138 (N_1138,In_492,In_1911);
nor U1139 (N_1139,In_1856,In_1522);
or U1140 (N_1140,In_1241,In_1912);
xor U1141 (N_1141,In_1665,In_1771);
xor U1142 (N_1142,In_693,In_749);
or U1143 (N_1143,In_171,In_381);
and U1144 (N_1144,In_1538,In_1058);
or U1145 (N_1145,In_1842,In_978);
or U1146 (N_1146,In_1051,In_1381);
xor U1147 (N_1147,In_1829,In_547);
and U1148 (N_1148,In_988,In_1577);
nor U1149 (N_1149,In_1375,In_1683);
xnor U1150 (N_1150,In_1212,In_1719);
xor U1151 (N_1151,In_1573,In_151);
nor U1152 (N_1152,In_1206,In_389);
nor U1153 (N_1153,In_54,In_1851);
xnor U1154 (N_1154,In_193,In_209);
xor U1155 (N_1155,In_867,In_731);
or U1156 (N_1156,In_569,In_1912);
xnor U1157 (N_1157,In_422,In_63);
or U1158 (N_1158,In_1051,In_164);
xnor U1159 (N_1159,In_729,In_51);
or U1160 (N_1160,In_1228,In_1781);
and U1161 (N_1161,In_700,In_1235);
xor U1162 (N_1162,In_1731,In_185);
nand U1163 (N_1163,In_1227,In_1549);
nor U1164 (N_1164,In_151,In_1056);
and U1165 (N_1165,In_38,In_1758);
xor U1166 (N_1166,In_448,In_1434);
or U1167 (N_1167,In_987,In_466);
nor U1168 (N_1168,In_1970,In_392);
nand U1169 (N_1169,In_1753,In_163);
xnor U1170 (N_1170,In_706,In_99);
nor U1171 (N_1171,In_1364,In_1060);
xor U1172 (N_1172,In_1478,In_1028);
nor U1173 (N_1173,In_979,In_1311);
nor U1174 (N_1174,In_1102,In_52);
and U1175 (N_1175,In_547,In_1867);
xor U1176 (N_1176,In_758,In_1068);
nand U1177 (N_1177,In_989,In_539);
or U1178 (N_1178,In_129,In_8);
xnor U1179 (N_1179,In_1484,In_914);
nor U1180 (N_1180,In_882,In_1569);
xnor U1181 (N_1181,In_772,In_1663);
and U1182 (N_1182,In_520,In_316);
nor U1183 (N_1183,In_1856,In_648);
xnor U1184 (N_1184,In_925,In_1447);
nor U1185 (N_1185,In_370,In_177);
xor U1186 (N_1186,In_1307,In_360);
or U1187 (N_1187,In_1178,In_780);
nand U1188 (N_1188,In_1851,In_361);
nor U1189 (N_1189,In_827,In_1846);
or U1190 (N_1190,In_384,In_578);
and U1191 (N_1191,In_1876,In_688);
nand U1192 (N_1192,In_609,In_1694);
xor U1193 (N_1193,In_1564,In_1210);
or U1194 (N_1194,In_103,In_195);
nor U1195 (N_1195,In_126,In_1819);
or U1196 (N_1196,In_1996,In_1502);
xnor U1197 (N_1197,In_1034,In_1403);
nand U1198 (N_1198,In_826,In_750);
or U1199 (N_1199,In_1870,In_56);
and U1200 (N_1200,In_455,In_777);
nand U1201 (N_1201,In_400,In_1782);
nor U1202 (N_1202,In_228,In_1033);
nor U1203 (N_1203,In_1265,In_1639);
and U1204 (N_1204,In_778,In_884);
and U1205 (N_1205,In_54,In_1932);
nor U1206 (N_1206,In_1728,In_1161);
nor U1207 (N_1207,In_845,In_1697);
nor U1208 (N_1208,In_1848,In_1279);
and U1209 (N_1209,In_324,In_44);
nor U1210 (N_1210,In_399,In_158);
nand U1211 (N_1211,In_463,In_562);
nand U1212 (N_1212,In_1625,In_637);
and U1213 (N_1213,In_1310,In_320);
xnor U1214 (N_1214,In_1143,In_795);
nor U1215 (N_1215,In_1986,In_1234);
nor U1216 (N_1216,In_900,In_1348);
nand U1217 (N_1217,In_990,In_489);
and U1218 (N_1218,In_1587,In_233);
and U1219 (N_1219,In_220,In_1534);
and U1220 (N_1220,In_1081,In_817);
and U1221 (N_1221,In_1675,In_587);
or U1222 (N_1222,In_1053,In_1811);
xnor U1223 (N_1223,In_686,In_1327);
nand U1224 (N_1224,In_1901,In_774);
nand U1225 (N_1225,In_1324,In_897);
xor U1226 (N_1226,In_1488,In_1218);
xnor U1227 (N_1227,In_1786,In_583);
nor U1228 (N_1228,In_1602,In_230);
nand U1229 (N_1229,In_301,In_1680);
xor U1230 (N_1230,In_449,In_1287);
and U1231 (N_1231,In_1141,In_1887);
or U1232 (N_1232,In_1918,In_1898);
nand U1233 (N_1233,In_1878,In_74);
and U1234 (N_1234,In_1861,In_1634);
nand U1235 (N_1235,In_228,In_1933);
nor U1236 (N_1236,In_182,In_947);
xnor U1237 (N_1237,In_894,In_1641);
and U1238 (N_1238,In_596,In_794);
and U1239 (N_1239,In_997,In_1228);
or U1240 (N_1240,In_634,In_43);
nand U1241 (N_1241,In_884,In_869);
nand U1242 (N_1242,In_110,In_204);
nor U1243 (N_1243,In_1515,In_193);
and U1244 (N_1244,In_635,In_134);
xnor U1245 (N_1245,In_1339,In_1857);
or U1246 (N_1246,In_122,In_219);
and U1247 (N_1247,In_573,In_1384);
xor U1248 (N_1248,In_1131,In_243);
nor U1249 (N_1249,In_1939,In_1882);
and U1250 (N_1250,In_16,In_14);
nand U1251 (N_1251,In_1687,In_1063);
xor U1252 (N_1252,In_1598,In_1966);
nor U1253 (N_1253,In_107,In_1294);
or U1254 (N_1254,In_680,In_1573);
xor U1255 (N_1255,In_1286,In_931);
or U1256 (N_1256,In_120,In_1364);
or U1257 (N_1257,In_300,In_590);
or U1258 (N_1258,In_969,In_685);
and U1259 (N_1259,In_106,In_1798);
nor U1260 (N_1260,In_499,In_1039);
xor U1261 (N_1261,In_260,In_255);
or U1262 (N_1262,In_362,In_932);
nand U1263 (N_1263,In_91,In_887);
nor U1264 (N_1264,In_1176,In_156);
nand U1265 (N_1265,In_511,In_625);
and U1266 (N_1266,In_1755,In_1047);
and U1267 (N_1267,In_1649,In_504);
and U1268 (N_1268,In_109,In_26);
nor U1269 (N_1269,In_1505,In_243);
and U1270 (N_1270,In_322,In_1718);
nand U1271 (N_1271,In_173,In_1645);
nor U1272 (N_1272,In_934,In_246);
xnor U1273 (N_1273,In_1208,In_1083);
or U1274 (N_1274,In_286,In_1510);
and U1275 (N_1275,In_69,In_140);
nor U1276 (N_1276,In_1280,In_1838);
and U1277 (N_1277,In_294,In_992);
nand U1278 (N_1278,In_1561,In_1539);
or U1279 (N_1279,In_1081,In_731);
nand U1280 (N_1280,In_340,In_792);
nor U1281 (N_1281,In_805,In_1840);
or U1282 (N_1282,In_254,In_1355);
nand U1283 (N_1283,In_618,In_412);
and U1284 (N_1284,In_659,In_971);
nor U1285 (N_1285,In_1889,In_222);
nor U1286 (N_1286,In_20,In_1977);
nor U1287 (N_1287,In_1380,In_1968);
or U1288 (N_1288,In_704,In_465);
nand U1289 (N_1289,In_404,In_1651);
or U1290 (N_1290,In_1836,In_331);
nor U1291 (N_1291,In_1292,In_1401);
nand U1292 (N_1292,In_1128,In_1486);
and U1293 (N_1293,In_1083,In_1510);
nor U1294 (N_1294,In_968,In_278);
nand U1295 (N_1295,In_1289,In_1591);
nand U1296 (N_1296,In_696,In_711);
nor U1297 (N_1297,In_94,In_434);
and U1298 (N_1298,In_908,In_914);
or U1299 (N_1299,In_133,In_613);
or U1300 (N_1300,In_1214,In_1812);
or U1301 (N_1301,In_1000,In_1540);
nor U1302 (N_1302,In_671,In_977);
nor U1303 (N_1303,In_1327,In_454);
xor U1304 (N_1304,In_1454,In_1809);
nand U1305 (N_1305,In_656,In_998);
xnor U1306 (N_1306,In_1153,In_939);
xor U1307 (N_1307,In_1947,In_1212);
or U1308 (N_1308,In_106,In_630);
nand U1309 (N_1309,In_1750,In_180);
or U1310 (N_1310,In_951,In_1663);
and U1311 (N_1311,In_411,In_796);
nor U1312 (N_1312,In_271,In_1303);
nand U1313 (N_1313,In_622,In_1083);
and U1314 (N_1314,In_576,In_1139);
xor U1315 (N_1315,In_1909,In_1099);
nor U1316 (N_1316,In_151,In_960);
nand U1317 (N_1317,In_16,In_1959);
or U1318 (N_1318,In_585,In_277);
xor U1319 (N_1319,In_1442,In_1143);
nand U1320 (N_1320,In_752,In_1994);
or U1321 (N_1321,In_537,In_916);
and U1322 (N_1322,In_163,In_1397);
and U1323 (N_1323,In_1586,In_1931);
or U1324 (N_1324,In_362,In_288);
and U1325 (N_1325,In_136,In_762);
and U1326 (N_1326,In_574,In_1088);
xnor U1327 (N_1327,In_1908,In_390);
or U1328 (N_1328,In_593,In_1415);
and U1329 (N_1329,In_172,In_1416);
nor U1330 (N_1330,In_768,In_1925);
nand U1331 (N_1331,In_1165,In_1995);
or U1332 (N_1332,In_1077,In_1336);
or U1333 (N_1333,In_1622,In_590);
or U1334 (N_1334,In_130,In_489);
xor U1335 (N_1335,In_721,In_455);
nor U1336 (N_1336,In_1852,In_348);
or U1337 (N_1337,In_1567,In_1888);
nand U1338 (N_1338,In_1463,In_175);
xnor U1339 (N_1339,In_1079,In_1685);
nor U1340 (N_1340,In_1874,In_1634);
xor U1341 (N_1341,In_1916,In_1567);
and U1342 (N_1342,In_1591,In_893);
nand U1343 (N_1343,In_916,In_107);
nand U1344 (N_1344,In_1875,In_231);
nor U1345 (N_1345,In_516,In_1111);
xor U1346 (N_1346,In_1809,In_1819);
or U1347 (N_1347,In_1592,In_1604);
or U1348 (N_1348,In_1979,In_841);
or U1349 (N_1349,In_367,In_386);
or U1350 (N_1350,In_445,In_1300);
nor U1351 (N_1351,In_115,In_938);
and U1352 (N_1352,In_425,In_525);
xor U1353 (N_1353,In_874,In_1608);
xor U1354 (N_1354,In_1328,In_558);
nand U1355 (N_1355,In_1990,In_1331);
xor U1356 (N_1356,In_281,In_713);
nor U1357 (N_1357,In_504,In_617);
nor U1358 (N_1358,In_1432,In_1558);
xnor U1359 (N_1359,In_374,In_1692);
nand U1360 (N_1360,In_1683,In_258);
xor U1361 (N_1361,In_1978,In_916);
nor U1362 (N_1362,In_776,In_1502);
or U1363 (N_1363,In_559,In_473);
and U1364 (N_1364,In_1267,In_884);
xor U1365 (N_1365,In_911,In_811);
or U1366 (N_1366,In_713,In_672);
or U1367 (N_1367,In_461,In_1469);
and U1368 (N_1368,In_1415,In_4);
or U1369 (N_1369,In_346,In_767);
xnor U1370 (N_1370,In_467,In_1007);
and U1371 (N_1371,In_671,In_1534);
xor U1372 (N_1372,In_150,In_157);
xor U1373 (N_1373,In_1165,In_661);
or U1374 (N_1374,In_1714,In_1077);
and U1375 (N_1375,In_1545,In_1030);
xor U1376 (N_1376,In_124,In_1248);
xor U1377 (N_1377,In_1958,In_278);
xor U1378 (N_1378,In_1125,In_1855);
nand U1379 (N_1379,In_1387,In_854);
or U1380 (N_1380,In_871,In_1936);
or U1381 (N_1381,In_1885,In_93);
xnor U1382 (N_1382,In_1038,In_535);
nand U1383 (N_1383,In_819,In_262);
xnor U1384 (N_1384,In_1433,In_576);
nor U1385 (N_1385,In_1805,In_404);
or U1386 (N_1386,In_1622,In_1548);
nand U1387 (N_1387,In_1859,In_962);
nor U1388 (N_1388,In_1316,In_1519);
nor U1389 (N_1389,In_1987,In_1394);
or U1390 (N_1390,In_1287,In_1255);
nor U1391 (N_1391,In_1339,In_984);
nand U1392 (N_1392,In_606,In_1423);
nand U1393 (N_1393,In_409,In_116);
and U1394 (N_1394,In_1457,In_960);
or U1395 (N_1395,In_356,In_1196);
xor U1396 (N_1396,In_1,In_1642);
xnor U1397 (N_1397,In_1841,In_1726);
or U1398 (N_1398,In_1387,In_1721);
xnor U1399 (N_1399,In_1796,In_1039);
or U1400 (N_1400,In_1781,In_1668);
and U1401 (N_1401,In_806,In_1153);
nor U1402 (N_1402,In_1504,In_637);
and U1403 (N_1403,In_421,In_817);
nand U1404 (N_1404,In_77,In_1370);
xnor U1405 (N_1405,In_1820,In_1287);
xnor U1406 (N_1406,In_812,In_951);
nand U1407 (N_1407,In_1847,In_542);
nor U1408 (N_1408,In_1268,In_1788);
nor U1409 (N_1409,In_1444,In_779);
nand U1410 (N_1410,In_1221,In_1513);
xnor U1411 (N_1411,In_1157,In_1035);
nand U1412 (N_1412,In_1994,In_1499);
xnor U1413 (N_1413,In_1542,In_804);
xor U1414 (N_1414,In_1514,In_1212);
nor U1415 (N_1415,In_450,In_1438);
nor U1416 (N_1416,In_416,In_552);
nand U1417 (N_1417,In_1554,In_1107);
and U1418 (N_1418,In_1192,In_436);
and U1419 (N_1419,In_19,In_1655);
and U1420 (N_1420,In_270,In_1453);
xnor U1421 (N_1421,In_191,In_72);
nand U1422 (N_1422,In_1011,In_633);
xor U1423 (N_1423,In_1077,In_1109);
nand U1424 (N_1424,In_460,In_94);
nand U1425 (N_1425,In_1150,In_1780);
nor U1426 (N_1426,In_546,In_1606);
or U1427 (N_1427,In_314,In_806);
nor U1428 (N_1428,In_1226,In_1093);
nor U1429 (N_1429,In_1760,In_1295);
or U1430 (N_1430,In_1256,In_498);
and U1431 (N_1431,In_642,In_108);
and U1432 (N_1432,In_1020,In_1419);
nand U1433 (N_1433,In_1143,In_1519);
and U1434 (N_1434,In_599,In_1081);
nor U1435 (N_1435,In_460,In_1989);
nand U1436 (N_1436,In_1612,In_1713);
or U1437 (N_1437,In_871,In_726);
xor U1438 (N_1438,In_837,In_1740);
nand U1439 (N_1439,In_1528,In_723);
and U1440 (N_1440,In_1942,In_1857);
or U1441 (N_1441,In_194,In_545);
or U1442 (N_1442,In_1039,In_362);
nand U1443 (N_1443,In_183,In_91);
xnor U1444 (N_1444,In_1024,In_208);
nor U1445 (N_1445,In_676,In_1357);
or U1446 (N_1446,In_869,In_697);
nor U1447 (N_1447,In_180,In_344);
or U1448 (N_1448,In_369,In_785);
and U1449 (N_1449,In_854,In_1523);
nor U1450 (N_1450,In_1576,In_46);
and U1451 (N_1451,In_1002,In_678);
xor U1452 (N_1452,In_742,In_603);
xor U1453 (N_1453,In_538,In_1184);
and U1454 (N_1454,In_592,In_266);
or U1455 (N_1455,In_825,In_1761);
xnor U1456 (N_1456,In_1328,In_45);
or U1457 (N_1457,In_966,In_14);
nand U1458 (N_1458,In_396,In_1106);
nor U1459 (N_1459,In_11,In_964);
or U1460 (N_1460,In_1757,In_1764);
or U1461 (N_1461,In_1313,In_1223);
or U1462 (N_1462,In_760,In_877);
or U1463 (N_1463,In_1431,In_108);
xnor U1464 (N_1464,In_491,In_1001);
and U1465 (N_1465,In_1138,In_1360);
nand U1466 (N_1466,In_892,In_1609);
nor U1467 (N_1467,In_1325,In_1766);
xor U1468 (N_1468,In_1533,In_375);
nor U1469 (N_1469,In_685,In_152);
and U1470 (N_1470,In_899,In_1969);
nor U1471 (N_1471,In_718,In_169);
and U1472 (N_1472,In_563,In_1243);
and U1473 (N_1473,In_763,In_1153);
and U1474 (N_1474,In_1468,In_353);
or U1475 (N_1475,In_515,In_1356);
and U1476 (N_1476,In_1221,In_912);
nor U1477 (N_1477,In_614,In_857);
xor U1478 (N_1478,In_1041,In_1209);
nand U1479 (N_1479,In_677,In_359);
and U1480 (N_1480,In_538,In_1350);
xnor U1481 (N_1481,In_639,In_1209);
nor U1482 (N_1482,In_932,In_831);
nand U1483 (N_1483,In_974,In_1647);
xor U1484 (N_1484,In_1543,In_443);
nor U1485 (N_1485,In_1414,In_645);
or U1486 (N_1486,In_1257,In_1212);
and U1487 (N_1487,In_725,In_1722);
xor U1488 (N_1488,In_1439,In_1712);
xor U1489 (N_1489,In_417,In_1278);
nor U1490 (N_1490,In_175,In_1244);
or U1491 (N_1491,In_2,In_421);
or U1492 (N_1492,In_1278,In_457);
xor U1493 (N_1493,In_32,In_26);
nor U1494 (N_1494,In_48,In_1126);
xor U1495 (N_1495,In_69,In_1399);
or U1496 (N_1496,In_32,In_1964);
nand U1497 (N_1497,In_1612,In_1043);
or U1498 (N_1498,In_1035,In_1829);
or U1499 (N_1499,In_1605,In_1108);
or U1500 (N_1500,In_72,In_1138);
nand U1501 (N_1501,In_690,In_1298);
or U1502 (N_1502,In_1449,In_1237);
or U1503 (N_1503,In_1137,In_1848);
or U1504 (N_1504,In_1836,In_436);
nand U1505 (N_1505,In_1000,In_541);
and U1506 (N_1506,In_794,In_449);
and U1507 (N_1507,In_1299,In_342);
and U1508 (N_1508,In_1247,In_1492);
nor U1509 (N_1509,In_1691,In_636);
nor U1510 (N_1510,In_1113,In_1619);
or U1511 (N_1511,In_688,In_300);
and U1512 (N_1512,In_983,In_1226);
xnor U1513 (N_1513,In_1196,In_280);
xnor U1514 (N_1514,In_1790,In_393);
nand U1515 (N_1515,In_760,In_1239);
and U1516 (N_1516,In_1037,In_1175);
or U1517 (N_1517,In_899,In_251);
nor U1518 (N_1518,In_1020,In_227);
xnor U1519 (N_1519,In_1648,In_1018);
nor U1520 (N_1520,In_941,In_1017);
or U1521 (N_1521,In_1517,In_565);
or U1522 (N_1522,In_1725,In_1125);
nand U1523 (N_1523,In_1174,In_1771);
xor U1524 (N_1524,In_85,In_1858);
and U1525 (N_1525,In_1367,In_1472);
and U1526 (N_1526,In_1517,In_1173);
xnor U1527 (N_1527,In_1383,In_1169);
nor U1528 (N_1528,In_1516,In_229);
nand U1529 (N_1529,In_1115,In_736);
nand U1530 (N_1530,In_1365,In_1221);
nand U1531 (N_1531,In_567,In_1426);
xor U1532 (N_1532,In_1423,In_1651);
or U1533 (N_1533,In_1914,In_405);
nor U1534 (N_1534,In_426,In_1592);
nor U1535 (N_1535,In_847,In_1376);
nand U1536 (N_1536,In_340,In_1042);
nor U1537 (N_1537,In_575,In_1514);
and U1538 (N_1538,In_1683,In_409);
nand U1539 (N_1539,In_1437,In_703);
nand U1540 (N_1540,In_1010,In_99);
nand U1541 (N_1541,In_508,In_379);
nor U1542 (N_1542,In_968,In_928);
nor U1543 (N_1543,In_735,In_561);
or U1544 (N_1544,In_901,In_1762);
nor U1545 (N_1545,In_1198,In_477);
nand U1546 (N_1546,In_544,In_17);
or U1547 (N_1547,In_848,In_1980);
and U1548 (N_1548,In_1490,In_116);
xor U1549 (N_1549,In_1523,In_892);
or U1550 (N_1550,In_611,In_1754);
nor U1551 (N_1551,In_1512,In_502);
or U1552 (N_1552,In_394,In_1941);
xnor U1553 (N_1553,In_713,In_1499);
or U1554 (N_1554,In_1892,In_808);
xnor U1555 (N_1555,In_355,In_1694);
nand U1556 (N_1556,In_995,In_880);
and U1557 (N_1557,In_213,In_882);
nand U1558 (N_1558,In_160,In_405);
xnor U1559 (N_1559,In_216,In_642);
nor U1560 (N_1560,In_1784,In_1487);
or U1561 (N_1561,In_950,In_809);
xor U1562 (N_1562,In_29,In_1736);
nand U1563 (N_1563,In_337,In_173);
or U1564 (N_1564,In_1744,In_276);
nor U1565 (N_1565,In_1488,In_512);
nand U1566 (N_1566,In_995,In_1892);
and U1567 (N_1567,In_326,In_1942);
xor U1568 (N_1568,In_783,In_577);
xnor U1569 (N_1569,In_784,In_86);
xnor U1570 (N_1570,In_1372,In_38);
and U1571 (N_1571,In_1667,In_1849);
xnor U1572 (N_1572,In_1935,In_485);
and U1573 (N_1573,In_1157,In_1790);
xor U1574 (N_1574,In_1210,In_737);
or U1575 (N_1575,In_1960,In_1915);
nand U1576 (N_1576,In_1005,In_1095);
nor U1577 (N_1577,In_1860,In_1185);
nor U1578 (N_1578,In_1142,In_773);
xor U1579 (N_1579,In_1240,In_1125);
and U1580 (N_1580,In_1323,In_393);
xnor U1581 (N_1581,In_1155,In_1919);
or U1582 (N_1582,In_911,In_890);
nand U1583 (N_1583,In_870,In_1351);
xnor U1584 (N_1584,In_1328,In_1742);
xnor U1585 (N_1585,In_72,In_104);
nand U1586 (N_1586,In_156,In_715);
nor U1587 (N_1587,In_1955,In_343);
xor U1588 (N_1588,In_1746,In_539);
xor U1589 (N_1589,In_98,In_1167);
nor U1590 (N_1590,In_1686,In_1622);
or U1591 (N_1591,In_790,In_1610);
xor U1592 (N_1592,In_232,In_1553);
xor U1593 (N_1593,In_235,In_291);
and U1594 (N_1594,In_1231,In_1483);
or U1595 (N_1595,In_525,In_187);
nor U1596 (N_1596,In_942,In_1078);
and U1597 (N_1597,In_1452,In_1388);
xnor U1598 (N_1598,In_276,In_1006);
nor U1599 (N_1599,In_972,In_270);
nand U1600 (N_1600,In_1054,In_43);
nor U1601 (N_1601,In_1070,In_467);
nor U1602 (N_1602,In_157,In_1947);
and U1603 (N_1603,In_1763,In_1881);
nor U1604 (N_1604,In_1328,In_547);
nand U1605 (N_1605,In_1286,In_1838);
and U1606 (N_1606,In_1379,In_1073);
and U1607 (N_1607,In_1614,In_1539);
nor U1608 (N_1608,In_1681,In_1267);
xnor U1609 (N_1609,In_1627,In_1096);
nand U1610 (N_1610,In_1548,In_1899);
nand U1611 (N_1611,In_1220,In_704);
or U1612 (N_1612,In_605,In_1315);
xnor U1613 (N_1613,In_678,In_97);
xnor U1614 (N_1614,In_1511,In_1851);
nand U1615 (N_1615,In_352,In_600);
xor U1616 (N_1616,In_1528,In_1570);
nand U1617 (N_1617,In_427,In_874);
nand U1618 (N_1618,In_604,In_1073);
xnor U1619 (N_1619,In_1045,In_1349);
and U1620 (N_1620,In_1601,In_1489);
or U1621 (N_1621,In_510,In_1520);
nor U1622 (N_1622,In_302,In_84);
nor U1623 (N_1623,In_1024,In_517);
nor U1624 (N_1624,In_366,In_549);
nand U1625 (N_1625,In_1214,In_649);
nor U1626 (N_1626,In_1927,In_282);
or U1627 (N_1627,In_749,In_1283);
or U1628 (N_1628,In_927,In_36);
xnor U1629 (N_1629,In_383,In_1860);
and U1630 (N_1630,In_1417,In_690);
and U1631 (N_1631,In_1513,In_766);
nor U1632 (N_1632,In_31,In_1888);
or U1633 (N_1633,In_298,In_1768);
and U1634 (N_1634,In_1154,In_369);
nand U1635 (N_1635,In_103,In_695);
or U1636 (N_1636,In_1893,In_1126);
nor U1637 (N_1637,In_1385,In_417);
xor U1638 (N_1638,In_1161,In_388);
nand U1639 (N_1639,In_929,In_73);
or U1640 (N_1640,In_111,In_207);
or U1641 (N_1641,In_1414,In_94);
nor U1642 (N_1642,In_1003,In_1960);
xor U1643 (N_1643,In_46,In_1516);
nand U1644 (N_1644,In_1525,In_154);
xor U1645 (N_1645,In_1839,In_688);
nand U1646 (N_1646,In_1468,In_162);
nand U1647 (N_1647,In_1821,In_1399);
and U1648 (N_1648,In_537,In_576);
or U1649 (N_1649,In_261,In_574);
and U1650 (N_1650,In_1953,In_1415);
and U1651 (N_1651,In_875,In_363);
nand U1652 (N_1652,In_957,In_1080);
and U1653 (N_1653,In_283,In_301);
nor U1654 (N_1654,In_1400,In_1676);
and U1655 (N_1655,In_460,In_254);
and U1656 (N_1656,In_103,In_1384);
nand U1657 (N_1657,In_443,In_1652);
and U1658 (N_1658,In_889,In_1895);
nor U1659 (N_1659,In_1113,In_1387);
and U1660 (N_1660,In_1135,In_893);
and U1661 (N_1661,In_1017,In_48);
or U1662 (N_1662,In_1719,In_1237);
or U1663 (N_1663,In_955,In_1352);
nand U1664 (N_1664,In_252,In_1081);
nor U1665 (N_1665,In_1739,In_1294);
xor U1666 (N_1666,In_800,In_136);
xnor U1667 (N_1667,In_1369,In_1564);
and U1668 (N_1668,In_1048,In_1280);
xnor U1669 (N_1669,In_1467,In_396);
nand U1670 (N_1670,In_1960,In_834);
or U1671 (N_1671,In_642,In_249);
xor U1672 (N_1672,In_1362,In_895);
or U1673 (N_1673,In_1336,In_1153);
nand U1674 (N_1674,In_559,In_646);
nor U1675 (N_1675,In_123,In_601);
nand U1676 (N_1676,In_1430,In_430);
nor U1677 (N_1677,In_1388,In_555);
and U1678 (N_1678,In_757,In_795);
and U1679 (N_1679,In_930,In_1536);
and U1680 (N_1680,In_1221,In_535);
and U1681 (N_1681,In_621,In_982);
nor U1682 (N_1682,In_1302,In_1523);
nor U1683 (N_1683,In_906,In_501);
and U1684 (N_1684,In_1817,In_1488);
xnor U1685 (N_1685,In_1142,In_398);
xnor U1686 (N_1686,In_521,In_1353);
or U1687 (N_1687,In_641,In_1059);
and U1688 (N_1688,In_1906,In_395);
or U1689 (N_1689,In_1295,In_1802);
nor U1690 (N_1690,In_1477,In_1270);
nor U1691 (N_1691,In_507,In_1191);
nand U1692 (N_1692,In_282,In_1955);
xnor U1693 (N_1693,In_1157,In_1651);
xor U1694 (N_1694,In_1012,In_51);
nand U1695 (N_1695,In_747,In_1025);
xor U1696 (N_1696,In_482,In_47);
nand U1697 (N_1697,In_1163,In_1921);
and U1698 (N_1698,In_838,In_1931);
and U1699 (N_1699,In_1216,In_1639);
xor U1700 (N_1700,In_869,In_115);
or U1701 (N_1701,In_767,In_112);
and U1702 (N_1702,In_107,In_14);
or U1703 (N_1703,In_1206,In_1003);
nand U1704 (N_1704,In_965,In_602);
and U1705 (N_1705,In_741,In_531);
or U1706 (N_1706,In_1983,In_507);
nand U1707 (N_1707,In_1773,In_1990);
or U1708 (N_1708,In_1144,In_1038);
or U1709 (N_1709,In_1225,In_600);
nor U1710 (N_1710,In_395,In_1958);
nor U1711 (N_1711,In_498,In_777);
nor U1712 (N_1712,In_27,In_1520);
or U1713 (N_1713,In_1366,In_313);
nor U1714 (N_1714,In_1754,In_1421);
nor U1715 (N_1715,In_1613,In_353);
nor U1716 (N_1716,In_573,In_298);
or U1717 (N_1717,In_1737,In_1804);
nand U1718 (N_1718,In_853,In_1393);
or U1719 (N_1719,In_1655,In_480);
nand U1720 (N_1720,In_273,In_533);
or U1721 (N_1721,In_702,In_1304);
nand U1722 (N_1722,In_699,In_346);
and U1723 (N_1723,In_400,In_252);
nor U1724 (N_1724,In_631,In_468);
nor U1725 (N_1725,In_307,In_1149);
xnor U1726 (N_1726,In_1866,In_836);
nand U1727 (N_1727,In_1012,In_1759);
xnor U1728 (N_1728,In_812,In_1459);
or U1729 (N_1729,In_72,In_893);
or U1730 (N_1730,In_754,In_426);
nand U1731 (N_1731,In_1703,In_1415);
xnor U1732 (N_1732,In_1930,In_497);
and U1733 (N_1733,In_1850,In_597);
nand U1734 (N_1734,In_1287,In_634);
nor U1735 (N_1735,In_1835,In_733);
and U1736 (N_1736,In_250,In_338);
xor U1737 (N_1737,In_362,In_828);
or U1738 (N_1738,In_336,In_50);
xor U1739 (N_1739,In_1037,In_393);
nor U1740 (N_1740,In_1770,In_419);
or U1741 (N_1741,In_140,In_141);
and U1742 (N_1742,In_301,In_1569);
and U1743 (N_1743,In_78,In_515);
nor U1744 (N_1744,In_288,In_1136);
nand U1745 (N_1745,In_1533,In_513);
nor U1746 (N_1746,In_650,In_935);
nor U1747 (N_1747,In_862,In_364);
nand U1748 (N_1748,In_465,In_628);
and U1749 (N_1749,In_1319,In_470);
and U1750 (N_1750,In_1226,In_343);
nand U1751 (N_1751,In_1625,In_1946);
xnor U1752 (N_1752,In_725,In_258);
and U1753 (N_1753,In_412,In_537);
or U1754 (N_1754,In_1061,In_1334);
nand U1755 (N_1755,In_860,In_1355);
nor U1756 (N_1756,In_755,In_206);
nor U1757 (N_1757,In_572,In_1527);
nand U1758 (N_1758,In_1581,In_1810);
or U1759 (N_1759,In_1010,In_1839);
xnor U1760 (N_1760,In_1665,In_946);
or U1761 (N_1761,In_1254,In_1307);
or U1762 (N_1762,In_1353,In_1004);
nand U1763 (N_1763,In_1393,In_700);
xor U1764 (N_1764,In_1028,In_1206);
nor U1765 (N_1765,In_362,In_1700);
nand U1766 (N_1766,In_1609,In_691);
or U1767 (N_1767,In_815,In_205);
or U1768 (N_1768,In_266,In_139);
nor U1769 (N_1769,In_225,In_621);
nor U1770 (N_1770,In_1804,In_896);
nor U1771 (N_1771,In_1825,In_1762);
or U1772 (N_1772,In_1532,In_1345);
or U1773 (N_1773,In_1088,In_1829);
and U1774 (N_1774,In_1148,In_1842);
and U1775 (N_1775,In_1783,In_376);
nand U1776 (N_1776,In_114,In_1318);
nor U1777 (N_1777,In_313,In_1776);
and U1778 (N_1778,In_263,In_1038);
xnor U1779 (N_1779,In_995,In_1504);
and U1780 (N_1780,In_764,In_536);
or U1781 (N_1781,In_782,In_1884);
or U1782 (N_1782,In_1571,In_1331);
and U1783 (N_1783,In_63,In_1372);
and U1784 (N_1784,In_438,In_1622);
and U1785 (N_1785,In_1408,In_1594);
nor U1786 (N_1786,In_1140,In_913);
nor U1787 (N_1787,In_735,In_1828);
nor U1788 (N_1788,In_1835,In_1652);
nand U1789 (N_1789,In_1337,In_142);
xor U1790 (N_1790,In_80,In_1806);
xnor U1791 (N_1791,In_1892,In_1038);
or U1792 (N_1792,In_1780,In_580);
and U1793 (N_1793,In_1103,In_628);
or U1794 (N_1794,In_1829,In_806);
and U1795 (N_1795,In_521,In_995);
nor U1796 (N_1796,In_275,In_770);
nand U1797 (N_1797,In_365,In_633);
or U1798 (N_1798,In_1601,In_65);
or U1799 (N_1799,In_261,In_1462);
nand U1800 (N_1800,In_1389,In_1874);
xor U1801 (N_1801,In_1296,In_793);
xnor U1802 (N_1802,In_41,In_250);
xnor U1803 (N_1803,In_726,In_1962);
xor U1804 (N_1804,In_305,In_1450);
xnor U1805 (N_1805,In_548,In_1561);
nand U1806 (N_1806,In_473,In_404);
or U1807 (N_1807,In_84,In_1312);
xnor U1808 (N_1808,In_1623,In_1502);
nor U1809 (N_1809,In_1314,In_743);
nor U1810 (N_1810,In_1315,In_22);
nand U1811 (N_1811,In_1421,In_1101);
nor U1812 (N_1812,In_1734,In_426);
nor U1813 (N_1813,In_128,In_331);
or U1814 (N_1814,In_1401,In_437);
and U1815 (N_1815,In_984,In_1720);
and U1816 (N_1816,In_983,In_593);
xor U1817 (N_1817,In_1431,In_1235);
and U1818 (N_1818,In_1986,In_1396);
or U1819 (N_1819,In_1259,In_77);
or U1820 (N_1820,In_1638,In_1491);
or U1821 (N_1821,In_690,In_1763);
or U1822 (N_1822,In_31,In_702);
xor U1823 (N_1823,In_613,In_751);
and U1824 (N_1824,In_621,In_1524);
nor U1825 (N_1825,In_55,In_1164);
nor U1826 (N_1826,In_1552,In_437);
and U1827 (N_1827,In_1529,In_1655);
and U1828 (N_1828,In_1474,In_947);
nand U1829 (N_1829,In_234,In_858);
nand U1830 (N_1830,In_986,In_705);
or U1831 (N_1831,In_444,In_244);
nand U1832 (N_1832,In_566,In_1571);
and U1833 (N_1833,In_849,In_541);
or U1834 (N_1834,In_1532,In_314);
nor U1835 (N_1835,In_1881,In_757);
nand U1836 (N_1836,In_582,In_1116);
and U1837 (N_1837,In_124,In_1010);
xor U1838 (N_1838,In_909,In_861);
nand U1839 (N_1839,In_1150,In_1701);
nand U1840 (N_1840,In_1913,In_308);
and U1841 (N_1841,In_287,In_161);
and U1842 (N_1842,In_804,In_980);
and U1843 (N_1843,In_1882,In_1421);
and U1844 (N_1844,In_739,In_1971);
and U1845 (N_1845,In_606,In_1228);
xnor U1846 (N_1846,In_1893,In_1041);
or U1847 (N_1847,In_1602,In_1165);
xnor U1848 (N_1848,In_794,In_906);
nor U1849 (N_1849,In_947,In_3);
and U1850 (N_1850,In_802,In_353);
nor U1851 (N_1851,In_473,In_944);
or U1852 (N_1852,In_1634,In_409);
and U1853 (N_1853,In_900,In_435);
or U1854 (N_1854,In_1048,In_701);
nand U1855 (N_1855,In_179,In_1044);
or U1856 (N_1856,In_1293,In_1586);
or U1857 (N_1857,In_759,In_1213);
xor U1858 (N_1858,In_885,In_588);
xor U1859 (N_1859,In_291,In_646);
or U1860 (N_1860,In_477,In_483);
nand U1861 (N_1861,In_561,In_1532);
xnor U1862 (N_1862,In_1440,In_882);
or U1863 (N_1863,In_605,In_434);
nor U1864 (N_1864,In_1298,In_734);
nor U1865 (N_1865,In_118,In_424);
nand U1866 (N_1866,In_820,In_1913);
xor U1867 (N_1867,In_1381,In_299);
nand U1868 (N_1868,In_1976,In_1376);
and U1869 (N_1869,In_930,In_1155);
or U1870 (N_1870,In_606,In_1003);
nand U1871 (N_1871,In_574,In_1639);
or U1872 (N_1872,In_188,In_1294);
xor U1873 (N_1873,In_471,In_576);
xnor U1874 (N_1874,In_246,In_11);
or U1875 (N_1875,In_23,In_1352);
and U1876 (N_1876,In_701,In_21);
nor U1877 (N_1877,In_137,In_425);
xor U1878 (N_1878,In_440,In_1119);
xnor U1879 (N_1879,In_847,In_1683);
xor U1880 (N_1880,In_998,In_1403);
xor U1881 (N_1881,In_1572,In_645);
nand U1882 (N_1882,In_791,In_675);
and U1883 (N_1883,In_1734,In_300);
and U1884 (N_1884,In_1699,In_1602);
nand U1885 (N_1885,In_140,In_113);
and U1886 (N_1886,In_729,In_1754);
xnor U1887 (N_1887,In_720,In_1502);
xnor U1888 (N_1888,In_368,In_1892);
nor U1889 (N_1889,In_1738,In_1080);
and U1890 (N_1890,In_379,In_1547);
or U1891 (N_1891,In_975,In_732);
and U1892 (N_1892,In_581,In_1632);
xor U1893 (N_1893,In_1205,In_381);
nand U1894 (N_1894,In_1533,In_1607);
and U1895 (N_1895,In_1766,In_840);
nor U1896 (N_1896,In_1903,In_959);
and U1897 (N_1897,In_347,In_424);
xnor U1898 (N_1898,In_1142,In_519);
and U1899 (N_1899,In_655,In_260);
nor U1900 (N_1900,In_1317,In_1782);
nand U1901 (N_1901,In_1142,In_27);
or U1902 (N_1902,In_1078,In_990);
nor U1903 (N_1903,In_162,In_31);
nor U1904 (N_1904,In_259,In_597);
or U1905 (N_1905,In_369,In_390);
nand U1906 (N_1906,In_946,In_642);
nor U1907 (N_1907,In_1764,In_405);
xor U1908 (N_1908,In_507,In_1770);
nand U1909 (N_1909,In_1714,In_1398);
nand U1910 (N_1910,In_499,In_408);
xnor U1911 (N_1911,In_328,In_201);
xor U1912 (N_1912,In_649,In_1003);
or U1913 (N_1913,In_1798,In_477);
xnor U1914 (N_1914,In_1102,In_516);
or U1915 (N_1915,In_1397,In_343);
and U1916 (N_1916,In_384,In_1549);
and U1917 (N_1917,In_1056,In_1081);
or U1918 (N_1918,In_971,In_1249);
and U1919 (N_1919,In_1032,In_433);
or U1920 (N_1920,In_818,In_1512);
xor U1921 (N_1921,In_1504,In_1633);
nand U1922 (N_1922,In_1223,In_1215);
and U1923 (N_1923,In_1048,In_71);
or U1924 (N_1924,In_47,In_1789);
nor U1925 (N_1925,In_1336,In_1211);
or U1926 (N_1926,In_392,In_141);
and U1927 (N_1927,In_1425,In_1275);
or U1928 (N_1928,In_1143,In_375);
or U1929 (N_1929,In_433,In_1763);
and U1930 (N_1930,In_869,In_1593);
nor U1931 (N_1931,In_1158,In_414);
or U1932 (N_1932,In_1891,In_372);
or U1933 (N_1933,In_150,In_742);
nand U1934 (N_1934,In_978,In_1583);
xnor U1935 (N_1935,In_1743,In_710);
nor U1936 (N_1936,In_1597,In_546);
xor U1937 (N_1937,In_670,In_898);
and U1938 (N_1938,In_1839,In_546);
or U1939 (N_1939,In_1311,In_289);
nor U1940 (N_1940,In_1678,In_1715);
nand U1941 (N_1941,In_396,In_548);
and U1942 (N_1942,In_1238,In_1891);
nand U1943 (N_1943,In_1663,In_51);
nand U1944 (N_1944,In_1740,In_1607);
or U1945 (N_1945,In_228,In_1577);
or U1946 (N_1946,In_1786,In_1024);
or U1947 (N_1947,In_592,In_1447);
xor U1948 (N_1948,In_542,In_328);
and U1949 (N_1949,In_681,In_1874);
or U1950 (N_1950,In_779,In_16);
nor U1951 (N_1951,In_330,In_1167);
nor U1952 (N_1952,In_1596,In_1613);
nand U1953 (N_1953,In_1010,In_1744);
nor U1954 (N_1954,In_891,In_1993);
nor U1955 (N_1955,In_569,In_1031);
xnor U1956 (N_1956,In_1414,In_1421);
and U1957 (N_1957,In_1643,In_1657);
nand U1958 (N_1958,In_625,In_668);
and U1959 (N_1959,In_1587,In_470);
xor U1960 (N_1960,In_1590,In_1223);
nor U1961 (N_1961,In_1347,In_1724);
or U1962 (N_1962,In_1629,In_1942);
or U1963 (N_1963,In_1221,In_1057);
xor U1964 (N_1964,In_767,In_747);
nand U1965 (N_1965,In_1447,In_1504);
nand U1966 (N_1966,In_1806,In_1880);
xnor U1967 (N_1967,In_157,In_1960);
nor U1968 (N_1968,In_573,In_1097);
and U1969 (N_1969,In_734,In_1035);
nand U1970 (N_1970,In_1104,In_1809);
nor U1971 (N_1971,In_160,In_1596);
nor U1972 (N_1972,In_1285,In_1950);
or U1973 (N_1973,In_662,In_1101);
nor U1974 (N_1974,In_1539,In_1012);
or U1975 (N_1975,In_815,In_707);
xnor U1976 (N_1976,In_299,In_151);
nor U1977 (N_1977,In_44,In_1233);
and U1978 (N_1978,In_251,In_328);
or U1979 (N_1979,In_572,In_894);
xnor U1980 (N_1980,In_1239,In_91);
nor U1981 (N_1981,In_1377,In_461);
xor U1982 (N_1982,In_835,In_1728);
nand U1983 (N_1983,In_1865,In_1390);
or U1984 (N_1984,In_811,In_244);
xor U1985 (N_1985,In_1673,In_723);
nor U1986 (N_1986,In_862,In_615);
xnor U1987 (N_1987,In_398,In_159);
or U1988 (N_1988,In_1632,In_1188);
nand U1989 (N_1989,In_813,In_761);
nand U1990 (N_1990,In_1700,In_1850);
or U1991 (N_1991,In_690,In_255);
nor U1992 (N_1992,In_950,In_128);
and U1993 (N_1993,In_1166,In_1031);
and U1994 (N_1994,In_1369,In_728);
nand U1995 (N_1995,In_1161,In_266);
xor U1996 (N_1996,In_576,In_762);
or U1997 (N_1997,In_337,In_1141);
or U1998 (N_1998,In_241,In_1999);
and U1999 (N_1999,In_1679,In_37);
xnor U2000 (N_2000,In_720,In_1917);
nand U2001 (N_2001,In_990,In_12);
xnor U2002 (N_2002,In_972,In_1018);
and U2003 (N_2003,In_1503,In_1629);
xnor U2004 (N_2004,In_1809,In_1450);
xor U2005 (N_2005,In_1326,In_1822);
or U2006 (N_2006,In_1892,In_1235);
nor U2007 (N_2007,In_1464,In_1990);
or U2008 (N_2008,In_30,In_1547);
and U2009 (N_2009,In_4,In_1772);
xor U2010 (N_2010,In_367,In_1028);
and U2011 (N_2011,In_460,In_1612);
xnor U2012 (N_2012,In_1343,In_764);
or U2013 (N_2013,In_1041,In_1664);
and U2014 (N_2014,In_323,In_211);
and U2015 (N_2015,In_1085,In_1159);
or U2016 (N_2016,In_1620,In_460);
xor U2017 (N_2017,In_595,In_1013);
or U2018 (N_2018,In_1,In_535);
nor U2019 (N_2019,In_674,In_1305);
xor U2020 (N_2020,In_1692,In_355);
xnor U2021 (N_2021,In_250,In_1834);
and U2022 (N_2022,In_1685,In_1113);
and U2023 (N_2023,In_815,In_170);
nor U2024 (N_2024,In_705,In_1235);
and U2025 (N_2025,In_662,In_227);
xnor U2026 (N_2026,In_1954,In_1763);
nor U2027 (N_2027,In_227,In_1323);
nor U2028 (N_2028,In_74,In_50);
and U2029 (N_2029,In_1284,In_399);
or U2030 (N_2030,In_56,In_163);
nand U2031 (N_2031,In_430,In_1682);
and U2032 (N_2032,In_1287,In_383);
and U2033 (N_2033,In_567,In_15);
or U2034 (N_2034,In_623,In_1698);
nand U2035 (N_2035,In_687,In_1417);
nor U2036 (N_2036,In_13,In_1055);
nor U2037 (N_2037,In_117,In_470);
and U2038 (N_2038,In_1790,In_596);
nor U2039 (N_2039,In_1017,In_1298);
nor U2040 (N_2040,In_1276,In_1073);
xnor U2041 (N_2041,In_626,In_1915);
nor U2042 (N_2042,In_730,In_1388);
xnor U2043 (N_2043,In_174,In_1457);
or U2044 (N_2044,In_677,In_1622);
and U2045 (N_2045,In_1512,In_1906);
and U2046 (N_2046,In_1865,In_1867);
nor U2047 (N_2047,In_293,In_1181);
xor U2048 (N_2048,In_1162,In_248);
or U2049 (N_2049,In_1374,In_780);
nor U2050 (N_2050,In_34,In_1148);
nand U2051 (N_2051,In_1883,In_475);
or U2052 (N_2052,In_952,In_841);
or U2053 (N_2053,In_326,In_955);
or U2054 (N_2054,In_42,In_648);
nor U2055 (N_2055,In_1533,In_1336);
and U2056 (N_2056,In_1710,In_1676);
nand U2057 (N_2057,In_1678,In_786);
or U2058 (N_2058,In_408,In_1601);
or U2059 (N_2059,In_981,In_1747);
nor U2060 (N_2060,In_850,In_9);
and U2061 (N_2061,In_753,In_1088);
and U2062 (N_2062,In_1561,In_1878);
or U2063 (N_2063,In_176,In_1445);
nand U2064 (N_2064,In_423,In_1051);
or U2065 (N_2065,In_1296,In_99);
nor U2066 (N_2066,In_1543,In_1757);
nand U2067 (N_2067,In_552,In_1075);
xnor U2068 (N_2068,In_900,In_1892);
nand U2069 (N_2069,In_1133,In_408);
or U2070 (N_2070,In_703,In_91);
nor U2071 (N_2071,In_1759,In_109);
nor U2072 (N_2072,In_1882,In_1587);
or U2073 (N_2073,In_746,In_1969);
xor U2074 (N_2074,In_936,In_1115);
nand U2075 (N_2075,In_602,In_95);
xnor U2076 (N_2076,In_507,In_1469);
nor U2077 (N_2077,In_938,In_1567);
or U2078 (N_2078,In_508,In_390);
or U2079 (N_2079,In_951,In_50);
nor U2080 (N_2080,In_1274,In_675);
and U2081 (N_2081,In_389,In_1033);
and U2082 (N_2082,In_1079,In_610);
nand U2083 (N_2083,In_565,In_1041);
xor U2084 (N_2084,In_1575,In_1409);
nand U2085 (N_2085,In_1681,In_13);
nand U2086 (N_2086,In_1700,In_1276);
and U2087 (N_2087,In_1513,In_1668);
xnor U2088 (N_2088,In_606,In_1664);
or U2089 (N_2089,In_583,In_315);
nand U2090 (N_2090,In_1420,In_914);
xnor U2091 (N_2091,In_1023,In_732);
nand U2092 (N_2092,In_846,In_1160);
xnor U2093 (N_2093,In_197,In_1448);
xor U2094 (N_2094,In_221,In_1658);
nand U2095 (N_2095,In_1382,In_78);
and U2096 (N_2096,In_1242,In_480);
nor U2097 (N_2097,In_786,In_894);
or U2098 (N_2098,In_279,In_17);
nand U2099 (N_2099,In_1041,In_1373);
and U2100 (N_2100,In_1866,In_1413);
and U2101 (N_2101,In_12,In_836);
xor U2102 (N_2102,In_1874,In_838);
nand U2103 (N_2103,In_505,In_656);
nand U2104 (N_2104,In_1540,In_1043);
nor U2105 (N_2105,In_49,In_1767);
nor U2106 (N_2106,In_243,In_644);
nor U2107 (N_2107,In_332,In_19);
xnor U2108 (N_2108,In_710,In_1338);
or U2109 (N_2109,In_1906,In_906);
and U2110 (N_2110,In_556,In_1953);
nor U2111 (N_2111,In_1631,In_163);
nand U2112 (N_2112,In_694,In_1406);
xnor U2113 (N_2113,In_517,In_1809);
or U2114 (N_2114,In_394,In_1292);
nor U2115 (N_2115,In_428,In_1228);
nand U2116 (N_2116,In_316,In_1022);
xor U2117 (N_2117,In_729,In_183);
nor U2118 (N_2118,In_477,In_696);
nand U2119 (N_2119,In_1762,In_1842);
xor U2120 (N_2120,In_560,In_77);
nor U2121 (N_2121,In_460,In_23);
or U2122 (N_2122,In_1743,In_496);
and U2123 (N_2123,In_1009,In_252);
and U2124 (N_2124,In_1317,In_214);
xnor U2125 (N_2125,In_1177,In_1453);
nor U2126 (N_2126,In_1068,In_736);
nor U2127 (N_2127,In_1234,In_116);
and U2128 (N_2128,In_212,In_578);
or U2129 (N_2129,In_468,In_1356);
xnor U2130 (N_2130,In_1046,In_1769);
xnor U2131 (N_2131,In_575,In_1852);
or U2132 (N_2132,In_1518,In_1393);
and U2133 (N_2133,In_1502,In_454);
and U2134 (N_2134,In_221,In_1410);
and U2135 (N_2135,In_452,In_851);
nand U2136 (N_2136,In_1719,In_1421);
nor U2137 (N_2137,In_167,In_754);
and U2138 (N_2138,In_736,In_1232);
nor U2139 (N_2139,In_581,In_221);
nor U2140 (N_2140,In_114,In_1825);
nand U2141 (N_2141,In_1739,In_631);
and U2142 (N_2142,In_87,In_1210);
nor U2143 (N_2143,In_922,In_1717);
nor U2144 (N_2144,In_1518,In_1326);
xnor U2145 (N_2145,In_1601,In_1117);
or U2146 (N_2146,In_426,In_1022);
nand U2147 (N_2147,In_957,In_1483);
or U2148 (N_2148,In_797,In_118);
or U2149 (N_2149,In_1997,In_593);
nand U2150 (N_2150,In_1512,In_438);
or U2151 (N_2151,In_529,In_394);
nor U2152 (N_2152,In_1291,In_1218);
nand U2153 (N_2153,In_200,In_404);
or U2154 (N_2154,In_1434,In_1191);
nor U2155 (N_2155,In_661,In_1907);
nand U2156 (N_2156,In_1996,In_1659);
and U2157 (N_2157,In_433,In_1513);
nor U2158 (N_2158,In_1104,In_1395);
or U2159 (N_2159,In_795,In_433);
nand U2160 (N_2160,In_826,In_632);
or U2161 (N_2161,In_904,In_751);
nand U2162 (N_2162,In_124,In_1832);
or U2163 (N_2163,In_1171,In_1972);
nor U2164 (N_2164,In_84,In_1056);
or U2165 (N_2165,In_1719,In_1572);
xor U2166 (N_2166,In_683,In_126);
nand U2167 (N_2167,In_1862,In_1855);
nor U2168 (N_2168,In_1942,In_1691);
nand U2169 (N_2169,In_1880,In_49);
and U2170 (N_2170,In_999,In_1080);
or U2171 (N_2171,In_978,In_121);
and U2172 (N_2172,In_861,In_389);
xnor U2173 (N_2173,In_1915,In_239);
or U2174 (N_2174,In_1355,In_1024);
or U2175 (N_2175,In_26,In_1271);
and U2176 (N_2176,In_927,In_694);
nor U2177 (N_2177,In_927,In_1968);
or U2178 (N_2178,In_1593,In_134);
or U2179 (N_2179,In_1612,In_1610);
nor U2180 (N_2180,In_1280,In_1572);
or U2181 (N_2181,In_103,In_39);
nor U2182 (N_2182,In_1072,In_992);
nand U2183 (N_2183,In_1055,In_1837);
and U2184 (N_2184,In_1070,In_1719);
or U2185 (N_2185,In_113,In_1607);
nand U2186 (N_2186,In_1832,In_669);
nor U2187 (N_2187,In_1806,In_862);
nor U2188 (N_2188,In_1131,In_927);
nor U2189 (N_2189,In_1424,In_1861);
or U2190 (N_2190,In_900,In_1400);
and U2191 (N_2191,In_40,In_907);
and U2192 (N_2192,In_1663,In_1630);
nor U2193 (N_2193,In_421,In_677);
or U2194 (N_2194,In_792,In_653);
xor U2195 (N_2195,In_10,In_1552);
or U2196 (N_2196,In_909,In_1375);
nand U2197 (N_2197,In_1947,In_908);
and U2198 (N_2198,In_871,In_702);
nor U2199 (N_2199,In_323,In_642);
and U2200 (N_2200,In_529,In_1385);
nand U2201 (N_2201,In_1138,In_822);
xor U2202 (N_2202,In_302,In_1001);
nand U2203 (N_2203,In_207,In_1495);
and U2204 (N_2204,In_805,In_506);
or U2205 (N_2205,In_1132,In_668);
and U2206 (N_2206,In_290,In_1265);
nand U2207 (N_2207,In_1142,In_926);
nor U2208 (N_2208,In_1434,In_499);
xnor U2209 (N_2209,In_482,In_1354);
xnor U2210 (N_2210,In_868,In_148);
and U2211 (N_2211,In_1902,In_581);
nor U2212 (N_2212,In_470,In_1922);
and U2213 (N_2213,In_226,In_1874);
or U2214 (N_2214,In_1011,In_95);
xnor U2215 (N_2215,In_430,In_654);
nand U2216 (N_2216,In_569,In_947);
nor U2217 (N_2217,In_903,In_409);
nor U2218 (N_2218,In_82,In_492);
or U2219 (N_2219,In_7,In_682);
or U2220 (N_2220,In_328,In_1830);
xor U2221 (N_2221,In_1391,In_565);
or U2222 (N_2222,In_14,In_1906);
xor U2223 (N_2223,In_628,In_888);
nand U2224 (N_2224,In_1681,In_1440);
nor U2225 (N_2225,In_309,In_1467);
and U2226 (N_2226,In_912,In_1230);
nor U2227 (N_2227,In_1106,In_122);
nor U2228 (N_2228,In_1869,In_680);
xnor U2229 (N_2229,In_1415,In_1032);
and U2230 (N_2230,In_1435,In_1887);
xor U2231 (N_2231,In_57,In_240);
and U2232 (N_2232,In_59,In_180);
xnor U2233 (N_2233,In_1705,In_1520);
nor U2234 (N_2234,In_1089,In_1977);
and U2235 (N_2235,In_1587,In_300);
or U2236 (N_2236,In_1602,In_229);
or U2237 (N_2237,In_1401,In_1596);
or U2238 (N_2238,In_1287,In_1936);
and U2239 (N_2239,In_1619,In_261);
nand U2240 (N_2240,In_634,In_351);
and U2241 (N_2241,In_1391,In_640);
xnor U2242 (N_2242,In_958,In_1617);
nand U2243 (N_2243,In_1043,In_1631);
or U2244 (N_2244,In_1445,In_1209);
and U2245 (N_2245,In_1127,In_1185);
nand U2246 (N_2246,In_912,In_834);
and U2247 (N_2247,In_744,In_580);
nor U2248 (N_2248,In_692,In_10);
and U2249 (N_2249,In_28,In_1300);
xnor U2250 (N_2250,In_1371,In_140);
or U2251 (N_2251,In_540,In_107);
or U2252 (N_2252,In_500,In_1024);
nor U2253 (N_2253,In_1556,In_1415);
nor U2254 (N_2254,In_1079,In_28);
and U2255 (N_2255,In_1575,In_1861);
or U2256 (N_2256,In_1188,In_1306);
and U2257 (N_2257,In_219,In_131);
nand U2258 (N_2258,In_1304,In_1913);
nand U2259 (N_2259,In_508,In_1996);
xor U2260 (N_2260,In_1333,In_370);
and U2261 (N_2261,In_1298,In_1142);
nor U2262 (N_2262,In_1520,In_1296);
nor U2263 (N_2263,In_1255,In_1337);
xor U2264 (N_2264,In_684,In_1357);
nand U2265 (N_2265,In_1,In_1546);
nand U2266 (N_2266,In_63,In_363);
nor U2267 (N_2267,In_1825,In_1330);
and U2268 (N_2268,In_1061,In_1250);
xor U2269 (N_2269,In_431,In_809);
and U2270 (N_2270,In_174,In_1491);
nand U2271 (N_2271,In_840,In_1516);
nor U2272 (N_2272,In_1837,In_1077);
nand U2273 (N_2273,In_1144,In_1316);
nor U2274 (N_2274,In_1895,In_743);
nor U2275 (N_2275,In_999,In_1717);
xnor U2276 (N_2276,In_121,In_1788);
or U2277 (N_2277,In_393,In_1126);
nand U2278 (N_2278,In_40,In_696);
or U2279 (N_2279,In_915,In_1366);
and U2280 (N_2280,In_1431,In_1808);
or U2281 (N_2281,In_826,In_1818);
nor U2282 (N_2282,In_775,In_923);
nand U2283 (N_2283,In_1957,In_313);
or U2284 (N_2284,In_1840,In_1535);
or U2285 (N_2285,In_1836,In_1802);
xnor U2286 (N_2286,In_1298,In_1617);
or U2287 (N_2287,In_432,In_1619);
nand U2288 (N_2288,In_901,In_1456);
nor U2289 (N_2289,In_247,In_1611);
or U2290 (N_2290,In_348,In_1046);
xor U2291 (N_2291,In_886,In_1344);
or U2292 (N_2292,In_1850,In_1723);
nand U2293 (N_2293,In_201,In_560);
or U2294 (N_2294,In_1316,In_1897);
and U2295 (N_2295,In_330,In_1363);
and U2296 (N_2296,In_742,In_1826);
xnor U2297 (N_2297,In_70,In_1260);
xnor U2298 (N_2298,In_757,In_213);
nor U2299 (N_2299,In_1066,In_578);
nor U2300 (N_2300,In_1160,In_1732);
nor U2301 (N_2301,In_1483,In_1951);
xnor U2302 (N_2302,In_1693,In_611);
nand U2303 (N_2303,In_1408,In_635);
nand U2304 (N_2304,In_1218,In_1809);
or U2305 (N_2305,In_506,In_1077);
xnor U2306 (N_2306,In_1087,In_1218);
xnor U2307 (N_2307,In_538,In_1058);
or U2308 (N_2308,In_750,In_211);
nor U2309 (N_2309,In_264,In_1054);
or U2310 (N_2310,In_1695,In_806);
nand U2311 (N_2311,In_147,In_1461);
or U2312 (N_2312,In_653,In_1254);
xnor U2313 (N_2313,In_38,In_1879);
and U2314 (N_2314,In_1855,In_870);
xor U2315 (N_2315,In_1337,In_1089);
and U2316 (N_2316,In_312,In_409);
nor U2317 (N_2317,In_663,In_268);
nor U2318 (N_2318,In_1728,In_1668);
and U2319 (N_2319,In_1939,In_372);
and U2320 (N_2320,In_385,In_1444);
xnor U2321 (N_2321,In_778,In_460);
or U2322 (N_2322,In_325,In_974);
and U2323 (N_2323,In_180,In_627);
xor U2324 (N_2324,In_37,In_979);
or U2325 (N_2325,In_725,In_573);
nand U2326 (N_2326,In_585,In_1071);
nand U2327 (N_2327,In_918,In_1182);
xor U2328 (N_2328,In_351,In_1074);
or U2329 (N_2329,In_1308,In_1234);
xor U2330 (N_2330,In_1272,In_1600);
nand U2331 (N_2331,In_1716,In_1161);
xor U2332 (N_2332,In_1547,In_1354);
xor U2333 (N_2333,In_841,In_1470);
nand U2334 (N_2334,In_1953,In_781);
nand U2335 (N_2335,In_222,In_1634);
nor U2336 (N_2336,In_1125,In_1185);
xnor U2337 (N_2337,In_741,In_1974);
or U2338 (N_2338,In_1167,In_248);
xnor U2339 (N_2339,In_696,In_915);
or U2340 (N_2340,In_1893,In_1336);
nor U2341 (N_2341,In_334,In_623);
nor U2342 (N_2342,In_307,In_1643);
xor U2343 (N_2343,In_241,In_926);
nand U2344 (N_2344,In_960,In_1213);
and U2345 (N_2345,In_1267,In_1622);
xnor U2346 (N_2346,In_738,In_1651);
and U2347 (N_2347,In_1975,In_752);
xor U2348 (N_2348,In_497,In_1660);
and U2349 (N_2349,In_1726,In_1431);
or U2350 (N_2350,In_1819,In_744);
xor U2351 (N_2351,In_1520,In_485);
nand U2352 (N_2352,In_564,In_308);
nand U2353 (N_2353,In_1422,In_1046);
and U2354 (N_2354,In_764,In_1191);
and U2355 (N_2355,In_281,In_315);
nor U2356 (N_2356,In_1804,In_1607);
nor U2357 (N_2357,In_1085,In_743);
or U2358 (N_2358,In_704,In_1133);
nor U2359 (N_2359,In_1634,In_158);
and U2360 (N_2360,In_1958,In_1720);
nor U2361 (N_2361,In_737,In_958);
nor U2362 (N_2362,In_925,In_1040);
nor U2363 (N_2363,In_1116,In_321);
nor U2364 (N_2364,In_1006,In_1019);
nor U2365 (N_2365,In_236,In_812);
nor U2366 (N_2366,In_600,In_909);
or U2367 (N_2367,In_1486,In_1487);
and U2368 (N_2368,In_1461,In_1659);
nor U2369 (N_2369,In_102,In_368);
nor U2370 (N_2370,In_1516,In_239);
or U2371 (N_2371,In_1586,In_1364);
or U2372 (N_2372,In_803,In_542);
nand U2373 (N_2373,In_1460,In_909);
and U2374 (N_2374,In_1009,In_1894);
nor U2375 (N_2375,In_1444,In_495);
or U2376 (N_2376,In_1928,In_1918);
or U2377 (N_2377,In_1743,In_623);
and U2378 (N_2378,In_1381,In_117);
and U2379 (N_2379,In_1111,In_1952);
and U2380 (N_2380,In_1668,In_1435);
xnor U2381 (N_2381,In_1731,In_1464);
xor U2382 (N_2382,In_1976,In_1219);
nor U2383 (N_2383,In_1193,In_1461);
nand U2384 (N_2384,In_1648,In_1046);
or U2385 (N_2385,In_93,In_247);
and U2386 (N_2386,In_1156,In_180);
xor U2387 (N_2387,In_1188,In_910);
nand U2388 (N_2388,In_755,In_1349);
nand U2389 (N_2389,In_1483,In_258);
nand U2390 (N_2390,In_533,In_806);
nor U2391 (N_2391,In_1019,In_225);
nand U2392 (N_2392,In_672,In_1671);
or U2393 (N_2393,In_1618,In_320);
and U2394 (N_2394,In_1067,In_796);
nor U2395 (N_2395,In_125,In_1167);
xor U2396 (N_2396,In_1604,In_568);
nor U2397 (N_2397,In_1110,In_939);
xnor U2398 (N_2398,In_1643,In_962);
or U2399 (N_2399,In_1287,In_725);
nand U2400 (N_2400,In_1181,In_181);
or U2401 (N_2401,In_0,In_1559);
and U2402 (N_2402,In_991,In_1250);
nand U2403 (N_2403,In_1627,In_57);
and U2404 (N_2404,In_22,In_231);
xnor U2405 (N_2405,In_10,In_1284);
and U2406 (N_2406,In_905,In_1630);
nor U2407 (N_2407,In_457,In_1097);
nand U2408 (N_2408,In_1983,In_1146);
nor U2409 (N_2409,In_1455,In_839);
and U2410 (N_2410,In_1300,In_478);
or U2411 (N_2411,In_82,In_1719);
xnor U2412 (N_2412,In_1269,In_683);
and U2413 (N_2413,In_84,In_1450);
or U2414 (N_2414,In_1966,In_1964);
nor U2415 (N_2415,In_800,In_355);
nor U2416 (N_2416,In_1545,In_530);
nor U2417 (N_2417,In_448,In_1400);
nor U2418 (N_2418,In_1719,In_1171);
nor U2419 (N_2419,In_856,In_1975);
or U2420 (N_2420,In_1972,In_1399);
or U2421 (N_2421,In_1061,In_1108);
and U2422 (N_2422,In_1908,In_934);
nor U2423 (N_2423,In_1382,In_1150);
or U2424 (N_2424,In_757,In_868);
and U2425 (N_2425,In_405,In_1847);
nor U2426 (N_2426,In_177,In_976);
nor U2427 (N_2427,In_261,In_1960);
xnor U2428 (N_2428,In_1132,In_569);
nor U2429 (N_2429,In_574,In_1245);
and U2430 (N_2430,In_305,In_442);
xnor U2431 (N_2431,In_1091,In_96);
nand U2432 (N_2432,In_747,In_1409);
xnor U2433 (N_2433,In_1998,In_1152);
or U2434 (N_2434,In_1999,In_1745);
or U2435 (N_2435,In_1967,In_1173);
xnor U2436 (N_2436,In_268,In_440);
and U2437 (N_2437,In_175,In_1466);
nand U2438 (N_2438,In_104,In_1598);
nand U2439 (N_2439,In_1048,In_270);
or U2440 (N_2440,In_1721,In_349);
xor U2441 (N_2441,In_1732,In_1977);
or U2442 (N_2442,In_237,In_991);
and U2443 (N_2443,In_658,In_1131);
nor U2444 (N_2444,In_1495,In_637);
and U2445 (N_2445,In_831,In_1762);
nor U2446 (N_2446,In_1265,In_1019);
nor U2447 (N_2447,In_890,In_823);
xor U2448 (N_2448,In_1175,In_1509);
xor U2449 (N_2449,In_331,In_1854);
or U2450 (N_2450,In_1245,In_818);
xnor U2451 (N_2451,In_904,In_486);
nor U2452 (N_2452,In_725,In_1224);
nor U2453 (N_2453,In_1005,In_1301);
and U2454 (N_2454,In_243,In_595);
or U2455 (N_2455,In_1053,In_558);
xor U2456 (N_2456,In_506,In_636);
or U2457 (N_2457,In_84,In_1179);
and U2458 (N_2458,In_255,In_679);
or U2459 (N_2459,In_1044,In_1277);
nand U2460 (N_2460,In_1543,In_1796);
and U2461 (N_2461,In_1266,In_1381);
nand U2462 (N_2462,In_898,In_549);
and U2463 (N_2463,In_1020,In_0);
xnor U2464 (N_2464,In_1586,In_1600);
xor U2465 (N_2465,In_901,In_929);
or U2466 (N_2466,In_530,In_545);
nor U2467 (N_2467,In_302,In_1959);
nand U2468 (N_2468,In_706,In_1660);
nand U2469 (N_2469,In_1757,In_664);
and U2470 (N_2470,In_89,In_1094);
nand U2471 (N_2471,In_946,In_1897);
and U2472 (N_2472,In_271,In_25);
xor U2473 (N_2473,In_1325,In_926);
and U2474 (N_2474,In_578,In_1982);
and U2475 (N_2475,In_1462,In_208);
nor U2476 (N_2476,In_1222,In_1241);
xnor U2477 (N_2477,In_1649,In_1268);
or U2478 (N_2478,In_1921,In_1337);
or U2479 (N_2479,In_440,In_869);
and U2480 (N_2480,In_1415,In_1740);
nand U2481 (N_2481,In_824,In_710);
and U2482 (N_2482,In_571,In_1277);
xnor U2483 (N_2483,In_1879,In_958);
or U2484 (N_2484,In_1074,In_344);
xor U2485 (N_2485,In_1087,In_900);
or U2486 (N_2486,In_512,In_1100);
or U2487 (N_2487,In_845,In_331);
nand U2488 (N_2488,In_834,In_606);
nand U2489 (N_2489,In_436,In_1642);
or U2490 (N_2490,In_328,In_1403);
or U2491 (N_2491,In_1982,In_862);
nor U2492 (N_2492,In_1064,In_1847);
nor U2493 (N_2493,In_1187,In_831);
or U2494 (N_2494,In_598,In_554);
xnor U2495 (N_2495,In_1888,In_522);
nand U2496 (N_2496,In_781,In_154);
and U2497 (N_2497,In_1864,In_890);
nand U2498 (N_2498,In_743,In_1898);
nor U2499 (N_2499,In_1147,In_1313);
and U2500 (N_2500,In_9,In_1188);
nand U2501 (N_2501,In_1001,In_1512);
nor U2502 (N_2502,In_1465,In_1082);
and U2503 (N_2503,In_1621,In_1175);
nand U2504 (N_2504,In_404,In_1285);
nor U2505 (N_2505,In_1003,In_1214);
and U2506 (N_2506,In_231,In_1579);
nand U2507 (N_2507,In_228,In_471);
and U2508 (N_2508,In_128,In_345);
xor U2509 (N_2509,In_1794,In_107);
or U2510 (N_2510,In_1671,In_759);
and U2511 (N_2511,In_1728,In_1536);
or U2512 (N_2512,In_752,In_1832);
xor U2513 (N_2513,In_1091,In_460);
xor U2514 (N_2514,In_1179,In_326);
or U2515 (N_2515,In_1279,In_956);
nand U2516 (N_2516,In_681,In_1233);
or U2517 (N_2517,In_1175,In_648);
nor U2518 (N_2518,In_1311,In_1503);
xor U2519 (N_2519,In_965,In_1079);
xor U2520 (N_2520,In_1420,In_1759);
and U2521 (N_2521,In_636,In_1215);
nand U2522 (N_2522,In_430,In_730);
xnor U2523 (N_2523,In_1772,In_179);
nand U2524 (N_2524,In_270,In_904);
xor U2525 (N_2525,In_1342,In_1828);
nand U2526 (N_2526,In_1311,In_1670);
xor U2527 (N_2527,In_1559,In_1938);
nand U2528 (N_2528,In_518,In_1360);
nor U2529 (N_2529,In_945,In_895);
nor U2530 (N_2530,In_1148,In_1272);
or U2531 (N_2531,In_62,In_363);
nor U2532 (N_2532,In_702,In_1804);
nand U2533 (N_2533,In_181,In_1427);
and U2534 (N_2534,In_1068,In_651);
or U2535 (N_2535,In_431,In_1719);
nand U2536 (N_2536,In_604,In_90);
and U2537 (N_2537,In_938,In_218);
and U2538 (N_2538,In_1299,In_1370);
and U2539 (N_2539,In_153,In_366);
or U2540 (N_2540,In_280,In_458);
nor U2541 (N_2541,In_1953,In_300);
and U2542 (N_2542,In_1699,In_331);
xor U2543 (N_2543,In_176,In_191);
or U2544 (N_2544,In_1214,In_1795);
nand U2545 (N_2545,In_1461,In_945);
and U2546 (N_2546,In_854,In_136);
nor U2547 (N_2547,In_23,In_1375);
nand U2548 (N_2548,In_1051,In_294);
or U2549 (N_2549,In_455,In_1930);
or U2550 (N_2550,In_1393,In_1398);
or U2551 (N_2551,In_1725,In_146);
and U2552 (N_2552,In_516,In_1034);
xor U2553 (N_2553,In_914,In_798);
and U2554 (N_2554,In_1076,In_953);
nand U2555 (N_2555,In_1218,In_104);
xnor U2556 (N_2556,In_104,In_1401);
or U2557 (N_2557,In_1472,In_1684);
nand U2558 (N_2558,In_453,In_82);
or U2559 (N_2559,In_1064,In_1494);
nor U2560 (N_2560,In_1875,In_430);
and U2561 (N_2561,In_342,In_129);
nor U2562 (N_2562,In_1466,In_762);
nand U2563 (N_2563,In_689,In_664);
xor U2564 (N_2564,In_1467,In_484);
nor U2565 (N_2565,In_892,In_1260);
xnor U2566 (N_2566,In_245,In_1787);
or U2567 (N_2567,In_556,In_659);
and U2568 (N_2568,In_1688,In_685);
and U2569 (N_2569,In_1788,In_1133);
or U2570 (N_2570,In_855,In_1411);
nor U2571 (N_2571,In_1452,In_404);
xor U2572 (N_2572,In_89,In_1980);
or U2573 (N_2573,In_601,In_1574);
and U2574 (N_2574,In_1178,In_532);
or U2575 (N_2575,In_817,In_192);
and U2576 (N_2576,In_495,In_1228);
xnor U2577 (N_2577,In_289,In_1361);
and U2578 (N_2578,In_896,In_1370);
and U2579 (N_2579,In_1598,In_363);
and U2580 (N_2580,In_1664,In_1169);
or U2581 (N_2581,In_1809,In_1555);
nor U2582 (N_2582,In_1728,In_1836);
nand U2583 (N_2583,In_1721,In_934);
and U2584 (N_2584,In_1403,In_404);
nor U2585 (N_2585,In_1979,In_1470);
nor U2586 (N_2586,In_1343,In_818);
or U2587 (N_2587,In_1389,In_457);
nor U2588 (N_2588,In_1401,In_571);
nand U2589 (N_2589,In_944,In_561);
nor U2590 (N_2590,In_1761,In_1030);
and U2591 (N_2591,In_1491,In_1837);
or U2592 (N_2592,In_1943,In_923);
nand U2593 (N_2593,In_549,In_498);
or U2594 (N_2594,In_40,In_422);
and U2595 (N_2595,In_1806,In_1542);
nand U2596 (N_2596,In_738,In_1591);
nand U2597 (N_2597,In_1697,In_123);
nand U2598 (N_2598,In_400,In_1215);
or U2599 (N_2599,In_924,In_1173);
and U2600 (N_2600,In_1080,In_1821);
and U2601 (N_2601,In_879,In_968);
nand U2602 (N_2602,In_1355,In_1363);
nand U2603 (N_2603,In_287,In_1525);
and U2604 (N_2604,In_1073,In_1109);
xor U2605 (N_2605,In_672,In_431);
and U2606 (N_2606,In_928,In_46);
nand U2607 (N_2607,In_1703,In_1531);
and U2608 (N_2608,In_1168,In_639);
and U2609 (N_2609,In_1864,In_978);
and U2610 (N_2610,In_433,In_299);
xor U2611 (N_2611,In_703,In_1435);
nand U2612 (N_2612,In_80,In_1829);
or U2613 (N_2613,In_1717,In_1798);
and U2614 (N_2614,In_342,In_14);
nand U2615 (N_2615,In_1530,In_1010);
nand U2616 (N_2616,In_53,In_1440);
or U2617 (N_2617,In_1287,In_1491);
nor U2618 (N_2618,In_818,In_1102);
nor U2619 (N_2619,In_1125,In_1054);
or U2620 (N_2620,In_1634,In_1170);
and U2621 (N_2621,In_5,In_630);
xnor U2622 (N_2622,In_444,In_591);
nand U2623 (N_2623,In_1410,In_1965);
and U2624 (N_2624,In_1717,In_1555);
or U2625 (N_2625,In_685,In_1480);
nand U2626 (N_2626,In_452,In_1949);
xnor U2627 (N_2627,In_1903,In_1488);
or U2628 (N_2628,In_34,In_206);
and U2629 (N_2629,In_38,In_1678);
xor U2630 (N_2630,In_421,In_410);
xnor U2631 (N_2631,In_1149,In_5);
xnor U2632 (N_2632,In_1552,In_685);
xnor U2633 (N_2633,In_39,In_970);
nand U2634 (N_2634,In_1824,In_1477);
and U2635 (N_2635,In_1582,In_1758);
nand U2636 (N_2636,In_100,In_1302);
xnor U2637 (N_2637,In_322,In_1595);
nor U2638 (N_2638,In_1936,In_562);
nand U2639 (N_2639,In_1190,In_1563);
nand U2640 (N_2640,In_364,In_1576);
xnor U2641 (N_2641,In_1495,In_1096);
nand U2642 (N_2642,In_81,In_1796);
xnor U2643 (N_2643,In_421,In_1444);
nand U2644 (N_2644,In_1849,In_839);
and U2645 (N_2645,In_861,In_1259);
nand U2646 (N_2646,In_1190,In_286);
nand U2647 (N_2647,In_180,In_721);
nor U2648 (N_2648,In_446,In_1905);
xnor U2649 (N_2649,In_927,In_707);
nor U2650 (N_2650,In_1906,In_1641);
nand U2651 (N_2651,In_1021,In_1404);
xor U2652 (N_2652,In_209,In_951);
nand U2653 (N_2653,In_320,In_1440);
and U2654 (N_2654,In_360,In_882);
nor U2655 (N_2655,In_333,In_126);
nand U2656 (N_2656,In_1512,In_300);
nand U2657 (N_2657,In_870,In_745);
or U2658 (N_2658,In_145,In_1960);
xnor U2659 (N_2659,In_822,In_922);
and U2660 (N_2660,In_1562,In_1403);
nor U2661 (N_2661,In_1638,In_1371);
nor U2662 (N_2662,In_1733,In_1046);
and U2663 (N_2663,In_1462,In_425);
xor U2664 (N_2664,In_421,In_252);
nand U2665 (N_2665,In_911,In_1703);
or U2666 (N_2666,In_806,In_1176);
nor U2667 (N_2667,In_742,In_183);
or U2668 (N_2668,In_200,In_345);
xnor U2669 (N_2669,In_1372,In_1551);
nor U2670 (N_2670,In_898,In_1179);
and U2671 (N_2671,In_1262,In_1841);
xnor U2672 (N_2672,In_332,In_1516);
nor U2673 (N_2673,In_1491,In_1217);
nor U2674 (N_2674,In_402,In_1297);
xnor U2675 (N_2675,In_1946,In_1750);
nand U2676 (N_2676,In_105,In_1823);
or U2677 (N_2677,In_1333,In_1943);
nor U2678 (N_2678,In_1163,In_258);
xor U2679 (N_2679,In_488,In_1566);
xnor U2680 (N_2680,In_445,In_1858);
and U2681 (N_2681,In_1168,In_184);
nand U2682 (N_2682,In_439,In_1275);
and U2683 (N_2683,In_932,In_968);
nor U2684 (N_2684,In_1763,In_1421);
or U2685 (N_2685,In_1166,In_667);
xor U2686 (N_2686,In_1546,In_1255);
and U2687 (N_2687,In_803,In_1976);
xor U2688 (N_2688,In_1176,In_1424);
or U2689 (N_2689,In_1326,In_385);
xnor U2690 (N_2690,In_1066,In_399);
nand U2691 (N_2691,In_727,In_1370);
and U2692 (N_2692,In_1414,In_1589);
nor U2693 (N_2693,In_1376,In_839);
and U2694 (N_2694,In_188,In_372);
nor U2695 (N_2695,In_510,In_1676);
xor U2696 (N_2696,In_1730,In_415);
nand U2697 (N_2697,In_1186,In_1074);
and U2698 (N_2698,In_1347,In_878);
xor U2699 (N_2699,In_1675,In_102);
or U2700 (N_2700,In_545,In_1587);
or U2701 (N_2701,In_143,In_871);
or U2702 (N_2702,In_1948,In_647);
nand U2703 (N_2703,In_1787,In_105);
nand U2704 (N_2704,In_1763,In_1547);
xor U2705 (N_2705,In_280,In_1724);
nor U2706 (N_2706,In_1831,In_1073);
or U2707 (N_2707,In_797,In_1431);
xnor U2708 (N_2708,In_226,In_994);
xnor U2709 (N_2709,In_635,In_1077);
nand U2710 (N_2710,In_1525,In_804);
or U2711 (N_2711,In_562,In_271);
nor U2712 (N_2712,In_1317,In_1687);
or U2713 (N_2713,In_1094,In_371);
or U2714 (N_2714,In_1559,In_1502);
nand U2715 (N_2715,In_1889,In_1987);
xnor U2716 (N_2716,In_1891,In_1894);
nand U2717 (N_2717,In_796,In_1908);
xnor U2718 (N_2718,In_203,In_97);
and U2719 (N_2719,In_437,In_690);
nand U2720 (N_2720,In_27,In_972);
nand U2721 (N_2721,In_302,In_59);
nand U2722 (N_2722,In_39,In_1431);
nor U2723 (N_2723,In_1092,In_1326);
xnor U2724 (N_2724,In_977,In_518);
nor U2725 (N_2725,In_617,In_1712);
nor U2726 (N_2726,In_1495,In_724);
or U2727 (N_2727,In_1021,In_134);
and U2728 (N_2728,In_1830,In_1839);
and U2729 (N_2729,In_941,In_1358);
or U2730 (N_2730,In_260,In_1032);
nor U2731 (N_2731,In_1038,In_898);
nor U2732 (N_2732,In_40,In_1852);
nor U2733 (N_2733,In_1592,In_1388);
nand U2734 (N_2734,In_109,In_1351);
and U2735 (N_2735,In_1653,In_100);
nand U2736 (N_2736,In_1383,In_1384);
xnor U2737 (N_2737,In_1004,In_418);
and U2738 (N_2738,In_331,In_865);
and U2739 (N_2739,In_869,In_1357);
nand U2740 (N_2740,In_357,In_433);
nor U2741 (N_2741,In_1726,In_1915);
or U2742 (N_2742,In_851,In_435);
nand U2743 (N_2743,In_1542,In_1679);
and U2744 (N_2744,In_74,In_1859);
nor U2745 (N_2745,In_980,In_1879);
nand U2746 (N_2746,In_1488,In_587);
and U2747 (N_2747,In_217,In_938);
or U2748 (N_2748,In_1158,In_1681);
nor U2749 (N_2749,In_81,In_1021);
nor U2750 (N_2750,In_1648,In_1177);
nor U2751 (N_2751,In_1165,In_612);
nor U2752 (N_2752,In_1940,In_1163);
xor U2753 (N_2753,In_1970,In_859);
nor U2754 (N_2754,In_8,In_1138);
or U2755 (N_2755,In_1694,In_1445);
and U2756 (N_2756,In_1358,In_779);
and U2757 (N_2757,In_141,In_493);
nand U2758 (N_2758,In_659,In_1602);
nor U2759 (N_2759,In_333,In_129);
or U2760 (N_2760,In_516,In_686);
and U2761 (N_2761,In_1750,In_1932);
xnor U2762 (N_2762,In_957,In_1838);
nand U2763 (N_2763,In_486,In_948);
nor U2764 (N_2764,In_1698,In_1914);
xor U2765 (N_2765,In_1856,In_358);
and U2766 (N_2766,In_1445,In_125);
and U2767 (N_2767,In_1907,In_1382);
nor U2768 (N_2768,In_627,In_388);
xor U2769 (N_2769,In_810,In_708);
nor U2770 (N_2770,In_1556,In_525);
and U2771 (N_2771,In_950,In_129);
nor U2772 (N_2772,In_1038,In_277);
or U2773 (N_2773,In_373,In_1337);
nor U2774 (N_2774,In_1078,In_1417);
xnor U2775 (N_2775,In_1393,In_381);
or U2776 (N_2776,In_1170,In_1779);
xor U2777 (N_2777,In_491,In_1522);
or U2778 (N_2778,In_1587,In_995);
xnor U2779 (N_2779,In_335,In_404);
and U2780 (N_2780,In_1730,In_1361);
nor U2781 (N_2781,In_1205,In_311);
xor U2782 (N_2782,In_558,In_170);
nand U2783 (N_2783,In_1054,In_547);
or U2784 (N_2784,In_1048,In_1813);
nand U2785 (N_2785,In_1845,In_875);
nand U2786 (N_2786,In_1222,In_852);
nand U2787 (N_2787,In_174,In_1443);
xnor U2788 (N_2788,In_1491,In_1480);
nor U2789 (N_2789,In_1637,In_590);
or U2790 (N_2790,In_286,In_1027);
or U2791 (N_2791,In_639,In_375);
nor U2792 (N_2792,In_1873,In_230);
and U2793 (N_2793,In_1007,In_212);
or U2794 (N_2794,In_1613,In_513);
xnor U2795 (N_2795,In_102,In_1026);
nor U2796 (N_2796,In_660,In_1166);
nor U2797 (N_2797,In_1892,In_281);
and U2798 (N_2798,In_990,In_899);
nand U2799 (N_2799,In_1361,In_402);
xor U2800 (N_2800,In_1298,In_1732);
nor U2801 (N_2801,In_650,In_903);
nand U2802 (N_2802,In_909,In_761);
nor U2803 (N_2803,In_718,In_482);
xnor U2804 (N_2804,In_223,In_615);
or U2805 (N_2805,In_1253,In_522);
and U2806 (N_2806,In_364,In_1113);
xor U2807 (N_2807,In_1167,In_1359);
and U2808 (N_2808,In_890,In_1565);
nand U2809 (N_2809,In_928,In_578);
xnor U2810 (N_2810,In_301,In_1546);
nor U2811 (N_2811,In_225,In_1512);
or U2812 (N_2812,In_439,In_695);
nand U2813 (N_2813,In_1524,In_1635);
or U2814 (N_2814,In_1809,In_1848);
and U2815 (N_2815,In_1034,In_1039);
and U2816 (N_2816,In_637,In_987);
or U2817 (N_2817,In_1890,In_56);
nand U2818 (N_2818,In_1368,In_431);
or U2819 (N_2819,In_230,In_458);
nand U2820 (N_2820,In_1555,In_764);
or U2821 (N_2821,In_199,In_253);
xor U2822 (N_2822,In_1705,In_354);
nand U2823 (N_2823,In_1204,In_1199);
or U2824 (N_2824,In_1578,In_222);
nor U2825 (N_2825,In_1346,In_850);
or U2826 (N_2826,In_745,In_1267);
nand U2827 (N_2827,In_842,In_1617);
nor U2828 (N_2828,In_1889,In_760);
and U2829 (N_2829,In_484,In_133);
nor U2830 (N_2830,In_1955,In_999);
and U2831 (N_2831,In_821,In_180);
nand U2832 (N_2832,In_1070,In_1037);
or U2833 (N_2833,In_1283,In_909);
nor U2834 (N_2834,In_822,In_497);
and U2835 (N_2835,In_1947,In_1370);
nor U2836 (N_2836,In_155,In_13);
or U2837 (N_2837,In_1512,In_7);
and U2838 (N_2838,In_863,In_981);
nand U2839 (N_2839,In_258,In_640);
nor U2840 (N_2840,In_1398,In_1843);
or U2841 (N_2841,In_1004,In_1855);
and U2842 (N_2842,In_1257,In_1012);
and U2843 (N_2843,In_1056,In_1852);
nand U2844 (N_2844,In_1650,In_285);
nand U2845 (N_2845,In_575,In_497);
and U2846 (N_2846,In_1879,In_1366);
and U2847 (N_2847,In_1947,In_1857);
xnor U2848 (N_2848,In_321,In_1570);
or U2849 (N_2849,In_1136,In_1794);
nor U2850 (N_2850,In_916,In_1808);
and U2851 (N_2851,In_1456,In_170);
or U2852 (N_2852,In_372,In_1366);
and U2853 (N_2853,In_277,In_151);
xnor U2854 (N_2854,In_538,In_1478);
xnor U2855 (N_2855,In_1556,In_633);
and U2856 (N_2856,In_360,In_685);
or U2857 (N_2857,In_552,In_1708);
nand U2858 (N_2858,In_1846,In_279);
and U2859 (N_2859,In_1682,In_1666);
xnor U2860 (N_2860,In_500,In_1160);
nand U2861 (N_2861,In_338,In_1338);
or U2862 (N_2862,In_1757,In_1429);
nor U2863 (N_2863,In_1350,In_579);
and U2864 (N_2864,In_796,In_116);
and U2865 (N_2865,In_356,In_1893);
or U2866 (N_2866,In_329,In_32);
and U2867 (N_2867,In_210,In_1679);
nor U2868 (N_2868,In_921,In_258);
xor U2869 (N_2869,In_1860,In_1532);
nand U2870 (N_2870,In_950,In_520);
nor U2871 (N_2871,In_311,In_1899);
and U2872 (N_2872,In_1526,In_1031);
xnor U2873 (N_2873,In_181,In_1274);
and U2874 (N_2874,In_1361,In_886);
and U2875 (N_2875,In_685,In_1244);
or U2876 (N_2876,In_194,In_1128);
nand U2877 (N_2877,In_1643,In_687);
nor U2878 (N_2878,In_893,In_1253);
or U2879 (N_2879,In_1522,In_39);
nand U2880 (N_2880,In_33,In_609);
and U2881 (N_2881,In_168,In_1063);
and U2882 (N_2882,In_1851,In_760);
nand U2883 (N_2883,In_1189,In_1762);
or U2884 (N_2884,In_1091,In_591);
nor U2885 (N_2885,In_610,In_969);
nor U2886 (N_2886,In_37,In_1600);
and U2887 (N_2887,In_1818,In_1708);
and U2888 (N_2888,In_1783,In_834);
xnor U2889 (N_2889,In_190,In_9);
nor U2890 (N_2890,In_1114,In_711);
xor U2891 (N_2891,In_1392,In_1648);
nand U2892 (N_2892,In_1355,In_1713);
nor U2893 (N_2893,In_744,In_343);
nor U2894 (N_2894,In_696,In_215);
or U2895 (N_2895,In_581,In_1339);
and U2896 (N_2896,In_767,In_360);
nand U2897 (N_2897,In_1602,In_733);
nand U2898 (N_2898,In_1662,In_596);
nor U2899 (N_2899,In_598,In_167);
nor U2900 (N_2900,In_1984,In_1517);
xor U2901 (N_2901,In_1341,In_987);
and U2902 (N_2902,In_1422,In_441);
and U2903 (N_2903,In_1166,In_577);
nor U2904 (N_2904,In_1552,In_851);
nand U2905 (N_2905,In_1666,In_990);
and U2906 (N_2906,In_411,In_590);
nand U2907 (N_2907,In_786,In_589);
nor U2908 (N_2908,In_1415,In_793);
nand U2909 (N_2909,In_251,In_1924);
and U2910 (N_2910,In_1285,In_603);
xnor U2911 (N_2911,In_285,In_742);
xnor U2912 (N_2912,In_1766,In_15);
and U2913 (N_2913,In_1527,In_384);
nand U2914 (N_2914,In_756,In_1871);
nor U2915 (N_2915,In_427,In_620);
and U2916 (N_2916,In_856,In_1240);
nor U2917 (N_2917,In_878,In_1141);
and U2918 (N_2918,In_710,In_1921);
xor U2919 (N_2919,In_1854,In_1711);
or U2920 (N_2920,In_1205,In_509);
nor U2921 (N_2921,In_1200,In_822);
nor U2922 (N_2922,In_1985,In_1641);
or U2923 (N_2923,In_1837,In_926);
xor U2924 (N_2924,In_1761,In_1837);
or U2925 (N_2925,In_973,In_557);
and U2926 (N_2926,In_356,In_628);
nand U2927 (N_2927,In_1273,In_1187);
nor U2928 (N_2928,In_806,In_837);
nand U2929 (N_2929,In_767,In_780);
xor U2930 (N_2930,In_1427,In_1761);
xor U2931 (N_2931,In_1884,In_1692);
or U2932 (N_2932,In_1978,In_1873);
and U2933 (N_2933,In_1938,In_612);
and U2934 (N_2934,In_845,In_1771);
xor U2935 (N_2935,In_642,In_122);
nand U2936 (N_2936,In_1052,In_32);
nor U2937 (N_2937,In_1485,In_1700);
nand U2938 (N_2938,In_936,In_157);
nor U2939 (N_2939,In_781,In_353);
nand U2940 (N_2940,In_1704,In_517);
nand U2941 (N_2941,In_1824,In_1735);
nand U2942 (N_2942,In_939,In_1565);
and U2943 (N_2943,In_1699,In_1231);
xnor U2944 (N_2944,In_336,In_627);
xnor U2945 (N_2945,In_112,In_1342);
nand U2946 (N_2946,In_1230,In_1048);
or U2947 (N_2947,In_1321,In_632);
nand U2948 (N_2948,In_223,In_1904);
xnor U2949 (N_2949,In_565,In_1652);
or U2950 (N_2950,In_415,In_816);
and U2951 (N_2951,In_1168,In_1946);
nor U2952 (N_2952,In_1315,In_1002);
and U2953 (N_2953,In_1243,In_1580);
and U2954 (N_2954,In_1195,In_1061);
and U2955 (N_2955,In_1551,In_1801);
or U2956 (N_2956,In_656,In_1439);
xnor U2957 (N_2957,In_883,In_983);
and U2958 (N_2958,In_1600,In_560);
xor U2959 (N_2959,In_1462,In_1401);
nand U2960 (N_2960,In_545,In_1030);
nor U2961 (N_2961,In_1652,In_259);
or U2962 (N_2962,In_1614,In_1175);
xor U2963 (N_2963,In_95,In_987);
and U2964 (N_2964,In_1179,In_1102);
and U2965 (N_2965,In_792,In_1451);
nand U2966 (N_2966,In_1358,In_1585);
nor U2967 (N_2967,In_1079,In_1194);
or U2968 (N_2968,In_250,In_1427);
or U2969 (N_2969,In_822,In_57);
or U2970 (N_2970,In_1766,In_1676);
or U2971 (N_2971,In_974,In_39);
nand U2972 (N_2972,In_1699,In_1674);
nand U2973 (N_2973,In_1746,In_1276);
xnor U2974 (N_2974,In_781,In_1212);
xnor U2975 (N_2975,In_868,In_144);
xnor U2976 (N_2976,In_1678,In_1942);
or U2977 (N_2977,In_1953,In_1567);
nand U2978 (N_2978,In_1306,In_1202);
or U2979 (N_2979,In_1572,In_1014);
nor U2980 (N_2980,In_1304,In_284);
xor U2981 (N_2981,In_48,In_1084);
nor U2982 (N_2982,In_837,In_681);
xnor U2983 (N_2983,In_690,In_343);
xor U2984 (N_2984,In_617,In_898);
nand U2985 (N_2985,In_386,In_867);
or U2986 (N_2986,In_1690,In_1027);
or U2987 (N_2987,In_181,In_463);
xnor U2988 (N_2988,In_1279,In_36);
xor U2989 (N_2989,In_699,In_1195);
or U2990 (N_2990,In_471,In_476);
nor U2991 (N_2991,In_1797,In_1182);
nor U2992 (N_2992,In_219,In_1567);
nand U2993 (N_2993,In_736,In_295);
nand U2994 (N_2994,In_11,In_1372);
and U2995 (N_2995,In_1178,In_31);
xnor U2996 (N_2996,In_1984,In_200);
nand U2997 (N_2997,In_955,In_255);
xnor U2998 (N_2998,In_1394,In_783);
nor U2999 (N_2999,In_467,In_1928);
nor U3000 (N_3000,In_292,In_1618);
xor U3001 (N_3001,In_1642,In_713);
and U3002 (N_3002,In_1681,In_1355);
or U3003 (N_3003,In_403,In_1739);
or U3004 (N_3004,In_333,In_973);
nand U3005 (N_3005,In_1962,In_1391);
nor U3006 (N_3006,In_799,In_1969);
nor U3007 (N_3007,In_1890,In_995);
nor U3008 (N_3008,In_93,In_501);
nor U3009 (N_3009,In_1651,In_89);
or U3010 (N_3010,In_1477,In_713);
nand U3011 (N_3011,In_1310,In_91);
nand U3012 (N_3012,In_1026,In_528);
or U3013 (N_3013,In_983,In_813);
nand U3014 (N_3014,In_833,In_1781);
nand U3015 (N_3015,In_1084,In_126);
nor U3016 (N_3016,In_1205,In_1384);
xnor U3017 (N_3017,In_1242,In_885);
and U3018 (N_3018,In_573,In_1295);
nand U3019 (N_3019,In_456,In_1555);
xnor U3020 (N_3020,In_1073,In_247);
and U3021 (N_3021,In_675,In_674);
or U3022 (N_3022,In_836,In_1635);
and U3023 (N_3023,In_212,In_234);
and U3024 (N_3024,In_64,In_1514);
or U3025 (N_3025,In_501,In_1571);
or U3026 (N_3026,In_44,In_1312);
nor U3027 (N_3027,In_548,In_1465);
or U3028 (N_3028,In_478,In_1419);
and U3029 (N_3029,In_1882,In_1336);
nor U3030 (N_3030,In_1139,In_1059);
nand U3031 (N_3031,In_160,In_326);
nand U3032 (N_3032,In_554,In_1337);
and U3033 (N_3033,In_237,In_1084);
or U3034 (N_3034,In_150,In_1951);
and U3035 (N_3035,In_733,In_121);
xor U3036 (N_3036,In_966,In_1803);
or U3037 (N_3037,In_266,In_1116);
xnor U3038 (N_3038,In_310,In_1268);
and U3039 (N_3039,In_1115,In_549);
xnor U3040 (N_3040,In_1343,In_1359);
nand U3041 (N_3041,In_1714,In_1887);
or U3042 (N_3042,In_840,In_1158);
and U3043 (N_3043,In_30,In_1655);
nand U3044 (N_3044,In_1403,In_990);
and U3045 (N_3045,In_1123,In_924);
or U3046 (N_3046,In_1539,In_640);
nand U3047 (N_3047,In_1915,In_1527);
and U3048 (N_3048,In_1907,In_789);
nand U3049 (N_3049,In_1979,In_1374);
and U3050 (N_3050,In_92,In_855);
xnor U3051 (N_3051,In_1276,In_925);
nand U3052 (N_3052,In_1630,In_1646);
and U3053 (N_3053,In_533,In_1128);
or U3054 (N_3054,In_1337,In_379);
or U3055 (N_3055,In_1471,In_1851);
nor U3056 (N_3056,In_1721,In_1824);
nor U3057 (N_3057,In_1518,In_1781);
xor U3058 (N_3058,In_604,In_685);
nor U3059 (N_3059,In_752,In_177);
and U3060 (N_3060,In_868,In_22);
xor U3061 (N_3061,In_1075,In_279);
nor U3062 (N_3062,In_307,In_724);
or U3063 (N_3063,In_1135,In_1277);
nand U3064 (N_3064,In_977,In_1648);
or U3065 (N_3065,In_1931,In_1029);
or U3066 (N_3066,In_384,In_774);
and U3067 (N_3067,In_631,In_1494);
or U3068 (N_3068,In_1107,In_767);
xor U3069 (N_3069,In_501,In_1029);
xor U3070 (N_3070,In_891,In_1891);
nor U3071 (N_3071,In_164,In_210);
xnor U3072 (N_3072,In_704,In_937);
nand U3073 (N_3073,In_1147,In_942);
nor U3074 (N_3074,In_128,In_9);
nor U3075 (N_3075,In_1297,In_1916);
nor U3076 (N_3076,In_1107,In_1886);
or U3077 (N_3077,In_538,In_95);
nor U3078 (N_3078,In_146,In_297);
nor U3079 (N_3079,In_1521,In_373);
nand U3080 (N_3080,In_1658,In_469);
and U3081 (N_3081,In_1142,In_975);
and U3082 (N_3082,In_350,In_1910);
nand U3083 (N_3083,In_908,In_609);
and U3084 (N_3084,In_705,In_172);
or U3085 (N_3085,In_1124,In_1953);
and U3086 (N_3086,In_333,In_1065);
nor U3087 (N_3087,In_1748,In_401);
xor U3088 (N_3088,In_9,In_1632);
xnor U3089 (N_3089,In_1914,In_739);
and U3090 (N_3090,In_1069,In_827);
or U3091 (N_3091,In_965,In_1042);
or U3092 (N_3092,In_1638,In_1270);
nor U3093 (N_3093,In_664,In_1954);
xor U3094 (N_3094,In_80,In_687);
xor U3095 (N_3095,In_1194,In_863);
xor U3096 (N_3096,In_1127,In_754);
or U3097 (N_3097,In_1879,In_405);
xnor U3098 (N_3098,In_855,In_744);
and U3099 (N_3099,In_351,In_1042);
and U3100 (N_3100,In_990,In_1524);
and U3101 (N_3101,In_1985,In_1353);
nor U3102 (N_3102,In_804,In_1772);
and U3103 (N_3103,In_1792,In_1624);
nand U3104 (N_3104,In_948,In_1768);
nand U3105 (N_3105,In_879,In_1295);
nor U3106 (N_3106,In_373,In_135);
xnor U3107 (N_3107,In_1994,In_1510);
and U3108 (N_3108,In_1732,In_308);
or U3109 (N_3109,In_1960,In_1697);
and U3110 (N_3110,In_1322,In_1042);
nand U3111 (N_3111,In_1109,In_494);
nand U3112 (N_3112,In_536,In_629);
xnor U3113 (N_3113,In_1645,In_1958);
nand U3114 (N_3114,In_1805,In_1235);
xor U3115 (N_3115,In_1572,In_54);
nand U3116 (N_3116,In_523,In_1000);
and U3117 (N_3117,In_1953,In_918);
or U3118 (N_3118,In_937,In_1963);
and U3119 (N_3119,In_1967,In_1943);
xor U3120 (N_3120,In_268,In_1748);
or U3121 (N_3121,In_509,In_1441);
or U3122 (N_3122,In_294,In_1715);
xor U3123 (N_3123,In_784,In_924);
nor U3124 (N_3124,In_1303,In_464);
and U3125 (N_3125,In_1109,In_1437);
and U3126 (N_3126,In_670,In_1106);
nand U3127 (N_3127,In_1813,In_133);
and U3128 (N_3128,In_1979,In_1251);
nor U3129 (N_3129,In_1913,In_191);
nand U3130 (N_3130,In_1560,In_736);
nor U3131 (N_3131,In_364,In_1226);
nor U3132 (N_3132,In_161,In_1361);
or U3133 (N_3133,In_245,In_1773);
or U3134 (N_3134,In_1616,In_1340);
nand U3135 (N_3135,In_681,In_910);
nand U3136 (N_3136,In_1659,In_1830);
and U3137 (N_3137,In_1838,In_1642);
xor U3138 (N_3138,In_1495,In_1398);
or U3139 (N_3139,In_368,In_678);
and U3140 (N_3140,In_744,In_1671);
and U3141 (N_3141,In_115,In_194);
or U3142 (N_3142,In_1600,In_270);
nor U3143 (N_3143,In_773,In_664);
and U3144 (N_3144,In_1332,In_1186);
xnor U3145 (N_3145,In_262,In_549);
and U3146 (N_3146,In_1441,In_853);
nand U3147 (N_3147,In_359,In_1995);
xnor U3148 (N_3148,In_1403,In_1261);
and U3149 (N_3149,In_376,In_261);
nand U3150 (N_3150,In_1328,In_1610);
nand U3151 (N_3151,In_53,In_400);
or U3152 (N_3152,In_1643,In_668);
and U3153 (N_3153,In_814,In_1632);
nand U3154 (N_3154,In_1344,In_1982);
and U3155 (N_3155,In_656,In_408);
or U3156 (N_3156,In_1697,In_1720);
xor U3157 (N_3157,In_923,In_584);
and U3158 (N_3158,In_3,In_1826);
and U3159 (N_3159,In_1115,In_643);
or U3160 (N_3160,In_1409,In_720);
xor U3161 (N_3161,In_1952,In_436);
xor U3162 (N_3162,In_1018,In_497);
or U3163 (N_3163,In_1588,In_1382);
or U3164 (N_3164,In_1921,In_700);
xor U3165 (N_3165,In_68,In_163);
xnor U3166 (N_3166,In_933,In_419);
nor U3167 (N_3167,In_71,In_37);
nor U3168 (N_3168,In_1391,In_1160);
nor U3169 (N_3169,In_1182,In_890);
and U3170 (N_3170,In_1839,In_754);
nor U3171 (N_3171,In_1256,In_108);
xor U3172 (N_3172,In_1081,In_38);
and U3173 (N_3173,In_1966,In_1494);
or U3174 (N_3174,In_1581,In_1945);
nand U3175 (N_3175,In_948,In_1258);
or U3176 (N_3176,In_665,In_1153);
and U3177 (N_3177,In_1007,In_1508);
and U3178 (N_3178,In_816,In_288);
and U3179 (N_3179,In_1362,In_264);
or U3180 (N_3180,In_1833,In_373);
or U3181 (N_3181,In_1116,In_1473);
nor U3182 (N_3182,In_1703,In_1972);
and U3183 (N_3183,In_664,In_1536);
xnor U3184 (N_3184,In_1803,In_369);
or U3185 (N_3185,In_134,In_472);
xnor U3186 (N_3186,In_1786,In_180);
and U3187 (N_3187,In_1229,In_1927);
nor U3188 (N_3188,In_850,In_316);
xnor U3189 (N_3189,In_261,In_271);
xnor U3190 (N_3190,In_827,In_373);
and U3191 (N_3191,In_1864,In_1420);
nand U3192 (N_3192,In_1990,In_1176);
nand U3193 (N_3193,In_1247,In_1276);
or U3194 (N_3194,In_1979,In_1689);
or U3195 (N_3195,In_165,In_34);
or U3196 (N_3196,In_514,In_441);
nor U3197 (N_3197,In_1916,In_62);
or U3198 (N_3198,In_1486,In_815);
nor U3199 (N_3199,In_860,In_1862);
and U3200 (N_3200,In_1872,In_1642);
and U3201 (N_3201,In_1385,In_776);
xnor U3202 (N_3202,In_1547,In_378);
nor U3203 (N_3203,In_1078,In_1779);
and U3204 (N_3204,In_1655,In_566);
nor U3205 (N_3205,In_194,In_162);
nor U3206 (N_3206,In_1191,In_436);
or U3207 (N_3207,In_1832,In_421);
and U3208 (N_3208,In_1018,In_85);
nor U3209 (N_3209,In_853,In_639);
and U3210 (N_3210,In_1765,In_527);
or U3211 (N_3211,In_1440,In_1547);
nand U3212 (N_3212,In_1351,In_1743);
or U3213 (N_3213,In_1075,In_1315);
xnor U3214 (N_3214,In_279,In_671);
nor U3215 (N_3215,In_4,In_1257);
nand U3216 (N_3216,In_1977,In_721);
or U3217 (N_3217,In_831,In_1055);
or U3218 (N_3218,In_271,In_793);
and U3219 (N_3219,In_1118,In_1371);
and U3220 (N_3220,In_898,In_1037);
nand U3221 (N_3221,In_1985,In_342);
or U3222 (N_3222,In_1224,In_824);
or U3223 (N_3223,In_736,In_1899);
or U3224 (N_3224,In_573,In_1914);
nor U3225 (N_3225,In_56,In_1924);
or U3226 (N_3226,In_1301,In_1492);
and U3227 (N_3227,In_404,In_184);
nand U3228 (N_3228,In_1418,In_1772);
nand U3229 (N_3229,In_1989,In_1863);
or U3230 (N_3230,In_828,In_401);
nand U3231 (N_3231,In_1492,In_1229);
nor U3232 (N_3232,In_653,In_608);
or U3233 (N_3233,In_822,In_524);
nand U3234 (N_3234,In_1696,In_1334);
and U3235 (N_3235,In_1871,In_897);
or U3236 (N_3236,In_1063,In_1326);
or U3237 (N_3237,In_1608,In_1425);
or U3238 (N_3238,In_817,In_1797);
or U3239 (N_3239,In_891,In_251);
and U3240 (N_3240,In_1872,In_1161);
or U3241 (N_3241,In_1792,In_492);
nand U3242 (N_3242,In_1748,In_472);
and U3243 (N_3243,In_150,In_1553);
and U3244 (N_3244,In_151,In_1016);
xor U3245 (N_3245,In_594,In_1086);
xor U3246 (N_3246,In_888,In_1265);
nor U3247 (N_3247,In_347,In_866);
nor U3248 (N_3248,In_1827,In_1789);
xnor U3249 (N_3249,In_1156,In_500);
and U3250 (N_3250,In_911,In_347);
and U3251 (N_3251,In_573,In_1843);
nand U3252 (N_3252,In_1451,In_1045);
nand U3253 (N_3253,In_1556,In_1921);
and U3254 (N_3254,In_86,In_1735);
xor U3255 (N_3255,In_668,In_871);
xor U3256 (N_3256,In_465,In_54);
or U3257 (N_3257,In_193,In_142);
xnor U3258 (N_3258,In_678,In_1110);
and U3259 (N_3259,In_940,In_1413);
nor U3260 (N_3260,In_99,In_95);
nor U3261 (N_3261,In_1978,In_983);
or U3262 (N_3262,In_909,In_1792);
nand U3263 (N_3263,In_579,In_801);
xor U3264 (N_3264,In_126,In_1793);
or U3265 (N_3265,In_1104,In_1055);
and U3266 (N_3266,In_898,In_590);
or U3267 (N_3267,In_1892,In_1988);
or U3268 (N_3268,In_1443,In_1668);
or U3269 (N_3269,In_1103,In_586);
and U3270 (N_3270,In_1812,In_409);
or U3271 (N_3271,In_439,In_1578);
and U3272 (N_3272,In_1496,In_442);
nand U3273 (N_3273,In_405,In_1880);
and U3274 (N_3274,In_1718,In_691);
nand U3275 (N_3275,In_1280,In_1346);
nor U3276 (N_3276,In_104,In_15);
and U3277 (N_3277,In_1594,In_1256);
or U3278 (N_3278,In_1621,In_404);
xnor U3279 (N_3279,In_1700,In_356);
xnor U3280 (N_3280,In_2,In_1390);
or U3281 (N_3281,In_575,In_1802);
nor U3282 (N_3282,In_178,In_1510);
nand U3283 (N_3283,In_1324,In_1798);
xor U3284 (N_3284,In_1493,In_1621);
nor U3285 (N_3285,In_164,In_1636);
and U3286 (N_3286,In_537,In_1606);
and U3287 (N_3287,In_1997,In_1137);
and U3288 (N_3288,In_772,In_318);
and U3289 (N_3289,In_1741,In_33);
or U3290 (N_3290,In_888,In_1285);
nand U3291 (N_3291,In_765,In_691);
and U3292 (N_3292,In_227,In_469);
and U3293 (N_3293,In_1553,In_652);
xor U3294 (N_3294,In_1395,In_14);
nor U3295 (N_3295,In_1227,In_463);
or U3296 (N_3296,In_56,In_838);
or U3297 (N_3297,In_930,In_1712);
nor U3298 (N_3298,In_476,In_667);
and U3299 (N_3299,In_495,In_1494);
nor U3300 (N_3300,In_1055,In_493);
nor U3301 (N_3301,In_1991,In_533);
xnor U3302 (N_3302,In_1033,In_1706);
nand U3303 (N_3303,In_725,In_175);
or U3304 (N_3304,In_881,In_1404);
or U3305 (N_3305,In_1719,In_1934);
xnor U3306 (N_3306,In_1221,In_133);
and U3307 (N_3307,In_983,In_1087);
or U3308 (N_3308,In_1304,In_1748);
nor U3309 (N_3309,In_483,In_1622);
or U3310 (N_3310,In_703,In_279);
nor U3311 (N_3311,In_1406,In_1138);
or U3312 (N_3312,In_1563,In_766);
xnor U3313 (N_3313,In_1580,In_297);
nor U3314 (N_3314,In_463,In_112);
and U3315 (N_3315,In_1345,In_1361);
nand U3316 (N_3316,In_95,In_1599);
nand U3317 (N_3317,In_316,In_750);
and U3318 (N_3318,In_352,In_629);
xnor U3319 (N_3319,In_254,In_819);
nor U3320 (N_3320,In_1129,In_1621);
xnor U3321 (N_3321,In_1582,In_1533);
and U3322 (N_3322,In_1293,In_848);
xor U3323 (N_3323,In_285,In_540);
nand U3324 (N_3324,In_1507,In_1602);
nor U3325 (N_3325,In_1809,In_1262);
and U3326 (N_3326,In_1814,In_1831);
and U3327 (N_3327,In_809,In_459);
or U3328 (N_3328,In_1016,In_1295);
nor U3329 (N_3329,In_267,In_955);
nor U3330 (N_3330,In_1083,In_85);
nand U3331 (N_3331,In_1626,In_382);
nor U3332 (N_3332,In_1539,In_1536);
nor U3333 (N_3333,In_1297,In_702);
xor U3334 (N_3334,In_1569,In_1635);
nor U3335 (N_3335,In_806,In_712);
nand U3336 (N_3336,In_830,In_512);
xor U3337 (N_3337,In_1636,In_995);
and U3338 (N_3338,In_1022,In_800);
and U3339 (N_3339,In_1810,In_627);
or U3340 (N_3340,In_1968,In_297);
or U3341 (N_3341,In_1751,In_946);
xnor U3342 (N_3342,In_1906,In_796);
or U3343 (N_3343,In_1788,In_560);
or U3344 (N_3344,In_214,In_1148);
or U3345 (N_3345,In_676,In_539);
nand U3346 (N_3346,In_1445,In_1606);
nor U3347 (N_3347,In_1590,In_425);
xnor U3348 (N_3348,In_469,In_1807);
xnor U3349 (N_3349,In_861,In_1042);
or U3350 (N_3350,In_905,In_257);
or U3351 (N_3351,In_255,In_744);
xor U3352 (N_3352,In_585,In_830);
nand U3353 (N_3353,In_808,In_1179);
nand U3354 (N_3354,In_11,In_1159);
or U3355 (N_3355,In_824,In_464);
xor U3356 (N_3356,In_688,In_1726);
and U3357 (N_3357,In_1281,In_690);
or U3358 (N_3358,In_625,In_1851);
nand U3359 (N_3359,In_147,In_952);
or U3360 (N_3360,In_389,In_1937);
or U3361 (N_3361,In_818,In_849);
nor U3362 (N_3362,In_1242,In_1776);
and U3363 (N_3363,In_1896,In_993);
or U3364 (N_3364,In_604,In_1649);
xnor U3365 (N_3365,In_1813,In_863);
nor U3366 (N_3366,In_1470,In_1932);
nor U3367 (N_3367,In_1870,In_119);
nand U3368 (N_3368,In_160,In_994);
xnor U3369 (N_3369,In_498,In_642);
xor U3370 (N_3370,In_1023,In_1122);
and U3371 (N_3371,In_1144,In_746);
nand U3372 (N_3372,In_148,In_137);
or U3373 (N_3373,In_452,In_1917);
nor U3374 (N_3374,In_1945,In_1889);
or U3375 (N_3375,In_1171,In_1519);
and U3376 (N_3376,In_1005,In_807);
and U3377 (N_3377,In_1025,In_126);
and U3378 (N_3378,In_948,In_499);
xor U3379 (N_3379,In_6,In_1575);
nand U3380 (N_3380,In_261,In_1010);
nand U3381 (N_3381,In_197,In_1955);
nor U3382 (N_3382,In_1815,In_908);
xnor U3383 (N_3383,In_1928,In_228);
xor U3384 (N_3384,In_1286,In_1118);
xnor U3385 (N_3385,In_127,In_873);
nor U3386 (N_3386,In_115,In_1432);
or U3387 (N_3387,In_1965,In_1188);
nand U3388 (N_3388,In_1063,In_1046);
nand U3389 (N_3389,In_1479,In_1914);
nand U3390 (N_3390,In_654,In_1837);
nand U3391 (N_3391,In_816,In_1033);
nor U3392 (N_3392,In_1894,In_1066);
or U3393 (N_3393,In_1333,In_1207);
or U3394 (N_3394,In_511,In_1388);
xor U3395 (N_3395,In_75,In_1433);
nor U3396 (N_3396,In_1912,In_1283);
nor U3397 (N_3397,In_853,In_218);
or U3398 (N_3398,In_246,In_1798);
xnor U3399 (N_3399,In_242,In_235);
nor U3400 (N_3400,In_926,In_233);
nand U3401 (N_3401,In_1002,In_121);
xor U3402 (N_3402,In_974,In_1128);
nand U3403 (N_3403,In_1420,In_384);
nor U3404 (N_3404,In_372,In_796);
xor U3405 (N_3405,In_425,In_1094);
nor U3406 (N_3406,In_56,In_787);
xnor U3407 (N_3407,In_1289,In_1106);
and U3408 (N_3408,In_54,In_1338);
nand U3409 (N_3409,In_1502,In_1018);
and U3410 (N_3410,In_725,In_695);
nand U3411 (N_3411,In_1104,In_79);
xor U3412 (N_3412,In_111,In_360);
nor U3413 (N_3413,In_47,In_860);
nor U3414 (N_3414,In_1862,In_996);
and U3415 (N_3415,In_839,In_916);
and U3416 (N_3416,In_758,In_1850);
nand U3417 (N_3417,In_241,In_396);
xor U3418 (N_3418,In_840,In_136);
nand U3419 (N_3419,In_645,In_338);
xnor U3420 (N_3420,In_1542,In_558);
and U3421 (N_3421,In_1798,In_610);
and U3422 (N_3422,In_1434,In_1889);
or U3423 (N_3423,In_998,In_1084);
nand U3424 (N_3424,In_18,In_1081);
nand U3425 (N_3425,In_1211,In_1094);
or U3426 (N_3426,In_301,In_1231);
and U3427 (N_3427,In_1585,In_1502);
and U3428 (N_3428,In_1973,In_726);
xnor U3429 (N_3429,In_606,In_1561);
or U3430 (N_3430,In_1061,In_173);
nand U3431 (N_3431,In_1567,In_1242);
or U3432 (N_3432,In_34,In_405);
nand U3433 (N_3433,In_1895,In_1940);
and U3434 (N_3434,In_1531,In_1601);
and U3435 (N_3435,In_1192,In_1328);
nor U3436 (N_3436,In_1253,In_808);
nand U3437 (N_3437,In_474,In_1389);
nand U3438 (N_3438,In_1856,In_1392);
nand U3439 (N_3439,In_1005,In_856);
nand U3440 (N_3440,In_930,In_96);
xor U3441 (N_3441,In_914,In_1958);
and U3442 (N_3442,In_1701,In_126);
or U3443 (N_3443,In_1102,In_80);
or U3444 (N_3444,In_92,In_308);
xor U3445 (N_3445,In_1948,In_1432);
nor U3446 (N_3446,In_1075,In_1778);
nor U3447 (N_3447,In_714,In_1759);
and U3448 (N_3448,In_1895,In_540);
or U3449 (N_3449,In_132,In_1728);
nand U3450 (N_3450,In_977,In_954);
nor U3451 (N_3451,In_1670,In_1465);
or U3452 (N_3452,In_392,In_1563);
nand U3453 (N_3453,In_237,In_545);
nor U3454 (N_3454,In_599,In_990);
nor U3455 (N_3455,In_1253,In_1497);
or U3456 (N_3456,In_608,In_1752);
nand U3457 (N_3457,In_497,In_423);
nand U3458 (N_3458,In_1881,In_1937);
and U3459 (N_3459,In_91,In_1918);
nand U3460 (N_3460,In_329,In_1320);
or U3461 (N_3461,In_518,In_319);
xor U3462 (N_3462,In_854,In_511);
nor U3463 (N_3463,In_689,In_436);
or U3464 (N_3464,In_1730,In_1965);
or U3465 (N_3465,In_1267,In_822);
xnor U3466 (N_3466,In_1242,In_1815);
and U3467 (N_3467,In_870,In_1610);
xor U3468 (N_3468,In_1808,In_1305);
nand U3469 (N_3469,In_951,In_1210);
nor U3470 (N_3470,In_720,In_1194);
xnor U3471 (N_3471,In_1162,In_390);
and U3472 (N_3472,In_615,In_534);
or U3473 (N_3473,In_1831,In_1200);
xor U3474 (N_3474,In_136,In_941);
nor U3475 (N_3475,In_732,In_830);
nor U3476 (N_3476,In_200,In_1811);
and U3477 (N_3477,In_1008,In_1511);
nor U3478 (N_3478,In_272,In_1111);
or U3479 (N_3479,In_1566,In_87);
and U3480 (N_3480,In_1878,In_1710);
nor U3481 (N_3481,In_1151,In_804);
nand U3482 (N_3482,In_31,In_205);
or U3483 (N_3483,In_1889,In_48);
or U3484 (N_3484,In_1547,In_1710);
and U3485 (N_3485,In_702,In_1714);
or U3486 (N_3486,In_1801,In_136);
nor U3487 (N_3487,In_163,In_813);
nand U3488 (N_3488,In_464,In_1922);
xor U3489 (N_3489,In_1378,In_1611);
nand U3490 (N_3490,In_1701,In_195);
or U3491 (N_3491,In_1136,In_672);
xnor U3492 (N_3492,In_868,In_522);
and U3493 (N_3493,In_1549,In_1474);
or U3494 (N_3494,In_1476,In_1821);
nor U3495 (N_3495,In_859,In_1232);
and U3496 (N_3496,In_181,In_1834);
xor U3497 (N_3497,In_1825,In_1806);
or U3498 (N_3498,In_1864,In_197);
xnor U3499 (N_3499,In_1263,In_547);
or U3500 (N_3500,In_1132,In_854);
nand U3501 (N_3501,In_1836,In_295);
and U3502 (N_3502,In_1237,In_1802);
xnor U3503 (N_3503,In_51,In_1451);
or U3504 (N_3504,In_1424,In_1566);
xor U3505 (N_3505,In_1832,In_5);
xnor U3506 (N_3506,In_1865,In_1221);
xor U3507 (N_3507,In_1029,In_192);
or U3508 (N_3508,In_999,In_1990);
or U3509 (N_3509,In_1797,In_1445);
nor U3510 (N_3510,In_1827,In_1980);
nor U3511 (N_3511,In_47,In_1413);
xnor U3512 (N_3512,In_795,In_1921);
nor U3513 (N_3513,In_1986,In_1286);
nor U3514 (N_3514,In_789,In_1798);
nand U3515 (N_3515,In_1921,In_952);
nand U3516 (N_3516,In_173,In_296);
nand U3517 (N_3517,In_1322,In_1946);
xor U3518 (N_3518,In_1011,In_346);
nand U3519 (N_3519,In_1988,In_1395);
nand U3520 (N_3520,In_1792,In_672);
nor U3521 (N_3521,In_612,In_1793);
xnor U3522 (N_3522,In_325,In_1485);
nand U3523 (N_3523,In_3,In_573);
xnor U3524 (N_3524,In_848,In_1382);
nand U3525 (N_3525,In_276,In_445);
or U3526 (N_3526,In_241,In_1035);
nor U3527 (N_3527,In_1866,In_1201);
xnor U3528 (N_3528,In_1861,In_1312);
or U3529 (N_3529,In_1724,In_1905);
nor U3530 (N_3530,In_1987,In_1482);
nor U3531 (N_3531,In_522,In_566);
xnor U3532 (N_3532,In_1882,In_1681);
or U3533 (N_3533,In_692,In_1498);
nor U3534 (N_3534,In_622,In_229);
and U3535 (N_3535,In_1744,In_1730);
xnor U3536 (N_3536,In_1095,In_1686);
nand U3537 (N_3537,In_23,In_609);
xnor U3538 (N_3538,In_47,In_776);
nor U3539 (N_3539,In_77,In_1315);
nor U3540 (N_3540,In_360,In_1754);
nor U3541 (N_3541,In_1691,In_441);
nor U3542 (N_3542,In_494,In_1447);
nor U3543 (N_3543,In_485,In_717);
or U3544 (N_3544,In_477,In_1578);
or U3545 (N_3545,In_1466,In_1327);
nor U3546 (N_3546,In_506,In_1091);
nor U3547 (N_3547,In_1338,In_228);
nand U3548 (N_3548,In_743,In_1315);
and U3549 (N_3549,In_494,In_1310);
nand U3550 (N_3550,In_1972,In_733);
xnor U3551 (N_3551,In_901,In_119);
and U3552 (N_3552,In_728,In_1120);
and U3553 (N_3553,In_1749,In_701);
nand U3554 (N_3554,In_1937,In_1637);
xor U3555 (N_3555,In_375,In_1255);
xor U3556 (N_3556,In_504,In_1377);
nand U3557 (N_3557,In_172,In_194);
xnor U3558 (N_3558,In_1985,In_1309);
nor U3559 (N_3559,In_180,In_525);
nor U3560 (N_3560,In_1038,In_1942);
and U3561 (N_3561,In_1634,In_534);
xnor U3562 (N_3562,In_1869,In_1537);
nor U3563 (N_3563,In_1673,In_42);
nand U3564 (N_3564,In_1477,In_1381);
and U3565 (N_3565,In_49,In_1947);
nand U3566 (N_3566,In_409,In_1195);
or U3567 (N_3567,In_999,In_1888);
and U3568 (N_3568,In_1639,In_182);
xor U3569 (N_3569,In_1941,In_280);
nand U3570 (N_3570,In_187,In_153);
or U3571 (N_3571,In_252,In_1496);
nand U3572 (N_3572,In_1667,In_1566);
nand U3573 (N_3573,In_394,In_654);
and U3574 (N_3574,In_473,In_1780);
xnor U3575 (N_3575,In_1980,In_1284);
nor U3576 (N_3576,In_301,In_1724);
xnor U3577 (N_3577,In_1926,In_1469);
and U3578 (N_3578,In_1890,In_1902);
nor U3579 (N_3579,In_1918,In_1951);
and U3580 (N_3580,In_1396,In_1697);
nor U3581 (N_3581,In_426,In_1820);
nand U3582 (N_3582,In_1075,In_1843);
xnor U3583 (N_3583,In_1753,In_658);
xor U3584 (N_3584,In_1943,In_1798);
nor U3585 (N_3585,In_699,In_1526);
xnor U3586 (N_3586,In_1592,In_32);
xnor U3587 (N_3587,In_305,In_1304);
nand U3588 (N_3588,In_954,In_667);
and U3589 (N_3589,In_1347,In_1387);
xor U3590 (N_3590,In_427,In_789);
xor U3591 (N_3591,In_1663,In_568);
and U3592 (N_3592,In_1920,In_394);
or U3593 (N_3593,In_1583,In_1733);
or U3594 (N_3594,In_1517,In_1391);
nor U3595 (N_3595,In_209,In_806);
xnor U3596 (N_3596,In_1145,In_9);
nand U3597 (N_3597,In_1012,In_774);
nand U3598 (N_3598,In_1667,In_1879);
nor U3599 (N_3599,In_11,In_318);
xnor U3600 (N_3600,In_1151,In_1266);
nand U3601 (N_3601,In_636,In_1122);
and U3602 (N_3602,In_316,In_262);
xor U3603 (N_3603,In_1229,In_23);
xnor U3604 (N_3604,In_218,In_397);
nand U3605 (N_3605,In_1402,In_1730);
nor U3606 (N_3606,In_1559,In_1624);
or U3607 (N_3607,In_1324,In_914);
nor U3608 (N_3608,In_1331,In_988);
or U3609 (N_3609,In_134,In_1943);
and U3610 (N_3610,In_1499,In_1202);
nand U3611 (N_3611,In_1385,In_1109);
nand U3612 (N_3612,In_1897,In_136);
xnor U3613 (N_3613,In_1551,In_200);
and U3614 (N_3614,In_1696,In_1518);
and U3615 (N_3615,In_1938,In_735);
nor U3616 (N_3616,In_928,In_1304);
nor U3617 (N_3617,In_77,In_1444);
and U3618 (N_3618,In_1799,In_653);
xnor U3619 (N_3619,In_851,In_1645);
nand U3620 (N_3620,In_632,In_1449);
and U3621 (N_3621,In_746,In_444);
xor U3622 (N_3622,In_1749,In_1082);
nand U3623 (N_3623,In_1319,In_899);
nor U3624 (N_3624,In_1229,In_422);
nor U3625 (N_3625,In_161,In_455);
xor U3626 (N_3626,In_1583,In_1342);
nand U3627 (N_3627,In_959,In_1819);
and U3628 (N_3628,In_1409,In_635);
nand U3629 (N_3629,In_1606,In_1097);
nand U3630 (N_3630,In_281,In_1286);
or U3631 (N_3631,In_306,In_1778);
xnor U3632 (N_3632,In_1902,In_111);
or U3633 (N_3633,In_1508,In_471);
or U3634 (N_3634,In_1355,In_1815);
nand U3635 (N_3635,In_1957,In_554);
and U3636 (N_3636,In_1237,In_566);
nor U3637 (N_3637,In_883,In_45);
nand U3638 (N_3638,In_278,In_414);
nor U3639 (N_3639,In_116,In_939);
and U3640 (N_3640,In_748,In_976);
nor U3641 (N_3641,In_1424,In_526);
xnor U3642 (N_3642,In_1180,In_1355);
nor U3643 (N_3643,In_1358,In_169);
and U3644 (N_3644,In_1353,In_1492);
xor U3645 (N_3645,In_39,In_1923);
xor U3646 (N_3646,In_167,In_1036);
and U3647 (N_3647,In_1939,In_279);
and U3648 (N_3648,In_484,In_1431);
and U3649 (N_3649,In_509,In_34);
and U3650 (N_3650,In_107,In_1845);
or U3651 (N_3651,In_827,In_125);
nand U3652 (N_3652,In_1533,In_544);
and U3653 (N_3653,In_326,In_1877);
xor U3654 (N_3654,In_1393,In_1729);
nand U3655 (N_3655,In_1317,In_1378);
nor U3656 (N_3656,In_1693,In_869);
xor U3657 (N_3657,In_1025,In_454);
or U3658 (N_3658,In_440,In_1048);
nand U3659 (N_3659,In_74,In_184);
or U3660 (N_3660,In_1299,In_1618);
and U3661 (N_3661,In_378,In_113);
xnor U3662 (N_3662,In_1196,In_944);
or U3663 (N_3663,In_1537,In_1739);
and U3664 (N_3664,In_62,In_1003);
nor U3665 (N_3665,In_1382,In_1209);
xor U3666 (N_3666,In_177,In_1804);
nor U3667 (N_3667,In_1396,In_527);
or U3668 (N_3668,In_814,In_1118);
nor U3669 (N_3669,In_220,In_589);
nand U3670 (N_3670,In_131,In_1620);
or U3671 (N_3671,In_1282,In_981);
xnor U3672 (N_3672,In_1778,In_893);
and U3673 (N_3673,In_1453,In_930);
or U3674 (N_3674,In_1924,In_1767);
and U3675 (N_3675,In_53,In_247);
or U3676 (N_3676,In_929,In_307);
or U3677 (N_3677,In_1973,In_785);
nor U3678 (N_3678,In_1227,In_851);
nand U3679 (N_3679,In_97,In_324);
and U3680 (N_3680,In_1140,In_1067);
xnor U3681 (N_3681,In_1131,In_1621);
and U3682 (N_3682,In_1892,In_1319);
nor U3683 (N_3683,In_1648,In_724);
nor U3684 (N_3684,In_763,In_497);
nand U3685 (N_3685,In_584,In_1728);
and U3686 (N_3686,In_596,In_190);
nand U3687 (N_3687,In_1610,In_349);
xor U3688 (N_3688,In_1893,In_1609);
xnor U3689 (N_3689,In_1610,In_1326);
nand U3690 (N_3690,In_1199,In_1873);
or U3691 (N_3691,In_404,In_1188);
or U3692 (N_3692,In_1312,In_1716);
or U3693 (N_3693,In_597,In_186);
nor U3694 (N_3694,In_1474,In_1769);
or U3695 (N_3695,In_752,In_163);
nor U3696 (N_3696,In_645,In_1742);
xor U3697 (N_3697,In_1182,In_1926);
nand U3698 (N_3698,In_1380,In_513);
and U3699 (N_3699,In_21,In_725);
or U3700 (N_3700,In_1548,In_1731);
nor U3701 (N_3701,In_586,In_739);
nor U3702 (N_3702,In_254,In_1864);
nor U3703 (N_3703,In_1743,In_612);
xor U3704 (N_3704,In_1390,In_61);
or U3705 (N_3705,In_1364,In_463);
and U3706 (N_3706,In_1088,In_1732);
and U3707 (N_3707,In_501,In_1997);
or U3708 (N_3708,In_1089,In_1296);
nor U3709 (N_3709,In_655,In_762);
nor U3710 (N_3710,In_1100,In_190);
nand U3711 (N_3711,In_723,In_1883);
nand U3712 (N_3712,In_48,In_797);
nor U3713 (N_3713,In_802,In_36);
nand U3714 (N_3714,In_1087,In_679);
xnor U3715 (N_3715,In_1420,In_821);
nor U3716 (N_3716,In_1425,In_1351);
nor U3717 (N_3717,In_507,In_1543);
xnor U3718 (N_3718,In_1926,In_877);
nor U3719 (N_3719,In_1628,In_1514);
or U3720 (N_3720,In_1983,In_363);
xor U3721 (N_3721,In_933,In_1409);
xor U3722 (N_3722,In_1849,In_660);
xor U3723 (N_3723,In_1954,In_311);
nand U3724 (N_3724,In_268,In_86);
nand U3725 (N_3725,In_1107,In_1076);
xor U3726 (N_3726,In_572,In_57);
nand U3727 (N_3727,In_1146,In_1543);
nand U3728 (N_3728,In_1226,In_1526);
nand U3729 (N_3729,In_453,In_762);
nor U3730 (N_3730,In_1308,In_1767);
nand U3731 (N_3731,In_1533,In_146);
or U3732 (N_3732,In_541,In_637);
or U3733 (N_3733,In_1084,In_110);
and U3734 (N_3734,In_257,In_44);
nor U3735 (N_3735,In_345,In_535);
xnor U3736 (N_3736,In_295,In_1596);
xnor U3737 (N_3737,In_226,In_187);
and U3738 (N_3738,In_560,In_1598);
nor U3739 (N_3739,In_1565,In_1167);
xnor U3740 (N_3740,In_42,In_906);
xnor U3741 (N_3741,In_1674,In_294);
nor U3742 (N_3742,In_946,In_747);
and U3743 (N_3743,In_1310,In_51);
and U3744 (N_3744,In_97,In_1401);
xor U3745 (N_3745,In_1931,In_1761);
nor U3746 (N_3746,In_898,In_1259);
nand U3747 (N_3747,In_148,In_399);
xnor U3748 (N_3748,In_201,In_70);
or U3749 (N_3749,In_529,In_1010);
nand U3750 (N_3750,In_1540,In_1552);
xor U3751 (N_3751,In_375,In_423);
nor U3752 (N_3752,In_1016,In_612);
and U3753 (N_3753,In_285,In_1264);
nor U3754 (N_3754,In_167,In_446);
nand U3755 (N_3755,In_1546,In_224);
and U3756 (N_3756,In_767,In_1283);
or U3757 (N_3757,In_1224,In_904);
or U3758 (N_3758,In_630,In_1155);
xor U3759 (N_3759,In_315,In_1756);
xnor U3760 (N_3760,In_216,In_1515);
xor U3761 (N_3761,In_393,In_155);
and U3762 (N_3762,In_867,In_1552);
nand U3763 (N_3763,In_913,In_108);
and U3764 (N_3764,In_799,In_1602);
or U3765 (N_3765,In_1923,In_1130);
or U3766 (N_3766,In_292,In_169);
nor U3767 (N_3767,In_1860,In_1792);
or U3768 (N_3768,In_1799,In_339);
nor U3769 (N_3769,In_1221,In_692);
nand U3770 (N_3770,In_927,In_346);
or U3771 (N_3771,In_1775,In_855);
xnor U3772 (N_3772,In_1636,In_453);
and U3773 (N_3773,In_1055,In_947);
xor U3774 (N_3774,In_1339,In_404);
and U3775 (N_3775,In_1925,In_171);
xnor U3776 (N_3776,In_1817,In_1644);
nor U3777 (N_3777,In_335,In_236);
or U3778 (N_3778,In_1471,In_1476);
nand U3779 (N_3779,In_1546,In_941);
and U3780 (N_3780,In_369,In_167);
nand U3781 (N_3781,In_227,In_1248);
nand U3782 (N_3782,In_760,In_1688);
and U3783 (N_3783,In_756,In_1689);
nand U3784 (N_3784,In_447,In_685);
nand U3785 (N_3785,In_667,In_983);
nand U3786 (N_3786,In_970,In_1844);
nand U3787 (N_3787,In_1999,In_1196);
xnor U3788 (N_3788,In_1200,In_682);
nand U3789 (N_3789,In_145,In_1299);
nand U3790 (N_3790,In_1624,In_687);
nor U3791 (N_3791,In_1023,In_695);
nor U3792 (N_3792,In_1746,In_1689);
nor U3793 (N_3793,In_706,In_1657);
nand U3794 (N_3794,In_1780,In_1803);
and U3795 (N_3795,In_1729,In_1961);
nor U3796 (N_3796,In_1679,In_1064);
and U3797 (N_3797,In_32,In_1155);
and U3798 (N_3798,In_1084,In_276);
or U3799 (N_3799,In_1539,In_1301);
and U3800 (N_3800,In_705,In_1119);
nand U3801 (N_3801,In_90,In_1172);
xor U3802 (N_3802,In_1958,In_517);
and U3803 (N_3803,In_175,In_1954);
xor U3804 (N_3804,In_1016,In_930);
and U3805 (N_3805,In_958,In_1799);
nor U3806 (N_3806,In_1827,In_1659);
nand U3807 (N_3807,In_873,In_1658);
nand U3808 (N_3808,In_824,In_1307);
and U3809 (N_3809,In_1608,In_529);
xor U3810 (N_3810,In_1964,In_394);
nand U3811 (N_3811,In_1121,In_227);
xnor U3812 (N_3812,In_259,In_910);
xor U3813 (N_3813,In_234,In_1353);
or U3814 (N_3814,In_1793,In_534);
nor U3815 (N_3815,In_1281,In_1229);
and U3816 (N_3816,In_988,In_1175);
or U3817 (N_3817,In_43,In_989);
xnor U3818 (N_3818,In_461,In_1035);
nor U3819 (N_3819,In_23,In_1909);
or U3820 (N_3820,In_1933,In_1527);
xnor U3821 (N_3821,In_1261,In_1669);
nand U3822 (N_3822,In_42,In_1745);
and U3823 (N_3823,In_1200,In_1815);
or U3824 (N_3824,In_1753,In_926);
and U3825 (N_3825,In_151,In_724);
xnor U3826 (N_3826,In_931,In_1084);
nand U3827 (N_3827,In_945,In_1578);
nand U3828 (N_3828,In_1096,In_304);
or U3829 (N_3829,In_1204,In_41);
nor U3830 (N_3830,In_1397,In_6);
xnor U3831 (N_3831,In_597,In_748);
xnor U3832 (N_3832,In_567,In_272);
or U3833 (N_3833,In_96,In_1142);
or U3834 (N_3834,In_254,In_690);
or U3835 (N_3835,In_1700,In_1845);
xnor U3836 (N_3836,In_534,In_805);
or U3837 (N_3837,In_1286,In_72);
xnor U3838 (N_3838,In_33,In_351);
xor U3839 (N_3839,In_1896,In_1472);
nor U3840 (N_3840,In_485,In_1840);
nand U3841 (N_3841,In_1453,In_1611);
nand U3842 (N_3842,In_1975,In_1566);
and U3843 (N_3843,In_110,In_1045);
and U3844 (N_3844,In_679,In_48);
nand U3845 (N_3845,In_744,In_1788);
xnor U3846 (N_3846,In_1966,In_1039);
nand U3847 (N_3847,In_738,In_52);
or U3848 (N_3848,In_1857,In_980);
nor U3849 (N_3849,In_1852,In_782);
and U3850 (N_3850,In_1472,In_1228);
and U3851 (N_3851,In_453,In_309);
nand U3852 (N_3852,In_1201,In_881);
nand U3853 (N_3853,In_571,In_1471);
nand U3854 (N_3854,In_848,In_1381);
and U3855 (N_3855,In_1995,In_1971);
nor U3856 (N_3856,In_1929,In_1361);
xnor U3857 (N_3857,In_1196,In_498);
or U3858 (N_3858,In_1049,In_1893);
or U3859 (N_3859,In_1261,In_1090);
xnor U3860 (N_3860,In_391,In_1762);
or U3861 (N_3861,In_736,In_42);
xnor U3862 (N_3862,In_1035,In_224);
xnor U3863 (N_3863,In_898,In_541);
nor U3864 (N_3864,In_1179,In_1822);
xor U3865 (N_3865,In_501,In_1025);
nor U3866 (N_3866,In_1002,In_1236);
and U3867 (N_3867,In_921,In_675);
nor U3868 (N_3868,In_1815,In_1840);
nor U3869 (N_3869,In_761,In_312);
and U3870 (N_3870,In_1243,In_1127);
nand U3871 (N_3871,In_246,In_838);
or U3872 (N_3872,In_1138,In_1504);
and U3873 (N_3873,In_409,In_922);
or U3874 (N_3874,In_1962,In_1495);
and U3875 (N_3875,In_586,In_384);
and U3876 (N_3876,In_1818,In_32);
xnor U3877 (N_3877,In_915,In_1377);
nand U3878 (N_3878,In_105,In_1625);
nand U3879 (N_3879,In_344,In_1809);
or U3880 (N_3880,In_960,In_476);
or U3881 (N_3881,In_1808,In_1606);
xor U3882 (N_3882,In_1640,In_327);
xnor U3883 (N_3883,In_42,In_1837);
and U3884 (N_3884,In_1880,In_1036);
nor U3885 (N_3885,In_38,In_1143);
or U3886 (N_3886,In_241,In_499);
or U3887 (N_3887,In_501,In_1518);
or U3888 (N_3888,In_1125,In_57);
xnor U3889 (N_3889,In_1630,In_1805);
nand U3890 (N_3890,In_864,In_1651);
xnor U3891 (N_3891,In_954,In_1781);
or U3892 (N_3892,In_892,In_348);
or U3893 (N_3893,In_1678,In_1487);
and U3894 (N_3894,In_1529,In_1054);
nand U3895 (N_3895,In_1428,In_1783);
xnor U3896 (N_3896,In_53,In_833);
and U3897 (N_3897,In_1868,In_1327);
and U3898 (N_3898,In_1053,In_1992);
or U3899 (N_3899,In_1375,In_889);
xnor U3900 (N_3900,In_1327,In_976);
nand U3901 (N_3901,In_1292,In_480);
nor U3902 (N_3902,In_629,In_568);
and U3903 (N_3903,In_256,In_867);
xor U3904 (N_3904,In_1003,In_1101);
or U3905 (N_3905,In_1834,In_449);
nand U3906 (N_3906,In_1717,In_1103);
and U3907 (N_3907,In_158,In_102);
nand U3908 (N_3908,In_918,In_882);
and U3909 (N_3909,In_646,In_258);
xor U3910 (N_3910,In_884,In_1669);
nand U3911 (N_3911,In_1857,In_63);
nor U3912 (N_3912,In_139,In_1489);
nand U3913 (N_3913,In_651,In_1321);
nand U3914 (N_3914,In_1994,In_1037);
and U3915 (N_3915,In_1733,In_23);
xnor U3916 (N_3916,In_1738,In_703);
or U3917 (N_3917,In_1822,In_349);
or U3918 (N_3918,In_1649,In_853);
or U3919 (N_3919,In_517,In_87);
xnor U3920 (N_3920,In_76,In_1454);
and U3921 (N_3921,In_723,In_89);
xnor U3922 (N_3922,In_674,In_74);
nor U3923 (N_3923,In_929,In_22);
and U3924 (N_3924,In_691,In_680);
nand U3925 (N_3925,In_809,In_1287);
xnor U3926 (N_3926,In_525,In_189);
nor U3927 (N_3927,In_441,In_1695);
nor U3928 (N_3928,In_69,In_55);
nor U3929 (N_3929,In_515,In_1332);
nand U3930 (N_3930,In_905,In_321);
nand U3931 (N_3931,In_1565,In_108);
nand U3932 (N_3932,In_1779,In_513);
nor U3933 (N_3933,In_1483,In_1458);
xor U3934 (N_3934,In_350,In_370);
nand U3935 (N_3935,In_146,In_837);
nor U3936 (N_3936,In_1506,In_744);
xnor U3937 (N_3937,In_807,In_1651);
and U3938 (N_3938,In_378,In_410);
nor U3939 (N_3939,In_1552,In_406);
and U3940 (N_3940,In_694,In_1575);
and U3941 (N_3941,In_1604,In_421);
xnor U3942 (N_3942,In_1282,In_2);
or U3943 (N_3943,In_556,In_1909);
nor U3944 (N_3944,In_1794,In_225);
xnor U3945 (N_3945,In_922,In_224);
and U3946 (N_3946,In_703,In_431);
and U3947 (N_3947,In_174,In_397);
or U3948 (N_3948,In_231,In_1535);
xor U3949 (N_3949,In_1434,In_405);
and U3950 (N_3950,In_1043,In_581);
nand U3951 (N_3951,In_148,In_768);
nor U3952 (N_3952,In_1215,In_1886);
or U3953 (N_3953,In_1147,In_1641);
xnor U3954 (N_3954,In_1864,In_146);
nor U3955 (N_3955,In_691,In_494);
and U3956 (N_3956,In_1125,In_1857);
xnor U3957 (N_3957,In_395,In_686);
nand U3958 (N_3958,In_714,In_1573);
xnor U3959 (N_3959,In_514,In_1783);
or U3960 (N_3960,In_1568,In_1742);
and U3961 (N_3961,In_553,In_454);
nor U3962 (N_3962,In_562,In_1373);
and U3963 (N_3963,In_1331,In_857);
nor U3964 (N_3964,In_1021,In_787);
nor U3965 (N_3965,In_1051,In_1982);
nor U3966 (N_3966,In_1835,In_876);
xor U3967 (N_3967,In_1785,In_1592);
nor U3968 (N_3968,In_1807,In_520);
nand U3969 (N_3969,In_1422,In_869);
xor U3970 (N_3970,In_1773,In_607);
and U3971 (N_3971,In_965,In_718);
nor U3972 (N_3972,In_1379,In_287);
and U3973 (N_3973,In_771,In_1474);
or U3974 (N_3974,In_1134,In_636);
or U3975 (N_3975,In_1269,In_784);
or U3976 (N_3976,In_1462,In_1152);
and U3977 (N_3977,In_1888,In_1371);
or U3978 (N_3978,In_712,In_1816);
nand U3979 (N_3979,In_1998,In_1074);
xnor U3980 (N_3980,In_1035,In_1996);
and U3981 (N_3981,In_840,In_483);
xor U3982 (N_3982,In_1210,In_312);
or U3983 (N_3983,In_1049,In_993);
xnor U3984 (N_3984,In_1544,In_159);
or U3985 (N_3985,In_1207,In_1992);
or U3986 (N_3986,In_142,In_1577);
or U3987 (N_3987,In_293,In_1062);
and U3988 (N_3988,In_565,In_1962);
nand U3989 (N_3989,In_1182,In_1985);
or U3990 (N_3990,In_1549,In_1871);
and U3991 (N_3991,In_752,In_49);
and U3992 (N_3992,In_6,In_1873);
xor U3993 (N_3993,In_1108,In_1346);
nand U3994 (N_3994,In_142,In_1113);
xnor U3995 (N_3995,In_598,In_534);
and U3996 (N_3996,In_477,In_849);
or U3997 (N_3997,In_350,In_373);
xnor U3998 (N_3998,In_1803,In_1644);
nor U3999 (N_3999,In_1387,In_1995);
nand U4000 (N_4000,In_1101,In_1802);
and U4001 (N_4001,In_1391,In_1961);
nand U4002 (N_4002,In_234,In_593);
nand U4003 (N_4003,In_962,In_1804);
and U4004 (N_4004,In_1790,In_917);
xor U4005 (N_4005,In_1643,In_659);
nand U4006 (N_4006,In_424,In_408);
nor U4007 (N_4007,In_137,In_279);
or U4008 (N_4008,In_794,In_1499);
nor U4009 (N_4009,In_536,In_1034);
nand U4010 (N_4010,In_617,In_584);
or U4011 (N_4011,In_1260,In_834);
nor U4012 (N_4012,In_1065,In_221);
xnor U4013 (N_4013,In_1510,In_1133);
xnor U4014 (N_4014,In_914,In_1507);
xor U4015 (N_4015,In_893,In_1997);
or U4016 (N_4016,In_437,In_1133);
xor U4017 (N_4017,In_1799,In_767);
nor U4018 (N_4018,In_1500,In_538);
nor U4019 (N_4019,In_1426,In_1678);
and U4020 (N_4020,In_1420,In_1600);
nand U4021 (N_4021,In_1741,In_691);
nor U4022 (N_4022,In_800,In_1353);
nand U4023 (N_4023,In_910,In_568);
nor U4024 (N_4024,In_318,In_204);
or U4025 (N_4025,In_1480,In_768);
and U4026 (N_4026,In_1413,In_644);
xnor U4027 (N_4027,In_1042,In_596);
xor U4028 (N_4028,In_1345,In_658);
and U4029 (N_4029,In_397,In_317);
and U4030 (N_4030,In_1936,In_1586);
or U4031 (N_4031,In_429,In_1092);
nor U4032 (N_4032,In_1731,In_630);
or U4033 (N_4033,In_1053,In_235);
xnor U4034 (N_4034,In_1492,In_430);
nand U4035 (N_4035,In_35,In_1738);
or U4036 (N_4036,In_1291,In_1469);
nor U4037 (N_4037,In_19,In_457);
nand U4038 (N_4038,In_94,In_1241);
xor U4039 (N_4039,In_1161,In_1931);
nor U4040 (N_4040,In_69,In_1476);
nand U4041 (N_4041,In_103,In_1795);
and U4042 (N_4042,In_1755,In_76);
xnor U4043 (N_4043,In_1982,In_262);
nand U4044 (N_4044,In_1911,In_1135);
nand U4045 (N_4045,In_1191,In_396);
nand U4046 (N_4046,In_1805,In_1312);
and U4047 (N_4047,In_1806,In_1848);
or U4048 (N_4048,In_1554,In_883);
or U4049 (N_4049,In_1066,In_1881);
or U4050 (N_4050,In_257,In_899);
nor U4051 (N_4051,In_1938,In_1994);
nor U4052 (N_4052,In_90,In_523);
xor U4053 (N_4053,In_1997,In_1948);
nand U4054 (N_4054,In_1873,In_942);
or U4055 (N_4055,In_312,In_1741);
xor U4056 (N_4056,In_485,In_1859);
nand U4057 (N_4057,In_1735,In_497);
nor U4058 (N_4058,In_1071,In_1197);
nor U4059 (N_4059,In_406,In_512);
or U4060 (N_4060,In_1160,In_1867);
and U4061 (N_4061,In_1562,In_1201);
and U4062 (N_4062,In_661,In_870);
and U4063 (N_4063,In_610,In_1792);
and U4064 (N_4064,In_1523,In_83);
nand U4065 (N_4065,In_505,In_1943);
or U4066 (N_4066,In_1691,In_1001);
nor U4067 (N_4067,In_1575,In_729);
nand U4068 (N_4068,In_1341,In_1226);
nor U4069 (N_4069,In_513,In_1667);
or U4070 (N_4070,In_1316,In_815);
nand U4071 (N_4071,In_1799,In_11);
nand U4072 (N_4072,In_19,In_1818);
nand U4073 (N_4073,In_1505,In_914);
nand U4074 (N_4074,In_1841,In_1820);
and U4075 (N_4075,In_842,In_1349);
xnor U4076 (N_4076,In_1922,In_346);
and U4077 (N_4077,In_79,In_1665);
and U4078 (N_4078,In_542,In_1397);
nor U4079 (N_4079,In_542,In_442);
and U4080 (N_4080,In_1810,In_1724);
and U4081 (N_4081,In_411,In_527);
nor U4082 (N_4082,In_128,In_1856);
and U4083 (N_4083,In_1069,In_1499);
and U4084 (N_4084,In_284,In_1505);
nor U4085 (N_4085,In_873,In_842);
nand U4086 (N_4086,In_1351,In_438);
and U4087 (N_4087,In_157,In_1374);
or U4088 (N_4088,In_623,In_1004);
nor U4089 (N_4089,In_432,In_1049);
and U4090 (N_4090,In_1253,In_821);
xnor U4091 (N_4091,In_1411,In_60);
nor U4092 (N_4092,In_845,In_1580);
nor U4093 (N_4093,In_1919,In_30);
nand U4094 (N_4094,In_1251,In_1814);
or U4095 (N_4095,In_834,In_88);
nor U4096 (N_4096,In_20,In_495);
and U4097 (N_4097,In_952,In_664);
nand U4098 (N_4098,In_1201,In_1016);
nand U4099 (N_4099,In_91,In_1466);
or U4100 (N_4100,In_1499,In_1177);
nand U4101 (N_4101,In_975,In_1216);
nand U4102 (N_4102,In_1120,In_1830);
or U4103 (N_4103,In_1823,In_440);
and U4104 (N_4104,In_495,In_1104);
nand U4105 (N_4105,In_420,In_1558);
nor U4106 (N_4106,In_1227,In_615);
nand U4107 (N_4107,In_365,In_762);
and U4108 (N_4108,In_991,In_288);
xor U4109 (N_4109,In_1960,In_551);
and U4110 (N_4110,In_1629,In_293);
nand U4111 (N_4111,In_1163,In_1919);
nor U4112 (N_4112,In_1123,In_465);
nor U4113 (N_4113,In_533,In_69);
xor U4114 (N_4114,In_1668,In_1303);
nor U4115 (N_4115,In_882,In_1037);
and U4116 (N_4116,In_1476,In_1059);
and U4117 (N_4117,In_1243,In_1963);
nor U4118 (N_4118,In_1129,In_1657);
and U4119 (N_4119,In_312,In_1229);
nand U4120 (N_4120,In_1011,In_74);
or U4121 (N_4121,In_1825,In_483);
nand U4122 (N_4122,In_763,In_1585);
nor U4123 (N_4123,In_938,In_922);
xor U4124 (N_4124,In_1623,In_1891);
or U4125 (N_4125,In_972,In_38);
and U4126 (N_4126,In_51,In_1403);
nand U4127 (N_4127,In_820,In_678);
nor U4128 (N_4128,In_788,In_712);
and U4129 (N_4129,In_1203,In_689);
nand U4130 (N_4130,In_1862,In_1675);
nor U4131 (N_4131,In_696,In_398);
xnor U4132 (N_4132,In_182,In_1379);
nor U4133 (N_4133,In_1817,In_1009);
and U4134 (N_4134,In_990,In_1676);
and U4135 (N_4135,In_530,In_463);
or U4136 (N_4136,In_1308,In_1697);
xnor U4137 (N_4137,In_42,In_1699);
nand U4138 (N_4138,In_318,In_54);
or U4139 (N_4139,In_1820,In_662);
nor U4140 (N_4140,In_456,In_1004);
nand U4141 (N_4141,In_163,In_652);
nor U4142 (N_4142,In_819,In_451);
nor U4143 (N_4143,In_494,In_355);
nand U4144 (N_4144,In_1554,In_618);
nor U4145 (N_4145,In_816,In_946);
nand U4146 (N_4146,In_1464,In_870);
xnor U4147 (N_4147,In_26,In_1354);
xnor U4148 (N_4148,In_617,In_733);
or U4149 (N_4149,In_32,In_1574);
nor U4150 (N_4150,In_1818,In_1175);
xnor U4151 (N_4151,In_368,In_776);
and U4152 (N_4152,In_938,In_150);
nor U4153 (N_4153,In_1453,In_1677);
nor U4154 (N_4154,In_290,In_1624);
nand U4155 (N_4155,In_1784,In_1701);
xor U4156 (N_4156,In_464,In_286);
and U4157 (N_4157,In_269,In_1439);
nand U4158 (N_4158,In_201,In_1730);
nand U4159 (N_4159,In_99,In_882);
nor U4160 (N_4160,In_935,In_308);
nor U4161 (N_4161,In_1812,In_1653);
or U4162 (N_4162,In_221,In_462);
nor U4163 (N_4163,In_1686,In_1588);
or U4164 (N_4164,In_1480,In_1300);
xor U4165 (N_4165,In_367,In_1306);
or U4166 (N_4166,In_1692,In_902);
xnor U4167 (N_4167,In_1260,In_1736);
and U4168 (N_4168,In_1532,In_1560);
xnor U4169 (N_4169,In_1423,In_1038);
and U4170 (N_4170,In_153,In_375);
nand U4171 (N_4171,In_632,In_1957);
nor U4172 (N_4172,In_931,In_1063);
nand U4173 (N_4173,In_1946,In_1402);
and U4174 (N_4174,In_807,In_859);
xnor U4175 (N_4175,In_224,In_442);
nand U4176 (N_4176,In_942,In_1146);
and U4177 (N_4177,In_1969,In_1609);
nand U4178 (N_4178,In_1085,In_633);
nor U4179 (N_4179,In_1118,In_833);
xor U4180 (N_4180,In_541,In_65);
nor U4181 (N_4181,In_819,In_1963);
xor U4182 (N_4182,In_784,In_1050);
nand U4183 (N_4183,In_509,In_282);
and U4184 (N_4184,In_965,In_1694);
xnor U4185 (N_4185,In_1548,In_1787);
or U4186 (N_4186,In_629,In_1604);
xor U4187 (N_4187,In_425,In_807);
and U4188 (N_4188,In_1005,In_235);
and U4189 (N_4189,In_257,In_1075);
or U4190 (N_4190,In_1373,In_266);
nor U4191 (N_4191,In_1031,In_1464);
xnor U4192 (N_4192,In_424,In_1841);
nor U4193 (N_4193,In_699,In_284);
or U4194 (N_4194,In_748,In_1824);
xnor U4195 (N_4195,In_1944,In_59);
and U4196 (N_4196,In_879,In_1255);
or U4197 (N_4197,In_1281,In_603);
and U4198 (N_4198,In_1034,In_1774);
nor U4199 (N_4199,In_1427,In_1438);
nand U4200 (N_4200,In_1774,In_1621);
or U4201 (N_4201,In_217,In_12);
or U4202 (N_4202,In_1904,In_1241);
or U4203 (N_4203,In_896,In_1551);
or U4204 (N_4204,In_1281,In_761);
or U4205 (N_4205,In_1318,In_261);
nand U4206 (N_4206,In_1864,In_417);
and U4207 (N_4207,In_1238,In_450);
nand U4208 (N_4208,In_971,In_1765);
xnor U4209 (N_4209,In_813,In_1661);
and U4210 (N_4210,In_1629,In_540);
nor U4211 (N_4211,In_1295,In_1384);
nand U4212 (N_4212,In_1567,In_727);
and U4213 (N_4213,In_1085,In_433);
and U4214 (N_4214,In_380,In_1024);
xnor U4215 (N_4215,In_1567,In_779);
nor U4216 (N_4216,In_543,In_1264);
or U4217 (N_4217,In_1752,In_716);
and U4218 (N_4218,In_1255,In_340);
and U4219 (N_4219,In_111,In_546);
nand U4220 (N_4220,In_925,In_116);
nand U4221 (N_4221,In_632,In_906);
or U4222 (N_4222,In_444,In_1265);
or U4223 (N_4223,In_1373,In_1732);
or U4224 (N_4224,In_731,In_1595);
nor U4225 (N_4225,In_1381,In_1916);
and U4226 (N_4226,In_1766,In_1219);
or U4227 (N_4227,In_649,In_1482);
or U4228 (N_4228,In_884,In_1006);
and U4229 (N_4229,In_1866,In_1795);
or U4230 (N_4230,In_1990,In_1860);
nor U4231 (N_4231,In_1464,In_1917);
and U4232 (N_4232,In_1726,In_998);
nor U4233 (N_4233,In_12,In_132);
nand U4234 (N_4234,In_1662,In_1679);
and U4235 (N_4235,In_1829,In_517);
nand U4236 (N_4236,In_1747,In_1484);
or U4237 (N_4237,In_233,In_1898);
or U4238 (N_4238,In_502,In_541);
and U4239 (N_4239,In_1158,In_1493);
or U4240 (N_4240,In_1037,In_447);
or U4241 (N_4241,In_249,In_1197);
xor U4242 (N_4242,In_1477,In_416);
nor U4243 (N_4243,In_936,In_1204);
or U4244 (N_4244,In_726,In_1147);
and U4245 (N_4245,In_1465,In_1327);
xnor U4246 (N_4246,In_1718,In_1494);
and U4247 (N_4247,In_453,In_1281);
xor U4248 (N_4248,In_1635,In_1814);
nor U4249 (N_4249,In_650,In_206);
nand U4250 (N_4250,In_442,In_79);
and U4251 (N_4251,In_1043,In_1624);
or U4252 (N_4252,In_6,In_1866);
or U4253 (N_4253,In_758,In_837);
or U4254 (N_4254,In_1333,In_569);
nand U4255 (N_4255,In_1176,In_27);
or U4256 (N_4256,In_354,In_251);
or U4257 (N_4257,In_1106,In_1019);
xor U4258 (N_4258,In_571,In_953);
or U4259 (N_4259,In_215,In_657);
or U4260 (N_4260,In_102,In_1527);
and U4261 (N_4261,In_236,In_1169);
nand U4262 (N_4262,In_966,In_1840);
nand U4263 (N_4263,In_933,In_1685);
xor U4264 (N_4264,In_892,In_1911);
nand U4265 (N_4265,In_202,In_414);
xor U4266 (N_4266,In_117,In_1661);
and U4267 (N_4267,In_222,In_1677);
xor U4268 (N_4268,In_1942,In_1375);
xnor U4269 (N_4269,In_882,In_1623);
xnor U4270 (N_4270,In_1303,In_1147);
or U4271 (N_4271,In_1319,In_1988);
xnor U4272 (N_4272,In_476,In_1836);
and U4273 (N_4273,In_1102,In_713);
nand U4274 (N_4274,In_979,In_803);
xor U4275 (N_4275,In_749,In_1623);
nand U4276 (N_4276,In_1432,In_1852);
and U4277 (N_4277,In_757,In_366);
nand U4278 (N_4278,In_240,In_1711);
xnor U4279 (N_4279,In_1091,In_1861);
xnor U4280 (N_4280,In_41,In_28);
or U4281 (N_4281,In_362,In_1788);
and U4282 (N_4282,In_1742,In_395);
nor U4283 (N_4283,In_216,In_375);
nand U4284 (N_4284,In_384,In_1926);
or U4285 (N_4285,In_729,In_542);
xnor U4286 (N_4286,In_528,In_1649);
nand U4287 (N_4287,In_1472,In_1355);
nor U4288 (N_4288,In_1325,In_827);
xnor U4289 (N_4289,In_1934,In_1804);
or U4290 (N_4290,In_1649,In_1428);
and U4291 (N_4291,In_348,In_717);
or U4292 (N_4292,In_1990,In_1868);
xnor U4293 (N_4293,In_1696,In_294);
or U4294 (N_4294,In_1983,In_1890);
or U4295 (N_4295,In_1700,In_957);
or U4296 (N_4296,In_1504,In_509);
or U4297 (N_4297,In_1773,In_1280);
and U4298 (N_4298,In_458,In_1220);
and U4299 (N_4299,In_1968,In_1232);
nand U4300 (N_4300,In_250,In_1113);
and U4301 (N_4301,In_1430,In_1738);
nor U4302 (N_4302,In_1651,In_1036);
and U4303 (N_4303,In_694,In_490);
xor U4304 (N_4304,In_1043,In_1332);
and U4305 (N_4305,In_1697,In_686);
nand U4306 (N_4306,In_1486,In_163);
xnor U4307 (N_4307,In_1634,In_678);
nor U4308 (N_4308,In_1996,In_1019);
nand U4309 (N_4309,In_693,In_1366);
or U4310 (N_4310,In_186,In_330);
nor U4311 (N_4311,In_1525,In_1750);
and U4312 (N_4312,In_1461,In_544);
nor U4313 (N_4313,In_1818,In_1145);
or U4314 (N_4314,In_242,In_155);
xor U4315 (N_4315,In_703,In_828);
xnor U4316 (N_4316,In_836,In_182);
or U4317 (N_4317,In_417,In_1352);
nor U4318 (N_4318,In_1173,In_1322);
nor U4319 (N_4319,In_854,In_337);
xnor U4320 (N_4320,In_1048,In_1111);
xnor U4321 (N_4321,In_1655,In_1219);
or U4322 (N_4322,In_1201,In_1319);
or U4323 (N_4323,In_1738,In_223);
xor U4324 (N_4324,In_1948,In_1435);
nor U4325 (N_4325,In_1863,In_1415);
and U4326 (N_4326,In_927,In_1240);
xor U4327 (N_4327,In_990,In_561);
xor U4328 (N_4328,In_1472,In_564);
nand U4329 (N_4329,In_177,In_259);
nor U4330 (N_4330,In_1645,In_1627);
nand U4331 (N_4331,In_780,In_1664);
or U4332 (N_4332,In_182,In_1703);
nand U4333 (N_4333,In_1870,In_1474);
xnor U4334 (N_4334,In_1901,In_1235);
nor U4335 (N_4335,In_1355,In_1372);
and U4336 (N_4336,In_1770,In_1774);
and U4337 (N_4337,In_146,In_1877);
nand U4338 (N_4338,In_788,In_182);
or U4339 (N_4339,In_1823,In_1918);
nand U4340 (N_4340,In_692,In_1116);
nand U4341 (N_4341,In_1981,In_1136);
xnor U4342 (N_4342,In_104,In_614);
nand U4343 (N_4343,In_1563,In_1491);
and U4344 (N_4344,In_135,In_356);
nor U4345 (N_4345,In_310,In_841);
or U4346 (N_4346,In_988,In_1836);
nor U4347 (N_4347,In_1049,In_1614);
nor U4348 (N_4348,In_1630,In_1902);
xnor U4349 (N_4349,In_521,In_1227);
nand U4350 (N_4350,In_179,In_509);
nand U4351 (N_4351,In_942,In_1379);
xor U4352 (N_4352,In_868,In_1676);
or U4353 (N_4353,In_1905,In_1775);
nor U4354 (N_4354,In_1698,In_380);
and U4355 (N_4355,In_948,In_240);
nand U4356 (N_4356,In_766,In_248);
or U4357 (N_4357,In_409,In_145);
nand U4358 (N_4358,In_318,In_1115);
xor U4359 (N_4359,In_221,In_122);
or U4360 (N_4360,In_950,In_690);
xnor U4361 (N_4361,In_1642,In_114);
nand U4362 (N_4362,In_1859,In_534);
and U4363 (N_4363,In_197,In_941);
nor U4364 (N_4364,In_221,In_1228);
and U4365 (N_4365,In_761,In_369);
nor U4366 (N_4366,In_541,In_1726);
nand U4367 (N_4367,In_1294,In_1765);
xnor U4368 (N_4368,In_1983,In_677);
xnor U4369 (N_4369,In_1935,In_303);
xnor U4370 (N_4370,In_225,In_44);
nand U4371 (N_4371,In_1374,In_1163);
or U4372 (N_4372,In_358,In_369);
xor U4373 (N_4373,In_540,In_1768);
and U4374 (N_4374,In_797,In_1670);
and U4375 (N_4375,In_1618,In_156);
nand U4376 (N_4376,In_21,In_1957);
or U4377 (N_4377,In_445,In_1349);
and U4378 (N_4378,In_159,In_1547);
and U4379 (N_4379,In_1990,In_1156);
nor U4380 (N_4380,In_138,In_478);
nor U4381 (N_4381,In_1115,In_1428);
xnor U4382 (N_4382,In_563,In_362);
or U4383 (N_4383,In_310,In_1738);
nor U4384 (N_4384,In_1239,In_1576);
nand U4385 (N_4385,In_1750,In_60);
nand U4386 (N_4386,In_103,In_1610);
nor U4387 (N_4387,In_1196,In_1586);
xnor U4388 (N_4388,In_871,In_695);
xor U4389 (N_4389,In_1916,In_409);
nand U4390 (N_4390,In_104,In_1719);
xnor U4391 (N_4391,In_1599,In_455);
nor U4392 (N_4392,In_1548,In_860);
nor U4393 (N_4393,In_1929,In_1740);
and U4394 (N_4394,In_1913,In_933);
or U4395 (N_4395,In_780,In_631);
xor U4396 (N_4396,In_841,In_366);
or U4397 (N_4397,In_1977,In_50);
xor U4398 (N_4398,In_238,In_1431);
nand U4399 (N_4399,In_1955,In_1171);
nand U4400 (N_4400,In_662,In_856);
xor U4401 (N_4401,In_309,In_1020);
nand U4402 (N_4402,In_1959,In_1683);
and U4403 (N_4403,In_643,In_1560);
xor U4404 (N_4404,In_1425,In_189);
nor U4405 (N_4405,In_631,In_1891);
or U4406 (N_4406,In_747,In_908);
nand U4407 (N_4407,In_924,In_727);
or U4408 (N_4408,In_1226,In_1563);
and U4409 (N_4409,In_901,In_1763);
nand U4410 (N_4410,In_1027,In_762);
or U4411 (N_4411,In_222,In_1646);
nand U4412 (N_4412,In_1001,In_381);
and U4413 (N_4413,In_1842,In_1839);
and U4414 (N_4414,In_152,In_185);
nand U4415 (N_4415,In_688,In_1060);
and U4416 (N_4416,In_515,In_243);
nand U4417 (N_4417,In_387,In_271);
and U4418 (N_4418,In_478,In_954);
nand U4419 (N_4419,In_1199,In_43);
nor U4420 (N_4420,In_1799,In_405);
or U4421 (N_4421,In_1265,In_593);
xnor U4422 (N_4422,In_1485,In_752);
or U4423 (N_4423,In_1448,In_503);
and U4424 (N_4424,In_95,In_404);
nand U4425 (N_4425,In_911,In_1298);
nand U4426 (N_4426,In_1983,In_1880);
nand U4427 (N_4427,In_1751,In_603);
nand U4428 (N_4428,In_649,In_627);
xor U4429 (N_4429,In_1648,In_192);
and U4430 (N_4430,In_925,In_729);
nor U4431 (N_4431,In_313,In_412);
and U4432 (N_4432,In_234,In_1229);
nand U4433 (N_4433,In_268,In_147);
and U4434 (N_4434,In_1300,In_1439);
nor U4435 (N_4435,In_1411,In_1650);
nor U4436 (N_4436,In_302,In_538);
or U4437 (N_4437,In_640,In_978);
or U4438 (N_4438,In_1515,In_348);
xor U4439 (N_4439,In_1648,In_46);
nor U4440 (N_4440,In_17,In_665);
and U4441 (N_4441,In_201,In_1614);
and U4442 (N_4442,In_1033,In_1010);
nor U4443 (N_4443,In_896,In_844);
or U4444 (N_4444,In_1163,In_1051);
xor U4445 (N_4445,In_1026,In_100);
nor U4446 (N_4446,In_1213,In_1652);
nor U4447 (N_4447,In_114,In_490);
nand U4448 (N_4448,In_838,In_1272);
or U4449 (N_4449,In_1194,In_919);
or U4450 (N_4450,In_1173,In_1851);
nand U4451 (N_4451,In_957,In_1533);
xor U4452 (N_4452,In_116,In_664);
or U4453 (N_4453,In_907,In_1821);
and U4454 (N_4454,In_1002,In_426);
and U4455 (N_4455,In_1686,In_1955);
and U4456 (N_4456,In_1515,In_721);
nand U4457 (N_4457,In_610,In_115);
and U4458 (N_4458,In_1807,In_1554);
xor U4459 (N_4459,In_848,In_1394);
nand U4460 (N_4460,In_1747,In_903);
nor U4461 (N_4461,In_15,In_805);
and U4462 (N_4462,In_1178,In_1081);
nand U4463 (N_4463,In_418,In_527);
nor U4464 (N_4464,In_1552,In_713);
nand U4465 (N_4465,In_778,In_1254);
nor U4466 (N_4466,In_1217,In_298);
nor U4467 (N_4467,In_240,In_1005);
nand U4468 (N_4468,In_188,In_1151);
and U4469 (N_4469,In_866,In_1033);
and U4470 (N_4470,In_1326,In_261);
nor U4471 (N_4471,In_1306,In_1964);
nand U4472 (N_4472,In_588,In_1194);
or U4473 (N_4473,In_1726,In_1315);
or U4474 (N_4474,In_1638,In_815);
nor U4475 (N_4475,In_407,In_925);
nand U4476 (N_4476,In_1699,In_1059);
and U4477 (N_4477,In_524,In_332);
xor U4478 (N_4478,In_1563,In_1800);
nand U4479 (N_4479,In_184,In_173);
nor U4480 (N_4480,In_1777,In_1724);
xnor U4481 (N_4481,In_1246,In_1625);
or U4482 (N_4482,In_1328,In_1189);
nand U4483 (N_4483,In_799,In_1129);
or U4484 (N_4484,In_13,In_160);
nand U4485 (N_4485,In_336,In_1268);
and U4486 (N_4486,In_1910,In_1142);
and U4487 (N_4487,In_6,In_1734);
or U4488 (N_4488,In_1610,In_1303);
or U4489 (N_4489,In_468,In_1964);
nand U4490 (N_4490,In_1332,In_893);
xnor U4491 (N_4491,In_1223,In_212);
or U4492 (N_4492,In_613,In_649);
or U4493 (N_4493,In_1356,In_1958);
nor U4494 (N_4494,In_21,In_1877);
nand U4495 (N_4495,In_46,In_393);
nand U4496 (N_4496,In_933,In_782);
nand U4497 (N_4497,In_432,In_1310);
xnor U4498 (N_4498,In_661,In_1383);
or U4499 (N_4499,In_606,In_1180);
nor U4500 (N_4500,In_1201,In_1696);
or U4501 (N_4501,In_435,In_1193);
nand U4502 (N_4502,In_261,In_1660);
xnor U4503 (N_4503,In_851,In_1614);
or U4504 (N_4504,In_1271,In_1774);
or U4505 (N_4505,In_1144,In_248);
nor U4506 (N_4506,In_1650,In_696);
xor U4507 (N_4507,In_622,In_1920);
nand U4508 (N_4508,In_365,In_634);
and U4509 (N_4509,In_479,In_1679);
nand U4510 (N_4510,In_1213,In_137);
and U4511 (N_4511,In_234,In_625);
nor U4512 (N_4512,In_348,In_1787);
xnor U4513 (N_4513,In_1806,In_1476);
or U4514 (N_4514,In_427,In_1520);
or U4515 (N_4515,In_798,In_762);
and U4516 (N_4516,In_622,In_1938);
and U4517 (N_4517,In_815,In_354);
xor U4518 (N_4518,In_379,In_382);
or U4519 (N_4519,In_1997,In_555);
nor U4520 (N_4520,In_1108,In_1000);
nor U4521 (N_4521,In_968,In_201);
and U4522 (N_4522,In_5,In_277);
or U4523 (N_4523,In_1957,In_67);
nor U4524 (N_4524,In_1106,In_65);
nor U4525 (N_4525,In_1289,In_1215);
nand U4526 (N_4526,In_379,In_937);
nand U4527 (N_4527,In_1895,In_75);
nand U4528 (N_4528,In_1917,In_343);
nand U4529 (N_4529,In_52,In_230);
or U4530 (N_4530,In_14,In_615);
and U4531 (N_4531,In_1506,In_1256);
nand U4532 (N_4532,In_487,In_1326);
and U4533 (N_4533,In_1064,In_36);
nand U4534 (N_4534,In_1884,In_1616);
or U4535 (N_4535,In_409,In_714);
nor U4536 (N_4536,In_981,In_1462);
xnor U4537 (N_4537,In_194,In_1509);
nand U4538 (N_4538,In_1681,In_1479);
nand U4539 (N_4539,In_1746,In_370);
nand U4540 (N_4540,In_1408,In_82);
or U4541 (N_4541,In_1016,In_133);
and U4542 (N_4542,In_455,In_1881);
or U4543 (N_4543,In_13,In_167);
and U4544 (N_4544,In_1750,In_1785);
or U4545 (N_4545,In_750,In_1635);
nand U4546 (N_4546,In_985,In_1195);
nor U4547 (N_4547,In_1118,In_454);
and U4548 (N_4548,In_325,In_771);
nand U4549 (N_4549,In_1836,In_1443);
or U4550 (N_4550,In_489,In_281);
nand U4551 (N_4551,In_1381,In_35);
nor U4552 (N_4552,In_479,In_922);
or U4553 (N_4553,In_551,In_1442);
xnor U4554 (N_4554,In_1278,In_1027);
or U4555 (N_4555,In_1590,In_1191);
or U4556 (N_4556,In_1463,In_638);
and U4557 (N_4557,In_77,In_1909);
nand U4558 (N_4558,In_257,In_1378);
or U4559 (N_4559,In_345,In_1753);
xnor U4560 (N_4560,In_907,In_1379);
nand U4561 (N_4561,In_505,In_1617);
nor U4562 (N_4562,In_510,In_1347);
or U4563 (N_4563,In_1465,In_1003);
nor U4564 (N_4564,In_117,In_238);
and U4565 (N_4565,In_35,In_957);
nand U4566 (N_4566,In_1605,In_3);
or U4567 (N_4567,In_1006,In_922);
and U4568 (N_4568,In_1358,In_609);
xor U4569 (N_4569,In_1609,In_1417);
and U4570 (N_4570,In_1801,In_1715);
and U4571 (N_4571,In_290,In_1694);
xor U4572 (N_4572,In_417,In_1718);
and U4573 (N_4573,In_1876,In_1915);
xor U4574 (N_4574,In_1107,In_1258);
nor U4575 (N_4575,In_1883,In_1085);
nor U4576 (N_4576,In_493,In_749);
and U4577 (N_4577,In_468,In_144);
or U4578 (N_4578,In_518,In_83);
and U4579 (N_4579,In_601,In_481);
nand U4580 (N_4580,In_519,In_466);
and U4581 (N_4581,In_333,In_398);
nor U4582 (N_4582,In_207,In_392);
nand U4583 (N_4583,In_1543,In_608);
xor U4584 (N_4584,In_1480,In_1334);
and U4585 (N_4585,In_1219,In_180);
nor U4586 (N_4586,In_420,In_145);
and U4587 (N_4587,In_1920,In_320);
or U4588 (N_4588,In_489,In_907);
nand U4589 (N_4589,In_261,In_1343);
nor U4590 (N_4590,In_1131,In_482);
and U4591 (N_4591,In_63,In_807);
nor U4592 (N_4592,In_1978,In_105);
or U4593 (N_4593,In_1964,In_1327);
or U4594 (N_4594,In_1951,In_271);
or U4595 (N_4595,In_725,In_426);
or U4596 (N_4596,In_573,In_202);
nor U4597 (N_4597,In_313,In_167);
nand U4598 (N_4598,In_528,In_20);
nand U4599 (N_4599,In_1664,In_556);
or U4600 (N_4600,In_757,In_1131);
nand U4601 (N_4601,In_1532,In_1023);
xnor U4602 (N_4602,In_637,In_221);
or U4603 (N_4603,In_1332,In_1478);
xor U4604 (N_4604,In_517,In_259);
and U4605 (N_4605,In_1271,In_166);
and U4606 (N_4606,In_1856,In_1307);
or U4607 (N_4607,In_1059,In_1691);
and U4608 (N_4608,In_1584,In_895);
and U4609 (N_4609,In_1605,In_551);
xnor U4610 (N_4610,In_149,In_1940);
or U4611 (N_4611,In_74,In_100);
and U4612 (N_4612,In_321,In_1156);
nor U4613 (N_4613,In_1211,In_1610);
xnor U4614 (N_4614,In_128,In_1705);
nand U4615 (N_4615,In_1774,In_1640);
nand U4616 (N_4616,In_1436,In_1241);
nor U4617 (N_4617,In_437,In_1216);
nor U4618 (N_4618,In_1322,In_551);
nand U4619 (N_4619,In_1311,In_1055);
or U4620 (N_4620,In_124,In_747);
or U4621 (N_4621,In_363,In_969);
nor U4622 (N_4622,In_1046,In_652);
nor U4623 (N_4623,In_1193,In_1492);
and U4624 (N_4624,In_87,In_1508);
and U4625 (N_4625,In_228,In_1764);
xnor U4626 (N_4626,In_1919,In_586);
nand U4627 (N_4627,In_1647,In_52);
or U4628 (N_4628,In_820,In_1329);
or U4629 (N_4629,In_611,In_1103);
nor U4630 (N_4630,In_896,In_1869);
xor U4631 (N_4631,In_1380,In_301);
xor U4632 (N_4632,In_298,In_639);
or U4633 (N_4633,In_765,In_1769);
nand U4634 (N_4634,In_260,In_941);
nand U4635 (N_4635,In_1717,In_177);
and U4636 (N_4636,In_1628,In_709);
and U4637 (N_4637,In_1638,In_307);
nor U4638 (N_4638,In_1691,In_148);
xor U4639 (N_4639,In_1793,In_1390);
or U4640 (N_4640,In_15,In_1783);
or U4641 (N_4641,In_1004,In_1499);
or U4642 (N_4642,In_222,In_304);
and U4643 (N_4643,In_1495,In_1118);
or U4644 (N_4644,In_1158,In_1556);
nor U4645 (N_4645,In_1413,In_80);
and U4646 (N_4646,In_1676,In_992);
xor U4647 (N_4647,In_1131,In_1067);
or U4648 (N_4648,In_1351,In_758);
nand U4649 (N_4649,In_1196,In_1972);
and U4650 (N_4650,In_1248,In_1091);
and U4651 (N_4651,In_1170,In_70);
or U4652 (N_4652,In_1061,In_1313);
nand U4653 (N_4653,In_1120,In_1259);
nand U4654 (N_4654,In_1759,In_1384);
or U4655 (N_4655,In_1379,In_1571);
nor U4656 (N_4656,In_1991,In_1734);
nand U4657 (N_4657,In_146,In_498);
nor U4658 (N_4658,In_1817,In_1258);
or U4659 (N_4659,In_538,In_1808);
xnor U4660 (N_4660,In_389,In_305);
nor U4661 (N_4661,In_385,In_561);
and U4662 (N_4662,In_467,In_66);
xnor U4663 (N_4663,In_1128,In_847);
and U4664 (N_4664,In_1758,In_665);
nand U4665 (N_4665,In_51,In_1508);
nand U4666 (N_4666,In_1516,In_1580);
nand U4667 (N_4667,In_826,In_190);
xor U4668 (N_4668,In_1614,In_267);
nor U4669 (N_4669,In_553,In_623);
and U4670 (N_4670,In_1075,In_128);
xor U4671 (N_4671,In_1312,In_413);
nand U4672 (N_4672,In_1602,In_1397);
or U4673 (N_4673,In_1032,In_327);
nand U4674 (N_4674,In_391,In_916);
nand U4675 (N_4675,In_1101,In_1551);
nand U4676 (N_4676,In_1663,In_1232);
xnor U4677 (N_4677,In_108,In_473);
and U4678 (N_4678,In_1330,In_1008);
or U4679 (N_4679,In_667,In_1038);
nor U4680 (N_4680,In_1376,In_1927);
nand U4681 (N_4681,In_1443,In_381);
nor U4682 (N_4682,In_730,In_633);
and U4683 (N_4683,In_557,In_1365);
nor U4684 (N_4684,In_810,In_530);
nor U4685 (N_4685,In_1846,In_473);
nor U4686 (N_4686,In_492,In_273);
xor U4687 (N_4687,In_1344,In_846);
and U4688 (N_4688,In_288,In_1359);
and U4689 (N_4689,In_1150,In_1627);
xor U4690 (N_4690,In_122,In_744);
xor U4691 (N_4691,In_155,In_129);
nor U4692 (N_4692,In_1275,In_68);
nor U4693 (N_4693,In_1190,In_1596);
xnor U4694 (N_4694,In_1594,In_797);
nor U4695 (N_4695,In_134,In_794);
nand U4696 (N_4696,In_628,In_1244);
nand U4697 (N_4697,In_1704,In_197);
nor U4698 (N_4698,In_463,In_174);
nor U4699 (N_4699,In_1539,In_1848);
and U4700 (N_4700,In_804,In_880);
or U4701 (N_4701,In_1589,In_1951);
nand U4702 (N_4702,In_253,In_1120);
or U4703 (N_4703,In_1962,In_1705);
or U4704 (N_4704,In_58,In_1258);
and U4705 (N_4705,In_893,In_1611);
xor U4706 (N_4706,In_1966,In_1912);
nand U4707 (N_4707,In_1904,In_1967);
nor U4708 (N_4708,In_1015,In_1386);
nand U4709 (N_4709,In_1442,In_881);
or U4710 (N_4710,In_1494,In_1045);
and U4711 (N_4711,In_1539,In_1673);
xor U4712 (N_4712,In_1771,In_1497);
xor U4713 (N_4713,In_753,In_1737);
nand U4714 (N_4714,In_1908,In_1367);
xor U4715 (N_4715,In_667,In_1394);
nor U4716 (N_4716,In_1099,In_300);
and U4717 (N_4717,In_896,In_826);
nor U4718 (N_4718,In_1955,In_1229);
nand U4719 (N_4719,In_350,In_1067);
and U4720 (N_4720,In_1324,In_1607);
and U4721 (N_4721,In_918,In_1173);
xnor U4722 (N_4722,In_434,In_1323);
or U4723 (N_4723,In_592,In_1218);
or U4724 (N_4724,In_381,In_1412);
xnor U4725 (N_4725,In_810,In_665);
and U4726 (N_4726,In_319,In_337);
nor U4727 (N_4727,In_573,In_338);
nor U4728 (N_4728,In_1519,In_487);
nor U4729 (N_4729,In_490,In_1667);
nor U4730 (N_4730,In_207,In_1967);
nand U4731 (N_4731,In_1101,In_1067);
and U4732 (N_4732,In_670,In_1650);
xor U4733 (N_4733,In_512,In_1575);
nand U4734 (N_4734,In_1573,In_1745);
nand U4735 (N_4735,In_867,In_1685);
xor U4736 (N_4736,In_1420,In_1787);
nor U4737 (N_4737,In_924,In_1357);
or U4738 (N_4738,In_1722,In_834);
nand U4739 (N_4739,In_597,In_1839);
xnor U4740 (N_4740,In_210,In_1017);
nor U4741 (N_4741,In_1917,In_687);
nand U4742 (N_4742,In_801,In_1396);
and U4743 (N_4743,In_174,In_1510);
or U4744 (N_4744,In_208,In_1443);
xnor U4745 (N_4745,In_981,In_1835);
nor U4746 (N_4746,In_136,In_1855);
and U4747 (N_4747,In_1030,In_239);
xnor U4748 (N_4748,In_1603,In_1175);
or U4749 (N_4749,In_752,In_1143);
xnor U4750 (N_4750,In_1841,In_284);
nor U4751 (N_4751,In_31,In_1781);
or U4752 (N_4752,In_1931,In_1297);
and U4753 (N_4753,In_499,In_1609);
or U4754 (N_4754,In_1706,In_258);
and U4755 (N_4755,In_1747,In_597);
nor U4756 (N_4756,In_36,In_788);
and U4757 (N_4757,In_1162,In_1330);
nand U4758 (N_4758,In_1818,In_118);
xnor U4759 (N_4759,In_965,In_919);
or U4760 (N_4760,In_1878,In_490);
or U4761 (N_4761,In_767,In_209);
nor U4762 (N_4762,In_197,In_1425);
nand U4763 (N_4763,In_1170,In_129);
and U4764 (N_4764,In_1405,In_1035);
and U4765 (N_4765,In_1662,In_1543);
nand U4766 (N_4766,In_1699,In_1616);
nand U4767 (N_4767,In_917,In_1505);
nor U4768 (N_4768,In_1434,In_1574);
nand U4769 (N_4769,In_948,In_1474);
nand U4770 (N_4770,In_1969,In_175);
and U4771 (N_4771,In_1438,In_715);
and U4772 (N_4772,In_1263,In_1861);
nand U4773 (N_4773,In_1381,In_1378);
nor U4774 (N_4774,In_111,In_169);
xor U4775 (N_4775,In_912,In_925);
or U4776 (N_4776,In_967,In_461);
and U4777 (N_4777,In_1702,In_1638);
and U4778 (N_4778,In_901,In_1150);
or U4779 (N_4779,In_1730,In_1539);
nor U4780 (N_4780,In_355,In_1822);
and U4781 (N_4781,In_1104,In_398);
nor U4782 (N_4782,In_710,In_1813);
nand U4783 (N_4783,In_567,In_1894);
and U4784 (N_4784,In_1895,In_967);
nor U4785 (N_4785,In_1462,In_703);
nand U4786 (N_4786,In_821,In_1618);
and U4787 (N_4787,In_1024,In_1134);
or U4788 (N_4788,In_117,In_1173);
or U4789 (N_4789,In_48,In_1160);
and U4790 (N_4790,In_1992,In_611);
or U4791 (N_4791,In_1201,In_40);
and U4792 (N_4792,In_191,In_614);
and U4793 (N_4793,In_1095,In_400);
nand U4794 (N_4794,In_1052,In_1065);
and U4795 (N_4795,In_1728,In_1966);
nor U4796 (N_4796,In_1878,In_591);
and U4797 (N_4797,In_820,In_921);
nand U4798 (N_4798,In_1247,In_1820);
nor U4799 (N_4799,In_1803,In_1213);
and U4800 (N_4800,In_1717,In_1426);
or U4801 (N_4801,In_44,In_1473);
and U4802 (N_4802,In_62,In_1933);
xnor U4803 (N_4803,In_497,In_483);
xnor U4804 (N_4804,In_88,In_1153);
xor U4805 (N_4805,In_1037,In_557);
and U4806 (N_4806,In_1812,In_1573);
xor U4807 (N_4807,In_354,In_301);
or U4808 (N_4808,In_1261,In_1846);
or U4809 (N_4809,In_724,In_46);
and U4810 (N_4810,In_1885,In_339);
nor U4811 (N_4811,In_813,In_1432);
nand U4812 (N_4812,In_1983,In_1836);
nand U4813 (N_4813,In_235,In_1254);
and U4814 (N_4814,In_1365,In_483);
or U4815 (N_4815,In_1165,In_806);
and U4816 (N_4816,In_826,In_913);
or U4817 (N_4817,In_899,In_175);
nand U4818 (N_4818,In_199,In_194);
nor U4819 (N_4819,In_1676,In_1875);
xnor U4820 (N_4820,In_556,In_568);
or U4821 (N_4821,In_867,In_1275);
nor U4822 (N_4822,In_1247,In_273);
nor U4823 (N_4823,In_879,In_133);
xnor U4824 (N_4824,In_1894,In_582);
nand U4825 (N_4825,In_328,In_647);
nand U4826 (N_4826,In_105,In_128);
and U4827 (N_4827,In_1779,In_1436);
nor U4828 (N_4828,In_1693,In_529);
or U4829 (N_4829,In_1214,In_1642);
nand U4830 (N_4830,In_1886,In_1847);
xor U4831 (N_4831,In_120,In_308);
nand U4832 (N_4832,In_941,In_227);
nor U4833 (N_4833,In_433,In_1932);
xnor U4834 (N_4834,In_108,In_757);
and U4835 (N_4835,In_200,In_1287);
or U4836 (N_4836,In_257,In_602);
xnor U4837 (N_4837,In_1375,In_292);
nor U4838 (N_4838,In_478,In_1010);
or U4839 (N_4839,In_128,In_87);
nor U4840 (N_4840,In_1861,In_502);
nand U4841 (N_4841,In_1702,In_370);
nand U4842 (N_4842,In_1177,In_1964);
nand U4843 (N_4843,In_1340,In_892);
and U4844 (N_4844,In_1491,In_957);
and U4845 (N_4845,In_287,In_1645);
xor U4846 (N_4846,In_956,In_1808);
nand U4847 (N_4847,In_1833,In_798);
and U4848 (N_4848,In_985,In_1615);
nand U4849 (N_4849,In_1701,In_1176);
nor U4850 (N_4850,In_1093,In_544);
nand U4851 (N_4851,In_258,In_1438);
xor U4852 (N_4852,In_220,In_20);
and U4853 (N_4853,In_1253,In_1207);
nor U4854 (N_4854,In_683,In_540);
and U4855 (N_4855,In_12,In_332);
nand U4856 (N_4856,In_1815,In_1482);
nand U4857 (N_4857,In_1061,In_1519);
nand U4858 (N_4858,In_1055,In_1096);
and U4859 (N_4859,In_1802,In_1937);
and U4860 (N_4860,In_1638,In_1312);
nand U4861 (N_4861,In_1595,In_1768);
or U4862 (N_4862,In_506,In_1038);
nand U4863 (N_4863,In_1826,In_1201);
and U4864 (N_4864,In_110,In_785);
nand U4865 (N_4865,In_475,In_495);
nand U4866 (N_4866,In_1205,In_1405);
or U4867 (N_4867,In_1602,In_441);
xnor U4868 (N_4868,In_859,In_633);
nand U4869 (N_4869,In_1937,In_889);
xor U4870 (N_4870,In_545,In_1240);
and U4871 (N_4871,In_1176,In_493);
nor U4872 (N_4872,In_1266,In_1592);
and U4873 (N_4873,In_1974,In_130);
or U4874 (N_4874,In_1614,In_1909);
xnor U4875 (N_4875,In_757,In_1246);
nand U4876 (N_4876,In_565,In_1405);
and U4877 (N_4877,In_1364,In_382);
xnor U4878 (N_4878,In_626,In_1029);
xor U4879 (N_4879,In_1429,In_1542);
xnor U4880 (N_4880,In_1460,In_1433);
nor U4881 (N_4881,In_438,In_1314);
nand U4882 (N_4882,In_581,In_758);
nor U4883 (N_4883,In_1771,In_588);
xor U4884 (N_4884,In_606,In_1488);
nand U4885 (N_4885,In_1812,In_344);
and U4886 (N_4886,In_1066,In_1941);
or U4887 (N_4887,In_1886,In_1993);
and U4888 (N_4888,In_256,In_780);
nor U4889 (N_4889,In_450,In_1232);
nand U4890 (N_4890,In_1032,In_1357);
xor U4891 (N_4891,In_1618,In_1301);
or U4892 (N_4892,In_1809,In_1461);
xor U4893 (N_4893,In_1512,In_854);
xnor U4894 (N_4894,In_697,In_1955);
or U4895 (N_4895,In_1922,In_325);
and U4896 (N_4896,In_1340,In_1612);
and U4897 (N_4897,In_1980,In_1449);
nand U4898 (N_4898,In_1645,In_744);
nand U4899 (N_4899,In_1379,In_331);
and U4900 (N_4900,In_1682,In_1547);
and U4901 (N_4901,In_1878,In_1939);
nor U4902 (N_4902,In_997,In_1874);
nor U4903 (N_4903,In_1374,In_1002);
xor U4904 (N_4904,In_632,In_71);
and U4905 (N_4905,In_1893,In_1534);
xnor U4906 (N_4906,In_1851,In_1373);
or U4907 (N_4907,In_806,In_448);
or U4908 (N_4908,In_1860,In_1940);
or U4909 (N_4909,In_371,In_1627);
nor U4910 (N_4910,In_381,In_1420);
and U4911 (N_4911,In_1947,In_917);
or U4912 (N_4912,In_884,In_1216);
xnor U4913 (N_4913,In_1844,In_1895);
nand U4914 (N_4914,In_898,In_990);
and U4915 (N_4915,In_227,In_1757);
or U4916 (N_4916,In_1460,In_1826);
or U4917 (N_4917,In_1261,In_581);
xor U4918 (N_4918,In_630,In_376);
and U4919 (N_4919,In_1542,In_1834);
nand U4920 (N_4920,In_923,In_841);
nand U4921 (N_4921,In_1168,In_1767);
nand U4922 (N_4922,In_1463,In_1977);
and U4923 (N_4923,In_1135,In_939);
or U4924 (N_4924,In_385,In_1409);
nor U4925 (N_4925,In_405,In_1241);
nor U4926 (N_4926,In_172,In_576);
xor U4927 (N_4927,In_59,In_456);
nand U4928 (N_4928,In_1021,In_903);
nand U4929 (N_4929,In_233,In_1206);
and U4930 (N_4930,In_1368,In_1177);
and U4931 (N_4931,In_1560,In_1205);
or U4932 (N_4932,In_165,In_1371);
nor U4933 (N_4933,In_1575,In_488);
xnor U4934 (N_4934,In_1707,In_1392);
nor U4935 (N_4935,In_988,In_657);
and U4936 (N_4936,In_1764,In_1183);
nand U4937 (N_4937,In_1406,In_872);
nor U4938 (N_4938,In_541,In_820);
or U4939 (N_4939,In_1220,In_314);
or U4940 (N_4940,In_1931,In_723);
and U4941 (N_4941,In_1708,In_262);
nand U4942 (N_4942,In_317,In_1021);
nor U4943 (N_4943,In_1783,In_1319);
nor U4944 (N_4944,In_1485,In_1674);
nand U4945 (N_4945,In_70,In_1252);
xnor U4946 (N_4946,In_473,In_370);
and U4947 (N_4947,In_583,In_739);
nand U4948 (N_4948,In_253,In_1698);
or U4949 (N_4949,In_157,In_1304);
xnor U4950 (N_4950,In_1992,In_49);
nand U4951 (N_4951,In_596,In_1989);
xnor U4952 (N_4952,In_1663,In_1990);
nor U4953 (N_4953,In_1272,In_1655);
and U4954 (N_4954,In_1875,In_139);
nor U4955 (N_4955,In_1855,In_1798);
nand U4956 (N_4956,In_1192,In_971);
xnor U4957 (N_4957,In_789,In_1972);
and U4958 (N_4958,In_20,In_1693);
or U4959 (N_4959,In_1145,In_220);
xor U4960 (N_4960,In_511,In_1457);
or U4961 (N_4961,In_1904,In_1613);
nor U4962 (N_4962,In_17,In_1981);
nor U4963 (N_4963,In_1184,In_743);
xor U4964 (N_4964,In_1472,In_1198);
nor U4965 (N_4965,In_1388,In_75);
xor U4966 (N_4966,In_1106,In_184);
or U4967 (N_4967,In_447,In_1724);
or U4968 (N_4968,In_1259,In_461);
xor U4969 (N_4969,In_1166,In_360);
and U4970 (N_4970,In_1367,In_1233);
and U4971 (N_4971,In_228,In_1985);
nand U4972 (N_4972,In_690,In_1943);
or U4973 (N_4973,In_303,In_783);
nand U4974 (N_4974,In_983,In_1275);
nand U4975 (N_4975,In_1940,In_1685);
nor U4976 (N_4976,In_840,In_1761);
or U4977 (N_4977,In_1952,In_1992);
and U4978 (N_4978,In_651,In_1159);
nor U4979 (N_4979,In_640,In_1556);
xnor U4980 (N_4980,In_1194,In_265);
nor U4981 (N_4981,In_589,In_1766);
nor U4982 (N_4982,In_173,In_1339);
nor U4983 (N_4983,In_415,In_1123);
xnor U4984 (N_4984,In_589,In_1659);
or U4985 (N_4985,In_1132,In_1896);
and U4986 (N_4986,In_1608,In_1806);
and U4987 (N_4987,In_836,In_1314);
xnor U4988 (N_4988,In_1986,In_149);
xnor U4989 (N_4989,In_16,In_248);
or U4990 (N_4990,In_1169,In_1528);
nor U4991 (N_4991,In_817,In_428);
xnor U4992 (N_4992,In_1571,In_662);
and U4993 (N_4993,In_1590,In_1562);
xor U4994 (N_4994,In_696,In_919);
xor U4995 (N_4995,In_489,In_1344);
nor U4996 (N_4996,In_1465,In_1645);
xnor U4997 (N_4997,In_925,In_807);
and U4998 (N_4998,In_1654,In_1774);
xor U4999 (N_4999,In_1773,In_378);
nand U5000 (N_5000,N_3180,N_3812);
and U5001 (N_5001,N_4901,N_4700);
or U5002 (N_5002,N_1239,N_3298);
nand U5003 (N_5003,N_560,N_1642);
nor U5004 (N_5004,N_2344,N_2783);
and U5005 (N_5005,N_4244,N_999);
and U5006 (N_5006,N_2802,N_2464);
nand U5007 (N_5007,N_3316,N_2608);
nor U5008 (N_5008,N_4705,N_3669);
and U5009 (N_5009,N_3544,N_1934);
xnor U5010 (N_5010,N_2226,N_356);
nand U5011 (N_5011,N_4608,N_4589);
nand U5012 (N_5012,N_4259,N_557);
nor U5013 (N_5013,N_2441,N_1389);
xnor U5014 (N_5014,N_4504,N_2716);
or U5015 (N_5015,N_1852,N_1218);
nand U5016 (N_5016,N_2057,N_1092);
and U5017 (N_5017,N_62,N_4405);
nand U5018 (N_5018,N_2805,N_1390);
nor U5019 (N_5019,N_4737,N_2247);
and U5020 (N_5020,N_124,N_706);
nand U5021 (N_5021,N_988,N_1974);
nor U5022 (N_5022,N_2378,N_3557);
nand U5023 (N_5023,N_3330,N_4824);
nor U5024 (N_5024,N_1299,N_3276);
nor U5025 (N_5025,N_2941,N_4751);
nand U5026 (N_5026,N_579,N_1941);
nand U5027 (N_5027,N_738,N_4435);
or U5028 (N_5028,N_4595,N_3204);
xor U5029 (N_5029,N_4518,N_187);
and U5030 (N_5030,N_1855,N_928);
or U5031 (N_5031,N_3525,N_2040);
or U5032 (N_5032,N_2328,N_1319);
or U5033 (N_5033,N_632,N_3810);
or U5034 (N_5034,N_1771,N_571);
and U5035 (N_5035,N_2159,N_3289);
nor U5036 (N_5036,N_2370,N_325);
and U5037 (N_5037,N_2277,N_1494);
xor U5038 (N_5038,N_2412,N_1425);
and U5039 (N_5039,N_4640,N_2659);
nand U5040 (N_5040,N_4269,N_1577);
xor U5041 (N_5041,N_4159,N_118);
or U5042 (N_5042,N_2272,N_1654);
xor U5043 (N_5043,N_1625,N_2036);
and U5044 (N_5044,N_2278,N_2947);
or U5045 (N_5045,N_2512,N_3621);
xor U5046 (N_5046,N_3697,N_3719);
nand U5047 (N_5047,N_1436,N_1076);
nand U5048 (N_5048,N_4695,N_610);
and U5049 (N_5049,N_3869,N_1265);
and U5050 (N_5050,N_1268,N_3964);
nand U5051 (N_5051,N_1809,N_2393);
or U5052 (N_5052,N_3391,N_4508);
nand U5053 (N_5053,N_2055,N_1971);
or U5054 (N_5054,N_4457,N_3256);
or U5055 (N_5055,N_4452,N_1854);
nand U5056 (N_5056,N_2688,N_2538);
and U5057 (N_5057,N_2715,N_722);
nor U5058 (N_5058,N_3124,N_4060);
or U5059 (N_5059,N_626,N_2958);
or U5060 (N_5060,N_2406,N_635);
nor U5061 (N_5061,N_3566,N_755);
nand U5062 (N_5062,N_530,N_574);
and U5063 (N_5063,N_354,N_4618);
and U5064 (N_5064,N_3632,N_64);
nand U5065 (N_5065,N_1048,N_2263);
xor U5066 (N_5066,N_1405,N_1245);
xor U5067 (N_5067,N_2911,N_162);
or U5068 (N_5068,N_4889,N_1392);
xnor U5069 (N_5069,N_1136,N_4651);
and U5070 (N_5070,N_751,N_1670);
and U5071 (N_5071,N_3677,N_615);
or U5072 (N_5072,N_1871,N_1116);
nand U5073 (N_5073,N_3793,N_695);
xnor U5074 (N_5074,N_921,N_4474);
nand U5075 (N_5075,N_1071,N_2139);
and U5076 (N_5076,N_2603,N_1369);
and U5077 (N_5077,N_980,N_1757);
xor U5078 (N_5078,N_3966,N_4963);
and U5079 (N_5079,N_3959,N_726);
nor U5080 (N_5080,N_17,N_1845);
nand U5081 (N_5081,N_4804,N_2616);
or U5082 (N_5082,N_4803,N_4795);
xor U5083 (N_5083,N_4682,N_3828);
or U5084 (N_5084,N_1468,N_2809);
and U5085 (N_5085,N_1763,N_3189);
or U5086 (N_5086,N_217,N_316);
nand U5087 (N_5087,N_4011,N_498);
or U5088 (N_5088,N_2791,N_4941);
nand U5089 (N_5089,N_2333,N_132);
xor U5090 (N_5090,N_2075,N_3929);
or U5091 (N_5091,N_3675,N_2231);
nor U5092 (N_5092,N_4334,N_2724);
or U5093 (N_5093,N_477,N_3548);
or U5094 (N_5094,N_3459,N_4880);
nor U5095 (N_5095,N_1001,N_2249);
xor U5096 (N_5096,N_4455,N_299);
nand U5097 (N_5097,N_4298,N_582);
or U5098 (N_5098,N_2801,N_1893);
or U5099 (N_5099,N_1953,N_1407);
or U5100 (N_5100,N_2868,N_328);
or U5101 (N_5101,N_4033,N_3443);
nand U5102 (N_5102,N_4570,N_2420);
xor U5103 (N_5103,N_2219,N_1185);
nor U5104 (N_5104,N_3775,N_4292);
or U5105 (N_5105,N_792,N_58);
nor U5106 (N_5106,N_3986,N_2651);
nor U5107 (N_5107,N_444,N_3427);
nand U5108 (N_5108,N_4460,N_549);
and U5109 (N_5109,N_1003,N_1960);
nand U5110 (N_5110,N_809,N_1754);
or U5111 (N_5111,N_838,N_1219);
nand U5112 (N_5112,N_2354,N_2854);
nor U5113 (N_5113,N_2371,N_1088);
xnor U5114 (N_5114,N_1844,N_4384);
xnor U5115 (N_5115,N_46,N_4337);
nor U5116 (N_5116,N_1469,N_1616);
and U5117 (N_5117,N_158,N_4161);
nor U5118 (N_5118,N_3378,N_3501);
or U5119 (N_5119,N_2921,N_257);
or U5120 (N_5120,N_810,N_4393);
nand U5121 (N_5121,N_3195,N_4850);
or U5122 (N_5122,N_4713,N_3015);
or U5123 (N_5123,N_3379,N_4120);
nor U5124 (N_5124,N_1879,N_4078);
nor U5125 (N_5125,N_1467,N_4732);
nand U5126 (N_5126,N_445,N_1169);
nand U5127 (N_5127,N_2508,N_3428);
and U5128 (N_5128,N_286,N_3310);
nand U5129 (N_5129,N_4984,N_3916);
or U5130 (N_5130,N_4774,N_4352);
xnor U5131 (N_5131,N_1899,N_1343);
xor U5132 (N_5132,N_1860,N_565);
and U5133 (N_5133,N_1207,N_1705);
nor U5134 (N_5134,N_1815,N_4173);
and U5135 (N_5135,N_1222,N_3908);
or U5136 (N_5136,N_600,N_1835);
nor U5137 (N_5137,N_2475,N_914);
nor U5138 (N_5138,N_3922,N_4162);
nand U5139 (N_5139,N_3996,N_3864);
nand U5140 (N_5140,N_2211,N_3232);
xor U5141 (N_5141,N_3612,N_265);
and U5142 (N_5142,N_732,N_198);
nor U5143 (N_5143,N_4262,N_1332);
and U5144 (N_5144,N_4953,N_2893);
xor U5145 (N_5145,N_3804,N_946);
xnor U5146 (N_5146,N_4468,N_2728);
nand U5147 (N_5147,N_4633,N_2201);
xnor U5148 (N_5148,N_3635,N_4872);
and U5149 (N_5149,N_1650,N_320);
nand U5150 (N_5150,N_4276,N_3291);
or U5151 (N_5151,N_2428,N_1171);
and U5152 (N_5152,N_1582,N_3944);
or U5153 (N_5153,N_929,N_3562);
xnor U5154 (N_5154,N_4375,N_3112);
and U5155 (N_5155,N_1931,N_1504);
or U5156 (N_5156,N_39,N_2114);
nor U5157 (N_5157,N_1984,N_3227);
nand U5158 (N_5158,N_3171,N_2647);
xor U5159 (N_5159,N_3845,N_3770);
or U5160 (N_5160,N_235,N_698);
xor U5161 (N_5161,N_2769,N_28);
nand U5162 (N_5162,N_2699,N_4197);
xor U5163 (N_5163,N_376,N_3269);
and U5164 (N_5164,N_1798,N_4693);
nor U5165 (N_5165,N_605,N_2117);
nor U5166 (N_5166,N_1359,N_515);
or U5167 (N_5167,N_1051,N_4707);
nand U5168 (N_5168,N_4184,N_1233);
nand U5169 (N_5169,N_387,N_3976);
and U5170 (N_5170,N_4561,N_2634);
nand U5171 (N_5171,N_3638,N_2712);
nor U5172 (N_5172,N_4502,N_1203);
or U5173 (N_5173,N_423,N_3216);
or U5174 (N_5174,N_2527,N_527);
or U5175 (N_5175,N_4841,N_4935);
nand U5176 (N_5176,N_2458,N_4621);
nand U5177 (N_5177,N_3346,N_1210);
nand U5178 (N_5178,N_2931,N_2734);
nand U5179 (N_5179,N_1270,N_2038);
nand U5180 (N_5180,N_394,N_1357);
and U5181 (N_5181,N_1613,N_4720);
or U5182 (N_5182,N_2661,N_761);
and U5183 (N_5183,N_2543,N_3312);
and U5184 (N_5184,N_2806,N_1340);
nor U5185 (N_5185,N_4106,N_4273);
or U5186 (N_5186,N_3871,N_3194);
nor U5187 (N_5187,N_1788,N_1635);
and U5188 (N_5188,N_1312,N_2838);
nor U5189 (N_5189,N_21,N_4088);
or U5190 (N_5190,N_4856,N_2704);
or U5191 (N_5191,N_2646,N_719);
and U5192 (N_5192,N_784,N_4532);
nand U5193 (N_5193,N_4839,N_712);
and U5194 (N_5194,N_944,N_2771);
and U5195 (N_5195,N_3678,N_708);
xor U5196 (N_5196,N_1621,N_2756);
or U5197 (N_5197,N_4081,N_3154);
nand U5198 (N_5198,N_3513,N_4085);
and U5199 (N_5199,N_4211,N_558);
and U5200 (N_5200,N_37,N_3756);
xor U5201 (N_5201,N_1975,N_1420);
xnor U5202 (N_5202,N_3229,N_4203);
xnor U5203 (N_5203,N_4849,N_4381);
nand U5204 (N_5204,N_2436,N_371);
or U5205 (N_5205,N_1111,N_4168);
and U5206 (N_5206,N_1243,N_3458);
nor U5207 (N_5207,N_1994,N_4109);
and U5208 (N_5208,N_2919,N_4045);
or U5209 (N_5209,N_1633,N_3345);
and U5210 (N_5210,N_2349,N_4221);
or U5211 (N_5211,N_49,N_2457);
and U5212 (N_5212,N_180,N_4882);
or U5213 (N_5213,N_4546,N_1505);
and U5214 (N_5214,N_4731,N_1646);
xnor U5215 (N_5215,N_1982,N_73);
nor U5216 (N_5216,N_1454,N_2070);
xor U5217 (N_5217,N_3784,N_3907);
or U5218 (N_5218,N_528,N_1099);
nor U5219 (N_5219,N_2024,N_4218);
nand U5220 (N_5220,N_2450,N_2929);
nor U5221 (N_5221,N_1373,N_3881);
nor U5222 (N_5222,N_786,N_4082);
nand U5223 (N_5223,N_1288,N_1933);
or U5224 (N_5224,N_1588,N_3438);
nand U5225 (N_5225,N_3333,N_228);
nand U5226 (N_5226,N_4727,N_138);
and U5227 (N_5227,N_4486,N_4741);
and U5228 (N_5228,N_4280,N_114);
and U5229 (N_5229,N_710,N_652);
xnor U5230 (N_5230,N_3064,N_3135);
xnor U5231 (N_5231,N_4353,N_3090);
xor U5232 (N_5232,N_3858,N_4412);
and U5233 (N_5233,N_4890,N_1247);
nand U5234 (N_5234,N_2439,N_44);
xor U5235 (N_5235,N_1719,N_4345);
nand U5236 (N_5236,N_770,N_4521);
nor U5237 (N_5237,N_2494,N_4637);
nor U5238 (N_5238,N_876,N_1710);
nand U5239 (N_5239,N_525,N_2162);
and U5240 (N_5240,N_2693,N_2510);
and U5241 (N_5241,N_3579,N_3146);
or U5242 (N_5242,N_127,N_827);
and U5243 (N_5243,N_967,N_2434);
xor U5244 (N_5244,N_4617,N_3898);
or U5245 (N_5245,N_862,N_998);
nor U5246 (N_5246,N_3471,N_985);
or U5247 (N_5247,N_904,N_936);
nand U5248 (N_5248,N_1301,N_1802);
nor U5249 (N_5249,N_847,N_3185);
nor U5250 (N_5250,N_2532,N_4287);
nor U5251 (N_5251,N_3868,N_844);
xor U5252 (N_5252,N_3165,N_1295);
xor U5253 (N_5253,N_2072,N_1221);
xor U5254 (N_5254,N_4138,N_4070);
or U5255 (N_5255,N_4285,N_1575);
or U5256 (N_5256,N_4158,N_1819);
nand U5257 (N_5257,N_2179,N_2111);
xor U5258 (N_5258,N_2968,N_2279);
and U5259 (N_5259,N_1784,N_2669);
nand U5260 (N_5260,N_2875,N_1568);
xnor U5261 (N_5261,N_2140,N_4860);
and U5262 (N_5262,N_3037,N_3550);
or U5263 (N_5263,N_4252,N_2748);
nor U5264 (N_5264,N_4464,N_850);
and U5265 (N_5265,N_830,N_3575);
nor U5266 (N_5266,N_4624,N_1351);
nor U5267 (N_5267,N_1033,N_4642);
nor U5268 (N_5268,N_3651,N_403);
nor U5269 (N_5269,N_1310,N_4654);
and U5270 (N_5270,N_2775,N_3574);
or U5271 (N_5271,N_1806,N_191);
and U5272 (N_5272,N_4821,N_4258);
or U5273 (N_5273,N_4628,N_3683);
nand U5274 (N_5274,N_4603,N_4937);
or U5275 (N_5275,N_2762,N_3702);
xor U5276 (N_5276,N_3570,N_2513);
and U5277 (N_5277,N_368,N_4746);
and U5278 (N_5278,N_3931,N_4555);
nor U5279 (N_5279,N_2779,N_3633);
or U5280 (N_5280,N_1032,N_3414);
or U5281 (N_5281,N_150,N_2687);
and U5282 (N_5282,N_4260,N_1403);
and U5283 (N_5283,N_1576,N_4805);
nor U5284 (N_5284,N_4433,N_1281);
and U5285 (N_5285,N_4372,N_2363);
and U5286 (N_5286,N_908,N_429);
xor U5287 (N_5287,N_2286,N_2718);
nand U5288 (N_5288,N_2877,N_3630);
and U5289 (N_5289,N_983,N_564);
xor U5290 (N_5290,N_2653,N_3958);
and U5291 (N_5291,N_4644,N_156);
and U5292 (N_5292,N_81,N_3581);
nor U5293 (N_5293,N_4369,N_1402);
xnor U5294 (N_5294,N_503,N_2817);
nor U5295 (N_5295,N_4869,N_2599);
and U5296 (N_5296,N_3887,N_3436);
and U5297 (N_5297,N_238,N_4611);
and U5298 (N_5298,N_3235,N_144);
and U5299 (N_5299,N_411,N_2684);
nor U5300 (N_5300,N_4750,N_2852);
and U5301 (N_5301,N_3540,N_1560);
or U5302 (N_5302,N_1132,N_2862);
or U5303 (N_5303,N_3610,N_1000);
xnor U5304 (N_5304,N_155,N_4302);
nor U5305 (N_5305,N_2421,N_3693);
and U5306 (N_5306,N_2053,N_2301);
or U5307 (N_5307,N_4745,N_4696);
or U5308 (N_5308,N_3698,N_4282);
nor U5309 (N_5309,N_288,N_2985);
xor U5310 (N_5310,N_4801,N_550);
xnor U5311 (N_5311,N_3382,N_4881);
xnor U5312 (N_5312,N_1018,N_3150);
nand U5313 (N_5313,N_3588,N_824);
nand U5314 (N_5314,N_3315,N_3854);
xor U5315 (N_5315,N_2061,N_3978);
xnor U5316 (N_5316,N_1927,N_909);
nand U5317 (N_5317,N_808,N_581);
and U5318 (N_5318,N_959,N_923);
and U5319 (N_5319,N_4049,N_4958);
and U5320 (N_5320,N_2473,N_2234);
nand U5321 (N_5321,N_4355,N_3704);
and U5322 (N_5322,N_4620,N_1063);
nand U5323 (N_5323,N_4847,N_3563);
and U5324 (N_5324,N_4398,N_1506);
nand U5325 (N_5325,N_1450,N_1829);
or U5326 (N_5326,N_4939,N_2845);
nand U5327 (N_5327,N_2296,N_3981);
nor U5328 (N_5328,N_398,N_545);
or U5329 (N_5329,N_4729,N_4017);
xnor U5330 (N_5330,N_2265,N_721);
xnor U5331 (N_5331,N_1325,N_483);
or U5332 (N_5332,N_4764,N_3118);
nand U5333 (N_5333,N_2180,N_3740);
nor U5334 (N_5334,N_280,N_3945);
nand U5335 (N_5335,N_4465,N_3460);
nand U5336 (N_5336,N_3254,N_1250);
nand U5337 (N_5337,N_4151,N_783);
or U5338 (N_5338,N_2853,N_3045);
or U5339 (N_5339,N_2666,N_1117);
nor U5340 (N_5340,N_1878,N_2976);
nand U5341 (N_5341,N_232,N_4782);
or U5342 (N_5342,N_2814,N_4264);
nor U5343 (N_5343,N_4386,N_701);
and U5344 (N_5344,N_3243,N_4572);
nor U5345 (N_5345,N_2992,N_4638);
xnor U5346 (N_5346,N_2639,N_3629);
and U5347 (N_5347,N_4816,N_3178);
xnor U5348 (N_5348,N_3499,N_2591);
xor U5349 (N_5349,N_287,N_330);
or U5350 (N_5350,N_1431,N_4975);
nor U5351 (N_5351,N_60,N_4212);
nand U5352 (N_5352,N_2184,N_1535);
or U5353 (N_5353,N_3558,N_4646);
xor U5354 (N_5354,N_2086,N_4722);
nand U5355 (N_5355,N_3634,N_2376);
nand U5356 (N_5356,N_2325,N_1424);
and U5357 (N_5357,N_757,N_1306);
xnor U5358 (N_5358,N_3301,N_1930);
xor U5359 (N_5359,N_1186,N_4970);
nor U5360 (N_5360,N_128,N_2143);
nand U5361 (N_5361,N_4916,N_1493);
or U5362 (N_5362,N_840,N_3322);
nor U5363 (N_5363,N_711,N_601);
nor U5364 (N_5364,N_3484,N_1198);
nand U5365 (N_5365,N_4960,N_4461);
or U5366 (N_5366,N_4793,N_3641);
xor U5367 (N_5367,N_4286,N_2673);
xnor U5368 (N_5368,N_4222,N_4016);
or U5369 (N_5369,N_750,N_2623);
nor U5370 (N_5370,N_2902,N_11);
xnor U5371 (N_5371,N_203,N_4594);
and U5372 (N_5372,N_2045,N_1160);
or U5373 (N_5373,N_227,N_1364);
and U5374 (N_5374,N_4471,N_657);
or U5375 (N_5375,N_2923,N_4419);
nand U5376 (N_5376,N_4267,N_2454);
nor U5377 (N_5377,N_1479,N_2088);
xnor U5378 (N_5378,N_1253,N_4323);
and U5379 (N_5379,N_392,N_2064);
or U5380 (N_5380,N_1767,N_2089);
nor U5381 (N_5381,N_3523,N_181);
nor U5382 (N_5382,N_2320,N_2396);
xnor U5383 (N_5383,N_3014,N_3771);
and U5384 (N_5384,N_4427,N_2268);
and U5385 (N_5385,N_3730,N_3405);
nor U5386 (N_5386,N_2135,N_1311);
nand U5387 (N_5387,N_3712,N_1913);
and U5388 (N_5388,N_1681,N_1362);
xnor U5389 (N_5389,N_588,N_3977);
or U5390 (N_5390,N_3913,N_4227);
and U5391 (N_5391,N_3524,N_1174);
or U5392 (N_5392,N_1327,N_4329);
xnor U5393 (N_5393,N_465,N_3426);
nor U5394 (N_5394,N_1110,N_3417);
xor U5395 (N_5395,N_795,N_1769);
nor U5396 (N_5396,N_369,N_4288);
or U5397 (N_5397,N_2105,N_1707);
nor U5398 (N_5398,N_2155,N_1715);
and U5399 (N_5399,N_1732,N_1985);
nand U5400 (N_5400,N_221,N_1138);
and U5401 (N_5401,N_2569,N_3902);
nand U5402 (N_5402,N_4180,N_2182);
or U5403 (N_5403,N_2721,N_2207);
nor U5404 (N_5404,N_3733,N_584);
or U5405 (N_5405,N_1759,N_4964);
and U5406 (N_5406,N_2364,N_2375);
nand U5407 (N_5407,N_4936,N_2306);
xnor U5408 (N_5408,N_540,N_4797);
nor U5409 (N_5409,N_1014,N_1330);
and U5410 (N_5410,N_3094,N_4668);
xor U5411 (N_5411,N_1685,N_2614);
nor U5412 (N_5412,N_2733,N_460);
or U5413 (N_5413,N_4991,N_139);
nand U5414 (N_5414,N_2492,N_1);
and U5415 (N_5415,N_3643,N_3324);
and U5416 (N_5416,N_4670,N_2767);
nor U5417 (N_5417,N_1915,N_4772);
nor U5418 (N_5418,N_3984,N_2670);
or U5419 (N_5419,N_1386,N_797);
xnor U5420 (N_5420,N_661,N_1495);
or U5421 (N_5421,N_3656,N_643);
nand U5422 (N_5422,N_2847,N_1697);
xnor U5423 (N_5423,N_979,N_4462);
xnor U5424 (N_5424,N_3852,N_991);
or U5425 (N_5425,N_2382,N_1512);
and U5426 (N_5426,N_4602,N_1030);
and U5427 (N_5427,N_3082,N_656);
nand U5428 (N_5428,N_3445,N_4765);
nand U5429 (N_5429,N_3421,N_3303);
nand U5430 (N_5430,N_633,N_3567);
nand U5431 (N_5431,N_3363,N_1649);
nor U5432 (N_5432,N_4548,N_2460);
nand U5433 (N_5433,N_4798,N_1224);
nand U5434 (N_5434,N_1881,N_1643);
or U5435 (N_5435,N_439,N_962);
and U5436 (N_5436,N_2795,N_2052);
nand U5437 (N_5437,N_2540,N_4906);
nor U5438 (N_5438,N_87,N_4056);
or U5439 (N_5439,N_4265,N_450);
or U5440 (N_5440,N_2648,N_2690);
and U5441 (N_5441,N_1282,N_1564);
nand U5442 (N_5442,N_2082,N_1241);
or U5443 (N_5443,N_4893,N_596);
and U5444 (N_5444,N_149,N_4526);
nor U5445 (N_5445,N_739,N_4758);
and U5446 (N_5446,N_2575,N_956);
or U5447 (N_5447,N_3163,N_4551);
or U5448 (N_5448,N_2595,N_723);
nor U5449 (N_5449,N_212,N_2336);
nor U5450 (N_5450,N_2257,N_513);
nor U5451 (N_5451,N_4819,N_1199);
nor U5452 (N_5452,N_3980,N_2427);
and U5453 (N_5453,N_4086,N_4808);
nand U5454 (N_5454,N_1531,N_2329);
and U5455 (N_5455,N_415,N_1602);
nand U5456 (N_5456,N_4364,N_1074);
nand U5457 (N_5457,N_2366,N_338);
or U5458 (N_5458,N_1413,N_2597);
and U5459 (N_5459,N_140,N_2107);
nand U5460 (N_5460,N_2635,N_1928);
or U5461 (N_5461,N_532,N_373);
and U5462 (N_5462,N_2292,N_3168);
or U5463 (N_5463,N_488,N_3925);
nand U5464 (N_5464,N_4796,N_4562);
or U5465 (N_5465,N_3372,N_1652);
and U5466 (N_5466,N_1070,N_3326);
and U5467 (N_5467,N_730,N_4092);
nor U5468 (N_5468,N_4556,N_972);
nand U5469 (N_5469,N_4600,N_717);
and U5470 (N_5470,N_1050,N_2908);
and U5471 (N_5471,N_529,N_806);
or U5472 (N_5472,N_2568,N_4466);
and U5473 (N_5473,N_2299,N_2585);
nand U5474 (N_5474,N_963,N_3824);
nand U5475 (N_5475,N_3463,N_512);
xor U5476 (N_5476,N_4525,N_725);
xnor U5477 (N_5477,N_3578,N_116);
and U5478 (N_5478,N_3297,N_1358);
or U5479 (N_5479,N_1886,N_1991);
nand U5480 (N_5480,N_84,N_3174);
and U5481 (N_5481,N_2878,N_2271);
xnor U5482 (N_5482,N_293,N_4202);
nand U5483 (N_5483,N_573,N_1713);
xnor U5484 (N_5484,N_4204,N_3341);
and U5485 (N_5485,N_3729,N_2520);
and U5486 (N_5486,N_1388,N_41);
or U5487 (N_5487,N_3988,N_602);
nor U5488 (N_5488,N_4601,N_75);
nand U5489 (N_5489,N_2642,N_586);
and U5490 (N_5490,N_1714,N_241);
nand U5491 (N_5491,N_506,N_1240);
xor U5492 (N_5492,N_957,N_1257);
or U5493 (N_5493,N_3745,N_0);
xnor U5494 (N_5494,N_3138,N_2840);
nand U5495 (N_5495,N_803,N_561);
nor U5496 (N_5496,N_3409,N_3273);
nand U5497 (N_5497,N_3295,N_1459);
and U5498 (N_5498,N_886,N_2945);
or U5499 (N_5499,N_871,N_2049);
xor U5500 (N_5500,N_3967,N_2887);
or U5501 (N_5501,N_2993,N_2130);
and U5502 (N_5502,N_3495,N_3939);
nand U5503 (N_5503,N_245,N_4981);
and U5504 (N_5504,N_4430,N_3726);
nand U5505 (N_5505,N_4789,N_546);
xnor U5506 (N_5506,N_497,N_1010);
nor U5507 (N_5507,N_1471,N_4191);
and U5508 (N_5508,N_1335,N_4683);
xnor U5509 (N_5509,N_1368,N_766);
or U5510 (N_5510,N_772,N_3965);
xor U5511 (N_5511,N_1414,N_4063);
xnor U5512 (N_5512,N_4498,N_38);
nand U5513 (N_5513,N_1511,N_1903);
nor U5514 (N_5514,N_3130,N_4385);
or U5515 (N_5515,N_1909,N_3078);
and U5516 (N_5516,N_1747,N_3522);
xnor U5517 (N_5517,N_1267,N_678);
and U5518 (N_5518,N_3342,N_1651);
xor U5519 (N_5519,N_360,N_3617);
or U5520 (N_5520,N_3777,N_222);
and U5521 (N_5521,N_2981,N_3863);
xnor U5522 (N_5522,N_1552,N_3175);
and U5523 (N_5523,N_3128,N_3311);
xor U5524 (N_5524,N_2035,N_3258);
nand U5525 (N_5525,N_4697,N_1733);
and U5526 (N_5526,N_3600,N_4490);
and U5527 (N_5527,N_3167,N_4884);
nand U5528 (N_5528,N_1205,N_625);
and U5529 (N_5529,N_2054,N_223);
or U5530 (N_5530,N_3096,N_2447);
and U5531 (N_5531,N_820,N_3387);
nor U5532 (N_5532,N_518,N_1382);
xor U5533 (N_5533,N_3769,N_1292);
or U5534 (N_5534,N_1374,N_2032);
nand U5535 (N_5535,N_1193,N_1487);
nand U5536 (N_5536,N_2391,N_1785);
nand U5537 (N_5537,N_3240,N_616);
and U5538 (N_5538,N_3754,N_4749);
nor U5539 (N_5539,N_4097,N_741);
xnor U5540 (N_5540,N_2110,N_2630);
or U5541 (N_5541,N_2864,N_3474);
nor U5542 (N_5542,N_1718,N_3158);
and U5543 (N_5543,N_731,N_3234);
xnor U5544 (N_5544,N_424,N_1170);
nor U5545 (N_5545,N_3721,N_427);
and U5546 (N_5546,N_2944,N_3126);
nand U5547 (N_5547,N_2821,N_822);
nor U5548 (N_5548,N_1967,N_2518);
nand U5549 (N_5549,N_2914,N_4201);
or U5550 (N_5550,N_2262,N_1557);
nor U5551 (N_5551,N_173,N_3644);
and U5552 (N_5552,N_1522,N_1700);
nand U5553 (N_5553,N_4156,N_2015);
nand U5554 (N_5554,N_2497,N_3450);
and U5555 (N_5555,N_2894,N_3862);
and U5556 (N_5556,N_3613,N_2019);
nand U5557 (N_5557,N_4395,N_4303);
and U5558 (N_5558,N_3,N_2503);
nand U5559 (N_5559,N_3136,N_1755);
nand U5560 (N_5560,N_4496,N_4420);
and U5561 (N_5561,N_1321,N_3571);
xor U5562 (N_5562,N_3856,N_4547);
xor U5563 (N_5563,N_1381,N_1480);
xnor U5564 (N_5564,N_195,N_428);
nand U5565 (N_5565,N_2675,N_1693);
nor U5566 (N_5566,N_3173,N_2986);
or U5567 (N_5567,N_4516,N_16);
and U5568 (N_5568,N_4721,N_1810);
or U5569 (N_5569,N_4718,N_3507);
nand U5570 (N_5570,N_4021,N_1384);
and U5571 (N_5571,N_541,N_1274);
xnor U5572 (N_5572,N_1079,N_851);
nor U5573 (N_5573,N_3963,N_4121);
nor U5574 (N_5574,N_3123,N_1691);
or U5575 (N_5575,N_3480,N_4535);
or U5576 (N_5576,N_3835,N_3498);
nand U5577 (N_5577,N_4684,N_2431);
xor U5578 (N_5578,N_3846,N_4896);
nand U5579 (N_5579,N_4025,N_493);
xor U5580 (N_5580,N_880,N_578);
or U5581 (N_5581,N_4359,N_4193);
xor U5582 (N_5582,N_4448,N_1291);
nand U5583 (N_5583,N_4910,N_4530);
or U5584 (N_5584,N_3468,N_4034);
nor U5585 (N_5585,N_1962,N_2332);
xor U5586 (N_5586,N_1726,N_361);
or U5587 (N_5587,N_2542,N_397);
or U5588 (N_5588,N_832,N_4389);
nand U5589 (N_5589,N_671,N_542);
or U5590 (N_5590,N_2157,N_4701);
xor U5591 (N_5591,N_679,N_1031);
nor U5592 (N_5592,N_267,N_1839);
and U5593 (N_5593,N_4631,N_3068);
or U5594 (N_5594,N_4463,N_689);
nor U5595 (N_5595,N_197,N_170);
xor U5596 (N_5596,N_1451,N_2984);
nor U5597 (N_5597,N_4778,N_3198);
nand U5598 (N_5598,N_4002,N_3305);
nor U5599 (N_5599,N_873,N_857);
or U5600 (N_5600,N_1594,N_4347);
nand U5601 (N_5601,N_4814,N_2283);
nor U5602 (N_5602,N_2148,N_2435);
or U5603 (N_5603,N_55,N_3636);
xor U5604 (N_5604,N_2731,N_4153);
xnor U5605 (N_5605,N_2886,N_1130);
and U5606 (N_5606,N_2395,N_1423);
nand U5607 (N_5607,N_1606,N_4100);
or U5608 (N_5608,N_520,N_496);
xor U5609 (N_5609,N_1302,N_4545);
or U5610 (N_5610,N_694,N_3992);
nor U5611 (N_5611,N_3073,N_4409);
nand U5612 (N_5612,N_753,N_1738);
nand U5613 (N_5613,N_2239,N_2657);
and U5614 (N_5614,N_3029,N_3587);
and U5615 (N_5615,N_4794,N_384);
or U5616 (N_5616,N_4406,N_2707);
nor U5617 (N_5617,N_973,N_2351);
xnor U5618 (N_5618,N_1867,N_4779);
nor U5619 (N_5619,N_2572,N_897);
or U5620 (N_5620,N_4136,N_1859);
and U5621 (N_5621,N_1745,N_734);
nand U5622 (N_5622,N_3147,N_1794);
nor U5623 (N_5623,N_2671,N_3200);
nor U5624 (N_5624,N_1435,N_4144);
nor U5625 (N_5625,N_3941,N_2844);
nand U5626 (N_5626,N_1189,N_2321);
and U5627 (N_5627,N_14,N_3773);
xor U5628 (N_5628,N_508,N_2511);
nor U5629 (N_5629,N_86,N_407);
xor U5630 (N_5630,N_2678,N_4708);
and U5631 (N_5631,N_2476,N_225);
nand U5632 (N_5632,N_97,N_3051);
nor U5633 (N_5633,N_2170,N_294);
and U5634 (N_5634,N_1489,N_4188);
nand U5635 (N_5635,N_4232,N_668);
nor U5636 (N_5636,N_2005,N_262);
xor U5637 (N_5637,N_1910,N_4581);
or U5638 (N_5638,N_802,N_773);
nor U5639 (N_5639,N_1023,N_4370);
and U5640 (N_5640,N_4519,N_1264);
and U5641 (N_5641,N_1923,N_1999);
and U5642 (N_5642,N_1348,N_3318);
nand U5643 (N_5643,N_4210,N_306);
and U5644 (N_5644,N_2726,N_3969);
or U5645 (N_5645,N_3528,N_2882);
nor U5646 (N_5646,N_2300,N_2823);
nand U5647 (N_5647,N_3736,N_2766);
nor U5648 (N_5648,N_4911,N_4289);
or U5649 (N_5649,N_4247,N_175);
nand U5650 (N_5650,N_3402,N_2936);
nand U5651 (N_5651,N_2871,N_4781);
xnor U5652 (N_5652,N_4434,N_648);
nor U5653 (N_5653,N_2810,N_2258);
nand U5654 (N_5654,N_2318,N_1862);
and U5655 (N_5655,N_2545,N_807);
nor U5656 (N_5656,N_279,N_4217);
nor U5657 (N_5657,N_4605,N_1825);
xor U5658 (N_5658,N_1586,N_4015);
xor U5659 (N_5659,N_1619,N_1801);
and U5660 (N_5660,N_3371,N_4128);
or U5661 (N_5661,N_4005,N_3095);
and U5662 (N_5662,N_3951,N_2146);
or U5663 (N_5663,N_1764,N_3410);
nand U5664 (N_5664,N_2060,N_3313);
and U5665 (N_5665,N_4902,N_3857);
or U5666 (N_5666,N_500,N_1075);
nor U5667 (N_5667,N_4174,N_4415);
and U5668 (N_5668,N_2830,N_3103);
nand U5669 (N_5669,N_4681,N_2786);
or U5670 (N_5670,N_1543,N_1113);
nor U5671 (N_5671,N_3673,N_247);
nor U5672 (N_5672,N_34,N_697);
nand U5673 (N_5673,N_202,N_1179);
xnor U5674 (N_5674,N_1856,N_892);
xnor U5675 (N_5675,N_192,N_2095);
nor U5676 (N_5676,N_2026,N_2906);
nand U5677 (N_5677,N_3743,N_882);
nand U5678 (N_5678,N_1486,N_4710);
or U5679 (N_5679,N_3626,N_4093);
nand U5680 (N_5680,N_4671,N_3870);
nor U5681 (N_5681,N_1408,N_2811);
and U5682 (N_5682,N_3211,N_3973);
and U5683 (N_5683,N_3547,N_4724);
nor U5684 (N_5684,N_4980,N_2963);
and U5685 (N_5685,N_3376,N_209);
nor U5686 (N_5686,N_816,N_2327);
xor U5687 (N_5687,N_3720,N_2033);
xor U5688 (N_5688,N_684,N_464);
xnor U5689 (N_5689,N_2761,N_1720);
nor U5690 (N_5690,N_4306,N_554);
nor U5691 (N_5691,N_1623,N_3645);
and U5692 (N_5692,N_2168,N_406);
or U5693 (N_5693,N_3652,N_3709);
nand U5694 (N_5694,N_434,N_1501);
nand U5695 (N_5695,N_248,N_3012);
and U5696 (N_5696,N_510,N_487);
nor U5697 (N_5697,N_867,N_1583);
nor U5698 (N_5698,N_4339,N_3503);
nor U5699 (N_5699,N_2142,N_3395);
nor U5700 (N_5700,N_2251,N_3920);
nand U5701 (N_5701,N_259,N_631);
or U5702 (N_5702,N_752,N_4150);
nand U5703 (N_5703,N_3667,N_4048);
xor U5704 (N_5704,N_2237,N_2863);
nand U5705 (N_5705,N_4650,N_3245);
nand U5706 (N_5706,N_3149,N_4152);
or U5707 (N_5707,N_326,N_2174);
nor U5708 (N_5708,N_1095,N_2073);
or U5709 (N_5709,N_1618,N_216);
and U5710 (N_5710,N_3794,N_2587);
nor U5711 (N_5711,N_618,N_2352);
nand U5712 (N_5712,N_3847,N_819);
nor U5713 (N_5713,N_629,N_3019);
xor U5714 (N_5714,N_1926,N_2956);
and U5715 (N_5715,N_3097,N_3020);
and U5716 (N_5716,N_3203,N_3456);
xor U5717 (N_5717,N_639,N_1695);
nor U5718 (N_5718,N_3866,N_2698);
or U5719 (N_5719,N_4178,N_4451);
or U5720 (N_5720,N_3714,N_448);
nand U5721 (N_5721,N_345,N_256);
xor U5722 (N_5722,N_1969,N_133);
nor U5723 (N_5723,N_4233,N_1355);
and U5724 (N_5724,N_1900,N_1698);
nand U5725 (N_5725,N_2658,N_4728);
nand U5726 (N_5726,N_901,N_2361);
or U5727 (N_5727,N_68,N_919);
nor U5728 (N_5728,N_1760,N_4024);
nand U5729 (N_5729,N_2013,N_1309);
and U5730 (N_5730,N_4743,N_1304);
or U5731 (N_5731,N_4643,N_3075);
nor U5732 (N_5732,N_4067,N_887);
nand U5733 (N_5733,N_4098,N_3415);
nor U5734 (N_5734,N_281,N_4008);
and U5735 (N_5735,N_2869,N_4848);
xnor U5736 (N_5736,N_3706,N_389);
xnor U5737 (N_5737,N_1795,N_2495);
and U5738 (N_5738,N_4844,N_3734);
xor U5739 (N_5739,N_975,N_1328);
and U5740 (N_5740,N_4733,N_20);
and U5741 (N_5741,N_1188,N_312);
and U5742 (N_5742,N_472,N_152);
nand U5743 (N_5743,N_4657,N_4878);
or U5744 (N_5744,N_3359,N_2144);
or U5745 (N_5745,N_1360,N_856);
or U5746 (N_5746,N_4686,N_2996);
xor U5747 (N_5747,N_4944,N_3035);
nor U5748 (N_5748,N_2297,N_3080);
nor U5749 (N_5749,N_4340,N_3972);
and U5750 (N_5750,N_1786,N_620);
nor U5751 (N_5751,N_4517,N_473);
nand U5752 (N_5752,N_2269,N_2829);
nor U5753 (N_5753,N_377,N_591);
and U5754 (N_5754,N_4503,N_568);
or U5755 (N_5755,N_3006,N_3515);
or U5756 (N_5756,N_3028,N_36);
xnor U5757 (N_5757,N_570,N_4058);
xor U5758 (N_5758,N_18,N_2695);
and U5759 (N_5759,N_2904,N_516);
or U5760 (N_5760,N_4553,N_3212);
nand U5761 (N_5761,N_968,N_4402);
xor U5762 (N_5762,N_4467,N_1052);
xor U5763 (N_5763,N_4342,N_981);
and U5764 (N_5764,N_899,N_1550);
and U5765 (N_5765,N_4079,N_1399);
xnor U5766 (N_5766,N_1244,N_4160);
xor U5767 (N_5767,N_3226,N_1005);
and U5768 (N_5768,N_4099,N_987);
nand U5769 (N_5769,N_2785,N_2660);
nor U5770 (N_5770,N_839,N_1978);
nor U5771 (N_5771,N_3098,N_2316);
or U5772 (N_5772,N_703,N_4514);
xnor U5773 (N_5773,N_4062,N_4622);
xor U5774 (N_5774,N_1181,N_4446);
xnor U5775 (N_5775,N_2252,N_3388);
and U5776 (N_5776,N_1073,N_1315);
and U5777 (N_5777,N_3529,N_1509);
xnor U5778 (N_5778,N_3530,N_2782);
nand U5779 (N_5779,N_4113,N_4312);
or U5780 (N_5780,N_4533,N_3059);
nand U5781 (N_5781,N_995,N_1847);
nor U5782 (N_5782,N_621,N_3596);
xnor U5783 (N_5783,N_4606,N_3027);
nor U5784 (N_5784,N_4295,N_2946);
xnor U5785 (N_5785,N_1541,N_2009);
xor U5786 (N_5786,N_1791,N_2037);
or U5787 (N_5787,N_419,N_3288);
nand U5788 (N_5788,N_4932,N_4275);
nand U5789 (N_5789,N_2592,N_3631);
xnor U5790 (N_5790,N_3886,N_492);
xor U5791 (N_5791,N_2090,N_4362);
xor U5792 (N_5792,N_1236,N_495);
xor U5793 (N_5793,N_2903,N_468);
nand U5794 (N_5794,N_3607,N_4744);
nand U5795 (N_5795,N_3660,N_2243);
nand U5796 (N_5796,N_2884,N_4540);
nand U5797 (N_5797,N_4392,N_2787);
nor U5798 (N_5798,N_142,N_2141);
xor U5799 (N_5799,N_3805,N_3874);
and U5800 (N_5800,N_702,N_1232);
nor U5801 (N_5801,N_4206,N_2681);
nor U5802 (N_5802,N_552,N_3599);
nor U5803 (N_5803,N_4513,N_474);
or U5804 (N_5804,N_3264,N_3739);
or U5805 (N_5805,N_1015,N_3011);
and U5806 (N_5806,N_3183,N_938);
xnor U5807 (N_5807,N_4112,N_244);
nor U5808 (N_5808,N_2334,N_3321);
nand U5809 (N_5809,N_1780,N_2169);
nor U5810 (N_5810,N_3830,N_1863);
nand U5811 (N_5811,N_3891,N_3900);
and U5812 (N_5812,N_2308,N_1055);
or U5813 (N_5813,N_4761,N_1884);
and U5814 (N_5814,N_1455,N_907);
nor U5815 (N_5815,N_3763,N_3533);
or U5816 (N_5816,N_402,N_2533);
and U5817 (N_5817,N_628,N_964);
nor U5818 (N_5818,N_309,N_1006);
and U5819 (N_5819,N_4236,N_3572);
nor U5820 (N_5820,N_2304,N_3889);
nand U5821 (N_5821,N_1590,N_4250);
and U5822 (N_5822,N_977,N_1090);
and U5823 (N_5823,N_3434,N_3646);
nand U5824 (N_5824,N_4652,N_1983);
nand U5825 (N_5825,N_4917,N_2478);
nand U5826 (N_5826,N_869,N_4031);
xnor U5827 (N_5827,N_1080,N_4832);
nand U5828 (N_5828,N_1885,N_1337);
xnor U5829 (N_5829,N_2360,N_2918);
xor U5830 (N_5830,N_3701,N_1391);
xor U5831 (N_5831,N_4114,N_292);
nand U5832 (N_5832,N_207,N_1404);
nand U5833 (N_5833,N_4931,N_457);
or U5834 (N_5834,N_2165,N_4075);
nor U5835 (N_5835,N_1009,N_2735);
nand U5836 (N_5836,N_3724,N_865);
nand U5837 (N_5837,N_250,N_932);
nor U5838 (N_5838,N_1307,N_425);
and U5839 (N_5839,N_1086,N_2703);
and U5840 (N_5840,N_4604,N_311);
nor U5841 (N_5841,N_553,N_3285);
xnor U5842 (N_5842,N_2189,N_955);
xnor U5843 (N_5843,N_1175,N_3531);
or U5844 (N_5844,N_1338,N_4170);
or U5845 (N_5845,N_4141,N_1026);
nand U5846 (N_5846,N_2025,N_3757);
or U5847 (N_5847,N_4123,N_2757);
and U5848 (N_5848,N_52,N_386);
nor U5849 (N_5849,N_3441,N_3818);
and U5850 (N_5850,N_823,N_481);
and U5851 (N_5851,N_4074,N_4068);
nand U5852 (N_5852,N_2108,N_4354);
xor U5853 (N_5853,N_3489,N_1148);
xor U5854 (N_5854,N_196,N_2502);
nand U5855 (N_5855,N_1154,N_3820);
xor U5856 (N_5856,N_4512,N_3137);
and U5857 (N_5857,N_126,N_682);
nor U5858 (N_5858,N_2459,N_3672);
and U5859 (N_5859,N_3995,N_1037);
xor U5860 (N_5860,N_3253,N_2643);
xnor U5861 (N_5861,N_2493,N_3787);
nor U5862 (N_5862,N_2896,N_1902);
or U5863 (N_5863,N_27,N_3911);
xnor U5864 (N_5864,N_3423,N_989);
or U5865 (N_5865,N_1842,N_1595);
or U5866 (N_5866,N_2150,N_1119);
nor U5867 (N_5867,N_4215,N_3597);
and U5868 (N_5868,N_1167,N_1437);
nor U5869 (N_5869,N_3374,N_2030);
and U5870 (N_5870,N_4026,N_2331);
nor U5871 (N_5871,N_556,N_4965);
nand U5872 (N_5872,N_304,N_4304);
or U5873 (N_5873,N_3089,N_1989);
xnor U5874 (N_5874,N_2177,N_902);
and U5875 (N_5875,N_4230,N_3519);
or U5876 (N_5876,N_2557,N_4360);
xnor U5877 (N_5877,N_2556,N_931);
nor U5878 (N_5878,N_215,N_4868);
or U5879 (N_5879,N_2732,N_442);
nor U5880 (N_5880,N_9,N_4515);
nor U5881 (N_5881,N_4951,N_3640);
xnor U5882 (N_5882,N_2433,N_3663);
nand U5883 (N_5883,N_2611,N_2624);
nand U5884 (N_5884,N_4055,N_2415);
or U5885 (N_5885,N_1433,N_2942);
and U5886 (N_5886,N_2600,N_942);
nand U5887 (N_5887,N_3549,N_2926);
nand U5888 (N_5888,N_2158,N_3025);
or U5889 (N_5889,N_1973,N_2101);
and U5890 (N_5890,N_3982,N_2195);
or U5891 (N_5891,N_1770,N_475);
nand U5892 (N_5892,N_815,N_2291);
nand U5893 (N_5893,N_2708,N_1818);
nand U5894 (N_5894,N_3044,N_2172);
and U5895 (N_5895,N_206,N_2676);
nor U5896 (N_5896,N_65,N_853);
xnor U5897 (N_5897,N_270,N_2392);
nand U5898 (N_5898,N_3717,N_1238);
or U5899 (N_5899,N_3224,N_2288);
xnor U5900 (N_5900,N_4537,N_4982);
nor U5901 (N_5901,N_1837,N_2565);
nand U5902 (N_5902,N_768,N_1127);
or U5903 (N_5903,N_3225,N_2584);
or U5904 (N_5904,N_935,N_347);
or U5905 (N_5905,N_4837,N_2190);
nor U5906 (N_5906,N_100,N_4812);
nor U5907 (N_5907,N_3609,N_3584);
xor U5908 (N_5908,N_480,N_4299);
or U5909 (N_5909,N_2173,N_2326);
or U5910 (N_5910,N_4903,N_2835);
xor U5911 (N_5911,N_4084,N_603);
xnor U5912 (N_5912,N_1375,N_785);
or U5913 (N_5913,N_146,N_4330);
nand U5914 (N_5914,N_4865,N_1584);
and U5915 (N_5915,N_4552,N_2043);
xnor U5916 (N_5916,N_4,N_3792);
or U5917 (N_5917,N_355,N_3657);
or U5918 (N_5918,N_4000,N_4317);
nor U5919 (N_5919,N_2723,N_1706);
and U5920 (N_5920,N_2960,N_1963);
nor U5921 (N_5921,N_3397,N_1082);
xor U5922 (N_5922,N_1699,N_297);
xor U5923 (N_5923,N_263,N_3166);
nor U5924 (N_5924,N_4432,N_4316);
or U5925 (N_5925,N_3715,N_1724);
xnor U5926 (N_5926,N_2560,N_4325);
and U5927 (N_5927,N_1042,N_4840);
xor U5928 (N_5928,N_1961,N_1831);
nor U5929 (N_5929,N_168,N_3244);
or U5930 (N_5930,N_3933,N_2136);
xnor U5931 (N_5931,N_57,N_4248);
nand U5932 (N_5932,N_2836,N_918);
nand U5933 (N_5933,N_1100,N_894);
nand U5934 (N_5934,N_4500,N_4196);
and U5935 (N_5935,N_79,N_4125);
nand U5936 (N_5936,N_466,N_4692);
xnor U5937 (N_5937,N_764,N_1849);
nor U5938 (N_5938,N_3849,N_2050);
nor U5939 (N_5939,N_3517,N_636);
nand U5940 (N_5940,N_421,N_2312);
or U5941 (N_5941,N_1028,N_4104);
or U5942 (N_5942,N_4855,N_3823);
nand U5943 (N_5943,N_1350,N_3233);
or U5944 (N_5944,N_4784,N_1120);
or U5945 (N_5945,N_4242,N_2380);
nand U5946 (N_5946,N_3393,N_3057);
and U5947 (N_5947,N_3449,N_641);
nor U5948 (N_5948,N_1363,N_3358);
xor U5949 (N_5949,N_2191,N_3205);
nor U5950 (N_5950,N_3591,N_3755);
nand U5951 (N_5951,N_3079,N_237);
nand U5952 (N_5952,N_2264,N_2029);
xor U5953 (N_5953,N_2094,N_3072);
xnor U5954 (N_5954,N_4040,N_1134);
or U5955 (N_5955,N_3552,N_352);
and U5956 (N_5956,N_1680,N_3210);
and U5957 (N_5957,N_934,N_976);
or U5958 (N_5958,N_1622,N_1952);
nor U5959 (N_5959,N_1458,N_4043);
or U5960 (N_5960,N_4484,N_2210);
xor U5961 (N_5961,N_135,N_4694);
and U5962 (N_5962,N_3375,N_1866);
nor U5963 (N_5963,N_1840,N_4703);
xnor U5964 (N_5964,N_3108,N_4182);
and U5965 (N_5965,N_3153,N_243);
and U5966 (N_5966,N_4523,N_1658);
xnor U5967 (N_5967,N_3467,N_3496);
nand U5968 (N_5968,N_4366,N_2152);
xnor U5969 (N_5969,N_2792,N_4587);
or U5970 (N_5970,N_4108,N_1737);
or U5971 (N_5971,N_4310,N_4071);
xor U5972 (N_5972,N_2358,N_2232);
nor U5973 (N_5973,N_1790,N_71);
nor U5974 (N_5974,N_4351,N_3543);
xor U5975 (N_5975,N_4835,N_1920);
xor U5976 (N_5976,N_1058,N_4813);
nand U5977 (N_5977,N_2154,N_4915);
nand U5978 (N_5978,N_1034,N_612);
nand U5979 (N_5979,N_4318,N_3408);
and U5980 (N_5980,N_315,N_2065);
or U5981 (N_5981,N_4053,N_4326);
nor U5982 (N_5982,N_482,N_1841);
and U5983 (N_5983,N_335,N_3266);
nand U5984 (N_5984,N_813,N_4578);
nor U5985 (N_5985,N_1639,N_2498);
xor U5986 (N_5986,N_2031,N_1140);
nand U5987 (N_5987,N_4485,N_3219);
or U5988 (N_5988,N_1426,N_2674);
xnor U5989 (N_5989,N_8,N_680);
nor U5990 (N_5990,N_1676,N_2954);
or U5991 (N_5991,N_2192,N_4249);
xor U5992 (N_5992,N_2953,N_2689);
nor U5993 (N_5993,N_2826,N_2682);
and U5994 (N_5994,N_1630,N_471);
and U5995 (N_5995,N_3993,N_3556);
and U5996 (N_5996,N_3299,N_494);
nor U5997 (N_5997,N_4319,N_3593);
and U5998 (N_5998,N_1640,N_2738);
or U5999 (N_5999,N_831,N_3586);
and U6000 (N_6000,N_1534,N_4311);
and U6001 (N_6001,N_3446,N_2725);
or U6002 (N_6002,N_3148,N_4487);
nor U6003 (N_6003,N_4927,N_7);
and U6004 (N_6004,N_3470,N_4135);
nand U6005 (N_6005,N_1461,N_1722);
nand U6006 (N_6006,N_829,N_3022);
nand U6007 (N_6007,N_2586,N_4183);
or U6008 (N_6008,N_1573,N_2346);
and U6009 (N_6009,N_1029,N_4223);
xnor U6010 (N_6010,N_1019,N_3347);
and U6011 (N_6011,N_4615,N_655);
xor U6012 (N_6012,N_595,N_1906);
nand U6013 (N_6013,N_4445,N_3386);
and U6014 (N_6014,N_598,N_1322);
nor U6015 (N_6015,N_1648,N_3919);
nand U6016 (N_6016,N_184,N_1546);
and U6017 (N_6017,N_422,N_2385);
and U6018 (N_6018,N_1460,N_3439);
nand U6019 (N_6019,N_1269,N_4842);
xor U6020 (N_6020,N_1657,N_2680);
nand U6021 (N_6021,N_3603,N_3758);
and U6022 (N_6022,N_4823,N_2516);
nand U6023 (N_6023,N_3001,N_2799);
and U6024 (N_6024,N_2323,N_1523);
and U6025 (N_6025,N_2311,N_2020);
nor U6026 (N_6026,N_1620,N_1415);
nor U6027 (N_6027,N_459,N_3520);
nand U6028 (N_6028,N_630,N_2235);
nand U6029 (N_6029,N_4788,N_954);
or U6030 (N_6030,N_763,N_2010);
xnor U6031 (N_6031,N_1540,N_3221);
and U6032 (N_6032,N_746,N_358);
nand U6033 (N_6033,N_4243,N_2197);
and U6034 (N_6034,N_3418,N_4968);
or U6035 (N_6035,N_3278,N_2808);
nand U6036 (N_6036,N_4623,N_4450);
nand U6037 (N_6037,N_1497,N_274);
or U6038 (N_6038,N_3354,N_4192);
or U6039 (N_6039,N_715,N_658);
nand U6040 (N_6040,N_1846,N_1508);
nand U6041 (N_6041,N_4256,N_4388);
and U6042 (N_6042,N_3105,N_324);
or U6043 (N_6043,N_4103,N_1889);
or U6044 (N_6044,N_4145,N_1477);
nor U6045 (N_6045,N_1869,N_3401);
xnor U6046 (N_6046,N_2705,N_4806);
nand U6047 (N_6047,N_3139,N_416);
nor U6048 (N_6048,N_2933,N_863);
and U6049 (N_6049,N_2039,N_3396);
nor U6050 (N_6050,N_3923,N_4769);
nand U6051 (N_6051,N_2822,N_2153);
nand U6052 (N_6052,N_3170,N_2613);
xnor U6053 (N_6053,N_1285,N_4072);
nor U6054 (N_6054,N_2067,N_1038);
xnor U6055 (N_6055,N_2580,N_2696);
xor U6056 (N_6056,N_1731,N_3659);
and U6057 (N_6057,N_4115,N_30);
and U6058 (N_6058,N_4723,N_1548);
nor U6059 (N_6059,N_1214,N_2295);
xor U6060 (N_6060,N_2737,N_834);
and U6061 (N_6061,N_1443,N_183);
nand U6062 (N_6062,N_3061,N_2490);
nand U6063 (N_6063,N_3152,N_3699);
nand U6064 (N_6064,N_4305,N_2951);
nand U6065 (N_6065,N_804,N_1361);
or U6066 (N_6066,N_4858,N_3485);
nor U6067 (N_6067,N_563,N_585);
or U6068 (N_6068,N_3055,N_4453);
and U6069 (N_6069,N_1585,N_2641);
nor U6070 (N_6070,N_1762,N_3048);
nand U6071 (N_6071,N_2289,N_3766);
nor U6072 (N_6072,N_3722,N_1756);
or U6073 (N_6073,N_3817,N_735);
and U6074 (N_6074,N_3350,N_251);
nand U6075 (N_6075,N_637,N_662);
or U6076 (N_6076,N_4712,N_1513);
nor U6077 (N_6077,N_2134,N_2602);
or U6078 (N_6078,N_2772,N_4776);
or U6079 (N_6079,N_939,N_4186);
xnor U6080 (N_6080,N_4431,N_393);
xnor U6081 (N_6081,N_2379,N_2217);
xor U6082 (N_6082,N_4591,N_1098);
nor U6083 (N_6083,N_2546,N_2453);
nand U6084 (N_6084,N_3654,N_2246);
or U6085 (N_6085,N_4336,N_1817);
or U6086 (N_6086,N_1462,N_2113);
and U6087 (N_6087,N_4612,N_3649);
and U6088 (N_6088,N_1465,N_3960);
nand U6089 (N_6089,N_1716,N_35);
and U6090 (N_6090,N_622,N_1223);
and U6091 (N_6091,N_3829,N_255);
xor U6092 (N_6092,N_3222,N_1547);
or U6093 (N_6093,N_2750,N_1293);
nand U6094 (N_6094,N_3559,N_59);
xnor U6095 (N_6095,N_3639,N_2470);
or U6096 (N_6096,N_3860,N_4786);
nor U6097 (N_6097,N_4059,N_3335);
xnor U6098 (N_6098,N_4122,N_2128);
or U6099 (N_6099,N_1197,N_4410);
nand U6100 (N_6100,N_2417,N_3813);
or U6101 (N_6101,N_210,N_3725);
or U6102 (N_6102,N_2939,N_2824);
xor U6103 (N_6103,N_1659,N_1025);
nor U6104 (N_6104,N_1660,N_2749);
and U6105 (N_6105,N_4171,N_4988);
nor U6106 (N_6106,N_1187,N_4942);
nor U6107 (N_6107,N_1377,N_4208);
and U6108 (N_6108,N_2081,N_1061);
xnor U6109 (N_6109,N_2843,N_3038);
or U6110 (N_6110,N_2573,N_4568);
nand U6111 (N_6111,N_4791,N_4101);
or U6112 (N_6112,N_4754,N_826);
xnor U6113 (N_6113,N_2935,N_1604);
or U6114 (N_6114,N_1234,N_2394);
nor U6115 (N_6115,N_4140,N_3928);
nor U6116 (N_6116,N_461,N_2972);
and U6117 (N_6117,N_4376,N_4437);
or U6118 (N_6118,N_4283,N_4726);
and U6119 (N_6119,N_3296,N_3282);
or U6120 (N_6120,N_1156,N_3077);
nand U6121 (N_6121,N_381,N_4894);
or U6122 (N_6122,N_937,N_1811);
or U6123 (N_6123,N_760,N_1083);
and U6124 (N_6124,N_3748,N_3509);
or U6125 (N_6125,N_4387,N_1476);
xnor U6126 (N_6126,N_4717,N_4126);
nor U6127 (N_6127,N_1277,N_614);
nor U6128 (N_6128,N_3688,N_125);
or U6129 (N_6129,N_551,N_3320);
and U6130 (N_6130,N_3328,N_1510);
xor U6131 (N_6131,N_4441,N_4948);
nand U6132 (N_6132,N_417,N_1258);
or U6133 (N_6133,N_860,N_1951);
and U6134 (N_6134,N_4972,N_3653);
xnor U6135 (N_6135,N_2691,N_3071);
or U6136 (N_6136,N_2858,N_1965);
and U6137 (N_6137,N_1516,N_2719);
or U6138 (N_6138,N_3539,N_1656);
or U6139 (N_6139,N_1263,N_2455);
or U6140 (N_6140,N_2525,N_4328);
and U6141 (N_6141,N_3121,N_3971);
and U6142 (N_6142,N_1448,N_1091);
nand U6143 (N_6143,N_2244,N_3265);
or U6144 (N_6144,N_1827,N_327);
or U6145 (N_6145,N_1394,N_1536);
and U6146 (N_6146,N_2873,N_2934);
nor U6147 (N_6147,N_4272,N_1229);
and U6148 (N_6148,N_4165,N_4167);
xnor U6149 (N_6149,N_1045,N_340);
or U6150 (N_6150,N_2920,N_383);
or U6151 (N_6151,N_2003,N_1345);
or U6152 (N_6152,N_2995,N_4662);
or U6153 (N_6153,N_587,N_4009);
or U6154 (N_6154,N_3953,N_2628);
or U6155 (N_6155,N_2870,N_3814);
nand U6156 (N_6156,N_357,N_3113);
nand U6157 (N_6157,N_242,N_1518);
or U6158 (N_6158,N_1353,N_378);
nand U6159 (N_6159,N_1828,N_1289);
nand U6160 (N_6160,N_3950,N_811);
or U6161 (N_6161,N_2927,N_290);
or U6162 (N_6162,N_93,N_3565);
xnor U6163 (N_6163,N_3447,N_2224);
nor U6164 (N_6164,N_2021,N_1104);
and U6165 (N_6165,N_2997,N_4698);
and U6166 (N_6166,N_3100,N_2381);
xor U6167 (N_6167,N_123,N_4087);
nand U6168 (N_6168,N_2469,N_3602);
xnor U6169 (N_6169,N_3802,N_2848);
xor U6170 (N_6170,N_2267,N_3689);
or U6171 (N_6171,N_89,N_4133);
nor U6172 (N_6172,N_1777,N_2881);
nor U6173 (N_6173,N_3737,N_3974);
nand U6174 (N_6174,N_4089,N_2730);
nor U6175 (N_6175,N_2571,N_1887);
and U6176 (N_6176,N_1131,N_3237);
and U6177 (N_6177,N_367,N_3164);
and U6178 (N_6178,N_4780,N_1581);
nor U6179 (N_6179,N_4914,N_1191);
xor U6180 (N_6180,N_700,N_2980);
and U6181 (N_6181,N_145,N_229);
xor U6182 (N_6182,N_4301,N_2897);
xor U6183 (N_6183,N_4922,N_1598);
or U6184 (N_6184,N_4199,N_3853);
nand U6185 (N_6185,N_2091,N_3527);
or U6186 (N_6186,N_3007,N_2526);
nor U6187 (N_6187,N_1624,N_3658);
nand U6188 (N_6188,N_66,N_446);
nor U6189 (N_6189,N_759,N_2593);
nand U6190 (N_6190,N_534,N_1318);
nor U6191 (N_6191,N_1916,N_4766);
nand U6192 (N_6192,N_2384,N_69);
and U6193 (N_6193,N_713,N_1942);
xnor U6194 (N_6194,N_2388,N_2213);
and U6195 (N_6195,N_254,N_246);
xnor U6196 (N_6196,N_4094,N_3561);
and U6197 (N_6197,N_1692,N_2367);
or U6198 (N_6198,N_2468,N_2622);
nand U6199 (N_6199,N_915,N_4961);
nor U6200 (N_6200,N_3087,N_45);
or U6201 (N_6201,N_3585,N_80);
nand U6202 (N_6202,N_2281,N_3448);
xnor U6203 (N_6203,N_716,N_4585);
xor U6204 (N_6204,N_1115,N_3618);
nand U6205 (N_6205,N_1765,N_2774);
xnor U6206 (N_6206,N_2205,N_3039);
xor U6207 (N_6207,N_4926,N_1190);
nor U6208 (N_6208,N_3493,N_821);
xor U6209 (N_6209,N_3109,N_1873);
xnor U6210 (N_6210,N_4422,N_2273);
or U6211 (N_6211,N_1629,N_1945);
xnor U6212 (N_6212,N_4039,N_2966);
and U6213 (N_6213,N_693,N_4983);
nor U6214 (N_6214,N_3466,N_3788);
or U6215 (N_6215,N_329,N_1481);
nand U6216 (N_6216,N_449,N_1708);
and U6217 (N_6217,N_2720,N_2777);
or U6218 (N_6218,N_1259,N_4660);
xnor U6219 (N_6219,N_3062,N_1814);
xor U6220 (N_6220,N_1452,N_490);
and U6221 (N_6221,N_837,N_4714);
and U6222 (N_6222,N_3361,N_665);
xnor U6223 (N_6223,N_1627,N_4962);
nor U6224 (N_6224,N_3942,N_4284);
nor U6225 (N_6225,N_505,N_883);
and U6226 (N_6226,N_2706,N_4817);
nand U6227 (N_6227,N_4706,N_4442);
xnor U6228 (N_6228,N_2574,N_4689);
xor U6229 (N_6229,N_3762,N_4073);
and U6230 (N_6230,N_1773,N_1141);
and U6231 (N_6231,N_1677,N_781);
or U6232 (N_6232,N_1365,N_2028);
nor U6233 (N_6233,N_3628,N_4164);
and U6234 (N_6234,N_1647,N_2118);
nand U6235 (N_6235,N_2373,N_4241);
xor U6236 (N_6236,N_1123,N_236);
and U6237 (N_6237,N_3131,N_3478);
xnor U6238 (N_6238,N_1572,N_2183);
xor U6239 (N_6239,N_2483,N_2355);
nand U6240 (N_6240,N_2841,N_2633);
xnor U6241 (N_6241,N_4543,N_4137);
nor U6242 (N_6242,N_3761,N_2885);
nor U6243 (N_6243,N_240,N_855);
and U6244 (N_6244,N_1694,N_208);
nor U6245 (N_6245,N_3279,N_966);
xnor U6246 (N_6246,N_2566,N_4130);
and U6247 (N_6247,N_2649,N_4959);
nor U6248 (N_6248,N_3497,N_4992);
xnor U6249 (N_6249,N_1936,N_2548);
nand U6250 (N_6250,N_4590,N_3655);
xor U6251 (N_6251,N_4549,N_2400);
or U6252 (N_6252,N_4898,N_1740);
nand U6253 (N_6253,N_3935,N_4767);
xnor U6254 (N_6254,N_2442,N_814);
or U6255 (N_6255,N_4888,N_160);
and U6256 (N_6256,N_3554,N_272);
and U6257 (N_6257,N_3490,N_2006);
or U6258 (N_6258,N_547,N_1527);
and U6259 (N_6259,N_2909,N_2116);
and U6260 (N_6260,N_4076,N_593);
xnor U6261 (N_6261,N_260,N_2507);
xor U6262 (N_6262,N_1410,N_1155);
nor U6263 (N_6263,N_3193,N_4687);
nor U6264 (N_6264,N_960,N_2925);
and U6265 (N_6265,N_930,N_1087);
nand U6266 (N_6266,N_1766,N_1085);
xnor U6267 (N_6267,N_1317,N_3157);
and U6268 (N_6268,N_342,N_1432);
nand U6269 (N_6269,N_4225,N_4268);
nor U6270 (N_6270,N_2650,N_765);
nor U6271 (N_6271,N_1401,N_4488);
and U6272 (N_6272,N_562,N_756);
and U6273 (N_6273,N_3260,N_186);
xnor U6274 (N_6274,N_1686,N_2672);
or U6275 (N_6275,N_3248,N_4871);
nor U6276 (N_6276,N_4149,N_2314);
nand U6277 (N_6277,N_3532,N_3506);
nor U6278 (N_6278,N_4609,N_1280);
and U6279 (N_6279,N_2357,N_2788);
nor U6280 (N_6280,N_2850,N_1376);
or U6281 (N_6281,N_4333,N_1194);
nand U6282 (N_6282,N_3404,N_1144);
and U6283 (N_6283,N_3093,N_2514);
xor U6284 (N_6284,N_1056,N_4251);
xnor U6285 (N_6285,N_218,N_2971);
nand U6286 (N_6286,N_3179,N_3272);
or U6287 (N_6287,N_1275,N_1894);
nand U6288 (N_6288,N_1152,N_677);
nand U6289 (N_6289,N_3088,N_2129);
or U6290 (N_6290,N_2187,N_4664);
and U6291 (N_6291,N_868,N_2917);
xnor U6292 (N_6292,N_2803,N_3475);
nor U6293 (N_6293,N_166,N_2937);
xnor U6294 (N_6294,N_370,N_538);
xnor U6295 (N_6295,N_2626,N_3521);
and U6296 (N_6296,N_2418,N_2214);
and U6297 (N_6297,N_3518,N_539);
xnor U6298 (N_6298,N_163,N_3782);
and U6299 (N_6299,N_2448,N_728);
xor U6300 (N_6300,N_2778,N_2874);
or U6301 (N_6301,N_2206,N_2230);
nand U6302 (N_6302,N_1416,N_4421);
xor U6303 (N_6303,N_1533,N_4997);
nor U6304 (N_6304,N_456,N_1297);
and U6305 (N_6305,N_1266,N_2567);
nand U6306 (N_6306,N_3791,N_4051);
xnor U6307 (N_6307,N_1378,N_1008);
and U6308 (N_6308,N_4014,N_3843);
or U6309 (N_6309,N_24,N_2700);
nor U6310 (N_6310,N_2562,N_436);
xor U6311 (N_6311,N_2175,N_4371);
xnor U6312 (N_6312,N_4626,N_1133);
and U6313 (N_6313,N_188,N_3694);
or U6314 (N_6314,N_2186,N_2969);
or U6315 (N_6315,N_3304,N_1664);
xnor U6316 (N_6316,N_2208,N_366);
and U6317 (N_6317,N_3214,N_470);
and U6318 (N_6318,N_2386,N_143);
or U6319 (N_6319,N_2215,N_4899);
nand U6320 (N_6320,N_303,N_1932);
and U6321 (N_6321,N_4827,N_699);
nor U6322 (N_6322,N_2751,N_2679);
nand U6323 (N_6323,N_3877,N_2466);
or U6324 (N_6324,N_1979,N_2612);
xnor U6325 (N_6325,N_4763,N_3832);
nor U6326 (N_6326,N_2794,N_1937);
and U6327 (N_6327,N_2256,N_499);
or U6328 (N_6328,N_1212,N_2023);
nand U6329 (N_6329,N_3482,N_3947);
and U6330 (N_6330,N_2702,N_924);
and U6331 (N_6331,N_4818,N_4830);
nand U6332 (N_6332,N_10,N_2411);
and U6333 (N_6333,N_2298,N_157);
nand U6334 (N_6334,N_3534,N_1768);
and U6335 (N_6335,N_2008,N_4885);
xor U6336 (N_6336,N_1044,N_3997);
or U6337 (N_6337,N_1683,N_200);
or U6338 (N_6338,N_780,N_4987);
nor U6339 (N_6339,N_1742,N_3798);
nand U6340 (N_6340,N_2547,N_4181);
xor U6341 (N_6341,N_1721,N_2227);
xnor U6342 (N_6342,N_1283,N_858);
or U6343 (N_6343,N_3855,N_1690);
nand U6344 (N_6344,N_2374,N_120);
or U6345 (N_6345,N_2377,N_1049);
nor U6346 (N_6346,N_3502,N_213);
xnor U6347 (N_6347,N_913,N_455);
or U6348 (N_6348,N_3053,N_2163);
nor U6349 (N_6349,N_4822,N_1145);
xnor U6350 (N_6350,N_22,N_1875);
nand U6351 (N_6351,N_2432,N_1286);
nand U6352 (N_6352,N_3344,N_4919);
or U6353 (N_6353,N_4064,N_1610);
nor U6354 (N_6354,N_925,N_848);
and U6355 (N_6355,N_4497,N_4449);
nor U6356 (N_6356,N_1102,N_3249);
nand U6357 (N_6357,N_3580,N_336);
nor U6358 (N_6358,N_3486,N_2790);
nand U6359 (N_6359,N_2259,N_2627);
xor U6360 (N_6360,N_109,N_4166);
nor U6361 (N_6361,N_2356,N_2022);
nor U6362 (N_6362,N_884,N_4649);
and U6363 (N_6363,N_4677,N_3666);
nor U6364 (N_6364,N_3481,N_2199);
nor U6365 (N_6365,N_2445,N_1950);
or U6366 (N_6366,N_1596,N_4538);
or U6367 (N_6367,N_1792,N_3765);
xnor U6368 (N_6368,N_1964,N_4489);
nor U6369 (N_6369,N_2422,N_1354);
or U6370 (N_6370,N_205,N_300);
or U6371 (N_6371,N_2099,N_613);
nor U6372 (N_6372,N_1484,N_4691);
nor U6373 (N_6373,N_1182,N_3332);
xor U6374 (N_6374,N_2467,N_796);
or U6375 (N_6375,N_2820,N_2973);
or U6376 (N_6376,N_1442,N_2368);
nor U6377 (N_6377,N_4277,N_3759);
and U6378 (N_6378,N_2664,N_2063);
nor U6379 (N_6379,N_4179,N_4394);
or U6380 (N_6380,N_3444,N_4377);
or U6381 (N_6381,N_3774,N_1062);
xor U6382 (N_6382,N_3742,N_1200);
or U6383 (N_6383,N_3512,N_2632);
and U6384 (N_6384,N_1201,N_337);
or U6385 (N_6385,N_1108,N_2062);
and U6386 (N_6386,N_3785,N_504);
nor U6387 (N_6387,N_1696,N_433);
nand U6388 (N_6388,N_2697,N_296);
and U6389 (N_6389,N_364,N_2149);
nand U6390 (N_6390,N_2932,N_4834);
and U6391 (N_6391,N_2488,N_647);
nor U6392 (N_6392,N_3454,N_3231);
xor U6393 (N_6393,N_4752,N_4414);
nand U6394 (N_6394,N_1824,N_990);
or U6395 (N_6395,N_2446,N_278);
nor U6396 (N_6396,N_4826,N_982);
nor U6397 (N_6397,N_4042,N_878);
and U6398 (N_6398,N_683,N_122);
or U6399 (N_6399,N_1252,N_4361);
and U6400 (N_6400,N_3716,N_390);
or U6401 (N_6401,N_380,N_4270);
and U6402 (N_6402,N_47,N_2080);
nand U6403 (N_6403,N_3885,N_544);
nand U6404 (N_6404,N_3283,N_1440);
xor U6405 (N_6405,N_4866,N_2588);
and U6406 (N_6406,N_3413,N_3187);
nor U6407 (N_6407,N_1972,N_161);
or U6408 (N_6408,N_51,N_3066);
nor U6409 (N_6409,N_4928,N_2856);
or U6410 (N_6410,N_3623,N_2656);
nand U6411 (N_6411,N_4416,N_2596);
xnor U6412 (N_6412,N_2123,N_3815);
nand U6413 (N_6413,N_72,N_4833);
xor U6414 (N_6414,N_2284,N_3104);
or U6415 (N_6415,N_4918,N_4592);
or U6416 (N_6416,N_4571,N_2200);
nor U6417 (N_6417,N_4675,N_1453);
nand U6418 (N_6418,N_1905,N_3710);
nand U6419 (N_6419,N_1173,N_2763);
and U6420 (N_6420,N_1012,N_4373);
xnor U6421 (N_6421,N_1892,N_4131);
xor U6422 (N_6422,N_4069,N_599);
nor U6423 (N_6423,N_3422,N_226);
xor U6424 (N_6424,N_4480,N_2399);
or U6425 (N_6425,N_961,N_2872);
or U6426 (N_6426,N_2747,N_4676);
xor U6427 (N_6427,N_3790,N_2305);
xnor U6428 (N_6428,N_3535,N_4588);
nor U6429 (N_6429,N_3582,N_3476);
nand U6430 (N_6430,N_3368,N_283);
xnor U6431 (N_6431,N_4176,N_644);
xnor U6432 (N_6432,N_2125,N_4246);
and U6433 (N_6433,N_4976,N_85);
nand U6434 (N_6434,N_164,N_233);
nor U6435 (N_6435,N_4293,N_4665);
nor U6436 (N_6436,N_3650,N_3674);
nor U6437 (N_6437,N_3357,N_1256);
xnor U6438 (N_6438,N_2722,N_2);
xor U6439 (N_6439,N_1986,N_3932);
and U6440 (N_6440,N_1287,N_2287);
or U6441 (N_6441,N_4846,N_2083);
and U6442 (N_6442,N_2132,N_147);
or U6443 (N_6443,N_31,N_1067);
nor U6444 (N_6444,N_2181,N_1021);
or U6445 (N_6445,N_2223,N_3703);
nand U6446 (N_6446,N_3302,N_501);
and U6447 (N_6447,N_1669,N_2745);
or U6448 (N_6448,N_1146,N_2451);
xnor U6449 (N_6449,N_3624,N_1329);
nor U6450 (N_6450,N_4627,N_3968);
or U6451 (N_6451,N_4338,N_438);
and U6452 (N_6452,N_1542,N_775);
nand U6453 (N_6453,N_3844,N_4300);
xor U6454 (N_6454,N_4913,N_1192);
or U6455 (N_6455,N_83,N_2524);
or U6456 (N_6456,N_2414,N_4321);
xnor U6457 (N_6457,N_1290,N_729);
and U6458 (N_6458,N_1313,N_4157);
or U6459 (N_6459,N_2655,N_2069);
xnor U6460 (N_6460,N_3750,N_1987);
nor U6461 (N_6461,N_2828,N_3381);
and U6462 (N_6462,N_3848,N_926);
xnor U6463 (N_6463,N_2307,N_3252);
nor U6464 (N_6464,N_4331,N_1367);
nor U6465 (N_6465,N_136,N_414);
or U6466 (N_6466,N_1105,N_4757);
nand U6467 (N_6467,N_3437,N_2343);
xor U6468 (N_6468,N_3215,N_2736);
nand U6469 (N_6469,N_2372,N_1888);
and U6470 (N_6470,N_4690,N_2987);
nor U6471 (N_6471,N_3872,N_3880);
xor U6472 (N_6472,N_4957,N_4800);
xnor U6473 (N_6473,N_4290,N_2452);
and U6474 (N_6474,N_2426,N_3851);
and U6475 (N_6475,N_559,N_891);
nand U6476 (N_6476,N_2922,N_4908);
nor U6477 (N_6477,N_12,N_1751);
xnor U6478 (N_6478,N_2888,N_2330);
and U6479 (N_6479,N_1472,N_1857);
xor U6480 (N_6480,N_1678,N_285);
nand U6481 (N_6481,N_1645,N_4879);
and U6482 (N_6482,N_3461,N_3838);
or U6483 (N_6483,N_769,N_1561);
nand U6484 (N_6484,N_1143,N_2485);
xor U6485 (N_6485,N_1797,N_2496);
xnor U6486 (N_6486,N_4725,N_2531);
nand U6487 (N_6487,N_4739,N_2515);
and U6488 (N_6488,N_94,N_1276);
and U6489 (N_6489,N_3142,N_3041);
or U6490 (N_6490,N_4639,N_3901);
xor U6491 (N_6491,N_2409,N_4032);
and U6492 (N_6492,N_3811,N_3186);
or U6493 (N_6493,N_2319,N_3199);
nand U6494 (N_6494,N_1558,N_3181);
and U6495 (N_6495,N_486,N_2804);
or U6496 (N_6496,N_2216,N_4314);
nand U6497 (N_6497,N_4567,N_2085);
nor U6498 (N_6498,N_1565,N_1632);
or U6499 (N_6499,N_3764,N_917);
and U6500 (N_6500,N_577,N_1579);
or U6501 (N_6501,N_4929,N_2640);
nor U6502 (N_6502,N_2582,N_696);
and U6503 (N_6503,N_1040,N_1064);
nand U6504 (N_6504,N_4709,N_1217);
nand U6505 (N_6505,N_4458,N_121);
nor U6506 (N_6506,N_1709,N_619);
or U6507 (N_6507,N_895,N_408);
nand U6508 (N_6508,N_2127,N_1128);
nand U6509 (N_6509,N_4820,N_3026);
nor U6510 (N_6510,N_3013,N_1157);
nor U6511 (N_6511,N_2758,N_1488);
xnor U6512 (N_6512,N_993,N_3776);
nor U6513 (N_6513,N_1457,N_3084);
xor U6514 (N_6514,N_2068,N_2857);
xor U6515 (N_6515,N_1668,N_4124);
or U6516 (N_6516,N_3294,N_4986);
nor U6517 (N_6517,N_791,N_3389);
or U6518 (N_6518,N_220,N_2260);
nor U6519 (N_6519,N_3718,N_1024);
nand U6520 (N_6520,N_3882,N_3070);
nor U6521 (N_6521,N_2242,N_3155);
nor U6522 (N_6522,N_388,N_467);
and U6523 (N_6523,N_4613,N_3955);
nor U6524 (N_6524,N_3573,N_137);
and U6525 (N_6525,N_3711,N_3682);
nor U6526 (N_6526,N_2523,N_3107);
xor U6527 (N_6527,N_575,N_3036);
and U6528 (N_6528,N_343,N_1977);
or U6529 (N_6529,N_3921,N_4228);
xor U6530 (N_6530,N_2383,N_673);
and U6531 (N_6531,N_4859,N_48);
xnor U6532 (N_6532,N_1439,N_4294);
or U6533 (N_6533,N_1163,N_3099);
xor U6534 (N_6534,N_1679,N_2581);
nand U6535 (N_6535,N_1323,N_1597);
nand U6536 (N_6536,N_3464,N_2876);
nor U6537 (N_6537,N_3117,N_2104);
or U6538 (N_6538,N_3822,N_1057);
xnor U6539 (N_6539,N_4440,N_479);
nand U6540 (N_6540,N_2544,N_4401);
and U6541 (N_6541,N_3337,N_4635);
or U6542 (N_6542,N_2437,N_4873);
nand U6543 (N_6543,N_2285,N_2982);
nand U6544 (N_6544,N_653,N_958);
or U6545 (N_6545,N_1242,N_2253);
nand U6546 (N_6546,N_1065,N_4998);
nor U6547 (N_6547,N_3120,N_3023);
and U6548 (N_6548,N_2714,N_4574);
xnor U6549 (N_6549,N_151,N_566);
nor U6550 (N_6550,N_3005,N_3159);
nor U6551 (N_6551,N_4857,N_1060);
and U6552 (N_6552,N_2625,N_2164);
or U6553 (N_6553,N_1907,N_2683);
nand U6554 (N_6554,N_634,N_3274);
nand U6555 (N_6555,N_3144,N_3679);
and U6556 (N_6556,N_2282,N_3116);
and U6557 (N_6557,N_911,N_2983);
and U6558 (N_6558,N_4077,N_4647);
or U6559 (N_6559,N_704,N_4423);
nand U6560 (N_6560,N_1789,N_3903);
and U6561 (N_6561,N_2477,N_1898);
or U6562 (N_6562,N_284,N_2663);
and U6563 (N_6563,N_2781,N_3016);
and U6564 (N_6564,N_3238,N_2389);
nor U6565 (N_6565,N_1002,N_4313);
xnor U6566 (N_6566,N_885,N_1667);
or U6567 (N_6567,N_3010,N_2797);
nor U6568 (N_6568,N_3505,N_1637);
and U6569 (N_6569,N_4426,N_1421);
nor U6570 (N_6570,N_2859,N_2837);
and U6571 (N_6571,N_1284,N_4447);
and U6572 (N_6572,N_271,N_2867);
or U6573 (N_6573,N_4037,N_1904);
xor U6574 (N_6574,N_758,N_3560);
or U6575 (N_6575,N_4408,N_1047);
and U6576 (N_6576,N_3380,N_1556);
nor U6577 (N_6577,N_1395,N_1216);
xnor U6578 (N_6578,N_3343,N_3789);
nor U6579 (N_6579,N_4550,N_2408);
xor U6580 (N_6580,N_1746,N_305);
nand U6581 (N_6581,N_2294,N_3074);
nand U6582 (N_6582,N_4263,N_3040);
or U6583 (N_6583,N_4054,N_1227);
xor U6584 (N_6584,N_4028,N_298);
and U6585 (N_6585,N_4308,N_1929);
xnor U6586 (N_6586,N_1370,N_4748);
and U6587 (N_6587,N_1741,N_3003);
xnor U6588 (N_6588,N_3111,N_4584);
nor U6589 (N_6589,N_1137,N_685);
and U6590 (N_6590,N_165,N_2665);
or U6591 (N_6591,N_3236,N_4470);
nand U6592 (N_6592,N_3259,N_3909);
nand U6593 (N_6593,N_888,N_4520);
nand U6594 (N_6594,N_1427,N_4522);
nand U6595 (N_6595,N_463,N_1578);
nand U6596 (N_6596,N_454,N_1383);
xor U6597 (N_6597,N_484,N_430);
xor U6598 (N_6598,N_3191,N_3209);
or U6599 (N_6599,N_3334,N_4736);
nand U6600 (N_6600,N_3340,N_2900);
nand U6601 (N_6601,N_4559,N_617);
and U6602 (N_6602,N_2860,N_331);
nand U6603 (N_6603,N_2014,N_1912);
nor U6604 (N_6604,N_1787,N_4905);
xor U6605 (N_6605,N_4999,N_2880);
xnor U6606 (N_6606,N_4491,N_1470);
or U6607 (N_6607,N_4632,N_2816);
xnor U6608 (N_6608,N_3962,N_1447);
nand U6609 (N_6609,N_4785,N_4996);
or U6610 (N_6610,N_1730,N_1441);
nor U6611 (N_6611,N_4382,N_517);
or U6612 (N_6612,N_675,N_2218);
xor U6613 (N_6613,N_4061,N_3000);
nor U6614 (N_6614,N_2245,N_903);
nor U6615 (N_6615,N_4399,N_1782);
xnor U6616 (N_6616,N_3384,N_4656);
nand U6617 (N_6617,N_604,N_1271);
nor U6618 (N_6618,N_817,N_385);
xnor U6619 (N_6619,N_4038,N_849);
and U6620 (N_6620,N_4012,N_1097);
xnor U6621 (N_6621,N_3290,N_2353);
or U6622 (N_6622,N_4494,N_2977);
and U6623 (N_6623,N_4648,N_3589);
xor U6624 (N_6624,N_451,N_2504);
nor U6625 (N_6625,N_3054,N_2694);
and U6626 (N_6626,N_4930,N_2924);
and U6627 (N_6627,N_3546,N_4904);
nand U6628 (N_6628,N_3192,N_4730);
nand U6629 (N_6629,N_1166,N_1172);
xor U6630 (N_6630,N_2793,N_4956);
or U6631 (N_6631,N_4083,N_3797);
nor U6632 (N_6632,N_4851,N_1877);
or U6633 (N_6633,N_2103,N_1980);
or U6634 (N_6634,N_420,N_199);
and U6635 (N_6635,N_1655,N_88);
or U6636 (N_6636,N_4575,N_2241);
and U6637 (N_6637,N_1901,N_3516);
or U6638 (N_6638,N_2907,N_339);
nor U6639 (N_6639,N_4577,N_2861);
nor U6640 (N_6640,N_193,N_1507);
and U6641 (N_6641,N_4541,N_3284);
nor U6642 (N_6642,N_2819,N_4383);
xor U6643 (N_6643,N_3021,N_4507);
or U6644 (N_6644,N_4255,N_800);
and U6645 (N_6645,N_3406,N_2474);
nor U6646 (N_6646,N_3339,N_1593);
or U6647 (N_6647,N_204,N_2486);
xor U6648 (N_6648,N_91,N_4886);
and U6649 (N_6649,N_4424,N_974);
nor U6650 (N_6650,N_2489,N_159);
xnor U6651 (N_6651,N_1039,N_310);
and U6652 (N_6652,N_1463,N_4116);
or U6653 (N_6653,N_4029,N_1734);
and U6654 (N_6654,N_2754,N_1054);
and U6655 (N_6655,N_3662,N_341);
xor U6656 (N_6656,N_4582,N_2654);
nand U6657 (N_6657,N_1385,N_4510);
nand U6658 (N_6658,N_3425,N_174);
and U6659 (N_6659,N_3182,N_313);
nand U6660 (N_6660,N_3768,N_3398);
nand U6661 (N_6661,N_2530,N_4853);
xor U6662 (N_6662,N_4877,N_3101);
and U6663 (N_6663,N_4023,N_1752);
nand U6664 (N_6664,N_1537,N_2449);
or U6665 (N_6665,N_3140,N_3876);
nand U6666 (N_6666,N_4438,N_4404);
or U6667 (N_6667,N_98,N_2151);
nor U6668 (N_6668,N_4678,N_970);
and U6669 (N_6669,N_642,N_3912);
nor U6670 (N_6670,N_1411,N_4747);
xor U6671 (N_6671,N_2796,N_1796);
nor U6672 (N_6672,N_78,N_1202);
xnor U6673 (N_6673,N_3956,N_4499);
nor U6674 (N_6674,N_4175,N_3781);
or U6675 (N_6675,N_3705,N_4052);
nor U6676 (N_6676,N_4324,N_3472);
and U6677 (N_6677,N_4895,N_2535);
and U6678 (N_6678,N_3878,N_2429);
nor U6679 (N_6679,N_2501,N_3833);
nor U6680 (N_6680,N_1159,N_1428);
nor U6681 (N_6681,N_4593,N_2832);
nor U6682 (N_6682,N_3819,N_3732);
xnor U6683 (N_6683,N_2609,N_4309);
xor U6684 (N_6684,N_3696,N_4257);
xor U6685 (N_6685,N_1041,N_289);
and U6686 (N_6686,N_3261,N_2519);
or U6687 (N_6687,N_1438,N_1139);
or U6688 (N_6688,N_1687,N_4870);
nand U6689 (N_6689,N_3452,N_418);
and U6690 (N_6690,N_537,N_1298);
xnor U6691 (N_6691,N_594,N_4281);
nand U6692 (N_6692,N_4266,N_940);
and U6693 (N_6693,N_812,N_572);
and U6694 (N_6694,N_709,N_1204);
xor U6695 (N_6695,N_253,N_447);
or U6696 (N_6696,N_2537,N_509);
or U6697 (N_6697,N_3999,N_4195);
xnor U6698 (N_6698,N_2236,N_3349);
xnor U6699 (N_6699,N_1168,N_927);
nor U6700 (N_6700,N_3537,N_1109);
and U6701 (N_6701,N_1178,N_2645);
and U6702 (N_6702,N_1911,N_1059);
xnor U6703 (N_6703,N_2952,N_4327);
or U6704 (N_6704,N_3934,N_2989);
xor U6705 (N_6705,N_920,N_2403);
and U6706 (N_6706,N_1591,N_535);
and U6707 (N_6707,N_2978,N_877);
and U6708 (N_6708,N_4674,N_4641);
and U6709 (N_6709,N_1611,N_589);
and U6710 (N_6710,N_321,N_3842);
xor U6711 (N_6711,N_302,N_4235);
nand U6712 (N_6712,N_1539,N_3457);
nand U6713 (N_6713,N_705,N_3267);
xor U6714 (N_6714,N_3488,N_4563);
or U6715 (N_6715,N_1320,N_4900);
xnor U6716 (N_6716,N_1449,N_1998);
or U6717 (N_6717,N_1393,N_736);
or U6718 (N_6718,N_405,N_4102);
xnor U6719 (N_6719,N_1196,N_833);
nor U6720 (N_6720,N_4524,N_2561);
nand U6721 (N_6721,N_1727,N_1485);
nor U6722 (N_6722,N_1935,N_4661);
nor U6723 (N_6723,N_33,N_3598);
or U6724 (N_6724,N_2949,N_1380);
or U6725 (N_6725,N_2491,N_2098);
xor U6726 (N_6726,N_3983,N_4132);
xnor U6727 (N_6727,N_2463,N_1823);
xnor U6728 (N_6728,N_4163,N_3590);
and U6729 (N_6729,N_99,N_1861);
and U6730 (N_6730,N_2930,N_2928);
nor U6731 (N_6731,N_4527,N_96);
nor U6732 (N_6732,N_1466,N_1626);
xor U6733 (N_6733,N_4887,N_2212);
and U6734 (N_6734,N_1078,N_4047);
nor U6735 (N_6735,N_3695,N_2000);
nand U6736 (N_6736,N_2955,N_1674);
nor U6737 (N_6737,N_3065,N_1883);
or U6738 (N_6738,N_1876,N_1628);
or U6739 (N_6739,N_3917,N_2784);
xnor U6740 (N_6740,N_4770,N_2348);
nor U6741 (N_6741,N_3161,N_4216);
or U6742 (N_6742,N_1122,N_1208);
or U6743 (N_6743,N_2563,N_3884);
nand U6744 (N_6744,N_2410,N_2109);
nor U6745 (N_6745,N_4349,N_1112);
nor U6746 (N_6746,N_4845,N_412);
nand U6747 (N_6747,N_3841,N_2717);
xnor U6748 (N_6748,N_4105,N_2892);
xnor U6749 (N_6749,N_4938,N_2487);
nor U6750 (N_6750,N_2759,N_767);
xnor U6751 (N_6751,N_718,N_2770);
or U6752 (N_6752,N_2505,N_778);
and U6753 (N_6753,N_1066,N_308);
xor U6754 (N_6754,N_4380,N_2965);
or U6755 (N_6755,N_624,N_4091);
nor U6756 (N_6756,N_1215,N_2017);
xor U6757 (N_6757,N_2051,N_4950);
or U6758 (N_6758,N_1799,N_4920);
xnor U6759 (N_6759,N_3806,N_3223);
nor U6760 (N_6760,N_1124,N_2741);
and U6761 (N_6761,N_2500,N_2943);
nand U6762 (N_6762,N_1688,N_4278);
or U6763 (N_6763,N_261,N_322);
or U6764 (N_6764,N_4755,N_4891);
nor U6765 (N_6765,N_3592,N_1592);
nor U6766 (N_6766,N_660,N_1324);
xnor U6767 (N_6767,N_4050,N_3307);
xor U6768 (N_6768,N_1689,N_3991);
or U6769 (N_6769,N_1816,N_1473);
and U6770 (N_6770,N_3433,N_2764);
xor U6771 (N_6771,N_906,N_95);
xor U6772 (N_6772,N_2552,N_2818);
or U6773 (N_6773,N_2988,N_3218);
nor U6774 (N_6774,N_949,N_2866);
and U6775 (N_6775,N_2404,N_3826);
nor U6776 (N_6776,N_523,N_4066);
nand U6777 (N_6777,N_1890,N_3239);
nor U6778 (N_6778,N_969,N_1526);
and U6779 (N_6779,N_1804,N_70);
nor U6780 (N_6780,N_2424,N_3620);
nor U6781 (N_6781,N_2522,N_1729);
nor U6782 (N_6782,N_3385,N_3975);
nand U6783 (N_6783,N_2901,N_432);
xor U6784 (N_6784,N_2991,N_1946);
nand U6785 (N_6785,N_3431,N_3510);
nor U6786 (N_6786,N_3615,N_1020);
nor U6787 (N_6787,N_3676,N_3430);
and U6788 (N_6788,N_3577,N_3081);
and U6789 (N_6789,N_3836,N_435);
or U6790 (N_6790,N_1743,N_2898);
and U6791 (N_6791,N_1262,N_670);
nor U6792 (N_6792,N_3595,N_2711);
nor U6793 (N_6793,N_3892,N_3050);
xor U6794 (N_6794,N_2752,N_2662);
nor U6795 (N_6795,N_2335,N_115);
nor U6796 (N_6796,N_3514,N_1896);
and U6797 (N_6797,N_1880,N_2975);
nand U6798 (N_6798,N_1843,N_3979);
and U6799 (N_6799,N_2776,N_2481);
nand U6800 (N_6800,N_583,N_3786);
or U6801 (N_6801,N_1296,N_105);
or U6802 (N_6802,N_1807,N_2729);
xnor U6803 (N_6803,N_3373,N_4172);
nor U6804 (N_6804,N_224,N_1865);
and U6805 (N_6805,N_458,N_676);
nand U6806 (N_6806,N_440,N_2092);
or U6807 (N_6807,N_4239,N_555);
xnor U6808 (N_6808,N_1106,N_462);
nor U6809 (N_6809,N_333,N_3994);
and U6810 (N_6810,N_2964,N_2059);
and U6811 (N_6811,N_1077,N_3594);
or U6812 (N_6812,N_4018,N_774);
or U6813 (N_6813,N_3910,N_4831);
nand U6814 (N_6814,N_681,N_1665);
nand U6815 (N_6815,N_2998,N_1666);
and U6816 (N_6816,N_2220,N_148);
nand U6817 (N_6817,N_2359,N_1736);
or U6818 (N_6818,N_650,N_2048);
or U6819 (N_6819,N_1429,N_108);
nand U6820 (N_6820,N_2161,N_399);
xnor U6821 (N_6821,N_3924,N_2147);
nor U6822 (N_6822,N_793,N_264);
nor U6823 (N_6823,N_4854,N_4279);
and U6824 (N_6824,N_3741,N_1158);
nor U6825 (N_6825,N_1532,N_307);
xor U6826 (N_6826,N_4809,N_1992);
nor U6827 (N_6827,N_859,N_1981);
or U6828 (N_6828,N_3690,N_4759);
nand U6829 (N_6829,N_879,N_846);
nand U6830 (N_6830,N_201,N_3989);
xnor U6831 (N_6831,N_2261,N_319);
and U6832 (N_6832,N_4365,N_2780);
or U6833 (N_6833,N_3648,N_3896);
and U6834 (N_6834,N_1895,N_4291);
xnor U6835 (N_6835,N_4403,N_3058);
xor U6836 (N_6836,N_1820,N_4655);
xor U6837 (N_6837,N_3952,N_2631);
and U6838 (N_6838,N_4946,N_4006);
xnor U6839 (N_6839,N_2709,N_171);
and U6840 (N_6840,N_688,N_2270);
nor U6841 (N_6841,N_2895,N_189);
or U6842 (N_6842,N_282,N_526);
xnor U6843 (N_6843,N_275,N_4046);
nor U6844 (N_6844,N_2046,N_2834);
xor U6845 (N_6845,N_3686,N_3032);
or U6846 (N_6846,N_4407,N_1673);
nand U6847 (N_6847,N_4454,N_4876);
or U6848 (N_6848,N_580,N_4715);
nand U6849 (N_6849,N_1444,N_1559);
xor U6850 (N_6850,N_1870,N_2443);
xor U6851 (N_6851,N_1704,N_2176);
nand U6852 (N_6852,N_3625,N_1150);
and U6853 (N_6853,N_2570,N_3429);
and U6854 (N_6854,N_4187,N_3687);
nand U6855 (N_6855,N_597,N_4425);
nor U6856 (N_6856,N_1371,N_531);
nor U6857 (N_6857,N_1068,N_805);
xor U6858 (N_6858,N_266,N_2097);
xnor U6859 (N_6859,N_2042,N_3314);
or U6860 (N_6860,N_854,N_1919);
xor U6861 (N_6861,N_1939,N_1349);
xor U6862 (N_6862,N_182,N_1101);
or U6863 (N_6863,N_2825,N_3145);
nand U6864 (N_6864,N_2815,N_3837);
and U6865 (N_6865,N_2079,N_3779);
xor U6866 (N_6866,N_3046,N_3366);
and U6867 (N_6867,N_4253,N_4554);
nor U6868 (N_6868,N_2948,N_965);
xor U6869 (N_6869,N_1046,N_1781);
nand U6870 (N_6870,N_1544,N_2096);
and U6871 (N_6871,N_3492,N_1761);
and U6872 (N_6872,N_2102,N_623);
nand U6873 (N_6873,N_32,N_395);
nand U6874 (N_6874,N_1036,N_2636);
nor U6875 (N_6875,N_4139,N_1434);
nor U6876 (N_6876,N_3241,N_1783);
nor U6877 (N_6877,N_789,N_649);
or U6878 (N_6878,N_2228,N_3156);
nor U6879 (N_6879,N_2250,N_4417);
nand U6880 (N_6880,N_1803,N_2755);
and U6881 (N_6881,N_4558,N_567);
and U6882 (N_6882,N_249,N_3348);
xnor U6883 (N_6883,N_841,N_1908);
nor U6884 (N_6884,N_1341,N_690);
or U6885 (N_6885,N_4428,N_2196);
xnor U6886 (N_6886,N_638,N_2618);
and U6887 (N_6887,N_437,N_3453);
and U6888 (N_6888,N_691,N_3728);
nand U6889 (N_6889,N_351,N_2087);
nand U6890 (N_6890,N_890,N_4495);
nor U6891 (N_6891,N_3825,N_4397);
nor U6892 (N_6892,N_1346,N_3970);
or U6893 (N_6893,N_3760,N_2509);
and U6894 (N_6894,N_3377,N_346);
nand U6895 (N_6895,N_3839,N_4734);
or U6896 (N_6896,N_1684,N_1013);
nor U6897 (N_6897,N_4307,N_2120);
and U6898 (N_6898,N_1703,N_4685);
and U6899 (N_6899,N_3275,N_3308);
and U6900 (N_6900,N_4036,N_2145);
and U6901 (N_6901,N_1671,N_1183);
nor U6902 (N_6902,N_1599,N_3946);
or U6903 (N_6903,N_659,N_3807);
and U6904 (N_6904,N_1851,N_3034);
or U6905 (N_6905,N_1490,N_3622);
nor U6906 (N_6906,N_4688,N_3494);
nor U6907 (N_6907,N_4238,N_2812);
or U6908 (N_6908,N_2541,N_1352);
nand U6909 (N_6909,N_2517,N_2579);
and U6910 (N_6910,N_771,N_3364);
nor U6911 (N_6911,N_2047,N_1614);
xor U6912 (N_6912,N_3927,N_350);
or U6913 (N_6913,N_119,N_1549);
or U6914 (N_6914,N_1826,N_4189);
nand U6915 (N_6915,N_3491,N_3394);
nand U6916 (N_6916,N_1955,N_4044);
xnor U6917 (N_6917,N_608,N_1149);
and U6918 (N_6918,N_1491,N_3904);
nand U6919 (N_6919,N_1151,N_2479);
and U6920 (N_6920,N_874,N_3247);
xnor U6921 (N_6921,N_4945,N_782);
nand U6922 (N_6922,N_3772,N_2115);
xor U6923 (N_6923,N_2743,N_4596);
nand U6924 (N_6924,N_4154,N_1958);
xor U6925 (N_6925,N_1995,N_777);
and U6926 (N_6926,N_3500,N_1089);
nand U6927 (N_6927,N_1093,N_106);
xor U6928 (N_6928,N_1748,N_4320);
nor U6929 (N_6929,N_511,N_3604);
xnor U6930 (N_6930,N_4711,N_5);
and U6931 (N_6931,N_1422,N_3271);
or U6932 (N_6932,N_3370,N_3250);
nor U6933 (N_6933,N_4634,N_4213);
xnor U6934 (N_6934,N_4509,N_469);
nand U6935 (N_6935,N_6,N_2322);
nand U6936 (N_6936,N_798,N_3608);
nand U6937 (N_6937,N_3850,N_3611);
xnor U6938 (N_6938,N_3076,N_453);
and U6939 (N_6939,N_2440,N_104);
or U6940 (N_6940,N_2121,N_4411);
or U6941 (N_6941,N_3504,N_3926);
nor U6942 (N_6942,N_2229,N_2462);
nor U6943 (N_6943,N_2137,N_4753);
and U6944 (N_6944,N_4967,N_1211);
or U6945 (N_6945,N_1661,N_1587);
nor U6946 (N_6946,N_1372,N_3207);
and U6947 (N_6947,N_3160,N_3938);
nor U6948 (N_6948,N_4630,N_4004);
and U6949 (N_6949,N_4231,N_2233);
nor U6950 (N_6950,N_353,N_4802);
nand U6951 (N_6951,N_4147,N_110);
xnor U6952 (N_6952,N_3681,N_1574);
nor U6953 (N_6953,N_1496,N_3865);
xor U6954 (N_6954,N_2610,N_1638);
and U6955 (N_6955,N_409,N_3526);
nor U6956 (N_6956,N_1662,N_4363);
nor U6957 (N_6957,N_1772,N_1948);
or U6958 (N_6958,N_1125,N_2528);
and U6959 (N_6959,N_651,N_1634);
xnor U6960 (N_6960,N_3060,N_3141);
or U6961 (N_6961,N_2362,N_666);
or U6962 (N_6962,N_950,N_4143);
or U6963 (N_6963,N_2865,N_4155);
xnor U6964 (N_6964,N_1220,N_514);
nand U6965 (N_6965,N_452,N_870);
nor U6966 (N_6966,N_3277,N_4501);
nor U6967 (N_6967,N_4107,N_1226);
xnor U6968 (N_6968,N_2302,N_1538);
nor U6969 (N_6969,N_4240,N_1379);
and U6970 (N_6970,N_2465,N_3664);
xor U6971 (N_6971,N_4013,N_3671);
nor U6972 (N_6972,N_4576,N_3873);
xor U6973 (N_6973,N_4799,N_4473);
nor U6974 (N_6974,N_4610,N_2617);
nand U6975 (N_6975,N_971,N_4477);
xor U6976 (N_6976,N_1822,N_4357);
or U6977 (N_6977,N_1607,N_4027);
and U6978 (N_6978,N_4118,N_4220);
nor U6979 (N_6979,N_1011,N_372);
and U6980 (N_6980,N_4949,N_524);
nand U6981 (N_6981,N_4940,N_1956);
xor U6982 (N_6982,N_502,N_4475);
or U6983 (N_6983,N_3262,N_3700);
and U6984 (N_6984,N_4995,N_947);
nor U6985 (N_6985,N_2913,N_2413);
xnor U6986 (N_6986,N_179,N_4599);
and U6987 (N_6987,N_1868,N_4921);
and U6988 (N_6988,N_4614,N_1569);
nor U6989 (N_6989,N_3293,N_943);
nand U6990 (N_6990,N_4829,N_1636);
xnor U6991 (N_6991,N_4679,N_818);
or U6992 (N_6992,N_1954,N_3287);
xor U6993 (N_6993,N_363,N_1519);
and U6994 (N_6994,N_3948,N_2225);
nand U6995 (N_6995,N_1701,N_1739);
and U6996 (N_6996,N_92,N_1300);
nor U6997 (N_6997,N_4897,N_4443);
or U6998 (N_6998,N_295,N_948);
nand U6999 (N_6999,N_2456,N_4469);
nand U7000 (N_7000,N_2425,N_2011);
nor U7001 (N_7001,N_3018,N_779);
nor U7002 (N_7002,N_3119,N_941);
or U7003 (N_7003,N_2074,N_3336);
xor U7004 (N_7004,N_3442,N_4479);
xnor U7005 (N_7005,N_737,N_1663);
or U7006 (N_7006,N_3292,N_4925);
nor U7007 (N_7007,N_1483,N_4379);
nor U7008 (N_7008,N_3867,N_1118);
nand U7009 (N_7009,N_801,N_3707);
or U7010 (N_7010,N_172,N_3043);
nand U7011 (N_7011,N_2962,N_2480);
nand U7012 (N_7012,N_2915,N_42);
or U7013 (N_7013,N_3169,N_2430);
and U7014 (N_7014,N_3731,N_1529);
xnor U7015 (N_7015,N_2559,N_489);
xor U7016 (N_7016,N_4341,N_4792);
nor U7017 (N_7017,N_4539,N_431);
nor U7018 (N_7018,N_3242,N_1478);
nor U7019 (N_7019,N_2350,N_852);
and U7020 (N_7020,N_3017,N_3190);
xnor U7021 (N_7021,N_1180,N_2979);
xnor U7022 (N_7022,N_1107,N_4864);
nor U7023 (N_7023,N_1464,N_2018);
nor U7024 (N_7024,N_1231,N_4200);
nand U7025 (N_7025,N_4127,N_1800);
nand U7026 (N_7026,N_3047,N_4934);
nand U7027 (N_7027,N_4760,N_1213);
nand U7028 (N_7028,N_1142,N_4237);
and U7029 (N_7029,N_3228,N_3723);
or U7030 (N_7030,N_61,N_1162);
and U7031 (N_7031,N_607,N_2554);
nor U7032 (N_7032,N_1135,N_1603);
nor U7033 (N_7033,N_2044,N_2753);
or U7034 (N_7034,N_4955,N_4274);
or U7035 (N_7035,N_2303,N_3985);
nand U7036 (N_7036,N_1562,N_4209);
nor U7037 (N_7037,N_3356,N_1921);
nand U7038 (N_7038,N_687,N_177);
nor U7039 (N_7039,N_2077,N_1456);
nand U7040 (N_7040,N_4943,N_3106);
xnor U7041 (N_7041,N_4807,N_3419);
nand U7042 (N_7042,N_4531,N_2001);
or U7043 (N_7043,N_3897,N_3083);
and U7044 (N_7044,N_4579,N_3957);
xnor U7045 (N_7045,N_1228,N_4843);
nand U7046 (N_7046,N_129,N_2967);
nand U7047 (N_7047,N_4374,N_4994);
xnor U7048 (N_7048,N_1521,N_359);
nor U7049 (N_7049,N_3708,N_67);
nor U7050 (N_7050,N_3780,N_744);
nand U7051 (N_7051,N_4344,N_3564);
and U7052 (N_7052,N_1711,N_1567);
xor U7053 (N_7053,N_1993,N_893);
or U7054 (N_7054,N_4573,N_2742);
nand U7055 (N_7055,N_4666,N_176);
and U7056 (N_7056,N_4985,N_50);
nor U7057 (N_7057,N_4702,N_536);
xnor U7058 (N_7058,N_1499,N_3738);
nand U7059 (N_7059,N_1808,N_2313);
nand U7060 (N_7060,N_76,N_2916);
nand U7061 (N_7061,N_548,N_2078);
and U7062 (N_7062,N_794,N_2536);
xnor U7063 (N_7063,N_4482,N_2324);
xnor U7064 (N_7064,N_4296,N_2607);
or U7065 (N_7065,N_2203,N_4096);
and U7066 (N_7066,N_1812,N_1545);
or U7067 (N_7067,N_3746,N_3360);
nor U7068 (N_7068,N_3619,N_276);
nand U7069 (N_7069,N_4332,N_113);
nor U7070 (N_7070,N_2310,N_4528);
and U7071 (N_7071,N_1366,N_3177);
nand U7072 (N_7072,N_1850,N_2668);
and U7073 (N_7073,N_2171,N_1344);
or U7074 (N_7074,N_4907,N_2550);
nor U7075 (N_7075,N_2012,N_905);
nor U7076 (N_7076,N_1617,N_4207);
xnor U7077 (N_7077,N_3213,N_4418);
nor U7078 (N_7078,N_2807,N_754);
and U7079 (N_7079,N_2558,N_1925);
nand U7080 (N_7080,N_4119,N_2521);
or U7081 (N_7081,N_2615,N_2883);
nand U7082 (N_7082,N_507,N_3331);
xnor U7083 (N_7083,N_2990,N_4742);
or U7084 (N_7084,N_3110,N_4194);
and U7085 (N_7085,N_2093,N_4828);
xor U7086 (N_7086,N_2416,N_986);
nor U7087 (N_7087,N_3642,N_211);
nand U7088 (N_7088,N_3637,N_1968);
nor U7089 (N_7089,N_825,N_4261);
or U7090 (N_7090,N_4185,N_2598);
nor U7091 (N_7091,N_787,N_4335);
nor U7092 (N_7092,N_4030,N_4536);
or U7093 (N_7093,N_4862,N_3353);
and U7094 (N_7094,N_994,N_1957);
and U7095 (N_7095,N_1184,N_3125);
nand U7096 (N_7096,N_4672,N_413);
nand U7097 (N_7097,N_2889,N_2423);
or U7098 (N_7098,N_4007,N_1702);
or U7099 (N_7099,N_4390,N_3796);
nand U7100 (N_7100,N_521,N_4142);
nor U7101 (N_7101,N_1035,N_1848);
or U7102 (N_7102,N_1922,N_4080);
xor U7103 (N_7103,N_4134,N_4636);
nor U7104 (N_7104,N_4544,N_3329);
nor U7105 (N_7105,N_4219,N_3133);
nor U7106 (N_7106,N_3306,N_1891);
xor U7107 (N_7107,N_3217,N_2209);
and U7108 (N_7108,N_3257,N_4110);
xor U7109 (N_7109,N_1251,N_2133);
nor U7110 (N_7110,N_4148,N_4653);
nor U7111 (N_7111,N_3102,N_3691);
nor U7112 (N_7112,N_1326,N_29);
nand U7113 (N_7113,N_4022,N_3680);
xor U7114 (N_7114,N_1775,N_2387);
or U7115 (N_7115,N_592,N_2027);
and U7116 (N_7116,N_2576,N_1750);
nand U7117 (N_7117,N_3961,N_74);
or U7118 (N_7118,N_4773,N_1970);
nand U7119 (N_7119,N_836,N_4892);
xnor U7120 (N_7120,N_2499,N_4598);
or U7121 (N_7121,N_843,N_4629);
nand U7122 (N_7122,N_1336,N_1515);
and U7123 (N_7123,N_4391,N_3808);
or U7124 (N_7124,N_3201,N_323);
nor U7125 (N_7125,N_4952,N_3990);
or U7126 (N_7126,N_3462,N_3861);
or U7127 (N_7127,N_2851,N_1235);
and U7128 (N_7128,N_1833,N_2957);
nand U7129 (N_7129,N_3270,N_4777);
nor U7130 (N_7130,N_1308,N_1129);
or U7131 (N_7131,N_3432,N_3127);
nor U7132 (N_7132,N_1474,N_3004);
nor U7133 (N_7133,N_2589,N_2831);
xor U7134 (N_7134,N_2034,N_3424);
xor U7135 (N_7135,N_3143,N_2016);
nand U7136 (N_7136,N_3954,N_3455);
nand U7137 (N_7137,N_743,N_2401);
or U7138 (N_7138,N_382,N_1612);
and U7139 (N_7139,N_1475,N_1517);
xor U7140 (N_7140,N_2347,N_1793);
xor U7141 (N_7141,N_2959,N_674);
or U7142 (N_7142,N_4483,N_740);
or U7143 (N_7143,N_4947,N_2138);
nor U7144 (N_7144,N_1004,N_1342);
nor U7145 (N_7145,N_1997,N_3551);
nand U7146 (N_7146,N_3831,N_1255);
nand U7147 (N_7147,N_1121,N_1412);
nand U7148 (N_7148,N_2813,N_3286);
nor U7149 (N_7149,N_4214,N_640);
nand U7150 (N_7150,N_4566,N_1864);
nand U7151 (N_7151,N_102,N_1126);
nand U7152 (N_7152,N_996,N_733);
nand U7153 (N_7153,N_543,N_952);
xnor U7154 (N_7154,N_1254,N_2407);
or U7155 (N_7155,N_4560,N_2126);
nor U7156 (N_7156,N_13,N_4977);
nor U7157 (N_7157,N_4979,N_277);
and U7158 (N_7158,N_3915,N_672);
or U7159 (N_7159,N_4810,N_3091);
and U7160 (N_7160,N_2398,N_3895);
or U7161 (N_7161,N_2131,N_4825);
nor U7162 (N_7162,N_3859,N_984);
nor U7163 (N_7163,N_724,N_1417);
xnor U7164 (N_7164,N_667,N_2402);
nand U7165 (N_7165,N_2621,N_2839);
and U7166 (N_7166,N_3906,N_2193);
nand U7167 (N_7167,N_2994,N_3206);
or U7168 (N_7168,N_3899,N_3875);
and U7169 (N_7169,N_1672,N_1589);
nand U7170 (N_7170,N_2564,N_1225);
xnor U7171 (N_7171,N_2266,N_3176);
nand U7172 (N_7172,N_485,N_3325);
xor U7173 (N_7173,N_1682,N_1605);
nand U7174 (N_7174,N_3542,N_4177);
nor U7175 (N_7175,N_4978,N_3403);
nor U7176 (N_7176,N_788,N_1007);
or U7177 (N_7177,N_26,N_2583);
nor U7178 (N_7178,N_1406,N_1949);
xnor U7179 (N_7179,N_1445,N_252);
xor U7180 (N_7180,N_4439,N_1400);
nor U7181 (N_7181,N_4198,N_2002);
nor U7182 (N_7182,N_2765,N_4912);
xor U7183 (N_7183,N_522,N_2339);
or U7184 (N_7184,N_2605,N_268);
or U7185 (N_7185,N_533,N_4838);
xor U7186 (N_7186,N_4234,N_2667);
and U7187 (N_7187,N_4534,N_2798);
and U7188 (N_7188,N_1600,N_2846);
nand U7189 (N_7189,N_3940,N_3801);
and U7190 (N_7190,N_43,N_2606);
nor U7191 (N_7191,N_4815,N_1753);
or U7192 (N_7192,N_3319,N_1555);
nand U7193 (N_7193,N_881,N_1176);
or U7194 (N_7194,N_4607,N_669);
or U7195 (N_7195,N_3031,N_112);
nor U7196 (N_7196,N_896,N_1114);
and U7197 (N_7197,N_866,N_3362);
and U7198 (N_7198,N_4506,N_443);
nor U7199 (N_7199,N_3049,N_1261);
xor U7200 (N_7200,N_1230,N_1419);
or U7201 (N_7201,N_77,N_3803);
or U7202 (N_7202,N_178,N_3086);
nand U7203 (N_7203,N_1248,N_1976);
xnor U7204 (N_7204,N_745,N_1303);
xnor U7205 (N_7205,N_4001,N_317);
nand U7206 (N_7206,N_1398,N_4493);
or U7207 (N_7207,N_4511,N_4529);
nor U7208 (N_7208,N_1675,N_1333);
nor U7209 (N_7209,N_391,N_1566);
and U7210 (N_7210,N_2365,N_3369);
nor U7211 (N_7211,N_3800,N_1924);
and U7212 (N_7212,N_3416,N_3616);
xor U7213 (N_7213,N_2534,N_1528);
nor U7214 (N_7214,N_2276,N_2482);
or U7215 (N_7215,N_714,N_3583);
and U7216 (N_7216,N_2345,N_4969);
xor U7217 (N_7217,N_3883,N_3541);
or U7218 (N_7218,N_4436,N_130);
or U7219 (N_7219,N_686,N_835);
nand U7220 (N_7220,N_1164,N_3890);
or U7221 (N_7221,N_1609,N_3987);
nand U7222 (N_7222,N_349,N_3263);
or U7223 (N_7223,N_2248,N_1195);
and U7224 (N_7224,N_410,N_2555);
nand U7225 (N_7225,N_2827,N_141);
xnor U7226 (N_7226,N_2833,N_348);
nand U7227 (N_7227,N_3905,N_19);
and U7228 (N_7228,N_362,N_2644);
or U7229 (N_7229,N_1069,N_4396);
xnor U7230 (N_7230,N_4663,N_3936);
xor U7231 (N_7231,N_3949,N_2084);
xor U7232 (N_7232,N_1153,N_3809);
nand U7233 (N_7233,N_828,N_3752);
or U7234 (N_7234,N_3713,N_2337);
nor U7235 (N_7235,N_3208,N_1482);
or U7236 (N_7236,N_396,N_3390);
nand U7237 (N_7237,N_2160,N_3024);
or U7238 (N_7238,N_90,N_2222);
nor U7239 (N_7239,N_1996,N_3056);
and U7240 (N_7240,N_1339,N_2910);
or U7241 (N_7241,N_3132,N_3052);
nand U7242 (N_7242,N_1022,N_1717);
nand U7243 (N_7243,N_1314,N_1917);
xor U7244 (N_7244,N_23,N_4699);
xor U7245 (N_7245,N_3351,N_3338);
xnor U7246 (N_7246,N_2912,N_3576);
and U7247 (N_7247,N_4658,N_2549);
or U7248 (N_7248,N_3727,N_2789);
nand U7249 (N_7249,N_1749,N_3367);
nand U7250 (N_7250,N_576,N_861);
nor U7251 (N_7251,N_1712,N_872);
and U7252 (N_7252,N_953,N_2594);
or U7253 (N_7253,N_748,N_2590);
nor U7254 (N_7254,N_3400,N_82);
xnor U7255 (N_7255,N_3783,N_3477);
or U7256 (N_7256,N_2341,N_3033);
nor U7257 (N_7257,N_1502,N_1897);
nor U7258 (N_7258,N_2637,N_2999);
xnor U7259 (N_7259,N_1988,N_2397);
and U7260 (N_7260,N_4716,N_1272);
nor U7261 (N_7261,N_4933,N_4852);
or U7262 (N_7262,N_4035,N_4569);
xnor U7263 (N_7263,N_1874,N_3317);
or U7264 (N_7264,N_2369,N_4659);
nand U7265 (N_7265,N_239,N_273);
xnor U7266 (N_7266,N_1725,N_1356);
or U7267 (N_7267,N_3383,N_1503);
nor U7268 (N_7268,N_1206,N_56);
and U7269 (N_7269,N_3352,N_2727);
or U7270 (N_7270,N_4095,N_2938);
and U7271 (N_7271,N_1858,N_4478);
nor U7272 (N_7272,N_1872,N_401);
or U7273 (N_7273,N_3536,N_4459);
xnor U7274 (N_7274,N_2342,N_4224);
nand U7275 (N_7275,N_4348,N_314);
xor U7276 (N_7276,N_491,N_2484);
xor U7277 (N_7277,N_1776,N_3300);
nor U7278 (N_7278,N_3473,N_1774);
nand U7279 (N_7279,N_727,N_2185);
and U7280 (N_7280,N_3009,N_1834);
or U7281 (N_7281,N_4836,N_692);
xor U7282 (N_7282,N_2240,N_4762);
nor U7283 (N_7283,N_654,N_3092);
nand U7284 (N_7284,N_2004,N_4771);
or U7285 (N_7285,N_3998,N_1387);
and U7286 (N_7286,N_291,N_3280);
nor U7287 (N_7287,N_3692,N_3684);
nor U7288 (N_7288,N_4254,N_3281);
or U7289 (N_7289,N_3553,N_1396);
and U7290 (N_7290,N_3002,N_4597);
or U7291 (N_7291,N_2578,N_194);
nor U7292 (N_7292,N_2713,N_1278);
or U7293 (N_7293,N_4787,N_4756);
nand U7294 (N_7294,N_978,N_4740);
or U7295 (N_7295,N_4586,N_3749);
nand U7296 (N_7296,N_4019,N_2167);
nand U7297 (N_7297,N_4625,N_4378);
and U7298 (N_7298,N_4226,N_318);
and U7299 (N_7299,N_426,N_404);
xor U7300 (N_7300,N_1492,N_4790);
xnor U7301 (N_7301,N_992,N_1331);
nor U7302 (N_7302,N_3162,N_334);
nand U7303 (N_7303,N_3816,N_2444);
or U7304 (N_7304,N_4476,N_4924);
and U7305 (N_7305,N_1249,N_1525);
xor U7306 (N_7306,N_1053,N_3888);
nor U7307 (N_7307,N_3914,N_1096);
nand U7308 (N_7308,N_1571,N_2058);
xor U7309 (N_7309,N_2577,N_4117);
nor U7310 (N_7310,N_3508,N_4667);
or U7311 (N_7311,N_4874,N_3511);
xnor U7312 (N_7312,N_3202,N_4413);
xnor U7313 (N_7313,N_2293,N_332);
or U7314 (N_7314,N_3568,N_2890);
or U7315 (N_7315,N_3412,N_1821);
xnor U7316 (N_7316,N_4315,N_375);
xnor U7317 (N_7317,N_3601,N_842);
and U7318 (N_7318,N_910,N_1305);
and U7319 (N_7319,N_1524,N_900);
nand U7320 (N_7320,N_3753,N_4875);
xor U7321 (N_7321,N_2744,N_3323);
or U7322 (N_7322,N_4923,N_365);
xnor U7323 (N_7323,N_4190,N_3122);
or U7324 (N_7324,N_3943,N_4271);
nor U7325 (N_7325,N_40,N_2317);
and U7326 (N_7326,N_4863,N_3893);
xnor U7327 (N_7327,N_4368,N_4564);
and U7328 (N_7328,N_3030,N_2438);
and U7329 (N_7329,N_2280,N_1641);
xnor U7330 (N_7330,N_2100,N_2472);
xor U7331 (N_7331,N_922,N_1940);
nor U7332 (N_7332,N_2198,N_1530);
xnor U7333 (N_7333,N_1615,N_4680);
nor U7334 (N_7334,N_2710,N_3555);
and U7335 (N_7335,N_3435,N_1853);
nor U7336 (N_7336,N_4129,N_742);
nand U7337 (N_7337,N_4229,N_2254);
nand U7338 (N_7338,N_3834,N_2106);
xor U7339 (N_7339,N_2855,N_645);
xnor U7340 (N_7340,N_945,N_2255);
or U7341 (N_7341,N_3487,N_2746);
and U7342 (N_7342,N_3085,N_646);
nand U7343 (N_7343,N_2773,N_1563);
nor U7344 (N_7344,N_3670,N_101);
or U7345 (N_7345,N_3744,N_2842);
or U7346 (N_7346,N_2461,N_4429);
nor U7347 (N_7347,N_1744,N_1758);
nand U7348 (N_7348,N_2390,N_1520);
nand U7349 (N_7349,N_1165,N_3309);
or U7350 (N_7350,N_169,N_2204);
xnor U7351 (N_7351,N_4297,N_1735);
xnor U7352 (N_7352,N_3735,N_258);
xnor U7353 (N_7353,N_4993,N_1959);
and U7354 (N_7354,N_1580,N_3937);
nor U7355 (N_7355,N_707,N_2950);
nor U7356 (N_7356,N_2539,N_3196);
nor U7357 (N_7357,N_63,N_4989);
nor U7358 (N_7358,N_4041,N_1944);
or U7359 (N_7359,N_2629,N_4619);
and U7360 (N_7360,N_2188,N_230);
and U7361 (N_7361,N_117,N_3614);
or U7362 (N_7362,N_1601,N_4010);
or U7363 (N_7363,N_1938,N_889);
and U7364 (N_7364,N_1072,N_3647);
nand U7365 (N_7365,N_2340,N_1498);
nand U7366 (N_7366,N_1631,N_4245);
nand U7367 (N_7367,N_997,N_1446);
nor U7368 (N_7368,N_3545,N_2315);
xnor U7369 (N_7369,N_4146,N_1551);
nand U7370 (N_7370,N_4472,N_749);
nand U7371 (N_7371,N_720,N_1966);
and U7372 (N_7372,N_898,N_4966);
and U7373 (N_7373,N_3569,N_4057);
and U7374 (N_7374,N_864,N_3627);
nor U7375 (N_7375,N_4973,N_2553);
xor U7376 (N_7376,N_1779,N_2879);
xor U7377 (N_7377,N_214,N_190);
xnor U7378 (N_7378,N_3795,N_2275);
xor U7379 (N_7379,N_3355,N_3114);
and U7380 (N_7380,N_933,N_2238);
xor U7381 (N_7381,N_4444,N_609);
and U7382 (N_7382,N_1813,N_3894);
xor U7383 (N_7383,N_1147,N_747);
or U7384 (N_7384,N_3469,N_2677);
or U7385 (N_7385,N_2768,N_3747);
xor U7386 (N_7386,N_219,N_951);
nor U7387 (N_7387,N_1316,N_2071);
nor U7388 (N_7388,N_2119,N_4974);
nor U7389 (N_7389,N_3685,N_2760);
nor U7390 (N_7390,N_2551,N_1094);
nand U7391 (N_7391,N_1728,N_3365);
or U7392 (N_7392,N_4768,N_111);
xnor U7393 (N_7393,N_3251,N_2041);
nor U7394 (N_7394,N_3129,N_153);
or U7395 (N_7395,N_3930,N_3465);
or U7396 (N_7396,N_4783,N_54);
xor U7397 (N_7397,N_2122,N_3063);
nand U7398 (N_7398,N_4356,N_344);
nor U7399 (N_7399,N_4400,N_1246);
and U7400 (N_7400,N_15,N_3538);
or U7401 (N_7401,N_107,N_1177);
xnor U7402 (N_7402,N_3879,N_1500);
nand U7403 (N_7403,N_3246,N_3451);
and U7404 (N_7404,N_4343,N_1918);
or U7405 (N_7405,N_2940,N_3268);
and U7406 (N_7406,N_2619,N_4669);
and U7407 (N_7407,N_2066,N_4735);
or U7408 (N_7408,N_4003,N_231);
nand U7409 (N_7409,N_611,N_3821);
and U7410 (N_7410,N_3479,N_441);
and U7411 (N_7411,N_1836,N_1943);
nand U7412 (N_7412,N_2405,N_4811);
and U7413 (N_7413,N_1838,N_762);
or U7414 (N_7414,N_1644,N_4738);
and U7415 (N_7415,N_4775,N_2221);
nand U7416 (N_7416,N_134,N_3767);
or U7417 (N_7417,N_3172,N_4090);
nand U7418 (N_7418,N_1805,N_2601);
xnor U7419 (N_7419,N_3134,N_4909);
xnor U7420 (N_7420,N_2471,N_1347);
nor U7421 (N_7421,N_2961,N_1409);
nor U7422 (N_7422,N_3483,N_269);
nor U7423 (N_7423,N_103,N_4350);
and U7424 (N_7424,N_1103,N_3606);
nor U7425 (N_7425,N_2685,N_2419);
or U7426 (N_7426,N_3220,N_1514);
or U7427 (N_7427,N_4322,N_3799);
nor U7428 (N_7428,N_4205,N_2849);
nand U7429 (N_7429,N_2290,N_3668);
or U7430 (N_7430,N_2620,N_569);
xor U7431 (N_7431,N_1084,N_2309);
nor U7432 (N_7432,N_1418,N_3399);
nor U7433 (N_7433,N_1043,N_1081);
and U7434 (N_7434,N_478,N_2800);
and U7435 (N_7435,N_3407,N_875);
or U7436 (N_7436,N_3778,N_1914);
and U7437 (N_7437,N_4481,N_53);
or U7438 (N_7438,N_2194,N_3751);
xor U7439 (N_7439,N_2899,N_627);
or U7440 (N_7440,N_1161,N_3661);
or U7441 (N_7441,N_3069,N_2970);
or U7442 (N_7442,N_4169,N_1608);
nand U7443 (N_7443,N_4883,N_4954);
nand U7444 (N_7444,N_1209,N_845);
xnor U7445 (N_7445,N_2652,N_519);
nor U7446 (N_7446,N_1882,N_25);
nor U7447 (N_7447,N_3840,N_1260);
xor U7448 (N_7448,N_4367,N_3230);
xnor U7449 (N_7449,N_2338,N_3827);
or U7450 (N_7450,N_167,N_1273);
and U7451 (N_7451,N_3188,N_2056);
or U7452 (N_7452,N_3420,N_1947);
and U7453 (N_7453,N_1990,N_1570);
and U7454 (N_7454,N_4580,N_3411);
nand U7455 (N_7455,N_4346,N_2905);
nand U7456 (N_7456,N_2506,N_4861);
or U7457 (N_7457,N_4505,N_1397);
and U7458 (N_7458,N_4583,N_2974);
nand U7459 (N_7459,N_4557,N_1294);
and U7460 (N_7460,N_590,N_131);
and U7461 (N_7461,N_1027,N_4020);
xor U7462 (N_7462,N_3184,N_3918);
nor U7463 (N_7463,N_606,N_2166);
and U7464 (N_7464,N_2638,N_4111);
nor U7465 (N_7465,N_185,N_476);
or U7466 (N_7466,N_2156,N_2124);
nand U7467 (N_7467,N_2112,N_2701);
or U7468 (N_7468,N_2178,N_4065);
nor U7469 (N_7469,N_3255,N_3392);
xnor U7470 (N_7470,N_374,N_1553);
xor U7471 (N_7471,N_3042,N_3197);
and U7472 (N_7472,N_2076,N_1334);
nor U7473 (N_7473,N_3008,N_1237);
xor U7474 (N_7474,N_2686,N_400);
xnor U7475 (N_7475,N_2891,N_4616);
xor U7476 (N_7476,N_1017,N_3151);
xnor U7477 (N_7477,N_3067,N_4645);
xnor U7478 (N_7478,N_2529,N_4492);
and U7479 (N_7479,N_4971,N_4990);
and U7480 (N_7480,N_1723,N_1279);
xnor U7481 (N_7481,N_379,N_1430);
xnor U7482 (N_7482,N_3327,N_2739);
xor U7483 (N_7483,N_1016,N_4719);
xnor U7484 (N_7484,N_154,N_234);
xor U7485 (N_7485,N_1554,N_4704);
xnor U7486 (N_7486,N_2604,N_1830);
nor U7487 (N_7487,N_4542,N_776);
nor U7488 (N_7488,N_2202,N_1832);
and U7489 (N_7489,N_2740,N_301);
nor U7490 (N_7490,N_912,N_4565);
and U7491 (N_7491,N_4456,N_3605);
nor U7492 (N_7492,N_790,N_4867);
nand U7493 (N_7493,N_3115,N_1653);
or U7494 (N_7494,N_4673,N_916);
and U7495 (N_7495,N_2274,N_799);
nand U7496 (N_7496,N_3440,N_664);
or U7497 (N_7497,N_1778,N_4358);
xor U7498 (N_7498,N_3665,N_2692);
nor U7499 (N_7499,N_2007,N_663);
nand U7500 (N_7500,N_2345,N_4878);
or U7501 (N_7501,N_3115,N_3043);
and U7502 (N_7502,N_2427,N_4660);
nor U7503 (N_7503,N_2265,N_4421);
xnor U7504 (N_7504,N_1351,N_393);
xnor U7505 (N_7505,N_3007,N_2781);
xor U7506 (N_7506,N_1821,N_3603);
xor U7507 (N_7507,N_4998,N_2852);
or U7508 (N_7508,N_3743,N_1696);
nand U7509 (N_7509,N_2092,N_2930);
xor U7510 (N_7510,N_1440,N_48);
or U7511 (N_7511,N_2597,N_2351);
xor U7512 (N_7512,N_2809,N_357);
nand U7513 (N_7513,N_4954,N_4248);
nand U7514 (N_7514,N_2562,N_413);
xnor U7515 (N_7515,N_2270,N_1733);
or U7516 (N_7516,N_2167,N_2329);
xnor U7517 (N_7517,N_1663,N_4314);
xnor U7518 (N_7518,N_593,N_613);
nor U7519 (N_7519,N_2074,N_2947);
xnor U7520 (N_7520,N_320,N_991);
xnor U7521 (N_7521,N_3913,N_3433);
nand U7522 (N_7522,N_4012,N_750);
nor U7523 (N_7523,N_3271,N_2147);
nand U7524 (N_7524,N_3006,N_2214);
and U7525 (N_7525,N_2479,N_3807);
nand U7526 (N_7526,N_463,N_1455);
nand U7527 (N_7527,N_2102,N_859);
and U7528 (N_7528,N_1479,N_4538);
and U7529 (N_7529,N_3687,N_4362);
or U7530 (N_7530,N_2688,N_2695);
or U7531 (N_7531,N_1068,N_3548);
xor U7532 (N_7532,N_2942,N_887);
xnor U7533 (N_7533,N_4437,N_1189);
nand U7534 (N_7534,N_1626,N_4471);
xor U7535 (N_7535,N_4228,N_3959);
or U7536 (N_7536,N_1871,N_513);
and U7537 (N_7537,N_4530,N_41);
and U7538 (N_7538,N_2202,N_1888);
or U7539 (N_7539,N_4789,N_487);
xor U7540 (N_7540,N_2044,N_2019);
xor U7541 (N_7541,N_2022,N_2148);
and U7542 (N_7542,N_2908,N_400);
and U7543 (N_7543,N_1404,N_4464);
nor U7544 (N_7544,N_3927,N_2845);
and U7545 (N_7545,N_1727,N_797);
nor U7546 (N_7546,N_2637,N_4088);
nor U7547 (N_7547,N_281,N_3550);
nand U7548 (N_7548,N_2557,N_849);
or U7549 (N_7549,N_4352,N_3831);
or U7550 (N_7550,N_1961,N_3963);
nand U7551 (N_7551,N_1231,N_2372);
nand U7552 (N_7552,N_3118,N_4973);
nand U7553 (N_7553,N_2583,N_2557);
or U7554 (N_7554,N_3980,N_102);
nand U7555 (N_7555,N_3663,N_3886);
and U7556 (N_7556,N_2922,N_1619);
or U7557 (N_7557,N_3834,N_1778);
xnor U7558 (N_7558,N_597,N_919);
and U7559 (N_7559,N_3744,N_4079);
nor U7560 (N_7560,N_147,N_3395);
nor U7561 (N_7561,N_1538,N_2526);
nand U7562 (N_7562,N_4320,N_191);
and U7563 (N_7563,N_4865,N_275);
xnor U7564 (N_7564,N_812,N_791);
nand U7565 (N_7565,N_1400,N_3069);
and U7566 (N_7566,N_1995,N_3212);
xor U7567 (N_7567,N_2025,N_2447);
nor U7568 (N_7568,N_2202,N_2042);
nand U7569 (N_7569,N_1980,N_3692);
nand U7570 (N_7570,N_2973,N_1313);
nand U7571 (N_7571,N_1947,N_1191);
and U7572 (N_7572,N_3684,N_3569);
and U7573 (N_7573,N_1833,N_4885);
and U7574 (N_7574,N_1410,N_4301);
nor U7575 (N_7575,N_341,N_1883);
and U7576 (N_7576,N_556,N_1280);
nor U7577 (N_7577,N_1024,N_3998);
or U7578 (N_7578,N_3752,N_3319);
xnor U7579 (N_7579,N_4244,N_3564);
xor U7580 (N_7580,N_796,N_1169);
or U7581 (N_7581,N_4670,N_1033);
nor U7582 (N_7582,N_46,N_3746);
nand U7583 (N_7583,N_3639,N_2181);
xnor U7584 (N_7584,N_3321,N_4930);
xor U7585 (N_7585,N_1668,N_3772);
nand U7586 (N_7586,N_4725,N_2713);
nand U7587 (N_7587,N_2946,N_394);
nor U7588 (N_7588,N_2078,N_4408);
nor U7589 (N_7589,N_775,N_4980);
xnor U7590 (N_7590,N_981,N_1914);
nand U7591 (N_7591,N_4410,N_108);
nand U7592 (N_7592,N_967,N_1171);
nand U7593 (N_7593,N_2298,N_834);
nor U7594 (N_7594,N_3528,N_4712);
or U7595 (N_7595,N_3484,N_1942);
xor U7596 (N_7596,N_2765,N_2324);
xnor U7597 (N_7597,N_1570,N_2111);
nand U7598 (N_7598,N_1645,N_942);
xor U7599 (N_7599,N_3429,N_797);
or U7600 (N_7600,N_1184,N_4710);
nand U7601 (N_7601,N_2672,N_1388);
xnor U7602 (N_7602,N_4090,N_2496);
or U7603 (N_7603,N_4325,N_576);
and U7604 (N_7604,N_4883,N_1010);
and U7605 (N_7605,N_3059,N_4569);
nor U7606 (N_7606,N_1370,N_1534);
xnor U7607 (N_7607,N_4019,N_311);
and U7608 (N_7608,N_1779,N_557);
and U7609 (N_7609,N_228,N_3562);
or U7610 (N_7610,N_1827,N_1224);
nor U7611 (N_7611,N_4677,N_4059);
and U7612 (N_7612,N_819,N_4837);
or U7613 (N_7613,N_3515,N_797);
or U7614 (N_7614,N_1902,N_2720);
nand U7615 (N_7615,N_169,N_2206);
and U7616 (N_7616,N_4095,N_4411);
nor U7617 (N_7617,N_4083,N_615);
nand U7618 (N_7618,N_1230,N_3217);
nor U7619 (N_7619,N_4465,N_3956);
nor U7620 (N_7620,N_3282,N_3069);
nor U7621 (N_7621,N_2562,N_3352);
or U7622 (N_7622,N_432,N_1775);
xnor U7623 (N_7623,N_3365,N_3912);
xnor U7624 (N_7624,N_2081,N_2144);
xor U7625 (N_7625,N_1909,N_707);
xnor U7626 (N_7626,N_4335,N_4907);
or U7627 (N_7627,N_4419,N_1019);
xnor U7628 (N_7628,N_1019,N_2632);
or U7629 (N_7629,N_3309,N_3434);
nor U7630 (N_7630,N_3964,N_4977);
nand U7631 (N_7631,N_2243,N_1322);
nand U7632 (N_7632,N_2652,N_3967);
or U7633 (N_7633,N_90,N_1805);
nand U7634 (N_7634,N_3301,N_3555);
xor U7635 (N_7635,N_3051,N_2950);
nand U7636 (N_7636,N_48,N_4592);
and U7637 (N_7637,N_1981,N_3417);
and U7638 (N_7638,N_3728,N_3256);
xnor U7639 (N_7639,N_1621,N_4369);
and U7640 (N_7640,N_4459,N_573);
nand U7641 (N_7641,N_2523,N_3081);
nor U7642 (N_7642,N_4715,N_1643);
nand U7643 (N_7643,N_4595,N_180);
nand U7644 (N_7644,N_4920,N_2011);
xnor U7645 (N_7645,N_4197,N_3329);
or U7646 (N_7646,N_1748,N_3790);
xnor U7647 (N_7647,N_4092,N_2435);
nor U7648 (N_7648,N_482,N_3603);
xnor U7649 (N_7649,N_2602,N_1060);
or U7650 (N_7650,N_1616,N_4610);
nand U7651 (N_7651,N_4797,N_3705);
xnor U7652 (N_7652,N_1852,N_3203);
nand U7653 (N_7653,N_3904,N_605);
or U7654 (N_7654,N_3543,N_921);
nand U7655 (N_7655,N_4260,N_4592);
or U7656 (N_7656,N_4984,N_288);
nand U7657 (N_7657,N_4014,N_3177);
nand U7658 (N_7658,N_2739,N_4876);
nor U7659 (N_7659,N_1281,N_4128);
xnor U7660 (N_7660,N_3156,N_3521);
nand U7661 (N_7661,N_1609,N_4698);
nor U7662 (N_7662,N_2647,N_187);
and U7663 (N_7663,N_4483,N_2994);
xor U7664 (N_7664,N_1045,N_354);
xor U7665 (N_7665,N_1373,N_4721);
nand U7666 (N_7666,N_3907,N_3559);
nor U7667 (N_7667,N_2249,N_4661);
nor U7668 (N_7668,N_1909,N_3237);
xnor U7669 (N_7669,N_2994,N_4803);
and U7670 (N_7670,N_2231,N_1503);
and U7671 (N_7671,N_2859,N_4164);
xnor U7672 (N_7672,N_4775,N_1847);
and U7673 (N_7673,N_540,N_3187);
xor U7674 (N_7674,N_2099,N_2244);
nand U7675 (N_7675,N_4698,N_1042);
nor U7676 (N_7676,N_3515,N_906);
xnor U7677 (N_7677,N_2125,N_4372);
nor U7678 (N_7678,N_3900,N_1366);
nand U7679 (N_7679,N_1207,N_3164);
xor U7680 (N_7680,N_310,N_3676);
nor U7681 (N_7681,N_3552,N_426);
nor U7682 (N_7682,N_1347,N_4588);
or U7683 (N_7683,N_917,N_3505);
nor U7684 (N_7684,N_272,N_3834);
or U7685 (N_7685,N_165,N_4734);
nor U7686 (N_7686,N_4083,N_2758);
nand U7687 (N_7687,N_2015,N_4025);
nand U7688 (N_7688,N_2130,N_2277);
nor U7689 (N_7689,N_189,N_3290);
or U7690 (N_7690,N_1565,N_2204);
xnor U7691 (N_7691,N_1390,N_1267);
nand U7692 (N_7692,N_1147,N_4638);
nand U7693 (N_7693,N_3129,N_3538);
xnor U7694 (N_7694,N_3266,N_2053);
xnor U7695 (N_7695,N_66,N_4822);
or U7696 (N_7696,N_4139,N_1108);
nor U7697 (N_7697,N_4504,N_3732);
xnor U7698 (N_7698,N_648,N_3764);
or U7699 (N_7699,N_3603,N_1329);
or U7700 (N_7700,N_4751,N_3737);
xor U7701 (N_7701,N_1258,N_1741);
xnor U7702 (N_7702,N_397,N_1007);
nand U7703 (N_7703,N_2444,N_1825);
xnor U7704 (N_7704,N_3083,N_2630);
or U7705 (N_7705,N_1062,N_452);
nand U7706 (N_7706,N_4906,N_3933);
and U7707 (N_7707,N_4919,N_2864);
nor U7708 (N_7708,N_3985,N_1623);
or U7709 (N_7709,N_2779,N_3047);
nor U7710 (N_7710,N_63,N_3581);
nand U7711 (N_7711,N_1960,N_583);
nor U7712 (N_7712,N_2005,N_589);
or U7713 (N_7713,N_2151,N_3705);
or U7714 (N_7714,N_1559,N_1613);
nand U7715 (N_7715,N_2056,N_4128);
nor U7716 (N_7716,N_2682,N_3928);
or U7717 (N_7717,N_3840,N_3855);
xor U7718 (N_7718,N_4925,N_3401);
xor U7719 (N_7719,N_2719,N_1153);
and U7720 (N_7720,N_3236,N_4290);
nor U7721 (N_7721,N_3248,N_3941);
and U7722 (N_7722,N_4045,N_2558);
nor U7723 (N_7723,N_337,N_4541);
nor U7724 (N_7724,N_4124,N_3299);
nand U7725 (N_7725,N_2468,N_905);
nor U7726 (N_7726,N_2458,N_1959);
and U7727 (N_7727,N_1349,N_3328);
or U7728 (N_7728,N_4063,N_2066);
or U7729 (N_7729,N_77,N_2181);
or U7730 (N_7730,N_318,N_987);
or U7731 (N_7731,N_3414,N_2527);
xor U7732 (N_7732,N_4437,N_2946);
and U7733 (N_7733,N_3413,N_2571);
and U7734 (N_7734,N_2319,N_3027);
and U7735 (N_7735,N_578,N_2261);
xnor U7736 (N_7736,N_3017,N_4666);
xnor U7737 (N_7737,N_3518,N_4484);
nor U7738 (N_7738,N_3334,N_77);
xor U7739 (N_7739,N_1071,N_3119);
xnor U7740 (N_7740,N_4536,N_4311);
or U7741 (N_7741,N_763,N_3275);
or U7742 (N_7742,N_2393,N_2141);
nor U7743 (N_7743,N_2230,N_4948);
nand U7744 (N_7744,N_2486,N_4906);
xnor U7745 (N_7745,N_1049,N_2292);
nor U7746 (N_7746,N_4538,N_3204);
or U7747 (N_7747,N_4174,N_4745);
xor U7748 (N_7748,N_2137,N_4450);
and U7749 (N_7749,N_4432,N_4559);
or U7750 (N_7750,N_2619,N_3252);
nor U7751 (N_7751,N_4032,N_3140);
and U7752 (N_7752,N_1576,N_1739);
nor U7753 (N_7753,N_3586,N_2850);
xnor U7754 (N_7754,N_1539,N_1610);
and U7755 (N_7755,N_3853,N_2622);
and U7756 (N_7756,N_1528,N_4803);
nand U7757 (N_7757,N_4660,N_3291);
and U7758 (N_7758,N_4796,N_709);
and U7759 (N_7759,N_445,N_2268);
nor U7760 (N_7760,N_3399,N_977);
nand U7761 (N_7761,N_921,N_2455);
or U7762 (N_7762,N_3463,N_4585);
xor U7763 (N_7763,N_1246,N_3403);
nor U7764 (N_7764,N_3611,N_4139);
nand U7765 (N_7765,N_2861,N_3758);
nor U7766 (N_7766,N_1405,N_1939);
nand U7767 (N_7767,N_4857,N_4149);
and U7768 (N_7768,N_2530,N_3522);
and U7769 (N_7769,N_3176,N_906);
and U7770 (N_7770,N_4133,N_1800);
or U7771 (N_7771,N_4185,N_903);
nor U7772 (N_7772,N_1788,N_1573);
nor U7773 (N_7773,N_4029,N_1846);
nand U7774 (N_7774,N_582,N_3082);
xnor U7775 (N_7775,N_3064,N_2460);
or U7776 (N_7776,N_1700,N_2523);
nor U7777 (N_7777,N_203,N_1025);
and U7778 (N_7778,N_3292,N_3302);
nor U7779 (N_7779,N_739,N_3786);
nor U7780 (N_7780,N_1066,N_3039);
nand U7781 (N_7781,N_590,N_4107);
nand U7782 (N_7782,N_4921,N_1052);
nor U7783 (N_7783,N_1349,N_1982);
nand U7784 (N_7784,N_3433,N_4752);
nor U7785 (N_7785,N_2611,N_4788);
xor U7786 (N_7786,N_653,N_4652);
nand U7787 (N_7787,N_2289,N_1250);
and U7788 (N_7788,N_2371,N_3091);
xor U7789 (N_7789,N_2122,N_3795);
nand U7790 (N_7790,N_3689,N_389);
xor U7791 (N_7791,N_957,N_775);
nor U7792 (N_7792,N_1093,N_2989);
nor U7793 (N_7793,N_2204,N_2405);
nor U7794 (N_7794,N_4760,N_1436);
nor U7795 (N_7795,N_3147,N_629);
nand U7796 (N_7796,N_1456,N_3488);
xnor U7797 (N_7797,N_1048,N_2966);
nand U7798 (N_7798,N_1458,N_1236);
nor U7799 (N_7799,N_1981,N_2260);
xor U7800 (N_7800,N_4257,N_4120);
xnor U7801 (N_7801,N_3655,N_2285);
and U7802 (N_7802,N_2225,N_1231);
or U7803 (N_7803,N_515,N_2569);
nor U7804 (N_7804,N_2015,N_4488);
nand U7805 (N_7805,N_3204,N_4766);
xor U7806 (N_7806,N_3666,N_3061);
and U7807 (N_7807,N_2274,N_4850);
or U7808 (N_7808,N_276,N_48);
or U7809 (N_7809,N_4638,N_4097);
and U7810 (N_7810,N_4311,N_4744);
nand U7811 (N_7811,N_2346,N_2614);
and U7812 (N_7812,N_3163,N_3723);
nor U7813 (N_7813,N_360,N_1951);
or U7814 (N_7814,N_4388,N_574);
xor U7815 (N_7815,N_4464,N_3106);
or U7816 (N_7816,N_3082,N_482);
and U7817 (N_7817,N_986,N_443);
and U7818 (N_7818,N_2181,N_3456);
or U7819 (N_7819,N_2916,N_4934);
and U7820 (N_7820,N_553,N_3236);
nand U7821 (N_7821,N_4185,N_137);
or U7822 (N_7822,N_4860,N_2009);
xor U7823 (N_7823,N_2178,N_4631);
or U7824 (N_7824,N_860,N_3481);
nand U7825 (N_7825,N_55,N_3734);
and U7826 (N_7826,N_2485,N_1504);
nor U7827 (N_7827,N_1097,N_3893);
and U7828 (N_7828,N_2293,N_1234);
or U7829 (N_7829,N_4360,N_467);
nor U7830 (N_7830,N_4364,N_3826);
nand U7831 (N_7831,N_165,N_2685);
or U7832 (N_7832,N_2073,N_3084);
and U7833 (N_7833,N_2654,N_565);
xnor U7834 (N_7834,N_1648,N_1787);
or U7835 (N_7835,N_1328,N_4086);
nand U7836 (N_7836,N_1548,N_2908);
or U7837 (N_7837,N_1286,N_3464);
nand U7838 (N_7838,N_3803,N_2901);
and U7839 (N_7839,N_2372,N_4286);
xnor U7840 (N_7840,N_499,N_1548);
and U7841 (N_7841,N_1680,N_3459);
nor U7842 (N_7842,N_473,N_3891);
xnor U7843 (N_7843,N_1861,N_4132);
nand U7844 (N_7844,N_2638,N_466);
xor U7845 (N_7845,N_4434,N_3652);
xnor U7846 (N_7846,N_1825,N_588);
xnor U7847 (N_7847,N_3100,N_2754);
nand U7848 (N_7848,N_4562,N_1844);
nand U7849 (N_7849,N_3769,N_3444);
or U7850 (N_7850,N_3483,N_1934);
xnor U7851 (N_7851,N_1166,N_1223);
nand U7852 (N_7852,N_3069,N_3664);
or U7853 (N_7853,N_3770,N_2926);
and U7854 (N_7854,N_733,N_2917);
nand U7855 (N_7855,N_4619,N_2368);
nor U7856 (N_7856,N_3148,N_2397);
nor U7857 (N_7857,N_3622,N_2871);
and U7858 (N_7858,N_2383,N_995);
nand U7859 (N_7859,N_984,N_280);
xnor U7860 (N_7860,N_2818,N_1580);
xnor U7861 (N_7861,N_4890,N_2437);
nor U7862 (N_7862,N_4311,N_4285);
or U7863 (N_7863,N_3859,N_315);
nand U7864 (N_7864,N_1309,N_428);
or U7865 (N_7865,N_4818,N_1277);
and U7866 (N_7866,N_3592,N_4037);
and U7867 (N_7867,N_1552,N_4203);
nand U7868 (N_7868,N_402,N_2203);
xnor U7869 (N_7869,N_2405,N_4612);
nor U7870 (N_7870,N_1190,N_2829);
nor U7871 (N_7871,N_3700,N_1578);
xor U7872 (N_7872,N_4236,N_3939);
and U7873 (N_7873,N_1573,N_4901);
or U7874 (N_7874,N_1587,N_1193);
xnor U7875 (N_7875,N_2395,N_3987);
and U7876 (N_7876,N_860,N_2716);
xnor U7877 (N_7877,N_4414,N_3865);
and U7878 (N_7878,N_1351,N_1707);
and U7879 (N_7879,N_854,N_27);
or U7880 (N_7880,N_4469,N_3361);
nand U7881 (N_7881,N_1637,N_2451);
nand U7882 (N_7882,N_720,N_4682);
nand U7883 (N_7883,N_3305,N_4473);
nor U7884 (N_7884,N_3841,N_3739);
nor U7885 (N_7885,N_2,N_83);
xnor U7886 (N_7886,N_3378,N_4043);
nand U7887 (N_7887,N_883,N_4265);
nand U7888 (N_7888,N_1201,N_4423);
nand U7889 (N_7889,N_648,N_2375);
or U7890 (N_7890,N_1720,N_2404);
nor U7891 (N_7891,N_4248,N_72);
or U7892 (N_7892,N_969,N_3253);
xor U7893 (N_7893,N_1980,N_165);
xnor U7894 (N_7894,N_1950,N_2592);
or U7895 (N_7895,N_450,N_3882);
and U7896 (N_7896,N_1045,N_1926);
or U7897 (N_7897,N_2624,N_307);
nor U7898 (N_7898,N_1775,N_3558);
nor U7899 (N_7899,N_3984,N_1750);
xor U7900 (N_7900,N_3039,N_1599);
and U7901 (N_7901,N_318,N_2562);
or U7902 (N_7902,N_1276,N_1469);
or U7903 (N_7903,N_3378,N_499);
nor U7904 (N_7904,N_4340,N_4421);
nand U7905 (N_7905,N_4795,N_3122);
nand U7906 (N_7906,N_3558,N_2845);
nand U7907 (N_7907,N_957,N_3055);
or U7908 (N_7908,N_2578,N_3734);
nand U7909 (N_7909,N_2658,N_908);
nor U7910 (N_7910,N_3733,N_1488);
nor U7911 (N_7911,N_647,N_877);
nand U7912 (N_7912,N_4682,N_2211);
xor U7913 (N_7913,N_3846,N_4271);
nor U7914 (N_7914,N_1564,N_931);
nand U7915 (N_7915,N_1863,N_4367);
and U7916 (N_7916,N_96,N_956);
nand U7917 (N_7917,N_3802,N_2988);
nand U7918 (N_7918,N_1591,N_4560);
xnor U7919 (N_7919,N_4563,N_1657);
and U7920 (N_7920,N_1815,N_4675);
xnor U7921 (N_7921,N_3386,N_1685);
xor U7922 (N_7922,N_3832,N_3113);
nor U7923 (N_7923,N_4169,N_4175);
nor U7924 (N_7924,N_1488,N_4606);
and U7925 (N_7925,N_4808,N_4693);
nor U7926 (N_7926,N_3840,N_2358);
nand U7927 (N_7927,N_2344,N_1475);
nor U7928 (N_7928,N_3318,N_2588);
nand U7929 (N_7929,N_4225,N_2017);
xnor U7930 (N_7930,N_1337,N_1919);
and U7931 (N_7931,N_3184,N_2289);
nor U7932 (N_7932,N_4526,N_1368);
nand U7933 (N_7933,N_3602,N_1347);
nand U7934 (N_7934,N_768,N_232);
nand U7935 (N_7935,N_1130,N_255);
and U7936 (N_7936,N_628,N_2761);
xnor U7937 (N_7937,N_2697,N_1612);
xor U7938 (N_7938,N_645,N_1106);
and U7939 (N_7939,N_1392,N_1847);
or U7940 (N_7940,N_4286,N_1787);
and U7941 (N_7941,N_208,N_3998);
nand U7942 (N_7942,N_428,N_4133);
xnor U7943 (N_7943,N_3685,N_1349);
and U7944 (N_7944,N_2631,N_3951);
nor U7945 (N_7945,N_1147,N_3785);
and U7946 (N_7946,N_2038,N_3498);
nor U7947 (N_7947,N_1519,N_4423);
and U7948 (N_7948,N_56,N_1280);
or U7949 (N_7949,N_4889,N_2807);
nand U7950 (N_7950,N_3314,N_56);
nor U7951 (N_7951,N_2448,N_2478);
xor U7952 (N_7952,N_3349,N_1158);
nor U7953 (N_7953,N_4191,N_3128);
and U7954 (N_7954,N_2245,N_1674);
xnor U7955 (N_7955,N_3214,N_2946);
and U7956 (N_7956,N_914,N_537);
nor U7957 (N_7957,N_2862,N_1778);
or U7958 (N_7958,N_4225,N_1234);
xor U7959 (N_7959,N_3827,N_1095);
and U7960 (N_7960,N_367,N_2086);
nor U7961 (N_7961,N_4290,N_1771);
nand U7962 (N_7962,N_3560,N_4498);
or U7963 (N_7963,N_1698,N_3364);
and U7964 (N_7964,N_4517,N_343);
or U7965 (N_7965,N_2840,N_409);
nor U7966 (N_7966,N_4745,N_3305);
nor U7967 (N_7967,N_2688,N_2289);
and U7968 (N_7968,N_3639,N_803);
nand U7969 (N_7969,N_813,N_3202);
or U7970 (N_7970,N_4603,N_109);
nor U7971 (N_7971,N_325,N_785);
nor U7972 (N_7972,N_1195,N_4082);
or U7973 (N_7973,N_974,N_1503);
and U7974 (N_7974,N_1102,N_4382);
and U7975 (N_7975,N_4482,N_116);
xnor U7976 (N_7976,N_123,N_719);
nor U7977 (N_7977,N_3354,N_2863);
xnor U7978 (N_7978,N_156,N_2024);
or U7979 (N_7979,N_2454,N_1079);
and U7980 (N_7980,N_402,N_1543);
xnor U7981 (N_7981,N_1144,N_727);
or U7982 (N_7982,N_2093,N_797);
xor U7983 (N_7983,N_2785,N_4947);
and U7984 (N_7984,N_1655,N_1990);
and U7985 (N_7985,N_1064,N_1405);
or U7986 (N_7986,N_1579,N_1758);
or U7987 (N_7987,N_3335,N_2046);
or U7988 (N_7988,N_4159,N_1165);
xnor U7989 (N_7989,N_1348,N_155);
and U7990 (N_7990,N_3155,N_1195);
or U7991 (N_7991,N_4654,N_4185);
xor U7992 (N_7992,N_1199,N_1943);
and U7993 (N_7993,N_4469,N_4241);
and U7994 (N_7994,N_3362,N_4574);
nor U7995 (N_7995,N_4938,N_1602);
or U7996 (N_7996,N_1234,N_4720);
nor U7997 (N_7997,N_3637,N_3585);
nand U7998 (N_7998,N_1523,N_2667);
xnor U7999 (N_7999,N_1759,N_2227);
nor U8000 (N_8000,N_1181,N_1612);
nand U8001 (N_8001,N_3428,N_3457);
or U8002 (N_8002,N_1903,N_3619);
and U8003 (N_8003,N_2036,N_1801);
nor U8004 (N_8004,N_634,N_1376);
and U8005 (N_8005,N_416,N_2445);
and U8006 (N_8006,N_4564,N_3969);
and U8007 (N_8007,N_3342,N_1562);
or U8008 (N_8008,N_2797,N_4108);
xor U8009 (N_8009,N_3949,N_3795);
and U8010 (N_8010,N_2484,N_3940);
xnor U8011 (N_8011,N_1442,N_610);
xnor U8012 (N_8012,N_392,N_3976);
and U8013 (N_8013,N_4621,N_3893);
nor U8014 (N_8014,N_552,N_3934);
nor U8015 (N_8015,N_2241,N_1436);
nor U8016 (N_8016,N_61,N_1807);
nand U8017 (N_8017,N_1114,N_4800);
nor U8018 (N_8018,N_875,N_4841);
nor U8019 (N_8019,N_3662,N_3130);
nand U8020 (N_8020,N_1059,N_4091);
nand U8021 (N_8021,N_4032,N_1538);
and U8022 (N_8022,N_874,N_779);
nor U8023 (N_8023,N_305,N_1505);
nand U8024 (N_8024,N_1448,N_1136);
and U8025 (N_8025,N_2323,N_2470);
or U8026 (N_8026,N_4873,N_3902);
nand U8027 (N_8027,N_3605,N_1064);
or U8028 (N_8028,N_305,N_3224);
and U8029 (N_8029,N_4989,N_3408);
nor U8030 (N_8030,N_2292,N_236);
xnor U8031 (N_8031,N_2456,N_1049);
nor U8032 (N_8032,N_3946,N_616);
or U8033 (N_8033,N_307,N_2296);
nor U8034 (N_8034,N_2843,N_3664);
or U8035 (N_8035,N_630,N_4755);
and U8036 (N_8036,N_4689,N_193);
nand U8037 (N_8037,N_3376,N_2383);
nand U8038 (N_8038,N_4677,N_1050);
nand U8039 (N_8039,N_3349,N_4042);
xnor U8040 (N_8040,N_4996,N_703);
or U8041 (N_8041,N_2799,N_3692);
xor U8042 (N_8042,N_1691,N_3033);
or U8043 (N_8043,N_491,N_2241);
xnor U8044 (N_8044,N_1232,N_1840);
xnor U8045 (N_8045,N_4876,N_2696);
nand U8046 (N_8046,N_4945,N_1016);
nor U8047 (N_8047,N_4938,N_4965);
and U8048 (N_8048,N_2932,N_4416);
and U8049 (N_8049,N_4838,N_2700);
xnor U8050 (N_8050,N_368,N_3027);
or U8051 (N_8051,N_4051,N_983);
nor U8052 (N_8052,N_3954,N_4911);
xnor U8053 (N_8053,N_3843,N_2375);
nor U8054 (N_8054,N_2627,N_392);
nor U8055 (N_8055,N_714,N_604);
nand U8056 (N_8056,N_695,N_4105);
nor U8057 (N_8057,N_4111,N_3537);
and U8058 (N_8058,N_2158,N_3801);
or U8059 (N_8059,N_564,N_1151);
xnor U8060 (N_8060,N_4246,N_2554);
xnor U8061 (N_8061,N_1203,N_4229);
nor U8062 (N_8062,N_1341,N_2959);
and U8063 (N_8063,N_2879,N_3081);
nand U8064 (N_8064,N_3458,N_3531);
nor U8065 (N_8065,N_4151,N_3996);
nor U8066 (N_8066,N_1428,N_3835);
or U8067 (N_8067,N_4884,N_981);
nor U8068 (N_8068,N_3704,N_3526);
and U8069 (N_8069,N_125,N_271);
xor U8070 (N_8070,N_1345,N_2137);
and U8071 (N_8071,N_1545,N_4338);
xor U8072 (N_8072,N_618,N_915);
xor U8073 (N_8073,N_3117,N_656);
nand U8074 (N_8074,N_1011,N_4039);
or U8075 (N_8075,N_1928,N_2613);
or U8076 (N_8076,N_2767,N_2860);
and U8077 (N_8077,N_975,N_3592);
xor U8078 (N_8078,N_256,N_1570);
and U8079 (N_8079,N_3193,N_4382);
and U8080 (N_8080,N_3740,N_4840);
xor U8081 (N_8081,N_3554,N_277);
nand U8082 (N_8082,N_3602,N_4447);
or U8083 (N_8083,N_4861,N_1334);
and U8084 (N_8084,N_2306,N_4305);
xor U8085 (N_8085,N_2209,N_863);
nor U8086 (N_8086,N_65,N_3459);
nor U8087 (N_8087,N_1513,N_985);
nand U8088 (N_8088,N_3433,N_1543);
nand U8089 (N_8089,N_3782,N_4163);
or U8090 (N_8090,N_3115,N_1099);
xnor U8091 (N_8091,N_4913,N_1724);
nand U8092 (N_8092,N_3886,N_4730);
nor U8093 (N_8093,N_1436,N_586);
and U8094 (N_8094,N_807,N_4435);
nand U8095 (N_8095,N_436,N_773);
and U8096 (N_8096,N_4637,N_751);
nand U8097 (N_8097,N_762,N_1875);
nor U8098 (N_8098,N_1285,N_1662);
nand U8099 (N_8099,N_1910,N_4482);
xor U8100 (N_8100,N_2420,N_4897);
xnor U8101 (N_8101,N_1539,N_3702);
and U8102 (N_8102,N_3741,N_3937);
or U8103 (N_8103,N_4594,N_4926);
and U8104 (N_8104,N_1868,N_1207);
or U8105 (N_8105,N_4374,N_2329);
or U8106 (N_8106,N_4272,N_4534);
or U8107 (N_8107,N_2387,N_141);
xor U8108 (N_8108,N_1828,N_2472);
and U8109 (N_8109,N_2628,N_1478);
nor U8110 (N_8110,N_320,N_2101);
nor U8111 (N_8111,N_2535,N_4325);
nor U8112 (N_8112,N_2344,N_3726);
xor U8113 (N_8113,N_1414,N_1190);
nand U8114 (N_8114,N_3440,N_1462);
nor U8115 (N_8115,N_161,N_856);
nor U8116 (N_8116,N_3690,N_1788);
and U8117 (N_8117,N_4647,N_4895);
or U8118 (N_8118,N_632,N_261);
or U8119 (N_8119,N_2365,N_1665);
xnor U8120 (N_8120,N_611,N_3887);
nor U8121 (N_8121,N_3706,N_921);
nand U8122 (N_8122,N_4017,N_1314);
nand U8123 (N_8123,N_497,N_4404);
and U8124 (N_8124,N_1709,N_1819);
or U8125 (N_8125,N_884,N_2722);
xor U8126 (N_8126,N_4776,N_327);
and U8127 (N_8127,N_1834,N_4200);
xnor U8128 (N_8128,N_4889,N_4205);
and U8129 (N_8129,N_2426,N_4168);
nor U8130 (N_8130,N_1442,N_331);
nand U8131 (N_8131,N_1870,N_699);
and U8132 (N_8132,N_4023,N_3806);
xnor U8133 (N_8133,N_46,N_3945);
nand U8134 (N_8134,N_3533,N_1508);
nand U8135 (N_8135,N_4975,N_1340);
xnor U8136 (N_8136,N_826,N_410);
nor U8137 (N_8137,N_4428,N_3048);
nand U8138 (N_8138,N_1752,N_4817);
or U8139 (N_8139,N_4,N_3677);
nor U8140 (N_8140,N_666,N_875);
xnor U8141 (N_8141,N_20,N_4069);
and U8142 (N_8142,N_3084,N_4086);
xnor U8143 (N_8143,N_936,N_3597);
nand U8144 (N_8144,N_3048,N_3045);
and U8145 (N_8145,N_4959,N_3577);
and U8146 (N_8146,N_4625,N_2649);
nor U8147 (N_8147,N_2194,N_178);
nand U8148 (N_8148,N_234,N_3267);
or U8149 (N_8149,N_1745,N_3220);
xnor U8150 (N_8150,N_3260,N_1584);
xnor U8151 (N_8151,N_2284,N_2736);
or U8152 (N_8152,N_4484,N_1818);
xnor U8153 (N_8153,N_1560,N_266);
nor U8154 (N_8154,N_229,N_2537);
nor U8155 (N_8155,N_3596,N_4999);
nand U8156 (N_8156,N_3540,N_1979);
xnor U8157 (N_8157,N_2642,N_573);
and U8158 (N_8158,N_1535,N_801);
xnor U8159 (N_8159,N_1087,N_1928);
xnor U8160 (N_8160,N_476,N_1123);
or U8161 (N_8161,N_1416,N_4067);
xor U8162 (N_8162,N_1647,N_1518);
and U8163 (N_8163,N_1331,N_1979);
or U8164 (N_8164,N_4302,N_209);
and U8165 (N_8165,N_763,N_2703);
nand U8166 (N_8166,N_1068,N_3012);
xnor U8167 (N_8167,N_4645,N_2159);
and U8168 (N_8168,N_2213,N_819);
or U8169 (N_8169,N_1160,N_2639);
nand U8170 (N_8170,N_3613,N_3114);
or U8171 (N_8171,N_628,N_3394);
or U8172 (N_8172,N_505,N_1036);
and U8173 (N_8173,N_4753,N_4127);
or U8174 (N_8174,N_3298,N_912);
nand U8175 (N_8175,N_2096,N_3189);
nand U8176 (N_8176,N_2729,N_4095);
nand U8177 (N_8177,N_4460,N_4937);
xnor U8178 (N_8178,N_3943,N_2245);
and U8179 (N_8179,N_837,N_2825);
nand U8180 (N_8180,N_1675,N_1373);
nor U8181 (N_8181,N_405,N_88);
xnor U8182 (N_8182,N_4373,N_4749);
nand U8183 (N_8183,N_4204,N_4720);
and U8184 (N_8184,N_4583,N_1434);
or U8185 (N_8185,N_4739,N_561);
nand U8186 (N_8186,N_3750,N_4596);
and U8187 (N_8187,N_2344,N_3776);
or U8188 (N_8188,N_1523,N_152);
or U8189 (N_8189,N_3235,N_4606);
nor U8190 (N_8190,N_303,N_4840);
nand U8191 (N_8191,N_4991,N_3096);
and U8192 (N_8192,N_3364,N_1797);
nand U8193 (N_8193,N_280,N_3740);
nor U8194 (N_8194,N_4443,N_1797);
and U8195 (N_8195,N_293,N_2837);
nor U8196 (N_8196,N_2631,N_2398);
or U8197 (N_8197,N_1768,N_3489);
xnor U8198 (N_8198,N_1508,N_3864);
and U8199 (N_8199,N_4017,N_4286);
nand U8200 (N_8200,N_621,N_4465);
or U8201 (N_8201,N_2224,N_1729);
nor U8202 (N_8202,N_4090,N_343);
xor U8203 (N_8203,N_1944,N_135);
nand U8204 (N_8204,N_4882,N_3818);
nand U8205 (N_8205,N_3348,N_180);
nor U8206 (N_8206,N_521,N_4364);
nand U8207 (N_8207,N_4960,N_1636);
nor U8208 (N_8208,N_3466,N_1750);
nand U8209 (N_8209,N_2835,N_3596);
xor U8210 (N_8210,N_2774,N_4596);
nand U8211 (N_8211,N_1306,N_3824);
and U8212 (N_8212,N_4643,N_2901);
xnor U8213 (N_8213,N_2000,N_649);
and U8214 (N_8214,N_2288,N_348);
and U8215 (N_8215,N_4302,N_517);
nor U8216 (N_8216,N_4301,N_1129);
xnor U8217 (N_8217,N_2735,N_820);
nand U8218 (N_8218,N_1789,N_4318);
and U8219 (N_8219,N_3650,N_4372);
and U8220 (N_8220,N_1057,N_3013);
nand U8221 (N_8221,N_3274,N_618);
nand U8222 (N_8222,N_491,N_3567);
nor U8223 (N_8223,N_4644,N_2728);
and U8224 (N_8224,N_4116,N_2662);
or U8225 (N_8225,N_3761,N_1368);
xnor U8226 (N_8226,N_3733,N_4819);
xor U8227 (N_8227,N_946,N_3230);
nand U8228 (N_8228,N_592,N_1708);
nand U8229 (N_8229,N_2440,N_2025);
and U8230 (N_8230,N_1941,N_1818);
xnor U8231 (N_8231,N_2537,N_1397);
and U8232 (N_8232,N_2515,N_4445);
nor U8233 (N_8233,N_2815,N_4364);
xnor U8234 (N_8234,N_1994,N_4971);
nor U8235 (N_8235,N_517,N_3014);
nor U8236 (N_8236,N_667,N_1805);
or U8237 (N_8237,N_4415,N_2892);
or U8238 (N_8238,N_4454,N_1040);
or U8239 (N_8239,N_4951,N_2784);
nand U8240 (N_8240,N_3314,N_690);
xnor U8241 (N_8241,N_4868,N_614);
xor U8242 (N_8242,N_192,N_3433);
nor U8243 (N_8243,N_1666,N_2515);
or U8244 (N_8244,N_3580,N_4999);
or U8245 (N_8245,N_4719,N_2791);
nor U8246 (N_8246,N_2446,N_715);
xor U8247 (N_8247,N_1458,N_382);
nor U8248 (N_8248,N_4248,N_3460);
or U8249 (N_8249,N_2280,N_3587);
xnor U8250 (N_8250,N_574,N_3664);
and U8251 (N_8251,N_2613,N_1624);
nand U8252 (N_8252,N_3171,N_2730);
xnor U8253 (N_8253,N_4083,N_4782);
and U8254 (N_8254,N_1252,N_3394);
nor U8255 (N_8255,N_2498,N_2679);
nand U8256 (N_8256,N_3763,N_2009);
or U8257 (N_8257,N_704,N_2961);
xor U8258 (N_8258,N_1502,N_760);
or U8259 (N_8259,N_3599,N_2965);
or U8260 (N_8260,N_3104,N_1069);
nand U8261 (N_8261,N_4958,N_1481);
nand U8262 (N_8262,N_2972,N_1724);
and U8263 (N_8263,N_1061,N_3780);
nand U8264 (N_8264,N_2672,N_2067);
and U8265 (N_8265,N_3386,N_4596);
and U8266 (N_8266,N_1951,N_3186);
nor U8267 (N_8267,N_1790,N_852);
xor U8268 (N_8268,N_2045,N_579);
nor U8269 (N_8269,N_534,N_1523);
xor U8270 (N_8270,N_3159,N_1530);
nor U8271 (N_8271,N_3527,N_2394);
and U8272 (N_8272,N_4114,N_1959);
nor U8273 (N_8273,N_2190,N_3225);
nand U8274 (N_8274,N_3610,N_1245);
or U8275 (N_8275,N_2616,N_2355);
nand U8276 (N_8276,N_503,N_2595);
xor U8277 (N_8277,N_2978,N_4712);
and U8278 (N_8278,N_2144,N_4196);
nand U8279 (N_8279,N_3968,N_4999);
nor U8280 (N_8280,N_4982,N_838);
and U8281 (N_8281,N_2912,N_4359);
xor U8282 (N_8282,N_2203,N_1792);
or U8283 (N_8283,N_610,N_2047);
nand U8284 (N_8284,N_3637,N_3310);
and U8285 (N_8285,N_3713,N_4916);
nand U8286 (N_8286,N_4502,N_2417);
and U8287 (N_8287,N_2782,N_2721);
and U8288 (N_8288,N_2960,N_281);
xor U8289 (N_8289,N_3047,N_1530);
nor U8290 (N_8290,N_3235,N_3165);
xor U8291 (N_8291,N_2678,N_1307);
xnor U8292 (N_8292,N_4018,N_342);
nand U8293 (N_8293,N_3272,N_3375);
xnor U8294 (N_8294,N_989,N_1173);
and U8295 (N_8295,N_2589,N_4589);
and U8296 (N_8296,N_4394,N_4340);
or U8297 (N_8297,N_3707,N_4747);
nand U8298 (N_8298,N_4550,N_4799);
or U8299 (N_8299,N_1406,N_1197);
nor U8300 (N_8300,N_4203,N_3448);
nand U8301 (N_8301,N_3674,N_2928);
and U8302 (N_8302,N_1941,N_1664);
nor U8303 (N_8303,N_3341,N_1529);
and U8304 (N_8304,N_3858,N_3635);
or U8305 (N_8305,N_2742,N_509);
nand U8306 (N_8306,N_1968,N_1697);
and U8307 (N_8307,N_2702,N_1795);
and U8308 (N_8308,N_61,N_422);
nand U8309 (N_8309,N_4968,N_3465);
nand U8310 (N_8310,N_2984,N_4880);
and U8311 (N_8311,N_4304,N_3243);
xor U8312 (N_8312,N_2568,N_1916);
nand U8313 (N_8313,N_428,N_4936);
and U8314 (N_8314,N_2870,N_1586);
and U8315 (N_8315,N_586,N_804);
or U8316 (N_8316,N_1014,N_2968);
or U8317 (N_8317,N_2950,N_801);
nor U8318 (N_8318,N_3151,N_926);
and U8319 (N_8319,N_3436,N_4552);
nor U8320 (N_8320,N_4205,N_4885);
nand U8321 (N_8321,N_32,N_3056);
or U8322 (N_8322,N_3067,N_1461);
and U8323 (N_8323,N_3611,N_4592);
or U8324 (N_8324,N_1089,N_4147);
nor U8325 (N_8325,N_3956,N_4380);
nor U8326 (N_8326,N_616,N_3549);
nand U8327 (N_8327,N_3368,N_2187);
and U8328 (N_8328,N_3888,N_4995);
and U8329 (N_8329,N_225,N_4418);
xnor U8330 (N_8330,N_2689,N_4844);
or U8331 (N_8331,N_4479,N_686);
nand U8332 (N_8332,N_3714,N_4212);
nor U8333 (N_8333,N_1979,N_3448);
nand U8334 (N_8334,N_3223,N_2024);
nor U8335 (N_8335,N_223,N_3842);
and U8336 (N_8336,N_3197,N_4277);
and U8337 (N_8337,N_1015,N_3077);
nor U8338 (N_8338,N_2140,N_2977);
xor U8339 (N_8339,N_3285,N_4219);
xnor U8340 (N_8340,N_477,N_1691);
xor U8341 (N_8341,N_854,N_4155);
nor U8342 (N_8342,N_399,N_3390);
xnor U8343 (N_8343,N_4383,N_3329);
or U8344 (N_8344,N_1004,N_1098);
and U8345 (N_8345,N_4643,N_1636);
and U8346 (N_8346,N_670,N_775);
xor U8347 (N_8347,N_3428,N_2648);
nor U8348 (N_8348,N_2303,N_1911);
nor U8349 (N_8349,N_1698,N_4450);
and U8350 (N_8350,N_4064,N_1166);
nand U8351 (N_8351,N_3583,N_2022);
nand U8352 (N_8352,N_465,N_318);
and U8353 (N_8353,N_2258,N_4302);
or U8354 (N_8354,N_4754,N_3006);
nor U8355 (N_8355,N_1453,N_2648);
nor U8356 (N_8356,N_237,N_4010);
xor U8357 (N_8357,N_3596,N_822);
xor U8358 (N_8358,N_1850,N_516);
nand U8359 (N_8359,N_4267,N_2849);
and U8360 (N_8360,N_3424,N_2632);
nor U8361 (N_8361,N_4074,N_1172);
nor U8362 (N_8362,N_1231,N_3037);
and U8363 (N_8363,N_4949,N_2933);
and U8364 (N_8364,N_2281,N_1839);
and U8365 (N_8365,N_469,N_1179);
or U8366 (N_8366,N_1044,N_4758);
and U8367 (N_8367,N_2366,N_2459);
xor U8368 (N_8368,N_1529,N_4658);
nor U8369 (N_8369,N_3661,N_3702);
nor U8370 (N_8370,N_317,N_1712);
nor U8371 (N_8371,N_3836,N_1144);
xnor U8372 (N_8372,N_3103,N_797);
or U8373 (N_8373,N_2157,N_3250);
xnor U8374 (N_8374,N_3484,N_2926);
or U8375 (N_8375,N_459,N_4706);
or U8376 (N_8376,N_2184,N_1930);
nand U8377 (N_8377,N_93,N_718);
nand U8378 (N_8378,N_1500,N_3450);
and U8379 (N_8379,N_2366,N_1086);
nor U8380 (N_8380,N_2289,N_781);
nand U8381 (N_8381,N_3987,N_4904);
or U8382 (N_8382,N_4131,N_1989);
or U8383 (N_8383,N_915,N_2515);
nand U8384 (N_8384,N_3861,N_3972);
nand U8385 (N_8385,N_3475,N_1143);
or U8386 (N_8386,N_1811,N_4154);
and U8387 (N_8387,N_1968,N_2440);
xnor U8388 (N_8388,N_4194,N_4291);
nor U8389 (N_8389,N_1955,N_181);
nand U8390 (N_8390,N_1727,N_1971);
or U8391 (N_8391,N_1029,N_3464);
or U8392 (N_8392,N_2532,N_2761);
nor U8393 (N_8393,N_4613,N_4701);
and U8394 (N_8394,N_1486,N_4927);
nand U8395 (N_8395,N_3041,N_1228);
nand U8396 (N_8396,N_933,N_4234);
xnor U8397 (N_8397,N_2518,N_2780);
and U8398 (N_8398,N_939,N_3751);
and U8399 (N_8399,N_4838,N_2119);
or U8400 (N_8400,N_356,N_4809);
nor U8401 (N_8401,N_4727,N_2525);
and U8402 (N_8402,N_2322,N_854);
or U8403 (N_8403,N_4557,N_110);
and U8404 (N_8404,N_3527,N_1048);
or U8405 (N_8405,N_891,N_3765);
and U8406 (N_8406,N_385,N_3672);
nor U8407 (N_8407,N_4315,N_4851);
or U8408 (N_8408,N_2824,N_4884);
and U8409 (N_8409,N_3642,N_1256);
nor U8410 (N_8410,N_1520,N_1424);
nor U8411 (N_8411,N_2935,N_4255);
or U8412 (N_8412,N_4109,N_2636);
nand U8413 (N_8413,N_1163,N_533);
or U8414 (N_8414,N_346,N_3922);
xnor U8415 (N_8415,N_2903,N_1800);
and U8416 (N_8416,N_3984,N_814);
nor U8417 (N_8417,N_2587,N_3450);
and U8418 (N_8418,N_4212,N_418);
and U8419 (N_8419,N_4422,N_991);
nand U8420 (N_8420,N_3044,N_1998);
nand U8421 (N_8421,N_4472,N_71);
and U8422 (N_8422,N_3175,N_1876);
and U8423 (N_8423,N_4346,N_2784);
nand U8424 (N_8424,N_4082,N_3774);
nor U8425 (N_8425,N_560,N_3942);
or U8426 (N_8426,N_2121,N_2963);
nor U8427 (N_8427,N_2388,N_78);
and U8428 (N_8428,N_961,N_4635);
xor U8429 (N_8429,N_2823,N_2581);
nand U8430 (N_8430,N_421,N_1793);
nor U8431 (N_8431,N_3018,N_3265);
and U8432 (N_8432,N_2261,N_3178);
xor U8433 (N_8433,N_4907,N_1604);
or U8434 (N_8434,N_4766,N_4697);
or U8435 (N_8435,N_388,N_1827);
nand U8436 (N_8436,N_315,N_189);
nand U8437 (N_8437,N_4412,N_3738);
nor U8438 (N_8438,N_311,N_4987);
nor U8439 (N_8439,N_2508,N_2779);
xnor U8440 (N_8440,N_1563,N_941);
or U8441 (N_8441,N_3225,N_508);
nor U8442 (N_8442,N_2094,N_97);
nor U8443 (N_8443,N_819,N_875);
and U8444 (N_8444,N_1150,N_402);
xnor U8445 (N_8445,N_3261,N_4246);
nand U8446 (N_8446,N_2245,N_2442);
nor U8447 (N_8447,N_3558,N_2906);
or U8448 (N_8448,N_1570,N_1749);
nor U8449 (N_8449,N_1886,N_4544);
nand U8450 (N_8450,N_263,N_2098);
nand U8451 (N_8451,N_3750,N_4866);
nor U8452 (N_8452,N_55,N_1902);
nor U8453 (N_8453,N_4965,N_3094);
nand U8454 (N_8454,N_3009,N_717);
and U8455 (N_8455,N_1253,N_2794);
and U8456 (N_8456,N_1733,N_2189);
nand U8457 (N_8457,N_4784,N_343);
or U8458 (N_8458,N_1599,N_2514);
or U8459 (N_8459,N_4071,N_1390);
xor U8460 (N_8460,N_1113,N_2279);
nor U8461 (N_8461,N_52,N_1255);
xor U8462 (N_8462,N_1327,N_499);
nand U8463 (N_8463,N_1156,N_2164);
nor U8464 (N_8464,N_1633,N_922);
xnor U8465 (N_8465,N_2726,N_4523);
nand U8466 (N_8466,N_1933,N_3103);
and U8467 (N_8467,N_1522,N_885);
nand U8468 (N_8468,N_4460,N_2793);
or U8469 (N_8469,N_2292,N_4868);
and U8470 (N_8470,N_323,N_2869);
nor U8471 (N_8471,N_47,N_3148);
xnor U8472 (N_8472,N_1391,N_4914);
nor U8473 (N_8473,N_389,N_4730);
xor U8474 (N_8474,N_4070,N_2125);
xor U8475 (N_8475,N_4375,N_2673);
nand U8476 (N_8476,N_2545,N_41);
nand U8477 (N_8477,N_3505,N_1899);
xor U8478 (N_8478,N_3865,N_4632);
xnor U8479 (N_8479,N_4720,N_1977);
or U8480 (N_8480,N_1200,N_4190);
or U8481 (N_8481,N_3956,N_1997);
xnor U8482 (N_8482,N_4304,N_4384);
xnor U8483 (N_8483,N_1558,N_2801);
xor U8484 (N_8484,N_4395,N_4846);
or U8485 (N_8485,N_2541,N_4233);
nor U8486 (N_8486,N_215,N_3337);
and U8487 (N_8487,N_2650,N_2867);
xor U8488 (N_8488,N_828,N_1996);
xnor U8489 (N_8489,N_3732,N_1613);
or U8490 (N_8490,N_2717,N_4080);
or U8491 (N_8491,N_1583,N_4331);
xnor U8492 (N_8492,N_2244,N_1861);
and U8493 (N_8493,N_4738,N_2293);
nand U8494 (N_8494,N_1089,N_2127);
nor U8495 (N_8495,N_3708,N_3861);
or U8496 (N_8496,N_4776,N_2314);
or U8497 (N_8497,N_4695,N_1760);
and U8498 (N_8498,N_393,N_4892);
nand U8499 (N_8499,N_1974,N_4053);
and U8500 (N_8500,N_4416,N_2151);
nor U8501 (N_8501,N_3885,N_4125);
nor U8502 (N_8502,N_1071,N_3991);
xor U8503 (N_8503,N_1884,N_3461);
and U8504 (N_8504,N_3765,N_1876);
and U8505 (N_8505,N_220,N_4501);
and U8506 (N_8506,N_3078,N_189);
and U8507 (N_8507,N_3924,N_4082);
or U8508 (N_8508,N_705,N_1097);
or U8509 (N_8509,N_88,N_2402);
nand U8510 (N_8510,N_576,N_4045);
nor U8511 (N_8511,N_1462,N_4794);
xor U8512 (N_8512,N_2704,N_2662);
nor U8513 (N_8513,N_4636,N_1625);
nand U8514 (N_8514,N_135,N_1581);
and U8515 (N_8515,N_3842,N_2511);
nor U8516 (N_8516,N_1557,N_2046);
xnor U8517 (N_8517,N_292,N_1785);
or U8518 (N_8518,N_4109,N_2714);
nand U8519 (N_8519,N_1324,N_994);
or U8520 (N_8520,N_1627,N_450);
and U8521 (N_8521,N_553,N_1199);
nor U8522 (N_8522,N_1957,N_3551);
nor U8523 (N_8523,N_4549,N_2705);
or U8524 (N_8524,N_4172,N_1944);
or U8525 (N_8525,N_3720,N_3483);
xor U8526 (N_8526,N_1603,N_2973);
and U8527 (N_8527,N_187,N_4759);
and U8528 (N_8528,N_2710,N_1980);
or U8529 (N_8529,N_3648,N_2438);
nand U8530 (N_8530,N_1352,N_2232);
nor U8531 (N_8531,N_2238,N_3522);
nand U8532 (N_8532,N_786,N_1177);
nand U8533 (N_8533,N_996,N_2279);
and U8534 (N_8534,N_4697,N_2640);
or U8535 (N_8535,N_4108,N_559);
and U8536 (N_8536,N_2517,N_2201);
or U8537 (N_8537,N_2151,N_3596);
nand U8538 (N_8538,N_2673,N_3989);
or U8539 (N_8539,N_1833,N_575);
and U8540 (N_8540,N_2550,N_2237);
nor U8541 (N_8541,N_3175,N_4377);
and U8542 (N_8542,N_374,N_4251);
nor U8543 (N_8543,N_4889,N_2287);
or U8544 (N_8544,N_3822,N_186);
nor U8545 (N_8545,N_1964,N_2432);
nor U8546 (N_8546,N_2380,N_684);
or U8547 (N_8547,N_2959,N_3106);
nand U8548 (N_8548,N_4909,N_4301);
and U8549 (N_8549,N_3558,N_1390);
nor U8550 (N_8550,N_758,N_3904);
nor U8551 (N_8551,N_3382,N_255);
xor U8552 (N_8552,N_4489,N_1921);
nor U8553 (N_8553,N_1355,N_4171);
xor U8554 (N_8554,N_1362,N_362);
xor U8555 (N_8555,N_2425,N_3137);
and U8556 (N_8556,N_4296,N_4026);
nand U8557 (N_8557,N_2106,N_2460);
or U8558 (N_8558,N_892,N_1119);
nor U8559 (N_8559,N_259,N_300);
or U8560 (N_8560,N_4983,N_919);
and U8561 (N_8561,N_628,N_3637);
or U8562 (N_8562,N_2664,N_2592);
xor U8563 (N_8563,N_2526,N_566);
nand U8564 (N_8564,N_3536,N_22);
nand U8565 (N_8565,N_3775,N_3849);
or U8566 (N_8566,N_3854,N_73);
and U8567 (N_8567,N_4156,N_3415);
and U8568 (N_8568,N_990,N_1175);
and U8569 (N_8569,N_3239,N_2837);
nand U8570 (N_8570,N_2302,N_1387);
xor U8571 (N_8571,N_1950,N_4991);
nor U8572 (N_8572,N_1752,N_1463);
nand U8573 (N_8573,N_4492,N_2079);
xor U8574 (N_8574,N_4558,N_677);
nor U8575 (N_8575,N_3068,N_3215);
nand U8576 (N_8576,N_435,N_1439);
and U8577 (N_8577,N_2331,N_4012);
and U8578 (N_8578,N_1752,N_2743);
nor U8579 (N_8579,N_1520,N_1075);
nand U8580 (N_8580,N_2621,N_4554);
nor U8581 (N_8581,N_151,N_2993);
xor U8582 (N_8582,N_3633,N_3801);
nor U8583 (N_8583,N_1498,N_516);
nand U8584 (N_8584,N_4108,N_1709);
nor U8585 (N_8585,N_3364,N_2462);
nor U8586 (N_8586,N_3180,N_1907);
and U8587 (N_8587,N_4059,N_4308);
xor U8588 (N_8588,N_3138,N_76);
nor U8589 (N_8589,N_499,N_819);
or U8590 (N_8590,N_1069,N_1856);
or U8591 (N_8591,N_2843,N_1088);
or U8592 (N_8592,N_2895,N_4944);
or U8593 (N_8593,N_4252,N_830);
nand U8594 (N_8594,N_3173,N_1679);
and U8595 (N_8595,N_4183,N_3668);
nand U8596 (N_8596,N_3329,N_1919);
nand U8597 (N_8597,N_978,N_3633);
and U8598 (N_8598,N_2871,N_2302);
nand U8599 (N_8599,N_1224,N_486);
and U8600 (N_8600,N_4692,N_339);
xnor U8601 (N_8601,N_3612,N_3659);
or U8602 (N_8602,N_357,N_1249);
and U8603 (N_8603,N_1137,N_1520);
or U8604 (N_8604,N_4363,N_3301);
nand U8605 (N_8605,N_1864,N_1922);
or U8606 (N_8606,N_3297,N_4186);
xnor U8607 (N_8607,N_1917,N_3955);
and U8608 (N_8608,N_2303,N_1577);
and U8609 (N_8609,N_2033,N_2468);
xor U8610 (N_8610,N_4601,N_1973);
and U8611 (N_8611,N_1877,N_1272);
and U8612 (N_8612,N_773,N_4698);
or U8613 (N_8613,N_4704,N_2510);
xor U8614 (N_8614,N_2700,N_1565);
and U8615 (N_8615,N_694,N_4098);
nor U8616 (N_8616,N_1826,N_382);
nand U8617 (N_8617,N_1822,N_2510);
xnor U8618 (N_8618,N_629,N_4120);
or U8619 (N_8619,N_2742,N_2221);
xor U8620 (N_8620,N_1063,N_506);
nor U8621 (N_8621,N_1460,N_4082);
xor U8622 (N_8622,N_2481,N_1134);
or U8623 (N_8623,N_139,N_2138);
or U8624 (N_8624,N_625,N_3385);
nand U8625 (N_8625,N_3383,N_2000);
or U8626 (N_8626,N_938,N_4393);
nand U8627 (N_8627,N_595,N_4711);
xnor U8628 (N_8628,N_4023,N_4725);
or U8629 (N_8629,N_2585,N_2717);
or U8630 (N_8630,N_797,N_4287);
nand U8631 (N_8631,N_1166,N_4848);
and U8632 (N_8632,N_2581,N_1294);
or U8633 (N_8633,N_713,N_1686);
nor U8634 (N_8634,N_3120,N_3015);
and U8635 (N_8635,N_2881,N_4185);
nand U8636 (N_8636,N_2648,N_2258);
nand U8637 (N_8637,N_1626,N_45);
and U8638 (N_8638,N_1821,N_3878);
or U8639 (N_8639,N_989,N_550);
and U8640 (N_8640,N_3882,N_4837);
nand U8641 (N_8641,N_1796,N_3730);
or U8642 (N_8642,N_1536,N_582);
nor U8643 (N_8643,N_2618,N_4370);
nand U8644 (N_8644,N_2888,N_2442);
nor U8645 (N_8645,N_3615,N_645);
and U8646 (N_8646,N_3102,N_2049);
nand U8647 (N_8647,N_4806,N_4788);
or U8648 (N_8648,N_1820,N_3674);
nor U8649 (N_8649,N_4651,N_3535);
or U8650 (N_8650,N_4240,N_3029);
and U8651 (N_8651,N_894,N_2708);
nand U8652 (N_8652,N_2127,N_1062);
nand U8653 (N_8653,N_3143,N_481);
and U8654 (N_8654,N_2132,N_1916);
and U8655 (N_8655,N_67,N_1315);
nand U8656 (N_8656,N_4344,N_3202);
nor U8657 (N_8657,N_1853,N_1525);
nor U8658 (N_8658,N_2392,N_3799);
xor U8659 (N_8659,N_290,N_4019);
or U8660 (N_8660,N_1840,N_4753);
or U8661 (N_8661,N_2436,N_4222);
nand U8662 (N_8662,N_4398,N_4468);
or U8663 (N_8663,N_937,N_1969);
or U8664 (N_8664,N_1658,N_102);
and U8665 (N_8665,N_3538,N_127);
xor U8666 (N_8666,N_3881,N_4296);
and U8667 (N_8667,N_4631,N_2313);
nand U8668 (N_8668,N_2295,N_330);
or U8669 (N_8669,N_4020,N_4015);
xor U8670 (N_8670,N_216,N_258);
nor U8671 (N_8671,N_2421,N_4990);
and U8672 (N_8672,N_3021,N_428);
nand U8673 (N_8673,N_3535,N_2162);
or U8674 (N_8674,N_494,N_3134);
and U8675 (N_8675,N_2187,N_4670);
nor U8676 (N_8676,N_1915,N_1763);
and U8677 (N_8677,N_1742,N_521);
or U8678 (N_8678,N_978,N_85);
or U8679 (N_8679,N_2947,N_2281);
nand U8680 (N_8680,N_1126,N_4125);
and U8681 (N_8681,N_2247,N_2495);
and U8682 (N_8682,N_3576,N_4043);
xnor U8683 (N_8683,N_1428,N_696);
xnor U8684 (N_8684,N_1032,N_2691);
nor U8685 (N_8685,N_2226,N_3190);
xor U8686 (N_8686,N_4530,N_3037);
and U8687 (N_8687,N_3561,N_2331);
nand U8688 (N_8688,N_1609,N_3966);
nor U8689 (N_8689,N_2128,N_3839);
xor U8690 (N_8690,N_1238,N_4822);
nor U8691 (N_8691,N_2150,N_4675);
nand U8692 (N_8692,N_2597,N_2920);
xor U8693 (N_8693,N_2519,N_3963);
nand U8694 (N_8694,N_1051,N_3306);
or U8695 (N_8695,N_3495,N_3909);
nand U8696 (N_8696,N_3227,N_4551);
xor U8697 (N_8697,N_3742,N_4476);
nor U8698 (N_8698,N_3683,N_1015);
xnor U8699 (N_8699,N_3879,N_707);
nand U8700 (N_8700,N_4603,N_1376);
nand U8701 (N_8701,N_1520,N_4101);
xor U8702 (N_8702,N_148,N_799);
and U8703 (N_8703,N_2327,N_592);
nand U8704 (N_8704,N_3628,N_4437);
xnor U8705 (N_8705,N_31,N_4384);
nand U8706 (N_8706,N_1534,N_3978);
and U8707 (N_8707,N_1738,N_4449);
xnor U8708 (N_8708,N_852,N_2189);
nor U8709 (N_8709,N_4582,N_4084);
nand U8710 (N_8710,N_1729,N_2736);
nand U8711 (N_8711,N_2275,N_2382);
nor U8712 (N_8712,N_981,N_3667);
nor U8713 (N_8713,N_3762,N_3741);
nor U8714 (N_8714,N_139,N_562);
nor U8715 (N_8715,N_1346,N_141);
and U8716 (N_8716,N_1254,N_1231);
and U8717 (N_8717,N_2342,N_3907);
nand U8718 (N_8718,N_710,N_3395);
or U8719 (N_8719,N_1082,N_565);
and U8720 (N_8720,N_4463,N_3967);
nor U8721 (N_8721,N_910,N_3881);
xnor U8722 (N_8722,N_2588,N_649);
or U8723 (N_8723,N_2191,N_3029);
nor U8724 (N_8724,N_1173,N_4871);
or U8725 (N_8725,N_2347,N_2080);
and U8726 (N_8726,N_2576,N_2653);
nor U8727 (N_8727,N_381,N_4379);
nand U8728 (N_8728,N_2734,N_629);
and U8729 (N_8729,N_42,N_1756);
or U8730 (N_8730,N_3163,N_108);
and U8731 (N_8731,N_2268,N_9);
or U8732 (N_8732,N_3041,N_979);
nand U8733 (N_8733,N_4646,N_3825);
xnor U8734 (N_8734,N_329,N_215);
and U8735 (N_8735,N_4375,N_3202);
and U8736 (N_8736,N_4163,N_4085);
nor U8737 (N_8737,N_3661,N_4772);
xor U8738 (N_8738,N_3242,N_4528);
xnor U8739 (N_8739,N_2709,N_677);
nand U8740 (N_8740,N_3191,N_3746);
and U8741 (N_8741,N_4085,N_2156);
or U8742 (N_8742,N_1339,N_1198);
xnor U8743 (N_8743,N_1737,N_2061);
nor U8744 (N_8744,N_167,N_3977);
xnor U8745 (N_8745,N_4737,N_3789);
and U8746 (N_8746,N_200,N_2266);
and U8747 (N_8747,N_201,N_1968);
nand U8748 (N_8748,N_1414,N_1952);
nand U8749 (N_8749,N_12,N_4917);
or U8750 (N_8750,N_4717,N_3032);
or U8751 (N_8751,N_1753,N_1892);
xor U8752 (N_8752,N_4374,N_1470);
nand U8753 (N_8753,N_148,N_4343);
or U8754 (N_8754,N_4333,N_1359);
and U8755 (N_8755,N_4984,N_3605);
and U8756 (N_8756,N_1725,N_1432);
nor U8757 (N_8757,N_620,N_4514);
nand U8758 (N_8758,N_4061,N_675);
and U8759 (N_8759,N_606,N_3580);
nand U8760 (N_8760,N_4230,N_332);
nor U8761 (N_8761,N_3578,N_2317);
xnor U8762 (N_8762,N_2372,N_2340);
or U8763 (N_8763,N_4515,N_1238);
nor U8764 (N_8764,N_3052,N_10);
nor U8765 (N_8765,N_4483,N_155);
xnor U8766 (N_8766,N_246,N_1294);
and U8767 (N_8767,N_3439,N_1620);
xnor U8768 (N_8768,N_588,N_2862);
nor U8769 (N_8769,N_2700,N_2154);
xor U8770 (N_8770,N_2810,N_1787);
xor U8771 (N_8771,N_4686,N_4486);
nor U8772 (N_8772,N_3590,N_4671);
nand U8773 (N_8773,N_4705,N_3240);
nand U8774 (N_8774,N_3772,N_2974);
nand U8775 (N_8775,N_4691,N_3897);
or U8776 (N_8776,N_4568,N_3475);
nand U8777 (N_8777,N_4998,N_3074);
xnor U8778 (N_8778,N_93,N_1224);
nand U8779 (N_8779,N_1472,N_972);
or U8780 (N_8780,N_4899,N_4247);
xor U8781 (N_8781,N_1770,N_4792);
and U8782 (N_8782,N_3550,N_2534);
nor U8783 (N_8783,N_1078,N_4890);
nand U8784 (N_8784,N_1106,N_1696);
and U8785 (N_8785,N_4201,N_1151);
or U8786 (N_8786,N_3457,N_4241);
nor U8787 (N_8787,N_299,N_4349);
xor U8788 (N_8788,N_4360,N_2326);
nor U8789 (N_8789,N_2422,N_4755);
nor U8790 (N_8790,N_3652,N_2034);
nor U8791 (N_8791,N_2941,N_4845);
and U8792 (N_8792,N_1276,N_4655);
nand U8793 (N_8793,N_4119,N_1130);
nand U8794 (N_8794,N_4829,N_4612);
nor U8795 (N_8795,N_4208,N_47);
nor U8796 (N_8796,N_1228,N_419);
nand U8797 (N_8797,N_3186,N_29);
xnor U8798 (N_8798,N_143,N_319);
or U8799 (N_8799,N_862,N_541);
xor U8800 (N_8800,N_2760,N_2342);
or U8801 (N_8801,N_2731,N_3632);
nand U8802 (N_8802,N_4108,N_1889);
or U8803 (N_8803,N_314,N_998);
or U8804 (N_8804,N_757,N_3847);
and U8805 (N_8805,N_2283,N_1810);
or U8806 (N_8806,N_2269,N_35);
nand U8807 (N_8807,N_914,N_398);
nor U8808 (N_8808,N_4062,N_703);
nor U8809 (N_8809,N_3100,N_3914);
or U8810 (N_8810,N_1217,N_2581);
or U8811 (N_8811,N_4762,N_998);
or U8812 (N_8812,N_4845,N_2738);
or U8813 (N_8813,N_1344,N_798);
xnor U8814 (N_8814,N_1705,N_761);
nand U8815 (N_8815,N_2837,N_1395);
or U8816 (N_8816,N_1519,N_1743);
nor U8817 (N_8817,N_871,N_2836);
xnor U8818 (N_8818,N_1574,N_1253);
nor U8819 (N_8819,N_2090,N_1797);
nor U8820 (N_8820,N_3953,N_2769);
nand U8821 (N_8821,N_3240,N_3888);
nand U8822 (N_8822,N_4026,N_1463);
and U8823 (N_8823,N_1795,N_766);
nand U8824 (N_8824,N_2309,N_3680);
nand U8825 (N_8825,N_202,N_2340);
xnor U8826 (N_8826,N_2831,N_1411);
and U8827 (N_8827,N_1410,N_2964);
nor U8828 (N_8828,N_270,N_1270);
nand U8829 (N_8829,N_21,N_3253);
nand U8830 (N_8830,N_3625,N_561);
or U8831 (N_8831,N_3734,N_4084);
or U8832 (N_8832,N_2138,N_1461);
or U8833 (N_8833,N_1336,N_4048);
nor U8834 (N_8834,N_1079,N_3011);
xnor U8835 (N_8835,N_2183,N_2087);
and U8836 (N_8836,N_3852,N_3765);
or U8837 (N_8837,N_2320,N_3235);
and U8838 (N_8838,N_1915,N_3739);
nand U8839 (N_8839,N_575,N_4864);
or U8840 (N_8840,N_860,N_1579);
nand U8841 (N_8841,N_3276,N_3503);
or U8842 (N_8842,N_2312,N_4130);
nand U8843 (N_8843,N_1395,N_3218);
xnor U8844 (N_8844,N_1851,N_189);
nor U8845 (N_8845,N_3964,N_3901);
nor U8846 (N_8846,N_2641,N_2403);
nor U8847 (N_8847,N_2461,N_42);
or U8848 (N_8848,N_1948,N_1560);
xor U8849 (N_8849,N_4805,N_1001);
xnor U8850 (N_8850,N_4888,N_2864);
or U8851 (N_8851,N_1550,N_4785);
or U8852 (N_8852,N_1569,N_1557);
nand U8853 (N_8853,N_344,N_4921);
and U8854 (N_8854,N_4579,N_1427);
xnor U8855 (N_8855,N_3789,N_284);
or U8856 (N_8856,N_3245,N_3916);
nand U8857 (N_8857,N_4864,N_3483);
xor U8858 (N_8858,N_359,N_304);
xor U8859 (N_8859,N_4788,N_1808);
nand U8860 (N_8860,N_4522,N_1934);
xor U8861 (N_8861,N_3380,N_3785);
nand U8862 (N_8862,N_3399,N_3908);
nor U8863 (N_8863,N_3048,N_2076);
xnor U8864 (N_8864,N_2481,N_1356);
or U8865 (N_8865,N_2275,N_4686);
and U8866 (N_8866,N_2628,N_3300);
nor U8867 (N_8867,N_4131,N_4052);
nor U8868 (N_8868,N_695,N_702);
and U8869 (N_8869,N_961,N_3022);
nand U8870 (N_8870,N_1886,N_1524);
nand U8871 (N_8871,N_513,N_1588);
and U8872 (N_8872,N_4611,N_4742);
xor U8873 (N_8873,N_3888,N_1127);
or U8874 (N_8874,N_2610,N_2877);
nand U8875 (N_8875,N_2278,N_3288);
nor U8876 (N_8876,N_561,N_3478);
nand U8877 (N_8877,N_3291,N_2936);
and U8878 (N_8878,N_184,N_640);
and U8879 (N_8879,N_4908,N_3297);
or U8880 (N_8880,N_3248,N_718);
nand U8881 (N_8881,N_2314,N_3646);
and U8882 (N_8882,N_4338,N_4977);
and U8883 (N_8883,N_3619,N_4675);
xnor U8884 (N_8884,N_2351,N_1032);
nor U8885 (N_8885,N_878,N_3043);
nor U8886 (N_8886,N_3162,N_3858);
xnor U8887 (N_8887,N_2371,N_1269);
nor U8888 (N_8888,N_4236,N_2605);
or U8889 (N_8889,N_1254,N_4130);
xnor U8890 (N_8890,N_3257,N_4237);
nand U8891 (N_8891,N_4485,N_2064);
xnor U8892 (N_8892,N_2478,N_3781);
or U8893 (N_8893,N_3438,N_613);
xor U8894 (N_8894,N_4025,N_1870);
and U8895 (N_8895,N_4739,N_3648);
nand U8896 (N_8896,N_2962,N_942);
or U8897 (N_8897,N_947,N_1019);
nor U8898 (N_8898,N_1470,N_558);
nor U8899 (N_8899,N_1885,N_512);
or U8900 (N_8900,N_4951,N_376);
nor U8901 (N_8901,N_175,N_1728);
or U8902 (N_8902,N_2010,N_4206);
nand U8903 (N_8903,N_3333,N_4232);
nor U8904 (N_8904,N_1215,N_4307);
xnor U8905 (N_8905,N_1320,N_1454);
xor U8906 (N_8906,N_3260,N_223);
nor U8907 (N_8907,N_3644,N_690);
nor U8908 (N_8908,N_2952,N_2817);
nand U8909 (N_8909,N_4573,N_558);
and U8910 (N_8910,N_788,N_2313);
and U8911 (N_8911,N_995,N_1495);
and U8912 (N_8912,N_4926,N_2054);
xor U8913 (N_8913,N_916,N_3647);
xor U8914 (N_8914,N_2958,N_4818);
and U8915 (N_8915,N_2856,N_1597);
and U8916 (N_8916,N_4709,N_4922);
nand U8917 (N_8917,N_3335,N_3763);
nor U8918 (N_8918,N_1802,N_2504);
or U8919 (N_8919,N_3169,N_4664);
or U8920 (N_8920,N_1792,N_4419);
and U8921 (N_8921,N_4694,N_3990);
or U8922 (N_8922,N_4482,N_1258);
or U8923 (N_8923,N_3484,N_800);
nand U8924 (N_8924,N_3245,N_510);
xor U8925 (N_8925,N_1201,N_214);
nor U8926 (N_8926,N_657,N_814);
xor U8927 (N_8927,N_2846,N_3175);
and U8928 (N_8928,N_1479,N_221);
xor U8929 (N_8929,N_2226,N_4845);
nand U8930 (N_8930,N_278,N_4954);
xor U8931 (N_8931,N_78,N_675);
or U8932 (N_8932,N_27,N_2163);
nor U8933 (N_8933,N_4164,N_309);
and U8934 (N_8934,N_1846,N_723);
or U8935 (N_8935,N_4650,N_3523);
and U8936 (N_8936,N_2376,N_1472);
nor U8937 (N_8937,N_3902,N_3761);
nor U8938 (N_8938,N_2922,N_3259);
or U8939 (N_8939,N_3746,N_2594);
and U8940 (N_8940,N_360,N_4229);
and U8941 (N_8941,N_1227,N_2754);
and U8942 (N_8942,N_1437,N_1937);
xnor U8943 (N_8943,N_2562,N_1);
nand U8944 (N_8944,N_2532,N_3278);
or U8945 (N_8945,N_223,N_2513);
and U8946 (N_8946,N_3639,N_123);
nand U8947 (N_8947,N_4231,N_1887);
xor U8948 (N_8948,N_3801,N_1058);
nand U8949 (N_8949,N_2259,N_1283);
or U8950 (N_8950,N_4483,N_1185);
nor U8951 (N_8951,N_3496,N_3291);
or U8952 (N_8952,N_2676,N_3947);
nor U8953 (N_8953,N_1660,N_4099);
or U8954 (N_8954,N_881,N_2397);
xor U8955 (N_8955,N_2061,N_4630);
nand U8956 (N_8956,N_3130,N_1679);
nand U8957 (N_8957,N_1676,N_4256);
nand U8958 (N_8958,N_2588,N_2031);
and U8959 (N_8959,N_2780,N_713);
and U8960 (N_8960,N_1867,N_3097);
nand U8961 (N_8961,N_3722,N_3417);
xnor U8962 (N_8962,N_2633,N_1014);
or U8963 (N_8963,N_253,N_3795);
nor U8964 (N_8964,N_1483,N_4523);
nand U8965 (N_8965,N_3130,N_1291);
nor U8966 (N_8966,N_187,N_376);
or U8967 (N_8967,N_4331,N_4036);
xnor U8968 (N_8968,N_4001,N_1939);
nand U8969 (N_8969,N_1802,N_1506);
nor U8970 (N_8970,N_1828,N_2971);
nor U8971 (N_8971,N_2619,N_4928);
and U8972 (N_8972,N_1384,N_2998);
or U8973 (N_8973,N_4793,N_4461);
nor U8974 (N_8974,N_576,N_4023);
xor U8975 (N_8975,N_2467,N_169);
xnor U8976 (N_8976,N_2414,N_4996);
xnor U8977 (N_8977,N_1807,N_583);
and U8978 (N_8978,N_528,N_4527);
nand U8979 (N_8979,N_2098,N_952);
or U8980 (N_8980,N_3359,N_3485);
nand U8981 (N_8981,N_2675,N_481);
nand U8982 (N_8982,N_532,N_119);
nand U8983 (N_8983,N_3524,N_4386);
and U8984 (N_8984,N_4159,N_418);
xnor U8985 (N_8985,N_1107,N_4283);
xnor U8986 (N_8986,N_2720,N_2286);
xor U8987 (N_8987,N_4408,N_443);
xnor U8988 (N_8988,N_259,N_2372);
nor U8989 (N_8989,N_4878,N_3378);
and U8990 (N_8990,N_2022,N_3098);
and U8991 (N_8991,N_3870,N_3214);
nor U8992 (N_8992,N_1817,N_116);
nand U8993 (N_8993,N_1137,N_4977);
nor U8994 (N_8994,N_1975,N_3509);
or U8995 (N_8995,N_2826,N_178);
and U8996 (N_8996,N_742,N_2164);
and U8997 (N_8997,N_4835,N_3339);
nor U8998 (N_8998,N_2363,N_1039);
nor U8999 (N_8999,N_661,N_4148);
and U9000 (N_9000,N_1521,N_2147);
and U9001 (N_9001,N_1011,N_3269);
or U9002 (N_9002,N_3517,N_3099);
nand U9003 (N_9003,N_4753,N_2901);
nor U9004 (N_9004,N_4754,N_684);
nand U9005 (N_9005,N_1129,N_2799);
xnor U9006 (N_9006,N_4464,N_3210);
and U9007 (N_9007,N_1721,N_1419);
nor U9008 (N_9008,N_3727,N_2559);
or U9009 (N_9009,N_2197,N_4176);
or U9010 (N_9010,N_1059,N_4645);
nand U9011 (N_9011,N_3449,N_319);
nor U9012 (N_9012,N_1909,N_4045);
nand U9013 (N_9013,N_1748,N_1925);
or U9014 (N_9014,N_3541,N_1231);
nor U9015 (N_9015,N_3809,N_10);
and U9016 (N_9016,N_1916,N_2106);
nand U9017 (N_9017,N_3723,N_883);
xor U9018 (N_9018,N_4787,N_579);
xor U9019 (N_9019,N_2378,N_3606);
xnor U9020 (N_9020,N_3711,N_3967);
and U9021 (N_9021,N_329,N_2906);
nor U9022 (N_9022,N_4387,N_4672);
xnor U9023 (N_9023,N_1698,N_1975);
or U9024 (N_9024,N_4911,N_370);
and U9025 (N_9025,N_16,N_2213);
or U9026 (N_9026,N_2868,N_4835);
xnor U9027 (N_9027,N_3806,N_2021);
nand U9028 (N_9028,N_4670,N_2308);
or U9029 (N_9029,N_1262,N_4598);
nand U9030 (N_9030,N_3565,N_2362);
xor U9031 (N_9031,N_2255,N_701);
xnor U9032 (N_9032,N_3062,N_1578);
xor U9033 (N_9033,N_4195,N_560);
nand U9034 (N_9034,N_3861,N_2261);
nor U9035 (N_9035,N_4365,N_1702);
nor U9036 (N_9036,N_869,N_456);
and U9037 (N_9037,N_1129,N_1101);
xor U9038 (N_9038,N_765,N_3137);
or U9039 (N_9039,N_1319,N_3585);
nand U9040 (N_9040,N_3062,N_2095);
or U9041 (N_9041,N_1128,N_2707);
xnor U9042 (N_9042,N_1459,N_4770);
nor U9043 (N_9043,N_4510,N_63);
and U9044 (N_9044,N_3696,N_430);
xor U9045 (N_9045,N_4338,N_1249);
nor U9046 (N_9046,N_4898,N_2544);
nor U9047 (N_9047,N_4196,N_1775);
xor U9048 (N_9048,N_2231,N_4063);
and U9049 (N_9049,N_2938,N_2665);
and U9050 (N_9050,N_4229,N_4629);
nand U9051 (N_9051,N_2350,N_2926);
nand U9052 (N_9052,N_3222,N_649);
and U9053 (N_9053,N_1267,N_3351);
nor U9054 (N_9054,N_2031,N_4294);
nor U9055 (N_9055,N_893,N_4189);
xor U9056 (N_9056,N_44,N_682);
nand U9057 (N_9057,N_3074,N_2641);
nand U9058 (N_9058,N_2954,N_3431);
or U9059 (N_9059,N_173,N_725);
and U9060 (N_9060,N_1855,N_2513);
nor U9061 (N_9061,N_4094,N_826);
nor U9062 (N_9062,N_3224,N_1312);
nand U9063 (N_9063,N_2157,N_1402);
xor U9064 (N_9064,N_3201,N_451);
xnor U9065 (N_9065,N_1921,N_2255);
and U9066 (N_9066,N_2277,N_100);
xor U9067 (N_9067,N_3132,N_3783);
and U9068 (N_9068,N_2692,N_3626);
or U9069 (N_9069,N_3342,N_1882);
xnor U9070 (N_9070,N_221,N_949);
nor U9071 (N_9071,N_1329,N_553);
and U9072 (N_9072,N_956,N_2486);
xor U9073 (N_9073,N_4408,N_1691);
nand U9074 (N_9074,N_4477,N_4297);
and U9075 (N_9075,N_1306,N_4653);
and U9076 (N_9076,N_4733,N_3389);
and U9077 (N_9077,N_1332,N_156);
xor U9078 (N_9078,N_1936,N_775);
or U9079 (N_9079,N_2296,N_4601);
and U9080 (N_9080,N_187,N_4062);
xor U9081 (N_9081,N_1063,N_3303);
nand U9082 (N_9082,N_1822,N_3964);
nand U9083 (N_9083,N_3332,N_1457);
xnor U9084 (N_9084,N_2866,N_4080);
nand U9085 (N_9085,N_3983,N_1501);
nor U9086 (N_9086,N_3761,N_2674);
and U9087 (N_9087,N_648,N_1791);
or U9088 (N_9088,N_440,N_3392);
nor U9089 (N_9089,N_2343,N_4282);
and U9090 (N_9090,N_3853,N_2931);
nand U9091 (N_9091,N_4018,N_2480);
nand U9092 (N_9092,N_671,N_1583);
or U9093 (N_9093,N_2938,N_1104);
nor U9094 (N_9094,N_4039,N_1496);
nand U9095 (N_9095,N_2607,N_52);
xor U9096 (N_9096,N_4197,N_282);
nor U9097 (N_9097,N_2409,N_488);
nor U9098 (N_9098,N_2278,N_4533);
and U9099 (N_9099,N_2893,N_1883);
xnor U9100 (N_9100,N_1518,N_927);
or U9101 (N_9101,N_4000,N_3080);
xnor U9102 (N_9102,N_3103,N_4004);
nand U9103 (N_9103,N_4381,N_535);
nor U9104 (N_9104,N_3289,N_3841);
and U9105 (N_9105,N_2160,N_3403);
xor U9106 (N_9106,N_511,N_835);
nor U9107 (N_9107,N_3620,N_94);
nand U9108 (N_9108,N_2253,N_1725);
xor U9109 (N_9109,N_1533,N_4485);
or U9110 (N_9110,N_2590,N_1434);
or U9111 (N_9111,N_1067,N_26);
nor U9112 (N_9112,N_1495,N_1576);
nor U9113 (N_9113,N_678,N_4085);
xor U9114 (N_9114,N_145,N_4047);
and U9115 (N_9115,N_1861,N_4640);
and U9116 (N_9116,N_110,N_45);
nand U9117 (N_9117,N_113,N_3238);
nor U9118 (N_9118,N_2443,N_4995);
or U9119 (N_9119,N_2089,N_4335);
nand U9120 (N_9120,N_3222,N_3175);
nand U9121 (N_9121,N_1484,N_1657);
or U9122 (N_9122,N_1639,N_4683);
or U9123 (N_9123,N_4439,N_2527);
xnor U9124 (N_9124,N_4744,N_1121);
or U9125 (N_9125,N_563,N_4660);
and U9126 (N_9126,N_2242,N_2998);
nor U9127 (N_9127,N_3492,N_2294);
or U9128 (N_9128,N_996,N_3635);
xnor U9129 (N_9129,N_1977,N_404);
and U9130 (N_9130,N_3469,N_2420);
and U9131 (N_9131,N_1759,N_3154);
xor U9132 (N_9132,N_498,N_1604);
nor U9133 (N_9133,N_4515,N_985);
or U9134 (N_9134,N_1478,N_4457);
or U9135 (N_9135,N_1331,N_941);
nor U9136 (N_9136,N_3645,N_2938);
or U9137 (N_9137,N_4470,N_2866);
nor U9138 (N_9138,N_2331,N_180);
nand U9139 (N_9139,N_1903,N_2230);
xor U9140 (N_9140,N_3972,N_4183);
xor U9141 (N_9141,N_4092,N_4488);
xor U9142 (N_9142,N_2899,N_2715);
or U9143 (N_9143,N_13,N_1586);
nand U9144 (N_9144,N_425,N_3337);
nand U9145 (N_9145,N_846,N_1099);
xor U9146 (N_9146,N_2628,N_4789);
or U9147 (N_9147,N_3846,N_4594);
and U9148 (N_9148,N_2469,N_881);
nand U9149 (N_9149,N_3537,N_4412);
and U9150 (N_9150,N_1153,N_2104);
or U9151 (N_9151,N_1583,N_3325);
nand U9152 (N_9152,N_1899,N_4759);
nand U9153 (N_9153,N_3672,N_1064);
and U9154 (N_9154,N_4752,N_918);
and U9155 (N_9155,N_2243,N_1840);
nand U9156 (N_9156,N_2752,N_224);
nand U9157 (N_9157,N_4533,N_1956);
nor U9158 (N_9158,N_2212,N_178);
and U9159 (N_9159,N_1835,N_551);
xor U9160 (N_9160,N_2627,N_1452);
xnor U9161 (N_9161,N_1723,N_2182);
xor U9162 (N_9162,N_3815,N_4735);
nor U9163 (N_9163,N_2156,N_516);
nor U9164 (N_9164,N_944,N_2360);
nor U9165 (N_9165,N_4265,N_4222);
and U9166 (N_9166,N_4686,N_1013);
xnor U9167 (N_9167,N_1292,N_2057);
nor U9168 (N_9168,N_1493,N_2948);
or U9169 (N_9169,N_2422,N_471);
nor U9170 (N_9170,N_3807,N_255);
xnor U9171 (N_9171,N_3447,N_1078);
nand U9172 (N_9172,N_1221,N_3574);
or U9173 (N_9173,N_4601,N_4559);
or U9174 (N_9174,N_3413,N_4661);
nand U9175 (N_9175,N_3837,N_3072);
and U9176 (N_9176,N_1011,N_4164);
and U9177 (N_9177,N_3151,N_1252);
nor U9178 (N_9178,N_2366,N_695);
and U9179 (N_9179,N_4875,N_1261);
or U9180 (N_9180,N_3828,N_666);
or U9181 (N_9181,N_4229,N_2125);
or U9182 (N_9182,N_3758,N_1810);
nand U9183 (N_9183,N_3908,N_3603);
and U9184 (N_9184,N_2302,N_3648);
nor U9185 (N_9185,N_1594,N_3347);
nor U9186 (N_9186,N_2860,N_529);
and U9187 (N_9187,N_312,N_567);
and U9188 (N_9188,N_1006,N_490);
and U9189 (N_9189,N_367,N_2564);
and U9190 (N_9190,N_2084,N_3899);
nand U9191 (N_9191,N_4042,N_4689);
and U9192 (N_9192,N_410,N_4623);
nor U9193 (N_9193,N_1015,N_3707);
nor U9194 (N_9194,N_3394,N_1759);
and U9195 (N_9195,N_3746,N_4864);
nand U9196 (N_9196,N_3594,N_586);
and U9197 (N_9197,N_4836,N_1175);
nor U9198 (N_9198,N_3450,N_286);
nor U9199 (N_9199,N_2724,N_2740);
xnor U9200 (N_9200,N_377,N_2347);
and U9201 (N_9201,N_1042,N_928);
or U9202 (N_9202,N_3809,N_667);
xor U9203 (N_9203,N_365,N_805);
nor U9204 (N_9204,N_2242,N_4942);
nand U9205 (N_9205,N_3582,N_1843);
nand U9206 (N_9206,N_1397,N_304);
nand U9207 (N_9207,N_1895,N_3809);
xor U9208 (N_9208,N_1565,N_4963);
nand U9209 (N_9209,N_4290,N_4820);
and U9210 (N_9210,N_3491,N_3367);
xnor U9211 (N_9211,N_1820,N_3403);
xor U9212 (N_9212,N_3856,N_945);
nand U9213 (N_9213,N_2453,N_2382);
and U9214 (N_9214,N_3486,N_2409);
nand U9215 (N_9215,N_2704,N_2265);
or U9216 (N_9216,N_2601,N_242);
xor U9217 (N_9217,N_2188,N_3335);
and U9218 (N_9218,N_1260,N_1145);
nand U9219 (N_9219,N_2471,N_2219);
and U9220 (N_9220,N_3304,N_296);
nor U9221 (N_9221,N_4386,N_1079);
nor U9222 (N_9222,N_1544,N_4308);
or U9223 (N_9223,N_1227,N_608);
and U9224 (N_9224,N_1650,N_215);
nor U9225 (N_9225,N_4550,N_4067);
nand U9226 (N_9226,N_4371,N_1083);
nor U9227 (N_9227,N_2237,N_3555);
and U9228 (N_9228,N_76,N_2608);
or U9229 (N_9229,N_3100,N_3691);
nand U9230 (N_9230,N_30,N_4113);
nor U9231 (N_9231,N_1210,N_4982);
nand U9232 (N_9232,N_1304,N_3524);
xnor U9233 (N_9233,N_4512,N_4644);
xor U9234 (N_9234,N_4198,N_4601);
or U9235 (N_9235,N_2813,N_3533);
nor U9236 (N_9236,N_927,N_4685);
xnor U9237 (N_9237,N_135,N_3926);
nand U9238 (N_9238,N_1687,N_3590);
nand U9239 (N_9239,N_4760,N_3933);
nor U9240 (N_9240,N_1930,N_32);
and U9241 (N_9241,N_294,N_4145);
xor U9242 (N_9242,N_3181,N_870);
nor U9243 (N_9243,N_513,N_2630);
and U9244 (N_9244,N_316,N_3370);
xnor U9245 (N_9245,N_3221,N_2463);
xnor U9246 (N_9246,N_1976,N_2847);
and U9247 (N_9247,N_1210,N_4940);
or U9248 (N_9248,N_3849,N_1276);
or U9249 (N_9249,N_2793,N_3118);
xor U9250 (N_9250,N_4007,N_4462);
nand U9251 (N_9251,N_1461,N_963);
or U9252 (N_9252,N_4859,N_4023);
xor U9253 (N_9253,N_1975,N_4125);
and U9254 (N_9254,N_2727,N_3768);
and U9255 (N_9255,N_3427,N_230);
xor U9256 (N_9256,N_2706,N_2799);
xnor U9257 (N_9257,N_3885,N_520);
xor U9258 (N_9258,N_4147,N_2074);
xor U9259 (N_9259,N_4094,N_1070);
and U9260 (N_9260,N_0,N_4861);
xnor U9261 (N_9261,N_3461,N_4336);
or U9262 (N_9262,N_1686,N_2689);
nor U9263 (N_9263,N_2498,N_3019);
xor U9264 (N_9264,N_4035,N_1293);
and U9265 (N_9265,N_4942,N_502);
xnor U9266 (N_9266,N_714,N_4143);
or U9267 (N_9267,N_4273,N_3901);
xnor U9268 (N_9268,N_3696,N_3582);
nor U9269 (N_9269,N_449,N_1377);
xnor U9270 (N_9270,N_4379,N_1930);
nand U9271 (N_9271,N_2870,N_4529);
nor U9272 (N_9272,N_4700,N_4144);
nand U9273 (N_9273,N_4063,N_635);
or U9274 (N_9274,N_96,N_2084);
or U9275 (N_9275,N_1940,N_3992);
xnor U9276 (N_9276,N_1250,N_2869);
xnor U9277 (N_9277,N_3993,N_1926);
nand U9278 (N_9278,N_1812,N_4974);
or U9279 (N_9279,N_3762,N_2692);
xnor U9280 (N_9280,N_150,N_3196);
or U9281 (N_9281,N_4940,N_2055);
nor U9282 (N_9282,N_1881,N_4528);
nand U9283 (N_9283,N_731,N_4816);
and U9284 (N_9284,N_2011,N_2321);
xor U9285 (N_9285,N_2174,N_3015);
xnor U9286 (N_9286,N_612,N_4665);
nand U9287 (N_9287,N_2210,N_2829);
xor U9288 (N_9288,N_1151,N_4017);
or U9289 (N_9289,N_4987,N_4628);
nand U9290 (N_9290,N_1253,N_3327);
or U9291 (N_9291,N_1301,N_86);
and U9292 (N_9292,N_1631,N_1795);
or U9293 (N_9293,N_2701,N_720);
nor U9294 (N_9294,N_1191,N_957);
xnor U9295 (N_9295,N_4422,N_1201);
or U9296 (N_9296,N_2553,N_4940);
or U9297 (N_9297,N_629,N_3269);
nand U9298 (N_9298,N_3160,N_404);
and U9299 (N_9299,N_348,N_4425);
nand U9300 (N_9300,N_411,N_3844);
nand U9301 (N_9301,N_403,N_2702);
nor U9302 (N_9302,N_3714,N_840);
nand U9303 (N_9303,N_4187,N_418);
nand U9304 (N_9304,N_1198,N_4995);
and U9305 (N_9305,N_1136,N_4866);
or U9306 (N_9306,N_360,N_870);
or U9307 (N_9307,N_548,N_4150);
xnor U9308 (N_9308,N_1731,N_3185);
xor U9309 (N_9309,N_1857,N_4950);
and U9310 (N_9310,N_4113,N_3110);
xnor U9311 (N_9311,N_4684,N_364);
or U9312 (N_9312,N_2275,N_32);
or U9313 (N_9313,N_1195,N_485);
nor U9314 (N_9314,N_143,N_3493);
nor U9315 (N_9315,N_2036,N_431);
or U9316 (N_9316,N_419,N_1818);
nor U9317 (N_9317,N_3897,N_2499);
xor U9318 (N_9318,N_3564,N_3887);
nor U9319 (N_9319,N_688,N_1478);
or U9320 (N_9320,N_1675,N_1608);
and U9321 (N_9321,N_3145,N_1970);
or U9322 (N_9322,N_149,N_3875);
and U9323 (N_9323,N_388,N_2430);
nor U9324 (N_9324,N_3138,N_1290);
xor U9325 (N_9325,N_4616,N_4019);
and U9326 (N_9326,N_2289,N_4115);
or U9327 (N_9327,N_4832,N_3741);
xor U9328 (N_9328,N_4165,N_1528);
nor U9329 (N_9329,N_1303,N_4631);
or U9330 (N_9330,N_4819,N_3550);
xnor U9331 (N_9331,N_4227,N_1003);
nor U9332 (N_9332,N_4914,N_3627);
xnor U9333 (N_9333,N_2712,N_1813);
and U9334 (N_9334,N_3737,N_2039);
or U9335 (N_9335,N_1521,N_3257);
or U9336 (N_9336,N_2576,N_1087);
nor U9337 (N_9337,N_4424,N_96);
xnor U9338 (N_9338,N_4298,N_4708);
nand U9339 (N_9339,N_879,N_1499);
nor U9340 (N_9340,N_798,N_1414);
and U9341 (N_9341,N_2796,N_1100);
xnor U9342 (N_9342,N_3128,N_247);
nor U9343 (N_9343,N_3761,N_4072);
nor U9344 (N_9344,N_1992,N_3802);
or U9345 (N_9345,N_4805,N_421);
nand U9346 (N_9346,N_1970,N_2195);
and U9347 (N_9347,N_1068,N_4267);
nor U9348 (N_9348,N_3882,N_2401);
and U9349 (N_9349,N_2951,N_2050);
xor U9350 (N_9350,N_2154,N_27);
and U9351 (N_9351,N_4594,N_1658);
nand U9352 (N_9352,N_4492,N_3355);
and U9353 (N_9353,N_3190,N_1482);
or U9354 (N_9354,N_591,N_3525);
or U9355 (N_9355,N_0,N_2018);
nor U9356 (N_9356,N_1730,N_4658);
nand U9357 (N_9357,N_4358,N_4575);
or U9358 (N_9358,N_1563,N_1371);
xor U9359 (N_9359,N_107,N_3489);
and U9360 (N_9360,N_2072,N_563);
nor U9361 (N_9361,N_3061,N_1935);
and U9362 (N_9362,N_3046,N_4313);
nor U9363 (N_9363,N_3580,N_2149);
nand U9364 (N_9364,N_3949,N_1885);
xnor U9365 (N_9365,N_2908,N_3612);
nand U9366 (N_9366,N_4875,N_3008);
nor U9367 (N_9367,N_1303,N_293);
nand U9368 (N_9368,N_3095,N_4105);
nor U9369 (N_9369,N_1632,N_4930);
or U9370 (N_9370,N_2922,N_564);
nor U9371 (N_9371,N_616,N_3796);
and U9372 (N_9372,N_252,N_3819);
nor U9373 (N_9373,N_4037,N_894);
and U9374 (N_9374,N_2896,N_3913);
and U9375 (N_9375,N_1024,N_4692);
nor U9376 (N_9376,N_2667,N_4468);
or U9377 (N_9377,N_2028,N_4925);
and U9378 (N_9378,N_709,N_831);
nand U9379 (N_9379,N_2772,N_3439);
xnor U9380 (N_9380,N_3987,N_78);
or U9381 (N_9381,N_4440,N_206);
and U9382 (N_9382,N_1159,N_4446);
and U9383 (N_9383,N_3027,N_4650);
and U9384 (N_9384,N_1735,N_4850);
or U9385 (N_9385,N_4817,N_2958);
and U9386 (N_9386,N_4096,N_4523);
xnor U9387 (N_9387,N_3261,N_2137);
nor U9388 (N_9388,N_656,N_1337);
and U9389 (N_9389,N_1419,N_4558);
and U9390 (N_9390,N_540,N_2948);
or U9391 (N_9391,N_2847,N_3467);
or U9392 (N_9392,N_1148,N_409);
nor U9393 (N_9393,N_1051,N_3344);
xor U9394 (N_9394,N_2905,N_3321);
xnor U9395 (N_9395,N_832,N_3473);
xor U9396 (N_9396,N_547,N_3379);
nand U9397 (N_9397,N_1876,N_1995);
or U9398 (N_9398,N_136,N_143);
or U9399 (N_9399,N_2013,N_3093);
or U9400 (N_9400,N_575,N_4997);
xor U9401 (N_9401,N_2558,N_4814);
or U9402 (N_9402,N_1192,N_2427);
and U9403 (N_9403,N_2538,N_1784);
xnor U9404 (N_9404,N_4904,N_1351);
nor U9405 (N_9405,N_862,N_4411);
nor U9406 (N_9406,N_2565,N_750);
nor U9407 (N_9407,N_727,N_1250);
or U9408 (N_9408,N_553,N_598);
or U9409 (N_9409,N_1206,N_3331);
nor U9410 (N_9410,N_4424,N_716);
or U9411 (N_9411,N_4498,N_2868);
and U9412 (N_9412,N_2330,N_3560);
nand U9413 (N_9413,N_2511,N_2299);
and U9414 (N_9414,N_1195,N_58);
and U9415 (N_9415,N_646,N_3470);
xnor U9416 (N_9416,N_3122,N_360);
and U9417 (N_9417,N_410,N_4920);
nand U9418 (N_9418,N_3472,N_3817);
nor U9419 (N_9419,N_4647,N_1215);
xor U9420 (N_9420,N_37,N_1127);
nand U9421 (N_9421,N_3025,N_627);
nor U9422 (N_9422,N_2771,N_1440);
or U9423 (N_9423,N_383,N_1466);
nor U9424 (N_9424,N_1655,N_1888);
xor U9425 (N_9425,N_1851,N_269);
and U9426 (N_9426,N_2009,N_1489);
nor U9427 (N_9427,N_4738,N_3517);
xor U9428 (N_9428,N_4373,N_4386);
nand U9429 (N_9429,N_805,N_3179);
nor U9430 (N_9430,N_3261,N_2432);
xor U9431 (N_9431,N_4707,N_1741);
and U9432 (N_9432,N_803,N_1084);
or U9433 (N_9433,N_2101,N_342);
or U9434 (N_9434,N_1621,N_1509);
xor U9435 (N_9435,N_1138,N_3110);
nor U9436 (N_9436,N_1083,N_2696);
xnor U9437 (N_9437,N_3339,N_3927);
xnor U9438 (N_9438,N_1437,N_444);
or U9439 (N_9439,N_0,N_2745);
and U9440 (N_9440,N_2491,N_2361);
xor U9441 (N_9441,N_551,N_2301);
xnor U9442 (N_9442,N_3327,N_4907);
nand U9443 (N_9443,N_923,N_78);
and U9444 (N_9444,N_2651,N_3888);
nand U9445 (N_9445,N_3371,N_1940);
nand U9446 (N_9446,N_4912,N_3804);
or U9447 (N_9447,N_4368,N_1378);
and U9448 (N_9448,N_2262,N_250);
nand U9449 (N_9449,N_3758,N_1911);
or U9450 (N_9450,N_3073,N_4479);
nand U9451 (N_9451,N_1039,N_3872);
or U9452 (N_9452,N_4039,N_3175);
or U9453 (N_9453,N_3934,N_4596);
nand U9454 (N_9454,N_2087,N_3695);
nor U9455 (N_9455,N_3437,N_3350);
and U9456 (N_9456,N_4451,N_4928);
nor U9457 (N_9457,N_3939,N_4616);
or U9458 (N_9458,N_4747,N_792);
xor U9459 (N_9459,N_4195,N_3642);
nor U9460 (N_9460,N_1645,N_146);
nand U9461 (N_9461,N_3306,N_2049);
or U9462 (N_9462,N_78,N_4770);
or U9463 (N_9463,N_1255,N_1196);
nor U9464 (N_9464,N_3168,N_2343);
nand U9465 (N_9465,N_2030,N_596);
or U9466 (N_9466,N_1811,N_1355);
xor U9467 (N_9467,N_3672,N_3941);
or U9468 (N_9468,N_3478,N_1324);
and U9469 (N_9469,N_1360,N_4532);
or U9470 (N_9470,N_2805,N_4948);
or U9471 (N_9471,N_2212,N_1481);
xnor U9472 (N_9472,N_1,N_709);
or U9473 (N_9473,N_1973,N_3240);
xnor U9474 (N_9474,N_786,N_3411);
nor U9475 (N_9475,N_4253,N_2582);
and U9476 (N_9476,N_1964,N_2519);
nor U9477 (N_9477,N_1231,N_1984);
xor U9478 (N_9478,N_3754,N_1700);
or U9479 (N_9479,N_4993,N_1656);
and U9480 (N_9480,N_2129,N_2714);
nand U9481 (N_9481,N_3597,N_2606);
or U9482 (N_9482,N_4350,N_3770);
and U9483 (N_9483,N_743,N_1872);
and U9484 (N_9484,N_3930,N_2417);
and U9485 (N_9485,N_2894,N_1252);
or U9486 (N_9486,N_2999,N_3088);
xor U9487 (N_9487,N_1816,N_2539);
nor U9488 (N_9488,N_4489,N_2455);
nor U9489 (N_9489,N_3368,N_1246);
and U9490 (N_9490,N_2681,N_1850);
nor U9491 (N_9491,N_1647,N_2233);
nand U9492 (N_9492,N_4639,N_2684);
nor U9493 (N_9493,N_617,N_483);
nand U9494 (N_9494,N_1171,N_2807);
and U9495 (N_9495,N_3768,N_176);
nand U9496 (N_9496,N_916,N_1643);
and U9497 (N_9497,N_3766,N_1562);
nand U9498 (N_9498,N_4382,N_684);
and U9499 (N_9499,N_3842,N_1660);
nand U9500 (N_9500,N_646,N_2747);
and U9501 (N_9501,N_2583,N_3902);
nor U9502 (N_9502,N_194,N_1557);
xor U9503 (N_9503,N_4006,N_2509);
nand U9504 (N_9504,N_2299,N_4133);
xor U9505 (N_9505,N_530,N_195);
or U9506 (N_9506,N_4094,N_4490);
or U9507 (N_9507,N_1364,N_2408);
xor U9508 (N_9508,N_3280,N_3136);
or U9509 (N_9509,N_3283,N_1845);
or U9510 (N_9510,N_2983,N_2608);
nand U9511 (N_9511,N_1444,N_678);
and U9512 (N_9512,N_628,N_1774);
xnor U9513 (N_9513,N_921,N_2679);
nor U9514 (N_9514,N_3810,N_720);
nor U9515 (N_9515,N_874,N_3928);
or U9516 (N_9516,N_3046,N_3767);
nor U9517 (N_9517,N_3088,N_1249);
nand U9518 (N_9518,N_230,N_3828);
or U9519 (N_9519,N_1680,N_4708);
or U9520 (N_9520,N_1898,N_2461);
and U9521 (N_9521,N_2609,N_2902);
xor U9522 (N_9522,N_2152,N_3753);
nor U9523 (N_9523,N_3977,N_4323);
xnor U9524 (N_9524,N_4393,N_4972);
nand U9525 (N_9525,N_3506,N_1292);
xnor U9526 (N_9526,N_482,N_3158);
nor U9527 (N_9527,N_4865,N_2621);
or U9528 (N_9528,N_1647,N_2966);
xor U9529 (N_9529,N_4926,N_1827);
nand U9530 (N_9530,N_294,N_1229);
and U9531 (N_9531,N_2948,N_516);
or U9532 (N_9532,N_683,N_3501);
xnor U9533 (N_9533,N_3255,N_2926);
nand U9534 (N_9534,N_3927,N_2467);
or U9535 (N_9535,N_4358,N_2230);
nor U9536 (N_9536,N_3103,N_1586);
xor U9537 (N_9537,N_1611,N_2474);
nor U9538 (N_9538,N_4924,N_4484);
nand U9539 (N_9539,N_2299,N_2827);
and U9540 (N_9540,N_4269,N_1108);
or U9541 (N_9541,N_861,N_176);
or U9542 (N_9542,N_4616,N_1034);
or U9543 (N_9543,N_2723,N_2807);
and U9544 (N_9544,N_4739,N_2412);
nor U9545 (N_9545,N_4083,N_3876);
or U9546 (N_9546,N_4253,N_2005);
nand U9547 (N_9547,N_4804,N_3509);
nor U9548 (N_9548,N_260,N_2901);
nor U9549 (N_9549,N_1988,N_2848);
and U9550 (N_9550,N_4826,N_1273);
and U9551 (N_9551,N_4334,N_4656);
xor U9552 (N_9552,N_1602,N_899);
nor U9553 (N_9553,N_1035,N_3348);
xor U9554 (N_9554,N_3464,N_4740);
and U9555 (N_9555,N_4459,N_2355);
xor U9556 (N_9556,N_494,N_2608);
nand U9557 (N_9557,N_2861,N_50);
xor U9558 (N_9558,N_3754,N_155);
or U9559 (N_9559,N_2014,N_539);
nor U9560 (N_9560,N_3942,N_133);
or U9561 (N_9561,N_2882,N_2962);
nand U9562 (N_9562,N_768,N_3753);
nand U9563 (N_9563,N_4000,N_2715);
nor U9564 (N_9564,N_467,N_1725);
and U9565 (N_9565,N_2544,N_4875);
nor U9566 (N_9566,N_1460,N_4939);
xor U9567 (N_9567,N_1168,N_1994);
nand U9568 (N_9568,N_2988,N_3058);
or U9569 (N_9569,N_3574,N_2849);
nor U9570 (N_9570,N_2734,N_1902);
and U9571 (N_9571,N_3264,N_129);
or U9572 (N_9572,N_2441,N_369);
nor U9573 (N_9573,N_2213,N_1528);
nand U9574 (N_9574,N_2305,N_2341);
and U9575 (N_9575,N_1327,N_3352);
or U9576 (N_9576,N_4634,N_1073);
nand U9577 (N_9577,N_3888,N_4608);
nand U9578 (N_9578,N_2613,N_3461);
nor U9579 (N_9579,N_3563,N_2332);
xnor U9580 (N_9580,N_2616,N_2055);
or U9581 (N_9581,N_3379,N_4734);
xor U9582 (N_9582,N_2418,N_3775);
xnor U9583 (N_9583,N_804,N_2480);
or U9584 (N_9584,N_3859,N_1129);
nand U9585 (N_9585,N_36,N_1400);
nor U9586 (N_9586,N_4662,N_3455);
nor U9587 (N_9587,N_1127,N_847);
nand U9588 (N_9588,N_591,N_2808);
nor U9589 (N_9589,N_3744,N_980);
nor U9590 (N_9590,N_3027,N_3433);
and U9591 (N_9591,N_4060,N_109);
or U9592 (N_9592,N_2386,N_2029);
and U9593 (N_9593,N_4117,N_2502);
nand U9594 (N_9594,N_2264,N_1512);
or U9595 (N_9595,N_4672,N_3211);
nor U9596 (N_9596,N_1104,N_4332);
nor U9597 (N_9597,N_2394,N_4350);
nor U9598 (N_9598,N_757,N_4808);
and U9599 (N_9599,N_3203,N_3442);
xor U9600 (N_9600,N_4245,N_2317);
xor U9601 (N_9601,N_1691,N_1367);
and U9602 (N_9602,N_3369,N_1585);
and U9603 (N_9603,N_2456,N_2028);
xnor U9604 (N_9604,N_2922,N_682);
nand U9605 (N_9605,N_2975,N_1299);
nand U9606 (N_9606,N_2340,N_4093);
nor U9607 (N_9607,N_3602,N_1365);
nand U9608 (N_9608,N_2480,N_2789);
nand U9609 (N_9609,N_4522,N_4427);
nor U9610 (N_9610,N_1105,N_2107);
nor U9611 (N_9611,N_1150,N_435);
or U9612 (N_9612,N_2549,N_3052);
or U9613 (N_9613,N_2072,N_1989);
xnor U9614 (N_9614,N_4451,N_2215);
and U9615 (N_9615,N_22,N_1602);
or U9616 (N_9616,N_2973,N_4135);
nand U9617 (N_9617,N_541,N_1474);
nand U9618 (N_9618,N_1105,N_3454);
nand U9619 (N_9619,N_1896,N_1656);
xnor U9620 (N_9620,N_3650,N_2308);
or U9621 (N_9621,N_1732,N_3413);
or U9622 (N_9622,N_3492,N_4387);
xor U9623 (N_9623,N_2377,N_1062);
and U9624 (N_9624,N_4358,N_3559);
nand U9625 (N_9625,N_321,N_3563);
or U9626 (N_9626,N_479,N_3235);
nand U9627 (N_9627,N_514,N_4699);
xor U9628 (N_9628,N_4049,N_4772);
nand U9629 (N_9629,N_3056,N_2849);
nor U9630 (N_9630,N_80,N_4049);
nor U9631 (N_9631,N_1815,N_2749);
nor U9632 (N_9632,N_158,N_356);
nor U9633 (N_9633,N_869,N_1835);
or U9634 (N_9634,N_3197,N_390);
or U9635 (N_9635,N_3533,N_3079);
and U9636 (N_9636,N_3463,N_4950);
nor U9637 (N_9637,N_2836,N_2405);
nand U9638 (N_9638,N_2677,N_4915);
and U9639 (N_9639,N_1901,N_3255);
nor U9640 (N_9640,N_4270,N_3531);
nand U9641 (N_9641,N_1095,N_3346);
xnor U9642 (N_9642,N_2560,N_4189);
and U9643 (N_9643,N_2502,N_717);
nand U9644 (N_9644,N_2555,N_4416);
and U9645 (N_9645,N_4277,N_3036);
and U9646 (N_9646,N_1827,N_2122);
xor U9647 (N_9647,N_4323,N_915);
xor U9648 (N_9648,N_4370,N_207);
nand U9649 (N_9649,N_2457,N_1831);
nor U9650 (N_9650,N_500,N_3822);
xor U9651 (N_9651,N_1732,N_2739);
or U9652 (N_9652,N_3559,N_2632);
nor U9653 (N_9653,N_3509,N_4861);
nor U9654 (N_9654,N_4796,N_1643);
and U9655 (N_9655,N_2068,N_1900);
nor U9656 (N_9656,N_4208,N_34);
xor U9657 (N_9657,N_1184,N_3906);
nand U9658 (N_9658,N_2721,N_1935);
nor U9659 (N_9659,N_670,N_3321);
xnor U9660 (N_9660,N_529,N_2353);
nor U9661 (N_9661,N_944,N_244);
xor U9662 (N_9662,N_2011,N_1629);
or U9663 (N_9663,N_598,N_4070);
xor U9664 (N_9664,N_4421,N_3325);
nand U9665 (N_9665,N_1691,N_3761);
nand U9666 (N_9666,N_3921,N_3814);
nor U9667 (N_9667,N_3737,N_359);
xnor U9668 (N_9668,N_1074,N_1445);
and U9669 (N_9669,N_1719,N_2762);
nand U9670 (N_9670,N_3145,N_1360);
or U9671 (N_9671,N_1011,N_4492);
nand U9672 (N_9672,N_4299,N_4274);
or U9673 (N_9673,N_2677,N_359);
or U9674 (N_9674,N_1290,N_2544);
xnor U9675 (N_9675,N_604,N_1025);
xor U9676 (N_9676,N_1078,N_1420);
nor U9677 (N_9677,N_154,N_3892);
nor U9678 (N_9678,N_1503,N_2661);
nand U9679 (N_9679,N_4475,N_3657);
nand U9680 (N_9680,N_854,N_4692);
xnor U9681 (N_9681,N_4141,N_2790);
nand U9682 (N_9682,N_1641,N_322);
nand U9683 (N_9683,N_2170,N_1240);
nor U9684 (N_9684,N_3106,N_2053);
or U9685 (N_9685,N_885,N_3883);
nand U9686 (N_9686,N_4968,N_1811);
and U9687 (N_9687,N_3201,N_1052);
xnor U9688 (N_9688,N_2560,N_2477);
and U9689 (N_9689,N_2315,N_2955);
nor U9690 (N_9690,N_507,N_2498);
and U9691 (N_9691,N_1373,N_560);
nor U9692 (N_9692,N_623,N_3528);
nor U9693 (N_9693,N_2494,N_3135);
xor U9694 (N_9694,N_3753,N_65);
and U9695 (N_9695,N_1531,N_1213);
nor U9696 (N_9696,N_4696,N_1317);
or U9697 (N_9697,N_3830,N_4587);
xnor U9698 (N_9698,N_3571,N_378);
and U9699 (N_9699,N_4111,N_2823);
or U9700 (N_9700,N_3838,N_689);
nand U9701 (N_9701,N_2967,N_975);
nand U9702 (N_9702,N_1204,N_3634);
nand U9703 (N_9703,N_4795,N_3326);
nor U9704 (N_9704,N_498,N_216);
xor U9705 (N_9705,N_2479,N_2569);
and U9706 (N_9706,N_3736,N_4424);
nor U9707 (N_9707,N_185,N_3318);
and U9708 (N_9708,N_1278,N_3151);
xor U9709 (N_9709,N_2267,N_4454);
or U9710 (N_9710,N_88,N_4825);
nor U9711 (N_9711,N_246,N_3885);
nor U9712 (N_9712,N_1590,N_1879);
xor U9713 (N_9713,N_4783,N_94);
xor U9714 (N_9714,N_1354,N_3605);
and U9715 (N_9715,N_398,N_53);
xor U9716 (N_9716,N_815,N_3134);
or U9717 (N_9717,N_3276,N_1994);
or U9718 (N_9718,N_4581,N_3723);
and U9719 (N_9719,N_2924,N_3888);
xnor U9720 (N_9720,N_2663,N_4312);
xnor U9721 (N_9721,N_2185,N_1411);
and U9722 (N_9722,N_248,N_4266);
xnor U9723 (N_9723,N_4195,N_3953);
nor U9724 (N_9724,N_3624,N_289);
nand U9725 (N_9725,N_365,N_4895);
xnor U9726 (N_9726,N_3594,N_2371);
and U9727 (N_9727,N_2735,N_91);
nor U9728 (N_9728,N_3813,N_1897);
nand U9729 (N_9729,N_4176,N_1308);
xnor U9730 (N_9730,N_1106,N_1490);
xnor U9731 (N_9731,N_2248,N_1914);
nand U9732 (N_9732,N_4849,N_194);
and U9733 (N_9733,N_1451,N_3061);
or U9734 (N_9734,N_1476,N_4566);
xor U9735 (N_9735,N_3013,N_2088);
nand U9736 (N_9736,N_2080,N_1127);
xor U9737 (N_9737,N_3479,N_549);
nand U9738 (N_9738,N_694,N_2113);
nor U9739 (N_9739,N_1967,N_853);
and U9740 (N_9740,N_1569,N_1647);
nor U9741 (N_9741,N_1021,N_2769);
nand U9742 (N_9742,N_318,N_1258);
xnor U9743 (N_9743,N_897,N_3160);
and U9744 (N_9744,N_1831,N_4644);
nand U9745 (N_9745,N_2490,N_4510);
xnor U9746 (N_9746,N_3846,N_3748);
and U9747 (N_9747,N_4286,N_2607);
or U9748 (N_9748,N_237,N_4007);
nand U9749 (N_9749,N_232,N_4880);
and U9750 (N_9750,N_677,N_1700);
or U9751 (N_9751,N_2984,N_97);
xor U9752 (N_9752,N_2038,N_3802);
and U9753 (N_9753,N_3546,N_1985);
nor U9754 (N_9754,N_3248,N_4272);
or U9755 (N_9755,N_1565,N_4876);
or U9756 (N_9756,N_2484,N_3110);
nor U9757 (N_9757,N_4658,N_2296);
and U9758 (N_9758,N_617,N_2897);
nand U9759 (N_9759,N_2086,N_9);
and U9760 (N_9760,N_3893,N_2204);
nand U9761 (N_9761,N_2626,N_3239);
or U9762 (N_9762,N_2752,N_1876);
nand U9763 (N_9763,N_4193,N_1635);
nor U9764 (N_9764,N_3843,N_87);
nand U9765 (N_9765,N_1616,N_1904);
or U9766 (N_9766,N_2693,N_2670);
or U9767 (N_9767,N_3853,N_1904);
nor U9768 (N_9768,N_1248,N_4607);
xnor U9769 (N_9769,N_4288,N_307);
xnor U9770 (N_9770,N_3891,N_353);
and U9771 (N_9771,N_1764,N_2072);
and U9772 (N_9772,N_2995,N_2494);
and U9773 (N_9773,N_1496,N_3272);
or U9774 (N_9774,N_3643,N_3009);
xnor U9775 (N_9775,N_3624,N_3230);
xnor U9776 (N_9776,N_4698,N_4714);
nor U9777 (N_9777,N_2365,N_720);
xor U9778 (N_9778,N_4383,N_1267);
and U9779 (N_9779,N_1886,N_2711);
or U9780 (N_9780,N_1611,N_2187);
xor U9781 (N_9781,N_1710,N_151);
xor U9782 (N_9782,N_2619,N_2951);
xnor U9783 (N_9783,N_1623,N_633);
nor U9784 (N_9784,N_1650,N_4573);
xor U9785 (N_9785,N_4575,N_3990);
and U9786 (N_9786,N_1111,N_1507);
and U9787 (N_9787,N_357,N_1704);
and U9788 (N_9788,N_3161,N_486);
and U9789 (N_9789,N_4913,N_1138);
nor U9790 (N_9790,N_162,N_4346);
nor U9791 (N_9791,N_3031,N_1240);
nor U9792 (N_9792,N_3426,N_2418);
or U9793 (N_9793,N_4135,N_1734);
or U9794 (N_9794,N_883,N_4110);
xor U9795 (N_9795,N_2405,N_3516);
or U9796 (N_9796,N_1072,N_3355);
nor U9797 (N_9797,N_3357,N_2944);
or U9798 (N_9798,N_2607,N_3946);
and U9799 (N_9799,N_441,N_3369);
and U9800 (N_9800,N_3886,N_1766);
and U9801 (N_9801,N_3740,N_4031);
nand U9802 (N_9802,N_4662,N_823);
or U9803 (N_9803,N_2899,N_3185);
nor U9804 (N_9804,N_4617,N_2614);
or U9805 (N_9805,N_455,N_1828);
nor U9806 (N_9806,N_873,N_4047);
xor U9807 (N_9807,N_4460,N_4004);
and U9808 (N_9808,N_4582,N_1499);
nor U9809 (N_9809,N_4909,N_2143);
nand U9810 (N_9810,N_2893,N_1793);
nor U9811 (N_9811,N_1628,N_152);
xnor U9812 (N_9812,N_4533,N_1556);
nand U9813 (N_9813,N_933,N_4271);
nand U9814 (N_9814,N_793,N_1845);
xnor U9815 (N_9815,N_4069,N_325);
or U9816 (N_9816,N_3651,N_362);
and U9817 (N_9817,N_29,N_2104);
nor U9818 (N_9818,N_4527,N_3863);
nand U9819 (N_9819,N_24,N_3026);
nor U9820 (N_9820,N_2762,N_4559);
nand U9821 (N_9821,N_4637,N_3271);
xor U9822 (N_9822,N_3146,N_1438);
nor U9823 (N_9823,N_1166,N_1717);
nand U9824 (N_9824,N_2635,N_3347);
xnor U9825 (N_9825,N_732,N_986);
or U9826 (N_9826,N_4509,N_2553);
xnor U9827 (N_9827,N_1143,N_3490);
nor U9828 (N_9828,N_997,N_3858);
nand U9829 (N_9829,N_401,N_991);
nor U9830 (N_9830,N_633,N_4637);
and U9831 (N_9831,N_3812,N_2774);
xor U9832 (N_9832,N_4572,N_3383);
nand U9833 (N_9833,N_2363,N_4161);
and U9834 (N_9834,N_705,N_1032);
and U9835 (N_9835,N_4752,N_3829);
and U9836 (N_9836,N_2950,N_469);
xor U9837 (N_9837,N_2862,N_1702);
nor U9838 (N_9838,N_3382,N_3259);
nand U9839 (N_9839,N_923,N_1923);
nor U9840 (N_9840,N_2468,N_3070);
nor U9841 (N_9841,N_4225,N_1682);
and U9842 (N_9842,N_2688,N_3960);
nand U9843 (N_9843,N_1247,N_3947);
nor U9844 (N_9844,N_4121,N_3555);
nor U9845 (N_9845,N_3812,N_3287);
or U9846 (N_9846,N_2169,N_2665);
nand U9847 (N_9847,N_3112,N_1807);
xor U9848 (N_9848,N_3602,N_1994);
or U9849 (N_9849,N_3007,N_488);
and U9850 (N_9850,N_1983,N_2579);
or U9851 (N_9851,N_415,N_3810);
nor U9852 (N_9852,N_670,N_2217);
and U9853 (N_9853,N_3296,N_3126);
or U9854 (N_9854,N_3961,N_4963);
nor U9855 (N_9855,N_2643,N_2003);
nor U9856 (N_9856,N_2440,N_4320);
nand U9857 (N_9857,N_4356,N_3990);
or U9858 (N_9858,N_1207,N_2142);
nor U9859 (N_9859,N_3795,N_3200);
nand U9860 (N_9860,N_4833,N_171);
and U9861 (N_9861,N_4022,N_216);
nand U9862 (N_9862,N_4597,N_3409);
xor U9863 (N_9863,N_1946,N_2806);
and U9864 (N_9864,N_1574,N_1437);
nand U9865 (N_9865,N_3159,N_3832);
and U9866 (N_9866,N_898,N_757);
xor U9867 (N_9867,N_222,N_2351);
nor U9868 (N_9868,N_3432,N_1232);
nor U9869 (N_9869,N_577,N_420);
or U9870 (N_9870,N_4464,N_3310);
and U9871 (N_9871,N_4674,N_593);
xor U9872 (N_9872,N_4157,N_4269);
or U9873 (N_9873,N_2246,N_1311);
nor U9874 (N_9874,N_1515,N_1213);
or U9875 (N_9875,N_2011,N_3524);
and U9876 (N_9876,N_1493,N_272);
nor U9877 (N_9877,N_458,N_1226);
nand U9878 (N_9878,N_267,N_3168);
nor U9879 (N_9879,N_2511,N_2810);
or U9880 (N_9880,N_3557,N_2092);
or U9881 (N_9881,N_3011,N_1056);
nand U9882 (N_9882,N_4261,N_4975);
and U9883 (N_9883,N_2849,N_4680);
nand U9884 (N_9884,N_3655,N_1153);
nor U9885 (N_9885,N_3797,N_3196);
and U9886 (N_9886,N_3903,N_4444);
or U9887 (N_9887,N_4739,N_1991);
xnor U9888 (N_9888,N_2669,N_4679);
and U9889 (N_9889,N_4249,N_3396);
nand U9890 (N_9890,N_28,N_2929);
or U9891 (N_9891,N_2633,N_1974);
or U9892 (N_9892,N_1159,N_3130);
xnor U9893 (N_9893,N_4074,N_2946);
and U9894 (N_9894,N_311,N_29);
nand U9895 (N_9895,N_390,N_4532);
xnor U9896 (N_9896,N_606,N_3826);
xnor U9897 (N_9897,N_760,N_4756);
nand U9898 (N_9898,N_3683,N_22);
nor U9899 (N_9899,N_1588,N_2599);
or U9900 (N_9900,N_1125,N_4956);
or U9901 (N_9901,N_3895,N_965);
xnor U9902 (N_9902,N_2220,N_4608);
xnor U9903 (N_9903,N_2306,N_1952);
nor U9904 (N_9904,N_4138,N_3612);
or U9905 (N_9905,N_1866,N_675);
and U9906 (N_9906,N_4598,N_1357);
xnor U9907 (N_9907,N_151,N_2907);
or U9908 (N_9908,N_4011,N_175);
and U9909 (N_9909,N_3414,N_2914);
nor U9910 (N_9910,N_4289,N_3806);
xnor U9911 (N_9911,N_3089,N_3169);
or U9912 (N_9912,N_4966,N_2647);
or U9913 (N_9913,N_4045,N_4049);
nor U9914 (N_9914,N_1388,N_3271);
nor U9915 (N_9915,N_3649,N_4227);
or U9916 (N_9916,N_4850,N_1111);
and U9917 (N_9917,N_339,N_3902);
nor U9918 (N_9918,N_2845,N_4080);
or U9919 (N_9919,N_1872,N_4061);
and U9920 (N_9920,N_4438,N_3883);
and U9921 (N_9921,N_4350,N_63);
nand U9922 (N_9922,N_4868,N_3765);
nand U9923 (N_9923,N_3817,N_1885);
and U9924 (N_9924,N_3858,N_1876);
xor U9925 (N_9925,N_1356,N_4590);
nor U9926 (N_9926,N_3089,N_596);
xnor U9927 (N_9927,N_4405,N_4223);
xor U9928 (N_9928,N_3257,N_4284);
nand U9929 (N_9929,N_3622,N_1628);
and U9930 (N_9930,N_365,N_3257);
or U9931 (N_9931,N_3142,N_3750);
and U9932 (N_9932,N_3980,N_4010);
and U9933 (N_9933,N_4818,N_3959);
nor U9934 (N_9934,N_12,N_2667);
nor U9935 (N_9935,N_1518,N_2323);
xnor U9936 (N_9936,N_1380,N_3152);
nand U9937 (N_9937,N_3920,N_1787);
nor U9938 (N_9938,N_3588,N_105);
nor U9939 (N_9939,N_1010,N_1648);
xnor U9940 (N_9940,N_284,N_1895);
or U9941 (N_9941,N_3459,N_3812);
or U9942 (N_9942,N_645,N_2431);
nand U9943 (N_9943,N_2920,N_1658);
xnor U9944 (N_9944,N_2649,N_4969);
or U9945 (N_9945,N_658,N_827);
xnor U9946 (N_9946,N_4211,N_2421);
or U9947 (N_9947,N_2664,N_4350);
xnor U9948 (N_9948,N_4254,N_4528);
or U9949 (N_9949,N_4468,N_4419);
or U9950 (N_9950,N_1544,N_873);
or U9951 (N_9951,N_2136,N_3230);
nand U9952 (N_9952,N_339,N_325);
nand U9953 (N_9953,N_1675,N_4188);
nor U9954 (N_9954,N_804,N_2399);
xor U9955 (N_9955,N_3266,N_896);
nor U9956 (N_9956,N_802,N_3781);
or U9957 (N_9957,N_4407,N_1630);
or U9958 (N_9958,N_2855,N_703);
xor U9959 (N_9959,N_3857,N_459);
nand U9960 (N_9960,N_344,N_4854);
nor U9961 (N_9961,N_4812,N_3152);
xor U9962 (N_9962,N_2607,N_3302);
nand U9963 (N_9963,N_1768,N_3695);
nand U9964 (N_9964,N_3578,N_2368);
or U9965 (N_9965,N_3129,N_4027);
nand U9966 (N_9966,N_2514,N_13);
xor U9967 (N_9967,N_2591,N_4535);
or U9968 (N_9968,N_2508,N_624);
nand U9969 (N_9969,N_3293,N_4058);
or U9970 (N_9970,N_47,N_2593);
nor U9971 (N_9971,N_1847,N_3698);
nor U9972 (N_9972,N_3743,N_3949);
nand U9973 (N_9973,N_3415,N_2165);
nand U9974 (N_9974,N_4036,N_4416);
and U9975 (N_9975,N_3984,N_1595);
and U9976 (N_9976,N_1299,N_1134);
and U9977 (N_9977,N_78,N_2533);
or U9978 (N_9978,N_4517,N_3071);
or U9979 (N_9979,N_3525,N_2676);
nand U9980 (N_9980,N_858,N_4939);
and U9981 (N_9981,N_3837,N_4222);
and U9982 (N_9982,N_3085,N_4953);
nor U9983 (N_9983,N_4434,N_2606);
or U9984 (N_9984,N_3682,N_1599);
or U9985 (N_9985,N_2882,N_3849);
xor U9986 (N_9986,N_1594,N_2181);
xor U9987 (N_9987,N_300,N_1157);
or U9988 (N_9988,N_2786,N_4944);
or U9989 (N_9989,N_511,N_817);
or U9990 (N_9990,N_1263,N_4216);
nand U9991 (N_9991,N_3316,N_4295);
or U9992 (N_9992,N_2244,N_2214);
nor U9993 (N_9993,N_4440,N_809);
xnor U9994 (N_9994,N_341,N_2196);
nand U9995 (N_9995,N_2755,N_339);
nand U9996 (N_9996,N_387,N_2173);
nor U9997 (N_9997,N_959,N_3608);
nor U9998 (N_9998,N_3294,N_988);
nor U9999 (N_9999,N_2801,N_4099);
nand U10000 (N_10000,N_8007,N_9630);
and U10001 (N_10001,N_5112,N_9597);
or U10002 (N_10002,N_8287,N_6463);
nand U10003 (N_10003,N_5336,N_7866);
xnor U10004 (N_10004,N_8405,N_7974);
or U10005 (N_10005,N_7590,N_8646);
nor U10006 (N_10006,N_7718,N_5761);
and U10007 (N_10007,N_6156,N_9123);
xor U10008 (N_10008,N_9897,N_7448);
nand U10009 (N_10009,N_8443,N_6360);
nor U10010 (N_10010,N_8300,N_6694);
xor U10011 (N_10011,N_8195,N_8347);
nand U10012 (N_10012,N_5174,N_5927);
nand U10013 (N_10013,N_7848,N_8217);
xnor U10014 (N_10014,N_9726,N_9909);
nand U10015 (N_10015,N_6622,N_6413);
or U10016 (N_10016,N_7834,N_5260);
xnor U10017 (N_10017,N_6551,N_5732);
nor U10018 (N_10018,N_7336,N_6461);
nand U10019 (N_10019,N_5291,N_7628);
nand U10020 (N_10020,N_7792,N_9942);
nor U10021 (N_10021,N_9814,N_5102);
nor U10022 (N_10022,N_9698,N_8201);
and U10023 (N_10023,N_7459,N_5481);
or U10024 (N_10024,N_5455,N_7329);
nand U10025 (N_10025,N_6897,N_9448);
or U10026 (N_10026,N_5380,N_6083);
nor U10027 (N_10027,N_5974,N_9585);
and U10028 (N_10028,N_8298,N_6733);
xor U10029 (N_10029,N_9756,N_5579);
nor U10030 (N_10030,N_7774,N_5632);
and U10031 (N_10031,N_6692,N_6742);
nor U10032 (N_10032,N_8952,N_9104);
nand U10033 (N_10033,N_5762,N_9154);
nor U10034 (N_10034,N_6944,N_5372);
or U10035 (N_10035,N_6184,N_9482);
nor U10036 (N_10036,N_8586,N_5705);
nor U10037 (N_10037,N_5898,N_9424);
and U10038 (N_10038,N_9758,N_6255);
nand U10039 (N_10039,N_9034,N_9927);
or U10040 (N_10040,N_6614,N_9061);
xor U10041 (N_10041,N_7141,N_7367);
nand U10042 (N_10042,N_7407,N_6318);
nor U10043 (N_10043,N_8553,N_6066);
or U10044 (N_10044,N_6535,N_5883);
nor U10045 (N_10045,N_6510,N_6289);
xor U10046 (N_10046,N_8481,N_9628);
or U10047 (N_10047,N_8808,N_5331);
xor U10048 (N_10048,N_8103,N_7871);
xnor U10049 (N_10049,N_8041,N_8827);
nand U10050 (N_10050,N_7476,N_9576);
nand U10051 (N_10051,N_9369,N_8514);
xnor U10052 (N_10052,N_5896,N_5303);
nand U10053 (N_10053,N_5866,N_7536);
nor U10054 (N_10054,N_6023,N_5595);
nor U10055 (N_10055,N_5129,N_8259);
and U10056 (N_10056,N_5633,N_5700);
nor U10057 (N_10057,N_9105,N_7402);
nor U10058 (N_10058,N_9910,N_7472);
nand U10059 (N_10059,N_7607,N_7066);
or U10060 (N_10060,N_5939,N_5061);
nor U10061 (N_10061,N_6630,N_9871);
and U10062 (N_10062,N_9640,N_8834);
nand U10063 (N_10063,N_8728,N_5493);
nor U10064 (N_10064,N_9226,N_7417);
nor U10065 (N_10065,N_6405,N_7559);
xnor U10066 (N_10066,N_8297,N_5111);
nor U10067 (N_10067,N_9944,N_8317);
xnor U10068 (N_10068,N_6383,N_8224);
nor U10069 (N_10069,N_9146,N_9738);
and U10070 (N_10070,N_6652,N_8561);
and U10071 (N_10071,N_6557,N_8526);
and U10072 (N_10072,N_8320,N_8450);
xor U10073 (N_10073,N_6749,N_6239);
nand U10074 (N_10074,N_5876,N_6588);
and U10075 (N_10075,N_7350,N_5279);
nand U10076 (N_10076,N_7038,N_5989);
xor U10077 (N_10077,N_7878,N_5919);
xor U10078 (N_10078,N_7556,N_6853);
nand U10079 (N_10079,N_6201,N_8638);
nor U10080 (N_10080,N_6218,N_6381);
xor U10081 (N_10081,N_9094,N_9418);
nor U10082 (N_10082,N_6299,N_8498);
and U10083 (N_10083,N_9109,N_7839);
xor U10084 (N_10084,N_7549,N_8092);
xor U10085 (N_10085,N_7130,N_7209);
or U10086 (N_10086,N_8322,N_9978);
or U10087 (N_10087,N_7493,N_9402);
or U10088 (N_10088,N_7423,N_9000);
nor U10089 (N_10089,N_8971,N_9318);
nor U10090 (N_10090,N_9158,N_5056);
nand U10091 (N_10091,N_9908,N_7680);
nor U10092 (N_10092,N_8896,N_8651);
and U10093 (N_10093,N_5949,N_8376);
nand U10094 (N_10094,N_9500,N_5987);
xnor U10095 (N_10095,N_7255,N_9149);
xor U10096 (N_10096,N_7847,N_7505);
nand U10097 (N_10097,N_6740,N_8953);
or U10098 (N_10098,N_7643,N_7452);
or U10099 (N_10099,N_9566,N_9579);
and U10100 (N_10100,N_7751,N_5826);
and U10101 (N_10101,N_6569,N_8951);
nand U10102 (N_10102,N_5857,N_8875);
nand U10103 (N_10103,N_6667,N_5489);
or U10104 (N_10104,N_6582,N_7431);
nand U10105 (N_10105,N_8886,N_8229);
xor U10106 (N_10106,N_8934,N_8010);
nor U10107 (N_10107,N_7308,N_6488);
or U10108 (N_10108,N_5284,N_5580);
and U10109 (N_10109,N_8147,N_7397);
nor U10110 (N_10110,N_8344,N_8199);
nor U10111 (N_10111,N_9413,N_6252);
xor U10112 (N_10112,N_7434,N_7158);
or U10113 (N_10113,N_6665,N_9567);
and U10114 (N_10114,N_5037,N_6715);
nand U10115 (N_10115,N_5335,N_5620);
xnor U10116 (N_10116,N_7796,N_5418);
nand U10117 (N_10117,N_9687,N_8282);
or U10118 (N_10118,N_5415,N_9182);
or U10119 (N_10119,N_7435,N_8751);
xor U10120 (N_10120,N_6000,N_9702);
xnor U10121 (N_10121,N_7801,N_8254);
or U10122 (N_10122,N_7770,N_6094);
xor U10123 (N_10123,N_5769,N_5009);
and U10124 (N_10124,N_6314,N_8962);
or U10125 (N_10125,N_9065,N_6202);
xnor U10126 (N_10126,N_6397,N_8558);
or U10127 (N_10127,N_5301,N_9936);
nor U10128 (N_10128,N_7877,N_7953);
nor U10129 (N_10129,N_9600,N_5094);
or U10130 (N_10130,N_5679,N_6936);
nand U10131 (N_10131,N_6596,N_6489);
or U10132 (N_10132,N_8079,N_7069);
nand U10133 (N_10133,N_9636,N_8505);
xor U10134 (N_10134,N_9218,N_5756);
or U10135 (N_10135,N_9537,N_5789);
nand U10136 (N_10136,N_7843,N_9818);
nor U10137 (N_10137,N_8266,N_7639);
nand U10138 (N_10138,N_7070,N_8303);
or U10139 (N_10139,N_9298,N_7723);
or U10140 (N_10140,N_6450,N_5315);
xnor U10141 (N_10141,N_9101,N_7132);
xnor U10142 (N_10142,N_6955,N_5109);
and U10143 (N_10143,N_6620,N_5381);
or U10144 (N_10144,N_6279,N_9623);
and U10145 (N_10145,N_5844,N_9442);
and U10146 (N_10146,N_6357,N_9121);
xor U10147 (N_10147,N_5449,N_9080);
or U10148 (N_10148,N_6361,N_9715);
or U10149 (N_10149,N_5736,N_5652);
nand U10150 (N_10150,N_6788,N_8197);
nor U10151 (N_10151,N_7778,N_9385);
nand U10152 (N_10152,N_6544,N_5773);
or U10153 (N_10153,N_5412,N_9992);
nand U10154 (N_10154,N_8495,N_6517);
and U10155 (N_10155,N_5634,N_6610);
nor U10156 (N_10156,N_6015,N_9898);
nand U10157 (N_10157,N_8114,N_5970);
xor U10158 (N_10158,N_5688,N_6248);
nand U10159 (N_10159,N_5858,N_5923);
or U10160 (N_10160,N_7880,N_5521);
and U10161 (N_10161,N_7173,N_7183);
and U10162 (N_10162,N_9139,N_5106);
or U10163 (N_10163,N_8527,N_6925);
xor U10164 (N_10164,N_8701,N_5695);
nor U10165 (N_10165,N_8679,N_5822);
nand U10166 (N_10166,N_8365,N_6457);
or U10167 (N_10167,N_8599,N_8183);
or U10168 (N_10168,N_6194,N_9042);
or U10169 (N_10169,N_6265,N_7623);
nor U10170 (N_10170,N_5911,N_7065);
and U10171 (N_10171,N_9358,N_8950);
xnor U10172 (N_10172,N_8148,N_7159);
nor U10173 (N_10173,N_6815,N_5630);
nand U10174 (N_10174,N_5388,N_5264);
xnor U10175 (N_10175,N_7300,N_7273);
xnor U10176 (N_10176,N_9841,N_7685);
nor U10177 (N_10177,N_5956,N_6057);
xor U10178 (N_10178,N_7389,N_5206);
xnor U10179 (N_10179,N_6053,N_5892);
xnor U10180 (N_10180,N_5780,N_6945);
and U10181 (N_10181,N_7468,N_8329);
nor U10182 (N_10182,N_7553,N_5877);
nor U10183 (N_10183,N_5431,N_6560);
nand U10184 (N_10184,N_7433,N_9221);
xor U10185 (N_10185,N_9453,N_9115);
and U10186 (N_10186,N_5364,N_5282);
or U10187 (N_10187,N_9980,N_7842);
and U10188 (N_10188,N_6783,N_6055);
nand U10189 (N_10189,N_9647,N_7032);
nand U10190 (N_10190,N_6563,N_8138);
or U10191 (N_10191,N_8268,N_8067);
and U10192 (N_10192,N_7694,N_8985);
xor U10193 (N_10193,N_7043,N_6542);
and U10194 (N_10194,N_8096,N_7802);
nor U10195 (N_10195,N_6567,N_7931);
or U10196 (N_10196,N_6878,N_5308);
or U10197 (N_10197,N_8131,N_8853);
nand U10198 (N_10198,N_7045,N_8018);
xor U10199 (N_10199,N_5066,N_6287);
and U10200 (N_10200,N_5712,N_6583);
nand U10201 (N_10201,N_8882,N_8885);
nand U10202 (N_10202,N_7289,N_7309);
or U10203 (N_10203,N_8351,N_9231);
or U10204 (N_10204,N_7487,N_5806);
or U10205 (N_10205,N_6346,N_7212);
or U10206 (N_10206,N_9704,N_5179);
xor U10207 (N_10207,N_5504,N_8039);
nand U10208 (N_10208,N_9331,N_8815);
nand U10209 (N_10209,N_6998,N_6837);
nor U10210 (N_10210,N_9663,N_8441);
and U10211 (N_10211,N_5880,N_8579);
nand U10212 (N_10212,N_8132,N_5398);
or U10213 (N_10213,N_8720,N_7907);
xor U10214 (N_10214,N_5680,N_5429);
xnor U10215 (N_10215,N_9799,N_9869);
or U10216 (N_10216,N_6136,N_6364);
nand U10217 (N_10217,N_8359,N_5678);
xor U10218 (N_10218,N_9718,N_7988);
and U10219 (N_10219,N_7884,N_6061);
nand U10220 (N_10220,N_5613,N_8639);
and U10221 (N_10221,N_7377,N_5104);
xnor U10222 (N_10222,N_9293,N_8105);
nor U10223 (N_10223,N_8629,N_7903);
nand U10224 (N_10224,N_9524,N_7742);
xor U10225 (N_10225,N_9510,N_5261);
nor U10226 (N_10226,N_7716,N_7291);
nand U10227 (N_10227,N_9862,N_6304);
nand U10228 (N_10228,N_5287,N_8472);
nor U10229 (N_10229,N_5859,N_6681);
nor U10230 (N_10230,N_9743,N_6787);
xor U10231 (N_10231,N_6391,N_9437);
or U10232 (N_10232,N_7322,N_7640);
or U10233 (N_10233,N_8683,N_9079);
or U10234 (N_10234,N_9404,N_9128);
xnor U10235 (N_10235,N_7138,N_7793);
nand U10236 (N_10236,N_9651,N_7337);
xnor U10237 (N_10237,N_9962,N_5224);
nand U10238 (N_10238,N_9100,N_6192);
and U10239 (N_10239,N_8657,N_7404);
nor U10240 (N_10240,N_6591,N_5592);
nor U10241 (N_10241,N_9465,N_6951);
xnor U10242 (N_10242,N_9801,N_9153);
nand U10243 (N_10243,N_8970,N_7485);
nor U10244 (N_10244,N_8642,N_5396);
nor U10245 (N_10245,N_9596,N_8417);
xnor U10246 (N_10246,N_8340,N_5399);
nand U10247 (N_10247,N_6024,N_5594);
xor U10248 (N_10248,N_6081,N_7196);
nor U10249 (N_10249,N_5997,N_8060);
xor U10250 (N_10250,N_5524,N_7677);
and U10251 (N_10251,N_8544,N_7438);
and U10252 (N_10252,N_6673,N_5186);
nand U10253 (N_10253,N_8880,N_8960);
and U10254 (N_10254,N_8273,N_6492);
or U10255 (N_10255,N_9710,N_6617);
nand U10256 (N_10256,N_9674,N_5792);
or U10257 (N_10257,N_8854,N_8125);
nor U10258 (N_10258,N_5363,N_8295);
and U10259 (N_10259,N_5092,N_9625);
nor U10260 (N_10260,N_9548,N_9706);
nor U10261 (N_10261,N_8097,N_9403);
or U10262 (N_10262,N_9430,N_6440);
nand U10263 (N_10263,N_7892,N_9682);
and U10264 (N_10264,N_8703,N_6608);
nor U10265 (N_10265,N_8852,N_8263);
nor U10266 (N_10266,N_7343,N_5059);
and U10267 (N_10267,N_5405,N_7693);
nand U10268 (N_10268,N_5435,N_6356);
or U10269 (N_10269,N_9297,N_6518);
nor U10270 (N_10270,N_6158,N_6827);
nand U10271 (N_10271,N_6281,N_5119);
and U10272 (N_10272,N_8164,N_7728);
or U10273 (N_10273,N_7018,N_5912);
or U10274 (N_10274,N_9302,N_6655);
and U10275 (N_10275,N_8725,N_6523);
nand U10276 (N_10276,N_9877,N_6179);
or U10277 (N_10277,N_8992,N_8850);
nand U10278 (N_10278,N_9744,N_8826);
nand U10279 (N_10279,N_7298,N_5465);
and U10280 (N_10280,N_6571,N_9638);
nand U10281 (N_10281,N_8784,N_5452);
xor U10282 (N_10282,N_6932,N_8972);
nor U10283 (N_10283,N_8672,N_5742);
nand U10284 (N_10284,N_9307,N_8063);
nand U10285 (N_10285,N_6394,N_8502);
or U10286 (N_10286,N_7027,N_6327);
and U10287 (N_10287,N_5306,N_9606);
xnor U10288 (N_10288,N_6266,N_8867);
xor U10289 (N_10289,N_9250,N_8400);
xnor U10290 (N_10290,N_8397,N_6999);
nand U10291 (N_10291,N_5842,N_7900);
nor U10292 (N_10292,N_8534,N_6033);
nor U10293 (N_10293,N_5181,N_8471);
xnor U10294 (N_10294,N_9283,N_8190);
nand U10295 (N_10295,N_5480,N_8941);
xnor U10296 (N_10296,N_5760,N_6819);
or U10297 (N_10297,N_6696,N_9435);
nor U10298 (N_10298,N_7233,N_8864);
xnor U10299 (N_10299,N_9714,N_7596);
xor U10300 (N_10300,N_8308,N_5784);
nand U10301 (N_10301,N_6766,N_8426);
nand U10302 (N_10302,N_7135,N_8621);
xor U10303 (N_10303,N_9243,N_7926);
nand U10304 (N_10304,N_9532,N_8496);
or U10305 (N_10305,N_7916,N_5525);
nor U10306 (N_10306,N_8754,N_6550);
nor U10307 (N_10307,N_9497,N_9048);
xor U10308 (N_10308,N_8899,N_5326);
or U10309 (N_10309,N_9050,N_6071);
and U10310 (N_10310,N_6721,N_9371);
xnor U10311 (N_10311,N_8723,N_6406);
and U10312 (N_10312,N_7840,N_5369);
xnor U10313 (N_10313,N_8588,N_6565);
nand U10314 (N_10314,N_9761,N_8036);
or U10315 (N_10315,N_6234,N_6553);
and U10316 (N_10316,N_7744,N_5038);
nand U10317 (N_10317,N_6091,N_6842);
xnor U10318 (N_10318,N_9905,N_6603);
or U10319 (N_10319,N_5627,N_7177);
xnor U10320 (N_10320,N_9914,N_5377);
nand U10321 (N_10321,N_7641,N_7029);
nand U10322 (N_10322,N_8492,N_8756);
and U10323 (N_10323,N_5341,N_9082);
xnor U10324 (N_10324,N_8153,N_5340);
and U10325 (N_10325,N_5672,N_9583);
or U10326 (N_10326,N_5016,N_9526);
xor U10327 (N_10327,N_6338,N_9560);
nand U10328 (N_10328,N_6166,N_7946);
xnor U10329 (N_10329,N_6931,N_7112);
or U10330 (N_10330,N_5740,N_7591);
or U10331 (N_10331,N_6683,N_7440);
xor U10332 (N_10332,N_8653,N_7126);
nor U10333 (N_10333,N_9310,N_9025);
nand U10334 (N_10334,N_7629,N_8069);
and U10335 (N_10335,N_8761,N_9794);
xor U10336 (N_10336,N_8293,N_9752);
xor U10337 (N_10337,N_6095,N_6367);
nor U10338 (N_10338,N_5086,N_8577);
nor U10339 (N_10339,N_8919,N_5026);
or U10340 (N_10340,N_7749,N_5755);
and U10341 (N_10341,N_6530,N_9261);
nand U10342 (N_10342,N_7063,N_7700);
xnor U10343 (N_10343,N_6212,N_6747);
nor U10344 (N_10344,N_9141,N_8944);
nand U10345 (N_10345,N_9843,N_8494);
or U10346 (N_10346,N_7672,N_6802);
or U10347 (N_10347,N_5607,N_5698);
and U10348 (N_10348,N_7058,N_7275);
or U10349 (N_10349,N_5660,N_9805);
xnor U10350 (N_10350,N_9290,N_6543);
nand U10351 (N_10351,N_5445,N_9299);
nor U10352 (N_10352,N_7481,N_8884);
xor U10353 (N_10353,N_7420,N_6839);
xor U10354 (N_10354,N_5664,N_5228);
and U10355 (N_10355,N_5983,N_8037);
nor U10356 (N_10356,N_9951,N_7030);
xor U10357 (N_10357,N_5601,N_6459);
nor U10358 (N_10358,N_5108,N_6816);
nor U10359 (N_10359,N_6691,N_9562);
or U10360 (N_10360,N_5915,N_8380);
and U10361 (N_10361,N_5235,N_5127);
xor U10362 (N_10362,N_6682,N_6240);
nor U10363 (N_10363,N_9728,N_7041);
xnor U10364 (N_10364,N_9975,N_7625);
nand U10365 (N_10365,N_5025,N_9938);
nand U10366 (N_10366,N_9713,N_5195);
or U10367 (N_10367,N_8830,N_6410);
xnor U10368 (N_10368,N_5558,N_7428);
nand U10369 (N_10369,N_8915,N_7996);
and U10370 (N_10370,N_7023,N_5598);
or U10371 (N_10371,N_8343,N_6908);
xor U10372 (N_10372,N_6592,N_8225);
nand U10373 (N_10373,N_7992,N_9495);
or U10374 (N_10374,N_6990,N_8978);
or U10375 (N_10375,N_9452,N_8996);
xnor U10376 (N_10376,N_5404,N_8401);
or U10377 (N_10377,N_6822,N_8666);
xnor U10378 (N_10378,N_9348,N_9570);
and U10379 (N_10379,N_7442,N_6589);
xnor U10380 (N_10380,N_8112,N_8810);
xor U10381 (N_10381,N_9601,N_6941);
nor U10382 (N_10382,N_5044,N_9166);
nand U10383 (N_10383,N_8011,N_6259);
xor U10384 (N_10384,N_7859,N_9943);
xnor U10385 (N_10385,N_9907,N_6835);
nand U10386 (N_10386,N_8937,N_8873);
nand U10387 (N_10387,N_5964,N_9396);
and U10388 (N_10388,N_7079,N_5669);
or U10389 (N_10389,N_8374,N_6199);
nand U10390 (N_10390,N_6409,N_6917);
xnor U10391 (N_10391,N_5426,N_8778);
xor U10392 (N_10392,N_7217,N_9895);
and U10393 (N_10393,N_8274,N_6757);
xor U10394 (N_10394,N_5014,N_6513);
or U10395 (N_10395,N_6145,N_7116);
xnor U10396 (N_10396,N_9904,N_9565);
or U10397 (N_10397,N_7581,N_8366);
or U10398 (N_10398,N_9444,N_9266);
nor U10399 (N_10399,N_5332,N_6422);
or U10400 (N_10400,N_5330,N_9813);
or U10401 (N_10401,N_6257,N_7583);
xor U10402 (N_10402,N_5374,N_6581);
xnor U10403 (N_10403,N_9828,N_9060);
nand U10404 (N_10404,N_5045,N_7824);
xor U10405 (N_10405,N_9865,N_7040);
and U10406 (N_10406,N_6408,N_6261);
nand U10407 (N_10407,N_6334,N_5820);
xnor U10408 (N_10408,N_7008,N_9339);
nand U10409 (N_10409,N_9125,N_7789);
or U10410 (N_10410,N_8319,N_6396);
or U10411 (N_10411,N_7817,N_5125);
nand U10412 (N_10412,N_7120,N_5670);
nor U10413 (N_10413,N_7514,N_7219);
nor U10414 (N_10414,N_6554,N_7664);
xor U10415 (N_10415,N_6800,N_9202);
xor U10416 (N_10416,N_5255,N_5123);
nor U10417 (N_10417,N_7649,N_7220);
or U10418 (N_10418,N_8444,N_6097);
nor U10419 (N_10419,N_5854,N_8969);
xor U10420 (N_10420,N_8154,N_8610);
nor U10421 (N_10421,N_5602,N_8708);
and U10422 (N_10422,N_7887,N_7797);
nor U10423 (N_10423,N_8115,N_8596);
xor U10424 (N_10424,N_7922,N_5548);
nand U10425 (N_10425,N_6432,N_7898);
or U10426 (N_10426,N_8608,N_6131);
nor U10427 (N_10427,N_6720,N_5873);
xor U10428 (N_10428,N_6549,N_9273);
xnor U10429 (N_10429,N_5031,N_9668);
nand U10430 (N_10430,N_8704,N_8332);
nor U10431 (N_10431,N_6995,N_8547);
nand U10432 (N_10432,N_7557,N_7633);
nor U10433 (N_10433,N_6627,N_5646);
nor U10434 (N_10434,N_6389,N_6796);
xnor U10435 (N_10435,N_8065,N_5370);
and U10436 (N_10436,N_5057,N_7371);
and U10437 (N_10437,N_6092,N_8580);
nor U10438 (N_10438,N_7737,N_6036);
and U10439 (N_10439,N_9083,N_8537);
nand U10440 (N_10440,N_9954,N_6585);
or U10441 (N_10441,N_6349,N_6121);
nor U10442 (N_10442,N_5074,N_5943);
or U10443 (N_10443,N_7381,N_6570);
or U10444 (N_10444,N_5673,N_9988);
or U10445 (N_10445,N_9120,N_5637);
and U10446 (N_10446,N_7053,N_8056);
or U10447 (N_10447,N_7624,N_9370);
and U10448 (N_10448,N_7686,N_5441);
xnor U10449 (N_10449,N_6102,N_9454);
nand U10450 (N_10450,N_7791,N_9447);
nor U10451 (N_10451,N_7967,N_6262);
and U10452 (N_10452,N_6431,N_5862);
xor U10453 (N_10453,N_8779,N_8803);
xor U10454 (N_10454,N_7998,N_6101);
and U10455 (N_10455,N_8981,N_8360);
nor U10456 (N_10456,N_5442,N_8030);
or U10457 (N_10457,N_5203,N_5611);
nor U10458 (N_10458,N_7709,N_9535);
nand U10459 (N_10459,N_8799,N_7940);
xor U10460 (N_10460,N_7021,N_8286);
or U10461 (N_10461,N_9229,N_7747);
nor U10462 (N_10462,N_9732,N_9882);
and U10463 (N_10463,N_5771,N_7787);
nand U10464 (N_10464,N_9263,N_9991);
xor U10465 (N_10465,N_7203,N_8304);
nand U10466 (N_10466,N_7644,N_6206);
nor U10467 (N_10467,N_7786,N_6484);
and U10468 (N_10468,N_8075,N_6512);
nand U10469 (N_10469,N_5468,N_5619);
and U10470 (N_10470,N_9705,N_5662);
xnor U10471 (N_10471,N_7010,N_7307);
nor U10472 (N_10472,N_9835,N_9508);
or U10473 (N_10473,N_6741,N_8513);
nand U10474 (N_10474,N_6045,N_9071);
nand U10475 (N_10475,N_5121,N_5804);
xor U10476 (N_10476,N_6111,N_8984);
or U10477 (N_10477,N_6601,N_5249);
and U10478 (N_10478,N_6828,N_6135);
xnor U10479 (N_10479,N_9451,N_7090);
nand U10480 (N_10480,N_5198,N_6548);
or U10481 (N_10481,N_9319,N_6105);
xnor U10482 (N_10482,N_6738,N_7568);
xor U10483 (N_10483,N_7175,N_7097);
and U10484 (N_10484,N_6729,N_9473);
nor U10485 (N_10485,N_8203,N_5077);
nor U10486 (N_10486,N_6298,N_6230);
and U10487 (N_10487,N_8175,N_6997);
nor U10488 (N_10488,N_7955,N_9730);
or U10489 (N_10489,N_5184,N_7531);
and U10490 (N_10490,N_8245,N_9832);
or U10491 (N_10491,N_8346,N_5827);
or U10492 (N_10492,N_8475,N_6452);
and U10493 (N_10493,N_6928,N_8363);
xor U10494 (N_10494,N_6967,N_8002);
and U10495 (N_10495,N_6175,N_6146);
xor U10496 (N_10496,N_9667,N_8939);
or U10497 (N_10497,N_7262,N_6223);
nand U10498 (N_10498,N_8729,N_6663);
or U10499 (N_10499,N_5200,N_5187);
nand U10500 (N_10500,N_7788,N_6233);
and U10501 (N_10501,N_9529,N_5350);
nor U10502 (N_10502,N_9772,N_9038);
nor U10503 (N_10503,N_8819,N_7124);
nor U10504 (N_10504,N_6744,N_7456);
nand U10505 (N_10505,N_5167,N_9431);
xnor U10506 (N_10506,N_5534,N_6286);
nand U10507 (N_10507,N_9327,N_8064);
nand U10508 (N_10508,N_5476,N_6502);
nor U10509 (N_10509,N_8959,N_7806);
xnor U10510 (N_10510,N_6495,N_8659);
nand U10511 (N_10511,N_9538,N_9249);
nor U10512 (N_10512,N_6678,N_6719);
nand U10513 (N_10513,N_8261,N_7000);
or U10514 (N_10514,N_6994,N_9866);
or U10515 (N_10515,N_9134,N_5810);
and U10516 (N_10516,N_9821,N_5356);
or U10517 (N_10517,N_9924,N_6467);
xnor U10518 (N_10518,N_8490,N_6244);
or U10519 (N_10519,N_8677,N_8240);
nand U10520 (N_10520,N_6618,N_9063);
or U10521 (N_10521,N_8872,N_5817);
xor U10522 (N_10522,N_7821,N_9851);
and U10523 (N_10523,N_5413,N_8179);
nand U10524 (N_10524,N_8349,N_9390);
xnor U10525 (N_10525,N_9819,N_9044);
nand U10526 (N_10526,N_7341,N_7147);
nand U10527 (N_10527,N_7885,N_7186);
and U10528 (N_10528,N_7102,N_9268);
nand U10529 (N_10529,N_9468,N_8822);
and U10530 (N_10530,N_6876,N_8160);
or U10531 (N_10531,N_6120,N_8795);
or U10532 (N_10532,N_7232,N_9365);
nor U10533 (N_10533,N_5265,N_5400);
nand U10534 (N_10534,N_5321,N_9414);
nand U10535 (N_10535,N_8008,N_5302);
nand U10536 (N_10536,N_9881,N_7195);
or U10537 (N_10537,N_6942,N_9615);
nand U10538 (N_10538,N_7961,N_6680);
nand U10539 (N_10539,N_9059,N_9655);
and U10540 (N_10540,N_5978,N_7836);
and U10541 (N_10541,N_9853,N_5828);
xor U10542 (N_10542,N_6311,N_6482);
xor U10543 (N_10543,N_8554,N_6813);
nor U10544 (N_10544,N_9353,N_5482);
nor U10545 (N_10545,N_8230,N_7332);
and U10546 (N_10546,N_9751,N_5644);
xnor U10547 (N_10547,N_5725,N_6671);
nor U10548 (N_10548,N_5948,N_5231);
xnor U10549 (N_10549,N_9621,N_7868);
xnor U10550 (N_10550,N_9325,N_8449);
and U10551 (N_10551,N_9543,N_5704);
nor U10552 (N_10552,N_9461,N_5357);
nand U10553 (N_10553,N_7704,N_9274);
xor U10554 (N_10554,N_8539,N_9490);
nand U10555 (N_10555,N_9703,N_5894);
nor U10556 (N_10556,N_6921,N_6737);
nand U10557 (N_10557,N_7987,N_9363);
and U10558 (N_10558,N_5596,N_9410);
nor U10559 (N_10559,N_5433,N_5342);
nand U10560 (N_10560,N_6520,N_9062);
nand U10561 (N_10561,N_7917,N_7263);
and U10562 (N_10562,N_7890,N_9934);
and U10563 (N_10563,N_6390,N_5779);
nor U10564 (N_10564,N_6593,N_6035);
or U10565 (N_10565,N_7106,N_8587);
nand U10566 (N_10566,N_6301,N_5499);
or U10567 (N_10567,N_5006,N_6605);
and U10568 (N_10568,N_7565,N_9419);
nand U10569 (N_10569,N_7560,N_9264);
nand U10570 (N_10570,N_7412,N_8152);
nor U10571 (N_10571,N_8042,N_8718);
or U10572 (N_10572,N_9998,N_9170);
xnor U10573 (N_10573,N_7034,N_9206);
nor U10574 (N_10574,N_8180,N_6752);
and U10575 (N_10575,N_6575,N_5367);
nand U10576 (N_10576,N_5214,N_6874);
nand U10577 (N_10577,N_9550,N_5355);
or U10578 (N_10578,N_8965,N_5737);
and U10579 (N_10579,N_8536,N_5313);
or U10580 (N_10580,N_5391,N_5692);
and U10581 (N_10581,N_8221,N_6190);
and U10582 (N_10582,N_7271,N_6370);
xor U10583 (N_10583,N_6873,N_7148);
or U10584 (N_10584,N_8606,N_7594);
or U10585 (N_10585,N_6499,N_9280);
nor U10586 (N_10586,N_7139,N_9970);
and U10587 (N_10587,N_7702,N_7668);
nor U10588 (N_10588,N_7290,N_8948);
or U10589 (N_10589,N_7429,N_7078);
nor U10590 (N_10590,N_5469,N_7608);
or U10591 (N_10591,N_6507,N_6910);
or U10592 (N_10592,N_8877,N_8540);
and U10593 (N_10593,N_7969,N_8173);
or U10594 (N_10594,N_9247,N_8545);
xnor U10595 (N_10595,N_6780,N_5141);
nor U10596 (N_10596,N_5414,N_9275);
xnor U10597 (N_10597,N_5194,N_5776);
and U10598 (N_10598,N_5176,N_9496);
nand U10599 (N_10599,N_6082,N_6188);
nand U10600 (N_10600,N_5132,N_9441);
nand U10601 (N_10601,N_5243,N_7011);
nand U10602 (N_10602,N_9748,N_9412);
nand U10603 (N_10603,N_7925,N_5572);
nor U10604 (N_10604,N_6666,N_7327);
or U10605 (N_10605,N_7865,N_5432);
nand U10606 (N_10606,N_5115,N_9069);
xnor U10607 (N_10607,N_8191,N_9831);
and U10608 (N_10608,N_7886,N_8993);
and U10609 (N_10609,N_5329,N_9676);
or U10610 (N_10610,N_6423,N_6730);
or U10611 (N_10611,N_5236,N_9278);
nand U10612 (N_10612,N_6833,N_6155);
or U10613 (N_10613,N_7837,N_6306);
or U10614 (N_10614,N_8936,N_8597);
and U10615 (N_10615,N_6472,N_8395);
or U10616 (N_10616,N_7086,N_8480);
nand U10617 (N_10617,N_7768,N_8082);
or U10618 (N_10618,N_6251,N_5182);
nor U10619 (N_10619,N_8829,N_7912);
or U10620 (N_10620,N_9028,N_7602);
and U10621 (N_10621,N_5814,N_6275);
and U10622 (N_10622,N_5298,N_7024);
nand U10623 (N_10623,N_8059,N_9085);
or U10624 (N_10624,N_9019,N_9234);
or U10625 (N_10625,N_5708,N_9296);
xnor U10626 (N_10626,N_7324,N_7490);
and U10627 (N_10627,N_7180,N_5735);
nand U10628 (N_10628,N_6070,N_6041);
and U10629 (N_10629,N_7932,N_7985);
nor U10630 (N_10630,N_7245,N_9917);
or U10631 (N_10631,N_8733,N_6660);
nor U10632 (N_10632,N_7477,N_9593);
and U10633 (N_10633,N_8766,N_8220);
or U10634 (N_10634,N_7676,N_5885);
xor U10635 (N_10635,N_8093,N_7167);
nand U10636 (N_10636,N_9786,N_8094);
nor U10637 (N_10637,N_6116,N_9400);
or U10638 (N_10638,N_5944,N_8234);
xor U10639 (N_10639,N_7393,N_6590);
xor U10640 (N_10640,N_8833,N_7782);
nor U10641 (N_10641,N_6748,N_9326);
nor U10642 (N_10642,N_9854,N_7100);
nand U10643 (N_10643,N_7897,N_8440);
or U10644 (N_10644,N_5640,N_9199);
nor U10645 (N_10645,N_8024,N_8654);
xor U10646 (N_10646,N_8661,N_9207);
xnor U10647 (N_10647,N_6509,N_7572);
nand U10648 (N_10648,N_6528,N_8313);
xnor U10649 (N_10649,N_9126,N_9624);
nor U10650 (N_10650,N_9287,N_7909);
and U10651 (N_10651,N_7819,N_7862);
nor U10652 (N_10652,N_9219,N_6867);
xnor U10653 (N_10653,N_5263,N_7082);
or U10654 (N_10654,N_8583,N_9868);
nor U10655 (N_10655,N_8504,N_7374);
and U10656 (N_10656,N_5205,N_5348);
or U10657 (N_10657,N_7051,N_9771);
or U10658 (N_10658,N_8057,N_5895);
xnor U10659 (N_10659,N_7669,N_7113);
and U10660 (N_10660,N_7178,N_9689);
nand U10661 (N_10661,N_7599,N_5775);
or U10662 (N_10662,N_8424,N_9252);
or U10663 (N_10663,N_7906,N_8614);
or U10664 (N_10664,N_7484,N_7703);
or U10665 (N_10665,N_7530,N_7665);
or U10666 (N_10666,N_8862,N_8572);
nand U10667 (N_10667,N_6189,N_7719);
nand U10668 (N_10668,N_5599,N_6746);
nor U10669 (N_10669,N_5285,N_7632);
nand U10670 (N_10670,N_7991,N_8506);
nand U10671 (N_10671,N_5543,N_8222);
and U10672 (N_10672,N_9333,N_9334);
nor U10673 (N_10673,N_7361,N_6402);
nor U10674 (N_10674,N_7651,N_7867);
nand U10675 (N_10675,N_9994,N_8804);
or U10676 (N_10676,N_6860,N_8595);
xnor U10677 (N_10677,N_7548,N_9573);
xor U10678 (N_10678,N_6037,N_7421);
nand U10679 (N_10679,N_5831,N_7314);
and U10680 (N_10680,N_5836,N_5511);
or U10681 (N_10681,N_7002,N_9332);
or U10682 (N_10682,N_6814,N_8127);
nand U10683 (N_10683,N_5135,N_8613);
xor U10684 (N_10684,N_9314,N_5910);
and U10685 (N_10685,N_6651,N_7270);
nor U10686 (N_10686,N_6529,N_9002);
nand U10687 (N_10687,N_5840,N_9322);
and U10688 (N_10688,N_5781,N_8119);
nand U10689 (N_10689,N_6340,N_8685);
and U10690 (N_10690,N_9033,N_6084);
nand U10691 (N_10691,N_7499,N_5641);
xnor U10692 (N_10692,N_7127,N_9066);
or U10693 (N_10693,N_5875,N_5318);
nor U10694 (N_10694,N_7841,N_6635);
nand U10695 (N_10695,N_7959,N_6458);
nor U10696 (N_10696,N_9780,N_8906);
xnor U10697 (N_10697,N_8212,N_5638);
nand U10698 (N_10698,N_8269,N_7214);
nor U10699 (N_10699,N_5386,N_7627);
and U10700 (N_10700,N_6823,N_7142);
nor U10701 (N_10701,N_7050,N_8213);
nor U10702 (N_10702,N_9940,N_5790);
nand U10703 (N_10703,N_5624,N_7820);
and U10704 (N_10704,N_7845,N_7753);
nand U10705 (N_10705,N_8687,N_5618);
and U10706 (N_10706,N_7697,N_5815);
and U10707 (N_10707,N_5190,N_7673);
nand U10708 (N_10708,N_9553,N_8218);
or U10709 (N_10709,N_8758,N_5981);
nand U10710 (N_10710,N_9657,N_7383);
xor U10711 (N_10711,N_9122,N_5498);
and U10712 (N_10712,N_5768,N_9572);
nand U10713 (N_10713,N_5130,N_5681);
nor U10714 (N_10714,N_9923,N_8702);
nor U10715 (N_10715,N_8626,N_9406);
nor U10716 (N_10716,N_6641,N_9790);
nor U10717 (N_10717,N_7949,N_9509);
nor U10718 (N_10718,N_8843,N_5479);
or U10719 (N_10719,N_8162,N_9681);
xnor U10720 (N_10720,N_5554,N_7683);
xnor U10721 (N_10721,N_9800,N_7432);
and U10722 (N_10722,N_9457,N_7465);
nand U10723 (N_10723,N_9378,N_9753);
nor U10724 (N_10724,N_6532,N_6141);
or U10725 (N_10725,N_8151,N_7520);
nand U10726 (N_10726,N_7750,N_8085);
xnor U10727 (N_10727,N_5210,N_6333);
nor U10728 (N_10728,N_7717,N_6250);
nand U10729 (N_10729,N_7571,N_6176);
and U10730 (N_10730,N_6919,N_9488);
or U10731 (N_10731,N_9384,N_9130);
nor U10732 (N_10732,N_6241,N_8887);
or U10733 (N_10733,N_9341,N_9906);
nor U10734 (N_10734,N_9747,N_7510);
xor U10735 (N_10735,N_6772,N_6698);
or U10736 (N_10736,N_5060,N_9253);
or U10737 (N_10737,N_8029,N_5178);
xnor U10738 (N_10738,N_8433,N_6602);
and U10739 (N_10739,N_5033,N_6991);
or U10740 (N_10740,N_6271,N_8788);
and U10741 (N_10741,N_9972,N_8905);
xnor U10742 (N_10742,N_8945,N_9254);
nand U10743 (N_10743,N_6043,N_8470);
or U10744 (N_10744,N_5703,N_5417);
and U10745 (N_10745,N_5696,N_9481);
nor U10746 (N_10746,N_9116,N_9008);
nand U10747 (N_10747,N_9281,N_8341);
or U10748 (N_10748,N_5080,N_9494);
nand U10749 (N_10749,N_5246,N_6753);
xor U10750 (N_10750,N_5458,N_8600);
and U10751 (N_10751,N_5666,N_9551);
nor U10752 (N_10752,N_8207,N_7618);
xor U10753 (N_10753,N_5034,N_7811);
nand U10754 (N_10754,N_6436,N_9587);
nand U10755 (N_10755,N_9335,N_7474);
xor U10756 (N_10756,N_5144,N_6485);
or U10757 (N_10757,N_7378,N_8446);
and U10758 (N_10758,N_5028,N_5947);
xnor U10759 (N_10759,N_5648,N_5850);
and U10760 (N_10760,N_6950,N_7150);
and U10761 (N_10761,N_8267,N_6167);
nor U10762 (N_10762,N_9416,N_8327);
or U10763 (N_10763,N_7509,N_7783);
or U10764 (N_10764,N_9644,N_7304);
nor U10765 (N_10765,N_5237,N_7168);
or U10766 (N_10766,N_5098,N_6859);
nor U10767 (N_10767,N_8427,N_8620);
nor U10768 (N_10768,N_9810,N_5984);
xor U10769 (N_10769,N_5616,N_7105);
nand U10770 (N_10770,N_7170,N_5715);
nand U10771 (N_10771,N_9629,N_5242);
xor U10772 (N_10772,N_5376,N_5727);
or U10773 (N_10773,N_5311,N_5832);
and U10774 (N_10774,N_8954,N_5752);
nor U10775 (N_10775,N_7014,N_7156);
or U10776 (N_10776,N_7288,N_7578);
and U10777 (N_10777,N_9097,N_8156);
nor U10778 (N_10778,N_5202,N_8503);
or U10779 (N_10779,N_5180,N_7121);
and U10780 (N_10780,N_6834,N_5635);
or U10781 (N_10781,N_6797,N_7206);
and U10782 (N_10782,N_5954,N_9428);
or U10783 (N_10783,N_9879,N_6285);
and U10784 (N_10784,N_5539,N_7286);
xor U10785 (N_10785,N_6508,N_5568);
nor U10786 (N_10786,N_5716,N_9659);
nand U10787 (N_10787,N_8876,N_9282);
or U10788 (N_10788,N_9475,N_8990);
and U10789 (N_10789,N_9620,N_6119);
or U10790 (N_10790,N_5684,N_9731);
nor U10791 (N_10791,N_7224,N_7975);
and U10792 (N_10792,N_9145,N_8288);
and U10793 (N_10793,N_7463,N_9032);
nand U10794 (N_10794,N_9552,N_7766);
or U10795 (N_10795,N_5448,N_9987);
nor U10796 (N_10796,N_8142,N_9329);
nand U10797 (N_10797,N_9040,N_9755);
or U10798 (N_10798,N_5397,N_8167);
and U10799 (N_10799,N_5829,N_5209);
nand U10800 (N_10800,N_7426,N_5651);
and U10801 (N_10801,N_9931,N_5998);
nor U10802 (N_10802,N_5100,N_8088);
nand U10803 (N_10803,N_6270,N_8251);
nand U10804 (N_10804,N_5244,N_5907);
nor U10805 (N_10805,N_7229,N_5658);
or U10806 (N_10806,N_8500,N_9997);
and U10807 (N_10807,N_9949,N_7052);
or U10808 (N_10808,N_5749,N_9641);
and U10809 (N_10809,N_8860,N_9530);
xnor U10810 (N_10810,N_9634,N_6351);
xor U10811 (N_10811,N_7483,N_5043);
nand U10812 (N_10812,N_6811,N_5514);
or U10813 (N_10813,N_5988,N_5217);
nor U10814 (N_10814,N_9479,N_5748);
nand U10815 (N_10815,N_7234,N_9709);
or U10816 (N_10816,N_5569,N_7881);
or U10817 (N_10817,N_6907,N_6366);
or U10818 (N_10818,N_9320,N_7725);
xor U10819 (N_10819,N_9586,N_8292);
xnor U10820 (N_10820,N_8126,N_7540);
and U10821 (N_10821,N_5714,N_9260);
nor U10822 (N_10822,N_7503,N_9688);
and U10823 (N_10823,N_7239,N_7133);
and U10824 (N_10824,N_9200,N_5220);
nand U10825 (N_10825,N_6840,N_6580);
xor U10826 (N_10826,N_6894,N_7104);
nor U10827 (N_10827,N_6377,N_7800);
nand U10828 (N_10828,N_5137,N_7853);
xor U10829 (N_10829,N_9722,N_9051);
xnor U10830 (N_10830,N_7457,N_6690);
nand U10831 (N_10831,N_7854,N_7470);
xnor U10832 (N_10832,N_8982,N_8656);
or U10833 (N_10833,N_7191,N_9876);
xnor U10834 (N_10834,N_6759,N_5593);
nand U10835 (N_10835,N_8186,N_6579);
xor U10836 (N_10836,N_6525,N_5022);
nand U10837 (N_10837,N_7424,N_8918);
nor U10838 (N_10838,N_6222,N_5021);
nor U10839 (N_10839,N_9078,N_9594);
xnor U10840 (N_10840,N_5322,N_9088);
or U10841 (N_10841,N_6040,N_6062);
xor U10842 (N_10842,N_9102,N_9035);
nor U10843 (N_10843,N_6172,N_6916);
nor U10844 (N_10844,N_9957,N_9446);
or U10845 (N_10845,N_8770,N_9196);
nand U10846 (N_10846,N_5239,N_5667);
or U10847 (N_10847,N_9616,N_9767);
or U10848 (N_10848,N_6703,N_9635);
nor U10849 (N_10849,N_8552,N_9357);
nand U10850 (N_10850,N_9837,N_5474);
and U10851 (N_10851,N_9073,N_8955);
xor U10852 (N_10852,N_6059,N_6979);
and U10853 (N_10853,N_8719,N_5314);
nor U10854 (N_10854,N_5917,N_7889);
xnor U10855 (N_10855,N_7251,N_9037);
nand U10856 (N_10856,N_9958,N_9872);
or U10857 (N_10857,N_7573,N_5720);
nor U10858 (N_10858,N_7760,N_8474);
xor U10859 (N_10859,N_8061,N_6808);
and U10860 (N_10860,N_8439,N_9176);
and U10861 (N_10861,N_8551,N_6885);
nand U10862 (N_10862,N_5276,N_6150);
or U10863 (N_10863,N_6294,N_5861);
nand U10864 (N_10864,N_7724,N_8477);
nand U10865 (N_10865,N_8226,N_5093);
or U10866 (N_10866,N_7221,N_9541);
nand U10867 (N_10867,N_7707,N_8275);
or U10868 (N_10868,N_9953,N_8658);
and U10869 (N_10869,N_8927,N_7757);
nand U10870 (N_10870,N_9893,N_7609);
nand U10871 (N_10871,N_8306,N_7390);
nor U10872 (N_10872,N_6096,N_7585);
nand U10873 (N_10873,N_5750,N_7075);
or U10874 (N_10874,N_6963,N_6923);
nor U10875 (N_10875,N_5550,N_7714);
xor U10876 (N_10876,N_6578,N_7558);
nor U10877 (N_10877,N_6029,N_7446);
or U10878 (N_10878,N_5621,N_5573);
and U10879 (N_10879,N_5751,N_7939);
nor U10880 (N_10880,N_7149,N_8515);
xnor U10881 (N_10881,N_7823,N_9815);
nand U10882 (N_10882,N_6920,N_9251);
nor U10883 (N_10883,N_9661,N_5011);
nor U10884 (N_10884,N_6280,N_9833);
and U10885 (N_10885,N_6722,N_6645);
and U10886 (N_10886,N_5535,N_7344);
xor U10887 (N_10887,N_9143,N_9575);
and U10888 (N_10888,N_5691,N_5394);
nor U10889 (N_10889,N_5483,N_7060);
and U10890 (N_10890,N_5886,N_7215);
xnor U10891 (N_10891,N_5856,N_8068);
xnor U10892 (N_10892,N_7733,N_8618);
or U10893 (N_10893,N_5575,N_9164);
nor U10894 (N_10894,N_5029,N_5300);
or U10895 (N_10895,N_8375,N_8264);
nand U10896 (N_10896,N_6974,N_7681);
nor U10897 (N_10897,N_6382,N_6085);
and U10898 (N_10898,N_6068,N_7579);
nand U10899 (N_10899,N_6208,N_7634);
or U10900 (N_10900,N_5252,N_7482);
nor U10901 (N_10901,N_6164,N_8377);
or U10902 (N_10902,N_8731,N_5959);
nand U10903 (N_10903,N_6378,N_7679);
or U10904 (N_10904,N_5072,N_6014);
xor U10905 (N_10905,N_7646,N_7352);
or U10906 (N_10906,N_6584,N_8387);
nand U10907 (N_10907,N_5275,N_6832);
and U10908 (N_10908,N_5958,N_9420);
or U10909 (N_10909,N_6676,N_7856);
nor U10910 (N_10910,N_5661,N_6147);
nand U10911 (N_10911,N_5934,N_5046);
or U10912 (N_10912,N_8394,N_7095);
and U10913 (N_10913,N_6964,N_7054);
xnor U10914 (N_10914,N_5101,N_8316);
or U10915 (N_10915,N_6398,N_6559);
nor U10916 (N_10916,N_5457,N_8564);
xnor U10917 (N_10917,N_6117,N_7722);
or U10918 (N_10918,N_7455,N_8837);
xor U10919 (N_10919,N_9075,N_6307);
nor U10920 (N_10920,N_6573,N_7515);
nor U10921 (N_10921,N_7409,N_7855);
and U10922 (N_10922,N_5428,N_7190);
nor U10923 (N_10923,N_5526,N_7965);
or U10924 (N_10924,N_7351,N_8533);
or U10925 (N_10925,N_8824,N_8655);
nand U10926 (N_10926,N_9336,N_9433);
or U10927 (N_10927,N_6007,N_7320);
nand U10928 (N_10928,N_8253,N_8081);
xnor U10929 (N_10929,N_6219,N_6433);
and U10930 (N_10930,N_9932,N_6069);
nand U10931 (N_10931,N_7944,N_6732);
and U10932 (N_10932,N_9417,N_8473);
nor U10933 (N_10933,N_7486,N_7460);
xor U10934 (N_10934,N_8623,N_6005);
and U10935 (N_10935,N_8130,N_5841);
nand U10936 (N_10936,N_6909,N_7171);
or U10937 (N_10937,N_9432,N_5110);
or U10938 (N_10938,N_5250,N_8021);
and U10939 (N_10939,N_8732,N_5385);
or U10940 (N_10940,N_5865,N_8023);
and U10941 (N_10941,N_8121,N_9746);
and U10942 (N_10942,N_6455,N_7566);
and U10943 (N_10943,N_5337,N_5068);
xor U10944 (N_10944,N_6392,N_9670);
or U10945 (N_10945,N_6900,N_6185);
xor U10946 (N_10946,N_6344,N_6444);
nor U10947 (N_10947,N_7734,N_9901);
nor U10948 (N_10948,N_8946,N_6658);
and U10949 (N_10949,N_7692,N_8797);
or U10950 (N_10950,N_7981,N_6320);
or U10951 (N_10951,N_6010,N_5574);
or U10952 (N_10952,N_9632,N_5196);
and U10953 (N_10953,N_5597,N_7642);
xor U10954 (N_10954,N_5802,N_5158);
and U10955 (N_10955,N_6773,N_7542);
and U10956 (N_10956,N_7035,N_5733);
and U10957 (N_10957,N_8947,N_5801);
xnor U10958 (N_10958,N_6711,N_7347);
or U10959 (N_10959,N_9588,N_8521);
and U10960 (N_10960,N_6473,N_5625);
nor U10961 (N_10961,N_5352,N_5324);
and U10962 (N_10962,N_7443,N_5346);
and U10963 (N_10963,N_6875,N_8956);
nand U10964 (N_10964,N_7883,N_5310);
nor U10965 (N_10965,N_5067,N_5191);
nor U10966 (N_10966,N_5924,N_9838);
or U10967 (N_10967,N_7525,N_7601);
nor U10968 (N_10968,N_7762,N_5852);
nand U10969 (N_10969,N_5517,N_7093);
nor U10970 (N_10970,N_6336,N_8294);
and U10971 (N_10971,N_6254,N_9184);
or U10972 (N_10972,N_8467,N_7199);
xnor U10973 (N_10973,N_6434,N_5821);
nand U10974 (N_10974,N_9822,N_8531);
xor U10975 (N_10975,N_6679,N_5296);
nand U10976 (N_10976,N_7269,N_7942);
xnor U10977 (N_10977,N_7595,N_5653);
nand U10978 (N_10978,N_5007,N_8847);
xnor U10979 (N_10979,N_7439,N_5764);
or U10980 (N_10980,N_9820,N_8735);
nand U10981 (N_10981,N_5234,N_8348);
nor U10982 (N_10982,N_9272,N_7282);
or U10983 (N_10983,N_8782,N_7611);
and U10984 (N_10984,N_9503,N_8413);
nor U10985 (N_10985,N_9259,N_7401);
or U10986 (N_10986,N_5408,N_8767);
and U10987 (N_10987,N_5054,N_8721);
nor U10988 (N_10988,N_6846,N_7555);
xnor U10989 (N_10989,N_7157,N_6806);
xor U10990 (N_10990,N_8420,N_6321);
nor U10991 (N_10991,N_8823,N_8323);
or U10992 (N_10992,N_7858,N_5126);
and U10993 (N_10993,N_8370,N_7891);
nand U10994 (N_10994,N_7830,N_6977);
or U10995 (N_10995,N_7645,N_7129);
nand U10996 (N_10996,N_5723,N_9708);
nand U10997 (N_10997,N_5803,N_7362);
nor U10998 (N_10998,N_6319,N_9294);
or U10999 (N_10999,N_6572,N_5212);
or U11000 (N_11000,N_9666,N_7977);
and U11001 (N_11001,N_8750,N_8107);
or U11002 (N_11002,N_8928,N_7995);
or U11003 (N_11003,N_9700,N_8333);
and U11004 (N_11004,N_6506,N_7242);
and U11005 (N_11005,N_8851,N_9165);
or U11006 (N_11006,N_7207,N_9612);
nand U11007 (N_11007,N_7617,N_9858);
nand U11008 (N_11008,N_5940,N_7293);
nor U11009 (N_11009,N_8861,N_8636);
nand U11010 (N_11010,N_5739,N_8140);
and U11011 (N_11011,N_6568,N_7799);
nor U11012 (N_11012,N_9173,N_8888);
xor U11013 (N_11013,N_7365,N_6863);
xnor U11014 (N_11014,N_5463,N_5930);
or U11015 (N_11015,N_5676,N_6870);
nand U11016 (N_11016,N_5603,N_7325);
xnor U11017 (N_11017,N_9072,N_8249);
xnor U11018 (N_11018,N_6152,N_6890);
and U11019 (N_11019,N_6237,N_8894);
or U11020 (N_11020,N_8706,N_8334);
nand U11021 (N_11021,N_9411,N_9262);
and U11022 (N_11022,N_7682,N_6597);
xor U11023 (N_11023,N_9680,N_7042);
nor U11024 (N_11024,N_6954,N_6144);
and U11025 (N_11025,N_5170,N_9077);
xnor U11026 (N_11026,N_5631,N_9981);
xor U11027 (N_11027,N_8410,N_5565);
nor U11028 (N_11028,N_6911,N_7197);
nand U11029 (N_11029,N_7194,N_5232);
xor U11030 (N_11030,N_9592,N_8076);
xor U11031 (N_11031,N_6456,N_9834);
nand U11032 (N_11032,N_8122,N_6474);
or U11033 (N_11033,N_8418,N_6022);
nand U11034 (N_11034,N_7888,N_6469);
or U11035 (N_11035,N_6586,N_5277);
and U11036 (N_11036,N_6013,N_6438);
nand U11037 (N_11037,N_8986,N_5269);
nor U11038 (N_11038,N_7805,N_8237);
nor U11039 (N_11039,N_8790,N_5172);
nand U11040 (N_11040,N_8752,N_7152);
xnor U11041 (N_11041,N_8461,N_6644);
xnor U11042 (N_11042,N_8257,N_8411);
xor U11043 (N_11043,N_9459,N_6871);
xnor U11044 (N_11044,N_8690,N_8419);
xnor U11045 (N_11045,N_5496,N_5963);
or U11046 (N_11046,N_7550,N_9845);
or U11047 (N_11047,N_9859,N_6211);
and U11048 (N_11048,N_6421,N_5928);
xor U11049 (N_11049,N_7254,N_6914);
or U11050 (N_11050,N_6180,N_9888);
nand U11051 (N_11051,N_6784,N_6982);
nand U11052 (N_11052,N_8149,N_5219);
nand U11053 (N_11053,N_5192,N_6718);
nor U11054 (N_11054,N_9513,N_9534);
or U11055 (N_11055,N_5783,N_9489);
nand U11056 (N_11056,N_7466,N_8507);
or U11057 (N_11057,N_8233,N_5459);
nor U11058 (N_11058,N_9602,N_9471);
nor U11059 (N_11059,N_9209,N_9679);
nor U11060 (N_11060,N_7816,N_5392);
xnor U11061 (N_11061,N_8211,N_6054);
nand U11062 (N_11062,N_8581,N_8339);
nor U11063 (N_11063,N_8310,N_8633);
and U11064 (N_11064,N_7294,N_8189);
xnor U11065 (N_11065,N_9222,N_5113);
nor U11066 (N_11066,N_6794,N_7238);
or U11067 (N_11067,N_6926,N_6012);
and U11068 (N_11068,N_9027,N_9783);
nor U11069 (N_11069,N_5807,N_5868);
xnor U11070 (N_11070,N_8184,N_8743);
and U11071 (N_11071,N_8863,N_7612);
and U11072 (N_11072,N_7074,N_5183);
or U11073 (N_11073,N_9584,N_8637);
nor U11074 (N_11074,N_6607,N_9577);
nor U11075 (N_11075,N_9968,N_5901);
or U11076 (N_11076,N_9982,N_8066);
nor U11077 (N_11077,N_7545,N_8143);
nand U11078 (N_11078,N_5818,N_5811);
nand U11079 (N_11079,N_7353,N_5157);
nand U11080 (N_11080,N_5610,N_9849);
or U11081 (N_11081,N_6699,N_8342);
nor U11082 (N_11082,N_5421,N_8592);
nand U11083 (N_11083,N_7552,N_7814);
and U11084 (N_11084,N_5797,N_8746);
or U11085 (N_11085,N_9985,N_8185);
nand U11086 (N_11086,N_5893,N_6122);
or U11087 (N_11087,N_7803,N_8457);
nand U11088 (N_11088,N_8345,N_9091);
nand U11089 (N_11089,N_8809,N_8671);
nand U11090 (N_11090,N_8812,N_6705);
xor U11091 (N_11091,N_5500,N_8680);
or U11092 (N_11092,N_9427,N_7009);
nor U11093 (N_11093,N_6629,N_6009);
nand U11094 (N_11094,N_8291,N_9487);
nand U11095 (N_11095,N_8315,N_5268);
xor U11096 (N_11096,N_9389,N_5439);
nor U11097 (N_11097,N_9377,N_8855);
and U11098 (N_11098,N_9757,N_7928);
and U11099 (N_11099,N_9181,N_5950);
and U11100 (N_11100,N_5032,N_5991);
or U11101 (N_11101,N_7334,N_6129);
or U11102 (N_11102,N_9067,N_8765);
nor U11103 (N_11103,N_9017,N_7475);
or U11104 (N_11104,N_9969,N_9765);
nand U11105 (N_11105,N_7598,N_5169);
or U11106 (N_11106,N_5270,N_5257);
and U11107 (N_11107,N_5462,N_6634);
nor U11108 (N_11108,N_9855,N_9693);
and U11109 (N_11109,N_5718,N_6831);
nand U11110 (N_11110,N_6403,N_8900);
nand U11111 (N_11111,N_7979,N_6417);
and U11112 (N_11112,N_6060,N_9022);
and U11113 (N_11113,N_8594,N_5966);
and U11114 (N_11114,N_6726,N_7306);
and U11115 (N_11115,N_6886,N_5711);
nor U11116 (N_11116,N_5096,N_9380);
nor U11117 (N_11117,N_7739,N_5443);
xor U11118 (N_11118,N_9836,N_9491);
xnor U11119 (N_11119,N_5977,N_6296);
or U11120 (N_11120,N_9823,N_6809);
xor U11121 (N_11121,N_8077,N_6952);
nor U11122 (N_11122,N_5366,N_8187);
and U11123 (N_11123,N_7125,N_5245);
or U11124 (N_11124,N_5547,N_5538);
or U11125 (N_11125,N_9582,N_9342);
or U11126 (N_11126,N_8781,N_8883);
nand U11127 (N_11127,N_9440,N_9549);
and U11128 (N_11128,N_9374,N_9456);
nor U11129 (N_11129,N_6313,N_8388);
nor U11130 (N_11130,N_6628,N_6290);
nor U11131 (N_11131,N_5334,N_6623);
xnor U11132 (N_11132,N_6659,N_8760);
xnor U11133 (N_11133,N_6197,N_9099);
nor U11134 (N_11134,N_5796,N_5419);
or U11135 (N_11135,N_6539,N_8983);
xor U11136 (N_11136,N_5248,N_5905);
nand U11137 (N_11137,N_8647,N_7076);
and U11138 (N_11138,N_5507,N_8713);
and U11139 (N_11139,N_9108,N_6404);
nand U11140 (N_11140,N_9127,N_6099);
and U11141 (N_11141,N_9140,N_9806);
or U11142 (N_11142,N_6662,N_8688);
nand U11143 (N_11143,N_7622,N_6868);
nor U11144 (N_11144,N_7342,N_6760);
and U11145 (N_11145,N_8818,N_7776);
nor U11146 (N_11146,N_8802,N_6899);
nor U11147 (N_11147,N_9194,N_6479);
nor U11148 (N_11148,N_5728,N_9285);
nand U11149 (N_11149,N_5975,N_6139);
and U11150 (N_11150,N_5990,N_6407);
nand U11151 (N_11151,N_6030,N_7192);
or U11152 (N_11152,N_5339,N_8932);
nor U11153 (N_11153,N_6767,N_9450);
nand U11154 (N_11154,N_6089,N_5654);
or U11155 (N_11155,N_8296,N_6905);
nor U11156 (N_11156,N_8764,N_9438);
and U11157 (N_11157,N_8025,N_9995);
or U11158 (N_11158,N_8309,N_6127);
nor U11159 (N_11159,N_9295,N_8022);
nand U11160 (N_11160,N_9662,N_9324);
xor U11161 (N_11161,N_8509,N_9279);
nor U11162 (N_11162,N_6109,N_6976);
nor U11163 (N_11163,N_9504,N_6100);
nand U11164 (N_11164,N_7764,N_6132);
nor U11165 (N_11165,N_9381,N_7857);
xnor U11166 (N_11166,N_8684,N_7835);
nand U11167 (N_11167,N_9599,N_5488);
or U11168 (N_11168,N_5710,N_7921);
nor U11169 (N_11169,N_7387,N_6527);
nand U11170 (N_11170,N_8892,N_6493);
and U11171 (N_11171,N_5918,N_9398);
nor U11172 (N_11172,N_6198,N_8745);
and U11173 (N_11173,N_5758,N_6672);
xor U11174 (N_11174,N_6476,N_7001);
and U11175 (N_11175,N_8116,N_9911);
and U11176 (N_11176,N_6067,N_7210);
nor U11177 (N_11177,N_5293,N_5744);
nor U11178 (N_11178,N_6656,N_9952);
or U11179 (N_11179,N_6639,N_5097);
nor U11180 (N_11180,N_6829,N_6393);
nand U11181 (N_11181,N_7091,N_5438);
xnor U11182 (N_11182,N_5003,N_9782);
nand U11183 (N_11183,N_8422,N_9269);
and U11184 (N_11184,N_5693,N_7296);
nand U11185 (N_11185,N_7523,N_8084);
xor U11186 (N_11186,N_8338,N_9918);
xnor U11187 (N_11187,N_7919,N_9787);
xnor U11188 (N_11188,N_5485,N_7730);
or U11189 (N_11189,N_9967,N_5855);
and U11190 (N_11190,N_5151,N_8828);
and U11191 (N_11191,N_5590,N_9707);
or U11192 (N_11192,N_9717,N_7620);
xor U11193 (N_11193,N_6242,N_5551);
or U11194 (N_11194,N_5048,N_7480);
nor U11195 (N_11195,N_8783,N_7328);
and U11196 (N_11196,N_5047,N_7015);
and U11197 (N_11197,N_7497,N_9580);
xor U11198 (N_11198,N_9742,N_7449);
or U11199 (N_11199,N_9436,N_6615);
nor U11200 (N_11200,N_5770,N_8739);
nor U11201 (N_11201,N_9795,N_6065);
xnor U11202 (N_11202,N_8139,N_7267);
nor U11203 (N_11203,N_6173,N_5772);
nand U11204 (N_11204,N_8166,N_8241);
nand U11205 (N_11205,N_7570,N_5027);
xnor U11206 (N_11206,N_5226,N_9113);
nand U11207 (N_11207,N_7647,N_9614);
nor U11208 (N_11208,N_8054,N_8881);
xnor U11209 (N_11209,N_6769,N_9885);
nand U11210 (N_11210,N_9963,N_6793);
nand U11211 (N_11211,N_5053,N_7166);
xnor U11212 (N_11212,N_6115,N_5347);
nand U11213 (N_11213,N_7059,N_6613);
and U11214 (N_11214,N_6847,N_6956);
nand U11215 (N_11215,N_6168,N_6915);
nand U11216 (N_11216,N_6595,N_8136);
and U11217 (N_11217,N_7441,N_6345);
and U11218 (N_11218,N_7338,N_9171);
and U11219 (N_11219,N_6792,N_5904);
nor U11220 (N_11220,N_9092,N_8262);
nand U11221 (N_11221,N_6210,N_5578);
and U11222 (N_11222,N_5843,N_7311);
nor U11223 (N_11223,N_5501,N_6225);
xor U11224 (N_11224,N_7920,N_8118);
xnor U11225 (N_11225,N_8487,N_8216);
and U11226 (N_11226,N_9338,N_7494);
nand U11227 (N_11227,N_9258,N_8270);
and U11228 (N_11228,N_9847,N_9238);
nand U11229 (N_11229,N_5437,N_9863);
xnor U11230 (N_11230,N_9664,N_5320);
and U11231 (N_11231,N_9469,N_8284);
xnor U11232 (N_11232,N_6545,N_5767);
or U11233 (N_11233,N_9046,N_7538);
and U11234 (N_11234,N_5518,N_6526);
nor U11235 (N_11235,N_7710,N_7918);
and U11236 (N_11236,N_5871,N_9093);
nand U11237 (N_11237,N_9581,N_5453);
nor U11238 (N_11238,N_7272,N_9277);
and U11239 (N_11239,N_6376,N_9913);
and U11240 (N_11240,N_9660,N_9734);
nor U11241 (N_11241,N_5393,N_9774);
or U11242 (N_11242,N_5582,N_5251);
xor U11243 (N_11243,N_6609,N_6359);
xor U11244 (N_11244,N_8062,N_9180);
nor U11245 (N_11245,N_8409,N_7256);
nand U11246 (N_11246,N_9267,N_9345);
nand U11247 (N_11247,N_5897,N_5657);
or U11248 (N_11248,N_7447,N_8622);
or U11249 (N_11249,N_6300,N_9425);
nor U11250 (N_11250,N_8964,N_7479);
and U11251 (N_11251,N_6906,N_7265);
xor U11252 (N_11252,N_7123,N_7109);
xnor U11253 (N_11253,N_7416,N_7185);
xor U11254 (N_11254,N_9941,N_6556);
or U11255 (N_11255,N_5140,N_8476);
nor U11256 (N_11256,N_9021,N_6826);
nand U11257 (N_11257,N_7973,N_9658);
and U11258 (N_11258,N_5193,N_9235);
or U11259 (N_11259,N_6269,N_5230);
nand U11260 (N_11260,N_8358,N_5173);
nand U11261 (N_11261,N_5208,N_9168);
and U11262 (N_11262,N_9891,N_9807);
xor U11263 (N_11263,N_7689,N_8775);
and U11264 (N_11264,N_5707,N_9915);
xnor U11265 (N_11265,N_9545,N_5211);
or U11266 (N_11266,N_8692,N_5932);
nor U11267 (N_11267,N_5349,N_9016);
nand U11268 (N_11268,N_9197,N_8049);
nor U11269 (N_11269,N_8926,N_5709);
xor U11270 (N_11270,N_8569,N_5747);
and U11271 (N_11271,N_5552,N_7504);
or U11272 (N_11272,N_5389,N_9719);
nand U11273 (N_11273,N_7061,N_9148);
nand U11274 (N_11274,N_5460,N_6268);
xnor U11275 (N_11275,N_9330,N_9054);
nand U11276 (N_11276,N_8631,N_7310);
and U11277 (N_11277,N_7301,N_7582);
nor U11278 (N_11278,N_5846,N_7500);
nand U11279 (N_11279,N_9216,N_9792);
nor U11280 (N_11280,N_7163,N_7527);
nand U11281 (N_11281,N_7990,N_7151);
and U11282 (N_11282,N_9364,N_8236);
nand U11283 (N_11283,N_8163,N_9388);
and U11284 (N_11284,N_5292,N_9407);
nor U11285 (N_11285,N_8133,N_7755);
and U11286 (N_11286,N_8559,N_7934);
or U11287 (N_11287,N_9458,N_9190);
and U11288 (N_11288,N_5008,N_6861);
or U11289 (N_11289,N_8696,N_8101);
nand U11290 (N_11290,N_5766,N_8726);
or U11291 (N_11291,N_9619,N_6325);
nand U11292 (N_11292,N_7706,N_7899);
nor U11293 (N_11293,N_6883,N_7081);
nor U11294 (N_11294,N_6226,N_6521);
xor U11295 (N_11295,N_9590,N_9484);
nor U11296 (N_11296,N_9257,N_7321);
and U11297 (N_11297,N_6466,N_5887);
and U11298 (N_11298,N_8415,N_8563);
or U11299 (N_11299,N_7652,N_7563);
and U11300 (N_11300,N_9043,N_7292);
xnor U11301 (N_11301,N_6273,N_5506);
nand U11302 (N_11302,N_8437,N_8794);
nor U11303 (N_11303,N_6016,N_7781);
and U11304 (N_11304,N_9653,N_6429);
xor U11305 (N_11305,N_8902,N_5450);
xor U11306 (N_11306,N_9754,N_7993);
or U11307 (N_11307,N_7017,N_5650);
or U11308 (N_11308,N_9359,N_7153);
nor U11309 (N_11309,N_9777,N_8836);
or U11310 (N_11310,N_5926,N_6216);
xnor U11311 (N_11311,N_7727,N_5216);
and U11312 (N_11312,N_9449,N_9947);
nand U11313 (N_11313,N_7458,N_7188);
or U11314 (N_11314,N_5845,N_5788);
or U11315 (N_11315,N_9429,N_5531);
nor U11316 (N_11316,N_8244,N_8640);
xor U11317 (N_11317,N_7376,N_7326);
xor U11318 (N_11318,N_9844,N_9023);
xnor U11319 (N_11319,N_6632,N_5030);
xor U11320 (N_11320,N_6229,N_7073);
and U11321 (N_11321,N_6001,N_9846);
or U11322 (N_11322,N_6751,N_8364);
or U11323 (N_11323,N_6426,N_5520);
nor U11324 (N_11324,N_8557,N_7189);
nor U11325 (N_11325,N_9654,N_6857);
xnor U11326 (N_11326,N_6078,N_5706);
or U11327 (N_11327,N_6948,N_8920);
nand U11328 (N_11328,N_9912,N_6953);
nand U11329 (N_11329,N_7227,N_5259);
and U11330 (N_11330,N_5171,N_5690);
and U11331 (N_11331,N_6511,N_7261);
xor U11332 (N_11332,N_5835,N_7305);
and U11333 (N_11333,N_6891,N_8090);
and U11334 (N_11334,N_9178,N_7057);
or U11335 (N_11335,N_8831,N_5813);
xnor U11336 (N_11336,N_9929,N_6049);
or U11337 (N_11337,N_6177,N_8434);
nand U11338 (N_11338,N_9470,N_7172);
and U11339 (N_11339,N_8402,N_5107);
xor U11340 (N_11340,N_6661,N_8710);
xnor U11341 (N_11341,N_8362,N_5849);
and U11342 (N_11342,N_6838,N_8123);
nand U11343 (N_11343,N_8890,N_8058);
nor U11344 (N_11344,N_6362,N_9245);
xnor U11345 (N_11345,N_9480,N_9499);
or U11346 (N_11346,N_7145,N_6470);
nand U11347 (N_11347,N_6312,N_8700);
or U11348 (N_11348,N_6125,N_6562);
or U11349 (N_11349,N_5063,N_7915);
and U11350 (N_11350,N_6516,N_6709);
or U11351 (N_11351,N_8356,N_8043);
or U11352 (N_11352,N_6762,N_8052);
nand U11353 (N_11353,N_5444,N_8177);
nor U11354 (N_11354,N_8491,N_7524);
or U11355 (N_11355,N_8188,N_9685);
and U11356 (N_11356,N_8598,N_8438);
nor U11357 (N_11357,N_9136,N_6962);
xnor U11358 (N_11358,N_5338,N_9124);
xnor U11359 (N_11359,N_5229,N_8223);
xor U11360 (N_11360,N_6807,N_8785);
nor U11361 (N_11361,N_9186,N_9711);
nand U11362 (N_11362,N_6372,N_8355);
or U11363 (N_11363,N_8493,N_5787);
nand U11364 (N_11364,N_6478,N_5951);
or U11365 (N_11365,N_9519,N_6631);
and U11366 (N_11366,N_9193,N_9177);
and U11367 (N_11367,N_7779,N_6118);
and U11368 (N_11368,N_5013,N_9925);
nand U11369 (N_11369,N_8464,N_5019);
or U11370 (N_11370,N_5390,N_8326);
and U11371 (N_11371,N_5384,N_6657);
and U11372 (N_11372,N_6088,N_5823);
or U11373 (N_11373,N_8352,N_6843);
nor U11374 (N_11374,N_5600,N_6754);
and U11375 (N_11375,N_9516,N_6889);
or U11376 (N_11376,N_9505,N_7517);
and U11377 (N_11377,N_5052,N_7615);
nand U11378 (N_11378,N_8086,N_6170);
nand U11379 (N_11379,N_6044,N_8378);
or U11380 (N_11380,N_6460,N_9776);
xnor U11381 (N_11381,N_6182,N_8176);
and U11382 (N_11382,N_7405,N_8368);
xnor U11383 (N_11383,N_5138,N_9137);
xnor U11384 (N_11384,N_5124,N_9478);
nand U11385 (N_11385,N_9030,N_9569);
nand U11386 (N_11386,N_8997,N_9699);
xnor U11387 (N_11387,N_5424,N_5800);
and U11388 (N_11388,N_8462,N_9498);
nor U11389 (N_11389,N_9959,N_5420);
nand U11390 (N_11390,N_8239,N_7037);
and U11391 (N_11391,N_7246,N_6642);
nor U11392 (N_11392,N_9603,N_7445);
or U11393 (N_11393,N_8276,N_5889);
nor U11394 (N_11394,N_9405,N_6151);
or U11395 (N_11395,N_5794,N_7413);
nor U11396 (N_11396,N_8458,N_9361);
nor U11397 (N_11397,N_8452,N_7055);
or U11398 (N_11398,N_6707,N_8576);
nor U11399 (N_11399,N_8100,N_6365);
nor U11400 (N_11400,N_7020,N_7894);
xor U11401 (N_11401,N_8643,N_6288);
and U11402 (N_11402,N_8357,N_7745);
nor U11403 (N_11403,N_5309,N_9397);
or U11404 (N_11404,N_9239,N_5615);
nand U11405 (N_11405,N_8738,N_6217);
or U11406 (N_11406,N_6704,N_6587);
nand U11407 (N_11407,N_8916,N_7533);
nand U11408 (N_11408,N_5837,N_5587);
xor U11409 (N_11409,N_8773,N_6371);
and U11410 (N_11410,N_6025,N_6810);
nand U11411 (N_11411,N_9315,N_8715);
and U11412 (N_11412,N_6200,N_8644);
nor U11413 (N_11413,N_5373,N_5973);
or U11414 (N_11414,N_8135,N_6181);
nand U11415 (N_11415,N_7631,N_7957);
xnor U11416 (N_11416,N_5406,N_6087);
nor U11417 (N_11417,N_8016,N_6178);
nand U11418 (N_11418,N_8321,N_9005);
xnor U11419 (N_11419,N_6329,N_5410);
nor U11420 (N_11420,N_5036,N_9015);
and U11421 (N_11421,N_9006,N_6191);
and U11422 (N_11422,N_9547,N_6577);
and U11423 (N_11423,N_9686,N_5001);
nor U11424 (N_11424,N_6123,N_6498);
xnor U11425 (N_11425,N_9211,N_5734);
xnor U11426 (N_11426,N_5466,N_5754);
nand U11427 (N_11427,N_6779,N_6006);
or U11428 (N_11428,N_6315,N_7005);
nand U11429 (N_11429,N_9977,N_8277);
xnor U11430 (N_11430,N_6090,N_8032);
nand U11431 (N_11431,N_7496,N_7103);
nand U11432 (N_11432,N_7736,N_8988);
and U11433 (N_11433,N_5848,N_6892);
and U11434 (N_11434,N_6183,N_8456);
nor U11435 (N_11435,N_7007,N_7241);
nand U11436 (N_11436,N_9889,N_7204);
and U11437 (N_11437,N_8210,N_5154);
nor U11438 (N_11438,N_8208,N_9618);
or U11439 (N_11439,N_9948,N_5085);
nor U11440 (N_11440,N_7516,N_9993);
nor U11441 (N_11441,N_7663,N_6227);
xor U11442 (N_11442,N_6844,N_6260);
and U11443 (N_11443,N_9527,N_9860);
nor U11444 (N_11444,N_7240,N_6047);
xnor U11445 (N_11445,N_5884,N_8204);
and U11446 (N_11446,N_9501,N_6818);
nand U11447 (N_11447,N_6864,N_7997);
and U11448 (N_11448,N_6353,N_7072);
xor U11449 (N_11449,N_5697,N_7430);
nand U11450 (N_11450,N_5497,N_5867);
nand U11451 (N_11451,N_8722,N_6138);
xor U11452 (N_11452,N_8772,N_8193);
nor U11453 (N_11453,N_6519,N_5454);
and U11454 (N_11454,N_5018,N_6379);
or U11455 (N_11455,N_5557,N_8774);
nand U11456 (N_11456,N_6231,N_9650);
xor U11457 (N_11457,N_6335,N_5609);
nand U11458 (N_11458,N_6700,N_9368);
nand U11459 (N_11459,N_8584,N_8698);
and U11460 (N_11460,N_6224,N_8998);
or U11461 (N_11461,N_7268,N_9939);
and U11462 (N_11462,N_8301,N_8977);
xnor U11463 (N_11463,N_9554,N_6399);
xor U11464 (N_11464,N_6228,N_5492);
or U11465 (N_11465,N_7913,N_7064);
nand U11466 (N_11466,N_5150,N_5765);
xor U11467 (N_11467,N_6415,N_8816);
nand U11468 (N_11468,N_7033,N_6790);
or U11469 (N_11469,N_6716,N_8938);
or U11470 (N_11470,N_8742,N_7205);
or U11471 (N_11471,N_5933,N_7597);
xor U11472 (N_11472,N_5833,N_5155);
nand U11473 (N_11473,N_8520,N_5353);
and U11474 (N_11474,N_8238,N_7828);
xor U11475 (N_11475,N_9003,N_5838);
or U11476 (N_11476,N_6984,N_8839);
nor U11477 (N_11477,N_5120,N_8695);
and U11478 (N_11478,N_6653,N_7831);
nor U11479 (N_11479,N_8660,N_6292);
and U11480 (N_11480,N_8565,N_9070);
nor U11481 (N_11481,N_5628,N_8603);
or U11482 (N_11482,N_9903,N_7635);
xor U11483 (N_11483,N_8335,N_7471);
nand U11484 (N_11484,N_5527,N_6032);
nand U11485 (N_11485,N_7077,N_6221);
xnor U11486 (N_11486,N_7257,N_7936);
nand U11487 (N_11487,N_8611,N_7958);
and U11488 (N_11488,N_5446,N_8874);
or U11489 (N_11489,N_7323,N_6026);
nand U11490 (N_11490,N_6888,N_5729);
nor U11491 (N_11491,N_6599,N_6256);
nand U11492 (N_11492,N_7720,N_9292);
and U11493 (N_11493,N_8840,N_8736);
nand U11494 (N_11494,N_6018,N_6038);
nand U11495 (N_11495,N_6350,N_5719);
nand U11496 (N_11496,N_5241,N_6801);
nor U11497 (N_11497,N_7923,N_9990);
xnor U11498 (N_11498,N_5741,N_8235);
xor U11499 (N_11499,N_6723,N_8757);
or U11500 (N_11500,N_5407,N_5515);
nand U11501 (N_11501,N_6989,N_6633);
xnor U11502 (N_11502,N_5247,N_7626);
xnor U11503 (N_11503,N_6604,N_7488);
or U11504 (N_11504,N_8047,N_7394);
or U11505 (N_11505,N_5655,N_8171);
and U11506 (N_11506,N_8412,N_8771);
nor U11507 (N_11507,N_6079,N_6282);
nand U11508 (N_11508,N_7765,N_6031);
xnor U11509 (N_11509,N_8478,N_8615);
or U11510 (N_11510,N_6785,N_9422);
and U11511 (N_11511,N_8913,N_8383);
xnor U11512 (N_11512,N_6496,N_5325);
xnor U11513 (N_11513,N_9826,N_6541);
nand U11514 (N_11514,N_9928,N_8423);
nand U11515 (N_11515,N_5233,N_7956);
nor U11516 (N_11516,N_9313,N_5145);
and U11517 (N_11517,N_6380,N_5937);
xnor U11518 (N_11518,N_9518,N_9631);
nor U11519 (N_11519,N_6195,N_7358);
nor U11520 (N_11520,N_6209,N_5581);
or U11521 (N_11521,N_8232,N_9649);
xnor U11522 (N_11522,N_5378,N_7826);
nand U11523 (N_11523,N_9210,N_5869);
nor U11524 (N_11524,N_7511,N_8445);
xor U11525 (N_11525,N_8786,N_5738);
nand U11526 (N_11526,N_9803,N_7534);
and U11527 (N_11527,N_7444,N_9857);
xnor U11528 (N_11528,N_8381,N_5049);
xnor U11529 (N_11529,N_6626,N_9811);
or U11530 (N_11530,N_5165,N_8535);
xnor U11531 (N_11531,N_7237,N_7056);
xnor U11532 (N_11532,N_9564,N_7731);
xor U11533 (N_11533,N_5588,N_7519);
nor U11534 (N_11534,N_7068,N_6143);
nor U11535 (N_11535,N_9874,N_8134);
and U11536 (N_11536,N_8194,N_8035);
and U11537 (N_11537,N_6913,N_5004);
xor U11538 (N_11538,N_8071,N_7489);
nand U11539 (N_11539,N_9528,N_7285);
xnor U11540 (N_11540,N_5982,N_5863);
nor U11541 (N_11541,N_8215,N_7372);
nand U11542 (N_11542,N_5073,N_5642);
and U11543 (N_11543,N_7879,N_9215);
nand U11544 (N_11544,N_9225,N_8128);
or U11545 (N_11545,N_8571,N_8080);
xnor U11546 (N_11546,N_5128,N_6781);
nand U11547 (N_11547,N_7852,N_9460);
xor U11548 (N_11548,N_5358,N_8454);
or U11549 (N_11549,N_9415,N_8159);
nor U11550 (N_11550,N_7355,N_8429);
xnor U11551 (N_11551,N_7422,N_7772);
nor U11552 (N_11552,N_6220,N_7813);
nand U11553 (N_11553,N_8289,N_5323);
nor U11554 (N_11554,N_9937,N_7732);
nand U11555 (N_11555,N_8849,N_9317);
xor U11556 (N_11556,N_6996,N_8285);
xnor U11557 (N_11557,N_9608,N_8451);
xnor U11558 (N_11558,N_7574,N_8485);
and U11559 (N_11559,N_8593,N_6500);
and U11560 (N_11560,N_5643,N_9973);
and U11561 (N_11561,N_6428,N_7391);
nor U11562 (N_11562,N_7317,N_7176);
nor U11563 (N_11563,N_9839,N_9476);
nor U11564 (N_11564,N_9678,N_6725);
xnor U11565 (N_11565,N_7775,N_7080);
nand U11566 (N_11566,N_9559,N_7543);
nor U11567 (N_11567,N_7044,N_6204);
and U11568 (N_11568,N_9024,N_8108);
xnor U11569 (N_11569,N_7658,N_8740);
nand U11570 (N_11570,N_7564,N_9684);
nand U11571 (N_11571,N_8582,N_9960);
xor U11572 (N_11572,N_5952,N_9486);
nand U11573 (N_11573,N_8858,N_5411);
nor U11574 (N_11574,N_8949,N_5133);
xnor U11575 (N_11575,N_9323,N_9031);
nor U11576 (N_11576,N_8428,N_7937);
nor U11577 (N_11577,N_9956,N_7211);
nor U11578 (N_11578,N_5503,N_8318);
nor U11579 (N_11579,N_8730,N_5015);
or U11580 (N_11580,N_5491,N_7315);
and U11581 (N_11581,N_5812,N_9595);
nand U11582 (N_11582,N_8602,N_5017);
or U11583 (N_11583,N_7136,N_9367);
xnor U11584 (N_11584,N_8768,N_6708);
and U11585 (N_11585,N_8548,N_5639);
and U11586 (N_11586,N_9607,N_5164);
and U11587 (N_11587,N_7164,N_8925);
nor U11588 (N_11588,N_5221,N_8372);
nor U11589 (N_11589,N_8205,N_7287);
and U11590 (N_11590,N_9291,N_9921);
nand U11591 (N_11591,N_5902,N_6243);
xnor U11592 (N_11592,N_8198,N_9241);
xnor U11593 (N_11593,N_7938,N_6236);
or U11594 (N_11594,N_5668,N_8120);
nand U11595 (N_11595,N_6643,N_8904);
or U11596 (N_11596,N_5713,N_9106);
nor U11597 (N_11597,N_7982,N_7948);
xor U11598 (N_11598,N_5570,N_6877);
nor U11599 (N_11599,N_9387,N_6352);
and U11600 (N_11600,N_5070,N_6537);
or U11601 (N_11601,N_7437,N_5774);
nand U11602 (N_11602,N_8098,N_6574);
and U11603 (N_11603,N_8868,N_7117);
nor U11604 (N_11604,N_7735,N_9768);
nor U11605 (N_11605,N_7414,N_5139);
or U11606 (N_11606,N_6624,N_7741);
nand U11607 (N_11607,N_9026,N_6764);
nand U11608 (N_11608,N_7146,N_7662);
and U11609 (N_11609,N_6324,N_9724);
nor U11610 (N_11610,N_9627,N_6534);
xnor U11611 (N_11611,N_9571,N_6750);
xor U11612 (N_11612,N_5223,N_6384);
nand U11613 (N_11613,N_7604,N_9525);
nor U11614 (N_11614,N_7019,N_6401);
xnor U11615 (N_11615,N_5343,N_6420);
or U11616 (N_11616,N_7562,N_7512);
and U11617 (N_11617,N_9760,N_9316);
or U11618 (N_11618,N_6154,N_9933);
and U11619 (N_11619,N_9270,N_9212);
xnor U11620 (N_11620,N_7384,N_9096);
nor U11621 (N_11621,N_9701,N_6114);
xor U11622 (N_11622,N_7231,N_6258);
nand U11623 (N_11623,N_6594,N_9399);
xor U11624 (N_11624,N_8796,N_7882);
nor U11625 (N_11625,N_5929,N_5472);
nand U11626 (N_11626,N_7874,N_7225);
nor U11627 (N_11627,N_5379,N_9466);
nand U11628 (N_11628,N_6782,N_6872);
nor U11629 (N_11629,N_9131,N_7359);
or U11630 (N_11630,N_7425,N_8787);
xnor U11631 (N_11631,N_8709,N_7825);
or U11632 (N_11632,N_6693,N_8003);
nand U11633 (N_11633,N_9598,N_5134);
nand U11634 (N_11634,N_6468,N_6975);
and U11635 (N_11635,N_5078,N_9883);
or U11636 (N_11636,N_9812,N_9922);
and U11637 (N_11637,N_8518,N_8607);
xnor U11638 (N_11638,N_6308,N_8897);
or U11639 (N_11639,N_9366,N_5786);
or U11640 (N_11640,N_8893,N_7748);
nand U11641 (N_11641,N_5743,N_5253);
or U11642 (N_11642,N_6232,N_7274);
or U11643 (N_11643,N_8838,N_7193);
and U11644 (N_11644,N_6758,N_7119);
nor U11645 (N_11645,N_6930,N_9001);
or U11646 (N_11646,N_6686,N_5079);
nor U11647 (N_11647,N_7223,N_5746);
or U11648 (N_11648,N_8281,N_6339);
nor U11649 (N_11649,N_5088,N_8716);
nand U11650 (N_11650,N_8435,N_6447);
and U11651 (N_11651,N_7829,N_7340);
nand U11652 (N_11652,N_7763,N_9522);
or U11653 (N_11653,N_6128,N_5864);
and U11654 (N_11654,N_8109,N_5117);
nor U11655 (N_11655,N_5577,N_6799);
or U11656 (N_11656,N_6830,N_6743);
nand U11657 (N_11657,N_7083,N_9214);
nor U11658 (N_11658,N_6108,N_5470);
and U11659 (N_11659,N_9695,N_8330);
or U11660 (N_11660,N_6449,N_5791);
xnor U11661 (N_11661,N_5986,N_5972);
or U11662 (N_11662,N_9873,N_6064);
nand U11663 (N_11663,N_5344,N_9514);
nor U11664 (N_11664,N_9020,N_9265);
xor U11665 (N_11665,N_7169,N_9646);
xor U11666 (N_11666,N_8083,N_8776);
or U11667 (N_11667,N_6107,N_7758);
and U11668 (N_11668,N_5955,N_8734);
nor U11669 (N_11669,N_8089,N_9386);
nor U11670 (N_11670,N_9609,N_9205);
xnor U11671 (N_11671,N_7616,N_5699);
and U11672 (N_11672,N_8510,N_9919);
xnor U11673 (N_11673,N_5240,N_9852);
or U11674 (N_11674,N_9408,N_6983);
and U11675 (N_11675,N_7861,N_5161);
xor U11676 (N_11676,N_6412,N_9979);
or U11677 (N_11677,N_5395,N_5160);
nor U11678 (N_11678,N_5361,N_9507);
nor U11679 (N_11679,N_9240,N_6253);
or U11680 (N_11680,N_8038,N_6278);
nand U11681 (N_11681,N_8393,N_7179);
xnor U11682 (N_11682,N_9198,N_6331);
or U11683 (N_11683,N_8331,N_5546);
xor U11684 (N_11684,N_6731,N_6918);
and U11685 (N_11685,N_8566,N_6017);
or U11686 (N_11686,N_7699,N_8681);
or U11687 (N_11687,N_7637,N_5683);
nand U11688 (N_11688,N_9462,N_8617);
xnor U11689 (N_11689,N_9759,N_5403);
nand U11690 (N_11690,N_7046,N_6303);
xor U11691 (N_11691,N_9542,N_6546);
nor U11692 (N_11692,N_9237,N_7972);
nor U11693 (N_11693,N_7675,N_8755);
nor U11694 (N_11694,N_9984,N_8353);
xor U11695 (N_11695,N_5508,N_9848);
nor U11696 (N_11696,N_8436,N_9648);
and U11697 (N_11697,N_7933,N_6771);
or U11698 (N_11698,N_7295,N_6052);
and U11699 (N_11699,N_5371,N_5071);
nor U11700 (N_11700,N_8727,N_5464);
nor U11701 (N_11701,N_5874,N_8174);
nand U11702 (N_11702,N_9788,N_7247);
or U11703 (N_11703,N_8099,N_8290);
and U11704 (N_11704,N_9463,N_9798);
xor U11705 (N_11705,N_9350,N_9376);
or U11706 (N_11706,N_7804,N_5213);
and U11707 (N_11707,N_8612,N_9103);
and U11708 (N_11708,N_5946,N_7605);
nor U11709 (N_11709,N_5402,N_8336);
xor U11710 (N_11710,N_9248,N_9288);
nor U11711 (N_11711,N_5383,N_8549);
nand U11712 (N_11712,N_9512,N_7025);
nor U11713 (N_11713,N_7339,N_7368);
and U11714 (N_11714,N_8178,N_8635);
nor U11715 (N_11715,N_7411,N_6246);
or U11716 (N_11716,N_5584,N_6901);
or U11717 (N_11717,N_8325,N_7952);
and U11718 (N_11718,N_7174,N_8307);
or U11719 (N_11719,N_9665,N_6598);
xor U11720 (N_11720,N_5163,N_6880);
nor U11721 (N_11721,N_8682,N_6072);
and U11722 (N_11722,N_7980,N_7427);
or U11723 (N_11723,N_9961,N_6347);
nor U11724 (N_11724,N_8158,N_7790);
nand U11725 (N_11725,N_9926,N_8337);
nor U11726 (N_11726,N_9671,N_8382);
and U11727 (N_11727,N_6163,N_8243);
or U11728 (N_11728,N_8479,N_9887);
or U11729 (N_11729,N_5065,N_6142);
xnor U11730 (N_11730,N_8841,N_7808);
and U11731 (N_11731,N_6419,N_8530);
or U11732 (N_11732,N_8912,N_5147);
nand U11733 (N_11733,N_9217,N_8421);
nor U11734 (N_11734,N_9118,N_9375);
nand U11735 (N_11735,N_5830,N_5701);
nand U11736 (N_11736,N_6825,N_6343);
xor U11737 (N_11737,N_8124,N_8931);
or U11738 (N_11738,N_5225,N_5890);
nor U11739 (N_11739,N_6795,N_7614);
nand U11740 (N_11740,N_7006,N_7863);
nand U11741 (N_11741,N_8609,N_9691);
xnor U11742 (N_11742,N_8870,N_5523);
or U11743 (N_11743,N_9546,N_6418);
xor U11744 (N_11744,N_8033,N_7521);
or U11745 (N_11745,N_5945,N_9945);
or U11746 (N_11746,N_8917,N_6969);
or U11747 (N_11747,N_5968,N_5816);
xnor U11748 (N_11748,N_7586,N_7695);
or U11749 (N_11749,N_6337,N_9568);
xnor U11750 (N_11750,N_5509,N_9520);
nor U11751 (N_11751,N_6735,N_7638);
nand U11752 (N_11752,N_9204,N_9009);
nand U11753 (N_11753,N_9161,N_5555);
or U11754 (N_11754,N_6851,N_6020);
or U11755 (N_11755,N_5333,N_6959);
or U11756 (N_11756,N_9521,N_8793);
and U11757 (N_11757,N_6756,N_6858);
and U11758 (N_11758,N_7386,N_8832);
nand U11759 (N_11759,N_7966,N_5475);
or U11760 (N_11760,N_9347,N_7356);
or U11761 (N_11761,N_5478,N_5979);
nand U11762 (N_11762,N_5860,N_7670);
or U11763 (N_11763,N_7115,N_8724);
nor U11764 (N_11764,N_7096,N_6836);
nand U11765 (N_11765,N_7085,N_8459);
nor U11766 (N_11766,N_6904,N_9183);
or U11767 (N_11767,N_5166,N_8165);
xor U11768 (N_11768,N_7281,N_7200);
and U11769 (N_11769,N_9036,N_7785);
or U11770 (N_11770,N_9340,N_8741);
nand U11771 (N_11771,N_9029,N_5717);
or U11772 (N_11772,N_9974,N_5024);
xor U11773 (N_11773,N_7469,N_9930);
and U11774 (N_11774,N_7278,N_9878);
nor U11775 (N_11775,N_8744,N_5971);
xor U11776 (N_11776,N_7087,N_5131);
xnor U11777 (N_11777,N_7049,N_8780);
nor U11778 (N_11778,N_8373,N_8280);
and U11779 (N_11779,N_5942,N_6451);
or U11780 (N_11780,N_7258,N_6896);
and U11781 (N_11781,N_7226,N_8072);
and U11782 (N_11782,N_5687,N_7849);
xnor U11783 (N_11783,N_6701,N_8922);
nor U11784 (N_11784,N_5591,N_5286);
nand U11785 (N_11785,N_5922,N_8031);
nand U11786 (N_11786,N_8391,N_8519);
nand U11787 (N_11787,N_8641,N_8560);
xnor U11788 (N_11788,N_6157,N_8453);
nand U11789 (N_11789,N_6425,N_9531);
and U11790 (N_11790,N_6805,N_7498);
nand U11791 (N_11791,N_7453,N_6965);
nand U11792 (N_11792,N_5020,N_5935);
xor U11793 (N_11793,N_6939,N_9163);
nor U11794 (N_11794,N_9793,N_9502);
xor U11795 (N_11795,N_9114,N_5114);
nor U11796 (N_11796,N_9950,N_5272);
or U11797 (N_11797,N_7978,N_7277);
nor U11798 (N_11798,N_9053,N_8196);
and U11799 (N_11799,N_9057,N_6912);
nand U11800 (N_11800,N_7218,N_6297);
and U11801 (N_11801,N_6798,N_9729);
xor U11802 (N_11802,N_6481,N_8737);
or U11803 (N_11803,N_7319,N_8390);
or U11804 (N_11804,N_9271,N_7419);
and U11805 (N_11805,N_7721,N_8013);
or U11806 (N_11806,N_9087,N_5993);
xnor U11807 (N_11807,N_6453,N_7198);
nor U11808 (N_11808,N_5146,N_7554);
or U11809 (N_11809,N_5035,N_5294);
xnor U11810 (N_11810,N_7551,N_9492);
nand U11811 (N_11811,N_8712,N_9802);
nand U11812 (N_11812,N_8717,N_8650);
or U11813 (N_11813,N_5851,N_8522);
nor U11814 (N_11814,N_7726,N_9741);
nand U11815 (N_11815,N_7283,N_9652);
or U11816 (N_11816,N_7507,N_8416);
or U11817 (N_11817,N_7818,N_6416);
nand U11818 (N_11818,N_6768,N_6161);
nor U11819 (N_11819,N_9421,N_5461);
or U11820 (N_11820,N_6008,N_7613);
and U11821 (N_11821,N_6697,N_8272);
nand U11822 (N_11822,N_5965,N_6929);
and U11823 (N_11823,N_5505,N_8871);
and U11824 (N_11824,N_9095,N_9965);
and U11825 (N_11825,N_8516,N_5425);
nor U11826 (N_11826,N_9563,N_7092);
and U11827 (N_11827,N_7299,N_8691);
or U11828 (N_11828,N_7363,N_8976);
and U11829 (N_11829,N_6850,N_5960);
nor U11830 (N_11830,N_5636,N_8911);
and U11831 (N_11831,N_6098,N_8006);
or U11832 (N_11832,N_5327,N_5090);
or U11833 (N_11833,N_6637,N_5516);
or U11834 (N_11834,N_6126,N_6149);
xor U11835 (N_11835,N_5512,N_7690);
xnor U11836 (N_11836,N_6791,N_6341);
nand U11837 (N_11837,N_7518,N_7279);
and U11838 (N_11838,N_9517,N_9796);
and U11839 (N_11839,N_8181,N_8619);
nand U11840 (N_11840,N_9613,N_9188);
nand U11841 (N_11841,N_7807,N_8910);
nand U11842 (N_11842,N_9737,N_7759);
nor U11843 (N_11843,N_8448,N_6981);
xor U11844 (N_11844,N_8966,N_7532);
nor U11845 (N_11845,N_8753,N_9809);
nor U11846 (N_11846,N_7924,N_8015);
xnor U11847 (N_11847,N_6765,N_6935);
and U11848 (N_11848,N_7408,N_5447);
and U11849 (N_11849,N_6669,N_9890);
nor U11850 (N_11850,N_7935,N_7712);
and U11851 (N_11851,N_8667,N_8889);
nor U11852 (N_11852,N_8525,N_5882);
and U11853 (N_11853,N_8389,N_9012);
nand U11854 (N_11854,N_6490,N_6540);
nor U11855 (N_11855,N_9643,N_6774);
nor U11856 (N_11856,N_5753,N_7701);
nor U11857 (N_11857,N_9355,N_7450);
and U11858 (N_11858,N_9816,N_7589);
nor U11859 (N_11859,N_8942,N_5677);
nor U11860 (N_11860,N_8051,N_6027);
or U11861 (N_11861,N_9394,N_7047);
and U11862 (N_11862,N_6612,N_5686);
nor U11863 (N_11863,N_7128,N_8591);
nor U11864 (N_11864,N_5000,N_7929);
nor U11865 (N_11865,N_7619,N_6106);
and U11866 (N_11866,N_7587,N_9966);
and U11867 (N_11867,N_7031,N_5103);
or U11868 (N_11868,N_6169,N_6477);
or U11869 (N_11869,N_8137,N_6961);
xor U11870 (N_11870,N_5936,N_7222);
and U11871 (N_11871,N_5798,N_9352);
nor U11872 (N_11872,N_8202,N_5387);
nor U11873 (N_11873,N_8014,N_9861);
nand U11874 (N_11874,N_9870,N_6968);
or U11875 (N_11875,N_6706,N_8247);
nand U11876 (N_11876,N_7593,N_8145);
xor U11877 (N_11877,N_9483,N_7187);
xnor U11878 (N_11878,N_5305,N_8546);
xnor U11879 (N_11879,N_6636,N_8050);
and U11880 (N_11880,N_8227,N_9558);
and U11881 (N_11881,N_7067,N_7567);
xor U11882 (N_11882,N_5142,N_8699);
nor U11883 (N_11883,N_6330,N_6531);
nand U11884 (N_11884,N_8814,N_7869);
and U11885 (N_11885,N_9555,N_9725);
and U11886 (N_11886,N_8141,N_6987);
and U11887 (N_11887,N_7366,N_8447);
or U11888 (N_11888,N_6063,N_5118);
and U11889 (N_11889,N_8792,N_7013);
xnor U11890 (N_11890,N_8508,N_5083);
or U11891 (N_11891,N_8645,N_9561);
xnor U11892 (N_11892,N_5069,N_8414);
nor U11893 (N_11893,N_5656,N_7506);
nor U11894 (N_11894,N_8908,N_5075);
nor U11895 (N_11895,N_6021,N_6841);
nor U11896 (N_11896,N_6988,N_8800);
or U11897 (N_11897,N_7266,N_5785);
nor U11898 (N_11898,N_5267,N_5916);
nor U11899 (N_11899,N_6882,N_5207);
nor U11900 (N_11900,N_8404,N_7812);
or U11901 (N_11901,N_6322,N_9983);
nand U11902 (N_11902,N_5041,N_9084);
and U11903 (N_11903,N_5422,N_8252);
xnor U11904 (N_11904,N_8312,N_5541);
nand U11905 (N_11905,N_8078,N_5540);
nor U11906 (N_11906,N_5289,N_8991);
nor U11907 (N_11907,N_9351,N_8157);
and U11908 (N_11908,N_9867,N_6677);
nor U11909 (N_11909,N_7385,N_9144);
nor U11910 (N_11910,N_6130,N_8935);
or U11911 (N_11911,N_8994,N_9642);
nor U11912 (N_11912,N_9362,N_7901);
nor U11913 (N_11913,N_5900,N_6654);
nand U11914 (N_11914,N_5689,N_9677);
nand U11915 (N_11915,N_9004,N_9192);
or U11916 (N_11916,N_9455,N_6621);
and U11917 (N_11917,N_8512,N_9692);
and U11918 (N_11918,N_9074,N_5222);
nor U11919 (N_11919,N_6514,N_6276);
and U11920 (N_11920,N_7584,N_9779);
xnor U11921 (N_11921,N_9996,N_9840);
nand U11922 (N_11922,N_7108,N_8759);
xnor U11923 (N_11923,N_9745,N_9778);
xnor U11924 (N_11924,N_8578,N_7844);
nand U11925 (N_11925,N_5058,N_5563);
xnor U11926 (N_11926,N_9055,N_7960);
xnor U11927 (N_11927,N_9556,N_5996);
or U11928 (N_11928,N_5319,N_9426);
and U11929 (N_11929,N_7905,N_7012);
and U11930 (N_11930,N_9152,N_6606);
and U11931 (N_11931,N_6160,N_6973);
nand U11932 (N_11932,N_7230,N_7235);
nand U11933 (N_11933,N_5659,N_8562);
xor U11934 (N_11934,N_8909,N_7754);
or U11935 (N_11935,N_6503,N_9303);
xnor U11936 (N_11936,N_5409,N_6295);
nand U11937 (N_11937,N_5763,N_8914);
and U11938 (N_11938,N_8901,N_8146);
and U11939 (N_11939,N_5148,N_9286);
xor U11940 (N_11940,N_9246,N_9300);
nand U11941 (N_11941,N_7603,N_8385);
or U11942 (N_11942,N_7403,N_7118);
or U11943 (N_11943,N_6437,N_8302);
or U11944 (N_11944,N_8999,N_5605);
xnor U11945 (N_11945,N_8879,N_6820);
or U11946 (N_11946,N_9393,N_5262);
xor U11947 (N_11947,N_9047,N_8979);
nor U11948 (N_11948,N_8169,N_8648);
xnor U11949 (N_11949,N_9696,N_5188);
and U11950 (N_11950,N_5042,N_7284);
and U11951 (N_11951,N_8219,N_9808);
or U11952 (N_11952,N_7436,N_7984);
xnor U11953 (N_11953,N_5938,N_8044);
nor U11954 (N_11954,N_7182,N_5040);
nor U11955 (N_11955,N_7107,N_7154);
or U11956 (N_11956,N_5757,N_5824);
and U11957 (N_11957,N_5903,N_9242);
xnor U11958 (N_11958,N_9086,N_7752);
xor U11959 (N_11959,N_5759,N_7660);
and U11960 (N_11960,N_6435,N_9610);
xnor U11961 (N_11961,N_9656,N_6552);
and U11962 (N_11962,N_9328,N_7451);
nor U11963 (N_11963,N_5536,N_7687);
nand U11964 (N_11964,N_6283,N_9157);
xnor U11965 (N_11965,N_8048,N_9633);
or U11966 (N_11966,N_8821,N_7099);
nor U11967 (N_11967,N_8846,N_5909);
xor U11968 (N_11968,N_6761,N_6903);
or U11969 (N_11969,N_7773,N_8017);
or U11970 (N_11970,N_6002,N_6625);
and U11971 (N_11971,N_9766,N_7373);
nor U11972 (N_11972,N_8689,N_8228);
nand U11973 (N_11973,N_9720,N_6277);
or U11974 (N_11974,N_7089,N_7927);
or U11975 (N_11975,N_5576,N_7535);
nand U11976 (N_11976,N_6776,N_8403);
or U11977 (N_11977,N_5839,N_8675);
nand U11978 (N_11978,N_8652,N_9672);
or U11979 (N_11979,N_9916,N_9775);
nand U11980 (N_11980,N_9039,N_5081);
xor U11981 (N_11981,N_6670,N_6494);
and U11982 (N_11982,N_7606,N_8555);
nor U11983 (N_11983,N_9379,N_9112);
xnor U11984 (N_11984,N_6714,N_6293);
or U11985 (N_11985,N_7003,N_7160);
nor U11986 (N_11986,N_7526,N_8248);
xor U11987 (N_11987,N_7264,N_6187);
nand U11988 (N_11988,N_9244,N_5062);
or U11989 (N_11989,N_8973,N_7454);
xnor U11990 (N_11990,N_5487,N_6972);
or U11991 (N_11991,N_6689,N_8601);
or U11992 (N_11992,N_7655,N_9135);
and U11993 (N_11993,N_9493,N_9236);
or U11994 (N_11994,N_5486,N_6238);
nor U11995 (N_11995,N_7954,N_9312);
xnor U11996 (N_11996,N_9506,N_8255);
nor U11997 (N_11997,N_8665,N_7908);
nand U11998 (N_11998,N_8206,N_5201);
nand U11999 (N_11999,N_5177,N_7253);
and U12000 (N_12000,N_8748,N_7746);
nor U12001 (N_12001,N_7561,N_9132);
nand U12002 (N_12002,N_9694,N_7872);
nand U12003 (N_12003,N_9172,N_5559);
or U12004 (N_12004,N_7513,N_6986);
or U12005 (N_12005,N_7794,N_9762);
and U12006 (N_12006,N_9539,N_6491);
and U12007 (N_12007,N_8020,N_5502);
or U12008 (N_12008,N_5254,N_5724);
nor U12009 (N_12009,N_5317,N_5316);
and U12010 (N_12010,N_6471,N_7648);
and U12011 (N_12011,N_7896,N_8820);
xnor U12012 (N_12012,N_5218,N_9989);
and U12013 (N_12013,N_7297,N_9337);
xnor U12014 (N_12014,N_5023,N_8497);
nand U12015 (N_12015,N_9255,N_6902);
and U12016 (N_12016,N_8053,N_6034);
or U12017 (N_12017,N_6992,N_8980);
and U12018 (N_12018,N_8278,N_9574);
and U12019 (N_12019,N_8957,N_9864);
xnor U12020 (N_12020,N_6441,N_5116);
xnor U12021 (N_12021,N_6736,N_8172);
xor U12022 (N_12022,N_5238,N_8182);
or U12023 (N_12023,N_7252,N_5694);
and U12024 (N_12024,N_6566,N_8511);
xor U12025 (N_12025,N_5012,N_5362);
or U12026 (N_12026,N_6561,N_7379);
xnor U12027 (N_12027,N_6960,N_6148);
nand U12028 (N_12028,N_7989,N_5795);
nor U12029 (N_12029,N_6564,N_6865);
and U12030 (N_12030,N_9076,N_7815);
and U12031 (N_12031,N_9068,N_8556);
and U12032 (N_12032,N_6724,N_6342);
xnor U12033 (N_12033,N_7084,N_6619);
or U12034 (N_12034,N_7364,N_5091);
or U12035 (N_12035,N_8663,N_8501);
nand U12036 (N_12036,N_9900,N_9739);
or U12037 (N_12037,N_8869,N_6110);
and U12038 (N_12038,N_6051,N_5925);
or U12039 (N_12039,N_9533,N_7318);
nor U12040 (N_12040,N_5649,N_5143);
xor U12041 (N_12041,N_5152,N_6003);
or U12042 (N_12042,N_6869,N_7134);
nor U12043 (N_12043,N_5941,N_8987);
or U12044 (N_12044,N_6073,N_6789);
nand U12045 (N_12045,N_7971,N_5805);
nor U12046 (N_12046,N_8628,N_5359);
nor U12047 (N_12047,N_7396,N_9804);
xnor U12048 (N_12048,N_7375,N_8465);
and U12049 (N_12049,N_6924,N_8019);
and U12050 (N_12050,N_5477,N_7945);
or U12051 (N_12051,N_8995,N_5351);
nor U12052 (N_12052,N_9256,N_8762);
xor U12053 (N_12053,N_9523,N_8711);
nor U12054 (N_12054,N_7678,N_8489);
or U12055 (N_12055,N_5175,N_6687);
xnor U12056 (N_12056,N_6505,N_6386);
xor U12057 (N_12057,N_7028,N_6354);
and U12058 (N_12058,N_6387,N_8466);
nand U12059 (N_12059,N_8432,N_8891);
nand U12060 (N_12060,N_6454,N_7688);
and U12061 (N_12061,N_9515,N_8538);
nor U12062 (N_12062,N_8813,N_5914);
nand U12063 (N_12063,N_7875,N_8311);
and U12064 (N_12064,N_5084,N_8110);
nand U12065 (N_12065,N_7335,N_8430);
nand U12066 (N_12066,N_8200,N_5440);
or U12067 (N_12067,N_9789,N_9578);
nor U12068 (N_12068,N_8627,N_7502);
and U12069 (N_12069,N_7382,N_9014);
nand U12070 (N_12070,N_6411,N_5149);
xor U12071 (N_12071,N_8625,N_7738);
and U12072 (N_12072,N_7983,N_6442);
nor U12073 (N_12073,N_9485,N_7388);
and U12074 (N_12074,N_6369,N_9764);
nor U12075 (N_12075,N_9360,N_8074);
and U12076 (N_12076,N_6786,N_9133);
xnor U12077 (N_12077,N_6879,N_7410);
nand U12078 (N_12078,N_8460,N_8769);
nor U12079 (N_12079,N_7541,N_6985);
nand U12080 (N_12080,N_6309,N_8328);
xnor U12081 (N_12081,N_7784,N_8486);
xnor U12082 (N_12082,N_6648,N_8961);
nor U12083 (N_12083,N_7048,N_6713);
or U12084 (N_12084,N_6688,N_9784);
nor U12085 (N_12085,N_9156,N_7140);
and U12086 (N_12086,N_5962,N_8924);
and U12087 (N_12087,N_8878,N_6947);
nand U12088 (N_12088,N_6536,N_7575);
nand U12089 (N_12089,N_6004,N_8386);
or U12090 (N_12090,N_9395,N_9346);
or U12091 (N_12091,N_9311,N_8674);
xnor U12092 (N_12092,N_7122,N_8789);
or U12093 (N_12093,N_9856,N_7213);
nand U12094 (N_12094,N_9356,N_5064);
xor U12095 (N_12095,N_8903,N_8399);
xnor U12096 (N_12096,N_7039,N_5283);
nand U12097 (N_12097,N_9208,N_8529);
or U12098 (N_12098,N_7761,N_8170);
nand U12099 (N_12099,N_6165,N_8283);
and U12100 (N_12100,N_7976,N_7941);
and U12101 (N_12101,N_7508,N_8299);
nand U12102 (N_12102,N_8524,N_6247);
xnor U12103 (N_12103,N_6640,N_5556);
nand U12104 (N_12104,N_5530,N_7838);
nand U12105 (N_12105,N_9373,N_5281);
and U12106 (N_12106,N_7756,N_5629);
nor U12107 (N_12107,N_9041,N_7833);
and U12108 (N_12108,N_5745,N_9605);
nor U12109 (N_12109,N_5571,N_6483);
nor U12110 (N_12110,N_7970,N_5921);
xnor U12111 (N_12111,N_6323,N_8314);
nand U12112 (N_12112,N_8482,N_9382);
or U12113 (N_12113,N_5010,N_9763);
nor U12114 (N_12114,N_5674,N_7691);
nand U12115 (N_12115,N_5583,N_9439);
nor U12116 (N_12116,N_6770,N_9220);
nand U12117 (N_12117,N_7202,N_6056);
or U12118 (N_12118,N_6887,N_8214);
nand U12119 (N_12119,N_8634,N_5522);
nand U12120 (N_12120,N_5122,N_9626);
or U12121 (N_12121,N_8040,N_5834);
nand U12122 (N_12122,N_5050,N_5808);
nor U12123 (N_12123,N_9434,N_7348);
xnor U12124 (N_12124,N_8001,N_6373);
xor U12125 (N_12125,N_6385,N_7592);
nand U12126 (N_12126,N_7276,N_6881);
nand U12127 (N_12127,N_8231,N_9117);
nand U12128 (N_12128,N_9669,N_5299);
and U12129 (N_12129,N_6267,N_5730);
xor U12130 (N_12130,N_6414,N_9639);
and U12131 (N_12131,N_6895,N_8499);
nand U12132 (N_12132,N_8662,N_7860);
nand U12133 (N_12133,N_6695,N_8589);
or U12134 (N_12134,N_5585,N_6205);
xor U12135 (N_12135,N_5197,N_5809);
nor U12136 (N_12136,N_7661,N_8630);
nand U12137 (N_12137,N_6080,N_7303);
xor U12138 (N_12138,N_8073,N_8455);
xor U12139 (N_12139,N_5545,N_8361);
and U12140 (N_12140,N_5375,N_5906);
or U12141 (N_12141,N_7780,N_8604);
or U12142 (N_12142,N_7846,N_6668);
nand U12143 (N_12143,N_6650,N_7827);
xor U12144 (N_12144,N_9511,N_6778);
and U12145 (N_12145,N_7280,N_5153);
and U12146 (N_12146,N_8678,N_5002);
nand U12147 (N_12147,N_8967,N_8406);
or U12148 (N_12148,N_5168,N_5532);
xor U12149 (N_12149,N_9089,N_8859);
nor U12150 (N_12150,N_7653,N_9284);
xnor U12151 (N_12151,N_6464,N_7914);
nand U12152 (N_12152,N_7684,N_9886);
and U12153 (N_12153,N_8921,N_6684);
or U12154 (N_12154,N_6443,N_6046);
nor U12155 (N_12155,N_7798,N_7415);
nor U12156 (N_12156,N_5312,N_9896);
nor U12157 (N_12157,N_8805,N_8669);
xor U12158 (N_12158,N_8250,N_5162);
nor U12159 (N_12159,N_7539,N_7822);
and U12160 (N_12160,N_9875,N_7962);
nor U12161 (N_12161,N_7101,N_8801);
nand U12162 (N_12162,N_8574,N_6845);
xnor U12163 (N_12163,N_8989,N_8087);
and U12164 (N_12164,N_7630,N_9540);
nor U12165 (N_12165,N_5726,N_8113);
or U12166 (N_12166,N_8034,N_8940);
or U12167 (N_12167,N_5544,N_9391);
nand U12168 (N_12168,N_7873,N_6162);
nand U12169 (N_12169,N_7636,N_5189);
or U12170 (N_12170,N_5495,N_7346);
xor U12171 (N_12171,N_9769,N_7098);
nand U12172 (N_12172,N_6685,N_7094);
and U12173 (N_12173,N_5382,N_6448);
and U12174 (N_12174,N_9712,N_9902);
xor U12175 (N_12175,N_7161,N_6817);
and U12176 (N_12176,N_6140,N_6316);
or U12177 (N_12177,N_8968,N_6777);
nor U12178 (N_12178,N_6649,N_5777);
nor U12179 (N_12179,N_8573,N_7462);
or U12180 (N_12180,N_5456,N_7850);
or U12181 (N_12181,N_7968,N_8469);
nor U12182 (N_12182,N_5560,N_6862);
or U12183 (N_12183,N_6093,N_5549);
nand U12184 (N_12184,N_5778,N_7729);
nor U12185 (N_12185,N_8923,N_7529);
and U12186 (N_12186,N_9185,N_7994);
and U12187 (N_12187,N_7666,N_7249);
nand U12188 (N_12188,N_7110,N_9344);
nor U12189 (N_12189,N_8279,N_9383);
or U12190 (N_12190,N_7659,N_5039);
nand U12191 (N_12191,N_7910,N_6475);
or U12192 (N_12192,N_9716,N_8817);
and U12193 (N_12193,N_6075,N_6958);
and U12194 (N_12194,N_5671,N_5290);
nand U12195 (N_12195,N_8807,N_7950);
nor U12196 (N_12196,N_5266,N_8825);
and U12197 (N_12197,N_7569,N_6355);
nand U12198 (N_12198,N_5722,N_8585);
or U12199 (N_12199,N_9443,N_5994);
and U12200 (N_12200,N_6940,N_9179);
xnor U12201 (N_12201,N_5564,N_8396);
nor U12202 (N_12202,N_5051,N_9191);
and U12203 (N_12203,N_7345,N_6824);
xor U12204 (N_12204,N_5345,N_7674);
and U12205 (N_12205,N_8763,N_5702);
or U12206 (N_12206,N_7260,N_6263);
or U12207 (N_12207,N_7228,N_9349);
or U12208 (N_12208,N_8664,N_9781);
and U12209 (N_12209,N_6755,N_5992);
or U12210 (N_12210,N_6848,N_6074);
nor U12211 (N_12211,N_5957,N_8371);
or U12212 (N_12212,N_9825,N_7713);
or U12213 (N_12213,N_6207,N_8168);
xnor U12214 (N_12214,N_9467,N_5215);
xor U12215 (N_12215,N_6374,N_6884);
or U12216 (N_12216,N_8693,N_8046);
nor U12217 (N_12217,N_6133,N_5416);
xnor U12218 (N_12218,N_9964,N_6465);
nand U12219 (N_12219,N_8379,N_9899);
and U12220 (N_12220,N_6515,N_6538);
xnor U12221 (N_12221,N_6745,N_6849);
xnor U12222 (N_12222,N_6291,N_7769);
nand U12223 (N_12223,N_8324,N_6039);
and U12224 (N_12224,N_8144,N_6856);
or U12225 (N_12225,N_5976,N_5881);
nor U12226 (N_12226,N_5622,N_9090);
xor U12227 (N_12227,N_8943,N_8898);
xnor U12228 (N_12228,N_7696,N_8528);
nand U12229 (N_12229,N_7809,N_9690);
xnor U12230 (N_12230,N_8354,N_6019);
nand U12231 (N_12231,N_6702,N_8209);
nand U12232 (N_12232,N_9401,N_6866);
and U12233 (N_12233,N_8673,N_5586);
and U12234 (N_12234,N_5608,N_5280);
or U12235 (N_12235,N_8842,N_8117);
xor U12236 (N_12236,N_7236,N_8192);
xor U12237 (N_12237,N_9107,N_5490);
xor U12238 (N_12238,N_5295,N_9892);
nor U12239 (N_12239,N_5076,N_5665);
or U12240 (N_12240,N_7312,N_6317);
or U12241 (N_12241,N_5731,N_5099);
xor U12242 (N_12242,N_6077,N_8694);
or U12243 (N_12243,N_9785,N_9321);
nand U12244 (N_12244,N_5256,N_5606);
and U12245 (N_12245,N_9201,N_9013);
nand U12246 (N_12246,N_8026,N_6274);
nor U12247 (N_12247,N_9817,N_5451);
nand U12248 (N_12248,N_7473,N_9827);
xor U12249 (N_12249,N_9150,N_9304);
nand U12250 (N_12250,N_5304,N_8543);
nand U12251 (N_12251,N_5494,N_9372);
nand U12252 (N_12252,N_7244,N_6938);
or U12253 (N_12253,N_7577,N_6048);
nor U12254 (N_12254,N_5872,N_8844);
nand U12255 (N_12255,N_9474,N_5087);
nor U12256 (N_12256,N_5484,N_6328);
nor U12257 (N_12257,N_5082,N_6616);
or U12258 (N_12258,N_5328,N_7316);
nand U12259 (N_12259,N_8104,N_5980);
nor U12260 (N_12260,N_6153,N_6524);
nand U12261 (N_12261,N_9675,N_7810);
nor U12262 (N_12262,N_7155,N_5533);
nand U12263 (N_12263,N_8707,N_6235);
xor U12264 (N_12264,N_7743,N_7767);
and U12265 (N_12265,N_5288,N_5005);
nor U12266 (N_12266,N_6104,N_6855);
nand U12267 (N_12267,N_6712,N_7062);
and U12268 (N_12268,N_6076,N_9477);
or U12269 (N_12269,N_5617,N_6497);
xor U12270 (N_12270,N_7250,N_9233);
xor U12271 (N_12271,N_5185,N_9309);
xnor U12272 (N_12272,N_7671,N_6480);
nand U12273 (N_12273,N_5782,N_6675);
nor U12274 (N_12274,N_8848,N_6086);
nor U12275 (N_12275,N_5931,N_5360);
or U12276 (N_12276,N_5105,N_5434);
or U12277 (N_12277,N_9052,N_9749);
xnor U12278 (N_12278,N_8866,N_6600);
xor U12279 (N_12279,N_9159,N_5307);
nor U12280 (N_12280,N_5136,N_7131);
or U12281 (N_12281,N_8242,N_9824);
nand U12282 (N_12282,N_7576,N_7491);
and U12283 (N_12283,N_8129,N_7964);
and U12284 (N_12284,N_5528,N_9637);
and U12285 (N_12285,N_9604,N_8857);
nand U12286 (N_12286,N_9999,N_8517);
nand U12287 (N_12287,N_5566,N_7369);
nand U12288 (N_12288,N_5853,N_9544);
nor U12289 (N_12289,N_8463,N_5614);
nor U12290 (N_12290,N_6501,N_5273);
and U12291 (N_12291,N_8523,N_6358);
nand U12292 (N_12292,N_7528,N_7876);
xnor U12293 (N_12293,N_7547,N_9276);
nor U12294 (N_12294,N_8407,N_8930);
or U12295 (N_12295,N_5204,N_6388);
xnor U12296 (N_12296,N_7184,N_9591);
nand U12297 (N_12297,N_7501,N_9589);
xor U12298 (N_12298,N_8102,N_6203);
nand U12299 (N_12299,N_9308,N_8095);
nor U12300 (N_12300,N_7654,N_6400);
or U12301 (N_12301,N_6710,N_9986);
xor U12302 (N_12302,N_9920,N_7370);
nor U12303 (N_12303,N_8791,N_8749);
or U12304 (N_12304,N_7963,N_7711);
nor U12305 (N_12305,N_7580,N_7650);
or U12306 (N_12306,N_6674,N_7656);
and U12307 (N_12307,N_8747,N_7698);
xnor U12308 (N_12308,N_8541,N_8624);
nand U12309 (N_12309,N_8798,N_8649);
or U12310 (N_12310,N_6980,N_9736);
nand U12311 (N_12311,N_8392,N_5589);
and U12312 (N_12312,N_6504,N_6305);
and U12313 (N_12313,N_7181,N_7004);
nand U12314 (N_12314,N_5427,N_6646);
nand U12315 (N_12315,N_7951,N_6113);
nand U12316 (N_12316,N_6446,N_8408);
nor U12317 (N_12317,N_8714,N_7395);
xnor U12318 (N_12318,N_9976,N_9723);
and U12319 (N_12319,N_6717,N_7357);
nand U12320 (N_12320,N_5567,N_5969);
nand U12321 (N_12321,N_9227,N_8550);
nand U12322 (N_12322,N_9098,N_6302);
xnor U12323 (N_12323,N_9740,N_5685);
and U12324 (N_12324,N_8111,N_8305);
nand U12325 (N_12325,N_6284,N_7302);
nand U12326 (N_12326,N_8425,N_7036);
and U12327 (N_12327,N_6611,N_6727);
and U12328 (N_12328,N_5953,N_6803);
and U12329 (N_12329,N_6739,N_6854);
nor U12330 (N_12330,N_8705,N_8012);
nor U12331 (N_12331,N_9174,N_7248);
nand U12332 (N_12332,N_5920,N_7930);
nor U12333 (N_12333,N_6922,N_7546);
and U12334 (N_12334,N_5529,N_8777);
xnor U12335 (N_12335,N_7999,N_8532);
xnor U12336 (N_12336,N_6486,N_6487);
xnor U12337 (N_12337,N_5156,N_8155);
nor U12338 (N_12338,N_6445,N_9162);
nand U12339 (N_12339,N_7902,N_7392);
xnor U12340 (N_12340,N_8686,N_7360);
nand U12341 (N_12341,N_7165,N_9018);
nand U12342 (N_12342,N_6898,N_8811);
and U12343 (N_12343,N_5278,N_9007);
nand U12344 (N_12344,N_5908,N_9727);
nand U12345 (N_12345,N_8929,N_7864);
xnor U12346 (N_12346,N_5471,N_9160);
and U12347 (N_12347,N_7621,N_6522);
nor U12348 (N_12348,N_9829,N_9049);
nand U12349 (N_12349,N_8907,N_8009);
and U12350 (N_12350,N_5961,N_9884);
xnor U12351 (N_12351,N_5985,N_9733);
nand U12352 (N_12352,N_7600,N_8027);
or U12353 (N_12353,N_5258,N_6249);
nor U12354 (N_12354,N_9773,N_5645);
xor U12355 (N_12355,N_6934,N_9850);
nor U12356 (N_12356,N_8000,N_9119);
nand U12357 (N_12357,N_7137,N_8350);
nand U12358 (N_12358,N_7588,N_8488);
and U12359 (N_12359,N_7399,N_6555);
xnor U12360 (N_12360,N_9306,N_8398);
xor U12361 (N_12361,N_6375,N_7243);
nor U12362 (N_12362,N_7400,N_8106);
nor U12363 (N_12363,N_6424,N_7406);
nor U12364 (N_12364,N_6664,N_8958);
nor U12365 (N_12365,N_6734,N_7114);
nor U12366 (N_12366,N_9011,N_6576);
nor U12367 (N_12367,N_7544,N_6430);
or U12368 (N_12368,N_9735,N_8271);
or U12369 (N_12369,N_6137,N_6852);
nor U12370 (N_12370,N_8542,N_9010);
and U12371 (N_12371,N_5513,N_8161);
or U12372 (N_12372,N_9971,N_7478);
xor U12373 (N_12373,N_5799,N_8895);
or U12374 (N_12374,N_7495,N_7947);
xnor U12375 (N_12375,N_8570,N_9228);
xor U12376 (N_12376,N_7313,N_7708);
xor U12377 (N_12377,N_6978,N_5663);
nor U12378 (N_12378,N_9147,N_5365);
nand U12379 (N_12379,N_8605,N_9110);
and U12380 (N_12380,N_7349,N_8670);
nand U12381 (N_12381,N_8005,N_9232);
nor U12382 (N_12382,N_5878,N_9195);
xnor U12383 (N_12383,N_7795,N_5561);
and U12384 (N_12384,N_7893,N_6893);
nand U12385 (N_12385,N_5967,N_9409);
and U12386 (N_12386,N_7071,N_6949);
or U12387 (N_12387,N_5542,N_5825);
xor U12388 (N_12388,N_5227,N_7216);
nand U12389 (N_12389,N_5401,N_8697);
xnor U12390 (N_12390,N_5473,N_8091);
or U12391 (N_12391,N_6971,N_6042);
nand U12392 (N_12392,N_9064,N_9472);
or U12393 (N_12393,N_5675,N_5888);
and U12394 (N_12394,N_6970,N_9423);
xnor U12395 (N_12395,N_7911,N_5271);
xor U12396 (N_12396,N_7667,N_9151);
nor U12397 (N_12397,N_6332,N_9289);
nor U12398 (N_12398,N_5430,N_7022);
or U12399 (N_12399,N_5562,N_6957);
nand U12400 (N_12400,N_5354,N_9770);
nand U12401 (N_12401,N_6050,N_6943);
or U12402 (N_12402,N_7144,N_8575);
nor U12403 (N_12403,N_9946,N_6214);
nand U12404 (N_12404,N_9791,N_9056);
nand U12405 (N_12405,N_8246,N_5891);
nand U12406 (N_12406,N_6427,N_9673);
xnor U12407 (N_12407,N_8590,N_9955);
nor U12408 (N_12408,N_6812,N_6245);
or U12409 (N_12409,N_6011,N_9935);
or U12410 (N_12410,N_9187,N_8028);
or U12411 (N_12411,N_5913,N_6171);
nor U12412 (N_12412,N_6368,N_6186);
nand U12413 (N_12413,N_7657,N_5436);
xnor U12414 (N_12414,N_7333,N_6028);
nor U12415 (N_12415,N_5721,N_8567);
xor U12416 (N_12416,N_7354,N_6775);
and U12417 (N_12417,N_9224,N_9230);
xor U12418 (N_12418,N_7464,N_5368);
xnor U12419 (N_12419,N_8845,N_6558);
nand U12420 (N_12420,N_8632,N_6103);
or U12421 (N_12421,N_6993,N_8676);
nand U12422 (N_12422,N_6533,N_8256);
or U12423 (N_12423,N_9617,N_9842);
xnor U12424 (N_12424,N_8616,N_8483);
nor U12425 (N_12425,N_6134,N_8865);
and U12426 (N_12426,N_9111,N_9880);
nor U12427 (N_12427,N_7986,N_7537);
and U12428 (N_12428,N_9081,N_5199);
xor U12429 (N_12429,N_5274,N_9611);
nor U12430 (N_12430,N_8835,N_8431);
nor U12431 (N_12431,N_6326,N_5467);
xor U12432 (N_12432,N_7259,N_9645);
and U12433 (N_12433,N_6728,N_8974);
nor U12434 (N_12434,N_6462,N_9045);
xnor U12435 (N_12435,N_9445,N_9305);
and U12436 (N_12436,N_6196,N_5095);
or U12437 (N_12437,N_7492,N_6395);
or U12438 (N_12438,N_7715,N_7771);
nor U12439 (N_12439,N_5612,N_5870);
nand U12440 (N_12440,N_5879,N_5604);
nand U12441 (N_12441,N_5089,N_9392);
xor U12442 (N_12442,N_9797,N_8004);
and U12443 (N_12443,N_8442,N_8568);
xnor U12444 (N_12444,N_6193,N_5626);
xor U12445 (N_12445,N_9622,N_7832);
nor U12446 (N_12446,N_6821,N_6112);
and U12447 (N_12447,N_9464,N_9354);
and U12448 (N_12448,N_5847,N_8975);
and U12449 (N_12449,N_8369,N_6638);
xor U12450 (N_12450,N_8963,N_6933);
nand U12451 (N_12451,N_5793,N_5819);
and U12452 (N_12452,N_6213,N_6946);
xnor U12453 (N_12453,N_7331,N_6966);
and U12454 (N_12454,N_7943,N_6763);
or U12455 (N_12455,N_7904,N_7851);
nand U12456 (N_12456,N_7088,N_7522);
xor U12457 (N_12457,N_8468,N_5995);
or U12458 (N_12458,N_7705,N_8258);
or U12459 (N_12459,N_7398,N_8668);
nand U12460 (N_12460,N_9138,N_8055);
or U12461 (N_12461,N_8367,N_7380);
and U12462 (N_12462,N_5553,N_7162);
or U12463 (N_12463,N_9213,N_9058);
and U12464 (N_12464,N_5519,N_7016);
nor U12465 (N_12465,N_7467,N_7143);
or U12466 (N_12466,N_7740,N_9175);
xor U12467 (N_12467,N_9169,N_7870);
nor U12468 (N_12468,N_6363,N_6124);
xor U12469 (N_12469,N_7111,N_8856);
or U12470 (N_12470,N_5999,N_6547);
nor U12471 (N_12471,N_5297,N_7895);
xnor U12472 (N_12472,N_9894,N_8933);
xnor U12473 (N_12473,N_6348,N_6272);
nand U12474 (N_12474,N_7461,N_8265);
xor U12475 (N_12475,N_7208,N_9189);
xnor U12476 (N_12476,N_5647,N_9343);
or U12477 (N_12477,N_6647,N_9142);
or U12478 (N_12478,N_7418,N_6937);
nand U12479 (N_12479,N_5055,N_5899);
or U12480 (N_12480,N_7330,N_5510);
nor U12481 (N_12481,N_9155,N_5423);
and U12482 (N_12482,N_9750,N_9167);
nor U12483 (N_12483,N_7201,N_5623);
nand U12484 (N_12484,N_6439,N_6804);
and U12485 (N_12485,N_9223,N_5682);
or U12486 (N_12486,N_8045,N_7026);
and U12487 (N_12487,N_9697,N_9536);
nand U12488 (N_12488,N_8484,N_9203);
and U12489 (N_12489,N_9129,N_7610);
or U12490 (N_12490,N_8384,N_9301);
nand U12491 (N_12491,N_5159,N_6159);
nor U12492 (N_12492,N_5537,N_9557);
nand U12493 (N_12493,N_9721,N_9830);
and U12494 (N_12494,N_8806,N_9683);
or U12495 (N_12495,N_6264,N_6310);
xnor U12496 (N_12496,N_8150,N_8260);
nor U12497 (N_12497,N_8070,N_6927);
nor U12498 (N_12498,N_6174,N_6058);
and U12499 (N_12499,N_6215,N_7777);
xor U12500 (N_12500,N_9268,N_8482);
xor U12501 (N_12501,N_9794,N_7240);
and U12502 (N_12502,N_6540,N_6246);
nand U12503 (N_12503,N_5322,N_8264);
and U12504 (N_12504,N_8826,N_5093);
or U12505 (N_12505,N_9351,N_5039);
and U12506 (N_12506,N_7360,N_5434);
or U12507 (N_12507,N_7100,N_7853);
nand U12508 (N_12508,N_6140,N_8065);
xor U12509 (N_12509,N_6392,N_5010);
nand U12510 (N_12510,N_6788,N_7567);
nor U12511 (N_12511,N_5431,N_5029);
and U12512 (N_12512,N_5395,N_7696);
nor U12513 (N_12513,N_9453,N_8538);
and U12514 (N_12514,N_8971,N_9066);
nor U12515 (N_12515,N_6015,N_6128);
and U12516 (N_12516,N_9547,N_6725);
xnor U12517 (N_12517,N_9580,N_5012);
xnor U12518 (N_12518,N_9487,N_6611);
nor U12519 (N_12519,N_8483,N_9720);
nand U12520 (N_12520,N_6790,N_9082);
nor U12521 (N_12521,N_8810,N_9240);
or U12522 (N_12522,N_8531,N_7304);
nor U12523 (N_12523,N_9281,N_9172);
and U12524 (N_12524,N_6230,N_7135);
nand U12525 (N_12525,N_8228,N_9323);
nand U12526 (N_12526,N_9993,N_5962);
nand U12527 (N_12527,N_6928,N_8418);
nand U12528 (N_12528,N_6011,N_7402);
nor U12529 (N_12529,N_9757,N_6812);
xor U12530 (N_12530,N_5703,N_9731);
or U12531 (N_12531,N_5929,N_8855);
nand U12532 (N_12532,N_7865,N_6571);
and U12533 (N_12533,N_9988,N_6389);
or U12534 (N_12534,N_9818,N_5102);
nor U12535 (N_12535,N_9145,N_5768);
or U12536 (N_12536,N_6506,N_8495);
and U12537 (N_12537,N_9111,N_5929);
nor U12538 (N_12538,N_8112,N_5762);
or U12539 (N_12539,N_8926,N_7135);
nor U12540 (N_12540,N_6786,N_7690);
nand U12541 (N_12541,N_6568,N_9196);
nor U12542 (N_12542,N_6760,N_9313);
or U12543 (N_12543,N_9146,N_6958);
nand U12544 (N_12544,N_8915,N_8530);
xnor U12545 (N_12545,N_5789,N_9427);
nand U12546 (N_12546,N_6520,N_5136);
nor U12547 (N_12547,N_9666,N_6811);
and U12548 (N_12548,N_8388,N_7693);
or U12549 (N_12549,N_6135,N_8599);
xnor U12550 (N_12550,N_6110,N_8925);
xor U12551 (N_12551,N_6929,N_9536);
and U12552 (N_12552,N_6864,N_8399);
nor U12553 (N_12553,N_9001,N_8810);
or U12554 (N_12554,N_9132,N_9413);
or U12555 (N_12555,N_9381,N_6130);
xor U12556 (N_12556,N_5884,N_9693);
or U12557 (N_12557,N_5666,N_6592);
xor U12558 (N_12558,N_9780,N_6205);
nor U12559 (N_12559,N_7293,N_6904);
xor U12560 (N_12560,N_8690,N_7707);
nor U12561 (N_12561,N_5270,N_6527);
nor U12562 (N_12562,N_7515,N_8963);
xnor U12563 (N_12563,N_6232,N_9158);
or U12564 (N_12564,N_5822,N_6221);
xnor U12565 (N_12565,N_6674,N_9702);
xor U12566 (N_12566,N_6896,N_8015);
and U12567 (N_12567,N_6262,N_8833);
xor U12568 (N_12568,N_8826,N_5305);
nor U12569 (N_12569,N_8303,N_9093);
and U12570 (N_12570,N_9932,N_9208);
nand U12571 (N_12571,N_9837,N_7459);
nor U12572 (N_12572,N_9048,N_8904);
nand U12573 (N_12573,N_9848,N_6369);
or U12574 (N_12574,N_6434,N_5583);
or U12575 (N_12575,N_9887,N_5945);
nand U12576 (N_12576,N_6118,N_6372);
nand U12577 (N_12577,N_8146,N_7317);
xor U12578 (N_12578,N_8999,N_6714);
and U12579 (N_12579,N_8503,N_9535);
xor U12580 (N_12580,N_9318,N_5973);
nand U12581 (N_12581,N_6469,N_6685);
nand U12582 (N_12582,N_7892,N_8676);
nand U12583 (N_12583,N_9462,N_8781);
or U12584 (N_12584,N_5616,N_7683);
nor U12585 (N_12585,N_5470,N_5563);
xor U12586 (N_12586,N_8194,N_6927);
and U12587 (N_12587,N_7957,N_6565);
nand U12588 (N_12588,N_9601,N_7397);
or U12589 (N_12589,N_9374,N_7720);
xnor U12590 (N_12590,N_7578,N_6759);
and U12591 (N_12591,N_5266,N_5396);
xor U12592 (N_12592,N_9151,N_9485);
nand U12593 (N_12593,N_7902,N_6137);
and U12594 (N_12594,N_6888,N_7854);
nor U12595 (N_12595,N_7437,N_6810);
xor U12596 (N_12596,N_6111,N_9133);
or U12597 (N_12597,N_5177,N_6768);
or U12598 (N_12598,N_5946,N_8894);
nand U12599 (N_12599,N_9482,N_6510);
xor U12600 (N_12600,N_7332,N_7277);
nor U12601 (N_12601,N_9131,N_5370);
nor U12602 (N_12602,N_9342,N_7407);
nor U12603 (N_12603,N_9453,N_8400);
or U12604 (N_12604,N_7172,N_8677);
nand U12605 (N_12605,N_7707,N_6472);
xnor U12606 (N_12606,N_6799,N_5737);
or U12607 (N_12607,N_8051,N_7180);
and U12608 (N_12608,N_7475,N_9563);
and U12609 (N_12609,N_7607,N_7462);
or U12610 (N_12610,N_8826,N_6093);
nor U12611 (N_12611,N_9790,N_9885);
and U12612 (N_12612,N_7855,N_8986);
nor U12613 (N_12613,N_8385,N_5096);
or U12614 (N_12614,N_5585,N_9262);
and U12615 (N_12615,N_6847,N_7237);
nor U12616 (N_12616,N_7817,N_7579);
nor U12617 (N_12617,N_5282,N_9336);
nor U12618 (N_12618,N_8225,N_5543);
xnor U12619 (N_12619,N_6049,N_7834);
nor U12620 (N_12620,N_7284,N_8975);
or U12621 (N_12621,N_6319,N_8391);
nor U12622 (N_12622,N_6322,N_5775);
and U12623 (N_12623,N_9230,N_6942);
or U12624 (N_12624,N_8599,N_6673);
or U12625 (N_12625,N_5969,N_9400);
nand U12626 (N_12626,N_7102,N_9942);
xor U12627 (N_12627,N_5328,N_6818);
or U12628 (N_12628,N_8943,N_8475);
or U12629 (N_12629,N_8657,N_6848);
nand U12630 (N_12630,N_6197,N_8319);
nand U12631 (N_12631,N_7440,N_6843);
nor U12632 (N_12632,N_6036,N_9498);
or U12633 (N_12633,N_5291,N_5898);
and U12634 (N_12634,N_8821,N_5968);
nor U12635 (N_12635,N_8413,N_9131);
xnor U12636 (N_12636,N_8824,N_6296);
nand U12637 (N_12637,N_9200,N_8798);
xor U12638 (N_12638,N_7334,N_6025);
nand U12639 (N_12639,N_5592,N_6631);
nor U12640 (N_12640,N_5234,N_8814);
and U12641 (N_12641,N_8616,N_6389);
nand U12642 (N_12642,N_7495,N_8601);
nor U12643 (N_12643,N_6847,N_6987);
nand U12644 (N_12644,N_8046,N_6678);
or U12645 (N_12645,N_6208,N_6851);
xnor U12646 (N_12646,N_9400,N_9846);
or U12647 (N_12647,N_7804,N_6825);
xor U12648 (N_12648,N_8867,N_5001);
nand U12649 (N_12649,N_8742,N_8694);
nor U12650 (N_12650,N_5935,N_6423);
and U12651 (N_12651,N_5235,N_7125);
and U12652 (N_12652,N_7116,N_8912);
nor U12653 (N_12653,N_8265,N_6548);
and U12654 (N_12654,N_7058,N_5412);
nand U12655 (N_12655,N_5460,N_6670);
or U12656 (N_12656,N_8248,N_8363);
or U12657 (N_12657,N_7125,N_8494);
xnor U12658 (N_12658,N_7680,N_5359);
and U12659 (N_12659,N_6143,N_7438);
nand U12660 (N_12660,N_5605,N_8022);
and U12661 (N_12661,N_8056,N_9283);
or U12662 (N_12662,N_6244,N_8686);
nor U12663 (N_12663,N_5008,N_8145);
nor U12664 (N_12664,N_8412,N_9072);
xor U12665 (N_12665,N_8530,N_9771);
nand U12666 (N_12666,N_9425,N_9963);
xor U12667 (N_12667,N_7882,N_8285);
or U12668 (N_12668,N_9769,N_9287);
and U12669 (N_12669,N_9687,N_8130);
and U12670 (N_12670,N_5111,N_5537);
xor U12671 (N_12671,N_8424,N_6596);
nand U12672 (N_12672,N_6433,N_8207);
nor U12673 (N_12673,N_5816,N_6681);
and U12674 (N_12674,N_7706,N_6903);
or U12675 (N_12675,N_8586,N_5944);
nor U12676 (N_12676,N_5754,N_6351);
xor U12677 (N_12677,N_5808,N_5810);
nand U12678 (N_12678,N_5312,N_9484);
and U12679 (N_12679,N_9606,N_8063);
and U12680 (N_12680,N_8481,N_9588);
and U12681 (N_12681,N_5745,N_7671);
or U12682 (N_12682,N_9605,N_5349);
nor U12683 (N_12683,N_8226,N_5470);
nor U12684 (N_12684,N_7660,N_6530);
nand U12685 (N_12685,N_5442,N_5699);
nand U12686 (N_12686,N_8305,N_5847);
nor U12687 (N_12687,N_9518,N_5287);
nand U12688 (N_12688,N_6056,N_9939);
nand U12689 (N_12689,N_8425,N_7367);
or U12690 (N_12690,N_7832,N_6724);
and U12691 (N_12691,N_9601,N_5789);
and U12692 (N_12692,N_9049,N_7471);
xnor U12693 (N_12693,N_9499,N_8140);
or U12694 (N_12694,N_7639,N_9776);
or U12695 (N_12695,N_9116,N_6707);
xnor U12696 (N_12696,N_9508,N_6604);
nand U12697 (N_12697,N_9229,N_6599);
xnor U12698 (N_12698,N_9924,N_8366);
xnor U12699 (N_12699,N_5481,N_7608);
nand U12700 (N_12700,N_5855,N_7898);
nand U12701 (N_12701,N_9242,N_7302);
or U12702 (N_12702,N_9240,N_7824);
and U12703 (N_12703,N_8392,N_8030);
and U12704 (N_12704,N_9248,N_7450);
or U12705 (N_12705,N_6585,N_9988);
xnor U12706 (N_12706,N_5884,N_9870);
xor U12707 (N_12707,N_6624,N_6160);
nor U12708 (N_12708,N_9741,N_6282);
nor U12709 (N_12709,N_8575,N_6811);
and U12710 (N_12710,N_9392,N_9776);
nor U12711 (N_12711,N_5843,N_5972);
xor U12712 (N_12712,N_8559,N_6977);
xnor U12713 (N_12713,N_9507,N_7710);
xor U12714 (N_12714,N_6640,N_5352);
or U12715 (N_12715,N_7611,N_5046);
and U12716 (N_12716,N_7808,N_5816);
nor U12717 (N_12717,N_9172,N_8433);
and U12718 (N_12718,N_5343,N_6888);
nor U12719 (N_12719,N_8193,N_6808);
and U12720 (N_12720,N_5360,N_6377);
nor U12721 (N_12721,N_9652,N_6051);
nand U12722 (N_12722,N_6690,N_8278);
and U12723 (N_12723,N_5553,N_7965);
or U12724 (N_12724,N_7182,N_7191);
or U12725 (N_12725,N_9780,N_5509);
nand U12726 (N_12726,N_8807,N_5955);
nor U12727 (N_12727,N_6134,N_7887);
or U12728 (N_12728,N_6924,N_5659);
or U12729 (N_12729,N_8549,N_6846);
or U12730 (N_12730,N_9839,N_7901);
xnor U12731 (N_12731,N_5598,N_8525);
or U12732 (N_12732,N_7389,N_7968);
or U12733 (N_12733,N_6162,N_5337);
nand U12734 (N_12734,N_9996,N_6015);
and U12735 (N_12735,N_9036,N_8276);
nor U12736 (N_12736,N_6641,N_9398);
xnor U12737 (N_12737,N_6835,N_9260);
and U12738 (N_12738,N_8207,N_8159);
and U12739 (N_12739,N_6688,N_6239);
xor U12740 (N_12740,N_6710,N_6344);
nand U12741 (N_12741,N_9558,N_8969);
nor U12742 (N_12742,N_7394,N_5785);
xor U12743 (N_12743,N_7861,N_8354);
and U12744 (N_12744,N_8415,N_6993);
nand U12745 (N_12745,N_5192,N_7212);
and U12746 (N_12746,N_6050,N_6257);
and U12747 (N_12747,N_8449,N_5600);
xor U12748 (N_12748,N_7385,N_7927);
xnor U12749 (N_12749,N_7441,N_8889);
xor U12750 (N_12750,N_7986,N_8647);
xor U12751 (N_12751,N_8695,N_8737);
xor U12752 (N_12752,N_8163,N_8275);
or U12753 (N_12753,N_9202,N_6308);
or U12754 (N_12754,N_7611,N_7748);
or U12755 (N_12755,N_9022,N_7007);
xor U12756 (N_12756,N_6043,N_5933);
nand U12757 (N_12757,N_8040,N_6676);
and U12758 (N_12758,N_6200,N_8124);
and U12759 (N_12759,N_8268,N_7309);
nor U12760 (N_12760,N_7598,N_8749);
xor U12761 (N_12761,N_8383,N_7092);
nand U12762 (N_12762,N_5635,N_6590);
xnor U12763 (N_12763,N_9850,N_9073);
xor U12764 (N_12764,N_6680,N_9173);
and U12765 (N_12765,N_8343,N_8635);
and U12766 (N_12766,N_6217,N_5204);
or U12767 (N_12767,N_5906,N_6621);
and U12768 (N_12768,N_5317,N_9233);
nor U12769 (N_12769,N_7274,N_8195);
or U12770 (N_12770,N_5082,N_5539);
or U12771 (N_12771,N_6253,N_9005);
nand U12772 (N_12772,N_8438,N_5777);
nor U12773 (N_12773,N_5886,N_7778);
or U12774 (N_12774,N_9070,N_6381);
and U12775 (N_12775,N_8769,N_5199);
or U12776 (N_12776,N_6343,N_6966);
and U12777 (N_12777,N_7440,N_6001);
or U12778 (N_12778,N_9829,N_7367);
and U12779 (N_12779,N_6159,N_8883);
or U12780 (N_12780,N_9091,N_6128);
nor U12781 (N_12781,N_7478,N_6574);
and U12782 (N_12782,N_8910,N_5966);
and U12783 (N_12783,N_9114,N_7075);
nor U12784 (N_12784,N_9530,N_9465);
or U12785 (N_12785,N_6750,N_7770);
xor U12786 (N_12786,N_6735,N_9181);
or U12787 (N_12787,N_9004,N_5147);
nor U12788 (N_12788,N_5682,N_9170);
or U12789 (N_12789,N_8834,N_7350);
xnor U12790 (N_12790,N_5621,N_9939);
and U12791 (N_12791,N_5835,N_9640);
and U12792 (N_12792,N_7994,N_6859);
nor U12793 (N_12793,N_6407,N_8123);
xnor U12794 (N_12794,N_7347,N_6842);
nand U12795 (N_12795,N_6212,N_9449);
and U12796 (N_12796,N_8363,N_5472);
and U12797 (N_12797,N_8929,N_8684);
nand U12798 (N_12798,N_9120,N_8300);
nor U12799 (N_12799,N_7235,N_9496);
nand U12800 (N_12800,N_8851,N_6598);
xnor U12801 (N_12801,N_9277,N_5859);
or U12802 (N_12802,N_7154,N_6332);
nand U12803 (N_12803,N_8202,N_9122);
nand U12804 (N_12804,N_7737,N_8244);
xnor U12805 (N_12805,N_7122,N_6534);
nand U12806 (N_12806,N_5835,N_6031);
nand U12807 (N_12807,N_7421,N_9251);
and U12808 (N_12808,N_6755,N_6456);
nor U12809 (N_12809,N_6150,N_5938);
nor U12810 (N_12810,N_5544,N_9160);
nand U12811 (N_12811,N_9678,N_9478);
nor U12812 (N_12812,N_7183,N_8419);
nand U12813 (N_12813,N_6748,N_6674);
or U12814 (N_12814,N_8089,N_8337);
nor U12815 (N_12815,N_6258,N_7338);
or U12816 (N_12816,N_7320,N_6392);
or U12817 (N_12817,N_8176,N_9428);
nor U12818 (N_12818,N_6289,N_5774);
nor U12819 (N_12819,N_8217,N_7450);
and U12820 (N_12820,N_9315,N_6252);
or U12821 (N_12821,N_6600,N_8366);
nand U12822 (N_12822,N_8147,N_6814);
nand U12823 (N_12823,N_6115,N_5795);
nand U12824 (N_12824,N_7095,N_5868);
nor U12825 (N_12825,N_5188,N_6078);
nand U12826 (N_12826,N_6019,N_8696);
and U12827 (N_12827,N_9753,N_5178);
xnor U12828 (N_12828,N_7537,N_9836);
xnor U12829 (N_12829,N_6710,N_5165);
or U12830 (N_12830,N_5310,N_9892);
nand U12831 (N_12831,N_5602,N_7580);
xnor U12832 (N_12832,N_6988,N_7860);
nor U12833 (N_12833,N_8714,N_6255);
nor U12834 (N_12834,N_5869,N_5010);
or U12835 (N_12835,N_9280,N_8298);
or U12836 (N_12836,N_5943,N_9605);
nor U12837 (N_12837,N_9981,N_9385);
nor U12838 (N_12838,N_6682,N_7491);
and U12839 (N_12839,N_6347,N_8308);
or U12840 (N_12840,N_7931,N_5014);
xnor U12841 (N_12841,N_9748,N_7594);
nand U12842 (N_12842,N_6307,N_6527);
xor U12843 (N_12843,N_9913,N_8825);
xnor U12844 (N_12844,N_8935,N_7278);
or U12845 (N_12845,N_7512,N_5278);
nor U12846 (N_12846,N_7304,N_8376);
nand U12847 (N_12847,N_6943,N_9150);
xor U12848 (N_12848,N_8709,N_6204);
xor U12849 (N_12849,N_8583,N_9452);
nor U12850 (N_12850,N_5325,N_5405);
and U12851 (N_12851,N_9372,N_5741);
nand U12852 (N_12852,N_9920,N_8675);
and U12853 (N_12853,N_9304,N_9395);
nor U12854 (N_12854,N_9668,N_8580);
nor U12855 (N_12855,N_9006,N_7453);
nor U12856 (N_12856,N_7446,N_6829);
and U12857 (N_12857,N_8433,N_5643);
or U12858 (N_12858,N_9109,N_6741);
nand U12859 (N_12859,N_7334,N_6007);
or U12860 (N_12860,N_8724,N_6787);
or U12861 (N_12861,N_7986,N_8322);
or U12862 (N_12862,N_7393,N_8071);
or U12863 (N_12863,N_5922,N_6445);
nor U12864 (N_12864,N_9916,N_8462);
and U12865 (N_12865,N_7086,N_5433);
and U12866 (N_12866,N_8599,N_8930);
or U12867 (N_12867,N_9459,N_5505);
xor U12868 (N_12868,N_8010,N_5436);
nand U12869 (N_12869,N_9349,N_8834);
and U12870 (N_12870,N_7066,N_6052);
xnor U12871 (N_12871,N_9259,N_8685);
xor U12872 (N_12872,N_5989,N_7921);
xnor U12873 (N_12873,N_5062,N_9608);
nand U12874 (N_12874,N_8981,N_8379);
nor U12875 (N_12875,N_5384,N_6291);
or U12876 (N_12876,N_6268,N_9774);
nand U12877 (N_12877,N_7124,N_7259);
nor U12878 (N_12878,N_9213,N_6351);
or U12879 (N_12879,N_6778,N_8593);
or U12880 (N_12880,N_9719,N_9000);
and U12881 (N_12881,N_5770,N_6848);
or U12882 (N_12882,N_5564,N_9185);
nor U12883 (N_12883,N_7420,N_8991);
and U12884 (N_12884,N_9180,N_5038);
or U12885 (N_12885,N_7276,N_7252);
or U12886 (N_12886,N_9813,N_7565);
nand U12887 (N_12887,N_7588,N_6677);
nor U12888 (N_12888,N_9231,N_5258);
and U12889 (N_12889,N_9358,N_6843);
nor U12890 (N_12890,N_8627,N_6407);
and U12891 (N_12891,N_9544,N_5028);
or U12892 (N_12892,N_5516,N_9374);
nor U12893 (N_12893,N_8696,N_6749);
nand U12894 (N_12894,N_7200,N_5368);
nor U12895 (N_12895,N_9427,N_5361);
xnor U12896 (N_12896,N_8309,N_8170);
nand U12897 (N_12897,N_6303,N_6575);
nor U12898 (N_12898,N_8771,N_7565);
xor U12899 (N_12899,N_9713,N_5717);
nand U12900 (N_12900,N_7871,N_6782);
nor U12901 (N_12901,N_6998,N_5862);
xnor U12902 (N_12902,N_6742,N_8531);
nand U12903 (N_12903,N_5042,N_6505);
nor U12904 (N_12904,N_6370,N_6516);
and U12905 (N_12905,N_5411,N_7979);
or U12906 (N_12906,N_5205,N_9535);
nor U12907 (N_12907,N_7829,N_8039);
or U12908 (N_12908,N_5313,N_9996);
and U12909 (N_12909,N_5895,N_9206);
and U12910 (N_12910,N_7858,N_6965);
nor U12911 (N_12911,N_9796,N_8986);
nor U12912 (N_12912,N_7707,N_7718);
nor U12913 (N_12913,N_6777,N_6673);
and U12914 (N_12914,N_9020,N_8759);
and U12915 (N_12915,N_9631,N_7613);
or U12916 (N_12916,N_7973,N_7919);
nor U12917 (N_12917,N_5491,N_8553);
nor U12918 (N_12918,N_5730,N_5757);
and U12919 (N_12919,N_6421,N_5795);
and U12920 (N_12920,N_8019,N_5403);
or U12921 (N_12921,N_8814,N_6493);
nand U12922 (N_12922,N_5062,N_9881);
xor U12923 (N_12923,N_7478,N_8026);
xnor U12924 (N_12924,N_6447,N_8130);
or U12925 (N_12925,N_9856,N_8432);
xnor U12926 (N_12926,N_5789,N_9226);
and U12927 (N_12927,N_8722,N_7803);
and U12928 (N_12928,N_7891,N_6106);
xnor U12929 (N_12929,N_5923,N_9743);
xnor U12930 (N_12930,N_8155,N_9654);
nor U12931 (N_12931,N_5046,N_6925);
xnor U12932 (N_12932,N_5674,N_8766);
xor U12933 (N_12933,N_9866,N_7820);
nor U12934 (N_12934,N_8030,N_9863);
xor U12935 (N_12935,N_9728,N_7405);
or U12936 (N_12936,N_6637,N_8866);
xnor U12937 (N_12937,N_9658,N_6052);
xor U12938 (N_12938,N_5234,N_6269);
or U12939 (N_12939,N_8645,N_6688);
nor U12940 (N_12940,N_5886,N_5316);
or U12941 (N_12941,N_6238,N_5951);
nand U12942 (N_12942,N_8546,N_5274);
nand U12943 (N_12943,N_8311,N_8365);
and U12944 (N_12944,N_5868,N_5514);
and U12945 (N_12945,N_6646,N_9032);
nand U12946 (N_12946,N_5661,N_9956);
xor U12947 (N_12947,N_8333,N_8536);
and U12948 (N_12948,N_5297,N_9659);
or U12949 (N_12949,N_8135,N_9861);
or U12950 (N_12950,N_6864,N_5382);
or U12951 (N_12951,N_6304,N_8284);
or U12952 (N_12952,N_7598,N_9470);
or U12953 (N_12953,N_6753,N_8830);
and U12954 (N_12954,N_5287,N_7175);
nor U12955 (N_12955,N_9500,N_9046);
nor U12956 (N_12956,N_9992,N_8585);
nor U12957 (N_12957,N_5920,N_6349);
nor U12958 (N_12958,N_9833,N_6112);
nor U12959 (N_12959,N_8177,N_5205);
xnor U12960 (N_12960,N_8977,N_5000);
nor U12961 (N_12961,N_6370,N_9267);
and U12962 (N_12962,N_6050,N_9433);
or U12963 (N_12963,N_9796,N_8249);
xor U12964 (N_12964,N_6652,N_5484);
nor U12965 (N_12965,N_9425,N_9164);
nand U12966 (N_12966,N_8507,N_6284);
xor U12967 (N_12967,N_8483,N_5893);
xor U12968 (N_12968,N_8011,N_5747);
or U12969 (N_12969,N_5995,N_7056);
xor U12970 (N_12970,N_9219,N_8189);
or U12971 (N_12971,N_9604,N_5098);
or U12972 (N_12972,N_6344,N_9780);
nor U12973 (N_12973,N_9789,N_6870);
xnor U12974 (N_12974,N_6302,N_7233);
nand U12975 (N_12975,N_8493,N_6272);
and U12976 (N_12976,N_7284,N_5632);
or U12977 (N_12977,N_9999,N_8694);
nand U12978 (N_12978,N_5978,N_5440);
and U12979 (N_12979,N_6422,N_9057);
nand U12980 (N_12980,N_5591,N_5283);
and U12981 (N_12981,N_8309,N_9770);
nand U12982 (N_12982,N_8906,N_8349);
or U12983 (N_12983,N_8281,N_5464);
and U12984 (N_12984,N_9268,N_5910);
nor U12985 (N_12985,N_7425,N_6131);
or U12986 (N_12986,N_5917,N_5286);
nand U12987 (N_12987,N_6529,N_8338);
xor U12988 (N_12988,N_8200,N_5344);
nand U12989 (N_12989,N_8686,N_6305);
xor U12990 (N_12990,N_7818,N_6682);
and U12991 (N_12991,N_7250,N_6965);
nor U12992 (N_12992,N_5833,N_5588);
or U12993 (N_12993,N_5341,N_9370);
nor U12994 (N_12994,N_9495,N_8011);
xnor U12995 (N_12995,N_9932,N_5256);
or U12996 (N_12996,N_5464,N_5358);
nor U12997 (N_12997,N_9394,N_5680);
or U12998 (N_12998,N_9698,N_6558);
nor U12999 (N_12999,N_8945,N_6505);
xnor U13000 (N_13000,N_8714,N_8788);
or U13001 (N_13001,N_5815,N_7681);
xor U13002 (N_13002,N_7377,N_8998);
xor U13003 (N_13003,N_5702,N_7372);
nand U13004 (N_13004,N_8769,N_9660);
nor U13005 (N_13005,N_5780,N_5382);
xnor U13006 (N_13006,N_9927,N_9587);
and U13007 (N_13007,N_9568,N_6884);
nor U13008 (N_13008,N_6330,N_8136);
xor U13009 (N_13009,N_5064,N_9772);
or U13010 (N_13010,N_7698,N_5224);
and U13011 (N_13011,N_9087,N_6507);
or U13012 (N_13012,N_5013,N_7451);
and U13013 (N_13013,N_5147,N_6272);
and U13014 (N_13014,N_9735,N_9084);
or U13015 (N_13015,N_9577,N_8586);
xnor U13016 (N_13016,N_7917,N_5492);
nor U13017 (N_13017,N_9583,N_6581);
xnor U13018 (N_13018,N_7327,N_5781);
or U13019 (N_13019,N_8905,N_9936);
or U13020 (N_13020,N_8848,N_7264);
nor U13021 (N_13021,N_5434,N_7325);
nand U13022 (N_13022,N_9580,N_7661);
xor U13023 (N_13023,N_9818,N_8409);
xor U13024 (N_13024,N_8857,N_7394);
nand U13025 (N_13025,N_5752,N_6199);
nand U13026 (N_13026,N_7225,N_8236);
and U13027 (N_13027,N_7632,N_6506);
or U13028 (N_13028,N_6995,N_7149);
nand U13029 (N_13029,N_6309,N_8973);
xor U13030 (N_13030,N_9985,N_6211);
and U13031 (N_13031,N_9530,N_5531);
nand U13032 (N_13032,N_9483,N_6818);
or U13033 (N_13033,N_9661,N_8343);
and U13034 (N_13034,N_7961,N_5479);
nor U13035 (N_13035,N_9251,N_7262);
or U13036 (N_13036,N_7585,N_6532);
xnor U13037 (N_13037,N_8377,N_5492);
nor U13038 (N_13038,N_5537,N_8540);
nand U13039 (N_13039,N_5983,N_6007);
nor U13040 (N_13040,N_5134,N_5680);
and U13041 (N_13041,N_5520,N_9379);
and U13042 (N_13042,N_6843,N_8497);
or U13043 (N_13043,N_5610,N_7432);
xnor U13044 (N_13044,N_5044,N_8636);
and U13045 (N_13045,N_6096,N_6952);
and U13046 (N_13046,N_6272,N_9169);
nand U13047 (N_13047,N_7003,N_8243);
xnor U13048 (N_13048,N_9942,N_8455);
nor U13049 (N_13049,N_7795,N_7270);
xnor U13050 (N_13050,N_8567,N_6693);
xnor U13051 (N_13051,N_9816,N_6768);
nand U13052 (N_13052,N_7243,N_9695);
or U13053 (N_13053,N_5223,N_9260);
xnor U13054 (N_13054,N_8553,N_5949);
and U13055 (N_13055,N_7885,N_5109);
nor U13056 (N_13056,N_6226,N_5105);
and U13057 (N_13057,N_7656,N_8849);
and U13058 (N_13058,N_5819,N_9983);
and U13059 (N_13059,N_8390,N_9188);
or U13060 (N_13060,N_5331,N_7839);
or U13061 (N_13061,N_7427,N_5168);
nand U13062 (N_13062,N_7847,N_5043);
and U13063 (N_13063,N_8831,N_7390);
and U13064 (N_13064,N_7048,N_6241);
and U13065 (N_13065,N_7554,N_6103);
and U13066 (N_13066,N_8890,N_8883);
and U13067 (N_13067,N_8881,N_7335);
or U13068 (N_13068,N_9525,N_9935);
xnor U13069 (N_13069,N_7107,N_7634);
nor U13070 (N_13070,N_9091,N_8490);
and U13071 (N_13071,N_7640,N_5102);
or U13072 (N_13072,N_8553,N_8794);
nor U13073 (N_13073,N_9022,N_7569);
or U13074 (N_13074,N_6451,N_9038);
and U13075 (N_13075,N_9646,N_6570);
xnor U13076 (N_13076,N_9069,N_8713);
and U13077 (N_13077,N_8547,N_8062);
nor U13078 (N_13078,N_5955,N_9603);
xor U13079 (N_13079,N_7053,N_8342);
or U13080 (N_13080,N_6065,N_5209);
nand U13081 (N_13081,N_5035,N_5098);
xor U13082 (N_13082,N_8259,N_8615);
nand U13083 (N_13083,N_7703,N_9870);
nand U13084 (N_13084,N_9486,N_6032);
and U13085 (N_13085,N_8533,N_7018);
and U13086 (N_13086,N_6716,N_9685);
nand U13087 (N_13087,N_7378,N_9863);
and U13088 (N_13088,N_9075,N_9240);
xor U13089 (N_13089,N_7717,N_5090);
and U13090 (N_13090,N_9657,N_7909);
nand U13091 (N_13091,N_8946,N_5712);
nand U13092 (N_13092,N_7821,N_9017);
or U13093 (N_13093,N_8303,N_8719);
xnor U13094 (N_13094,N_9347,N_5687);
xor U13095 (N_13095,N_9259,N_8782);
or U13096 (N_13096,N_8644,N_9958);
xor U13097 (N_13097,N_5875,N_7104);
nor U13098 (N_13098,N_8103,N_7651);
nor U13099 (N_13099,N_5819,N_7115);
xor U13100 (N_13100,N_5842,N_6080);
nor U13101 (N_13101,N_6529,N_7579);
nor U13102 (N_13102,N_9437,N_8391);
xnor U13103 (N_13103,N_9522,N_9295);
nand U13104 (N_13104,N_6831,N_9221);
xor U13105 (N_13105,N_6707,N_6817);
xor U13106 (N_13106,N_5210,N_7336);
xnor U13107 (N_13107,N_7374,N_6038);
xor U13108 (N_13108,N_9670,N_7882);
nor U13109 (N_13109,N_5005,N_9473);
or U13110 (N_13110,N_8753,N_9305);
xnor U13111 (N_13111,N_9714,N_8382);
nand U13112 (N_13112,N_9576,N_9454);
and U13113 (N_13113,N_5275,N_7776);
or U13114 (N_13114,N_9071,N_6318);
and U13115 (N_13115,N_9386,N_8177);
xnor U13116 (N_13116,N_8331,N_7857);
and U13117 (N_13117,N_8757,N_7132);
or U13118 (N_13118,N_8480,N_8370);
and U13119 (N_13119,N_8925,N_9319);
nand U13120 (N_13120,N_8044,N_6685);
nor U13121 (N_13121,N_9168,N_6498);
and U13122 (N_13122,N_7843,N_8759);
nor U13123 (N_13123,N_9371,N_9857);
and U13124 (N_13124,N_9974,N_7009);
and U13125 (N_13125,N_9422,N_7154);
nor U13126 (N_13126,N_8866,N_7350);
or U13127 (N_13127,N_8751,N_8986);
nor U13128 (N_13128,N_8340,N_5005);
xor U13129 (N_13129,N_6295,N_5185);
and U13130 (N_13130,N_8294,N_5630);
xor U13131 (N_13131,N_8863,N_7704);
or U13132 (N_13132,N_8831,N_8838);
nand U13133 (N_13133,N_7919,N_6261);
or U13134 (N_13134,N_7248,N_7645);
nand U13135 (N_13135,N_6827,N_9085);
or U13136 (N_13136,N_8189,N_9395);
nand U13137 (N_13137,N_8216,N_6386);
and U13138 (N_13138,N_8315,N_6465);
nor U13139 (N_13139,N_5833,N_8919);
nor U13140 (N_13140,N_6166,N_8068);
nor U13141 (N_13141,N_7315,N_6596);
nand U13142 (N_13142,N_7821,N_6142);
nand U13143 (N_13143,N_5230,N_7693);
or U13144 (N_13144,N_6647,N_7509);
nand U13145 (N_13145,N_9628,N_8175);
xnor U13146 (N_13146,N_8676,N_5225);
nor U13147 (N_13147,N_6841,N_6001);
or U13148 (N_13148,N_8644,N_8803);
nor U13149 (N_13149,N_8984,N_8842);
nor U13150 (N_13150,N_7814,N_9165);
nand U13151 (N_13151,N_5203,N_6804);
nand U13152 (N_13152,N_5139,N_5516);
and U13153 (N_13153,N_6116,N_5730);
nor U13154 (N_13154,N_6544,N_7799);
nand U13155 (N_13155,N_8783,N_8926);
nor U13156 (N_13156,N_8887,N_9642);
or U13157 (N_13157,N_7458,N_7634);
nand U13158 (N_13158,N_5751,N_6738);
xnor U13159 (N_13159,N_7457,N_5498);
or U13160 (N_13160,N_9342,N_7183);
nor U13161 (N_13161,N_9584,N_9180);
or U13162 (N_13162,N_7899,N_5314);
or U13163 (N_13163,N_5874,N_5338);
nand U13164 (N_13164,N_6045,N_6034);
nand U13165 (N_13165,N_9746,N_8245);
nand U13166 (N_13166,N_8357,N_8485);
xor U13167 (N_13167,N_8899,N_6645);
nor U13168 (N_13168,N_5095,N_8173);
nor U13169 (N_13169,N_7011,N_5968);
nor U13170 (N_13170,N_8902,N_9512);
nand U13171 (N_13171,N_5784,N_5935);
and U13172 (N_13172,N_6828,N_6599);
nor U13173 (N_13173,N_6117,N_5873);
and U13174 (N_13174,N_9077,N_7369);
or U13175 (N_13175,N_9606,N_5156);
or U13176 (N_13176,N_7527,N_7688);
xnor U13177 (N_13177,N_5904,N_6031);
and U13178 (N_13178,N_9797,N_8529);
nand U13179 (N_13179,N_9097,N_6390);
and U13180 (N_13180,N_6034,N_8544);
and U13181 (N_13181,N_8951,N_5145);
nand U13182 (N_13182,N_9176,N_8547);
nor U13183 (N_13183,N_8460,N_5977);
xor U13184 (N_13184,N_7473,N_7212);
xnor U13185 (N_13185,N_5209,N_5682);
or U13186 (N_13186,N_5593,N_8595);
or U13187 (N_13187,N_9524,N_9342);
or U13188 (N_13188,N_5212,N_6776);
xor U13189 (N_13189,N_5908,N_9555);
or U13190 (N_13190,N_7923,N_8342);
nand U13191 (N_13191,N_6483,N_7045);
nand U13192 (N_13192,N_5505,N_5214);
xnor U13193 (N_13193,N_5771,N_6701);
xor U13194 (N_13194,N_9865,N_9278);
nor U13195 (N_13195,N_9727,N_8626);
or U13196 (N_13196,N_7039,N_6092);
xor U13197 (N_13197,N_9975,N_9918);
and U13198 (N_13198,N_7648,N_8440);
or U13199 (N_13199,N_8863,N_5211);
and U13200 (N_13200,N_5104,N_8048);
or U13201 (N_13201,N_7341,N_5897);
nand U13202 (N_13202,N_8040,N_6413);
xnor U13203 (N_13203,N_6968,N_6326);
xnor U13204 (N_13204,N_6339,N_7920);
nor U13205 (N_13205,N_7974,N_8303);
and U13206 (N_13206,N_8146,N_9644);
and U13207 (N_13207,N_6632,N_6484);
or U13208 (N_13208,N_7182,N_6847);
and U13209 (N_13209,N_7636,N_5289);
xnor U13210 (N_13210,N_9660,N_7121);
xnor U13211 (N_13211,N_5659,N_5539);
xor U13212 (N_13212,N_8110,N_7076);
xor U13213 (N_13213,N_6838,N_7636);
xor U13214 (N_13214,N_6997,N_8348);
nand U13215 (N_13215,N_7119,N_6135);
and U13216 (N_13216,N_8571,N_9570);
or U13217 (N_13217,N_9142,N_7441);
and U13218 (N_13218,N_5802,N_5723);
and U13219 (N_13219,N_8475,N_6408);
or U13220 (N_13220,N_7487,N_7032);
xor U13221 (N_13221,N_8018,N_5673);
and U13222 (N_13222,N_5112,N_9534);
nand U13223 (N_13223,N_6284,N_6379);
and U13224 (N_13224,N_7473,N_7878);
xor U13225 (N_13225,N_9720,N_9129);
or U13226 (N_13226,N_6167,N_8218);
nor U13227 (N_13227,N_7834,N_8396);
xnor U13228 (N_13228,N_5458,N_7827);
and U13229 (N_13229,N_9076,N_7850);
xor U13230 (N_13230,N_6913,N_8339);
nand U13231 (N_13231,N_9667,N_7617);
and U13232 (N_13232,N_9653,N_8975);
nor U13233 (N_13233,N_5975,N_9883);
or U13234 (N_13234,N_8560,N_9816);
xnor U13235 (N_13235,N_8599,N_5276);
nor U13236 (N_13236,N_9286,N_5086);
or U13237 (N_13237,N_8347,N_7791);
or U13238 (N_13238,N_6675,N_5310);
xor U13239 (N_13239,N_8985,N_5086);
xnor U13240 (N_13240,N_7838,N_7081);
or U13241 (N_13241,N_6843,N_6217);
or U13242 (N_13242,N_6785,N_8006);
nand U13243 (N_13243,N_8344,N_8686);
or U13244 (N_13244,N_9254,N_7900);
or U13245 (N_13245,N_9603,N_6523);
xor U13246 (N_13246,N_7456,N_8712);
and U13247 (N_13247,N_5013,N_8369);
nor U13248 (N_13248,N_5705,N_5641);
or U13249 (N_13249,N_8923,N_9138);
or U13250 (N_13250,N_8367,N_8600);
xnor U13251 (N_13251,N_8702,N_7552);
nand U13252 (N_13252,N_6464,N_8164);
nand U13253 (N_13253,N_8760,N_6147);
xor U13254 (N_13254,N_9143,N_5222);
nor U13255 (N_13255,N_7287,N_9423);
or U13256 (N_13256,N_7303,N_7029);
and U13257 (N_13257,N_5468,N_8516);
nor U13258 (N_13258,N_8042,N_8566);
nor U13259 (N_13259,N_9889,N_6006);
nor U13260 (N_13260,N_6931,N_7929);
or U13261 (N_13261,N_6612,N_9135);
or U13262 (N_13262,N_5451,N_8111);
and U13263 (N_13263,N_6818,N_9120);
nand U13264 (N_13264,N_8138,N_5012);
and U13265 (N_13265,N_7754,N_8215);
nand U13266 (N_13266,N_6323,N_8811);
or U13267 (N_13267,N_8172,N_7252);
or U13268 (N_13268,N_9224,N_6750);
xnor U13269 (N_13269,N_7376,N_7739);
and U13270 (N_13270,N_8942,N_5219);
and U13271 (N_13271,N_5468,N_7591);
nand U13272 (N_13272,N_5856,N_8539);
xnor U13273 (N_13273,N_7944,N_6489);
xor U13274 (N_13274,N_5232,N_5104);
and U13275 (N_13275,N_5385,N_5510);
nor U13276 (N_13276,N_9859,N_9332);
nor U13277 (N_13277,N_5920,N_9150);
nand U13278 (N_13278,N_5680,N_8197);
and U13279 (N_13279,N_9215,N_6590);
nand U13280 (N_13280,N_6687,N_9050);
or U13281 (N_13281,N_6001,N_5529);
xnor U13282 (N_13282,N_6665,N_7393);
and U13283 (N_13283,N_5157,N_7716);
or U13284 (N_13284,N_6989,N_7916);
nand U13285 (N_13285,N_5448,N_5135);
xnor U13286 (N_13286,N_8716,N_5714);
nand U13287 (N_13287,N_9178,N_9311);
xor U13288 (N_13288,N_7599,N_6252);
nand U13289 (N_13289,N_7881,N_6123);
nand U13290 (N_13290,N_6140,N_5285);
xnor U13291 (N_13291,N_8563,N_5885);
xnor U13292 (N_13292,N_6041,N_8863);
xnor U13293 (N_13293,N_5857,N_5724);
xnor U13294 (N_13294,N_6360,N_6090);
and U13295 (N_13295,N_8975,N_9966);
nor U13296 (N_13296,N_9960,N_5038);
nor U13297 (N_13297,N_5162,N_8976);
xnor U13298 (N_13298,N_5010,N_6031);
and U13299 (N_13299,N_9726,N_9225);
and U13300 (N_13300,N_6268,N_5840);
or U13301 (N_13301,N_8647,N_7066);
nor U13302 (N_13302,N_8501,N_9631);
xor U13303 (N_13303,N_9357,N_5265);
or U13304 (N_13304,N_6488,N_9077);
or U13305 (N_13305,N_6972,N_7431);
nor U13306 (N_13306,N_7796,N_5841);
nand U13307 (N_13307,N_9124,N_6636);
xor U13308 (N_13308,N_8198,N_7653);
nor U13309 (N_13309,N_6705,N_7128);
xor U13310 (N_13310,N_7050,N_5651);
xnor U13311 (N_13311,N_6956,N_7568);
nand U13312 (N_13312,N_7736,N_5543);
nand U13313 (N_13313,N_7499,N_8572);
nand U13314 (N_13314,N_5451,N_7843);
nand U13315 (N_13315,N_6225,N_8459);
and U13316 (N_13316,N_8807,N_7356);
nor U13317 (N_13317,N_8956,N_6655);
or U13318 (N_13318,N_5058,N_6281);
nand U13319 (N_13319,N_7208,N_9670);
nor U13320 (N_13320,N_7109,N_6378);
xnor U13321 (N_13321,N_6516,N_7280);
nand U13322 (N_13322,N_5607,N_6744);
xor U13323 (N_13323,N_9902,N_7547);
nor U13324 (N_13324,N_7714,N_5053);
or U13325 (N_13325,N_5453,N_8424);
and U13326 (N_13326,N_6533,N_5374);
and U13327 (N_13327,N_7492,N_8298);
xor U13328 (N_13328,N_6518,N_5024);
and U13329 (N_13329,N_8237,N_7045);
or U13330 (N_13330,N_8170,N_5321);
nand U13331 (N_13331,N_6906,N_5540);
nand U13332 (N_13332,N_8810,N_7791);
and U13333 (N_13333,N_8811,N_8184);
and U13334 (N_13334,N_9649,N_9311);
or U13335 (N_13335,N_8427,N_9085);
xnor U13336 (N_13336,N_7519,N_8822);
or U13337 (N_13337,N_6424,N_8257);
or U13338 (N_13338,N_7210,N_9355);
xnor U13339 (N_13339,N_7759,N_5495);
nand U13340 (N_13340,N_7255,N_9551);
or U13341 (N_13341,N_9585,N_5970);
nor U13342 (N_13342,N_8410,N_6431);
nor U13343 (N_13343,N_8016,N_5000);
and U13344 (N_13344,N_9352,N_6152);
and U13345 (N_13345,N_8484,N_5563);
xor U13346 (N_13346,N_7857,N_5792);
or U13347 (N_13347,N_6730,N_7831);
or U13348 (N_13348,N_9570,N_6787);
nor U13349 (N_13349,N_6605,N_6551);
and U13350 (N_13350,N_6085,N_9720);
or U13351 (N_13351,N_5994,N_8307);
and U13352 (N_13352,N_5066,N_8916);
nand U13353 (N_13353,N_9564,N_8425);
xnor U13354 (N_13354,N_8083,N_5941);
xnor U13355 (N_13355,N_7447,N_7272);
or U13356 (N_13356,N_8838,N_8026);
nand U13357 (N_13357,N_9200,N_6295);
nor U13358 (N_13358,N_9159,N_6593);
or U13359 (N_13359,N_7973,N_7135);
xnor U13360 (N_13360,N_7112,N_6941);
nand U13361 (N_13361,N_6411,N_8515);
nand U13362 (N_13362,N_8175,N_8935);
nand U13363 (N_13363,N_6547,N_9852);
nand U13364 (N_13364,N_7232,N_6172);
nor U13365 (N_13365,N_8400,N_7871);
nand U13366 (N_13366,N_8021,N_7942);
nor U13367 (N_13367,N_7358,N_8460);
or U13368 (N_13368,N_7316,N_6017);
or U13369 (N_13369,N_8024,N_5458);
and U13370 (N_13370,N_5650,N_9189);
nand U13371 (N_13371,N_5425,N_5638);
or U13372 (N_13372,N_7107,N_6608);
and U13373 (N_13373,N_7644,N_7782);
and U13374 (N_13374,N_5661,N_9706);
nand U13375 (N_13375,N_7892,N_7162);
xor U13376 (N_13376,N_6898,N_6382);
nor U13377 (N_13377,N_6178,N_8674);
and U13378 (N_13378,N_9437,N_8989);
nor U13379 (N_13379,N_7265,N_7095);
nor U13380 (N_13380,N_5152,N_6915);
or U13381 (N_13381,N_5635,N_7664);
and U13382 (N_13382,N_7700,N_8156);
or U13383 (N_13383,N_6947,N_5989);
nand U13384 (N_13384,N_6990,N_5598);
and U13385 (N_13385,N_8885,N_5786);
nor U13386 (N_13386,N_6649,N_9037);
nor U13387 (N_13387,N_8911,N_9808);
or U13388 (N_13388,N_7062,N_9999);
nand U13389 (N_13389,N_6605,N_7040);
nand U13390 (N_13390,N_9530,N_5841);
nor U13391 (N_13391,N_5892,N_9539);
and U13392 (N_13392,N_5451,N_7454);
nand U13393 (N_13393,N_6074,N_9117);
or U13394 (N_13394,N_6951,N_9758);
or U13395 (N_13395,N_6730,N_9774);
xnor U13396 (N_13396,N_5372,N_9559);
or U13397 (N_13397,N_7594,N_9786);
nor U13398 (N_13398,N_9599,N_9746);
nor U13399 (N_13399,N_7494,N_7072);
nor U13400 (N_13400,N_6138,N_7210);
xor U13401 (N_13401,N_7064,N_8860);
nand U13402 (N_13402,N_9098,N_6033);
and U13403 (N_13403,N_5403,N_6082);
nor U13404 (N_13404,N_7132,N_6158);
and U13405 (N_13405,N_6812,N_5673);
nor U13406 (N_13406,N_8973,N_5353);
and U13407 (N_13407,N_8999,N_8204);
and U13408 (N_13408,N_7671,N_8969);
and U13409 (N_13409,N_5532,N_6796);
or U13410 (N_13410,N_9718,N_7987);
xnor U13411 (N_13411,N_7678,N_9435);
and U13412 (N_13412,N_7177,N_6832);
nand U13413 (N_13413,N_7562,N_9255);
and U13414 (N_13414,N_7758,N_9961);
nand U13415 (N_13415,N_9773,N_5307);
or U13416 (N_13416,N_7830,N_9049);
xnor U13417 (N_13417,N_9472,N_6294);
xnor U13418 (N_13418,N_9519,N_7463);
or U13419 (N_13419,N_5069,N_8544);
nor U13420 (N_13420,N_6173,N_6156);
and U13421 (N_13421,N_5183,N_6589);
and U13422 (N_13422,N_7410,N_7469);
and U13423 (N_13423,N_9798,N_8258);
nor U13424 (N_13424,N_9803,N_8388);
nor U13425 (N_13425,N_9941,N_5379);
nand U13426 (N_13426,N_9765,N_9299);
nand U13427 (N_13427,N_5045,N_7310);
or U13428 (N_13428,N_7504,N_7186);
xor U13429 (N_13429,N_5537,N_8293);
xnor U13430 (N_13430,N_7654,N_8016);
nor U13431 (N_13431,N_8233,N_6165);
nand U13432 (N_13432,N_6658,N_7671);
and U13433 (N_13433,N_7698,N_8841);
and U13434 (N_13434,N_5006,N_7866);
and U13435 (N_13435,N_8444,N_9181);
nor U13436 (N_13436,N_9754,N_7972);
nor U13437 (N_13437,N_6439,N_5604);
nand U13438 (N_13438,N_8277,N_8000);
xor U13439 (N_13439,N_6878,N_8568);
nand U13440 (N_13440,N_5131,N_8334);
xnor U13441 (N_13441,N_9345,N_6586);
xor U13442 (N_13442,N_6964,N_9478);
nor U13443 (N_13443,N_7888,N_5413);
xnor U13444 (N_13444,N_7144,N_8594);
nor U13445 (N_13445,N_5081,N_8991);
xor U13446 (N_13446,N_6168,N_5454);
or U13447 (N_13447,N_7569,N_8480);
nor U13448 (N_13448,N_7856,N_8895);
xor U13449 (N_13449,N_6556,N_8377);
and U13450 (N_13450,N_7642,N_7081);
nand U13451 (N_13451,N_8450,N_5068);
nand U13452 (N_13452,N_5208,N_8708);
xnor U13453 (N_13453,N_9499,N_6560);
and U13454 (N_13454,N_5754,N_7897);
or U13455 (N_13455,N_8245,N_6215);
or U13456 (N_13456,N_9357,N_8249);
xor U13457 (N_13457,N_6332,N_9937);
nor U13458 (N_13458,N_9905,N_9783);
or U13459 (N_13459,N_6568,N_6458);
xnor U13460 (N_13460,N_9617,N_7997);
and U13461 (N_13461,N_7584,N_7737);
xnor U13462 (N_13462,N_8077,N_7718);
xor U13463 (N_13463,N_8530,N_7640);
nor U13464 (N_13464,N_6224,N_6261);
or U13465 (N_13465,N_9455,N_8051);
xnor U13466 (N_13466,N_6376,N_5075);
or U13467 (N_13467,N_7609,N_7756);
xnor U13468 (N_13468,N_9515,N_8429);
and U13469 (N_13469,N_9486,N_5801);
nand U13470 (N_13470,N_5859,N_8700);
or U13471 (N_13471,N_9848,N_8185);
and U13472 (N_13472,N_8174,N_8775);
or U13473 (N_13473,N_7539,N_8033);
or U13474 (N_13474,N_6285,N_9771);
xnor U13475 (N_13475,N_9534,N_9929);
nor U13476 (N_13476,N_8832,N_7061);
or U13477 (N_13477,N_7732,N_9085);
xnor U13478 (N_13478,N_7195,N_6565);
or U13479 (N_13479,N_5097,N_6724);
nor U13480 (N_13480,N_6863,N_5097);
nand U13481 (N_13481,N_5139,N_5493);
and U13482 (N_13482,N_8797,N_6142);
nand U13483 (N_13483,N_5592,N_7504);
and U13484 (N_13484,N_6335,N_5422);
and U13485 (N_13485,N_6924,N_8512);
nor U13486 (N_13486,N_8836,N_6497);
nand U13487 (N_13487,N_6495,N_6854);
or U13488 (N_13488,N_5269,N_5366);
and U13489 (N_13489,N_8909,N_9620);
and U13490 (N_13490,N_8926,N_5383);
or U13491 (N_13491,N_8413,N_7437);
and U13492 (N_13492,N_5797,N_5176);
and U13493 (N_13493,N_9337,N_7835);
nand U13494 (N_13494,N_7799,N_6170);
xor U13495 (N_13495,N_8742,N_9702);
and U13496 (N_13496,N_8334,N_7169);
and U13497 (N_13497,N_5675,N_6304);
nor U13498 (N_13498,N_6114,N_7731);
and U13499 (N_13499,N_7787,N_9021);
nor U13500 (N_13500,N_8125,N_9355);
and U13501 (N_13501,N_6832,N_5115);
nor U13502 (N_13502,N_8923,N_6398);
or U13503 (N_13503,N_9986,N_5220);
nand U13504 (N_13504,N_5797,N_8015);
or U13505 (N_13505,N_9921,N_7042);
nor U13506 (N_13506,N_9881,N_5105);
and U13507 (N_13507,N_5992,N_5254);
and U13508 (N_13508,N_7095,N_9489);
or U13509 (N_13509,N_7074,N_8047);
or U13510 (N_13510,N_7798,N_9786);
nor U13511 (N_13511,N_5067,N_5199);
or U13512 (N_13512,N_8425,N_8851);
nand U13513 (N_13513,N_5144,N_5431);
nand U13514 (N_13514,N_9902,N_5892);
or U13515 (N_13515,N_6951,N_9508);
xor U13516 (N_13516,N_9102,N_7234);
xor U13517 (N_13517,N_9402,N_5149);
and U13518 (N_13518,N_6639,N_5562);
and U13519 (N_13519,N_7289,N_7039);
and U13520 (N_13520,N_9878,N_7418);
xor U13521 (N_13521,N_8099,N_8007);
xor U13522 (N_13522,N_6775,N_6684);
and U13523 (N_13523,N_6901,N_9923);
and U13524 (N_13524,N_6313,N_9548);
and U13525 (N_13525,N_6150,N_5499);
or U13526 (N_13526,N_8876,N_6873);
or U13527 (N_13527,N_8784,N_5461);
and U13528 (N_13528,N_8560,N_7884);
or U13529 (N_13529,N_7245,N_5870);
nor U13530 (N_13530,N_5879,N_8101);
nor U13531 (N_13531,N_8407,N_5994);
and U13532 (N_13532,N_9371,N_6946);
or U13533 (N_13533,N_8487,N_7096);
nand U13534 (N_13534,N_7250,N_7613);
nor U13535 (N_13535,N_7973,N_8422);
and U13536 (N_13536,N_6028,N_9136);
xor U13537 (N_13537,N_6118,N_7397);
nand U13538 (N_13538,N_6509,N_7193);
nor U13539 (N_13539,N_5512,N_6604);
nor U13540 (N_13540,N_7796,N_5050);
nand U13541 (N_13541,N_9606,N_9503);
nor U13542 (N_13542,N_6216,N_9804);
nor U13543 (N_13543,N_8443,N_9486);
xor U13544 (N_13544,N_6308,N_9605);
nor U13545 (N_13545,N_7987,N_8015);
nor U13546 (N_13546,N_5718,N_8031);
or U13547 (N_13547,N_7269,N_6423);
xor U13548 (N_13548,N_9362,N_6023);
or U13549 (N_13549,N_7636,N_7900);
or U13550 (N_13550,N_7034,N_8322);
nand U13551 (N_13551,N_8211,N_8898);
nor U13552 (N_13552,N_8332,N_6053);
and U13553 (N_13553,N_7129,N_8745);
nor U13554 (N_13554,N_5435,N_9563);
xor U13555 (N_13555,N_7479,N_5854);
xnor U13556 (N_13556,N_5775,N_6088);
and U13557 (N_13557,N_8965,N_9313);
nor U13558 (N_13558,N_9630,N_5490);
and U13559 (N_13559,N_5064,N_8491);
or U13560 (N_13560,N_8807,N_6246);
xnor U13561 (N_13561,N_8499,N_5700);
nand U13562 (N_13562,N_5942,N_6463);
or U13563 (N_13563,N_5627,N_7601);
and U13564 (N_13564,N_6862,N_5536);
xor U13565 (N_13565,N_6957,N_9325);
nand U13566 (N_13566,N_8145,N_7027);
nor U13567 (N_13567,N_6527,N_8241);
nor U13568 (N_13568,N_5144,N_7756);
and U13569 (N_13569,N_6320,N_7103);
and U13570 (N_13570,N_8322,N_6336);
and U13571 (N_13571,N_5681,N_6459);
xor U13572 (N_13572,N_9047,N_9432);
xnor U13573 (N_13573,N_8496,N_5251);
nand U13574 (N_13574,N_5739,N_5763);
and U13575 (N_13575,N_6863,N_5294);
xor U13576 (N_13576,N_7175,N_8705);
nor U13577 (N_13577,N_6973,N_5466);
xor U13578 (N_13578,N_9086,N_7108);
and U13579 (N_13579,N_9610,N_6758);
or U13580 (N_13580,N_8112,N_6113);
or U13581 (N_13581,N_7393,N_7641);
nor U13582 (N_13582,N_7603,N_9851);
xnor U13583 (N_13583,N_7757,N_6946);
nor U13584 (N_13584,N_6619,N_5163);
and U13585 (N_13585,N_7543,N_7455);
xnor U13586 (N_13586,N_6877,N_7881);
xnor U13587 (N_13587,N_6192,N_9307);
and U13588 (N_13588,N_9919,N_6583);
nand U13589 (N_13589,N_7534,N_7128);
xnor U13590 (N_13590,N_6454,N_9971);
and U13591 (N_13591,N_7067,N_9853);
nor U13592 (N_13592,N_8830,N_6484);
nor U13593 (N_13593,N_8444,N_5871);
nor U13594 (N_13594,N_5540,N_9308);
and U13595 (N_13595,N_8775,N_9598);
xnor U13596 (N_13596,N_8228,N_7358);
xnor U13597 (N_13597,N_5114,N_9806);
xnor U13598 (N_13598,N_9677,N_7472);
nand U13599 (N_13599,N_9964,N_8484);
or U13600 (N_13600,N_8893,N_8922);
or U13601 (N_13601,N_6583,N_5950);
and U13602 (N_13602,N_8373,N_9101);
or U13603 (N_13603,N_7385,N_9933);
nor U13604 (N_13604,N_8707,N_6415);
nor U13605 (N_13605,N_8182,N_7292);
nor U13606 (N_13606,N_6377,N_7834);
nand U13607 (N_13607,N_7743,N_9582);
or U13608 (N_13608,N_6718,N_9992);
xnor U13609 (N_13609,N_5361,N_9855);
nand U13610 (N_13610,N_6481,N_5098);
or U13611 (N_13611,N_9107,N_6249);
nor U13612 (N_13612,N_9796,N_6666);
xnor U13613 (N_13613,N_7600,N_9666);
xnor U13614 (N_13614,N_7264,N_9448);
and U13615 (N_13615,N_8339,N_5815);
or U13616 (N_13616,N_6017,N_5989);
xor U13617 (N_13617,N_7285,N_7830);
nor U13618 (N_13618,N_9962,N_9999);
nand U13619 (N_13619,N_8860,N_9123);
or U13620 (N_13620,N_6773,N_8880);
xnor U13621 (N_13621,N_7827,N_5917);
xnor U13622 (N_13622,N_6423,N_9218);
or U13623 (N_13623,N_9263,N_6860);
or U13624 (N_13624,N_7509,N_9715);
or U13625 (N_13625,N_7995,N_5902);
xnor U13626 (N_13626,N_8996,N_5503);
or U13627 (N_13627,N_6893,N_8632);
nor U13628 (N_13628,N_5142,N_5662);
or U13629 (N_13629,N_8275,N_5180);
and U13630 (N_13630,N_9586,N_5458);
and U13631 (N_13631,N_6713,N_7549);
xnor U13632 (N_13632,N_5239,N_9609);
xnor U13633 (N_13633,N_7462,N_8893);
or U13634 (N_13634,N_5493,N_9567);
and U13635 (N_13635,N_7304,N_6605);
or U13636 (N_13636,N_9878,N_9897);
nand U13637 (N_13637,N_9037,N_5547);
nand U13638 (N_13638,N_5463,N_6714);
or U13639 (N_13639,N_6395,N_9039);
nand U13640 (N_13640,N_8703,N_6930);
nand U13641 (N_13641,N_5546,N_8606);
nand U13642 (N_13642,N_6144,N_9985);
and U13643 (N_13643,N_7245,N_8718);
or U13644 (N_13644,N_8096,N_5540);
xor U13645 (N_13645,N_5931,N_8712);
and U13646 (N_13646,N_5999,N_5057);
or U13647 (N_13647,N_5212,N_8604);
nand U13648 (N_13648,N_8299,N_9810);
and U13649 (N_13649,N_8898,N_8000);
xor U13650 (N_13650,N_8266,N_9832);
xnor U13651 (N_13651,N_6516,N_7407);
nand U13652 (N_13652,N_7451,N_6127);
or U13653 (N_13653,N_5496,N_8715);
nor U13654 (N_13654,N_7292,N_5654);
xnor U13655 (N_13655,N_8891,N_5300);
nor U13656 (N_13656,N_7843,N_7884);
or U13657 (N_13657,N_8691,N_6262);
nor U13658 (N_13658,N_6864,N_8227);
and U13659 (N_13659,N_6652,N_6564);
nor U13660 (N_13660,N_7620,N_5334);
and U13661 (N_13661,N_9487,N_9760);
xor U13662 (N_13662,N_8026,N_5752);
xor U13663 (N_13663,N_5284,N_9064);
nor U13664 (N_13664,N_6857,N_9765);
or U13665 (N_13665,N_8152,N_6684);
nor U13666 (N_13666,N_9377,N_5939);
nand U13667 (N_13667,N_7939,N_9645);
and U13668 (N_13668,N_5857,N_9478);
nor U13669 (N_13669,N_9854,N_6691);
xnor U13670 (N_13670,N_5085,N_5956);
xor U13671 (N_13671,N_7551,N_5189);
or U13672 (N_13672,N_8610,N_6130);
nor U13673 (N_13673,N_9356,N_7808);
or U13674 (N_13674,N_5844,N_6583);
or U13675 (N_13675,N_9830,N_9086);
xnor U13676 (N_13676,N_9976,N_5339);
or U13677 (N_13677,N_8593,N_8783);
xor U13678 (N_13678,N_9252,N_7748);
xnor U13679 (N_13679,N_7612,N_9174);
or U13680 (N_13680,N_5499,N_7103);
nor U13681 (N_13681,N_7058,N_6553);
nand U13682 (N_13682,N_6210,N_6913);
xor U13683 (N_13683,N_9064,N_7462);
and U13684 (N_13684,N_8178,N_7368);
xnor U13685 (N_13685,N_7485,N_7626);
nand U13686 (N_13686,N_7684,N_7080);
or U13687 (N_13687,N_7787,N_6642);
nand U13688 (N_13688,N_8454,N_7113);
nand U13689 (N_13689,N_7698,N_8630);
and U13690 (N_13690,N_9449,N_6581);
nor U13691 (N_13691,N_9653,N_9837);
nor U13692 (N_13692,N_6659,N_5705);
or U13693 (N_13693,N_8609,N_9405);
xnor U13694 (N_13694,N_6889,N_5863);
nand U13695 (N_13695,N_9159,N_6438);
xor U13696 (N_13696,N_6848,N_9863);
nor U13697 (N_13697,N_7601,N_8229);
nand U13698 (N_13698,N_6838,N_6297);
nand U13699 (N_13699,N_5468,N_9458);
and U13700 (N_13700,N_8395,N_5188);
nand U13701 (N_13701,N_9222,N_6870);
and U13702 (N_13702,N_6500,N_8243);
nand U13703 (N_13703,N_9185,N_9010);
and U13704 (N_13704,N_8090,N_7773);
nand U13705 (N_13705,N_5747,N_9046);
xor U13706 (N_13706,N_8470,N_8145);
nand U13707 (N_13707,N_7789,N_6745);
nor U13708 (N_13708,N_9326,N_5404);
or U13709 (N_13709,N_6767,N_5619);
nor U13710 (N_13710,N_5683,N_8243);
and U13711 (N_13711,N_9803,N_7933);
nand U13712 (N_13712,N_9198,N_5098);
nor U13713 (N_13713,N_5347,N_8375);
nand U13714 (N_13714,N_7475,N_6741);
nand U13715 (N_13715,N_6475,N_5352);
xnor U13716 (N_13716,N_7584,N_8391);
or U13717 (N_13717,N_6059,N_9739);
xor U13718 (N_13718,N_5027,N_8480);
nor U13719 (N_13719,N_9343,N_6439);
nor U13720 (N_13720,N_7419,N_6915);
nor U13721 (N_13721,N_9568,N_7246);
and U13722 (N_13722,N_6562,N_5633);
nor U13723 (N_13723,N_8236,N_5407);
and U13724 (N_13724,N_9385,N_6481);
xnor U13725 (N_13725,N_9431,N_5075);
nor U13726 (N_13726,N_6247,N_7965);
or U13727 (N_13727,N_8635,N_9900);
xnor U13728 (N_13728,N_7581,N_5648);
and U13729 (N_13729,N_5842,N_6893);
nor U13730 (N_13730,N_6418,N_6722);
or U13731 (N_13731,N_8647,N_8488);
and U13732 (N_13732,N_8234,N_7169);
xnor U13733 (N_13733,N_8363,N_7209);
or U13734 (N_13734,N_8397,N_7891);
xnor U13735 (N_13735,N_6925,N_6022);
and U13736 (N_13736,N_9955,N_7074);
xor U13737 (N_13737,N_9230,N_6260);
xor U13738 (N_13738,N_8488,N_9525);
and U13739 (N_13739,N_9629,N_9964);
or U13740 (N_13740,N_8851,N_5827);
nand U13741 (N_13741,N_7323,N_5812);
or U13742 (N_13742,N_8464,N_6343);
and U13743 (N_13743,N_8291,N_7115);
nand U13744 (N_13744,N_5973,N_7211);
nand U13745 (N_13745,N_5703,N_8138);
and U13746 (N_13746,N_7020,N_8566);
nor U13747 (N_13747,N_5916,N_9209);
and U13748 (N_13748,N_6732,N_5832);
and U13749 (N_13749,N_9106,N_6214);
nor U13750 (N_13750,N_7184,N_7281);
nor U13751 (N_13751,N_9200,N_7844);
nor U13752 (N_13752,N_8244,N_5293);
and U13753 (N_13753,N_6230,N_5258);
nor U13754 (N_13754,N_6871,N_9645);
or U13755 (N_13755,N_9741,N_6457);
nor U13756 (N_13756,N_9607,N_5135);
or U13757 (N_13757,N_5101,N_9095);
nand U13758 (N_13758,N_7912,N_5717);
nand U13759 (N_13759,N_9025,N_5738);
or U13760 (N_13760,N_9287,N_7028);
or U13761 (N_13761,N_5755,N_8207);
or U13762 (N_13762,N_7083,N_6594);
xor U13763 (N_13763,N_5598,N_6798);
and U13764 (N_13764,N_7367,N_8152);
or U13765 (N_13765,N_8002,N_8022);
nand U13766 (N_13766,N_5376,N_9352);
nand U13767 (N_13767,N_6492,N_9361);
nand U13768 (N_13768,N_9791,N_9778);
and U13769 (N_13769,N_9952,N_8240);
nor U13770 (N_13770,N_6024,N_5505);
nand U13771 (N_13771,N_8545,N_9530);
xnor U13772 (N_13772,N_7098,N_6868);
xor U13773 (N_13773,N_7407,N_9528);
or U13774 (N_13774,N_9048,N_8023);
or U13775 (N_13775,N_5634,N_9349);
and U13776 (N_13776,N_9343,N_6167);
or U13777 (N_13777,N_5796,N_5726);
nand U13778 (N_13778,N_8623,N_5807);
or U13779 (N_13779,N_8031,N_8090);
nor U13780 (N_13780,N_6403,N_5016);
or U13781 (N_13781,N_7836,N_8669);
nand U13782 (N_13782,N_5864,N_5445);
nor U13783 (N_13783,N_7411,N_9569);
or U13784 (N_13784,N_5903,N_7621);
or U13785 (N_13785,N_6717,N_6908);
xor U13786 (N_13786,N_9598,N_5439);
or U13787 (N_13787,N_6312,N_7069);
nor U13788 (N_13788,N_6063,N_7255);
nor U13789 (N_13789,N_7621,N_8185);
nor U13790 (N_13790,N_6440,N_8583);
or U13791 (N_13791,N_8649,N_5815);
xnor U13792 (N_13792,N_5132,N_9464);
or U13793 (N_13793,N_6910,N_7835);
and U13794 (N_13794,N_8151,N_8701);
or U13795 (N_13795,N_9513,N_8154);
nand U13796 (N_13796,N_7577,N_5241);
nand U13797 (N_13797,N_6712,N_8998);
nand U13798 (N_13798,N_7372,N_7947);
nand U13799 (N_13799,N_8747,N_7094);
or U13800 (N_13800,N_9355,N_9836);
nor U13801 (N_13801,N_6089,N_6768);
xnor U13802 (N_13802,N_8550,N_8629);
and U13803 (N_13803,N_5546,N_5603);
and U13804 (N_13804,N_9154,N_8054);
or U13805 (N_13805,N_6947,N_5327);
nand U13806 (N_13806,N_5286,N_9817);
or U13807 (N_13807,N_9199,N_8952);
xor U13808 (N_13808,N_5537,N_7946);
and U13809 (N_13809,N_6729,N_5292);
and U13810 (N_13810,N_8375,N_5328);
xor U13811 (N_13811,N_7867,N_6758);
xnor U13812 (N_13812,N_7575,N_6160);
nand U13813 (N_13813,N_7756,N_9013);
xnor U13814 (N_13814,N_9248,N_7388);
or U13815 (N_13815,N_6475,N_9894);
nand U13816 (N_13816,N_8316,N_6084);
nand U13817 (N_13817,N_6746,N_7982);
nand U13818 (N_13818,N_8428,N_6545);
or U13819 (N_13819,N_5697,N_6652);
nand U13820 (N_13820,N_6595,N_8670);
and U13821 (N_13821,N_8791,N_6438);
nand U13822 (N_13822,N_5154,N_5544);
nor U13823 (N_13823,N_6730,N_5231);
nor U13824 (N_13824,N_7601,N_5907);
xor U13825 (N_13825,N_7335,N_6188);
or U13826 (N_13826,N_6795,N_9919);
xnor U13827 (N_13827,N_5849,N_9682);
xor U13828 (N_13828,N_5309,N_6423);
nor U13829 (N_13829,N_8905,N_5891);
nor U13830 (N_13830,N_5512,N_8244);
nor U13831 (N_13831,N_8839,N_9685);
nand U13832 (N_13832,N_7980,N_8962);
nand U13833 (N_13833,N_9325,N_8125);
xor U13834 (N_13834,N_8297,N_8128);
nor U13835 (N_13835,N_5510,N_7568);
and U13836 (N_13836,N_5164,N_7518);
nor U13837 (N_13837,N_5966,N_9529);
and U13838 (N_13838,N_6415,N_9374);
nand U13839 (N_13839,N_6406,N_6836);
nor U13840 (N_13840,N_7262,N_5417);
or U13841 (N_13841,N_7179,N_5178);
nand U13842 (N_13842,N_5012,N_6342);
xnor U13843 (N_13843,N_7364,N_6792);
nor U13844 (N_13844,N_5052,N_8503);
nor U13845 (N_13845,N_8777,N_7787);
nor U13846 (N_13846,N_8545,N_8868);
or U13847 (N_13847,N_8808,N_8181);
nor U13848 (N_13848,N_7417,N_8436);
nor U13849 (N_13849,N_7465,N_8691);
or U13850 (N_13850,N_6519,N_9112);
xnor U13851 (N_13851,N_9374,N_5619);
xnor U13852 (N_13852,N_7693,N_8443);
or U13853 (N_13853,N_6057,N_6802);
nand U13854 (N_13854,N_8733,N_6102);
or U13855 (N_13855,N_9789,N_5418);
xnor U13856 (N_13856,N_5300,N_5997);
and U13857 (N_13857,N_9182,N_9015);
nand U13858 (N_13858,N_5893,N_9396);
and U13859 (N_13859,N_7638,N_7490);
xnor U13860 (N_13860,N_8297,N_8376);
nand U13861 (N_13861,N_5696,N_9748);
nand U13862 (N_13862,N_6777,N_8499);
nor U13863 (N_13863,N_8299,N_9570);
and U13864 (N_13864,N_7430,N_7248);
or U13865 (N_13865,N_5335,N_7826);
xor U13866 (N_13866,N_9884,N_6648);
and U13867 (N_13867,N_8352,N_6174);
xor U13868 (N_13868,N_7168,N_7061);
or U13869 (N_13869,N_7299,N_9377);
or U13870 (N_13870,N_5650,N_5186);
nor U13871 (N_13871,N_6748,N_8276);
and U13872 (N_13872,N_9027,N_7344);
nor U13873 (N_13873,N_7747,N_8009);
and U13874 (N_13874,N_6946,N_9798);
nand U13875 (N_13875,N_5559,N_6278);
or U13876 (N_13876,N_9252,N_8819);
or U13877 (N_13877,N_5017,N_8732);
nand U13878 (N_13878,N_8723,N_7964);
nand U13879 (N_13879,N_5693,N_5015);
nor U13880 (N_13880,N_9822,N_9164);
or U13881 (N_13881,N_5654,N_6507);
nand U13882 (N_13882,N_9466,N_8202);
or U13883 (N_13883,N_9432,N_8644);
and U13884 (N_13884,N_8182,N_6401);
nand U13885 (N_13885,N_6145,N_8598);
or U13886 (N_13886,N_9480,N_7148);
and U13887 (N_13887,N_6954,N_7469);
nor U13888 (N_13888,N_9115,N_8528);
and U13889 (N_13889,N_5207,N_5885);
and U13890 (N_13890,N_9155,N_9209);
nand U13891 (N_13891,N_7280,N_5346);
nor U13892 (N_13892,N_6397,N_9621);
xor U13893 (N_13893,N_7119,N_9311);
xor U13894 (N_13894,N_6161,N_5864);
xor U13895 (N_13895,N_8841,N_9440);
xnor U13896 (N_13896,N_9680,N_5602);
xnor U13897 (N_13897,N_6093,N_6399);
nor U13898 (N_13898,N_9890,N_9687);
and U13899 (N_13899,N_6248,N_8474);
nor U13900 (N_13900,N_9356,N_9775);
and U13901 (N_13901,N_8530,N_6392);
xor U13902 (N_13902,N_8269,N_5470);
or U13903 (N_13903,N_7092,N_6325);
and U13904 (N_13904,N_5818,N_5595);
and U13905 (N_13905,N_8207,N_9035);
or U13906 (N_13906,N_9413,N_9565);
or U13907 (N_13907,N_7953,N_8976);
nand U13908 (N_13908,N_8973,N_8478);
or U13909 (N_13909,N_9883,N_7789);
or U13910 (N_13910,N_9321,N_7732);
nand U13911 (N_13911,N_6785,N_6769);
nand U13912 (N_13912,N_9605,N_8682);
or U13913 (N_13913,N_7141,N_9115);
nand U13914 (N_13914,N_5403,N_5518);
nand U13915 (N_13915,N_7162,N_9137);
and U13916 (N_13916,N_8097,N_5876);
or U13917 (N_13917,N_9734,N_8972);
nand U13918 (N_13918,N_8278,N_8681);
xor U13919 (N_13919,N_5459,N_8715);
and U13920 (N_13920,N_6564,N_5598);
nand U13921 (N_13921,N_8922,N_7745);
or U13922 (N_13922,N_6648,N_5869);
or U13923 (N_13923,N_7363,N_6880);
nor U13924 (N_13924,N_5328,N_9823);
xnor U13925 (N_13925,N_5240,N_9695);
xnor U13926 (N_13926,N_9625,N_6218);
nand U13927 (N_13927,N_6656,N_6272);
xor U13928 (N_13928,N_7882,N_7464);
nor U13929 (N_13929,N_9628,N_8061);
xnor U13930 (N_13930,N_6615,N_9782);
nor U13931 (N_13931,N_7673,N_8241);
or U13932 (N_13932,N_8551,N_8788);
and U13933 (N_13933,N_6235,N_8400);
nor U13934 (N_13934,N_6093,N_7635);
and U13935 (N_13935,N_7289,N_9809);
or U13936 (N_13936,N_5673,N_9148);
xnor U13937 (N_13937,N_6276,N_8115);
or U13938 (N_13938,N_5160,N_9877);
and U13939 (N_13939,N_9088,N_5288);
nand U13940 (N_13940,N_8811,N_7291);
and U13941 (N_13941,N_7466,N_8960);
nand U13942 (N_13942,N_5851,N_8110);
and U13943 (N_13943,N_5528,N_6280);
or U13944 (N_13944,N_5941,N_6597);
xnor U13945 (N_13945,N_7097,N_8019);
and U13946 (N_13946,N_5279,N_8348);
nand U13947 (N_13947,N_5880,N_6024);
nand U13948 (N_13948,N_5453,N_7703);
and U13949 (N_13949,N_5261,N_7634);
xor U13950 (N_13950,N_7014,N_9292);
nor U13951 (N_13951,N_6982,N_6831);
nand U13952 (N_13952,N_8202,N_8914);
and U13953 (N_13953,N_5420,N_7867);
or U13954 (N_13954,N_7117,N_7606);
nor U13955 (N_13955,N_7949,N_5859);
nand U13956 (N_13956,N_9175,N_8479);
nor U13957 (N_13957,N_6131,N_5208);
nand U13958 (N_13958,N_7620,N_7959);
nor U13959 (N_13959,N_8987,N_6051);
and U13960 (N_13960,N_5046,N_6639);
xor U13961 (N_13961,N_7379,N_8068);
nor U13962 (N_13962,N_9912,N_9044);
or U13963 (N_13963,N_9936,N_5562);
or U13964 (N_13964,N_5826,N_7499);
nand U13965 (N_13965,N_8181,N_9279);
and U13966 (N_13966,N_7926,N_7603);
nand U13967 (N_13967,N_6981,N_6097);
nor U13968 (N_13968,N_6781,N_5690);
and U13969 (N_13969,N_9361,N_7889);
or U13970 (N_13970,N_8540,N_9749);
or U13971 (N_13971,N_6747,N_5018);
xor U13972 (N_13972,N_7536,N_6284);
xnor U13973 (N_13973,N_9867,N_5430);
nor U13974 (N_13974,N_6338,N_6730);
xnor U13975 (N_13975,N_6157,N_8885);
and U13976 (N_13976,N_7487,N_8197);
or U13977 (N_13977,N_7780,N_6853);
xnor U13978 (N_13978,N_8605,N_7345);
and U13979 (N_13979,N_7596,N_8227);
xnor U13980 (N_13980,N_9472,N_5543);
nor U13981 (N_13981,N_6819,N_9900);
nor U13982 (N_13982,N_7869,N_9813);
or U13983 (N_13983,N_6815,N_5812);
nand U13984 (N_13984,N_5394,N_6088);
or U13985 (N_13985,N_8198,N_5067);
or U13986 (N_13986,N_6751,N_9020);
xor U13987 (N_13987,N_8931,N_9975);
nand U13988 (N_13988,N_5468,N_6222);
nor U13989 (N_13989,N_7550,N_8683);
xnor U13990 (N_13990,N_8453,N_9050);
or U13991 (N_13991,N_7794,N_7199);
or U13992 (N_13992,N_7799,N_6081);
xnor U13993 (N_13993,N_9645,N_8519);
and U13994 (N_13994,N_9045,N_9606);
or U13995 (N_13995,N_5690,N_5225);
nand U13996 (N_13996,N_8629,N_9156);
xnor U13997 (N_13997,N_5059,N_9812);
xor U13998 (N_13998,N_8725,N_8554);
nor U13999 (N_13999,N_5901,N_9908);
and U14000 (N_14000,N_9025,N_6958);
or U14001 (N_14001,N_7343,N_9357);
or U14002 (N_14002,N_8068,N_5176);
nor U14003 (N_14003,N_5329,N_6272);
and U14004 (N_14004,N_5573,N_7146);
nand U14005 (N_14005,N_7258,N_5750);
or U14006 (N_14006,N_5749,N_9979);
or U14007 (N_14007,N_8146,N_8722);
xor U14008 (N_14008,N_9398,N_9031);
nand U14009 (N_14009,N_7971,N_6675);
and U14010 (N_14010,N_9187,N_8984);
nand U14011 (N_14011,N_7264,N_5009);
and U14012 (N_14012,N_8786,N_6172);
and U14013 (N_14013,N_9270,N_8347);
and U14014 (N_14014,N_5398,N_5963);
xor U14015 (N_14015,N_6910,N_7962);
and U14016 (N_14016,N_6587,N_6647);
xor U14017 (N_14017,N_8259,N_5518);
nand U14018 (N_14018,N_8716,N_7252);
nor U14019 (N_14019,N_5338,N_7648);
or U14020 (N_14020,N_6241,N_6462);
or U14021 (N_14021,N_8462,N_6148);
or U14022 (N_14022,N_9535,N_8980);
xnor U14023 (N_14023,N_9230,N_9746);
or U14024 (N_14024,N_5158,N_6972);
xnor U14025 (N_14025,N_8017,N_5540);
nor U14026 (N_14026,N_7090,N_5869);
nand U14027 (N_14027,N_5047,N_7677);
and U14028 (N_14028,N_6220,N_7366);
xor U14029 (N_14029,N_9763,N_8312);
nor U14030 (N_14030,N_8084,N_5882);
and U14031 (N_14031,N_6492,N_9804);
nor U14032 (N_14032,N_5523,N_9127);
or U14033 (N_14033,N_8744,N_8677);
and U14034 (N_14034,N_6134,N_8392);
xnor U14035 (N_14035,N_8508,N_8597);
and U14036 (N_14036,N_5660,N_5546);
xnor U14037 (N_14037,N_8022,N_6021);
nand U14038 (N_14038,N_9518,N_5721);
or U14039 (N_14039,N_9718,N_9107);
xor U14040 (N_14040,N_6857,N_9534);
and U14041 (N_14041,N_7063,N_5245);
and U14042 (N_14042,N_6250,N_7695);
nand U14043 (N_14043,N_6921,N_5676);
and U14044 (N_14044,N_7738,N_6291);
or U14045 (N_14045,N_8636,N_5258);
xor U14046 (N_14046,N_7003,N_7884);
and U14047 (N_14047,N_6477,N_9250);
and U14048 (N_14048,N_7281,N_7129);
nor U14049 (N_14049,N_5154,N_8023);
and U14050 (N_14050,N_6472,N_5154);
nand U14051 (N_14051,N_5156,N_7957);
nor U14052 (N_14052,N_7006,N_7433);
nor U14053 (N_14053,N_6630,N_8468);
and U14054 (N_14054,N_5367,N_8400);
and U14055 (N_14055,N_9072,N_9898);
nor U14056 (N_14056,N_5638,N_7416);
or U14057 (N_14057,N_5849,N_9084);
or U14058 (N_14058,N_8735,N_5814);
and U14059 (N_14059,N_9155,N_6076);
nand U14060 (N_14060,N_6702,N_7508);
xnor U14061 (N_14061,N_7815,N_6960);
and U14062 (N_14062,N_6328,N_7150);
xnor U14063 (N_14063,N_7349,N_5687);
xnor U14064 (N_14064,N_6075,N_7805);
xor U14065 (N_14065,N_9691,N_6731);
and U14066 (N_14066,N_7885,N_8241);
or U14067 (N_14067,N_9928,N_9302);
xnor U14068 (N_14068,N_5904,N_7477);
and U14069 (N_14069,N_9166,N_8467);
or U14070 (N_14070,N_5348,N_6014);
nor U14071 (N_14071,N_9568,N_7627);
and U14072 (N_14072,N_8999,N_5439);
nand U14073 (N_14073,N_6129,N_6672);
or U14074 (N_14074,N_7278,N_6280);
nand U14075 (N_14075,N_5662,N_7935);
or U14076 (N_14076,N_6460,N_9115);
nor U14077 (N_14077,N_8610,N_9044);
or U14078 (N_14078,N_5197,N_8881);
nor U14079 (N_14079,N_5342,N_6163);
nand U14080 (N_14080,N_6499,N_9078);
or U14081 (N_14081,N_8488,N_5899);
nor U14082 (N_14082,N_5506,N_9026);
and U14083 (N_14083,N_8796,N_9088);
or U14084 (N_14084,N_9264,N_6406);
nor U14085 (N_14085,N_7157,N_9880);
and U14086 (N_14086,N_7432,N_7732);
xor U14087 (N_14087,N_6869,N_6312);
nand U14088 (N_14088,N_6893,N_9478);
xor U14089 (N_14089,N_8073,N_7150);
and U14090 (N_14090,N_7918,N_9568);
or U14091 (N_14091,N_5915,N_8201);
and U14092 (N_14092,N_8291,N_9323);
nor U14093 (N_14093,N_9567,N_7832);
xor U14094 (N_14094,N_9965,N_8744);
nor U14095 (N_14095,N_5638,N_8170);
or U14096 (N_14096,N_9445,N_7263);
or U14097 (N_14097,N_7595,N_7439);
xnor U14098 (N_14098,N_8289,N_6219);
nand U14099 (N_14099,N_8203,N_9223);
nor U14100 (N_14100,N_6600,N_8755);
xor U14101 (N_14101,N_8747,N_9211);
or U14102 (N_14102,N_7688,N_8891);
or U14103 (N_14103,N_6846,N_6003);
nand U14104 (N_14104,N_8601,N_6144);
nor U14105 (N_14105,N_6319,N_6072);
nand U14106 (N_14106,N_8679,N_8301);
nor U14107 (N_14107,N_6239,N_8959);
nor U14108 (N_14108,N_6214,N_9602);
nand U14109 (N_14109,N_7242,N_9683);
nand U14110 (N_14110,N_6120,N_5542);
and U14111 (N_14111,N_9442,N_9630);
xor U14112 (N_14112,N_7747,N_6306);
nor U14113 (N_14113,N_5239,N_7821);
nand U14114 (N_14114,N_6986,N_6450);
nand U14115 (N_14115,N_6510,N_8830);
xnor U14116 (N_14116,N_9981,N_8865);
or U14117 (N_14117,N_7455,N_9306);
or U14118 (N_14118,N_5184,N_9180);
or U14119 (N_14119,N_7615,N_9217);
nand U14120 (N_14120,N_6156,N_5709);
or U14121 (N_14121,N_5517,N_7090);
nand U14122 (N_14122,N_5542,N_7719);
and U14123 (N_14123,N_8630,N_9485);
nor U14124 (N_14124,N_7224,N_7633);
or U14125 (N_14125,N_9151,N_5546);
nor U14126 (N_14126,N_6214,N_6332);
or U14127 (N_14127,N_5605,N_6807);
or U14128 (N_14128,N_7881,N_8628);
xnor U14129 (N_14129,N_5356,N_8735);
and U14130 (N_14130,N_5193,N_7080);
and U14131 (N_14131,N_6636,N_7453);
and U14132 (N_14132,N_7706,N_9662);
and U14133 (N_14133,N_5803,N_8532);
or U14134 (N_14134,N_9513,N_7873);
xnor U14135 (N_14135,N_5143,N_5107);
xnor U14136 (N_14136,N_8204,N_6824);
and U14137 (N_14137,N_9397,N_6090);
or U14138 (N_14138,N_6272,N_9072);
nand U14139 (N_14139,N_8094,N_9327);
or U14140 (N_14140,N_8483,N_8096);
nor U14141 (N_14141,N_9973,N_6847);
or U14142 (N_14142,N_6306,N_8934);
and U14143 (N_14143,N_9011,N_7585);
and U14144 (N_14144,N_8572,N_6034);
nand U14145 (N_14145,N_6893,N_7604);
nor U14146 (N_14146,N_6008,N_7765);
nand U14147 (N_14147,N_7535,N_9450);
nor U14148 (N_14148,N_9286,N_7396);
or U14149 (N_14149,N_5954,N_8448);
nor U14150 (N_14150,N_5462,N_9760);
nand U14151 (N_14151,N_9533,N_7576);
xnor U14152 (N_14152,N_9504,N_6148);
xor U14153 (N_14153,N_8693,N_6183);
nand U14154 (N_14154,N_8655,N_8552);
nor U14155 (N_14155,N_8637,N_8264);
or U14156 (N_14156,N_6108,N_7259);
nor U14157 (N_14157,N_5221,N_8156);
xnor U14158 (N_14158,N_6202,N_8734);
or U14159 (N_14159,N_6579,N_8041);
or U14160 (N_14160,N_9415,N_6803);
nand U14161 (N_14161,N_8578,N_9475);
nand U14162 (N_14162,N_6620,N_8596);
nor U14163 (N_14163,N_6385,N_9479);
or U14164 (N_14164,N_8315,N_9095);
nor U14165 (N_14165,N_8110,N_5514);
nand U14166 (N_14166,N_7419,N_9282);
or U14167 (N_14167,N_9905,N_9634);
nor U14168 (N_14168,N_7284,N_8626);
and U14169 (N_14169,N_7761,N_7514);
nor U14170 (N_14170,N_5469,N_6112);
and U14171 (N_14171,N_5261,N_7563);
and U14172 (N_14172,N_7371,N_5628);
nor U14173 (N_14173,N_5711,N_8631);
xor U14174 (N_14174,N_8819,N_6351);
or U14175 (N_14175,N_7267,N_5710);
nand U14176 (N_14176,N_8452,N_8851);
nand U14177 (N_14177,N_6831,N_7174);
and U14178 (N_14178,N_7343,N_9962);
or U14179 (N_14179,N_7246,N_9314);
nand U14180 (N_14180,N_9488,N_7356);
and U14181 (N_14181,N_6901,N_8065);
xor U14182 (N_14182,N_9313,N_6813);
nor U14183 (N_14183,N_8029,N_8049);
nand U14184 (N_14184,N_8446,N_9307);
xnor U14185 (N_14185,N_7118,N_6827);
xor U14186 (N_14186,N_5675,N_5681);
and U14187 (N_14187,N_8366,N_9836);
xnor U14188 (N_14188,N_6762,N_8631);
nand U14189 (N_14189,N_8663,N_5407);
nand U14190 (N_14190,N_7747,N_7502);
or U14191 (N_14191,N_7957,N_7068);
nand U14192 (N_14192,N_7469,N_9379);
nor U14193 (N_14193,N_8631,N_7634);
or U14194 (N_14194,N_9639,N_7001);
nor U14195 (N_14195,N_7928,N_9522);
xor U14196 (N_14196,N_7363,N_7698);
nand U14197 (N_14197,N_7000,N_7296);
and U14198 (N_14198,N_6272,N_5698);
xnor U14199 (N_14199,N_8445,N_7660);
nor U14200 (N_14200,N_7660,N_7586);
or U14201 (N_14201,N_7478,N_6256);
or U14202 (N_14202,N_6549,N_6383);
nand U14203 (N_14203,N_8194,N_8710);
nand U14204 (N_14204,N_8647,N_6990);
nand U14205 (N_14205,N_7702,N_8999);
or U14206 (N_14206,N_6036,N_5827);
or U14207 (N_14207,N_5891,N_7548);
nor U14208 (N_14208,N_7364,N_8352);
xor U14209 (N_14209,N_6332,N_8349);
nor U14210 (N_14210,N_9073,N_5302);
or U14211 (N_14211,N_8590,N_6721);
or U14212 (N_14212,N_7749,N_8146);
xor U14213 (N_14213,N_5355,N_9054);
nand U14214 (N_14214,N_6452,N_6325);
and U14215 (N_14215,N_6230,N_9301);
and U14216 (N_14216,N_8033,N_7184);
or U14217 (N_14217,N_7782,N_7430);
nand U14218 (N_14218,N_9555,N_8618);
nand U14219 (N_14219,N_9456,N_6061);
and U14220 (N_14220,N_6690,N_6965);
xor U14221 (N_14221,N_5991,N_8373);
nor U14222 (N_14222,N_9372,N_5773);
nor U14223 (N_14223,N_9248,N_6478);
xor U14224 (N_14224,N_9862,N_8509);
nor U14225 (N_14225,N_8821,N_9357);
xnor U14226 (N_14226,N_9587,N_9399);
xor U14227 (N_14227,N_5944,N_5006);
or U14228 (N_14228,N_7479,N_8035);
and U14229 (N_14229,N_9141,N_6033);
or U14230 (N_14230,N_9001,N_9156);
or U14231 (N_14231,N_9167,N_7334);
and U14232 (N_14232,N_6948,N_9387);
and U14233 (N_14233,N_9853,N_8214);
or U14234 (N_14234,N_5216,N_7751);
nand U14235 (N_14235,N_5767,N_9496);
or U14236 (N_14236,N_5638,N_9859);
xor U14237 (N_14237,N_5588,N_9736);
xnor U14238 (N_14238,N_7270,N_7371);
xor U14239 (N_14239,N_6490,N_9710);
or U14240 (N_14240,N_5905,N_8455);
and U14241 (N_14241,N_5562,N_5393);
xnor U14242 (N_14242,N_7888,N_9247);
and U14243 (N_14243,N_9794,N_5243);
and U14244 (N_14244,N_7845,N_7764);
nand U14245 (N_14245,N_6978,N_6385);
xor U14246 (N_14246,N_5814,N_8412);
and U14247 (N_14247,N_5570,N_7918);
xnor U14248 (N_14248,N_8976,N_7860);
and U14249 (N_14249,N_6701,N_6118);
nor U14250 (N_14250,N_6744,N_5790);
or U14251 (N_14251,N_9166,N_7743);
or U14252 (N_14252,N_5493,N_5832);
xnor U14253 (N_14253,N_8453,N_7731);
or U14254 (N_14254,N_9798,N_6436);
xnor U14255 (N_14255,N_8904,N_5156);
nor U14256 (N_14256,N_5742,N_5435);
xnor U14257 (N_14257,N_9632,N_8354);
nand U14258 (N_14258,N_9962,N_8437);
and U14259 (N_14259,N_9543,N_9557);
nor U14260 (N_14260,N_6118,N_6206);
nand U14261 (N_14261,N_8835,N_9098);
and U14262 (N_14262,N_7054,N_5678);
nor U14263 (N_14263,N_8943,N_9363);
nor U14264 (N_14264,N_6020,N_6500);
and U14265 (N_14265,N_8300,N_5737);
or U14266 (N_14266,N_6532,N_6424);
xor U14267 (N_14267,N_9236,N_8753);
nand U14268 (N_14268,N_6119,N_5744);
nor U14269 (N_14269,N_8811,N_8424);
nand U14270 (N_14270,N_7872,N_8658);
xnor U14271 (N_14271,N_5129,N_6060);
nor U14272 (N_14272,N_8978,N_5519);
or U14273 (N_14273,N_9306,N_9435);
xor U14274 (N_14274,N_6963,N_7375);
or U14275 (N_14275,N_7377,N_6609);
nand U14276 (N_14276,N_7111,N_9275);
nor U14277 (N_14277,N_8145,N_5458);
nor U14278 (N_14278,N_8385,N_6383);
nor U14279 (N_14279,N_8798,N_6293);
xnor U14280 (N_14280,N_8752,N_9536);
xnor U14281 (N_14281,N_8468,N_7794);
nand U14282 (N_14282,N_9329,N_9356);
or U14283 (N_14283,N_9454,N_7028);
nand U14284 (N_14284,N_8322,N_7249);
nand U14285 (N_14285,N_8668,N_8618);
and U14286 (N_14286,N_8784,N_8089);
nand U14287 (N_14287,N_9618,N_7612);
xor U14288 (N_14288,N_9640,N_7149);
and U14289 (N_14289,N_6824,N_7601);
nand U14290 (N_14290,N_8833,N_7749);
or U14291 (N_14291,N_5339,N_8326);
nand U14292 (N_14292,N_9937,N_5897);
nand U14293 (N_14293,N_7244,N_6922);
nand U14294 (N_14294,N_8587,N_5515);
and U14295 (N_14295,N_6574,N_8004);
or U14296 (N_14296,N_6680,N_9686);
nand U14297 (N_14297,N_8822,N_5305);
nand U14298 (N_14298,N_8404,N_7670);
or U14299 (N_14299,N_9843,N_8322);
nor U14300 (N_14300,N_8374,N_9350);
nor U14301 (N_14301,N_8144,N_7250);
nand U14302 (N_14302,N_8934,N_5994);
nand U14303 (N_14303,N_7774,N_5719);
and U14304 (N_14304,N_9538,N_9074);
xor U14305 (N_14305,N_8913,N_5866);
nor U14306 (N_14306,N_6272,N_5721);
or U14307 (N_14307,N_9822,N_5354);
nand U14308 (N_14308,N_6068,N_6982);
and U14309 (N_14309,N_5911,N_6394);
xnor U14310 (N_14310,N_6257,N_6251);
nand U14311 (N_14311,N_5201,N_9824);
nand U14312 (N_14312,N_5418,N_8534);
nor U14313 (N_14313,N_8022,N_5014);
and U14314 (N_14314,N_6397,N_7403);
nor U14315 (N_14315,N_9183,N_6074);
nor U14316 (N_14316,N_6141,N_8603);
nor U14317 (N_14317,N_8573,N_7960);
or U14318 (N_14318,N_7051,N_6903);
nor U14319 (N_14319,N_6170,N_9511);
and U14320 (N_14320,N_7403,N_5377);
nand U14321 (N_14321,N_6396,N_9477);
or U14322 (N_14322,N_5375,N_5299);
nand U14323 (N_14323,N_6580,N_5711);
nand U14324 (N_14324,N_6228,N_6829);
nand U14325 (N_14325,N_6592,N_7543);
or U14326 (N_14326,N_6518,N_5319);
and U14327 (N_14327,N_7219,N_5847);
nor U14328 (N_14328,N_6280,N_9161);
nor U14329 (N_14329,N_5688,N_6731);
nor U14330 (N_14330,N_7298,N_7842);
nand U14331 (N_14331,N_5609,N_5352);
and U14332 (N_14332,N_9196,N_8962);
nor U14333 (N_14333,N_5595,N_5954);
and U14334 (N_14334,N_7533,N_6939);
nand U14335 (N_14335,N_9823,N_5559);
nand U14336 (N_14336,N_8518,N_8243);
and U14337 (N_14337,N_9437,N_6228);
nand U14338 (N_14338,N_6550,N_9451);
nand U14339 (N_14339,N_5790,N_7422);
nor U14340 (N_14340,N_6448,N_5054);
xnor U14341 (N_14341,N_7882,N_7045);
nand U14342 (N_14342,N_5878,N_9368);
and U14343 (N_14343,N_5048,N_6135);
nor U14344 (N_14344,N_6795,N_7523);
nor U14345 (N_14345,N_6356,N_5746);
or U14346 (N_14346,N_7400,N_9597);
nor U14347 (N_14347,N_6812,N_5927);
nand U14348 (N_14348,N_7349,N_9191);
or U14349 (N_14349,N_7603,N_9141);
xor U14350 (N_14350,N_9701,N_7310);
or U14351 (N_14351,N_8231,N_5764);
and U14352 (N_14352,N_8116,N_9931);
xor U14353 (N_14353,N_8804,N_7239);
nand U14354 (N_14354,N_9010,N_6878);
nand U14355 (N_14355,N_8066,N_6382);
xnor U14356 (N_14356,N_9020,N_9610);
nor U14357 (N_14357,N_6567,N_8004);
xor U14358 (N_14358,N_7779,N_6946);
nand U14359 (N_14359,N_7798,N_5286);
and U14360 (N_14360,N_5046,N_6592);
xor U14361 (N_14361,N_9293,N_8969);
and U14362 (N_14362,N_9280,N_7452);
nand U14363 (N_14363,N_7023,N_7439);
nor U14364 (N_14364,N_8721,N_7636);
or U14365 (N_14365,N_6080,N_6863);
nor U14366 (N_14366,N_7977,N_6291);
or U14367 (N_14367,N_9266,N_5007);
or U14368 (N_14368,N_6208,N_5401);
nor U14369 (N_14369,N_6761,N_6950);
and U14370 (N_14370,N_7543,N_9536);
or U14371 (N_14371,N_9783,N_8436);
or U14372 (N_14372,N_8531,N_6184);
xnor U14373 (N_14373,N_9959,N_8027);
xnor U14374 (N_14374,N_5015,N_7759);
or U14375 (N_14375,N_5715,N_8965);
and U14376 (N_14376,N_7226,N_7282);
and U14377 (N_14377,N_6681,N_9254);
nand U14378 (N_14378,N_9698,N_7378);
nor U14379 (N_14379,N_8152,N_6628);
nor U14380 (N_14380,N_8792,N_7094);
nand U14381 (N_14381,N_7181,N_9871);
or U14382 (N_14382,N_8934,N_6448);
and U14383 (N_14383,N_5981,N_8214);
or U14384 (N_14384,N_9848,N_7021);
xor U14385 (N_14385,N_9783,N_6127);
nor U14386 (N_14386,N_5206,N_8165);
nand U14387 (N_14387,N_7828,N_7944);
nand U14388 (N_14388,N_5621,N_6121);
and U14389 (N_14389,N_6694,N_6760);
and U14390 (N_14390,N_9174,N_9299);
nor U14391 (N_14391,N_9356,N_5185);
nand U14392 (N_14392,N_9634,N_8262);
nor U14393 (N_14393,N_6210,N_6442);
nor U14394 (N_14394,N_5331,N_5002);
xor U14395 (N_14395,N_8287,N_7476);
nand U14396 (N_14396,N_7417,N_5160);
nor U14397 (N_14397,N_5504,N_9174);
or U14398 (N_14398,N_7246,N_7404);
nand U14399 (N_14399,N_5622,N_7313);
and U14400 (N_14400,N_9713,N_9714);
or U14401 (N_14401,N_8446,N_8934);
nor U14402 (N_14402,N_9468,N_5177);
and U14403 (N_14403,N_6337,N_7458);
xnor U14404 (N_14404,N_9520,N_5177);
xnor U14405 (N_14405,N_6374,N_8709);
and U14406 (N_14406,N_7420,N_5102);
and U14407 (N_14407,N_5576,N_7279);
xnor U14408 (N_14408,N_5886,N_5426);
xnor U14409 (N_14409,N_6042,N_6583);
nor U14410 (N_14410,N_7596,N_5405);
and U14411 (N_14411,N_6252,N_7417);
xor U14412 (N_14412,N_5175,N_9911);
xor U14413 (N_14413,N_6359,N_7126);
and U14414 (N_14414,N_7280,N_6208);
nand U14415 (N_14415,N_7627,N_8960);
nor U14416 (N_14416,N_7587,N_8316);
and U14417 (N_14417,N_8056,N_8001);
and U14418 (N_14418,N_6631,N_8478);
or U14419 (N_14419,N_7023,N_7529);
nand U14420 (N_14420,N_5642,N_6502);
nor U14421 (N_14421,N_9181,N_9052);
xor U14422 (N_14422,N_9705,N_6962);
or U14423 (N_14423,N_5697,N_9596);
or U14424 (N_14424,N_8325,N_9891);
xnor U14425 (N_14425,N_7103,N_8060);
nor U14426 (N_14426,N_8857,N_9150);
nor U14427 (N_14427,N_6040,N_5651);
or U14428 (N_14428,N_6012,N_9343);
and U14429 (N_14429,N_8632,N_7197);
nand U14430 (N_14430,N_8264,N_9525);
and U14431 (N_14431,N_6286,N_8416);
or U14432 (N_14432,N_5765,N_8387);
or U14433 (N_14433,N_8389,N_8668);
nor U14434 (N_14434,N_9232,N_6791);
nor U14435 (N_14435,N_8822,N_6737);
or U14436 (N_14436,N_5957,N_7195);
and U14437 (N_14437,N_7604,N_7961);
or U14438 (N_14438,N_8125,N_9564);
and U14439 (N_14439,N_5766,N_6347);
or U14440 (N_14440,N_5265,N_9630);
or U14441 (N_14441,N_6625,N_7161);
and U14442 (N_14442,N_8259,N_5092);
nand U14443 (N_14443,N_6114,N_5653);
and U14444 (N_14444,N_5565,N_8773);
xor U14445 (N_14445,N_6516,N_7297);
nor U14446 (N_14446,N_7214,N_6845);
nor U14447 (N_14447,N_7543,N_6815);
nand U14448 (N_14448,N_9279,N_9364);
or U14449 (N_14449,N_9824,N_5488);
or U14450 (N_14450,N_6290,N_5488);
and U14451 (N_14451,N_9453,N_8869);
or U14452 (N_14452,N_7499,N_5871);
nor U14453 (N_14453,N_9531,N_5692);
nor U14454 (N_14454,N_6144,N_5455);
nor U14455 (N_14455,N_8959,N_7515);
nor U14456 (N_14456,N_7360,N_7846);
nor U14457 (N_14457,N_8703,N_6685);
or U14458 (N_14458,N_9091,N_6029);
and U14459 (N_14459,N_6953,N_9376);
nand U14460 (N_14460,N_6175,N_9052);
xor U14461 (N_14461,N_7428,N_5980);
or U14462 (N_14462,N_9840,N_8163);
nand U14463 (N_14463,N_7332,N_8602);
or U14464 (N_14464,N_7409,N_9817);
nand U14465 (N_14465,N_9159,N_6030);
xnor U14466 (N_14466,N_8230,N_9072);
or U14467 (N_14467,N_9699,N_7594);
xnor U14468 (N_14468,N_7353,N_9810);
xnor U14469 (N_14469,N_9861,N_7395);
nand U14470 (N_14470,N_7357,N_6722);
and U14471 (N_14471,N_9438,N_7970);
and U14472 (N_14472,N_9141,N_7987);
xnor U14473 (N_14473,N_8333,N_9169);
xor U14474 (N_14474,N_6440,N_6444);
nor U14475 (N_14475,N_6576,N_8657);
or U14476 (N_14476,N_6319,N_8652);
xnor U14477 (N_14477,N_7614,N_9116);
and U14478 (N_14478,N_7144,N_9303);
xnor U14479 (N_14479,N_5056,N_5124);
and U14480 (N_14480,N_5771,N_5247);
and U14481 (N_14481,N_6801,N_6382);
or U14482 (N_14482,N_5996,N_5181);
xor U14483 (N_14483,N_9493,N_7709);
nand U14484 (N_14484,N_7133,N_6697);
or U14485 (N_14485,N_7555,N_5381);
or U14486 (N_14486,N_8487,N_5056);
nand U14487 (N_14487,N_8444,N_7907);
nor U14488 (N_14488,N_9576,N_7620);
nor U14489 (N_14489,N_7307,N_5854);
xnor U14490 (N_14490,N_8977,N_9657);
nor U14491 (N_14491,N_9756,N_6003);
nor U14492 (N_14492,N_8910,N_5956);
nand U14493 (N_14493,N_8591,N_8876);
xor U14494 (N_14494,N_5749,N_8112);
or U14495 (N_14495,N_5109,N_7865);
nor U14496 (N_14496,N_8377,N_6519);
and U14497 (N_14497,N_8396,N_8845);
nand U14498 (N_14498,N_6347,N_9941);
nand U14499 (N_14499,N_5398,N_7726);
or U14500 (N_14500,N_8024,N_9220);
and U14501 (N_14501,N_9535,N_9717);
and U14502 (N_14502,N_7245,N_9417);
xnor U14503 (N_14503,N_7837,N_5580);
or U14504 (N_14504,N_8239,N_6094);
nor U14505 (N_14505,N_9773,N_8937);
xnor U14506 (N_14506,N_7800,N_7509);
or U14507 (N_14507,N_8253,N_5381);
or U14508 (N_14508,N_9426,N_8764);
and U14509 (N_14509,N_8600,N_5448);
nor U14510 (N_14510,N_8394,N_9338);
nor U14511 (N_14511,N_6727,N_9057);
and U14512 (N_14512,N_8036,N_9443);
xnor U14513 (N_14513,N_7377,N_8537);
and U14514 (N_14514,N_8765,N_9330);
xor U14515 (N_14515,N_8948,N_7504);
xor U14516 (N_14516,N_5958,N_8345);
nor U14517 (N_14517,N_9482,N_8673);
or U14518 (N_14518,N_5156,N_5326);
nor U14519 (N_14519,N_6061,N_7873);
or U14520 (N_14520,N_6255,N_6538);
or U14521 (N_14521,N_9189,N_5165);
or U14522 (N_14522,N_9696,N_8809);
xnor U14523 (N_14523,N_5778,N_7164);
nor U14524 (N_14524,N_9261,N_6145);
xor U14525 (N_14525,N_8336,N_8504);
or U14526 (N_14526,N_6038,N_9247);
nand U14527 (N_14527,N_9861,N_8720);
nand U14528 (N_14528,N_9044,N_8801);
nor U14529 (N_14529,N_7823,N_8425);
nor U14530 (N_14530,N_6764,N_5176);
nand U14531 (N_14531,N_5400,N_6257);
nor U14532 (N_14532,N_8782,N_8063);
xnor U14533 (N_14533,N_8397,N_8536);
and U14534 (N_14534,N_5638,N_9516);
nor U14535 (N_14535,N_6825,N_7006);
and U14536 (N_14536,N_5311,N_5817);
and U14537 (N_14537,N_8068,N_8445);
xor U14538 (N_14538,N_7635,N_7395);
nor U14539 (N_14539,N_9946,N_7837);
nand U14540 (N_14540,N_6907,N_6556);
nand U14541 (N_14541,N_8027,N_5855);
nand U14542 (N_14542,N_7341,N_6389);
or U14543 (N_14543,N_9678,N_7837);
or U14544 (N_14544,N_5410,N_9652);
and U14545 (N_14545,N_7796,N_7915);
nor U14546 (N_14546,N_9975,N_5480);
nor U14547 (N_14547,N_6138,N_8205);
nor U14548 (N_14548,N_8702,N_6359);
or U14549 (N_14549,N_6046,N_8731);
or U14550 (N_14550,N_6460,N_5450);
or U14551 (N_14551,N_8013,N_7269);
and U14552 (N_14552,N_8086,N_9694);
nor U14553 (N_14553,N_5251,N_8964);
and U14554 (N_14554,N_6917,N_6651);
nor U14555 (N_14555,N_8439,N_6969);
and U14556 (N_14556,N_5565,N_7805);
nor U14557 (N_14557,N_7400,N_7477);
or U14558 (N_14558,N_8041,N_9103);
nor U14559 (N_14559,N_5339,N_9725);
or U14560 (N_14560,N_5792,N_5529);
and U14561 (N_14561,N_6315,N_6358);
or U14562 (N_14562,N_9561,N_9729);
and U14563 (N_14563,N_9362,N_7793);
or U14564 (N_14564,N_9295,N_5979);
and U14565 (N_14565,N_5030,N_9819);
and U14566 (N_14566,N_9389,N_6307);
and U14567 (N_14567,N_6484,N_5789);
nand U14568 (N_14568,N_5497,N_8474);
nor U14569 (N_14569,N_6852,N_6255);
xnor U14570 (N_14570,N_8057,N_6232);
nor U14571 (N_14571,N_9659,N_9182);
and U14572 (N_14572,N_7324,N_6457);
or U14573 (N_14573,N_7471,N_5065);
and U14574 (N_14574,N_7691,N_9380);
nand U14575 (N_14575,N_8529,N_9373);
and U14576 (N_14576,N_6848,N_9413);
nand U14577 (N_14577,N_6943,N_8793);
xnor U14578 (N_14578,N_7027,N_7311);
or U14579 (N_14579,N_8690,N_9968);
xor U14580 (N_14580,N_5774,N_6942);
or U14581 (N_14581,N_5327,N_8294);
and U14582 (N_14582,N_9748,N_5125);
nand U14583 (N_14583,N_7896,N_5553);
xnor U14584 (N_14584,N_6712,N_8043);
nand U14585 (N_14585,N_6761,N_6915);
xor U14586 (N_14586,N_5704,N_6974);
xnor U14587 (N_14587,N_8161,N_6173);
xor U14588 (N_14588,N_9102,N_9424);
nor U14589 (N_14589,N_8954,N_8970);
xor U14590 (N_14590,N_6150,N_6745);
and U14591 (N_14591,N_6980,N_7119);
nor U14592 (N_14592,N_7444,N_8044);
and U14593 (N_14593,N_5341,N_7617);
nor U14594 (N_14594,N_7115,N_5557);
and U14595 (N_14595,N_6381,N_9823);
xnor U14596 (N_14596,N_9997,N_7475);
or U14597 (N_14597,N_7078,N_9601);
xor U14598 (N_14598,N_9831,N_8752);
nand U14599 (N_14599,N_5635,N_8496);
and U14600 (N_14600,N_7211,N_9201);
or U14601 (N_14601,N_9532,N_9612);
xor U14602 (N_14602,N_7879,N_6262);
nand U14603 (N_14603,N_5894,N_9495);
and U14604 (N_14604,N_9727,N_8533);
nand U14605 (N_14605,N_7963,N_9735);
or U14606 (N_14606,N_7218,N_6025);
nor U14607 (N_14607,N_6688,N_7669);
nand U14608 (N_14608,N_6832,N_9398);
xnor U14609 (N_14609,N_9447,N_9212);
or U14610 (N_14610,N_5998,N_5434);
or U14611 (N_14611,N_9727,N_6719);
xor U14612 (N_14612,N_6463,N_5197);
xor U14613 (N_14613,N_5283,N_9727);
nor U14614 (N_14614,N_9050,N_6761);
or U14615 (N_14615,N_9503,N_6427);
or U14616 (N_14616,N_9192,N_6631);
or U14617 (N_14617,N_5987,N_6115);
or U14618 (N_14618,N_9416,N_8435);
nor U14619 (N_14619,N_5543,N_6429);
nand U14620 (N_14620,N_6780,N_9904);
or U14621 (N_14621,N_9734,N_8893);
xor U14622 (N_14622,N_5062,N_7630);
nand U14623 (N_14623,N_6348,N_5594);
and U14624 (N_14624,N_6847,N_8526);
xor U14625 (N_14625,N_9834,N_5834);
or U14626 (N_14626,N_8076,N_5083);
nor U14627 (N_14627,N_5610,N_6121);
xor U14628 (N_14628,N_8261,N_5824);
xor U14629 (N_14629,N_6627,N_8167);
nand U14630 (N_14630,N_9589,N_8087);
xnor U14631 (N_14631,N_8879,N_5122);
and U14632 (N_14632,N_7833,N_5274);
nor U14633 (N_14633,N_6268,N_5081);
nor U14634 (N_14634,N_7245,N_5017);
xnor U14635 (N_14635,N_8088,N_9136);
nand U14636 (N_14636,N_9625,N_9701);
or U14637 (N_14637,N_5666,N_9937);
nand U14638 (N_14638,N_6103,N_9047);
or U14639 (N_14639,N_7786,N_7867);
xor U14640 (N_14640,N_7540,N_5372);
xnor U14641 (N_14641,N_9657,N_6894);
and U14642 (N_14642,N_8327,N_5616);
or U14643 (N_14643,N_7001,N_5890);
nor U14644 (N_14644,N_8136,N_5815);
nor U14645 (N_14645,N_6802,N_5493);
nor U14646 (N_14646,N_8679,N_8994);
and U14647 (N_14647,N_5477,N_5584);
or U14648 (N_14648,N_6079,N_6900);
nand U14649 (N_14649,N_8581,N_7790);
and U14650 (N_14650,N_6294,N_6581);
nor U14651 (N_14651,N_5025,N_9969);
nor U14652 (N_14652,N_6780,N_5164);
or U14653 (N_14653,N_7848,N_8667);
nand U14654 (N_14654,N_8713,N_5250);
nor U14655 (N_14655,N_8874,N_5044);
nor U14656 (N_14656,N_8124,N_7988);
nor U14657 (N_14657,N_6530,N_9595);
nand U14658 (N_14658,N_7328,N_5969);
xor U14659 (N_14659,N_5761,N_9222);
nor U14660 (N_14660,N_6990,N_8224);
nor U14661 (N_14661,N_5700,N_5619);
nand U14662 (N_14662,N_6899,N_7535);
nand U14663 (N_14663,N_7995,N_5527);
and U14664 (N_14664,N_5157,N_7747);
nand U14665 (N_14665,N_7482,N_8629);
or U14666 (N_14666,N_6232,N_8749);
nor U14667 (N_14667,N_9296,N_7799);
nand U14668 (N_14668,N_8241,N_6913);
nor U14669 (N_14669,N_8376,N_6882);
xor U14670 (N_14670,N_5831,N_5862);
nor U14671 (N_14671,N_7381,N_9879);
nand U14672 (N_14672,N_5471,N_8773);
nor U14673 (N_14673,N_6865,N_8300);
or U14674 (N_14674,N_9517,N_9855);
xor U14675 (N_14675,N_9978,N_9845);
and U14676 (N_14676,N_9462,N_7352);
and U14677 (N_14677,N_8741,N_7378);
xnor U14678 (N_14678,N_7717,N_7140);
nand U14679 (N_14679,N_8377,N_6515);
xnor U14680 (N_14680,N_6103,N_7073);
or U14681 (N_14681,N_9741,N_9958);
and U14682 (N_14682,N_6483,N_9520);
nand U14683 (N_14683,N_6649,N_5595);
nor U14684 (N_14684,N_8253,N_8881);
nor U14685 (N_14685,N_6695,N_8962);
xor U14686 (N_14686,N_8821,N_5115);
xor U14687 (N_14687,N_5644,N_8949);
or U14688 (N_14688,N_7268,N_6938);
nor U14689 (N_14689,N_5446,N_5250);
and U14690 (N_14690,N_9310,N_5005);
or U14691 (N_14691,N_8391,N_6547);
or U14692 (N_14692,N_6530,N_9594);
and U14693 (N_14693,N_5621,N_9662);
and U14694 (N_14694,N_6080,N_9265);
or U14695 (N_14695,N_8820,N_7616);
and U14696 (N_14696,N_5666,N_9526);
or U14697 (N_14697,N_7142,N_6643);
or U14698 (N_14698,N_5150,N_9162);
and U14699 (N_14699,N_8248,N_5245);
nand U14700 (N_14700,N_5509,N_6169);
nor U14701 (N_14701,N_5543,N_8577);
nand U14702 (N_14702,N_5190,N_9761);
and U14703 (N_14703,N_6090,N_8255);
nand U14704 (N_14704,N_6321,N_6986);
nor U14705 (N_14705,N_6402,N_8815);
nand U14706 (N_14706,N_7524,N_6963);
and U14707 (N_14707,N_7880,N_7372);
nand U14708 (N_14708,N_8972,N_6480);
and U14709 (N_14709,N_8210,N_5670);
or U14710 (N_14710,N_7641,N_5121);
xor U14711 (N_14711,N_9459,N_7960);
nor U14712 (N_14712,N_5584,N_6334);
xor U14713 (N_14713,N_9258,N_9622);
or U14714 (N_14714,N_7819,N_9361);
xnor U14715 (N_14715,N_5274,N_5107);
and U14716 (N_14716,N_6808,N_6305);
and U14717 (N_14717,N_7531,N_9596);
xnor U14718 (N_14718,N_5455,N_9510);
or U14719 (N_14719,N_5798,N_5614);
and U14720 (N_14720,N_8623,N_5622);
xnor U14721 (N_14721,N_5838,N_9792);
or U14722 (N_14722,N_7191,N_5402);
nand U14723 (N_14723,N_8039,N_9460);
xor U14724 (N_14724,N_7208,N_8954);
nand U14725 (N_14725,N_9165,N_6692);
nor U14726 (N_14726,N_9858,N_7802);
and U14727 (N_14727,N_6911,N_5855);
nor U14728 (N_14728,N_8166,N_6578);
or U14729 (N_14729,N_8142,N_9364);
nand U14730 (N_14730,N_7419,N_8287);
nand U14731 (N_14731,N_5637,N_7630);
nor U14732 (N_14732,N_5401,N_8097);
and U14733 (N_14733,N_6365,N_8613);
xor U14734 (N_14734,N_7065,N_9093);
or U14735 (N_14735,N_5119,N_6434);
or U14736 (N_14736,N_5926,N_8328);
and U14737 (N_14737,N_7814,N_8634);
and U14738 (N_14738,N_9370,N_9505);
or U14739 (N_14739,N_9166,N_5046);
nand U14740 (N_14740,N_8438,N_7385);
or U14741 (N_14741,N_5364,N_9827);
or U14742 (N_14742,N_5535,N_7950);
xnor U14743 (N_14743,N_5189,N_5039);
nor U14744 (N_14744,N_5173,N_7942);
xnor U14745 (N_14745,N_6669,N_5202);
nor U14746 (N_14746,N_8422,N_5663);
and U14747 (N_14747,N_7036,N_6806);
nand U14748 (N_14748,N_5451,N_6301);
and U14749 (N_14749,N_6241,N_7535);
and U14750 (N_14750,N_5452,N_6272);
nor U14751 (N_14751,N_6821,N_6593);
nor U14752 (N_14752,N_5891,N_6652);
and U14753 (N_14753,N_7912,N_5756);
xnor U14754 (N_14754,N_7908,N_6344);
xnor U14755 (N_14755,N_7553,N_5558);
nand U14756 (N_14756,N_5637,N_6510);
or U14757 (N_14757,N_6556,N_6134);
or U14758 (N_14758,N_5084,N_7036);
or U14759 (N_14759,N_9127,N_6218);
and U14760 (N_14760,N_9653,N_5891);
or U14761 (N_14761,N_8413,N_6827);
nor U14762 (N_14762,N_5421,N_8037);
nor U14763 (N_14763,N_7479,N_8946);
or U14764 (N_14764,N_8447,N_6476);
nand U14765 (N_14765,N_8014,N_7682);
nor U14766 (N_14766,N_8340,N_9815);
nand U14767 (N_14767,N_9039,N_8010);
xor U14768 (N_14768,N_5400,N_8250);
and U14769 (N_14769,N_7740,N_8702);
nor U14770 (N_14770,N_9378,N_9097);
and U14771 (N_14771,N_8744,N_7874);
nor U14772 (N_14772,N_9779,N_6890);
nand U14773 (N_14773,N_5814,N_7293);
or U14774 (N_14774,N_9492,N_5549);
and U14775 (N_14775,N_9329,N_9198);
nand U14776 (N_14776,N_8367,N_5738);
nor U14777 (N_14777,N_8283,N_9406);
and U14778 (N_14778,N_5046,N_5368);
and U14779 (N_14779,N_5561,N_9263);
or U14780 (N_14780,N_9386,N_5513);
and U14781 (N_14781,N_9844,N_7988);
and U14782 (N_14782,N_5540,N_5522);
or U14783 (N_14783,N_5955,N_9039);
nand U14784 (N_14784,N_9487,N_6270);
xnor U14785 (N_14785,N_5103,N_6319);
nand U14786 (N_14786,N_5885,N_7783);
nor U14787 (N_14787,N_7926,N_5010);
xor U14788 (N_14788,N_6835,N_7633);
nor U14789 (N_14789,N_9038,N_5953);
xnor U14790 (N_14790,N_7343,N_6939);
or U14791 (N_14791,N_9373,N_6691);
or U14792 (N_14792,N_5212,N_6236);
xor U14793 (N_14793,N_5967,N_8712);
or U14794 (N_14794,N_8633,N_8202);
nor U14795 (N_14795,N_5118,N_6081);
xnor U14796 (N_14796,N_6696,N_9819);
or U14797 (N_14797,N_8869,N_8688);
xnor U14798 (N_14798,N_9300,N_7828);
nor U14799 (N_14799,N_9657,N_7013);
or U14800 (N_14800,N_6277,N_7687);
nor U14801 (N_14801,N_7395,N_5499);
nor U14802 (N_14802,N_5169,N_8149);
nand U14803 (N_14803,N_9590,N_6348);
and U14804 (N_14804,N_5033,N_5432);
nand U14805 (N_14805,N_7586,N_9639);
or U14806 (N_14806,N_5467,N_8400);
xor U14807 (N_14807,N_5083,N_7561);
nand U14808 (N_14808,N_8928,N_8908);
xnor U14809 (N_14809,N_5712,N_8558);
xor U14810 (N_14810,N_8693,N_5525);
xor U14811 (N_14811,N_6272,N_5208);
nand U14812 (N_14812,N_7351,N_7319);
xor U14813 (N_14813,N_5165,N_8449);
nand U14814 (N_14814,N_5561,N_8877);
nand U14815 (N_14815,N_5086,N_7363);
nand U14816 (N_14816,N_9191,N_8900);
nor U14817 (N_14817,N_8942,N_7357);
and U14818 (N_14818,N_7577,N_8304);
nand U14819 (N_14819,N_6226,N_7729);
nor U14820 (N_14820,N_7801,N_6572);
and U14821 (N_14821,N_7687,N_7293);
nand U14822 (N_14822,N_5236,N_9251);
nor U14823 (N_14823,N_7451,N_7993);
or U14824 (N_14824,N_7288,N_7348);
or U14825 (N_14825,N_7305,N_7773);
nand U14826 (N_14826,N_6051,N_7628);
nor U14827 (N_14827,N_6038,N_8639);
nand U14828 (N_14828,N_8143,N_6274);
nand U14829 (N_14829,N_9423,N_6335);
nor U14830 (N_14830,N_9672,N_7912);
and U14831 (N_14831,N_6304,N_9400);
xnor U14832 (N_14832,N_5168,N_9896);
and U14833 (N_14833,N_6102,N_5800);
xnor U14834 (N_14834,N_9366,N_8007);
or U14835 (N_14835,N_9121,N_8149);
and U14836 (N_14836,N_7071,N_5211);
nand U14837 (N_14837,N_7332,N_5308);
or U14838 (N_14838,N_7199,N_5734);
nand U14839 (N_14839,N_8497,N_7212);
or U14840 (N_14840,N_5114,N_9586);
and U14841 (N_14841,N_8348,N_7651);
nor U14842 (N_14842,N_8621,N_9065);
or U14843 (N_14843,N_8712,N_7969);
nand U14844 (N_14844,N_9160,N_5837);
or U14845 (N_14845,N_6512,N_5967);
and U14846 (N_14846,N_9469,N_5905);
xnor U14847 (N_14847,N_8289,N_5685);
nand U14848 (N_14848,N_5723,N_7729);
xor U14849 (N_14849,N_7973,N_5694);
xnor U14850 (N_14850,N_9448,N_7312);
or U14851 (N_14851,N_6565,N_9281);
nand U14852 (N_14852,N_8548,N_5429);
or U14853 (N_14853,N_6511,N_8268);
nand U14854 (N_14854,N_5636,N_7361);
or U14855 (N_14855,N_6449,N_6140);
xnor U14856 (N_14856,N_9467,N_9011);
xnor U14857 (N_14857,N_9294,N_8370);
xor U14858 (N_14858,N_9084,N_6508);
xnor U14859 (N_14859,N_6112,N_6389);
or U14860 (N_14860,N_6756,N_7114);
and U14861 (N_14861,N_9833,N_9319);
xor U14862 (N_14862,N_8410,N_8068);
xnor U14863 (N_14863,N_5361,N_7321);
xnor U14864 (N_14864,N_9620,N_5729);
or U14865 (N_14865,N_8878,N_8240);
and U14866 (N_14866,N_8662,N_9990);
or U14867 (N_14867,N_7099,N_6789);
nand U14868 (N_14868,N_8936,N_6618);
or U14869 (N_14869,N_6983,N_7181);
nor U14870 (N_14870,N_9530,N_9302);
nand U14871 (N_14871,N_7563,N_7909);
and U14872 (N_14872,N_9622,N_5644);
xnor U14873 (N_14873,N_7711,N_7123);
or U14874 (N_14874,N_7339,N_8844);
and U14875 (N_14875,N_7645,N_9915);
and U14876 (N_14876,N_6422,N_9138);
nand U14877 (N_14877,N_7901,N_5239);
xor U14878 (N_14878,N_7959,N_9773);
nand U14879 (N_14879,N_7309,N_8731);
or U14880 (N_14880,N_7345,N_9064);
xor U14881 (N_14881,N_7879,N_5449);
or U14882 (N_14882,N_9976,N_7097);
and U14883 (N_14883,N_9630,N_8118);
nor U14884 (N_14884,N_8765,N_7107);
or U14885 (N_14885,N_7282,N_5465);
nor U14886 (N_14886,N_7471,N_6977);
xor U14887 (N_14887,N_8621,N_7906);
or U14888 (N_14888,N_5602,N_9470);
nor U14889 (N_14889,N_9151,N_6079);
and U14890 (N_14890,N_6381,N_9239);
or U14891 (N_14891,N_6062,N_9591);
nand U14892 (N_14892,N_5962,N_9108);
and U14893 (N_14893,N_8145,N_7408);
xnor U14894 (N_14894,N_9753,N_7591);
nand U14895 (N_14895,N_5870,N_5800);
or U14896 (N_14896,N_9276,N_7539);
nor U14897 (N_14897,N_7648,N_6357);
nand U14898 (N_14898,N_5088,N_7548);
nor U14899 (N_14899,N_5197,N_5309);
xnor U14900 (N_14900,N_7066,N_6846);
nand U14901 (N_14901,N_8665,N_9067);
or U14902 (N_14902,N_9076,N_6775);
or U14903 (N_14903,N_8692,N_5962);
nand U14904 (N_14904,N_7786,N_5848);
nand U14905 (N_14905,N_8088,N_5392);
and U14906 (N_14906,N_6993,N_6704);
nand U14907 (N_14907,N_5310,N_6205);
nand U14908 (N_14908,N_5585,N_8659);
nor U14909 (N_14909,N_8247,N_6471);
and U14910 (N_14910,N_9287,N_5823);
or U14911 (N_14911,N_7513,N_5585);
and U14912 (N_14912,N_9851,N_9041);
and U14913 (N_14913,N_8886,N_5310);
and U14914 (N_14914,N_5131,N_6907);
xnor U14915 (N_14915,N_5425,N_5749);
or U14916 (N_14916,N_8758,N_7672);
and U14917 (N_14917,N_8163,N_5066);
xor U14918 (N_14918,N_9273,N_8816);
xnor U14919 (N_14919,N_6886,N_9041);
nor U14920 (N_14920,N_7560,N_9241);
and U14921 (N_14921,N_9156,N_6720);
or U14922 (N_14922,N_5942,N_9145);
xor U14923 (N_14923,N_7231,N_9896);
and U14924 (N_14924,N_5395,N_9304);
or U14925 (N_14925,N_6323,N_8311);
and U14926 (N_14926,N_5745,N_9899);
nand U14927 (N_14927,N_6418,N_9502);
nor U14928 (N_14928,N_7214,N_5077);
nor U14929 (N_14929,N_9037,N_5142);
nand U14930 (N_14930,N_6700,N_8648);
nand U14931 (N_14931,N_7657,N_5853);
or U14932 (N_14932,N_7678,N_9284);
xnor U14933 (N_14933,N_5785,N_9996);
nor U14934 (N_14934,N_7743,N_9677);
xor U14935 (N_14935,N_6466,N_9292);
and U14936 (N_14936,N_9561,N_7047);
xnor U14937 (N_14937,N_9827,N_9175);
and U14938 (N_14938,N_7847,N_5256);
or U14939 (N_14939,N_7677,N_6712);
nor U14940 (N_14940,N_9233,N_7971);
xnor U14941 (N_14941,N_7181,N_5317);
xor U14942 (N_14942,N_7572,N_9481);
nor U14943 (N_14943,N_6592,N_9646);
nor U14944 (N_14944,N_5145,N_9283);
nor U14945 (N_14945,N_9944,N_7365);
or U14946 (N_14946,N_9908,N_8508);
or U14947 (N_14947,N_6793,N_6681);
xnor U14948 (N_14948,N_9403,N_9048);
or U14949 (N_14949,N_7232,N_7705);
and U14950 (N_14950,N_8001,N_7061);
xor U14951 (N_14951,N_9543,N_6774);
and U14952 (N_14952,N_9590,N_6880);
nor U14953 (N_14953,N_8428,N_9989);
and U14954 (N_14954,N_8290,N_6751);
nand U14955 (N_14955,N_5415,N_5214);
nand U14956 (N_14956,N_7776,N_7458);
nor U14957 (N_14957,N_9066,N_6148);
nor U14958 (N_14958,N_5734,N_9667);
nor U14959 (N_14959,N_8130,N_5979);
and U14960 (N_14960,N_7956,N_5984);
or U14961 (N_14961,N_9122,N_6308);
and U14962 (N_14962,N_7413,N_5052);
xor U14963 (N_14963,N_9931,N_8981);
or U14964 (N_14964,N_6292,N_8784);
and U14965 (N_14965,N_7473,N_5696);
or U14966 (N_14966,N_9113,N_7465);
or U14967 (N_14967,N_5498,N_8898);
and U14968 (N_14968,N_5274,N_7556);
nand U14969 (N_14969,N_6970,N_9981);
nor U14970 (N_14970,N_5238,N_7925);
nor U14971 (N_14971,N_9504,N_5618);
nor U14972 (N_14972,N_7988,N_6339);
and U14973 (N_14973,N_5752,N_6653);
or U14974 (N_14974,N_6324,N_5484);
and U14975 (N_14975,N_8652,N_5545);
nand U14976 (N_14976,N_9163,N_5234);
xor U14977 (N_14977,N_7030,N_6370);
nand U14978 (N_14978,N_8272,N_7277);
and U14979 (N_14979,N_8382,N_6849);
and U14980 (N_14980,N_5993,N_9938);
and U14981 (N_14981,N_6988,N_8182);
nand U14982 (N_14982,N_5278,N_8105);
or U14983 (N_14983,N_8042,N_6411);
and U14984 (N_14984,N_9046,N_5729);
nand U14985 (N_14985,N_5294,N_6574);
nand U14986 (N_14986,N_7429,N_7116);
nor U14987 (N_14987,N_7318,N_6947);
xor U14988 (N_14988,N_5521,N_9226);
nand U14989 (N_14989,N_9063,N_5683);
nor U14990 (N_14990,N_8256,N_5543);
or U14991 (N_14991,N_6969,N_8205);
or U14992 (N_14992,N_9585,N_5034);
and U14993 (N_14993,N_8270,N_8550);
and U14994 (N_14994,N_6997,N_7243);
xnor U14995 (N_14995,N_8826,N_7945);
or U14996 (N_14996,N_8073,N_7170);
xnor U14997 (N_14997,N_9842,N_7354);
or U14998 (N_14998,N_5181,N_5138);
nand U14999 (N_14999,N_6971,N_5597);
nand U15000 (N_15000,N_13999,N_11398);
and U15001 (N_15001,N_13866,N_14409);
and U15002 (N_15002,N_12822,N_10376);
xnor U15003 (N_15003,N_12853,N_14463);
xnor U15004 (N_15004,N_13328,N_14018);
xnor U15005 (N_15005,N_13822,N_14001);
xor U15006 (N_15006,N_12071,N_11101);
or U15007 (N_15007,N_10388,N_14902);
nand U15008 (N_15008,N_12885,N_12030);
nor U15009 (N_15009,N_13269,N_10967);
nand U15010 (N_15010,N_14461,N_12864);
xnor U15011 (N_15011,N_10992,N_12743);
or U15012 (N_15012,N_11200,N_13386);
or U15013 (N_15013,N_14655,N_10979);
nand U15014 (N_15014,N_12462,N_11401);
nand U15015 (N_15015,N_14381,N_13112);
and U15016 (N_15016,N_13945,N_11237);
or U15017 (N_15017,N_12664,N_11329);
nand U15018 (N_15018,N_13399,N_13816);
xnor U15019 (N_15019,N_14485,N_11457);
and U15020 (N_15020,N_10447,N_10123);
nor U15021 (N_15021,N_10427,N_12389);
and U15022 (N_15022,N_14193,N_12940);
xor U15023 (N_15023,N_11198,N_13082);
xor U15024 (N_15024,N_13201,N_13874);
nand U15025 (N_15025,N_11183,N_10189);
or U15026 (N_15026,N_12975,N_14512);
and U15027 (N_15027,N_11671,N_10135);
and U15028 (N_15028,N_13780,N_10499);
or U15029 (N_15029,N_11925,N_12816);
and U15030 (N_15030,N_10477,N_12114);
or U15031 (N_15031,N_10625,N_13955);
and U15032 (N_15032,N_10698,N_11432);
xor U15033 (N_15033,N_10888,N_13211);
or U15034 (N_15034,N_14804,N_10849);
nor U15035 (N_15035,N_13752,N_10103);
nand U15036 (N_15036,N_13544,N_13693);
nor U15037 (N_15037,N_12970,N_14363);
and U15038 (N_15038,N_13690,N_14423);
nor U15039 (N_15039,N_13712,N_11632);
nor U15040 (N_15040,N_14360,N_13204);
nor U15041 (N_15041,N_14375,N_10090);
or U15042 (N_15042,N_10913,N_14402);
nor U15043 (N_15043,N_14337,N_14931);
nand U15044 (N_15044,N_13965,N_12798);
and U15045 (N_15045,N_11738,N_14755);
xnor U15046 (N_15046,N_12536,N_13247);
or U15047 (N_15047,N_13340,N_13276);
nand U15048 (N_15048,N_13393,N_12554);
and U15049 (N_15049,N_14087,N_10915);
and U15050 (N_15050,N_10786,N_11240);
nor U15051 (N_15051,N_13427,N_13251);
xnor U15052 (N_15052,N_11438,N_13238);
nand U15053 (N_15053,N_12806,N_10776);
or U15054 (N_15054,N_12006,N_12882);
or U15055 (N_15055,N_12989,N_11212);
and U15056 (N_15056,N_13703,N_10880);
xnor U15057 (N_15057,N_13107,N_12920);
nand U15058 (N_15058,N_13715,N_12364);
nand U15059 (N_15059,N_14333,N_10951);
and U15060 (N_15060,N_10164,N_10016);
xnor U15061 (N_15061,N_14564,N_13319);
or U15062 (N_15062,N_13080,N_14951);
and U15063 (N_15063,N_12715,N_13264);
and U15064 (N_15064,N_10702,N_13883);
nor U15065 (N_15065,N_12847,N_12767);
xnor U15066 (N_15066,N_13627,N_14208);
nor U15067 (N_15067,N_13597,N_14326);
nor U15068 (N_15068,N_10464,N_11260);
and U15069 (N_15069,N_11355,N_13587);
nand U15070 (N_15070,N_13392,N_10287);
nor U15071 (N_15071,N_11096,N_13293);
xnor U15072 (N_15072,N_11687,N_14594);
nor U15073 (N_15073,N_12826,N_11667);
or U15074 (N_15074,N_11711,N_14657);
nor U15075 (N_15075,N_12420,N_10645);
nor U15076 (N_15076,N_10817,N_13020);
nand U15077 (N_15077,N_14444,N_11822);
nor U15078 (N_15078,N_11487,N_12180);
nor U15079 (N_15079,N_13259,N_11326);
nand U15080 (N_15080,N_12145,N_12582);
nor U15081 (N_15081,N_11187,N_14611);
or U15082 (N_15082,N_11518,N_13330);
and U15083 (N_15083,N_11106,N_14926);
or U15084 (N_15084,N_12884,N_13362);
nand U15085 (N_15085,N_10032,N_11416);
and U15086 (N_15086,N_10610,N_13061);
and U15087 (N_15087,N_14453,N_12903);
nor U15088 (N_15088,N_13709,N_10219);
nand U15089 (N_15089,N_10833,N_14276);
nand U15090 (N_15090,N_11128,N_13058);
nor U15091 (N_15091,N_13434,N_10803);
nor U15092 (N_15092,N_12883,N_10401);
nor U15093 (N_15093,N_13696,N_10836);
nor U15094 (N_15094,N_14012,N_11344);
nand U15095 (N_15095,N_11454,N_12500);
or U15096 (N_15096,N_12445,N_11215);
xor U15097 (N_15097,N_14542,N_14278);
nand U15098 (N_15098,N_10601,N_12363);
xnor U15099 (N_15099,N_12993,N_10630);
or U15100 (N_15100,N_14458,N_14960);
nand U15101 (N_15101,N_12906,N_10246);
or U15102 (N_15102,N_11074,N_10166);
or U15103 (N_15103,N_13173,N_10064);
nor U15104 (N_15104,N_13086,N_13667);
nand U15105 (N_15105,N_12540,N_11390);
or U15106 (N_15106,N_11273,N_10999);
or U15107 (N_15107,N_14364,N_14996);
nor U15108 (N_15108,N_14867,N_10357);
nand U15109 (N_15109,N_10983,N_11455);
and U15110 (N_15110,N_14451,N_13441);
nand U15111 (N_15111,N_11626,N_14273);
nand U15112 (N_15112,N_11916,N_11895);
xnor U15113 (N_15113,N_10087,N_11970);
and U15114 (N_15114,N_14620,N_14894);
and U15115 (N_15115,N_13047,N_10536);
nor U15116 (N_15116,N_13761,N_12466);
and U15117 (N_15117,N_10538,N_11782);
nor U15118 (N_15118,N_14380,N_14006);
or U15119 (N_15119,N_10091,N_11542);
and U15120 (N_15120,N_14190,N_14993);
or U15121 (N_15121,N_12168,N_12497);
nor U15122 (N_15122,N_11206,N_12605);
nor U15123 (N_15123,N_13605,N_10043);
xor U15124 (N_15124,N_13215,N_11075);
nand U15125 (N_15125,N_10775,N_14302);
nand U15126 (N_15126,N_14492,N_11793);
or U15127 (N_15127,N_12014,N_14039);
and U15128 (N_15128,N_14147,N_10758);
or U15129 (N_15129,N_10738,N_11290);
or U15130 (N_15130,N_12714,N_10877);
or U15131 (N_15131,N_13950,N_10522);
and U15132 (N_15132,N_14370,N_10764);
xor U15133 (N_15133,N_11189,N_11691);
or U15134 (N_15134,N_11866,N_11930);
and U15135 (N_15135,N_14650,N_12679);
and U15136 (N_15136,N_14315,N_10067);
and U15137 (N_15137,N_10424,N_14917);
and U15138 (N_15138,N_12656,N_10885);
nand U15139 (N_15139,N_10117,N_14102);
or U15140 (N_15140,N_12710,N_14774);
nor U15141 (N_15141,N_12307,N_10021);
or U15142 (N_15142,N_14879,N_11689);
and U15143 (N_15143,N_13856,N_10220);
nand U15144 (N_15144,N_13042,N_14435);
nor U15145 (N_15145,N_14590,N_14271);
nand U15146 (N_15146,N_12593,N_14311);
nand U15147 (N_15147,N_11571,N_14119);
or U15148 (N_15148,N_10856,N_13579);
nor U15149 (N_15149,N_11351,N_12378);
nor U15150 (N_15150,N_13472,N_10864);
xnor U15151 (N_15151,N_14694,N_11717);
xnor U15152 (N_15152,N_11127,N_10286);
nor U15153 (N_15153,N_10453,N_11041);
nor U15154 (N_15154,N_14167,N_14881);
nand U15155 (N_15155,N_13758,N_13754);
xnor U15156 (N_15156,N_10070,N_14297);
xor U15157 (N_15157,N_14216,N_13174);
xnor U15158 (N_15158,N_10523,N_12692);
nand U15159 (N_15159,N_11712,N_11214);
nand U15160 (N_15160,N_13474,N_11250);
nand U15161 (N_15161,N_11978,N_10819);
and U15162 (N_15162,N_12653,N_12726);
xnor U15163 (N_15163,N_11479,N_13638);
nand U15164 (N_15164,N_11406,N_10598);
nand U15165 (N_15165,N_13523,N_13998);
and U15166 (N_15166,N_14214,N_10696);
nor U15167 (N_15167,N_13845,N_13734);
or U15168 (N_15168,N_10027,N_11044);
xnor U15169 (N_15169,N_14464,N_10188);
nand U15170 (N_15170,N_13982,N_14303);
or U15171 (N_15171,N_14267,N_14390);
and U15172 (N_15172,N_13223,N_12665);
or U15173 (N_15173,N_12248,N_12918);
or U15174 (N_15174,N_12097,N_10129);
xor U15175 (N_15175,N_14796,N_11072);
xnor U15176 (N_15176,N_11262,N_14396);
and U15177 (N_15177,N_14225,N_11057);
or U15178 (N_15178,N_12400,N_11425);
nand U15179 (N_15179,N_12428,N_10485);
nor U15180 (N_15180,N_13286,N_13622);
and U15181 (N_15181,N_12407,N_12240);
or U15182 (N_15182,N_12325,N_14729);
nand U15183 (N_15183,N_12844,N_10660);
and U15184 (N_15184,N_10642,N_13275);
nor U15185 (N_15185,N_12241,N_13806);
or U15186 (N_15186,N_12104,N_10431);
xor U15187 (N_15187,N_12217,N_11734);
or U15188 (N_15188,N_12251,N_11790);
or U15189 (N_15189,N_14395,N_10059);
xor U15190 (N_15190,N_12837,N_11472);
or U15191 (N_15191,N_10311,N_13193);
or U15192 (N_15192,N_13954,N_10600);
xnor U15193 (N_15193,N_14983,N_13561);
nand U15194 (N_15194,N_12132,N_11062);
xor U15195 (N_15195,N_10560,N_11405);
nor U15196 (N_15196,N_11115,N_13594);
xor U15197 (N_15197,N_12062,N_11634);
xor U15198 (N_15198,N_11028,N_14771);
xor U15199 (N_15199,N_14721,N_14106);
nor U15200 (N_15200,N_14747,N_13175);
and U15201 (N_15201,N_14582,N_13202);
xor U15202 (N_15202,N_13987,N_11500);
or U15203 (N_15203,N_12629,N_13565);
xnor U15204 (N_15204,N_13819,N_11474);
xor U15205 (N_15205,N_14070,N_14124);
xnor U15206 (N_15206,N_10524,N_13531);
nand U15207 (N_15207,N_10667,N_14838);
nand U15208 (N_15208,N_14571,N_13847);
nand U15209 (N_15209,N_11141,N_11340);
nand U15210 (N_15210,N_10230,N_10476);
nor U15211 (N_15211,N_10301,N_12173);
or U15212 (N_15212,N_11478,N_11102);
or U15213 (N_15213,N_14263,N_14616);
and U15214 (N_15214,N_11919,N_11533);
nor U15215 (N_15215,N_12449,N_13048);
or U15216 (N_15216,N_13871,N_13070);
xnor U15217 (N_15217,N_13469,N_13731);
or U15218 (N_15218,N_11315,N_14946);
nor U15219 (N_15219,N_10735,N_13583);
or U15220 (N_15220,N_13801,N_10386);
or U15221 (N_15221,N_10868,N_12453);
xnor U15222 (N_15222,N_10903,N_10873);
and U15223 (N_15223,N_12245,N_13180);
nand U15224 (N_15224,N_13763,N_11413);
xor U15225 (N_15225,N_14189,N_12136);
nand U15226 (N_15226,N_12327,N_11373);
or U15227 (N_15227,N_10841,N_10394);
nor U15228 (N_15228,N_13039,N_10143);
and U15229 (N_15229,N_12817,N_14172);
or U15230 (N_15230,N_10916,N_14743);
nand U15231 (N_15231,N_13558,N_14356);
xor U15232 (N_15232,N_10297,N_11664);
or U15233 (N_15233,N_13069,N_10118);
xnor U15234 (N_15234,N_13268,N_13348);
xor U15235 (N_15235,N_10369,N_11251);
or U15236 (N_15236,N_12133,N_10520);
xnor U15237 (N_15237,N_14568,N_12519);
nor U15238 (N_15238,N_11374,N_10508);
or U15239 (N_15239,N_10761,N_13835);
xnor U15240 (N_15240,N_10403,N_13050);
nand U15241 (N_15241,N_12463,N_14839);
or U15242 (N_15242,N_12652,N_12698);
nor U15243 (N_15243,N_12057,N_10283);
nand U15244 (N_15244,N_13864,N_14929);
nor U15245 (N_15245,N_12976,N_14678);
nor U15246 (N_15246,N_10549,N_11180);
and U15247 (N_15247,N_14666,N_13971);
nand U15248 (N_15248,N_14196,N_11951);
xnor U15249 (N_15249,N_14258,N_10025);
or U15250 (N_15250,N_11610,N_14572);
and U15251 (N_15251,N_14977,N_13098);
nor U15252 (N_15252,N_11991,N_11055);
and U15253 (N_15253,N_10878,N_12399);
nand U15254 (N_15254,N_13718,N_14352);
or U15255 (N_15255,N_14502,N_13074);
xor U15256 (N_15256,N_14751,N_12394);
or U15257 (N_15257,N_12712,N_10104);
or U15258 (N_15258,N_12748,N_10715);
or U15259 (N_15259,N_13220,N_13036);
xnor U15260 (N_15260,N_14872,N_12915);
or U15261 (N_15261,N_14766,N_11625);
nor U15262 (N_15262,N_14093,N_14832);
xnor U15263 (N_15263,N_11331,N_12103);
or U15264 (N_15264,N_11674,N_11155);
xor U15265 (N_15265,N_14702,N_14534);
nand U15266 (N_15266,N_14324,N_10593);
or U15267 (N_15267,N_10334,N_11651);
and U15268 (N_15268,N_11143,N_13697);
nand U15269 (N_15269,N_10838,N_14135);
and U15270 (N_15270,N_14210,N_14596);
nor U15271 (N_15271,N_11371,N_12728);
nand U15272 (N_15272,N_14159,N_13993);
or U15273 (N_15273,N_12659,N_10919);
nor U15274 (N_15274,N_14095,N_11134);
nor U15275 (N_15275,N_13942,N_12213);
xor U15276 (N_15276,N_10402,N_13366);
and U15277 (N_15277,N_13191,N_13342);
or U15278 (N_15278,N_11224,N_11567);
nor U15279 (N_15279,N_13480,N_11439);
nor U15280 (N_15280,N_11507,N_13899);
nor U15281 (N_15281,N_12082,N_13821);
and U15282 (N_15282,N_13009,N_11252);
xor U15283 (N_15283,N_11071,N_10602);
nor U15284 (N_15284,N_10443,N_12904);
xor U15285 (N_15285,N_12015,N_12231);
xnor U15286 (N_15286,N_11482,N_14111);
and U15287 (N_15287,N_14520,N_10668);
and U15288 (N_15288,N_10678,N_10718);
xnor U15289 (N_15289,N_14178,N_11116);
nand U15290 (N_15290,N_11085,N_11993);
xnor U15291 (N_15291,N_13290,N_12452);
and U15292 (N_15292,N_13903,N_11157);
xor U15293 (N_15293,N_12633,N_13357);
nor U15294 (N_15294,N_10559,N_11268);
or U15295 (N_15295,N_11238,N_14280);
nand U15296 (N_15296,N_12049,N_12539);
nand U15297 (N_15297,N_12160,N_11733);
nand U15298 (N_15298,N_14430,N_10177);
or U15299 (N_15299,N_12396,N_13504);
or U15300 (N_15300,N_12064,N_14875);
xor U15301 (N_15301,N_12668,N_14962);
or U15302 (N_15302,N_11806,N_13165);
and U15303 (N_15303,N_14217,N_11977);
xor U15304 (N_15304,N_12306,N_13094);
xor U15305 (N_15305,N_10886,N_10943);
and U15306 (N_15306,N_12894,N_11988);
xor U15307 (N_15307,N_14516,N_14933);
or U15308 (N_15308,N_11126,N_14448);
xnor U15309 (N_15309,N_14897,N_11575);
nor U15310 (N_15310,N_14126,N_10440);
and U15311 (N_15311,N_13485,N_14110);
and U15312 (N_15312,N_13155,N_12723);
nand U15313 (N_15313,N_10907,N_11657);
xor U15314 (N_15314,N_14412,N_12654);
nand U15315 (N_15315,N_12948,N_10362);
or U15316 (N_15316,N_10451,N_13507);
and U15317 (N_15317,N_14914,N_14293);
and U15318 (N_15318,N_14882,N_13887);
xor U15319 (N_15319,N_13875,N_13656);
nor U15320 (N_15320,N_10210,N_11468);
nand U15321 (N_15321,N_14846,N_14699);
nor U15322 (N_15322,N_10596,N_14811);
or U15323 (N_15323,N_11595,N_12171);
nor U15324 (N_15324,N_10428,N_11515);
nand U15325 (N_15325,N_12867,N_11872);
nor U15326 (N_15326,N_14792,N_14338);
or U15327 (N_15327,N_11746,N_12812);
or U15328 (N_15328,N_12274,N_12427);
and U15329 (N_15329,N_10018,N_14248);
nand U15330 (N_15330,N_10013,N_12148);
and U15331 (N_15331,N_14849,N_12107);
nand U15332 (N_15332,N_13836,N_14294);
nand U15333 (N_15333,N_12571,N_10222);
and U15334 (N_15334,N_11152,N_11483);
xnor U15335 (N_15335,N_11807,N_12416);
and U15336 (N_15336,N_13534,N_10304);
and U15337 (N_15337,N_12998,N_12968);
nand U15338 (N_15338,N_12780,N_12919);
xor U15339 (N_15339,N_10808,N_12786);
xnor U15340 (N_15340,N_11636,N_11713);
xor U15341 (N_15341,N_14062,N_10434);
and U15342 (N_15342,N_12525,N_14022);
or U15343 (N_15343,N_11714,N_13486);
nor U15344 (N_15344,N_11752,N_13858);
nor U15345 (N_15345,N_14861,N_11678);
nor U15346 (N_15346,N_10727,N_13820);
or U15347 (N_15347,N_13225,N_11559);
or U15348 (N_15348,N_14250,N_14096);
nor U15349 (N_15349,N_10194,N_13440);
and U15350 (N_15350,N_12163,N_10924);
and U15351 (N_15351,N_10521,N_12549);
nor U15352 (N_15352,N_14470,N_10557);
nand U15353 (N_15353,N_10482,N_13040);
or U15354 (N_15354,N_10479,N_10934);
or U15355 (N_15355,N_13444,N_14007);
nand U15356 (N_15356,N_11317,N_11555);
nand U15357 (N_15357,N_14975,N_13332);
xor U15358 (N_15358,N_11441,N_13519);
and U15359 (N_15359,N_14915,N_13272);
nand U15360 (N_15360,N_12166,N_14529);
nand U15361 (N_15361,N_14685,N_12944);
nor U15362 (N_15362,N_11799,N_10211);
xor U15363 (N_15363,N_14887,N_13224);
nor U15364 (N_15364,N_12016,N_11794);
or U15365 (N_15365,N_10842,N_14223);
and U15366 (N_15366,N_10797,N_11148);
xor U15367 (N_15367,N_14094,N_11700);
and U15368 (N_15368,N_14489,N_14599);
nand U15369 (N_15369,N_14369,N_14733);
nand U15370 (N_15370,N_10707,N_11572);
nor U15371 (N_15371,N_11829,N_10708);
and U15372 (N_15372,N_10778,N_11066);
or U15373 (N_15373,N_10689,N_14296);
xnor U15374 (N_15374,N_14232,N_11186);
xnor U15375 (N_15375,N_12598,N_13126);
or U15376 (N_15376,N_14530,N_10539);
or U15377 (N_15377,N_11810,N_12156);
nor U15378 (N_15378,N_13008,N_13572);
nor U15379 (N_15379,N_12935,N_10850);
nor U15380 (N_15380,N_13234,N_14506);
and U15381 (N_15381,N_13068,N_10266);
xor U15382 (N_15382,N_13571,N_10497);
and U15383 (N_15383,N_10950,N_10504);
nand U15384 (N_15384,N_10406,N_12913);
nand U15385 (N_15385,N_12486,N_14635);
and U15386 (N_15386,N_12784,N_10973);
or U15387 (N_15387,N_13203,N_10316);
or U15388 (N_15388,N_13028,N_10320);
nand U15389 (N_15389,N_13218,N_10081);
or U15390 (N_15390,N_13621,N_12290);
xnor U15391 (N_15391,N_13928,N_11628);
nor U15392 (N_15392,N_12476,N_11918);
and U15393 (N_15393,N_12567,N_10370);
xor U15394 (N_15394,N_13729,N_14531);
and U15395 (N_15395,N_12475,N_13181);
or U15396 (N_15396,N_13510,N_14361);
xor U15397 (N_15397,N_11909,N_11048);
nand U15398 (N_15398,N_14675,N_10325);
or U15399 (N_15399,N_12969,N_11497);
nor U15400 (N_15400,N_14127,N_14254);
or U15401 (N_15401,N_13650,N_13166);
or U15402 (N_15402,N_10429,N_11934);
or U15403 (N_15403,N_14667,N_10410);
and U15404 (N_15404,N_10754,N_13460);
xnor U15405 (N_15405,N_14078,N_12119);
or U15406 (N_15406,N_11360,N_14921);
and U15407 (N_15407,N_13862,N_13018);
xnor U15408 (N_15408,N_12761,N_13807);
nand U15409 (N_15409,N_11284,N_13598);
or U15410 (N_15410,N_10237,N_11861);
nand U15411 (N_15411,N_12293,N_12966);
and U15412 (N_15412,N_12996,N_12927);
xor U15413 (N_15413,N_11650,N_11121);
and U15414 (N_15414,N_14477,N_13412);
nor U15415 (N_15415,N_13445,N_14040);
nor U15416 (N_15416,N_12259,N_13209);
or U15417 (N_15417,N_10692,N_14578);
xnor U15418 (N_15418,N_12724,N_12950);
and U15419 (N_15419,N_11655,N_12058);
xnor U15420 (N_15420,N_11865,N_10659);
nor U15421 (N_15421,N_13250,N_14060);
and U15422 (N_15422,N_11429,N_14362);
and U15423 (N_15423,N_11837,N_10638);
or U15424 (N_15424,N_12887,N_13576);
xor U15425 (N_15425,N_14756,N_10231);
or U15426 (N_15426,N_13610,N_14630);
xor U15427 (N_15427,N_10132,N_11588);
and U15428 (N_15428,N_10806,N_12455);
or U15429 (N_15429,N_10444,N_12342);
or U15430 (N_15430,N_13795,N_11675);
xnor U15431 (N_15431,N_12308,N_10567);
or U15432 (N_15432,N_11409,N_13505);
nand U15433 (N_15433,N_11508,N_12794);
nand U15434 (N_15434,N_13137,N_14490);
or U15435 (N_15435,N_14515,N_14026);
nor U15436 (N_15436,N_11471,N_13450);
or U15437 (N_15437,N_11410,N_13185);
nor U15438 (N_15438,N_13035,N_11614);
and U15439 (N_15439,N_14035,N_13302);
nor U15440 (N_15440,N_13162,N_10858);
xnor U15441 (N_15441,N_12003,N_13213);
and U15442 (N_15442,N_14622,N_13732);
xor U15443 (N_15443,N_13979,N_13741);
and U15444 (N_15444,N_10425,N_13897);
nor U15445 (N_15445,N_14943,N_12023);
nand U15446 (N_15446,N_12279,N_14129);
nand U15447 (N_15447,N_14950,N_13421);
nor U15448 (N_15448,N_13377,N_10382);
nor U15449 (N_15449,N_14858,N_13593);
nor U15450 (N_15450,N_14257,N_11910);
or U15451 (N_15451,N_10512,N_10739);
xor U15452 (N_15452,N_14964,N_12199);
xnor U15453 (N_15453,N_14603,N_10187);
nor U15454 (N_15454,N_13685,N_13194);
nor U15455 (N_15455,N_14373,N_12541);
and U15456 (N_15456,N_11905,N_13435);
nor U15457 (N_15457,N_11608,N_14998);
or U15458 (N_15458,N_12220,N_12219);
nor U15459 (N_15459,N_12155,N_12451);
nand U15460 (N_15460,N_11192,N_10768);
nor U15461 (N_15461,N_14191,N_13532);
and U15462 (N_15462,N_12291,N_12739);
and U15463 (N_15463,N_12305,N_10161);
xnor U15464 (N_15464,N_11368,N_13674);
xnor U15465 (N_15465,N_10458,N_10473);
nand U15466 (N_15466,N_10221,N_10605);
xor U15467 (N_15467,N_11505,N_10996);
or U15468 (N_15468,N_14549,N_13829);
xor U15469 (N_15469,N_14313,N_12182);
nor U15470 (N_15470,N_11286,N_11556);
and U15471 (N_15471,N_12526,N_11431);
nand U15472 (N_15472,N_11694,N_12843);
and U15473 (N_15473,N_13492,N_10650);
and U15474 (N_15474,N_10564,N_10652);
xnor U15475 (N_15475,N_13724,N_12807);
nor U15476 (N_15476,N_12146,N_12411);
or U15477 (N_15477,N_14118,N_12147);
nand U15478 (N_15478,N_13996,N_12845);
xnor U15479 (N_15479,N_13298,N_12052);
nor U15480 (N_15480,N_11249,N_10899);
xor U15481 (N_15481,N_12223,N_11639);
xor U15482 (N_15482,N_12878,N_14883);
and U15483 (N_15483,N_10454,N_11568);
and U15484 (N_15484,N_10599,N_10395);
nor U15485 (N_15485,N_12460,N_14160);
and U15486 (N_15486,N_10379,N_12441);
and U15487 (N_15487,N_11851,N_10953);
nor U15488 (N_15488,N_12745,N_12765);
nand U15489 (N_15489,N_12754,N_14857);
nor U15490 (N_15490,N_12628,N_13292);
nand U15491 (N_15491,N_14826,N_11226);
or U15492 (N_15492,N_10383,N_13818);
nor U15493 (N_15493,N_10204,N_13358);
and U15494 (N_15494,N_11956,N_11773);
nand U15495 (N_15495,N_11422,N_10818);
xnor U15496 (N_15496,N_10576,N_12939);
nand U15497 (N_15497,N_13465,N_10227);
and U15498 (N_15498,N_12932,N_14498);
nor U15499 (N_15499,N_12189,N_11528);
or U15500 (N_15500,N_10271,N_12135);
xnor U15501 (N_15501,N_13351,N_12749);
or U15502 (N_15502,N_10619,N_14670);
xor U15503 (N_15503,N_10044,N_10178);
nor U15504 (N_15504,N_14000,N_13721);
nor U15505 (N_15505,N_10314,N_13071);
xor U15506 (N_15506,N_13848,N_12564);
nor U15507 (N_15507,N_10156,N_13477);
and U15508 (N_15508,N_10683,N_12208);
and U15509 (N_15509,N_12090,N_13163);
nand U15510 (N_15510,N_14610,N_14871);
nand U15511 (N_15511,N_14357,N_14455);
and U15512 (N_15512,N_11976,N_13533);
nand U15513 (N_15513,N_14074,N_12169);
nor U15514 (N_15514,N_13285,N_11530);
nor U15515 (N_15515,N_10618,N_14563);
or U15516 (N_15516,N_11424,N_10085);
nand U15517 (N_15517,N_12489,N_14884);
nor U15518 (N_15518,N_11514,N_13432);
nor U15519 (N_15519,N_13426,N_13616);
or U15520 (N_15520,N_10065,N_10985);
nor U15521 (N_15521,N_10046,N_10348);
nor U15522 (N_15522,N_14949,N_14801);
nor U15523 (N_15523,N_10871,N_13810);
xnor U15524 (N_15524,N_12320,N_11301);
or U15525 (N_15525,N_10197,N_14561);
nand U15526 (N_15526,N_10912,N_14619);
or U15527 (N_15527,N_14770,N_12127);
nand U15528 (N_15528,N_10920,N_11613);
nand U15529 (N_15529,N_10274,N_10009);
xor U15530 (N_15530,N_11463,N_12143);
and U15531 (N_15531,N_12448,N_10948);
nand U15532 (N_15532,N_13514,N_11370);
xnor U15533 (N_15533,N_11011,N_14776);
xor U15534 (N_15534,N_14965,N_14999);
or U15535 (N_15535,N_12684,N_14179);
and U15536 (N_15536,N_14525,N_14144);
xor U15537 (N_15537,N_11881,N_14696);
and U15538 (N_15538,N_13057,N_10131);
nand U15539 (N_15539,N_11236,N_10062);
and U15540 (N_15540,N_12093,N_12404);
and U15541 (N_15541,N_13384,N_14404);
nor U15542 (N_15542,N_10782,N_11949);
and U15543 (N_15543,N_12644,N_12863);
xnor U15544 (N_15544,N_13737,N_13869);
or U15545 (N_15545,N_13096,N_14305);
xnor U15546 (N_15546,N_10795,N_11112);
nand U15547 (N_15547,N_10097,N_13684);
nand U15548 (N_15548,N_12693,N_10991);
or U15549 (N_15549,N_10285,N_14708);
or U15550 (N_15550,N_11117,N_11384);
and U15551 (N_15551,N_14501,N_11965);
xnor U15552 (N_15552,N_12008,N_14320);
nand U15553 (N_15553,N_11648,N_12557);
xnor U15554 (N_15554,N_12938,N_10927);
or U15555 (N_15555,N_10976,N_12849);
nor U15556 (N_15556,N_13545,N_14941);
or U15557 (N_15557,N_14973,N_11216);
nand U15558 (N_15558,N_10055,N_13488);
nand U15559 (N_15559,N_11338,N_13401);
and U15560 (N_15560,N_14579,N_11059);
xnor U15561 (N_15561,N_14346,N_10686);
and U15562 (N_15562,N_12717,N_11231);
and U15563 (N_15563,N_11120,N_10573);
xor U15564 (N_15564,N_11885,N_13755);
nand U15565 (N_15565,N_14222,N_10998);
nor U15566 (N_15566,N_14438,N_10284);
xor U15567 (N_15567,N_11942,N_12979);
xnor U15568 (N_15568,N_14301,N_14827);
nor U15569 (N_15569,N_11926,N_13267);
or U15570 (N_15570,N_11311,N_12188);
xor U15571 (N_15571,N_13361,N_10665);
and U15572 (N_15572,N_10162,N_14986);
and U15573 (N_15573,N_12271,N_12286);
xor U15574 (N_15574,N_12861,N_10695);
and U15575 (N_15575,N_12854,N_10248);
and U15576 (N_15576,N_12756,N_13817);
nand U15577 (N_15577,N_11645,N_12496);
nand U15578 (N_15578,N_11103,N_11523);
xnor U15579 (N_15579,N_11423,N_12253);
xnor U15580 (N_15580,N_10407,N_11707);
nand U15581 (N_15581,N_12128,N_14137);
and U15582 (N_15582,N_10039,N_12035);
nand U15583 (N_15583,N_11476,N_13063);
nor U15584 (N_15584,N_12908,N_14809);
and U15585 (N_15585,N_11907,N_11299);
xnor U15586 (N_15586,N_14633,N_13778);
nand U15587 (N_15587,N_12921,N_13760);
xor U15588 (N_15588,N_10298,N_12473);
xor U15589 (N_15589,N_14231,N_11270);
nand U15590 (N_15590,N_14428,N_13024);
and U15591 (N_15591,N_13145,N_12434);
xor U15592 (N_15592,N_12575,N_11688);
nor U15593 (N_15593,N_10080,N_10603);
xnor U15594 (N_15594,N_14281,N_14574);
nor U15595 (N_15595,N_13857,N_11743);
and U15596 (N_15596,N_13805,N_10422);
nand U15597 (N_15597,N_14669,N_12838);
xnor U15598 (N_15598,N_12116,N_13479);
or U15599 (N_15599,N_12360,N_13462);
xor U15600 (N_15600,N_11092,N_11972);
nor U15601 (N_15601,N_11723,N_14880);
or U15602 (N_15602,N_14605,N_13612);
xor U15603 (N_15603,N_13840,N_14930);
or U15604 (N_15604,N_13639,N_14647);
xor U15605 (N_15605,N_12905,N_14471);
xnor U15606 (N_15606,N_11933,N_13258);
xnor U15607 (N_15607,N_11652,N_12926);
and U15608 (N_15608,N_12298,N_10397);
xor U15609 (N_15609,N_10957,N_14156);
nor U15610 (N_15610,N_13146,N_11780);
nand U15611 (N_15611,N_10537,N_12524);
or U15612 (N_15612,N_13844,N_12314);
or U15613 (N_15613,N_12690,N_14976);
nor U15614 (N_15614,N_12689,N_10050);
xnor U15615 (N_15615,N_12955,N_10988);
nor U15616 (N_15616,N_13908,N_11825);
and U15617 (N_15617,N_10942,N_10180);
nor U15618 (N_15618,N_12392,N_14814);
or U15619 (N_15619,N_13615,N_12187);
and U15620 (N_15620,N_12572,N_10014);
nor U15621 (N_15621,N_13345,N_11981);
xnor U15622 (N_15622,N_13849,N_11167);
xor U15623 (N_15623,N_13517,N_12545);
xor U15624 (N_15624,N_11715,N_13284);
nand U15625 (N_15625,N_11010,N_10970);
nor U15626 (N_15626,N_14090,N_10848);
nor U15627 (N_15627,N_14194,N_11114);
xor U15628 (N_15628,N_12587,N_10543);
and U15629 (N_15629,N_12439,N_11159);
xor U15630 (N_15630,N_14152,N_14325);
nand U15631 (N_15631,N_10812,N_12183);
or U15632 (N_15632,N_14744,N_10932);
nand U15633 (N_15633,N_13962,N_10396);
nand U15634 (N_15634,N_12161,N_12467);
nand U15635 (N_15635,N_10518,N_11144);
nor U15636 (N_15636,N_14886,N_10720);
or U15637 (N_15637,N_10887,N_14913);
xor U15638 (N_15638,N_14658,N_14604);
nor U15639 (N_15639,N_14785,N_12468);
nand U15640 (N_15640,N_10460,N_11932);
and U15641 (N_15641,N_13296,N_10632);
and U15642 (N_15642,N_12782,N_10811);
nand U15643 (N_15643,N_14259,N_10896);
or U15644 (N_15644,N_10218,N_10098);
nor U15645 (N_15645,N_12408,N_14953);
xnor U15646 (N_15646,N_13349,N_14030);
xor U15647 (N_15647,N_13045,N_13881);
xor U15648 (N_15648,N_12914,N_10083);
and U15649 (N_15649,N_12393,N_10313);
nor U15650 (N_15650,N_10214,N_10420);
nand U15651 (N_15651,N_12098,N_14252);
xnor U15652 (N_15652,N_11466,N_11615);
nand U15653 (N_15653,N_10317,N_11150);
nand U15654 (N_15654,N_10206,N_14546);
nor U15655 (N_15655,N_13105,N_10580);
nor U15656 (N_15656,N_11963,N_11435);
and U15657 (N_15657,N_12680,N_10209);
nand U15658 (N_15658,N_11903,N_12424);
or U15659 (N_15659,N_10302,N_14805);
xor U15660 (N_15660,N_10371,N_12112);
or U15661 (N_15661,N_13511,N_13952);
or U15662 (N_15662,N_13280,N_11809);
xor U15663 (N_15663,N_14992,N_12129);
or U15664 (N_15664,N_13481,N_13915);
nand U15665 (N_15665,N_13313,N_11193);
and U15666 (N_15666,N_12310,N_10267);
or U15667 (N_15667,N_14845,N_13265);
xnor U15668 (N_15668,N_13750,N_14940);
nor U15669 (N_15669,N_11884,N_13242);
nor U15670 (N_15670,N_11465,N_14283);
and U15671 (N_15671,N_13689,N_12421);
and U15672 (N_15672,N_13464,N_11870);
or U15673 (N_15673,N_13992,N_14469);
xnor U15674 (N_15674,N_10611,N_12075);
nand U15675 (N_15675,N_13859,N_10446);
or U15676 (N_15676,N_14056,N_10481);
and U15677 (N_15677,N_10861,N_14077);
and U15678 (N_15678,N_11285,N_13744);
and U15679 (N_15679,N_11283,N_12125);
nor U15680 (N_15680,N_11975,N_13052);
nor U15681 (N_15681,N_14932,N_14387);
xor U15682 (N_15682,N_13007,N_14608);
and U15683 (N_15683,N_13437,N_12872);
xnor U15684 (N_15684,N_13350,N_10509);
and U15685 (N_15685,N_12909,N_10989);
nor U15686 (N_15686,N_10006,N_10426);
or U15687 (N_15687,N_10011,N_14677);
or U15688 (N_15688,N_12624,N_10022);
or U15689 (N_15689,N_11166,N_10941);
and U15690 (N_15690,N_10163,N_10116);
nand U15691 (N_15691,N_10929,N_11722);
and U15692 (N_15692,N_13431,N_11164);
nor U15693 (N_15693,N_11365,N_14407);
or U15694 (N_15694,N_12830,N_12270);
and U15695 (N_15695,N_14705,N_10828);
and U15696 (N_15696,N_10914,N_12102);
or U15697 (N_15697,N_14995,N_14331);
xnor U15698 (N_15698,N_14038,N_12985);
nand U15699 (N_15699,N_10949,N_12170);
nand U15700 (N_15700,N_13665,N_11452);
nor U15701 (N_15701,N_11201,N_11397);
nand U15702 (N_15702,N_13704,N_11637);
and U15703 (N_15703,N_14730,N_12612);
or U15704 (N_15704,N_14474,N_14922);
and U15705 (N_15705,N_13994,N_14233);
and U15706 (N_15706,N_14537,N_12356);
xor U15707 (N_15707,N_12821,N_13785);
nand U15708 (N_15708,N_12077,N_11584);
and U15709 (N_15709,N_13217,N_14649);
xnor U15710 (N_15710,N_10042,N_12622);
nor U15711 (N_15711,N_13159,N_13143);
or U15712 (N_15712,N_10663,N_11381);
or U15713 (N_15713,N_14982,N_14173);
and U15714 (N_15714,N_10898,N_12391);
nor U15715 (N_15715,N_14199,N_14779);
or U15716 (N_15716,N_14437,N_13506);
and U15717 (N_15717,N_11022,N_11443);
nor U15718 (N_15718,N_13365,N_10829);
nand U15719 (N_15719,N_10608,N_12300);
xnor U15720 (N_15720,N_14146,N_12774);
or U15721 (N_15721,N_13937,N_13974);
and U15722 (N_15722,N_14299,N_13283);
and U15723 (N_15723,N_13680,N_12447);
nor U15724 (N_15724,N_10724,N_13198);
or U15725 (N_15725,N_13214,N_10077);
or U15726 (N_15726,N_12716,N_11816);
nor U15727 (N_15727,N_11546,N_10069);
nand U15728 (N_15728,N_13662,N_11047);
nand U15729 (N_15729,N_12444,N_11122);
nand U15730 (N_15730,N_13046,N_12063);
nand U15731 (N_15731,N_11385,N_14764);
and U15732 (N_15732,N_11305,N_13929);
nor U15733 (N_15733,N_11860,N_12937);
and U15734 (N_15734,N_12362,N_10489);
nand U15735 (N_15735,N_10449,N_13387);
xnor U15736 (N_15736,N_10472,N_12172);
xor U15737 (N_15737,N_12422,N_10507);
or U15738 (N_15738,N_13228,N_10264);
and U15739 (N_15739,N_13617,N_12042);
nor U15740 (N_15740,N_10900,N_11579);
nor U15741 (N_15741,N_10514,N_11132);
and U15742 (N_15742,N_14336,N_13142);
nor U15743 (N_15743,N_11481,N_10251);
nand U15744 (N_15744,N_10581,N_14803);
and U15745 (N_15745,N_10793,N_12076);
and U15746 (N_15746,N_11369,N_12144);
or U15747 (N_15747,N_11361,N_13783);
or U15748 (N_15748,N_10092,N_13005);
nand U15749 (N_15749,N_14136,N_10653);
xor U15750 (N_15750,N_11038,N_14452);
and U15751 (N_15751,N_14581,N_13030);
nand U15752 (N_15752,N_14113,N_11163);
or U15753 (N_15753,N_10366,N_13197);
and U15754 (N_15754,N_12319,N_11968);
nor U15755 (N_15755,N_11440,N_13733);
xor U15756 (N_15756,N_14786,N_12639);
nor U15757 (N_15757,N_13490,N_10258);
xnor U15758 (N_15758,N_11876,N_11662);
nor U15759 (N_15759,N_14005,N_11617);
nand U15760 (N_15760,N_10361,N_12292);
nor U15761 (N_15761,N_14784,N_10101);
nor U15762 (N_15762,N_12376,N_10354);
nor U15763 (N_15763,N_14737,N_10517);
and U15764 (N_15764,N_13631,N_12409);
xnor U15765 (N_15765,N_12007,N_11736);
and U15766 (N_15766,N_11551,N_13855);
or U15767 (N_15767,N_13206,N_10241);
or U15768 (N_15768,N_12401,N_13740);
or U15769 (N_15769,N_14413,N_11769);
nand U15770 (N_15770,N_11094,N_12550);
and U15771 (N_15771,N_11267,N_10906);
or U15772 (N_15772,N_12091,N_13725);
xnor U15773 (N_15773,N_12209,N_10994);
xor U15774 (N_15774,N_11668,N_13051);
and U15775 (N_15775,N_10028,N_10854);
xor U15776 (N_15776,N_13793,N_14433);
nand U15777 (N_15777,N_11052,N_14580);
xnor U15778 (N_15778,N_14789,N_11569);
xor U15779 (N_15779,N_10703,N_10041);
or U15780 (N_15780,N_10433,N_10840);
nor U15781 (N_15781,N_12301,N_10033);
and U15782 (N_15782,N_12699,N_10170);
or U15783 (N_15783,N_11845,N_12406);
nand U15784 (N_15784,N_11775,N_10959);
and U15785 (N_15785,N_10530,N_14327);
and U15786 (N_15786,N_13122,N_12933);
nand U15787 (N_15787,N_13552,N_11129);
or U15788 (N_15788,N_11345,N_11695);
and U15789 (N_15789,N_12859,N_11529);
nand U15790 (N_15790,N_10228,N_13119);
and U15791 (N_15791,N_12483,N_10003);
nand U15792 (N_15792,N_10119,N_12113);
and U15793 (N_15793,N_14550,N_11053);
or U15794 (N_15794,N_13727,N_11412);
nor U15795 (N_15795,N_14835,N_14083);
or U15796 (N_15796,N_11363,N_13977);
and U15797 (N_15797,N_13263,N_12491);
and U15798 (N_15798,N_12831,N_10295);
nor U15799 (N_15799,N_10052,N_10254);
nand U15800 (N_15800,N_13891,N_12402);
or U15801 (N_15801,N_10020,N_11253);
and U15802 (N_15802,N_12729,N_13158);
or U15803 (N_15803,N_12616,N_10622);
or U15804 (N_15804,N_13619,N_11380);
nor U15805 (N_15805,N_14101,N_13315);
xor U15806 (N_15806,N_13411,N_11263);
and U15807 (N_15807,N_11939,N_11749);
nand U15808 (N_15808,N_10110,N_11151);
nor U15809 (N_15809,N_13326,N_12024);
and U15810 (N_15810,N_13909,N_11629);
nand U15811 (N_15811,N_12686,N_10045);
xnor U15812 (N_15812,N_11350,N_14041);
nand U15813 (N_15813,N_10277,N_14691);
or U15814 (N_15814,N_11592,N_13187);
xnor U15815 (N_15815,N_10993,N_13027);
and U15816 (N_15816,N_10389,N_10669);
xnor U15817 (N_15817,N_14759,N_11781);
xnor U15818 (N_15818,N_10001,N_10269);
nand U15819 (N_15819,N_10205,N_11922);
nor U15820 (N_15820,N_14676,N_12586);
and U15821 (N_15821,N_13385,N_14638);
nand U15822 (N_15822,N_13723,N_11083);
or U15823 (N_15823,N_14004,N_13629);
or U15824 (N_15824,N_14107,N_10419);
nand U15825 (N_15825,N_12403,N_12663);
and U15826 (N_15826,N_12795,N_14543);
nor U15827 (N_15827,N_11288,N_11924);
and U15828 (N_15828,N_10784,N_12836);
nand U15829 (N_15829,N_11853,N_14429);
xnor U15830 (N_15830,N_10766,N_12337);
and U15831 (N_15831,N_11767,N_14539);
xor U15832 (N_15832,N_14767,N_12383);
xor U15833 (N_15833,N_10635,N_12681);
or U15834 (N_15834,N_11417,N_14300);
and U15835 (N_15835,N_13931,N_14800);
xnor U15836 (N_15836,N_12026,N_14625);
xor U15837 (N_15837,N_11469,N_13554);
nand U15838 (N_15838,N_10796,N_10240);
nand U15839 (N_15839,N_10852,N_10649);
nor U15840 (N_15840,N_11658,N_14028);
nor U15841 (N_15841,N_10546,N_10881);
nor U15842 (N_15842,N_14679,N_14227);
nor U15843 (N_15843,N_10186,N_10655);
and U15844 (N_15844,N_10331,N_12433);
xnor U15845 (N_15845,N_14162,N_11950);
xnor U15846 (N_15846,N_11104,N_11998);
or U15847 (N_15847,N_10802,N_14139);
or U15848 (N_15848,N_13331,N_14899);
and U15849 (N_15849,N_13823,N_10496);
xor U15850 (N_15850,N_14704,N_10273);
xnor U15851 (N_15851,N_10725,N_12562);
or U15852 (N_15852,N_13653,N_10722);
nand U15853 (N_15853,N_13839,N_14188);
or U15854 (N_15854,N_11420,N_11407);
xor U15855 (N_15855,N_10409,N_11254);
and U15856 (N_15856,N_12576,N_10207);
or U15857 (N_15857,N_11154,N_14080);
or U15858 (N_15858,N_14241,N_10093);
or U15859 (N_15859,N_11901,N_14496);
nand U15860 (N_15860,N_12506,N_13841);
and U15861 (N_15861,N_13730,N_14406);
or U15862 (N_15862,N_14761,N_12719);
and U15863 (N_15863,N_12157,N_14521);
xnor U15864 (N_15864,N_13919,N_12590);
nand U15865 (N_15865,N_12606,N_11874);
nor U15866 (N_15866,N_10673,N_11086);
nor U15867 (N_15867,N_10445,N_11182);
nand U15868 (N_15868,N_13019,N_11944);
and U15869 (N_15869,N_14629,N_13687);
and U15870 (N_15870,N_12011,N_13749);
and U15871 (N_15871,N_11999,N_14533);
xnor U15872 (N_15872,N_11631,N_14230);
and U15873 (N_15873,N_13966,N_11230);
nand U15874 (N_15874,N_13352,N_14256);
nand U15875 (N_15875,N_11635,N_10519);
nand U15876 (N_15876,N_10662,N_11377);
xnor U15877 (N_15877,N_12910,N_14526);
nand U15878 (N_15878,N_14116,N_13513);
nand U15879 (N_15879,N_13424,N_14709);
or U15880 (N_15880,N_12552,N_12994);
or U15881 (N_15881,N_11547,N_14651);
nand U15882 (N_15882,N_12381,N_11064);
and U15883 (N_15883,N_12152,N_12931);
nor U15884 (N_15884,N_14032,N_13141);
nor U15885 (N_15885,N_13882,N_13927);
xor U15886 (N_15886,N_13487,N_13403);
nor U15887 (N_15887,N_14092,N_10455);
nor U15888 (N_15888,N_11485,N_13232);
xor U15889 (N_15889,N_11550,N_12126);
or U15890 (N_15890,N_11506,N_12038);
or U15891 (N_15891,N_12043,N_13688);
nand U15892 (N_15892,N_13600,N_14797);
nor U15893 (N_15893,N_11756,N_14808);
nand U15894 (N_15894,N_11213,N_12951);
or U15895 (N_15895,N_12981,N_12099);
nor U15896 (N_15896,N_11118,N_10570);
nand U15897 (N_15897,N_11480,N_11681);
nand U15898 (N_15898,N_13406,N_14916);
nor U15899 (N_15899,N_11957,N_11403);
nand U15900 (N_15900,N_14644,N_14765);
xnor U15901 (N_15901,N_10971,N_12852);
xnor U15902 (N_15902,N_12201,N_14480);
xor U15903 (N_15903,N_14184,N_12630);
xnor U15904 (N_15904,N_12667,N_13015);
nand U15905 (N_15905,N_10544,N_14242);
nor U15906 (N_15906,N_10335,N_13973);
or U15907 (N_15907,N_13642,N_11776);
xnor U15908 (N_15908,N_10905,N_13524);
nor U15909 (N_15909,N_12815,N_10368);
nor U15910 (N_15910,N_13341,N_10687);
and U15911 (N_15911,N_13984,N_11783);
xnor U15912 (N_15912,N_13400,N_12446);
xor U15913 (N_15913,N_10387,N_12986);
or U15914 (N_15914,N_13092,N_12255);
nand U15915 (N_15915,N_10372,N_10731);
and U15916 (N_15916,N_11923,N_14822);
nand U15917 (N_15917,N_11109,N_14168);
nor U15918 (N_15918,N_14711,N_10247);
xor U15919 (N_15919,N_11032,N_11908);
nor U15920 (N_15920,N_13936,N_14439);
or U15921 (N_15921,N_11552,N_10716);
xor U15922 (N_15922,N_11077,N_14054);
and U15923 (N_15923,N_14426,N_11765);
or U15924 (N_15924,N_11510,N_13566);
nand U15925 (N_15925,N_11896,N_12495);
or U15926 (N_15926,N_12005,N_13879);
nor U15927 (N_15927,N_14115,N_10235);
nor U15928 (N_15928,N_10751,N_10336);
nor U15929 (N_15929,N_11513,N_10928);
nor U15930 (N_15930,N_14552,N_14665);
and U15931 (N_15931,N_11084,N_13079);
and U15932 (N_15932,N_12351,N_10324);
xnor U15933 (N_15933,N_14348,N_13316);
nand U15934 (N_15934,N_10592,N_13404);
nand U15935 (N_15935,N_10771,N_13933);
nor U15936 (N_15936,N_12174,N_13324);
and U15937 (N_15937,N_13779,N_13262);
xor U15938 (N_15938,N_12614,N_10275);
nand U15939 (N_15939,N_12565,N_10615);
and U15940 (N_15940,N_13522,N_12085);
xnor U15941 (N_15941,N_12193,N_12964);
and U15942 (N_15942,N_13772,N_14169);
nand U15943 (N_15943,N_10350,N_11037);
xnor U15944 (N_15944,N_10261,N_14358);
nor U15945 (N_15945,N_11081,N_13661);
xor U15946 (N_15946,N_14114,N_14286);
nand U15947 (N_15947,N_11188,N_14154);
xor U15948 (N_15948,N_12262,N_13087);
xnor U15949 (N_15949,N_11840,N_10233);
nor U15950 (N_15950,N_13978,N_10679);
xor U15951 (N_15951,N_12150,N_13390);
or U15952 (N_15952,N_10182,N_11527);
or U15953 (N_15953,N_11181,N_12142);
xor U15954 (N_15954,N_13698,N_12385);
and U15955 (N_15955,N_10770,N_11012);
nand U15956 (N_15956,N_12802,N_10631);
xnor U15957 (N_15957,N_10185,N_11018);
nor U15958 (N_15958,N_10327,N_13053);
xnor U15959 (N_15959,N_10730,N_11821);
nand U15960 (N_15960,N_13414,N_12295);
and U15961 (N_15961,N_14794,N_10794);
nand U15962 (N_15962,N_11257,N_14908);
and U15963 (N_15963,N_14592,N_12084);
xnor U15964 (N_15964,N_12060,N_13282);
xor U15965 (N_15965,N_10938,N_11185);
xnor U15966 (N_15966,N_12930,N_11069);
nand U15967 (N_15967,N_10257,N_14957);
nor U15968 (N_15968,N_13054,N_13646);
nor U15969 (N_15969,N_14668,N_10289);
nor U15970 (N_15970,N_14748,N_12012);
nand U15971 (N_15971,N_14726,N_14186);
nor U15972 (N_15972,N_12429,N_11372);
xnor U15973 (N_15973,N_13208,N_13777);
xnor U15974 (N_15974,N_13133,N_13614);
xor U15975 (N_15975,N_12706,N_13212);
xor U15976 (N_15976,N_10202,N_11258);
and U15977 (N_15977,N_13016,N_12809);
nor U15978 (N_15978,N_10884,N_12159);
nand U15979 (N_15979,N_10288,N_14717);
or U15980 (N_15980,N_14165,N_11660);
nor U15981 (N_15981,N_11450,N_14585);
and U15982 (N_15982,N_13620,N_10502);
or U15983 (N_15983,N_13327,N_13254);
or U15984 (N_15984,N_10323,N_14420);
nand U15985 (N_15985,N_13521,N_14275);
nor U15986 (N_15986,N_14646,N_10096);
or U15987 (N_15987,N_13636,N_11107);
or U15988 (N_15988,N_11033,N_12896);
or U15989 (N_15989,N_12708,N_11004);
or U15990 (N_15990,N_12520,N_11969);
or U15991 (N_15991,N_13260,N_12200);
xnor U15992 (N_15992,N_12370,N_14852);
and U15993 (N_15993,N_11279,N_10183);
nand U15994 (N_15994,N_14247,N_13182);
nand U15995 (N_15995,N_13183,N_12101);
xor U15996 (N_15996,N_11194,N_12344);
xor U15997 (N_15997,N_11009,N_10480);
and U15998 (N_15998,N_10358,N_13289);
nor U15999 (N_15999,N_11050,N_12207);
and U16000 (N_16000,N_13370,N_11023);
or U16001 (N_16001,N_12522,N_12678);
xnor U16002 (N_16002,N_14344,N_10404);
xnor U16003 (N_16003,N_13726,N_11725);
xnor U16004 (N_16004,N_13484,N_14029);
nand U16005 (N_16005,N_13055,N_14499);
xor U16006 (N_16006,N_12415,N_10105);
nor U16007 (N_16007,N_10365,N_10337);
and U16008 (N_16008,N_12138,N_10734);
nand U16009 (N_16009,N_13473,N_10540);
xor U16010 (N_16010,N_10495,N_11994);
xor U16011 (N_16011,N_10597,N_14688);
nand U16012 (N_16012,N_12432,N_10099);
nand U16013 (N_16013,N_11223,N_11883);
or U16014 (N_16014,N_10591,N_14213);
and U16015 (N_16015,N_12682,N_12869);
xor U16016 (N_16016,N_11158,N_13115);
or U16017 (N_16017,N_12443,N_13278);
nand U16018 (N_16018,N_13125,N_10726);
nand U16019 (N_16019,N_14746,N_13920);
and U16020 (N_16020,N_13679,N_11911);
and U16021 (N_16021,N_10822,N_11887);
and U16022 (N_16022,N_14343,N_13060);
nand U16023 (N_16023,N_14714,N_11003);
xor U16024 (N_16024,N_10846,N_11088);
or U16025 (N_16025,N_11828,N_12094);
or U16026 (N_16026,N_13520,N_12829);
and U16027 (N_16027,N_12176,N_13100);
or U16028 (N_16028,N_13567,N_11867);
or U16029 (N_16029,N_13151,N_13804);
nor U16030 (N_16030,N_14862,N_13694);
and U16031 (N_16031,N_11784,N_10990);
and U16032 (N_16032,N_10122,N_11962);
or U16033 (N_16033,N_13419,N_11512);
nor U16034 (N_16034,N_10319,N_10181);
nor U16035 (N_16035,N_11719,N_10975);
and U16036 (N_16036,N_13809,N_12140);
nand U16037 (N_16037,N_11272,N_12260);
or U16038 (N_16038,N_10569,N_14099);
or U16039 (N_16039,N_10534,N_10023);
nor U16040 (N_16040,N_11291,N_13611);
xor U16041 (N_16041,N_10626,N_11785);
and U16042 (N_16042,N_14076,N_14869);
xor U16043 (N_16043,N_12482,N_10579);
nand U16044 (N_16044,N_11729,N_14394);
xnor U16045 (N_16045,N_12303,N_12078);
xor U16046 (N_16046,N_14517,N_10814);
and U16047 (N_16047,N_14994,N_12646);
and U16048 (N_16048,N_11947,N_13156);
xor U16049 (N_16049,N_12973,N_10617);
or U16050 (N_16050,N_11418,N_14618);
and U16051 (N_16051,N_11974,N_11720);
nand U16052 (N_16052,N_11649,N_14661);
nand U16053 (N_16053,N_10215,N_12340);
nor U16054 (N_16054,N_14595,N_10484);
xor U16055 (N_16055,N_14482,N_14219);
and U16056 (N_16056,N_13503,N_10478);
nor U16057 (N_16057,N_11082,N_11669);
nand U16058 (N_16058,N_13606,N_10329);
nor U16059 (N_16059,N_12508,N_13759);
xnor U16060 (N_16060,N_10743,N_13439);
nand U16061 (N_16061,N_12805,N_11156);
nand U16062 (N_16062,N_10922,N_10079);
xnor U16063 (N_16063,N_10717,N_14697);
nor U16064 (N_16064,N_12379,N_11693);
xor U16065 (N_16065,N_13154,N_10769);
nor U16066 (N_16066,N_10684,N_11680);
and U16067 (N_16067,N_13496,N_12758);
xor U16068 (N_16068,N_12753,N_10714);
xor U16069 (N_16069,N_13673,N_13389);
or U16070 (N_16070,N_13200,N_14434);
and U16071 (N_16071,N_11244,N_14948);
xor U16072 (N_16072,N_10853,N_14215);
xor U16073 (N_16073,N_14583,N_13699);
and U16074 (N_16074,N_13960,N_11414);
or U16075 (N_16075,N_11462,N_10308);
and U16076 (N_16076,N_14969,N_12053);
or U16077 (N_16077,N_12361,N_14237);
nor U16078 (N_16078,N_13604,N_11888);
and U16079 (N_16079,N_14736,N_13969);
or U16080 (N_16080,N_11593,N_14445);
nand U16081 (N_16081,N_14615,N_14815);
nor U16082 (N_16082,N_11815,N_12744);
nor U16083 (N_16083,N_13388,N_13959);
or U16084 (N_16084,N_11739,N_12569);
nor U16085 (N_16085,N_13334,N_12345);
xor U16086 (N_16086,N_14974,N_10529);
xnor U16087 (N_16087,N_14540,N_14816);
xnor U16088 (N_16088,N_10680,N_12302);
nand U16089 (N_16089,N_12238,N_14010);
and U16090 (N_16090,N_11227,N_13309);
nor U16091 (N_16091,N_14084,N_11941);
and U16092 (N_16092,N_10048,N_10457);
nor U16093 (N_16093,N_14624,N_11906);
xor U16094 (N_16094,N_11195,N_13607);
xnor U16095 (N_16095,N_14143,N_12736);
or U16096 (N_16096,N_10646,N_14253);
xor U16097 (N_16097,N_13743,N_12339);
nor U16098 (N_16098,N_12898,N_13963);
xor U16099 (N_16099,N_13888,N_12881);
xnor U16100 (N_16100,N_11278,N_10931);
and U16101 (N_16101,N_11630,N_10270);
nor U16102 (N_16102,N_10908,N_10594);
nand U16103 (N_16103,N_12258,N_11852);
nor U16104 (N_16104,N_10349,N_14284);
xnor U16105 (N_16105,N_10641,N_10745);
nand U16106 (N_16106,N_12212,N_14097);
xor U16107 (N_16107,N_14997,N_13307);
and U16108 (N_16108,N_10063,N_11786);
and U16109 (N_16109,N_12111,N_11008);
nand U16110 (N_16110,N_12691,N_14209);
nor U16111 (N_16111,N_13796,N_12591);
nor U16112 (N_16112,N_14422,N_11747);
and U16113 (N_16113,N_11805,N_10321);
nand U16114 (N_16114,N_10892,N_13085);
nand U16115 (N_16115,N_10015,N_10347);
nor U16116 (N_16116,N_13010,N_13569);
nand U16117 (N_16117,N_10595,N_10516);
or U16118 (N_16118,N_14961,N_10825);
or U16119 (N_16119,N_13176,N_13457);
nor U16120 (N_16120,N_12730,N_13153);
and U16121 (N_16121,N_12618,N_11142);
nor U16122 (N_16122,N_11348,N_10125);
xor U16123 (N_16123,N_14164,N_11357);
xor U16124 (N_16124,N_12479,N_12703);
nor U16125 (N_16125,N_13169,N_12769);
nor U16126 (N_16126,N_14141,N_10057);
xnor U16127 (N_16127,N_14906,N_14245);
xnor U16128 (N_16128,N_11005,N_12722);
and U16129 (N_16129,N_11312,N_13923);
and U16130 (N_16130,N_12558,N_12709);
and U16131 (N_16131,N_10658,N_11878);
nand U16132 (N_16132,N_13802,N_13548);
xor U16133 (N_16133,N_14312,N_13675);
nor U16134 (N_16134,N_14322,N_13618);
and U16135 (N_16135,N_11808,N_10902);
or U16136 (N_16136,N_14522,N_14475);
nor U16137 (N_16137,N_10693,N_13669);
and U16138 (N_16138,N_14240,N_11899);
nor U16139 (N_16139,N_10883,N_13356);
nand U16140 (N_16140,N_14928,N_14036);
xor U16141 (N_16141,N_13354,N_14802);
nand U16142 (N_16142,N_14308,N_11953);
xnor U16143 (N_16143,N_13516,N_13336);
and U16144 (N_16144,N_14494,N_13216);
or U16145 (N_16145,N_11587,N_13782);
or U16146 (N_16146,N_13144,N_10561);
xor U16147 (N_16147,N_10790,N_11204);
nor U16148 (N_16148,N_11605,N_14952);
nand U16149 (N_16149,N_12589,N_10000);
xor U16150 (N_16150,N_13318,N_11966);
or U16151 (N_16151,N_13792,N_10986);
nor U16152 (N_16152,N_13916,N_12755);
and U16153 (N_16153,N_12925,N_10310);
xnor U16154 (N_16154,N_11387,N_12059);
and U16155 (N_16155,N_14557,N_13808);
and U16156 (N_16156,N_14355,N_14306);
nor U16157 (N_16157,N_13538,N_11777);
nor U16158 (N_16158,N_13310,N_11509);
nand U16159 (N_16159,N_14660,N_14255);
nor U16160 (N_16160,N_13396,N_10416);
or U16161 (N_16161,N_14689,N_12046);
xor U16162 (N_16162,N_12033,N_12505);
nand U16163 (N_16163,N_10268,N_13338);
xor U16164 (N_16164,N_11616,N_13422);
xnor U16165 (N_16165,N_13415,N_12924);
or U16166 (N_16166,N_14775,N_10837);
or U16167 (N_16167,N_14386,N_12317);
or U16168 (N_16168,N_14234,N_13983);
nor U16169 (N_16169,N_13167,N_11190);
nand U16170 (N_16170,N_10053,N_11731);
nand U16171 (N_16171,N_13241,N_14100);
nor U16172 (N_16172,N_12888,N_14073);
and U16173 (N_16173,N_10528,N_11111);
nand U16174 (N_16174,N_14903,N_13797);
nor U16175 (N_16175,N_13127,N_13592);
nor U16176 (N_16176,N_12181,N_10262);
nand U16177 (N_16177,N_14518,N_14523);
nor U16178 (N_16178,N_14671,N_12775);
and U16179 (N_16179,N_13044,N_11758);
nand U16180 (N_16180,N_14291,N_13770);
or U16181 (N_16181,N_10584,N_12366);
and U16182 (N_16182,N_13235,N_14200);
or U16183 (N_16183,N_14937,N_10084);
xor U16184 (N_16184,N_11024,N_12438);
or U16185 (N_16185,N_13410,N_14472);
or U16186 (N_16186,N_12184,N_13308);
and U16187 (N_16187,N_14220,N_14166);
nor U16188 (N_16188,N_10140,N_11855);
nand U16189 (N_16189,N_13031,N_13588);
and U16190 (N_16190,N_11255,N_13088);
nand U16191 (N_16191,N_13123,N_14683);
and U16192 (N_16192,N_14484,N_13281);
xnor U16193 (N_16193,N_10713,N_11757);
nor U16194 (N_16194,N_14889,N_14972);
and U16195 (N_16195,N_14443,N_12232);
nor U16196 (N_16196,N_13131,N_10772);
and U16197 (N_16197,N_13106,N_14013);
and U16198 (N_16198,N_10609,N_10510);
nor U16199 (N_16199,N_11294,N_14085);
or U16200 (N_16200,N_14098,N_12472);
nor U16201 (N_16201,N_13456,N_14378);
nand U16202 (N_16202,N_10807,N_12670);
nor U16203 (N_16203,N_13425,N_13397);
and U16204 (N_16204,N_14198,N_14153);
and U16205 (N_16205,N_12694,N_12546);
or U16206 (N_16206,N_12397,N_13641);
nand U16207 (N_16207,N_11292,N_12760);
nand U16208 (N_16208,N_11545,N_13438);
nand U16209 (N_16209,N_11210,N_12988);
or U16210 (N_16210,N_10089,N_11001);
nor U16211 (N_16211,N_11802,N_13245);
xor U16212 (N_16212,N_14980,N_13574);
xor U16213 (N_16213,N_12874,N_13573);
or U16214 (N_16214,N_11772,N_12787);
xor U16215 (N_16215,N_14440,N_11197);
nor U16216 (N_16216,N_12972,N_11728);
xnor U16217 (N_16217,N_11054,N_11307);
and U16218 (N_16218,N_14567,N_13940);
xor U16219 (N_16219,N_11308,N_13297);
nor U16220 (N_16220,N_12952,N_12115);
nor U16221 (N_16221,N_14449,N_10875);
nand U16222 (N_16222,N_12083,N_14151);
xnor U16223 (N_16223,N_11123,N_12704);
xor U16224 (N_16224,N_12808,N_14432);
nand U16225 (N_16225,N_10643,N_10760);
xnor U16226 (N_16226,N_10469,N_11058);
xnor U16227 (N_16227,N_10562,N_10843);
nand U16228 (N_16228,N_12318,N_12561);
and U16229 (N_16229,N_13249,N_14740);
nor U16230 (N_16230,N_12430,N_12492);
and U16231 (N_16231,N_10226,N_12687);
nand U16232 (N_16232,N_10657,N_10503);
xnor U16233 (N_16233,N_13873,N_13791);
nand U16234 (N_16234,N_13526,N_10292);
nor U16235 (N_16235,N_13939,N_10113);
and U16236 (N_16236,N_13171,N_14778);
and U16237 (N_16237,N_13902,N_14924);
nor U16238 (N_16238,N_13288,N_13003);
nand U16239 (N_16239,N_12601,N_14015);
nor U16240 (N_16240,N_13394,N_10548);
xor U16241 (N_16241,N_13312,N_11745);
and U16242 (N_16242,N_13584,N_14260);
or U16243 (N_16243,N_14613,N_14659);
and U16244 (N_16244,N_14185,N_10405);
nand U16245 (N_16245,N_14896,N_14701);
xor U16246 (N_16246,N_13843,N_11801);
nor U16247 (N_16247,N_11179,N_14130);
and U16248 (N_16248,N_13483,N_12529);
or U16249 (N_16249,N_12490,N_10309);
and U16250 (N_16250,N_13192,N_12649);
xnor U16251 (N_16251,N_13781,N_11287);
nand U16252 (N_16252,N_10377,N_12027);
and U16253 (N_16253,N_14640,N_12167);
nor U16254 (N_16254,N_13271,N_12117);
nand U16255 (N_16255,N_12532,N_10082);
nor U16256 (N_16256,N_13773,N_13651);
or U16257 (N_16257,N_12257,N_11233);
nor U16258 (N_16258,N_12256,N_11404);
and U16259 (N_16259,N_12281,N_13547);
xnor U16260 (N_16260,N_11316,N_13138);
nor U16261 (N_16261,N_10107,N_11880);
nand U16262 (N_16262,N_13905,N_14844);
or U16263 (N_16263,N_14891,N_13113);
nand U16264 (N_16264,N_11314,N_13335);
nand U16265 (N_16265,N_11234,N_13114);
nand U16266 (N_16266,N_12456,N_14047);
and U16267 (N_16267,N_13957,N_12880);
nor U16268 (N_16268,N_10568,N_14374);
xnor U16269 (N_16269,N_14710,N_12353);
xor U16270 (N_16270,N_10299,N_13728);
nand U16271 (N_16271,N_11654,N_11061);
nand U16272 (N_16272,N_11386,N_14984);
or U16273 (N_16273,N_10574,N_14180);
and U16274 (N_16274,N_11269,N_11750);
xor U16275 (N_16275,N_14828,N_11955);
and U16276 (N_16276,N_13735,N_12105);
nor U16277 (N_16277,N_12537,N_12768);
or U16278 (N_16278,N_11318,N_13135);
xor U16279 (N_16279,N_13001,N_10834);
xnor U16280 (N_16280,N_14133,N_13964);
nand U16281 (N_16281,N_14864,N_10762);
nand U16282 (N_16282,N_13599,N_13466);
or U16283 (N_16283,N_14853,N_11503);
and U16284 (N_16284,N_10933,N_12611);
or U16285 (N_16285,N_10342,N_13240);
or U16286 (N_16286,N_13374,N_13764);
or U16287 (N_16287,N_13033,N_10345);
xor U16288 (N_16288,N_13495,N_14203);
xnor U16289 (N_16289,N_11264,N_11768);
or U16290 (N_16290,N_13471,N_11346);
nand U16291 (N_16291,N_14968,N_12205);
or U16292 (N_16292,N_12583,N_12856);
xor U16293 (N_16293,N_10373,N_12651);
nor U16294 (N_16294,N_11666,N_14295);
xor U16295 (N_16295,N_14500,N_11692);
nand U16296 (N_16296,N_12912,N_13831);
or U16297 (N_16297,N_14161,N_13076);
xor U16298 (N_16298,N_12315,N_11531);
nand U16299 (N_16299,N_12631,N_13850);
and U16300 (N_16300,N_14712,N_14885);
xor U16301 (N_16301,N_12485,N_11589);
nor U16302 (N_16302,N_13372,N_13355);
nor U16303 (N_16303,N_12900,N_10421);
and U16304 (N_16304,N_12372,N_10106);
or U16305 (N_16305,N_13951,N_10876);
nor U16306 (N_16306,N_11869,N_10925);
xnor U16307 (N_16307,N_10149,N_13157);
nand U16308 (N_16308,N_11511,N_13407);
nand U16309 (N_16309,N_12675,N_10088);
nand U16310 (N_16310,N_12068,N_13222);
xnor U16311 (N_16311,N_12999,N_12074);
xnor U16312 (N_16312,N_14249,N_12056);
or U16313 (N_16313,N_14398,N_13681);
nor U16314 (N_16314,N_10753,N_10551);
and U16315 (N_16315,N_14269,N_14120);
nand U16316 (N_16316,N_11349,N_12733);
xor U16317 (N_16317,N_14586,N_13556);
or U16318 (N_16318,N_12777,N_12875);
nand U16319 (N_16319,N_14063,N_14365);
and U16320 (N_16320,N_12221,N_14460);
and U16321 (N_16321,N_10322,N_11607);
or U16322 (N_16322,N_13815,N_14140);
nand U16323 (N_16323,N_10779,N_14339);
nor U16324 (N_16324,N_11434,N_12596);
nor U16325 (N_16325,N_10705,N_11992);
xor U16326 (N_16326,N_10863,N_10176);
nand U16327 (N_16327,N_11873,N_12335);
and U16328 (N_16328,N_13132,N_10995);
or U16329 (N_16329,N_14359,N_13775);
nor U16330 (N_16330,N_12275,N_10234);
nor U16331 (N_16331,N_13585,N_12892);
xnor U16332 (N_16332,N_14656,N_10666);
nand U16333 (N_16333,N_14780,N_13602);
nand U16334 (N_16334,N_13317,N_12470);
nand U16335 (N_16335,N_11727,N_14034);
and U16336 (N_16336,N_12820,N_12632);
nor U16337 (N_16337,N_14454,N_14681);
xor U16338 (N_16338,N_11456,N_12165);
xor U16339 (N_16339,N_14843,N_11020);
and U16340 (N_16340,N_11598,N_11889);
or U16341 (N_16341,N_11362,N_12650);
and U16342 (N_16342,N_10086,N_10511);
nor U16343 (N_16343,N_14105,N_10223);
nand U16344 (N_16344,N_14427,N_13720);
nand U16345 (N_16345,N_13670,N_12130);
xor U16346 (N_16346,N_12547,N_10167);
and U16347 (N_16347,N_12800,N_14684);
xnor U16348 (N_16348,N_10374,N_11139);
nand U16349 (N_16349,N_14459,N_11400);
nand U16350 (N_16350,N_13664,N_12516);
nor U16351 (N_16351,N_13702,N_11105);
nand U16352 (N_16352,N_14048,N_11735);
or U16353 (N_16353,N_10583,N_10977);
and U16354 (N_16354,N_13613,N_12080);
xor U16355 (N_16355,N_12987,N_11341);
nor U16356 (N_16356,N_14963,N_10800);
xnor U16357 (N_16357,N_10921,N_12246);
nand U16358 (N_16358,N_14870,N_11954);
xnor U16359 (N_16359,N_13766,N_11334);
nor U16360 (N_16360,N_11864,N_13121);
xnor U16361 (N_16361,N_12941,N_14641);
and U16362 (N_16362,N_10438,N_13091);
or U16363 (N_16363,N_11276,N_12846);
xor U16364 (N_16364,N_10047,N_10944);
xor U16365 (N_16365,N_11178,N_10757);
xor U16366 (N_16366,N_14109,N_11426);
nor U16367 (N_16367,N_14788,N_13910);
xnor U16368 (N_16368,N_10535,N_12527);
xnor U16369 (N_16369,N_12737,N_12354);
xor U16370 (N_16370,N_11653,N_12288);
or U16371 (N_16371,N_11644,N_10483);
and U16372 (N_16372,N_12984,N_12740);
xnor U16373 (N_16373,N_10831,N_13452);
or U16374 (N_16374,N_14868,N_10157);
or U16375 (N_16375,N_14760,N_14019);
xor U16376 (N_16376,N_13491,N_12426);
nor U16377 (N_16377,N_13442,N_13748);
or U16378 (N_16378,N_13803,N_13564);
nor U16379 (N_16379,N_13287,N_11289);
nor U16380 (N_16380,N_10777,N_14576);
nand U16381 (N_16381,N_12216,N_12597);
and U16382 (N_16382,N_12211,N_11814);
nor U16383 (N_16383,N_11526,N_12978);
nor U16384 (N_16384,N_10909,N_14122);
nand U16385 (N_16385,N_10364,N_13364);
or U16386 (N_16386,N_14720,N_12322);
nand U16387 (N_16387,N_10196,N_12280);
nor U16388 (N_16388,N_13002,N_14648);
nand U16389 (N_16389,N_13578,N_11583);
nand U16390 (N_16390,N_10541,N_13248);
nor U16391 (N_16391,N_11266,N_11663);
nor U16392 (N_16392,N_10408,N_13373);
xor U16393 (N_16393,N_11219,N_13103);
xnor U16394 (N_16394,N_11504,N_12643);
or U16395 (N_16395,N_11313,N_10917);
nand U16396 (N_16396,N_12031,N_14457);
nor U16397 (N_16397,N_12419,N_10676);
xnor U16398 (N_16398,N_12956,N_12732);
and U16399 (N_16399,N_13913,N_12134);
xor U16400 (N_16400,N_13066,N_12751);
xnor U16401 (N_16401,N_10870,N_11256);
nor U16402 (N_16402,N_12542,N_12041);
and U16403 (N_16403,N_10767,N_10586);
or U16404 (N_16404,N_14014,N_13630);
or U16405 (N_16405,N_12153,N_14555);
nand U16406 (N_16406,N_12265,N_13918);
and U16407 (N_16407,N_13102,N_11566);
nor U16408 (N_16408,N_13540,N_12348);
and U16409 (N_16409,N_13753,N_14855);
nor U16410 (N_16410,N_14910,N_12788);
nor U16411 (N_16411,N_10154,N_14384);
xor U16412 (N_16412,N_11448,N_11539);
or U16413 (N_16413,N_11176,N_13059);
nand U16414 (N_16414,N_14566,N_14318);
nand U16415 (N_16415,N_13991,N_11990);
and U16416 (N_16416,N_13188,N_12131);
and U16417 (N_16417,N_11447,N_12635);
and U16418 (N_16418,N_10437,N_14967);
nor U16419 (N_16419,N_14628,N_11848);
xor U16420 (N_16420,N_12982,N_10670);
and U16421 (N_16421,N_12513,N_10142);
or U16422 (N_16422,N_12677,N_10897);
nand U16423 (N_16423,N_11359,N_14925);
or U16424 (N_16424,N_10217,N_11110);
nor U16425 (N_16425,N_14664,N_13900);
or U16426 (N_16426,N_13985,N_11656);
and U16427 (N_16427,N_12022,N_14860);
xnor U16428 (N_16428,N_13590,N_11124);
nor U16429 (N_16429,N_14718,N_10947);
nand U16430 (N_16430,N_10690,N_12282);
nand U16431 (N_16431,N_12224,N_14447);
nor U16432 (N_16432,N_10049,N_11927);
and U16433 (N_16433,N_11891,N_12963);
xnor U16434 (N_16434,N_10588,N_14865);
and U16435 (N_16435,N_10506,N_14123);
xnor U16436 (N_16436,N_11641,N_13912);
or U16437 (N_16437,N_13938,N_14934);
or U16438 (N_16438,N_11724,N_13395);
or U16439 (N_16439,N_14824,N_11080);
nor U16440 (N_16440,N_14866,N_12096);
nand U16441 (N_16441,N_14601,N_10385);
or U16442 (N_16442,N_12175,N_13663);
nand U16443 (N_16443,N_10244,N_13347);
xor U16444 (N_16444,N_14551,N_14134);
nand U16445 (N_16445,N_10058,N_14289);
nand U16446 (N_16446,N_10542,N_14617);
nor U16447 (N_16447,N_13889,N_12959);
xnor U16448 (N_16448,N_12047,N_12814);
nand U16449 (N_16449,N_10987,N_13502);
nor U16450 (N_16450,N_10700,N_11659);
or U16451 (N_16451,N_12029,N_13130);
and U16452 (N_16452,N_12833,N_11445);
nor U16453 (N_16453,N_14020,N_12380);
nand U16454 (N_16454,N_11961,N_12735);
nand U16455 (N_16455,N_10141,N_10585);
or U16456 (N_16456,N_11561,N_10911);
nor U16457 (N_16457,N_10378,N_10120);
nor U16458 (N_16458,N_13314,N_14991);
and U16459 (N_16459,N_14128,N_12498);
nor U16460 (N_16460,N_13941,N_13990);
or U16461 (N_16461,N_11721,N_13461);
nor U16462 (N_16462,N_11984,N_11175);
or U16463 (N_16463,N_12218,N_14279);
nand U16464 (N_16464,N_10958,N_14687);
and U16465 (N_16465,N_13644,N_14393);
or U16466 (N_16466,N_12018,N_10552);
and U16467 (N_16467,N_13826,N_12304);
or U16468 (N_16468,N_12530,N_12487);
and U16469 (N_16469,N_11517,N_12899);
xnor U16470 (N_16470,N_13559,N_13409);
nor U16471 (N_16471,N_12474,N_14171);
nor U16472 (N_16472,N_10417,N_11846);
and U16473 (N_16473,N_12273,N_10553);
nand U16474 (N_16474,N_14183,N_13391);
and U16475 (N_16475,N_10351,N_13111);
nand U16476 (N_16476,N_12544,N_12585);
or U16477 (N_16477,N_10491,N_12871);
xnor U16478 (N_16478,N_13837,N_12895);
nor U16479 (N_16479,N_10007,N_10100);
nand U16480 (N_16480,N_11683,N_14825);
or U16481 (N_16481,N_10008,N_14724);
xor U16482 (N_16482,N_12334,N_10109);
xnor U16483 (N_16483,N_10525,N_12902);
nand U16484 (N_16484,N_13893,N_11396);
nor U16485 (N_16485,N_10936,N_12548);
nor U16486 (N_16486,N_14923,N_13790);
nand U16487 (N_16487,N_12610,N_10450);
nor U16488 (N_16488,N_10037,N_13595);
nand U16489 (N_16489,N_11937,N_13417);
nor U16490 (N_16490,N_13117,N_12328);
or U16491 (N_16491,N_11196,N_14626);
or U16492 (N_16492,N_12001,N_12660);
and U16493 (N_16493,N_12528,N_12752);
nand U16494 (N_16494,N_13886,N_13186);
and U16495 (N_16495,N_13205,N_11217);
and U16496 (N_16496,N_12405,N_12645);
and U16497 (N_16497,N_13255,N_12488);
or U16498 (N_16498,N_10781,N_14783);
and U16499 (N_16499,N_11174,N_10616);
and U16500 (N_16500,N_12079,N_13535);
xor U16501 (N_16501,N_14468,N_13762);
or U16502 (N_16502,N_12233,N_14410);
nor U16503 (N_16503,N_11800,N_11356);
or U16504 (N_16504,N_12759,N_10681);
nor U16505 (N_16505,N_10330,N_14349);
xor U16506 (N_16506,N_14236,N_11040);
or U16507 (N_16507,N_14009,N_11446);
nor U16508 (N_16508,N_13832,N_10889);
xor U16509 (N_16509,N_11826,N_11554);
xnor U16510 (N_16510,N_13860,N_11488);
or U16511 (N_16511,N_10294,N_13237);
xnor U16512 (N_16512,N_12268,N_11670);
or U16513 (N_16513,N_12493,N_10076);
and U16514 (N_16514,N_11762,N_14673);
and U16515 (N_16515,N_14329,N_14749);
and U16516 (N_16516,N_10279,N_12781);
nand U16517 (N_16517,N_10571,N_11408);
xor U16518 (N_16518,N_13647,N_14787);
and U16519 (N_16519,N_13553,N_12263);
nor U16520 (N_16520,N_13075,N_10706);
or U16521 (N_16521,N_12783,N_11298);
xnor U16522 (N_16522,N_14272,N_14466);
and U16523 (N_16523,N_11495,N_11986);
nand U16524 (N_16524,N_10432,N_12065);
nor U16525 (N_16525,N_14104,N_14662);
or U16526 (N_16526,N_13353,N_10747);
nor U16527 (N_16527,N_14955,N_14837);
and U16528 (N_16528,N_14510,N_11921);
and U16529 (N_16529,N_10656,N_12626);
and U16530 (N_16530,N_14205,N_10391);
xnor U16531 (N_16531,N_11484,N_11558);
xor U16532 (N_16532,N_12600,N_12570);
xor U16533 (N_16533,N_12028,N_10175);
nor U16534 (N_16534,N_14415,N_12515);
nand U16535 (N_16535,N_13904,N_10139);
nor U16536 (N_16536,N_10978,N_13634);
nor U16537 (N_16537,N_11501,N_13608);
and U16538 (N_16538,N_12512,N_14497);
and U16539 (N_16539,N_13379,N_14781);
or U16540 (N_16540,N_11827,N_11191);
or U16541 (N_16541,N_10375,N_13101);
nor U16542 (N_16542,N_14532,N_12423);
nand U16543 (N_16543,N_11464,N_10318);
and U16544 (N_16544,N_10126,N_10565);
and U16545 (N_16545,N_10965,N_13947);
nor U16546 (N_16546,N_10960,N_13402);
nor U16547 (N_16547,N_12164,N_13551);
xor U16548 (N_16548,N_12696,N_10291);
nand U16549 (N_16549,N_13700,N_14345);
nand U16550 (N_16550,N_10360,N_12458);
nand U16551 (N_16551,N_10972,N_10671);
xor U16552 (N_16552,N_11239,N_14602);
xnor U16553 (N_16553,N_12036,N_13089);
nor U16554 (N_16554,N_11095,N_10017);
and U16555 (N_16555,N_14149,N_14491);
and U16556 (N_16556,N_12000,N_13512);
nand U16557 (N_16557,N_12818,N_11281);
nor U16558 (N_16558,N_13478,N_11323);
or U16559 (N_16559,N_14821,N_12813);
or U16560 (N_16560,N_14810,N_13529);
nand U16561 (N_16561,N_13266,N_13953);
and U16562 (N_16562,N_12514,N_13581);
or U16563 (N_16563,N_13536,N_13632);
and U16564 (N_16564,N_14597,N_12359);
and U16565 (N_16565,N_10746,N_11379);
nor U16566 (N_16566,N_14330,N_12247);
xnor U16567 (N_16567,N_11309,N_14382);
nor U16568 (N_16568,N_10821,N_12721);
or U16569 (N_16569,N_13501,N_13333);
and U16570 (N_16570,N_14851,N_13067);
and U16571 (N_16571,N_12374,N_11938);
nor U16572 (N_16572,N_11243,N_10010);
and U16573 (N_16573,N_12695,N_12347);
nand U16574 (N_16574,N_13231,N_10253);
nor U16575 (N_16575,N_14918,N_14024);
or U16576 (N_16576,N_11265,N_13376);
or U16577 (N_16577,N_14978,N_11333);
and U16578 (N_16578,N_13838,N_13861);
nor U16579 (N_16579,N_10930,N_11014);
or U16580 (N_16580,N_12599,N_14288);
nand U16581 (N_16581,N_11553,N_13322);
or U16582 (N_16582,N_12352,N_14854);
xnor U16583 (N_16583,N_13894,N_13363);
and U16584 (N_16584,N_12284,N_14723);
xor U16585 (N_16585,N_14527,N_12615);
nand U16586 (N_16586,N_13924,N_14587);
and U16587 (N_16587,N_14519,N_12789);
xnor U16588 (N_16588,N_11564,N_12139);
xor U16589 (N_16589,N_14769,N_12911);
xnor U16590 (N_16590,N_10721,N_10532);
or U16591 (N_16591,N_13623,N_14988);
xnor U16592 (N_16592,N_14031,N_11812);
xnor U16593 (N_16593,N_10029,N_14768);
xnor U16594 (N_16594,N_11557,N_12707);
nand U16595 (N_16595,N_13776,N_10533);
xnor U16596 (N_16596,N_13321,N_10488);
and U16597 (N_16597,N_13539,N_12563);
xnor U16598 (N_16598,N_12862,N_13914);
nor U16599 (N_16599,N_10160,N_12658);
xor U16600 (N_16600,N_13956,N_11337);
nor U16601 (N_16601,N_14371,N_12272);
nand U16602 (N_16602,N_11835,N_13870);
xor U16603 (N_16603,N_14639,N_12936);
xor U16604 (N_16604,N_13383,N_10151);
or U16605 (N_16605,N_14340,N_10891);
xnor U16606 (N_16606,N_11078,N_12278);
nand U16607 (N_16607,N_10648,N_12560);
xor U16608 (N_16608,N_14052,N_11570);
nor U16609 (N_16609,N_12995,N_10809);
xor U16610 (N_16610,N_10620,N_11437);
nor U16611 (N_16611,N_14643,N_14900);
nor U16612 (N_16612,N_14874,N_13000);
nand U16613 (N_16613,N_11753,N_11902);
nor U16614 (N_16614,N_14738,N_12511);
xor U16615 (N_16615,N_14959,N_13853);
nand U16616 (N_16616,N_11209,N_12507);
xor U16617 (N_16617,N_10102,N_12124);
or U16618 (N_16618,N_13120,N_10114);
nor U16619 (N_16619,N_13375,N_10624);
nand U16620 (N_16620,N_12727,N_10075);
nand U16621 (N_16621,N_14739,N_14584);
or U16622 (N_16622,N_11677,N_11838);
xor U16623 (N_16623,N_12672,N_12534);
nand U16624 (N_16624,N_12763,N_10832);
xor U16625 (N_16625,N_11045,N_13458);
nor U16626 (N_16626,N_12227,N_13291);
xnor U16627 (N_16627,N_12215,N_11113);
xnor U16628 (N_16628,N_10340,N_10664);
and U16629 (N_16629,N_11293,N_12386);
and U16630 (N_16630,N_11958,N_14627);
nor U16631 (N_16631,N_10399,N_13813);
nor U16632 (N_16632,N_10060,N_13178);
and U16633 (N_16633,N_14536,N_10232);
and U16634 (N_16634,N_13925,N_11494);
and U16635 (N_16635,N_12202,N_14383);
nor U16636 (N_16636,N_13747,N_12338);
nand U16637 (N_16637,N_12613,N_11718);
nand U16638 (N_16638,N_11839,N_10229);
nor U16639 (N_16639,N_13041,N_11229);
or U16640 (N_16640,N_13708,N_14777);
nand U16641 (N_16641,N_13643,N_12796);
nand U16642 (N_16642,N_13751,N_11376);
nor U16643 (N_16643,N_10918,N_13591);
and U16644 (N_16644,N_12414,N_14703);
nor U16645 (N_16645,N_14088,N_11740);
nand U16646 (N_16646,N_10071,N_10893);
nand U16647 (N_16647,N_10577,N_10633);
and U16648 (N_16648,N_10072,N_10968);
xor U16649 (N_16649,N_11627,N_12588);
and U16650 (N_16650,N_13988,N_14239);
and U16651 (N_16651,N_13430,N_13295);
nand U16652 (N_16652,N_14637,N_10296);
or U16653 (N_16653,N_14347,N_13655);
or U16654 (N_16654,N_13344,N_11996);
or U16655 (N_16655,N_14892,N_11296);
xnor U16656 (N_16656,N_13895,N_10208);
nor U16657 (N_16657,N_10256,N_14686);
and U16658 (N_16658,N_11461,N_13500);
nor U16659 (N_16659,N_11863,N_11006);
nand U16660 (N_16660,N_14462,N_13104);
and U16661 (N_16661,N_12799,N_12296);
or U16662 (N_16662,N_10260,N_14754);
or U16663 (N_16663,N_14873,N_11597);
nand U16664 (N_16664,N_11031,N_12465);
or U16665 (N_16665,N_11890,N_13378);
or U16666 (N_16666,N_12521,N_14112);
nor U16667 (N_16667,N_11766,N_14841);
nor U16668 (N_16668,N_10341,N_10026);
nand U16669 (N_16669,N_12336,N_13788);
and U16670 (N_16670,N_10621,N_14966);
or U16671 (N_16671,N_14061,N_10801);
or U16672 (N_16672,N_11979,N_10239);
nor U16673 (N_16673,N_12197,N_10290);
or U16674 (N_16674,N_13459,N_12481);
nand U16675 (N_16675,N_14046,N_12194);
nand U16676 (N_16676,N_11764,N_14351);
and U16677 (N_16677,N_13658,N_12766);
nor U16678 (N_16678,N_13164,N_13463);
or U16679 (N_16679,N_12287,N_10866);
and U16680 (N_16680,N_13454,N_12608);
or U16681 (N_16681,N_11642,N_10827);
nand U16682 (N_16682,N_12971,N_11138);
xnor U16683 (N_16683,N_11153,N_10168);
xnor U16684 (N_16684,N_11759,N_12141);
xor U16685 (N_16685,N_10441,N_13719);
or U16686 (N_16686,N_13448,N_11868);
and U16687 (N_16687,N_11935,N_12243);
or U16688 (N_16688,N_11199,N_12326);
or U16689 (N_16689,N_10677,N_12823);
and U16690 (N_16690,N_11847,N_11067);
or U16691 (N_16691,N_14391,N_11322);
nand U16692 (N_16692,N_11089,N_14314);
nand U16693 (N_16693,N_13885,N_12700);
nand U16694 (N_16694,N_10326,N_12953);
and U16695 (N_16695,N_11304,N_10572);
nor U16696 (N_16696,N_12934,N_12321);
xor U16697 (N_16697,N_10002,N_13294);
nand U16698 (N_16698,N_12398,N_13199);
or U16699 (N_16699,N_10647,N_12577);
and U16700 (N_16700,N_14023,N_10418);
nand U16701 (N_16701,N_13834,N_10578);
and U16702 (N_16702,N_13179,N_10982);
nor U16703 (N_16703,N_13482,N_14927);
xor U16704 (N_16704,N_14575,N_11751);
and U16705 (N_16705,N_10498,N_12203);
xnor U16706 (N_16706,N_10380,N_12333);
xnor U16707 (N_16707,N_14473,N_13932);
or U16708 (N_16708,N_10068,N_13038);
or U16709 (N_16709,N_11399,N_14298);
xor U16710 (N_16710,N_12067,N_13011);
nor U16711 (N_16711,N_13081,N_13494);
xnor U16712 (N_16712,N_12555,N_12044);
xor U16713 (N_16713,N_13907,N_14758);
or U16714 (N_16714,N_10688,N_13329);
xnor U16715 (N_16715,N_14513,N_11421);
nor U16716 (N_16716,N_11051,N_10115);
nand U16717 (N_16717,N_14150,N_14385);
or U16718 (N_16718,N_11242,N_13274);
xnor U16719 (N_16719,N_12418,N_13025);
nor U16720 (N_16720,N_12324,N_12469);
xnor U16721 (N_16721,N_13136,N_14600);
or U16722 (N_16722,N_12459,N_13515);
nor U16723 (N_16723,N_11205,N_14606);
or U16724 (N_16724,N_14431,N_11830);
nand U16725 (N_16725,N_11496,N_12741);
nand U16726 (N_16726,N_10865,N_12581);
nor U16727 (N_16727,N_12584,N_12824);
nand U16728 (N_16728,N_13980,N_11882);
and U16729 (N_16729,N_12657,N_14207);
or U16730 (N_16730,N_14690,N_12834);
xor U16731 (N_16731,N_13022,N_13878);
and U16732 (N_16732,N_10894,N_14290);
and U16733 (N_16733,N_13369,N_11070);
xnor U16734 (N_16734,N_14535,N_14598);
nand U16735 (N_16735,N_14876,N_11091);
nor U16736 (N_16736,N_11389,N_10148);
xnor U16737 (N_16737,N_11701,N_14282);
nor U16738 (N_16738,N_14418,N_13423);
and U16739 (N_16739,N_12790,N_14367);
nand U16740 (N_16740,N_10466,N_11730);
xor U16741 (N_16741,N_10074,N_10969);
and U16742 (N_16742,N_10835,N_10356);
and U16743 (N_16743,N_12990,N_13652);
nor U16744 (N_16744,N_13270,N_12072);
or U16745 (N_16745,N_11520,N_14829);
nand U16746 (N_16746,N_13170,N_14065);
nand U16747 (N_16747,N_11119,N_13084);
and U16748 (N_16748,N_13736,N_13635);
or U16749 (N_16749,N_10172,N_13946);
nor U16750 (N_16750,N_12713,N_13149);
xnor U16751 (N_16751,N_14945,N_13429);
nand U16752 (N_16752,N_10862,N_12676);
or U16753 (N_16753,N_10728,N_14197);
nand U16754 (N_16754,N_13306,N_13722);
nor U16755 (N_16755,N_13930,N_13575);
and U16756 (N_16756,N_14224,N_12210);
or U16757 (N_16757,N_11177,N_12464);
nand U16758 (N_16758,N_12417,N_10195);
nand U16759 (N_16759,N_12332,N_12499);
or U16760 (N_16760,N_10712,N_12627);
and U16761 (N_16761,N_11218,N_13880);
nand U16762 (N_16762,N_11894,N_13299);
nor U16763 (N_16763,N_13596,N_13325);
and U16764 (N_16764,N_13083,N_10030);
xnor U16765 (N_16765,N_12848,N_14177);
or U16766 (N_16766,N_14607,N_12825);
nor U16767 (N_16767,N_13475,N_12535);
nor U16768 (N_16768,N_10547,N_10212);
and U16769 (N_16769,N_11225,N_13468);
xnor U16770 (N_16770,N_11548,N_14366);
xor U16771 (N_16771,N_10411,N_14103);
nor U16772 (N_16772,N_14732,N_13433);
nand U16773 (N_16773,N_10582,N_14243);
nor U16774 (N_16774,N_14072,N_11027);
xor U16775 (N_16775,N_10031,N_12960);
xor U16776 (N_16776,N_13420,N_10872);
xnor U16777 (N_16777,N_14898,N_11843);
nor U16778 (N_16778,N_11449,N_12025);
or U16779 (N_16779,N_13628,N_14830);
and U16780 (N_16780,N_13099,N_13746);
or U16781 (N_16781,N_10955,N_11643);
nor U16782 (N_16782,N_10004,N_12269);
and U16783 (N_16783,N_14614,N_10869);
and U16784 (N_16784,N_13682,N_12501);
and U16785 (N_16785,N_11708,N_13768);
and U16786 (N_16786,N_11521,N_14560);
xnor U16787 (N_16787,N_12860,N_11302);
nor U16788 (N_16788,N_11914,N_12776);
or U16789 (N_16789,N_14834,N_14544);
or U16790 (N_16790,N_11383,N_14377);
xnor U16791 (N_16791,N_11893,N_12309);
nand U16792 (N_16792,N_11021,N_14424);
nor U16793 (N_16793,N_13901,N_13811);
xor U16794 (N_16794,N_11108,N_11241);
nand U16795 (N_16795,N_11502,N_13771);
nand U16796 (N_16796,N_13997,N_13603);
xnor U16797 (N_16797,N_10710,N_10587);
or U16798 (N_16798,N_10238,N_13525);
or U16799 (N_16799,N_11415,N_10300);
or U16800 (N_16800,N_12702,N_10184);
and U16801 (N_16801,N_13049,N_10737);
or U16802 (N_16802,N_12294,N_14970);
nand U16803 (N_16803,N_12040,N_14157);
or U16804 (N_16804,N_12661,N_11875);
xor U16805 (N_16805,N_11804,N_12442);
or U16806 (N_16806,N_12832,N_12283);
xnor U16807 (N_16807,N_14481,N_11971);
nand U16808 (N_16808,N_13195,N_11943);
and U16809 (N_16809,N_12081,N_11684);
nand U16810 (N_16810,N_13678,N_11836);
or U16811 (N_16811,N_14057,N_10390);
nand U16812 (N_16812,N_11710,N_13256);
nand U16813 (N_16813,N_13012,N_10823);
or U16814 (N_16814,N_14727,N_14309);
nor U16815 (N_16815,N_12425,N_13892);
nand U16816 (N_16816,N_10505,N_10810);
xnor U16817 (N_16817,N_11980,N_12242);
nand U16818 (N_16818,N_11492,N_11016);
nor U16819 (N_16819,N_10939,N_14693);
nand U16820 (N_16820,N_10826,N_11586);
nor U16821 (N_16821,N_13863,N_13056);
and U16822 (N_16822,N_10259,N_12051);
nand U16823 (N_16823,N_14905,N_12086);
nand U16824 (N_16824,N_11560,N_12277);
xnor U16825 (N_16825,N_11172,N_14368);
nand U16826 (N_16826,N_10882,N_13917);
nand U16827 (N_16827,N_13110,N_10250);
nand U16828 (N_16828,N_14138,N_14706);
or U16829 (N_16829,N_12121,N_13339);
nor U16830 (N_16830,N_11886,N_11207);
or U16831 (N_16831,N_14392,N_12034);
xnor U16832 (N_16832,N_11858,N_12746);
nand U16833 (N_16833,N_10333,N_13851);
or U16834 (N_16834,N_14069,N_14479);
xor U16835 (N_16835,N_11149,N_13943);
and U16836 (N_16836,N_13095,N_10024);
xnor U16837 (N_16837,N_11771,N_14244);
nand U16838 (N_16838,N_14071,N_11600);
and U16839 (N_16839,N_12355,N_10127);
or U16840 (N_16840,N_13489,N_13017);
nand U16841 (N_16841,N_14524,N_13827);
or U16842 (N_16842,N_10265,N_14086);
nand U16843 (N_16843,N_10353,N_10694);
and U16844 (N_16844,N_14938,N_12313);
nor U16845 (N_16845,N_10732,N_11391);
nand U16846 (N_16846,N_10604,N_12048);
or U16847 (N_16847,N_10152,N_12237);
xor U16848 (N_16848,N_14108,N_10384);
xor U16849 (N_16849,N_12636,N_13814);
xnor U16850 (N_16850,N_13253,N_12764);
nand U16851 (N_16851,N_14806,N_10962);
nor U16852 (N_16852,N_13774,N_14229);
nor U16853 (N_16853,N_14421,N_11576);
and U16854 (N_16854,N_12671,N_14935);
and U16855 (N_16855,N_14238,N_12870);
or U16856 (N_16856,N_14734,N_10640);
xnor U16857 (N_16857,N_12773,N_11606);
or U16858 (N_16858,N_12917,N_10034);
nand U16859 (N_16859,N_11703,N_11162);
and U16860 (N_16860,N_10315,N_14082);
or U16861 (N_16861,N_10787,N_10278);
or U16862 (N_16862,N_14155,N_11879);
and U16863 (N_16863,N_14820,N_11920);
nor U16864 (N_16864,N_13418,N_12868);
or U16865 (N_16865,N_13568,N_10415);
and U16866 (N_16866,N_11940,N_13756);
nor U16867 (N_16867,N_10352,N_12329);
nor U16868 (N_16868,N_12236,N_13582);
nand U16869 (N_16869,N_13601,N_12991);
nor U16870 (N_16870,N_13745,N_12092);
or U16871 (N_16871,N_13787,N_14091);
and U16872 (N_16872,N_12267,N_12662);
nor U16873 (N_16873,N_10783,N_11709);
nand U16874 (N_16874,N_12234,N_12772);
xnor U16875 (N_16875,N_10359,N_12395);
nor U16876 (N_16876,N_13077,N_12087);
xor U16877 (N_16877,N_14505,N_12578);
or U16878 (N_16878,N_13229,N_12461);
and U16879 (N_16879,N_14790,N_11203);
or U16880 (N_16880,N_10860,N_10243);
and U16881 (N_16881,N_13184,N_10171);
nor U16882 (N_16882,N_14877,N_11698);
and U16883 (N_16883,N_13825,N_12192);
nand U16884 (N_16884,N_12477,N_12673);
and U16885 (N_16885,N_14725,N_10839);
nor U16886 (N_16886,N_10272,N_12039);
nor U16887 (N_16887,N_11232,N_11541);
xor U16888 (N_16888,N_10674,N_13695);
or U16889 (N_16889,N_14692,N_10774);
and U16890 (N_16890,N_13337,N_10200);
xnor U16891 (N_16891,N_14553,N_10733);
nor U16892 (N_16892,N_13236,N_10134);
or U16893 (N_16893,N_13701,N_11638);
and U16894 (N_16894,N_13654,N_10744);
nand U16895 (N_16895,N_12791,N_11788);
xnor U16896 (N_16896,N_11779,N_10740);
nand U16897 (N_16897,N_11682,N_14265);
nor U16898 (N_16898,N_11618,N_11491);
xnor U16899 (N_16899,N_12177,N_10759);
nor U16900 (N_16900,N_12538,N_14350);
nor U16901 (N_16901,N_14731,N_13824);
nor U16902 (N_16902,N_10691,N_11877);
and U16903 (N_16903,N_11612,N_14066);
and U16904 (N_16904,N_11427,N_10550);
or U16905 (N_16905,N_12471,N_12793);
and U16906 (N_16906,N_12718,N_12509);
nor U16907 (N_16907,N_14847,N_12997);
xor U16908 (N_16908,N_14044,N_13949);
nand U16909 (N_16909,N_11964,N_14570);
nand U16910 (N_16910,N_13589,N_11339);
nor U16911 (N_16911,N_11135,N_12010);
and U16912 (N_16912,N_10442,N_11065);
nand U16913 (N_16913,N_12804,N_12266);
and U16914 (N_16914,N_11271,N_12436);
nor U16915 (N_16915,N_10165,N_11419);
nor U16916 (N_16916,N_14654,N_11676);
nand U16917 (N_16917,N_10566,N_11303);
xnor U16918 (N_16918,N_13975,N_12225);
nand U16919 (N_16919,N_14121,N_14334);
nand U16920 (N_16920,N_14979,N_12828);
xnor U16921 (N_16921,N_11620,N_13323);
and U16922 (N_16922,N_13078,N_14456);
nand U16923 (N_16923,N_11565,N_11573);
xor U16924 (N_16924,N_11026,N_10392);
nor U16925 (N_16925,N_14504,N_14508);
nor U16926 (N_16926,N_12069,N_11489);
and U16927 (N_16927,N_14285,N_13784);
nand U16928 (N_16928,N_11433,N_13128);
xor U16929 (N_16929,N_12579,N_10554);
and U16930 (N_16930,N_14321,N_10474);
nor U16931 (N_16931,N_13633,N_12191);
or U16932 (N_16932,N_12050,N_10487);
nor U16933 (N_16933,N_10475,N_11228);
xor U16934 (N_16934,N_12779,N_11857);
nand U16935 (N_16935,N_10137,N_11833);
nor U16936 (N_16936,N_13148,N_11029);
xnor U16937 (N_16937,N_10494,N_10155);
nor U16938 (N_16938,N_11679,N_14842);
or U16939 (N_16939,N_12750,N_12803);
nor U16940 (N_16940,N_10108,N_10697);
nand U16941 (N_16941,N_12120,N_14556);
or U16942 (N_16942,N_11017,N_13043);
nand U16943 (N_16943,N_12602,N_11811);
nand U16944 (N_16944,N_10935,N_14682);
nor U16945 (N_16945,N_11034,N_14399);
nor U16946 (N_16946,N_14663,N_13300);
and U16947 (N_16947,N_13637,N_11948);
nor U16948 (N_16948,N_13660,N_12559);
or U16949 (N_16949,N_12957,N_10095);
and U16950 (N_16950,N_10575,N_10792);
nor U16951 (N_16951,N_12323,N_10997);
and U16952 (N_16952,N_13360,N_10201);
nand U16953 (N_16953,N_10056,N_10332);
and U16954 (N_16954,N_14907,N_11519);
nor U16955 (N_16955,N_11601,N_12916);
xnor U16956 (N_16956,N_13884,N_12070);
nor U16957 (N_16957,N_11330,N_10493);
xnor U16958 (N_16958,N_10124,N_14813);
xor U16959 (N_16959,N_12890,N_14262);
or U16960 (N_16960,N_10639,N_13304);
or U16961 (N_16961,N_10556,N_12261);
xnor U16962 (N_16962,N_14987,N_14850);
or U16963 (N_16963,N_11295,N_11532);
xor U16964 (N_16964,N_13072,N_12118);
nor U16965 (N_16965,N_11549,N_11328);
and U16966 (N_16966,N_14901,N_11594);
or U16967 (N_16967,N_13380,N_10459);
or U16968 (N_16968,N_14936,N_12734);
xnor U16969 (N_16969,N_14158,N_13252);
nor U16970 (N_16970,N_12349,N_11544);
nand U16971 (N_16971,N_11498,N_10094);
or U16972 (N_16972,N_10855,N_11774);
xor U16973 (N_16973,N_14379,N_11093);
xnor U16974 (N_16974,N_13626,N_14131);
xnor U16975 (N_16975,N_12230,N_14904);
or U16976 (N_16976,N_13872,N_13948);
nor U16977 (N_16977,N_13303,N_12373);
xor U16978 (N_16978,N_10966,N_13911);
and U16979 (N_16979,N_14593,N_12178);
or U16980 (N_16980,N_12877,N_14985);
nor U16981 (N_16981,N_13577,N_14514);
xnor U16982 (N_16982,N_11850,N_14323);
xor U16983 (N_16983,N_12819,N_12901);
xnor U16984 (N_16984,N_12797,N_11699);
or U16985 (N_16985,N_14947,N_10224);
and U16986 (N_16986,N_10138,N_10146);
or U16987 (N_16987,N_12603,N_14840);
or U16988 (N_16988,N_11347,N_12108);
xor U16989 (N_16989,N_13097,N_11321);
nor U16990 (N_16990,N_14989,N_11854);
nor U16991 (N_16991,N_13189,N_10452);
nand U16992 (N_16992,N_11945,N_10729);
nand U16993 (N_16993,N_12222,N_13645);
and U16994 (N_16994,N_12922,N_14548);
nand U16995 (N_16995,N_13926,N_11792);
or U16996 (N_16996,N_10558,N_13029);
nor U16997 (N_16997,N_10367,N_11098);
nor U16998 (N_16998,N_10623,N_12943);
nand U16999 (N_16999,N_11336,N_10830);
nand U17000 (N_17000,N_12365,N_11145);
and U17001 (N_17001,N_12839,N_13769);
nand U17002 (N_17002,N_13846,N_11342);
nand U17003 (N_17003,N_14317,N_13550);
and U17004 (N_17004,N_10061,N_13967);
and U17005 (N_17005,N_14170,N_11582);
nor U17006 (N_17006,N_13833,N_13549);
nand U17007 (N_17007,N_12369,N_10307);
nor U17008 (N_17008,N_12810,N_14037);
nand U17009 (N_17009,N_10946,N_10051);
and U17010 (N_17010,N_13711,N_13476);
xor U17011 (N_17011,N_11470,N_11602);
nand U17012 (N_17012,N_11742,N_10430);
nor U17013 (N_17013,N_13499,N_12595);
and U17014 (N_17014,N_14403,N_12367);
or U17015 (N_17015,N_12510,N_10461);
nand U17016 (N_17016,N_14181,N_11222);
and U17017 (N_17017,N_14745,N_11325);
nor U17018 (N_17018,N_11789,N_12162);
or U17019 (N_17019,N_11849,N_12556);
nor U17020 (N_17020,N_14417,N_13006);
nor U17021 (N_17021,N_10078,N_11862);
nand U17022 (N_17022,N_10173,N_12965);
and U17023 (N_17023,N_13706,N_12954);
or U17024 (N_17024,N_11622,N_11904);
and U17025 (N_17025,N_10393,N_12066);
xnor U17026 (N_17026,N_14264,N_12866);
xnor U17027 (N_17027,N_10701,N_12617);
nand U17028 (N_17028,N_11543,N_12962);
or U17029 (N_17029,N_10153,N_14467);
nor U17030 (N_17030,N_11842,N_10824);
nor U17031 (N_17031,N_14195,N_10012);
xnor U17032 (N_17032,N_13830,N_12198);
nand U17033 (N_17033,N_11744,N_10651);
xnor U17034 (N_17034,N_10263,N_13190);
nand U17035 (N_17035,N_11211,N_14228);
nor U17036 (N_17036,N_11039,N_13705);
and U17037 (N_17037,N_12980,N_10280);
nand U17038 (N_17038,N_12249,N_11035);
nand U17039 (N_17039,N_10305,N_10513);
and U17040 (N_17040,N_14045,N_11574);
and U17041 (N_17041,N_11169,N_13707);
nor U17042 (N_17042,N_12625,N_14836);
nand U17043 (N_17043,N_13757,N_11580);
xor U17044 (N_17044,N_11537,N_12851);
or U17045 (N_17045,N_12543,N_14757);
or U17046 (N_17046,N_12891,N_11147);
nand U17047 (N_17047,N_12835,N_12949);
nand U17048 (N_17048,N_14328,N_13221);
nand U17049 (N_17049,N_13509,N_10112);
nand U17050 (N_17050,N_10159,N_13446);
nor U17051 (N_17051,N_13493,N_10216);
and U17052 (N_17052,N_11686,N_10901);
nand U17053 (N_17053,N_13129,N_11460);
and U17054 (N_17054,N_10984,N_10213);
and U17055 (N_17055,N_11046,N_10038);
nand U17056 (N_17056,N_14920,N_11647);
nor U17057 (N_17057,N_12961,N_13093);
nor U17058 (N_17058,N_14763,N_12250);
xnor U17059 (N_17059,N_13273,N_10637);
nor U17060 (N_17060,N_11146,N_11324);
nor U17061 (N_17061,N_11451,N_12683);
nor U17062 (N_17062,N_13244,N_14632);
xor U17063 (N_17063,N_13246,N_12450);
or U17064 (N_17064,N_11856,N_11834);
or U17065 (N_17065,N_14831,N_10711);
and U17066 (N_17066,N_11430,N_10763);
xor U17067 (N_17067,N_14890,N_14017);
nand U17068 (N_17068,N_14441,N_11596);
and U17069 (N_17069,N_14049,N_12343);
xnor U17070 (N_17070,N_12553,N_10851);
nor U17071 (N_17071,N_10005,N_12410);
xor U17072 (N_17072,N_14895,N_14742);
or U17073 (N_17073,N_11000,N_10465);
or U17074 (N_17074,N_12928,N_14059);
nor U17075 (N_17075,N_10910,N_11352);
nor U17076 (N_17076,N_11221,N_13413);
and U17077 (N_17077,N_14287,N_10682);
and U17078 (N_17078,N_10672,N_13958);
or U17079 (N_17079,N_12857,N_14541);
or U17080 (N_17080,N_11803,N_13542);
nor U17081 (N_17081,N_14719,N_13233);
or U17082 (N_17082,N_11173,N_12958);
or U17083 (N_17083,N_14335,N_14859);
and U17084 (N_17084,N_13717,N_13543);
nor U17085 (N_17085,N_14175,N_12858);
nor U17086 (N_17086,N_11280,N_12792);
or U17087 (N_17087,N_13470,N_11335);
or U17088 (N_17088,N_10486,N_12523);
and U17089 (N_17089,N_12021,N_13562);
nor U17090 (N_17090,N_13497,N_10798);
xnor U17091 (N_17091,N_10436,N_14652);
xor U17092 (N_17092,N_13416,N_10736);
nor U17093 (N_17093,N_13172,N_12778);
xor U17094 (N_17094,N_11704,N_14503);
and U17095 (N_17095,N_13023,N_11165);
nand U17096 (N_17096,N_14478,N_10130);
nor U17097 (N_17097,N_14067,N_12228);
or U17098 (N_17098,N_10144,N_11705);
nor U17099 (N_17099,N_11248,N_14008);
nor U17100 (N_17100,N_11604,N_10249);
or U17101 (N_17101,N_14274,N_13671);
or U17102 (N_17102,N_12642,N_11898);
nand U17103 (N_17103,N_12923,N_11917);
and U17104 (N_17104,N_11130,N_14042);
and U17105 (N_17105,N_14817,N_13968);
nor U17106 (N_17106,N_12533,N_14958);
and U17107 (N_17107,N_14050,N_10413);
nand U17108 (N_17108,N_12195,N_10344);
nor U17109 (N_17109,N_11748,N_14799);
nand U17110 (N_17110,N_14261,N_10400);
or U17111 (N_17111,N_10756,N_10742);
or U17112 (N_17112,N_13368,N_10685);
or U17113 (N_17113,N_13714,N_14713);
or U17114 (N_17114,N_10199,N_12061);
nor U17115 (N_17115,N_11516,N_14089);
and U17116 (N_17116,N_12648,N_10363);
nor U17117 (N_17117,N_13683,N_11395);
nor U17118 (N_17118,N_13691,N_14981);
nor U17119 (N_17119,N_12330,N_13279);
nand U17120 (N_17120,N_12299,N_10035);
and U17121 (N_17121,N_10192,N_10066);
xnor U17122 (N_17122,N_12073,N_13609);
xnor U17123 (N_17123,N_14591,N_14319);
nand U17124 (N_17124,N_12641,N_10414);
and U17125 (N_17125,N_11959,N_14509);
or U17126 (N_17126,N_10179,N_14856);
and U17127 (N_17127,N_14577,N_13367);
or U17128 (N_17128,N_12731,N_10956);
xor U17129 (N_17129,N_13428,N_13868);
xnor U17130 (N_17130,N_11818,N_12244);
nor U17131 (N_17131,N_13557,N_14304);
or U17132 (N_17132,N_14507,N_11310);
or U17133 (N_17133,N_11760,N_11797);
nand U17134 (N_17134,N_14125,N_12382);
xor U17135 (N_17135,N_11458,N_13906);
and U17136 (N_17136,N_14695,N_10492);
xnor U17137 (N_17137,N_12977,N_10281);
or U17138 (N_17138,N_13343,N_12517);
nor U17139 (N_17139,N_11099,N_10952);
nor U17140 (N_17140,N_11090,N_11540);
or U17141 (N_17141,N_14436,N_10815);
nor U17142 (N_17142,N_14310,N_12312);
or U17143 (N_17143,N_12204,N_11985);
and U17144 (N_17144,N_13877,N_14307);
or U17145 (N_17145,N_11646,N_12017);
xnor U17146 (N_17146,N_10463,N_13555);
nand U17147 (N_17147,N_11915,N_11133);
xnor U17148 (N_17148,N_11685,N_10255);
xnor U17149 (N_17149,N_12551,N_12431);
and U17150 (N_17150,N_13064,N_11928);
or U17151 (N_17151,N_12013,N_12454);
nand U17152 (N_17152,N_12316,N_13226);
nor U17153 (N_17153,N_14174,N_10627);
and U17154 (N_17154,N_10500,N_11332);
or U17155 (N_17155,N_10501,N_13305);
and U17156 (N_17156,N_10859,N_13580);
nor U17157 (N_17157,N_11202,N_11049);
and U17158 (N_17158,N_14942,N_11912);
and U17159 (N_17159,N_12531,N_14634);
and U17160 (N_17160,N_12705,N_12457);
nand U17161 (N_17161,N_14053,N_13586);
and U17162 (N_17162,N_11184,N_14735);
nor U17163 (N_17163,N_13257,N_11161);
or U17164 (N_17164,N_14642,N_14762);
or U17165 (N_17165,N_12110,N_12377);
nor U17166 (N_17166,N_13382,N_14716);
and U17167 (N_17167,N_11137,N_14003);
or U17168 (N_17168,N_12357,N_13219);
nor U17169 (N_17169,N_11140,N_10749);
or U17170 (N_17170,N_12154,N_12720);
and U17171 (N_17171,N_11073,N_12413);
nand U17172 (N_17172,N_14268,N_14226);
nor U17173 (N_17173,N_12095,N_12566);
and U17174 (N_17174,N_11599,N_10203);
and U17175 (N_17175,N_12412,N_12285);
xor U17176 (N_17176,N_11436,N_10874);
xnor U17177 (N_17177,N_10338,N_10412);
and U17178 (N_17178,N_11473,N_14653);
or U17179 (N_17179,N_13625,N_11929);
nor U17180 (N_17180,N_11087,N_12435);
and U17181 (N_17181,N_11060,N_11536);
xnor U17182 (N_17182,N_14425,N_10490);
xor U17183 (N_17183,N_11168,N_11609);
xnor U17184 (N_17184,N_12947,N_14251);
nor U17185 (N_17185,N_12666,N_12239);
nor U17186 (N_17186,N_10355,N_10805);
nor U17187 (N_17187,N_12311,N_12484);
nor U17188 (N_17188,N_11208,N_13021);
or U17189 (N_17189,N_13812,N_13467);
and U17190 (N_17190,N_13986,N_13865);
nor U17191 (N_17191,N_11761,N_12619);
nand U17192 (N_17192,N_11696,N_11817);
nor U17193 (N_17193,N_13742,N_11590);
and U17194 (N_17194,N_12478,N_10844);
xnor U17195 (N_17195,N_11015,N_12889);
nor U17196 (N_17196,N_14483,N_11726);
xnor U17197 (N_17197,N_11871,N_14565);
nor U17198 (N_17198,N_14631,N_12688);
nor U17199 (N_17199,N_13261,N_14043);
and U17200 (N_17200,N_12004,N_11097);
nand U17201 (N_17201,N_13710,N_14389);
or U17202 (N_17202,N_11261,N_10661);
nor U17203 (N_17203,N_14145,N_12992);
xor U17204 (N_17204,N_10765,N_14486);
xor U17205 (N_17205,N_11859,N_11538);
or U17206 (N_17206,N_10133,N_13546);
or U17207 (N_17207,N_13800,N_14909);
xor U17208 (N_17208,N_13359,N_12123);
and U17209 (N_17209,N_10799,N_11036);
xnor U17210 (N_17210,N_11603,N_10879);
or U17211 (N_17211,N_14211,N_11897);
nand U17212 (N_17212,N_10423,N_14266);
nand U17213 (N_17213,N_13528,N_14573);
nor U17214 (N_17214,N_10111,N_12697);
nand U17215 (N_17215,N_10435,N_12088);
xnor U17216 (N_17216,N_13004,N_10785);
and U17217 (N_17217,N_14332,N_11068);
and U17218 (N_17218,N_11282,N_11477);
nor U17219 (N_17219,N_12647,N_14823);
xor U17220 (N_17220,N_10252,N_13876);
and U17221 (N_17221,N_11702,N_14419);
or U17222 (N_17222,N_11063,N_14645);
or U17223 (N_17223,N_11378,N_13090);
nand U17224 (N_17224,N_12897,N_10755);
xnor U17225 (N_17225,N_11354,N_10293);
or U17226 (N_17226,N_12609,N_12738);
and U17227 (N_17227,N_10867,N_12019);
nand U17228 (N_17228,N_10471,N_14246);
nor U17229 (N_17229,N_12580,N_11499);
nand U17230 (N_17230,N_12503,N_10634);
and U17231 (N_17231,N_14400,N_11076);
nor U17232 (N_17232,N_11823,N_14212);
nand U17233 (N_17233,N_14715,N_10788);
or U17234 (N_17234,N_12592,N_14218);
xor U17235 (N_17235,N_11486,N_11056);
or U17236 (N_17236,N_11973,N_11535);
nor U17237 (N_17237,N_11983,N_10981);
nand U17238 (N_17238,N_10276,N_13981);
nand U17239 (N_17239,N_10752,N_13716);
xnor U17240 (N_17240,N_10780,N_11043);
xnor U17241 (N_17241,N_14401,N_11522);
nand U17242 (N_17242,N_14388,N_10974);
nand U17243 (N_17243,N_14939,N_14192);
nand U17244 (N_17244,N_11995,N_10036);
or U17245 (N_17245,N_13408,N_10748);
and U17246 (N_17246,N_11819,N_14442);
nand U17247 (N_17247,N_10964,N_11770);
or U17248 (N_17248,N_13443,N_13160);
xnor U17249 (N_17249,N_10612,N_12983);
nand U17250 (N_17250,N_10614,N_10448);
xnor U17251 (N_17251,N_14674,N_11732);
nor U17252 (N_17252,N_11320,N_12742);
or U17253 (N_17253,N_14132,N_13139);
and U17254 (N_17254,N_14569,N_14487);
and U17255 (N_17255,N_13970,N_14187);
and U17256 (N_17256,N_14117,N_11795);
xnor U17257 (N_17257,N_11274,N_12494);
xnor U17258 (N_17258,N_13739,N_10121);
nor U17259 (N_17259,N_11160,N_12757);
or U17260 (N_17260,N_11297,N_12179);
or U17261 (N_17261,N_13014,N_14893);
and U17262 (N_17262,N_14623,N_10709);
nor U17263 (N_17263,N_12604,N_10923);
xnor U17264 (N_17264,N_14270,N_14176);
xor U17265 (N_17265,N_12387,N_11392);
nand U17266 (N_17266,N_11577,N_10198);
nand U17267 (N_17267,N_13898,N_13311);
nor U17268 (N_17268,N_14221,N_13794);
nand U17269 (N_17269,N_12106,N_10439);
xor U17270 (N_17270,N_13161,N_14722);
nor U17271 (N_17271,N_11019,N_14793);
xor U17272 (N_17272,N_11796,N_13944);
or U17273 (N_17273,N_10306,N_12893);
nand U17274 (N_17274,N_11787,N_13239);
and U17275 (N_17275,N_10526,N_12185);
nand U17276 (N_17276,N_14277,N_14342);
xnor U17277 (N_17277,N_13560,N_11997);
xnor U17278 (N_17278,N_13026,N_11665);
and U17279 (N_17279,N_11136,N_11798);
nand U17280 (N_17280,N_12518,N_12502);
and U17281 (N_17281,N_13541,N_12122);
nor U17282 (N_17282,N_12358,N_12827);
nand U17283 (N_17283,N_12785,N_11936);
nand U17284 (N_17284,N_11931,N_14750);
xnor U17285 (N_17285,N_14588,N_12390);
nor U17286 (N_17286,N_11131,N_10346);
nor U17287 (N_17287,N_10628,N_12655);
or U17288 (N_17288,N_11987,N_13168);
xnor U17289 (N_17289,N_14354,N_14411);
and U17290 (N_17290,N_10675,N_13961);
nor U17291 (N_17291,N_12850,N_11690);
nor U17292 (N_17292,N_13765,N_13570);
nor U17293 (N_17293,N_14025,N_14201);
and U17294 (N_17294,N_10470,N_12009);
or U17295 (N_17295,N_13207,N_11442);
or U17296 (N_17296,N_12801,N_12037);
xnor U17297 (N_17297,N_12621,N_11813);
and U17298 (N_17298,N_14446,N_14495);
or U17299 (N_17299,N_14405,N_12967);
and U17300 (N_17300,N_13798,N_13686);
nand U17301 (N_17301,N_11832,N_13676);
nor U17302 (N_17302,N_12375,N_10242);
nand U17303 (N_17303,N_14051,N_10845);
nand U17304 (N_17304,N_13277,N_14707);
or U17305 (N_17305,N_11672,N_10954);
xnor U17306 (N_17306,N_12907,N_10926);
or U17307 (N_17307,N_12840,N_11002);
or U17308 (N_17308,N_10820,N_13799);
or U17309 (N_17309,N_10636,N_11428);
xnor U17310 (N_17310,N_13852,N_11493);
xor U17311 (N_17311,N_13346,N_11820);
nor U17312 (N_17312,N_13890,N_14954);
nand U17313 (N_17313,N_13453,N_14559);
xnor U17314 (N_17314,N_14476,N_12289);
nand U17315 (N_17315,N_13922,N_11247);
nand U17316 (N_17316,N_14011,N_10629);
and U17317 (N_17317,N_11755,N_11013);
nor U17318 (N_17318,N_13118,N_14819);
nor U17319 (N_17319,N_11382,N_13657);
nand U17320 (N_17320,N_10150,N_11763);
and U17321 (N_17321,N_13789,N_14878);
nand U17322 (N_17322,N_12637,N_12942);
nor U17323 (N_17323,N_12388,N_12054);
xor U17324 (N_17324,N_10895,N_10456);
nand U17325 (N_17325,N_12574,N_12480);
and U17326 (N_17326,N_14058,N_13210);
xnor U17327 (N_17327,N_11125,N_10147);
and U17328 (N_17328,N_13449,N_13995);
or U17329 (N_17329,N_10158,N_12876);
nor U17330 (N_17330,N_11741,N_14397);
or U17331 (N_17331,N_11913,N_11490);
nor U17332 (N_17332,N_13109,N_14202);
nor U17333 (N_17333,N_12634,N_14636);
or U17334 (N_17334,N_12879,N_11353);
or U17335 (N_17335,N_11946,N_14944);
and U17336 (N_17336,N_12685,N_12747);
or U17337 (N_17337,N_11364,N_13498);
and U17338 (N_17338,N_14204,N_13301);
xor U17339 (N_17339,N_12841,N_14562);
nand U17340 (N_17340,N_11967,N_13508);
nor U17341 (N_17341,N_11591,N_13935);
and U17342 (N_17342,N_14609,N_11661);
or U17343 (N_17343,N_14055,N_13934);
nand U17344 (N_17344,N_10073,N_14612);
nand U17345 (N_17345,N_10467,N_10515);
or U17346 (N_17346,N_12206,N_12669);
and U17347 (N_17347,N_12711,N_12186);
nor U17348 (N_17348,N_12623,N_12771);
and U17349 (N_17349,N_10128,N_11343);
nand U17350 (N_17350,N_10191,N_12770);
nand U17351 (N_17351,N_14807,N_11079);
and U17352 (N_17352,N_11525,N_11716);
or U17353 (N_17353,N_14741,N_13854);
nor U17354 (N_17354,N_10398,N_13640);
or U17355 (N_17355,N_12811,N_10773);
nand U17356 (N_17356,N_10937,N_12226);
nand U17357 (N_17357,N_12842,N_11697);
and U17358 (N_17358,N_14773,N_14545);
and U17359 (N_17359,N_12620,N_12594);
nand U17360 (N_17360,N_11778,N_11844);
nand U17361 (N_17361,N_12371,N_13062);
or U17362 (N_17362,N_11393,N_11411);
and U17363 (N_17363,N_13677,N_11831);
nor U17364 (N_17364,N_10750,N_13116);
or U17365 (N_17365,N_11562,N_12346);
nand U17366 (N_17366,N_12252,N_13828);
or U17367 (N_17367,N_14027,N_14990);
and U17368 (N_17368,N_13989,N_13659);
nor U17369 (N_17369,N_13134,N_10190);
xor U17370 (N_17370,N_14971,N_11989);
and U17371 (N_17371,N_12190,N_12573);
nor U17372 (N_17372,N_12214,N_10339);
xnor U17373 (N_17373,N_12368,N_10723);
or U17374 (N_17374,N_12235,N_12002);
or U17375 (N_17375,N_14812,N_11245);
nor U17376 (N_17376,N_14148,N_12945);
xnor U17377 (N_17377,N_14450,N_14016);
nand U17378 (N_17378,N_11025,N_11754);
nand U17379 (N_17379,N_11892,N_10847);
nand U17380 (N_17380,N_12341,N_11581);
xor U17381 (N_17381,N_10699,N_13976);
nand U17382 (N_17382,N_13013,N_14353);
xor U17383 (N_17383,N_10312,N_13563);
xor U17384 (N_17384,N_11366,N_12886);
xor U17385 (N_17385,N_10589,N_13152);
and U17386 (N_17386,N_14752,N_12674);
nand U17387 (N_17387,N_10328,N_10343);
xnor U17388 (N_17388,N_11534,N_11623);
xor U17389 (N_17389,N_14863,N_10381);
nand U17390 (N_17390,N_12568,N_14292);
xnor U17391 (N_17391,N_12638,N_11524);
nor U17392 (N_17392,N_10468,N_14538);
and U17393 (N_17393,N_13972,N_12149);
and U17394 (N_17394,N_13032,N_13147);
and U17395 (N_17395,N_10963,N_14621);
nand U17396 (N_17396,N_11467,N_10040);
and U17397 (N_17397,N_13140,N_13842);
nor U17398 (N_17398,N_11578,N_10563);
nand U17399 (N_17399,N_11367,N_11841);
or U17400 (N_17400,N_13666,N_13767);
or U17401 (N_17401,N_14848,N_13405);
or U17402 (N_17402,N_11275,N_14033);
nor U17403 (N_17403,N_10245,N_10654);
and U17404 (N_17404,N_14728,N_14672);
nor U17405 (N_17405,N_11402,N_12297);
xnor U17406 (N_17406,N_11611,N_10590);
nand U17407 (N_17407,N_13648,N_11171);
and U17408 (N_17408,N_10704,N_11277);
and U17409 (N_17409,N_13150,N_10303);
nor U17410 (N_17410,N_10980,N_13196);
or U17411 (N_17411,N_11259,N_14068);
nand U17412 (N_17412,N_14416,N_12437);
or U17413 (N_17413,N_12701,N_11394);
nor U17414 (N_17414,N_11388,N_13527);
nor U17415 (N_17415,N_11633,N_13896);
xnor U17416 (N_17416,N_13073,N_14316);
nand U17417 (N_17417,N_12045,N_11619);
nand U17418 (N_17418,N_12350,N_10857);
xnor U17419 (N_17419,N_12440,N_14956);
nand U17420 (N_17420,N_14698,N_14488);
and U17421 (N_17421,N_12865,N_13455);
nor U17422 (N_17422,N_11624,N_12946);
xor U17423 (N_17423,N_14465,N_11375);
and U17424 (N_17424,N_11030,N_11300);
xnor U17425 (N_17425,N_12158,N_14376);
or U17426 (N_17426,N_13124,N_12089);
xor U17427 (N_17427,N_14341,N_10890);
xor U17428 (N_17428,N_10054,N_11791);
nor U17429 (N_17429,N_14753,N_13034);
xnor U17430 (N_17430,N_12974,N_10940);
and U17431 (N_17431,N_13381,N_11459);
and U17432 (N_17432,N_14818,N_11960);
or U17433 (N_17433,N_10813,N_12607);
nor U17434 (N_17434,N_11706,N_10945);
and U17435 (N_17435,N_12109,N_14021);
and U17436 (N_17436,N_13518,N_10145);
or U17437 (N_17437,N_12331,N_12929);
nand U17438 (N_17438,N_10644,N_14235);
xor U17439 (N_17439,N_10791,N_14163);
and U17440 (N_17440,N_14075,N_13243);
and U17441 (N_17441,N_11100,N_13537);
and U17442 (N_17442,N_11737,N_11246);
xnor U17443 (N_17443,N_12725,N_10613);
nor U17444 (N_17444,N_10136,N_14079);
nor U17445 (N_17445,N_13177,N_14554);
or U17446 (N_17446,N_12504,N_11220);
xor U17447 (N_17447,N_14547,N_13867);
nor U17448 (N_17448,N_11824,N_13447);
nand U17449 (N_17449,N_12151,N_12264);
or U17450 (N_17450,N_12855,N_13436);
xnor U17451 (N_17451,N_14493,N_11327);
nand U17452 (N_17452,N_12276,N_13672);
xor U17453 (N_17453,N_14528,N_11007);
nor U17454 (N_17454,N_12254,N_13786);
or U17455 (N_17455,N_13227,N_10555);
and U17456 (N_17456,N_11673,N_10282);
xor U17457 (N_17457,N_11982,N_13738);
or U17458 (N_17458,N_13451,N_14791);
nor U17459 (N_17459,N_12100,N_13108);
nor U17460 (N_17460,N_11235,N_10225);
nand U17461 (N_17461,N_11952,N_13713);
or U17462 (N_17462,N_14558,N_12020);
and U17463 (N_17463,N_11621,N_12137);
nor U17464 (N_17464,N_13530,N_10719);
nor U17465 (N_17465,N_14142,N_12384);
nand U17466 (N_17466,N_12229,N_11640);
xnor U17467 (N_17467,N_14182,N_10462);
and U17468 (N_17468,N_14798,N_10174);
and U17469 (N_17469,N_14772,N_10193);
nor U17470 (N_17470,N_11453,N_10961);
nor U17471 (N_17471,N_14782,N_11170);
or U17472 (N_17472,N_13624,N_10741);
xnor U17473 (N_17473,N_14700,N_13230);
xor U17474 (N_17474,N_12032,N_14511);
xnor U17475 (N_17475,N_13921,N_12762);
or U17476 (N_17476,N_11475,N_14888);
xor U17477 (N_17477,N_10531,N_14680);
or U17478 (N_17478,N_13398,N_13371);
xnor U17479 (N_17479,N_11900,N_11444);
xor U17480 (N_17480,N_12055,N_12873);
and U17481 (N_17481,N_14919,N_10236);
or U17482 (N_17482,N_10607,N_10904);
nor U17483 (N_17483,N_13692,N_14795);
or U17484 (N_17484,N_10804,N_14414);
or U17485 (N_17485,N_12196,N_10019);
nor U17486 (N_17486,N_14833,N_11563);
nor U17487 (N_17487,N_14589,N_12640);
and U17488 (N_17488,N_10816,N_11358);
nand U17489 (N_17489,N_10789,N_14081);
xnor U17490 (N_17490,N_13065,N_14912);
nand U17491 (N_17491,N_13320,N_10169);
xor U17492 (N_17492,N_10606,N_14206);
or U17493 (N_17493,N_10527,N_13668);
nand U17494 (N_17494,N_11306,N_14408);
nor U17495 (N_17495,N_14911,N_13037);
xnor U17496 (N_17496,N_13649,N_10545);
nand U17497 (N_17497,N_14002,N_11319);
xor U17498 (N_17498,N_11042,N_14372);
nor U17499 (N_17499,N_14064,N_11585);
nor U17500 (N_17500,N_14601,N_11983);
and U17501 (N_17501,N_13045,N_14628);
or U17502 (N_17502,N_13701,N_11874);
or U17503 (N_17503,N_12291,N_12659);
nor U17504 (N_17504,N_11863,N_12850);
nor U17505 (N_17505,N_14357,N_12877);
xor U17506 (N_17506,N_10260,N_10603);
nand U17507 (N_17507,N_12774,N_13373);
nor U17508 (N_17508,N_13822,N_12772);
xnor U17509 (N_17509,N_11532,N_10441);
nand U17510 (N_17510,N_11401,N_14926);
and U17511 (N_17511,N_11554,N_14903);
nor U17512 (N_17512,N_13630,N_10566);
nand U17513 (N_17513,N_12405,N_13177);
or U17514 (N_17514,N_10591,N_14597);
xor U17515 (N_17515,N_11128,N_10946);
or U17516 (N_17516,N_12170,N_11961);
nor U17517 (N_17517,N_10463,N_12608);
nand U17518 (N_17518,N_14181,N_14828);
nand U17519 (N_17519,N_12578,N_12088);
nand U17520 (N_17520,N_13223,N_13230);
nand U17521 (N_17521,N_14867,N_11771);
xor U17522 (N_17522,N_13978,N_12167);
or U17523 (N_17523,N_10408,N_13781);
or U17524 (N_17524,N_13465,N_10594);
or U17525 (N_17525,N_11099,N_12186);
xnor U17526 (N_17526,N_10184,N_11399);
nand U17527 (N_17527,N_13255,N_12959);
xnor U17528 (N_17528,N_10275,N_13033);
or U17529 (N_17529,N_11538,N_10966);
or U17530 (N_17530,N_10958,N_12302);
nand U17531 (N_17531,N_10798,N_10117);
or U17532 (N_17532,N_11248,N_11798);
or U17533 (N_17533,N_12781,N_14333);
nor U17534 (N_17534,N_11186,N_10138);
nand U17535 (N_17535,N_14918,N_10513);
nor U17536 (N_17536,N_11044,N_11209);
and U17537 (N_17537,N_14954,N_11673);
xnor U17538 (N_17538,N_11816,N_10320);
nor U17539 (N_17539,N_11898,N_14231);
and U17540 (N_17540,N_11447,N_12477);
nor U17541 (N_17541,N_14853,N_13545);
and U17542 (N_17542,N_12451,N_10928);
xor U17543 (N_17543,N_11973,N_10397);
nand U17544 (N_17544,N_10772,N_13795);
nor U17545 (N_17545,N_13479,N_11529);
or U17546 (N_17546,N_14140,N_10786);
xnor U17547 (N_17547,N_14006,N_10846);
or U17548 (N_17548,N_10517,N_14488);
and U17549 (N_17549,N_11775,N_11433);
xor U17550 (N_17550,N_12195,N_11965);
xnor U17551 (N_17551,N_10758,N_13080);
nor U17552 (N_17552,N_10196,N_13860);
xnor U17553 (N_17553,N_10452,N_13957);
nand U17554 (N_17554,N_10998,N_14523);
and U17555 (N_17555,N_12946,N_12521);
nand U17556 (N_17556,N_11696,N_12281);
xor U17557 (N_17557,N_12466,N_10744);
or U17558 (N_17558,N_12885,N_14340);
nor U17559 (N_17559,N_14217,N_12486);
or U17560 (N_17560,N_12878,N_13595);
nor U17561 (N_17561,N_13257,N_10877);
or U17562 (N_17562,N_14735,N_14681);
nand U17563 (N_17563,N_14286,N_11961);
xnor U17564 (N_17564,N_14586,N_10860);
and U17565 (N_17565,N_13011,N_13619);
xor U17566 (N_17566,N_12519,N_14917);
and U17567 (N_17567,N_11170,N_14810);
nor U17568 (N_17568,N_11311,N_11435);
and U17569 (N_17569,N_11016,N_13034);
or U17570 (N_17570,N_13860,N_13616);
or U17571 (N_17571,N_10648,N_13072);
nand U17572 (N_17572,N_12679,N_12851);
and U17573 (N_17573,N_13738,N_14392);
nand U17574 (N_17574,N_13531,N_11390);
nor U17575 (N_17575,N_13107,N_14886);
xnor U17576 (N_17576,N_10093,N_12869);
xnor U17577 (N_17577,N_14346,N_13966);
xor U17578 (N_17578,N_12991,N_12443);
xor U17579 (N_17579,N_12033,N_14550);
or U17580 (N_17580,N_12291,N_13074);
nor U17581 (N_17581,N_14044,N_14617);
and U17582 (N_17582,N_11931,N_10295);
and U17583 (N_17583,N_11834,N_13479);
nor U17584 (N_17584,N_12115,N_13588);
and U17585 (N_17585,N_12279,N_14158);
or U17586 (N_17586,N_14842,N_11031);
or U17587 (N_17587,N_13642,N_12246);
and U17588 (N_17588,N_13522,N_11886);
nor U17589 (N_17589,N_11665,N_12011);
nor U17590 (N_17590,N_11922,N_12157);
nor U17591 (N_17591,N_11205,N_10896);
nor U17592 (N_17592,N_14353,N_11427);
or U17593 (N_17593,N_13651,N_13406);
nor U17594 (N_17594,N_11184,N_10992);
xnor U17595 (N_17595,N_10499,N_13579);
nor U17596 (N_17596,N_12232,N_11259);
nand U17597 (N_17597,N_10350,N_13378);
xor U17598 (N_17598,N_14334,N_12571);
nand U17599 (N_17599,N_14538,N_10862);
nand U17600 (N_17600,N_13301,N_12877);
or U17601 (N_17601,N_10351,N_14399);
and U17602 (N_17602,N_10516,N_10716);
xor U17603 (N_17603,N_12220,N_11733);
nor U17604 (N_17604,N_14725,N_10918);
or U17605 (N_17605,N_11727,N_14156);
or U17606 (N_17606,N_11058,N_10520);
xor U17607 (N_17607,N_14291,N_11450);
xor U17608 (N_17608,N_14387,N_14704);
and U17609 (N_17609,N_14095,N_10428);
and U17610 (N_17610,N_12476,N_11284);
xor U17611 (N_17611,N_14524,N_13905);
nand U17612 (N_17612,N_14472,N_11472);
nand U17613 (N_17613,N_14890,N_10565);
xnor U17614 (N_17614,N_13410,N_13553);
nor U17615 (N_17615,N_11093,N_11946);
nand U17616 (N_17616,N_14597,N_10876);
nand U17617 (N_17617,N_14355,N_11132);
xor U17618 (N_17618,N_11028,N_13751);
or U17619 (N_17619,N_13162,N_12842);
xnor U17620 (N_17620,N_11060,N_11196);
and U17621 (N_17621,N_10053,N_11730);
xnor U17622 (N_17622,N_12323,N_14626);
and U17623 (N_17623,N_14149,N_11973);
nand U17624 (N_17624,N_11895,N_13605);
or U17625 (N_17625,N_11563,N_11319);
xor U17626 (N_17626,N_10211,N_12094);
nor U17627 (N_17627,N_10855,N_10698);
xor U17628 (N_17628,N_12286,N_12423);
and U17629 (N_17629,N_13988,N_13581);
nand U17630 (N_17630,N_14772,N_14890);
xor U17631 (N_17631,N_11737,N_11072);
nor U17632 (N_17632,N_13992,N_14462);
or U17633 (N_17633,N_11814,N_12365);
nand U17634 (N_17634,N_11405,N_14734);
and U17635 (N_17635,N_13480,N_14131);
and U17636 (N_17636,N_10211,N_13482);
xnor U17637 (N_17637,N_13813,N_10854);
nor U17638 (N_17638,N_12032,N_14217);
and U17639 (N_17639,N_12084,N_10985);
or U17640 (N_17640,N_11085,N_11340);
and U17641 (N_17641,N_10817,N_12995);
nor U17642 (N_17642,N_12148,N_14682);
xnor U17643 (N_17643,N_10785,N_12605);
xnor U17644 (N_17644,N_10038,N_11930);
or U17645 (N_17645,N_12279,N_12657);
or U17646 (N_17646,N_10311,N_12622);
nand U17647 (N_17647,N_13810,N_11136);
nor U17648 (N_17648,N_10618,N_10787);
and U17649 (N_17649,N_10611,N_11161);
and U17650 (N_17650,N_11695,N_12082);
nand U17651 (N_17651,N_11203,N_10567);
nor U17652 (N_17652,N_13895,N_13379);
xor U17653 (N_17653,N_12495,N_12278);
nand U17654 (N_17654,N_12297,N_10767);
or U17655 (N_17655,N_10788,N_13027);
or U17656 (N_17656,N_10706,N_12242);
nand U17657 (N_17657,N_14514,N_11800);
xnor U17658 (N_17658,N_10079,N_14003);
or U17659 (N_17659,N_12054,N_13669);
nor U17660 (N_17660,N_13782,N_13457);
xnor U17661 (N_17661,N_10809,N_12421);
and U17662 (N_17662,N_14737,N_13848);
and U17663 (N_17663,N_10148,N_11957);
xor U17664 (N_17664,N_13096,N_14348);
xnor U17665 (N_17665,N_13611,N_13899);
nand U17666 (N_17666,N_14415,N_12679);
nor U17667 (N_17667,N_11046,N_10725);
nor U17668 (N_17668,N_14455,N_12378);
xnor U17669 (N_17669,N_13721,N_14867);
and U17670 (N_17670,N_10881,N_10463);
xnor U17671 (N_17671,N_11966,N_10406);
or U17672 (N_17672,N_13501,N_11180);
nor U17673 (N_17673,N_11662,N_12688);
and U17674 (N_17674,N_11891,N_12757);
and U17675 (N_17675,N_12595,N_14476);
and U17676 (N_17676,N_11166,N_13511);
and U17677 (N_17677,N_14166,N_10009);
or U17678 (N_17678,N_12389,N_11219);
xor U17679 (N_17679,N_14505,N_12391);
or U17680 (N_17680,N_10438,N_14024);
nor U17681 (N_17681,N_13288,N_14724);
and U17682 (N_17682,N_13138,N_13056);
and U17683 (N_17683,N_11796,N_12748);
or U17684 (N_17684,N_11810,N_12008);
and U17685 (N_17685,N_13829,N_11690);
and U17686 (N_17686,N_10245,N_13741);
nor U17687 (N_17687,N_11872,N_10803);
nor U17688 (N_17688,N_13495,N_11021);
xor U17689 (N_17689,N_11825,N_12102);
and U17690 (N_17690,N_13492,N_12290);
nor U17691 (N_17691,N_11908,N_13313);
and U17692 (N_17692,N_11818,N_14634);
or U17693 (N_17693,N_14257,N_12943);
nor U17694 (N_17694,N_11934,N_10218);
xnor U17695 (N_17695,N_12136,N_11961);
or U17696 (N_17696,N_14324,N_11352);
nand U17697 (N_17697,N_11560,N_11838);
nand U17698 (N_17698,N_12322,N_14941);
xor U17699 (N_17699,N_10871,N_12451);
nand U17700 (N_17700,N_13279,N_10751);
nor U17701 (N_17701,N_10805,N_12820);
and U17702 (N_17702,N_14905,N_13511);
nand U17703 (N_17703,N_13303,N_11298);
xnor U17704 (N_17704,N_14439,N_12709);
nand U17705 (N_17705,N_10805,N_14020);
nor U17706 (N_17706,N_10025,N_10817);
or U17707 (N_17707,N_11731,N_11544);
xnor U17708 (N_17708,N_10466,N_12009);
xor U17709 (N_17709,N_13849,N_11017);
or U17710 (N_17710,N_10013,N_10186);
and U17711 (N_17711,N_13507,N_13960);
xor U17712 (N_17712,N_12296,N_11499);
and U17713 (N_17713,N_13359,N_14789);
or U17714 (N_17714,N_13204,N_12973);
nor U17715 (N_17715,N_14009,N_13332);
or U17716 (N_17716,N_10223,N_13002);
nor U17717 (N_17717,N_13479,N_14712);
nor U17718 (N_17718,N_12668,N_11581);
nor U17719 (N_17719,N_10799,N_10246);
nand U17720 (N_17720,N_11458,N_11354);
and U17721 (N_17721,N_14292,N_12960);
nand U17722 (N_17722,N_11123,N_11080);
nor U17723 (N_17723,N_11823,N_11845);
and U17724 (N_17724,N_13032,N_11186);
or U17725 (N_17725,N_11258,N_14846);
nand U17726 (N_17726,N_10375,N_13561);
or U17727 (N_17727,N_10725,N_12751);
nor U17728 (N_17728,N_11427,N_13356);
xor U17729 (N_17729,N_11553,N_10774);
nand U17730 (N_17730,N_11956,N_10297);
and U17731 (N_17731,N_12683,N_10721);
nand U17732 (N_17732,N_10890,N_14138);
nand U17733 (N_17733,N_11457,N_10157);
or U17734 (N_17734,N_11813,N_14818);
nand U17735 (N_17735,N_12396,N_10011);
nand U17736 (N_17736,N_13758,N_11367);
nand U17737 (N_17737,N_11801,N_12035);
nand U17738 (N_17738,N_10309,N_14325);
or U17739 (N_17739,N_13117,N_14562);
nand U17740 (N_17740,N_12891,N_13359);
or U17741 (N_17741,N_10617,N_10084);
nand U17742 (N_17742,N_11909,N_11659);
nand U17743 (N_17743,N_10104,N_14937);
and U17744 (N_17744,N_11151,N_13105);
and U17745 (N_17745,N_14824,N_12358);
nand U17746 (N_17746,N_10458,N_10500);
and U17747 (N_17747,N_10022,N_13758);
nand U17748 (N_17748,N_14477,N_10148);
nor U17749 (N_17749,N_10221,N_13245);
nand U17750 (N_17750,N_11973,N_12585);
and U17751 (N_17751,N_10371,N_14116);
nand U17752 (N_17752,N_12270,N_11831);
and U17753 (N_17753,N_13988,N_11256);
nand U17754 (N_17754,N_13975,N_13714);
and U17755 (N_17755,N_11288,N_12858);
and U17756 (N_17756,N_13645,N_12204);
nor U17757 (N_17757,N_12431,N_10843);
or U17758 (N_17758,N_12656,N_11338);
nand U17759 (N_17759,N_12270,N_12907);
xnor U17760 (N_17760,N_13591,N_11931);
nand U17761 (N_17761,N_13908,N_10242);
or U17762 (N_17762,N_11633,N_11607);
or U17763 (N_17763,N_12116,N_10815);
nor U17764 (N_17764,N_14736,N_10625);
xnor U17765 (N_17765,N_10728,N_12377);
and U17766 (N_17766,N_13445,N_10231);
nand U17767 (N_17767,N_12212,N_13796);
nand U17768 (N_17768,N_14063,N_11719);
nor U17769 (N_17769,N_14019,N_13334);
xor U17770 (N_17770,N_12440,N_10575);
xor U17771 (N_17771,N_12520,N_10310);
nor U17772 (N_17772,N_14340,N_14418);
nand U17773 (N_17773,N_13425,N_14160);
or U17774 (N_17774,N_13302,N_13132);
or U17775 (N_17775,N_14500,N_10358);
nand U17776 (N_17776,N_13997,N_10348);
xor U17777 (N_17777,N_11340,N_11912);
and U17778 (N_17778,N_14848,N_10673);
xnor U17779 (N_17779,N_12523,N_11328);
xnor U17780 (N_17780,N_14840,N_14570);
nand U17781 (N_17781,N_14495,N_13479);
nor U17782 (N_17782,N_12580,N_11752);
nand U17783 (N_17783,N_10483,N_10841);
xnor U17784 (N_17784,N_14145,N_10964);
xnor U17785 (N_17785,N_14651,N_11114);
xor U17786 (N_17786,N_13478,N_12697);
nand U17787 (N_17787,N_14561,N_10694);
xor U17788 (N_17788,N_14809,N_14768);
xor U17789 (N_17789,N_11289,N_13834);
or U17790 (N_17790,N_14092,N_13124);
xor U17791 (N_17791,N_11971,N_13459);
nor U17792 (N_17792,N_13688,N_10780);
and U17793 (N_17793,N_10811,N_13947);
nor U17794 (N_17794,N_10234,N_14757);
nand U17795 (N_17795,N_11742,N_14150);
xor U17796 (N_17796,N_12980,N_14441);
nand U17797 (N_17797,N_14684,N_12528);
xnor U17798 (N_17798,N_10222,N_12340);
nor U17799 (N_17799,N_14463,N_12893);
or U17800 (N_17800,N_13268,N_10580);
xnor U17801 (N_17801,N_11969,N_10167);
and U17802 (N_17802,N_14901,N_11596);
or U17803 (N_17803,N_11121,N_11918);
and U17804 (N_17804,N_14934,N_10618);
nor U17805 (N_17805,N_10759,N_12120);
nand U17806 (N_17806,N_11543,N_14667);
nor U17807 (N_17807,N_12065,N_14809);
nor U17808 (N_17808,N_11895,N_12836);
nand U17809 (N_17809,N_14571,N_10933);
and U17810 (N_17810,N_13797,N_13900);
or U17811 (N_17811,N_13987,N_14336);
and U17812 (N_17812,N_13365,N_10211);
or U17813 (N_17813,N_14754,N_13246);
nor U17814 (N_17814,N_13343,N_12950);
nand U17815 (N_17815,N_14892,N_12186);
nand U17816 (N_17816,N_10849,N_12826);
and U17817 (N_17817,N_13812,N_10138);
or U17818 (N_17818,N_11050,N_10754);
nor U17819 (N_17819,N_14083,N_14371);
xor U17820 (N_17820,N_10738,N_11513);
or U17821 (N_17821,N_14090,N_14582);
nor U17822 (N_17822,N_13707,N_11853);
and U17823 (N_17823,N_13976,N_14868);
and U17824 (N_17824,N_12153,N_11208);
nand U17825 (N_17825,N_14022,N_10923);
or U17826 (N_17826,N_12069,N_12099);
nand U17827 (N_17827,N_11845,N_11060);
nor U17828 (N_17828,N_10755,N_11484);
xor U17829 (N_17829,N_10013,N_10783);
and U17830 (N_17830,N_13626,N_11100);
or U17831 (N_17831,N_10896,N_12276);
or U17832 (N_17832,N_13124,N_12908);
and U17833 (N_17833,N_12866,N_10727);
nor U17834 (N_17834,N_11614,N_13832);
and U17835 (N_17835,N_12381,N_14512);
xor U17836 (N_17836,N_10389,N_14945);
nand U17837 (N_17837,N_11606,N_13079);
or U17838 (N_17838,N_10351,N_10289);
and U17839 (N_17839,N_14219,N_13409);
and U17840 (N_17840,N_13433,N_11200);
nand U17841 (N_17841,N_11641,N_13756);
nand U17842 (N_17842,N_12422,N_12857);
and U17843 (N_17843,N_13698,N_13738);
xnor U17844 (N_17844,N_12002,N_14740);
nor U17845 (N_17845,N_11531,N_10842);
xor U17846 (N_17846,N_12719,N_11400);
nor U17847 (N_17847,N_11153,N_14300);
nor U17848 (N_17848,N_11589,N_10242);
or U17849 (N_17849,N_14283,N_14030);
nor U17850 (N_17850,N_12329,N_13370);
xnor U17851 (N_17851,N_12389,N_13595);
or U17852 (N_17852,N_10803,N_14974);
nor U17853 (N_17853,N_13020,N_11239);
xnor U17854 (N_17854,N_10330,N_14848);
and U17855 (N_17855,N_12683,N_12196);
or U17856 (N_17856,N_12310,N_10280);
and U17857 (N_17857,N_10758,N_12542);
nor U17858 (N_17858,N_14147,N_11198);
nor U17859 (N_17859,N_10452,N_14186);
or U17860 (N_17860,N_13399,N_11960);
and U17861 (N_17861,N_13541,N_12996);
nor U17862 (N_17862,N_11087,N_14610);
nor U17863 (N_17863,N_14782,N_14480);
or U17864 (N_17864,N_11294,N_13781);
and U17865 (N_17865,N_13880,N_11967);
xor U17866 (N_17866,N_14092,N_10776);
nand U17867 (N_17867,N_14916,N_14181);
or U17868 (N_17868,N_13636,N_10519);
or U17869 (N_17869,N_14933,N_14212);
or U17870 (N_17870,N_13501,N_10918);
and U17871 (N_17871,N_11535,N_14145);
or U17872 (N_17872,N_12016,N_13086);
nand U17873 (N_17873,N_11858,N_14343);
nand U17874 (N_17874,N_10179,N_12854);
or U17875 (N_17875,N_11268,N_12000);
or U17876 (N_17876,N_10026,N_10851);
nor U17877 (N_17877,N_13316,N_12519);
xor U17878 (N_17878,N_14007,N_12299);
nand U17879 (N_17879,N_13130,N_12755);
or U17880 (N_17880,N_10740,N_10714);
or U17881 (N_17881,N_10221,N_12390);
and U17882 (N_17882,N_14125,N_11697);
or U17883 (N_17883,N_12849,N_14885);
xor U17884 (N_17884,N_11260,N_13300);
or U17885 (N_17885,N_11660,N_14393);
or U17886 (N_17886,N_13875,N_13418);
nand U17887 (N_17887,N_12749,N_11429);
nor U17888 (N_17888,N_12281,N_12833);
xnor U17889 (N_17889,N_11807,N_11666);
or U17890 (N_17890,N_11192,N_10356);
nor U17891 (N_17891,N_13712,N_14331);
nand U17892 (N_17892,N_10168,N_13452);
or U17893 (N_17893,N_11133,N_11737);
nor U17894 (N_17894,N_14807,N_11511);
or U17895 (N_17895,N_14703,N_10788);
nand U17896 (N_17896,N_14821,N_14890);
or U17897 (N_17897,N_13450,N_13627);
or U17898 (N_17898,N_12988,N_14815);
nor U17899 (N_17899,N_14004,N_12578);
and U17900 (N_17900,N_10087,N_13718);
or U17901 (N_17901,N_13296,N_10532);
nor U17902 (N_17902,N_12633,N_11541);
xnor U17903 (N_17903,N_12237,N_13801);
nand U17904 (N_17904,N_10582,N_13953);
xor U17905 (N_17905,N_10610,N_10222);
nand U17906 (N_17906,N_11472,N_13760);
nand U17907 (N_17907,N_13106,N_10759);
nor U17908 (N_17908,N_13761,N_12789);
xnor U17909 (N_17909,N_14426,N_10335);
nor U17910 (N_17910,N_10521,N_11213);
nor U17911 (N_17911,N_11818,N_13644);
or U17912 (N_17912,N_10463,N_12610);
xor U17913 (N_17913,N_14393,N_14445);
or U17914 (N_17914,N_14856,N_10012);
nand U17915 (N_17915,N_12761,N_11030);
xor U17916 (N_17916,N_11554,N_11020);
nand U17917 (N_17917,N_14725,N_13631);
nor U17918 (N_17918,N_11196,N_13266);
and U17919 (N_17919,N_12056,N_13718);
nand U17920 (N_17920,N_13720,N_11375);
nor U17921 (N_17921,N_11016,N_14764);
or U17922 (N_17922,N_10758,N_12218);
xor U17923 (N_17923,N_10493,N_11482);
xor U17924 (N_17924,N_10957,N_11442);
and U17925 (N_17925,N_10588,N_14260);
and U17926 (N_17926,N_10046,N_10724);
and U17927 (N_17927,N_10206,N_13207);
nand U17928 (N_17928,N_14564,N_10470);
xnor U17929 (N_17929,N_13332,N_13495);
nor U17930 (N_17930,N_10478,N_13528);
nor U17931 (N_17931,N_10650,N_13970);
nor U17932 (N_17932,N_13733,N_11613);
xnor U17933 (N_17933,N_13212,N_13229);
nor U17934 (N_17934,N_11277,N_13437);
or U17935 (N_17935,N_14033,N_13797);
or U17936 (N_17936,N_11829,N_13763);
and U17937 (N_17937,N_12686,N_11806);
or U17938 (N_17938,N_14174,N_11256);
nor U17939 (N_17939,N_13834,N_11500);
or U17940 (N_17940,N_13672,N_13006);
and U17941 (N_17941,N_13374,N_10368);
nand U17942 (N_17942,N_10091,N_14479);
nor U17943 (N_17943,N_13923,N_12501);
and U17944 (N_17944,N_12778,N_12293);
nand U17945 (N_17945,N_14521,N_10771);
and U17946 (N_17946,N_11932,N_12501);
or U17947 (N_17947,N_13576,N_13848);
nor U17948 (N_17948,N_10550,N_13059);
nor U17949 (N_17949,N_14553,N_14269);
nor U17950 (N_17950,N_11465,N_13069);
or U17951 (N_17951,N_12658,N_13427);
nor U17952 (N_17952,N_11642,N_12354);
and U17953 (N_17953,N_14796,N_12115);
xnor U17954 (N_17954,N_13613,N_10332);
nand U17955 (N_17955,N_12083,N_12262);
nor U17956 (N_17956,N_11908,N_11674);
nor U17957 (N_17957,N_14870,N_14254);
and U17958 (N_17958,N_14093,N_10486);
or U17959 (N_17959,N_11131,N_13309);
xor U17960 (N_17960,N_11862,N_12322);
and U17961 (N_17961,N_10366,N_14345);
nand U17962 (N_17962,N_13746,N_12625);
xnor U17963 (N_17963,N_10952,N_13877);
nand U17964 (N_17964,N_14054,N_13701);
nor U17965 (N_17965,N_13170,N_11544);
and U17966 (N_17966,N_11582,N_13365);
and U17967 (N_17967,N_12331,N_12313);
nand U17968 (N_17968,N_10615,N_10766);
or U17969 (N_17969,N_13694,N_12198);
or U17970 (N_17970,N_11234,N_13011);
nand U17971 (N_17971,N_12087,N_10741);
or U17972 (N_17972,N_13594,N_13200);
nand U17973 (N_17973,N_14719,N_11529);
or U17974 (N_17974,N_13843,N_12958);
nor U17975 (N_17975,N_10667,N_13625);
or U17976 (N_17976,N_13615,N_13256);
nor U17977 (N_17977,N_10267,N_12109);
and U17978 (N_17978,N_11233,N_13129);
nand U17979 (N_17979,N_12035,N_12636);
nor U17980 (N_17980,N_14513,N_14289);
and U17981 (N_17981,N_12175,N_13563);
or U17982 (N_17982,N_12593,N_13328);
and U17983 (N_17983,N_14580,N_14283);
and U17984 (N_17984,N_10269,N_13317);
or U17985 (N_17985,N_11452,N_10953);
or U17986 (N_17986,N_12531,N_11693);
nor U17987 (N_17987,N_13184,N_11813);
nor U17988 (N_17988,N_10079,N_11503);
or U17989 (N_17989,N_11527,N_14015);
nand U17990 (N_17990,N_10116,N_11486);
or U17991 (N_17991,N_13633,N_13013);
or U17992 (N_17992,N_10858,N_14619);
or U17993 (N_17993,N_12146,N_12736);
and U17994 (N_17994,N_13766,N_10022);
and U17995 (N_17995,N_14608,N_13820);
and U17996 (N_17996,N_10808,N_11025);
or U17997 (N_17997,N_13821,N_13759);
or U17998 (N_17998,N_11464,N_14635);
and U17999 (N_17999,N_14747,N_11642);
nor U18000 (N_18000,N_10764,N_11058);
and U18001 (N_18001,N_10421,N_13947);
or U18002 (N_18002,N_13548,N_13963);
or U18003 (N_18003,N_14028,N_11004);
nor U18004 (N_18004,N_14324,N_12496);
xor U18005 (N_18005,N_11327,N_13523);
nor U18006 (N_18006,N_11576,N_13014);
xnor U18007 (N_18007,N_12895,N_10484);
nand U18008 (N_18008,N_14987,N_10820);
nor U18009 (N_18009,N_11280,N_10999);
xor U18010 (N_18010,N_11690,N_10707);
and U18011 (N_18011,N_14198,N_11301);
and U18012 (N_18012,N_14615,N_14340);
nor U18013 (N_18013,N_12052,N_14515);
nand U18014 (N_18014,N_13022,N_14995);
nor U18015 (N_18015,N_10410,N_14359);
xor U18016 (N_18016,N_14583,N_13791);
nand U18017 (N_18017,N_14857,N_11343);
or U18018 (N_18018,N_13472,N_12001);
or U18019 (N_18019,N_11135,N_10678);
nand U18020 (N_18020,N_12902,N_13781);
nor U18021 (N_18021,N_14541,N_14568);
or U18022 (N_18022,N_10400,N_14791);
and U18023 (N_18023,N_13259,N_10173);
or U18024 (N_18024,N_14499,N_10908);
xnor U18025 (N_18025,N_10727,N_11847);
xor U18026 (N_18026,N_11808,N_10121);
or U18027 (N_18027,N_11363,N_11584);
xnor U18028 (N_18028,N_13186,N_12118);
nor U18029 (N_18029,N_13693,N_10709);
or U18030 (N_18030,N_12332,N_11879);
xor U18031 (N_18031,N_12964,N_11068);
or U18032 (N_18032,N_12675,N_11534);
nor U18033 (N_18033,N_11696,N_12019);
xnor U18034 (N_18034,N_11159,N_10245);
nor U18035 (N_18035,N_11372,N_14902);
or U18036 (N_18036,N_11503,N_12567);
and U18037 (N_18037,N_10292,N_11835);
or U18038 (N_18038,N_14868,N_11419);
nand U18039 (N_18039,N_14826,N_11147);
xor U18040 (N_18040,N_13171,N_14434);
or U18041 (N_18041,N_14817,N_14689);
or U18042 (N_18042,N_10170,N_13080);
nor U18043 (N_18043,N_13133,N_13201);
nor U18044 (N_18044,N_12825,N_14612);
xor U18045 (N_18045,N_11091,N_13347);
or U18046 (N_18046,N_13520,N_14032);
and U18047 (N_18047,N_10594,N_14161);
or U18048 (N_18048,N_11857,N_14270);
xor U18049 (N_18049,N_14651,N_12457);
xnor U18050 (N_18050,N_11508,N_14811);
xor U18051 (N_18051,N_12040,N_12449);
and U18052 (N_18052,N_12851,N_10369);
and U18053 (N_18053,N_12676,N_10429);
or U18054 (N_18054,N_11481,N_12744);
xor U18055 (N_18055,N_10747,N_11024);
xnor U18056 (N_18056,N_14910,N_10360);
nor U18057 (N_18057,N_14407,N_13585);
xnor U18058 (N_18058,N_11126,N_14912);
nand U18059 (N_18059,N_13592,N_11173);
nand U18060 (N_18060,N_11349,N_11916);
nor U18061 (N_18061,N_13561,N_13558);
nor U18062 (N_18062,N_14672,N_12833);
nand U18063 (N_18063,N_13651,N_11920);
xnor U18064 (N_18064,N_12781,N_10592);
nor U18065 (N_18065,N_13386,N_13754);
xor U18066 (N_18066,N_13134,N_12361);
and U18067 (N_18067,N_10970,N_10279);
xor U18068 (N_18068,N_13156,N_12630);
and U18069 (N_18069,N_10429,N_14516);
and U18070 (N_18070,N_11238,N_10664);
or U18071 (N_18071,N_11413,N_12354);
nor U18072 (N_18072,N_14306,N_14567);
nand U18073 (N_18073,N_10174,N_12777);
nand U18074 (N_18074,N_12525,N_11959);
and U18075 (N_18075,N_13599,N_10145);
and U18076 (N_18076,N_14418,N_10111);
nor U18077 (N_18077,N_10771,N_12653);
nor U18078 (N_18078,N_10215,N_14517);
nand U18079 (N_18079,N_11612,N_14732);
nor U18080 (N_18080,N_10730,N_12623);
or U18081 (N_18081,N_14405,N_10573);
nor U18082 (N_18082,N_10993,N_11308);
or U18083 (N_18083,N_14100,N_11584);
nor U18084 (N_18084,N_13618,N_11692);
and U18085 (N_18085,N_11519,N_12158);
nand U18086 (N_18086,N_11920,N_14956);
nand U18087 (N_18087,N_14182,N_14050);
nand U18088 (N_18088,N_10211,N_13400);
and U18089 (N_18089,N_13718,N_11710);
xor U18090 (N_18090,N_10418,N_12278);
and U18091 (N_18091,N_13706,N_12472);
nor U18092 (N_18092,N_13636,N_13227);
xnor U18093 (N_18093,N_10688,N_12216);
nor U18094 (N_18094,N_12611,N_11894);
nand U18095 (N_18095,N_14375,N_12723);
nand U18096 (N_18096,N_14672,N_13133);
xor U18097 (N_18097,N_11854,N_10844);
nand U18098 (N_18098,N_11612,N_13880);
or U18099 (N_18099,N_14069,N_14693);
nand U18100 (N_18100,N_11739,N_13326);
and U18101 (N_18101,N_13455,N_12159);
nand U18102 (N_18102,N_12171,N_10508);
and U18103 (N_18103,N_14029,N_10015);
nor U18104 (N_18104,N_14777,N_12750);
and U18105 (N_18105,N_11248,N_13482);
and U18106 (N_18106,N_11808,N_12146);
nand U18107 (N_18107,N_11467,N_14785);
nand U18108 (N_18108,N_14043,N_14437);
xor U18109 (N_18109,N_12570,N_13561);
nor U18110 (N_18110,N_10623,N_10486);
nand U18111 (N_18111,N_14362,N_12324);
nand U18112 (N_18112,N_10288,N_11010);
or U18113 (N_18113,N_11155,N_13738);
or U18114 (N_18114,N_10729,N_13467);
or U18115 (N_18115,N_11792,N_14912);
nand U18116 (N_18116,N_13912,N_12946);
and U18117 (N_18117,N_12090,N_11526);
or U18118 (N_18118,N_10269,N_13553);
nor U18119 (N_18119,N_13893,N_12347);
or U18120 (N_18120,N_12534,N_12949);
nand U18121 (N_18121,N_12628,N_12806);
nand U18122 (N_18122,N_13315,N_10611);
xor U18123 (N_18123,N_14455,N_14439);
nand U18124 (N_18124,N_13984,N_12861);
nor U18125 (N_18125,N_12196,N_14333);
and U18126 (N_18126,N_11956,N_10163);
or U18127 (N_18127,N_12036,N_11340);
nand U18128 (N_18128,N_14967,N_14073);
and U18129 (N_18129,N_11043,N_13770);
nor U18130 (N_18130,N_13356,N_12009);
and U18131 (N_18131,N_11507,N_11986);
xor U18132 (N_18132,N_12388,N_10862);
nor U18133 (N_18133,N_10158,N_11694);
nor U18134 (N_18134,N_12360,N_12146);
and U18135 (N_18135,N_12711,N_10069);
or U18136 (N_18136,N_13434,N_13755);
xor U18137 (N_18137,N_10790,N_14296);
nand U18138 (N_18138,N_10861,N_11971);
nand U18139 (N_18139,N_12592,N_11831);
xor U18140 (N_18140,N_12558,N_14183);
or U18141 (N_18141,N_13755,N_14621);
xor U18142 (N_18142,N_12589,N_10784);
or U18143 (N_18143,N_13783,N_11691);
xor U18144 (N_18144,N_10391,N_11565);
xor U18145 (N_18145,N_10652,N_10982);
nor U18146 (N_18146,N_10150,N_13099);
nand U18147 (N_18147,N_13594,N_10093);
or U18148 (N_18148,N_13083,N_14765);
and U18149 (N_18149,N_13837,N_14054);
nor U18150 (N_18150,N_12003,N_14977);
nor U18151 (N_18151,N_10922,N_12549);
or U18152 (N_18152,N_12478,N_13792);
nand U18153 (N_18153,N_11679,N_14553);
nand U18154 (N_18154,N_13353,N_10150);
or U18155 (N_18155,N_10841,N_12371);
xnor U18156 (N_18156,N_12941,N_13400);
nand U18157 (N_18157,N_13154,N_10929);
nand U18158 (N_18158,N_14084,N_11720);
nand U18159 (N_18159,N_10082,N_12827);
xor U18160 (N_18160,N_14251,N_11034);
or U18161 (N_18161,N_12279,N_13653);
nor U18162 (N_18162,N_12072,N_12551);
xor U18163 (N_18163,N_11996,N_11162);
and U18164 (N_18164,N_12697,N_12818);
nor U18165 (N_18165,N_10315,N_13302);
nand U18166 (N_18166,N_13420,N_12421);
xnor U18167 (N_18167,N_13754,N_10547);
nor U18168 (N_18168,N_10159,N_10446);
or U18169 (N_18169,N_12673,N_14993);
and U18170 (N_18170,N_12556,N_12687);
or U18171 (N_18171,N_10227,N_11009);
xnor U18172 (N_18172,N_14324,N_14022);
xnor U18173 (N_18173,N_12309,N_14322);
and U18174 (N_18174,N_11673,N_12648);
or U18175 (N_18175,N_11239,N_13079);
or U18176 (N_18176,N_12999,N_11422);
or U18177 (N_18177,N_11400,N_12087);
nor U18178 (N_18178,N_11509,N_13283);
and U18179 (N_18179,N_11017,N_13841);
or U18180 (N_18180,N_10591,N_14426);
nor U18181 (N_18181,N_12987,N_14763);
nand U18182 (N_18182,N_11489,N_11275);
nor U18183 (N_18183,N_10838,N_14037);
or U18184 (N_18184,N_12655,N_10265);
nand U18185 (N_18185,N_11682,N_13624);
xor U18186 (N_18186,N_12007,N_11481);
or U18187 (N_18187,N_14576,N_11352);
and U18188 (N_18188,N_13669,N_12464);
or U18189 (N_18189,N_12440,N_11235);
nor U18190 (N_18190,N_11122,N_14352);
nand U18191 (N_18191,N_12478,N_11776);
xnor U18192 (N_18192,N_13223,N_10364);
and U18193 (N_18193,N_14854,N_14640);
or U18194 (N_18194,N_11759,N_10700);
xnor U18195 (N_18195,N_12894,N_11289);
and U18196 (N_18196,N_10122,N_11118);
nand U18197 (N_18197,N_12298,N_12608);
and U18198 (N_18198,N_13731,N_12331);
or U18199 (N_18199,N_11003,N_13829);
or U18200 (N_18200,N_12376,N_13915);
xor U18201 (N_18201,N_11149,N_14669);
or U18202 (N_18202,N_12315,N_14913);
and U18203 (N_18203,N_12106,N_13698);
nor U18204 (N_18204,N_13783,N_12660);
nor U18205 (N_18205,N_13316,N_14400);
nor U18206 (N_18206,N_11844,N_11245);
and U18207 (N_18207,N_13615,N_10509);
nand U18208 (N_18208,N_12811,N_11076);
or U18209 (N_18209,N_10356,N_14512);
nand U18210 (N_18210,N_14622,N_10439);
or U18211 (N_18211,N_12599,N_10596);
nor U18212 (N_18212,N_11433,N_10342);
or U18213 (N_18213,N_12463,N_14669);
xnor U18214 (N_18214,N_11611,N_10262);
and U18215 (N_18215,N_14858,N_10797);
or U18216 (N_18216,N_10072,N_12606);
nor U18217 (N_18217,N_14579,N_13587);
xnor U18218 (N_18218,N_13699,N_12041);
nor U18219 (N_18219,N_12401,N_12859);
or U18220 (N_18220,N_12935,N_14461);
nand U18221 (N_18221,N_14735,N_13338);
xnor U18222 (N_18222,N_13111,N_14638);
or U18223 (N_18223,N_10241,N_10343);
or U18224 (N_18224,N_12121,N_10380);
xnor U18225 (N_18225,N_11622,N_13405);
nand U18226 (N_18226,N_10147,N_13603);
nor U18227 (N_18227,N_10031,N_11248);
nor U18228 (N_18228,N_10658,N_14915);
nor U18229 (N_18229,N_13450,N_11628);
or U18230 (N_18230,N_13206,N_14842);
nand U18231 (N_18231,N_11539,N_10934);
and U18232 (N_18232,N_14347,N_11118);
xor U18233 (N_18233,N_11357,N_11094);
xor U18234 (N_18234,N_12983,N_11758);
nor U18235 (N_18235,N_12445,N_12079);
and U18236 (N_18236,N_14061,N_10632);
or U18237 (N_18237,N_14941,N_11470);
and U18238 (N_18238,N_12304,N_13108);
nor U18239 (N_18239,N_10397,N_13756);
nand U18240 (N_18240,N_13642,N_11013);
xnor U18241 (N_18241,N_11619,N_11246);
or U18242 (N_18242,N_12809,N_14096);
xnor U18243 (N_18243,N_12130,N_11563);
nand U18244 (N_18244,N_11979,N_12316);
or U18245 (N_18245,N_10230,N_12422);
and U18246 (N_18246,N_11670,N_13401);
xor U18247 (N_18247,N_14795,N_12293);
and U18248 (N_18248,N_14764,N_10004);
or U18249 (N_18249,N_10072,N_10159);
and U18250 (N_18250,N_11840,N_12977);
nand U18251 (N_18251,N_14316,N_11453);
xnor U18252 (N_18252,N_13473,N_13700);
or U18253 (N_18253,N_13409,N_10542);
nor U18254 (N_18254,N_12720,N_12906);
nand U18255 (N_18255,N_11467,N_10881);
or U18256 (N_18256,N_12947,N_14577);
nand U18257 (N_18257,N_10861,N_11065);
nor U18258 (N_18258,N_13484,N_11877);
or U18259 (N_18259,N_13048,N_11216);
nand U18260 (N_18260,N_11386,N_11180);
or U18261 (N_18261,N_12214,N_13515);
nor U18262 (N_18262,N_13307,N_13398);
xnor U18263 (N_18263,N_14570,N_13123);
xor U18264 (N_18264,N_14275,N_14882);
nor U18265 (N_18265,N_12368,N_13584);
and U18266 (N_18266,N_10368,N_10575);
xor U18267 (N_18267,N_11606,N_12641);
and U18268 (N_18268,N_12616,N_14904);
or U18269 (N_18269,N_14648,N_13935);
and U18270 (N_18270,N_10083,N_13203);
nor U18271 (N_18271,N_13360,N_10901);
nand U18272 (N_18272,N_14016,N_13515);
and U18273 (N_18273,N_14647,N_10948);
or U18274 (N_18274,N_11770,N_12022);
and U18275 (N_18275,N_10274,N_13579);
xnor U18276 (N_18276,N_13751,N_12871);
or U18277 (N_18277,N_12974,N_14642);
nor U18278 (N_18278,N_14408,N_11416);
nor U18279 (N_18279,N_11909,N_12462);
nand U18280 (N_18280,N_13162,N_14891);
nor U18281 (N_18281,N_11387,N_13540);
xor U18282 (N_18282,N_14409,N_12193);
and U18283 (N_18283,N_10766,N_12823);
and U18284 (N_18284,N_12490,N_14820);
nand U18285 (N_18285,N_13124,N_10374);
or U18286 (N_18286,N_13438,N_14295);
xnor U18287 (N_18287,N_12931,N_12634);
xor U18288 (N_18288,N_10035,N_14441);
nand U18289 (N_18289,N_11481,N_11304);
nand U18290 (N_18290,N_14186,N_11433);
or U18291 (N_18291,N_14508,N_13132);
or U18292 (N_18292,N_10514,N_13022);
and U18293 (N_18293,N_11906,N_12274);
and U18294 (N_18294,N_14725,N_11395);
xnor U18295 (N_18295,N_12944,N_11228);
nand U18296 (N_18296,N_10218,N_14275);
or U18297 (N_18297,N_11534,N_14987);
xnor U18298 (N_18298,N_11147,N_14353);
nand U18299 (N_18299,N_14852,N_11795);
xor U18300 (N_18300,N_11578,N_12979);
xnor U18301 (N_18301,N_14522,N_12837);
or U18302 (N_18302,N_13443,N_12457);
nor U18303 (N_18303,N_10245,N_11836);
xor U18304 (N_18304,N_13199,N_10425);
nand U18305 (N_18305,N_14759,N_11741);
and U18306 (N_18306,N_11720,N_11796);
xor U18307 (N_18307,N_14397,N_11750);
and U18308 (N_18308,N_14391,N_10230);
and U18309 (N_18309,N_14095,N_13855);
or U18310 (N_18310,N_11658,N_11037);
xnor U18311 (N_18311,N_11983,N_13978);
nand U18312 (N_18312,N_11223,N_10444);
and U18313 (N_18313,N_12821,N_12972);
nand U18314 (N_18314,N_11488,N_11513);
nor U18315 (N_18315,N_14213,N_11880);
and U18316 (N_18316,N_14396,N_13184);
or U18317 (N_18317,N_11637,N_11233);
nor U18318 (N_18318,N_10229,N_12389);
nand U18319 (N_18319,N_13214,N_13560);
nor U18320 (N_18320,N_10025,N_12711);
or U18321 (N_18321,N_12643,N_10267);
nor U18322 (N_18322,N_12204,N_14818);
nand U18323 (N_18323,N_13225,N_12423);
and U18324 (N_18324,N_13358,N_11355);
xor U18325 (N_18325,N_10734,N_11935);
nor U18326 (N_18326,N_10383,N_13176);
nand U18327 (N_18327,N_13336,N_14895);
xor U18328 (N_18328,N_10298,N_11142);
and U18329 (N_18329,N_13230,N_13039);
nor U18330 (N_18330,N_12665,N_10547);
and U18331 (N_18331,N_13128,N_11711);
nor U18332 (N_18332,N_14881,N_14585);
nand U18333 (N_18333,N_13868,N_11925);
and U18334 (N_18334,N_11371,N_12571);
nor U18335 (N_18335,N_12388,N_12144);
and U18336 (N_18336,N_14712,N_13946);
nor U18337 (N_18337,N_11684,N_10402);
xor U18338 (N_18338,N_13679,N_14019);
or U18339 (N_18339,N_11223,N_11131);
or U18340 (N_18340,N_10649,N_10870);
and U18341 (N_18341,N_14490,N_14256);
xnor U18342 (N_18342,N_12734,N_11592);
nand U18343 (N_18343,N_12413,N_10459);
nor U18344 (N_18344,N_12649,N_12015);
and U18345 (N_18345,N_10408,N_14704);
xor U18346 (N_18346,N_10216,N_14558);
and U18347 (N_18347,N_13493,N_10726);
xnor U18348 (N_18348,N_12325,N_14976);
and U18349 (N_18349,N_13100,N_11085);
xor U18350 (N_18350,N_13541,N_10625);
nor U18351 (N_18351,N_11407,N_11219);
or U18352 (N_18352,N_10248,N_11289);
or U18353 (N_18353,N_13016,N_13945);
nand U18354 (N_18354,N_10338,N_13851);
and U18355 (N_18355,N_12488,N_11963);
nand U18356 (N_18356,N_10257,N_14338);
xor U18357 (N_18357,N_14040,N_12408);
nor U18358 (N_18358,N_11848,N_12411);
nand U18359 (N_18359,N_14469,N_12855);
nand U18360 (N_18360,N_10564,N_13170);
and U18361 (N_18361,N_10129,N_11841);
xnor U18362 (N_18362,N_13538,N_13130);
xnor U18363 (N_18363,N_13652,N_13923);
nand U18364 (N_18364,N_10247,N_10226);
or U18365 (N_18365,N_13655,N_11310);
nand U18366 (N_18366,N_10799,N_14679);
and U18367 (N_18367,N_14562,N_12059);
xor U18368 (N_18368,N_11832,N_10590);
nor U18369 (N_18369,N_14807,N_12206);
and U18370 (N_18370,N_12146,N_14856);
and U18371 (N_18371,N_12591,N_10940);
nand U18372 (N_18372,N_11559,N_11945);
nor U18373 (N_18373,N_11326,N_11009);
and U18374 (N_18374,N_12982,N_11762);
nor U18375 (N_18375,N_10144,N_12055);
xor U18376 (N_18376,N_10328,N_12355);
or U18377 (N_18377,N_14886,N_14756);
xor U18378 (N_18378,N_14971,N_11924);
xor U18379 (N_18379,N_13714,N_13049);
and U18380 (N_18380,N_12982,N_11870);
xor U18381 (N_18381,N_11343,N_12959);
and U18382 (N_18382,N_10179,N_13112);
nand U18383 (N_18383,N_11948,N_11203);
nor U18384 (N_18384,N_13822,N_13481);
xor U18385 (N_18385,N_12073,N_14176);
and U18386 (N_18386,N_10388,N_10368);
or U18387 (N_18387,N_11688,N_10344);
nand U18388 (N_18388,N_14363,N_14771);
nand U18389 (N_18389,N_10229,N_12100);
or U18390 (N_18390,N_11538,N_12156);
nor U18391 (N_18391,N_14334,N_10437);
nor U18392 (N_18392,N_14665,N_13474);
and U18393 (N_18393,N_13168,N_14789);
nor U18394 (N_18394,N_10819,N_14566);
and U18395 (N_18395,N_11232,N_14732);
and U18396 (N_18396,N_10713,N_11404);
or U18397 (N_18397,N_14839,N_14010);
and U18398 (N_18398,N_10335,N_10206);
and U18399 (N_18399,N_12136,N_10826);
and U18400 (N_18400,N_10233,N_11789);
or U18401 (N_18401,N_11322,N_11952);
xor U18402 (N_18402,N_14068,N_14074);
or U18403 (N_18403,N_13258,N_14717);
nand U18404 (N_18404,N_12161,N_10069);
nand U18405 (N_18405,N_12774,N_13159);
and U18406 (N_18406,N_12158,N_11466);
nand U18407 (N_18407,N_14976,N_12628);
xnor U18408 (N_18408,N_12721,N_13099);
and U18409 (N_18409,N_14254,N_11207);
or U18410 (N_18410,N_13389,N_13299);
nor U18411 (N_18411,N_12114,N_11435);
and U18412 (N_18412,N_10131,N_11564);
or U18413 (N_18413,N_12402,N_10755);
xnor U18414 (N_18414,N_13256,N_12066);
or U18415 (N_18415,N_11744,N_14442);
nand U18416 (N_18416,N_13075,N_13780);
xnor U18417 (N_18417,N_13947,N_14749);
and U18418 (N_18418,N_10299,N_10173);
nor U18419 (N_18419,N_14148,N_12415);
nand U18420 (N_18420,N_14644,N_13196);
nand U18421 (N_18421,N_11643,N_10458);
xor U18422 (N_18422,N_11078,N_13290);
nor U18423 (N_18423,N_11768,N_11498);
or U18424 (N_18424,N_14711,N_14456);
xor U18425 (N_18425,N_12048,N_13131);
or U18426 (N_18426,N_13439,N_14671);
nor U18427 (N_18427,N_12425,N_13610);
and U18428 (N_18428,N_11720,N_13757);
nor U18429 (N_18429,N_13305,N_12485);
and U18430 (N_18430,N_14038,N_10520);
xor U18431 (N_18431,N_11904,N_12448);
nor U18432 (N_18432,N_12679,N_12351);
nor U18433 (N_18433,N_13787,N_11845);
xnor U18434 (N_18434,N_12635,N_12012);
nor U18435 (N_18435,N_12674,N_12527);
and U18436 (N_18436,N_14608,N_14396);
or U18437 (N_18437,N_14242,N_10828);
and U18438 (N_18438,N_13034,N_13717);
xnor U18439 (N_18439,N_11286,N_14483);
and U18440 (N_18440,N_11316,N_11332);
or U18441 (N_18441,N_12373,N_13727);
and U18442 (N_18442,N_11433,N_10787);
xor U18443 (N_18443,N_14452,N_10775);
xnor U18444 (N_18444,N_11911,N_10905);
or U18445 (N_18445,N_13324,N_11203);
xnor U18446 (N_18446,N_14584,N_13576);
nor U18447 (N_18447,N_10222,N_13445);
nor U18448 (N_18448,N_14296,N_14719);
and U18449 (N_18449,N_13992,N_14900);
xnor U18450 (N_18450,N_10679,N_11851);
nand U18451 (N_18451,N_13105,N_12865);
and U18452 (N_18452,N_10894,N_13343);
xnor U18453 (N_18453,N_12003,N_11316);
nor U18454 (N_18454,N_11384,N_11674);
and U18455 (N_18455,N_12927,N_11332);
and U18456 (N_18456,N_14354,N_11637);
and U18457 (N_18457,N_11094,N_14574);
xnor U18458 (N_18458,N_14333,N_14145);
nand U18459 (N_18459,N_10545,N_12812);
xnor U18460 (N_18460,N_10457,N_11011);
nor U18461 (N_18461,N_13376,N_13250);
nand U18462 (N_18462,N_11151,N_11026);
xnor U18463 (N_18463,N_10338,N_10421);
xor U18464 (N_18464,N_12625,N_10428);
xor U18465 (N_18465,N_12485,N_12175);
nor U18466 (N_18466,N_13516,N_10604);
nand U18467 (N_18467,N_11946,N_13995);
or U18468 (N_18468,N_10546,N_14214);
xor U18469 (N_18469,N_14213,N_13351);
or U18470 (N_18470,N_10566,N_14785);
and U18471 (N_18471,N_14840,N_11430);
and U18472 (N_18472,N_12579,N_11284);
xor U18473 (N_18473,N_13844,N_14313);
xnor U18474 (N_18474,N_13740,N_14356);
or U18475 (N_18475,N_11990,N_14787);
nand U18476 (N_18476,N_11289,N_13893);
nor U18477 (N_18477,N_10278,N_10198);
nor U18478 (N_18478,N_12061,N_12911);
nor U18479 (N_18479,N_12948,N_11250);
and U18480 (N_18480,N_12334,N_12593);
nor U18481 (N_18481,N_12634,N_13116);
or U18482 (N_18482,N_13823,N_10415);
xnor U18483 (N_18483,N_12038,N_12144);
nor U18484 (N_18484,N_13311,N_10741);
xor U18485 (N_18485,N_13142,N_10502);
and U18486 (N_18486,N_13441,N_12429);
nor U18487 (N_18487,N_12396,N_12187);
nor U18488 (N_18488,N_12208,N_12550);
nand U18489 (N_18489,N_10982,N_12220);
nand U18490 (N_18490,N_11231,N_10640);
nor U18491 (N_18491,N_11257,N_10820);
and U18492 (N_18492,N_13817,N_14848);
or U18493 (N_18493,N_10552,N_11678);
nor U18494 (N_18494,N_12876,N_14069);
or U18495 (N_18495,N_10943,N_12669);
nand U18496 (N_18496,N_14430,N_10832);
nand U18497 (N_18497,N_10133,N_10327);
and U18498 (N_18498,N_13509,N_10420);
or U18499 (N_18499,N_11905,N_10771);
xnor U18500 (N_18500,N_13735,N_11048);
xnor U18501 (N_18501,N_14873,N_11461);
nand U18502 (N_18502,N_11729,N_12331);
xnor U18503 (N_18503,N_13263,N_13410);
or U18504 (N_18504,N_10662,N_13050);
nand U18505 (N_18505,N_14243,N_11412);
and U18506 (N_18506,N_11770,N_13277);
xor U18507 (N_18507,N_11531,N_13358);
nand U18508 (N_18508,N_13422,N_11487);
or U18509 (N_18509,N_13058,N_10240);
and U18510 (N_18510,N_12548,N_13854);
or U18511 (N_18511,N_13907,N_12842);
and U18512 (N_18512,N_11875,N_10362);
or U18513 (N_18513,N_14601,N_13590);
or U18514 (N_18514,N_12034,N_14424);
or U18515 (N_18515,N_10604,N_12793);
or U18516 (N_18516,N_11452,N_14087);
nor U18517 (N_18517,N_13960,N_11473);
nand U18518 (N_18518,N_11088,N_11725);
or U18519 (N_18519,N_11529,N_14368);
or U18520 (N_18520,N_10803,N_12211);
or U18521 (N_18521,N_14020,N_10422);
and U18522 (N_18522,N_11562,N_13068);
or U18523 (N_18523,N_10234,N_10298);
nand U18524 (N_18524,N_13611,N_11357);
nand U18525 (N_18525,N_11981,N_10965);
nor U18526 (N_18526,N_13659,N_11011);
and U18527 (N_18527,N_14591,N_10567);
and U18528 (N_18528,N_14276,N_11088);
nor U18529 (N_18529,N_10134,N_12294);
or U18530 (N_18530,N_12085,N_10409);
or U18531 (N_18531,N_10728,N_11298);
or U18532 (N_18532,N_11288,N_11133);
xor U18533 (N_18533,N_12366,N_14670);
and U18534 (N_18534,N_14633,N_13438);
nand U18535 (N_18535,N_14968,N_13688);
nand U18536 (N_18536,N_13937,N_11640);
xor U18537 (N_18537,N_10849,N_12650);
nor U18538 (N_18538,N_13773,N_10501);
xor U18539 (N_18539,N_13516,N_13443);
nand U18540 (N_18540,N_14377,N_11890);
nand U18541 (N_18541,N_14136,N_12075);
xnor U18542 (N_18542,N_10097,N_10626);
and U18543 (N_18543,N_12322,N_12967);
xor U18544 (N_18544,N_13385,N_14923);
xnor U18545 (N_18545,N_14336,N_13557);
xor U18546 (N_18546,N_10288,N_14767);
nand U18547 (N_18547,N_12835,N_10754);
or U18548 (N_18548,N_12252,N_10951);
xnor U18549 (N_18549,N_11479,N_13538);
and U18550 (N_18550,N_13587,N_12739);
and U18551 (N_18551,N_10616,N_11029);
or U18552 (N_18552,N_10726,N_14389);
or U18553 (N_18553,N_10529,N_11183);
or U18554 (N_18554,N_12584,N_14662);
and U18555 (N_18555,N_12423,N_14372);
nor U18556 (N_18556,N_13222,N_14713);
or U18557 (N_18557,N_12665,N_14190);
xnor U18558 (N_18558,N_10200,N_12046);
nor U18559 (N_18559,N_14469,N_13510);
nor U18560 (N_18560,N_14978,N_14081);
or U18561 (N_18561,N_14116,N_11561);
nand U18562 (N_18562,N_14592,N_13076);
and U18563 (N_18563,N_14888,N_11208);
nor U18564 (N_18564,N_11070,N_13776);
nor U18565 (N_18565,N_10145,N_13172);
nor U18566 (N_18566,N_12211,N_11981);
nand U18567 (N_18567,N_13594,N_12925);
nor U18568 (N_18568,N_13735,N_11300);
nor U18569 (N_18569,N_14760,N_14365);
nand U18570 (N_18570,N_13951,N_14477);
nand U18571 (N_18571,N_11259,N_12637);
and U18572 (N_18572,N_14900,N_11852);
or U18573 (N_18573,N_13849,N_13451);
and U18574 (N_18574,N_13682,N_11527);
nand U18575 (N_18575,N_10585,N_13885);
and U18576 (N_18576,N_10962,N_14488);
xor U18577 (N_18577,N_14404,N_13535);
and U18578 (N_18578,N_12035,N_14133);
xnor U18579 (N_18579,N_10249,N_12056);
and U18580 (N_18580,N_14458,N_14481);
or U18581 (N_18581,N_11537,N_11793);
xor U18582 (N_18582,N_14012,N_11861);
nor U18583 (N_18583,N_12938,N_11651);
nor U18584 (N_18584,N_11734,N_10054);
xnor U18585 (N_18585,N_14894,N_10922);
xor U18586 (N_18586,N_10663,N_11868);
and U18587 (N_18587,N_10894,N_12897);
nand U18588 (N_18588,N_11827,N_10558);
or U18589 (N_18589,N_14788,N_14838);
and U18590 (N_18590,N_12340,N_11946);
xor U18591 (N_18591,N_12205,N_13341);
nor U18592 (N_18592,N_14488,N_14907);
or U18593 (N_18593,N_12638,N_12793);
nor U18594 (N_18594,N_14534,N_14269);
and U18595 (N_18595,N_10917,N_12567);
nand U18596 (N_18596,N_10402,N_14505);
nand U18597 (N_18597,N_13623,N_14311);
and U18598 (N_18598,N_14295,N_13746);
nand U18599 (N_18599,N_14697,N_13620);
or U18600 (N_18600,N_14980,N_12883);
nor U18601 (N_18601,N_11417,N_13643);
nand U18602 (N_18602,N_14928,N_13290);
xnor U18603 (N_18603,N_13993,N_13931);
and U18604 (N_18604,N_11046,N_11814);
nor U18605 (N_18605,N_11279,N_14876);
and U18606 (N_18606,N_13074,N_10055);
or U18607 (N_18607,N_11738,N_10952);
or U18608 (N_18608,N_12814,N_11439);
and U18609 (N_18609,N_12422,N_14168);
and U18610 (N_18610,N_13617,N_10367);
and U18611 (N_18611,N_14090,N_11263);
nand U18612 (N_18612,N_12627,N_10402);
nor U18613 (N_18613,N_12981,N_13541);
or U18614 (N_18614,N_12044,N_12991);
and U18615 (N_18615,N_13908,N_12606);
nand U18616 (N_18616,N_10508,N_13777);
or U18617 (N_18617,N_11493,N_14537);
and U18618 (N_18618,N_13753,N_12534);
xor U18619 (N_18619,N_12263,N_12970);
nand U18620 (N_18620,N_11214,N_11768);
xnor U18621 (N_18621,N_10019,N_11728);
or U18622 (N_18622,N_10430,N_13859);
nand U18623 (N_18623,N_14856,N_10044);
nand U18624 (N_18624,N_11548,N_11962);
nand U18625 (N_18625,N_12093,N_14540);
nand U18626 (N_18626,N_12997,N_10037);
or U18627 (N_18627,N_10814,N_11667);
nand U18628 (N_18628,N_10379,N_11411);
nand U18629 (N_18629,N_11235,N_10573);
nor U18630 (N_18630,N_13537,N_12573);
xor U18631 (N_18631,N_12738,N_12223);
and U18632 (N_18632,N_13247,N_13210);
or U18633 (N_18633,N_14856,N_12404);
nand U18634 (N_18634,N_13045,N_10685);
or U18635 (N_18635,N_10000,N_12181);
and U18636 (N_18636,N_11549,N_14959);
or U18637 (N_18637,N_14340,N_12558);
nor U18638 (N_18638,N_11718,N_14179);
or U18639 (N_18639,N_10761,N_11889);
xnor U18640 (N_18640,N_13929,N_10839);
xnor U18641 (N_18641,N_12545,N_12042);
and U18642 (N_18642,N_11322,N_12051);
and U18643 (N_18643,N_14670,N_12959);
and U18644 (N_18644,N_13910,N_13129);
nor U18645 (N_18645,N_14916,N_13505);
xnor U18646 (N_18646,N_14009,N_14532);
nor U18647 (N_18647,N_11563,N_14230);
nand U18648 (N_18648,N_13504,N_11233);
xor U18649 (N_18649,N_10571,N_13542);
nand U18650 (N_18650,N_10574,N_13496);
and U18651 (N_18651,N_13894,N_12603);
or U18652 (N_18652,N_13531,N_10535);
and U18653 (N_18653,N_14359,N_12019);
and U18654 (N_18654,N_14468,N_11238);
nor U18655 (N_18655,N_14539,N_10850);
nand U18656 (N_18656,N_14469,N_13952);
xor U18657 (N_18657,N_11764,N_12313);
xor U18658 (N_18658,N_14730,N_12076);
nand U18659 (N_18659,N_13907,N_13829);
nor U18660 (N_18660,N_11561,N_14441);
and U18661 (N_18661,N_11419,N_14577);
and U18662 (N_18662,N_14377,N_12734);
xnor U18663 (N_18663,N_11388,N_10087);
nor U18664 (N_18664,N_13998,N_11351);
or U18665 (N_18665,N_11216,N_14987);
xnor U18666 (N_18666,N_11595,N_11941);
nand U18667 (N_18667,N_11158,N_13505);
or U18668 (N_18668,N_11784,N_14106);
nor U18669 (N_18669,N_11831,N_12597);
and U18670 (N_18670,N_11778,N_11386);
or U18671 (N_18671,N_14875,N_14137);
xnor U18672 (N_18672,N_10012,N_12870);
nor U18673 (N_18673,N_14861,N_12155);
or U18674 (N_18674,N_10248,N_12749);
nor U18675 (N_18675,N_14255,N_13297);
nand U18676 (N_18676,N_13320,N_14640);
nor U18677 (N_18677,N_12188,N_13573);
nand U18678 (N_18678,N_10178,N_13758);
xor U18679 (N_18679,N_13501,N_14336);
nor U18680 (N_18680,N_12969,N_10110);
or U18681 (N_18681,N_12247,N_13838);
and U18682 (N_18682,N_10319,N_10495);
nand U18683 (N_18683,N_10322,N_11031);
nand U18684 (N_18684,N_13491,N_14838);
or U18685 (N_18685,N_14370,N_14452);
nor U18686 (N_18686,N_11692,N_10951);
xnor U18687 (N_18687,N_12261,N_13384);
or U18688 (N_18688,N_12609,N_12589);
and U18689 (N_18689,N_12369,N_12112);
nand U18690 (N_18690,N_12437,N_12164);
nor U18691 (N_18691,N_13480,N_14370);
xnor U18692 (N_18692,N_12180,N_12528);
nand U18693 (N_18693,N_14131,N_11154);
xnor U18694 (N_18694,N_11659,N_12470);
and U18695 (N_18695,N_14844,N_13886);
and U18696 (N_18696,N_11044,N_14817);
nor U18697 (N_18697,N_10486,N_10396);
and U18698 (N_18698,N_11682,N_13523);
nand U18699 (N_18699,N_12963,N_12495);
or U18700 (N_18700,N_13991,N_10358);
and U18701 (N_18701,N_14545,N_11881);
xor U18702 (N_18702,N_11118,N_14471);
nand U18703 (N_18703,N_13805,N_10846);
nor U18704 (N_18704,N_13149,N_14393);
or U18705 (N_18705,N_10358,N_10523);
nand U18706 (N_18706,N_12779,N_14393);
nor U18707 (N_18707,N_11561,N_13772);
nand U18708 (N_18708,N_13791,N_12555);
and U18709 (N_18709,N_12032,N_13544);
nand U18710 (N_18710,N_12905,N_13068);
nor U18711 (N_18711,N_12049,N_13126);
xnor U18712 (N_18712,N_10742,N_13343);
and U18713 (N_18713,N_12342,N_14793);
xnor U18714 (N_18714,N_14638,N_14818);
nor U18715 (N_18715,N_12674,N_12129);
xor U18716 (N_18716,N_13104,N_14344);
or U18717 (N_18717,N_10642,N_14880);
xnor U18718 (N_18718,N_13645,N_14115);
xnor U18719 (N_18719,N_10708,N_12187);
and U18720 (N_18720,N_14622,N_14585);
nand U18721 (N_18721,N_10533,N_13034);
nand U18722 (N_18722,N_12958,N_13717);
or U18723 (N_18723,N_11246,N_14919);
and U18724 (N_18724,N_11508,N_14339);
xnor U18725 (N_18725,N_14279,N_14425);
xnor U18726 (N_18726,N_10499,N_12940);
or U18727 (N_18727,N_14984,N_14531);
nor U18728 (N_18728,N_13239,N_10870);
nor U18729 (N_18729,N_11335,N_14706);
nor U18730 (N_18730,N_10533,N_10175);
or U18731 (N_18731,N_10413,N_14435);
nand U18732 (N_18732,N_13675,N_14735);
nor U18733 (N_18733,N_10515,N_13998);
xor U18734 (N_18734,N_13398,N_12581);
nor U18735 (N_18735,N_12780,N_14634);
or U18736 (N_18736,N_10834,N_13058);
and U18737 (N_18737,N_13059,N_12832);
nor U18738 (N_18738,N_12712,N_12623);
nand U18739 (N_18739,N_12640,N_10993);
xnor U18740 (N_18740,N_14357,N_11429);
nand U18741 (N_18741,N_12270,N_13088);
or U18742 (N_18742,N_13023,N_11000);
or U18743 (N_18743,N_11198,N_12097);
or U18744 (N_18744,N_14723,N_11554);
or U18745 (N_18745,N_12201,N_11105);
or U18746 (N_18746,N_13129,N_12951);
nand U18747 (N_18747,N_12977,N_13883);
nand U18748 (N_18748,N_10127,N_13442);
or U18749 (N_18749,N_13737,N_12780);
nor U18750 (N_18750,N_13756,N_11781);
nand U18751 (N_18751,N_10113,N_11738);
nor U18752 (N_18752,N_13657,N_10243);
nand U18753 (N_18753,N_12252,N_14636);
nand U18754 (N_18754,N_11011,N_12994);
or U18755 (N_18755,N_10944,N_12537);
nand U18756 (N_18756,N_12450,N_14459);
nand U18757 (N_18757,N_11496,N_13474);
xor U18758 (N_18758,N_12518,N_13751);
xor U18759 (N_18759,N_14726,N_14563);
or U18760 (N_18760,N_12115,N_13178);
xnor U18761 (N_18761,N_12424,N_12956);
nor U18762 (N_18762,N_13747,N_13631);
nor U18763 (N_18763,N_12931,N_10017);
nand U18764 (N_18764,N_14105,N_12090);
nand U18765 (N_18765,N_14761,N_13482);
nand U18766 (N_18766,N_14415,N_12615);
or U18767 (N_18767,N_10558,N_11551);
and U18768 (N_18768,N_12558,N_10945);
and U18769 (N_18769,N_12985,N_13735);
and U18770 (N_18770,N_11978,N_14052);
or U18771 (N_18771,N_11730,N_13347);
or U18772 (N_18772,N_11275,N_11466);
nand U18773 (N_18773,N_13660,N_10786);
nand U18774 (N_18774,N_14169,N_12188);
nor U18775 (N_18775,N_13455,N_14279);
and U18776 (N_18776,N_14054,N_14237);
nor U18777 (N_18777,N_10649,N_12405);
nor U18778 (N_18778,N_10581,N_10899);
nor U18779 (N_18779,N_12338,N_11106);
nand U18780 (N_18780,N_12913,N_12674);
nand U18781 (N_18781,N_11095,N_12074);
nor U18782 (N_18782,N_14743,N_11793);
or U18783 (N_18783,N_10345,N_11057);
nor U18784 (N_18784,N_10835,N_10914);
and U18785 (N_18785,N_10786,N_14026);
nand U18786 (N_18786,N_13864,N_14592);
or U18787 (N_18787,N_11770,N_12812);
nor U18788 (N_18788,N_14411,N_10755);
xnor U18789 (N_18789,N_10984,N_12382);
and U18790 (N_18790,N_13739,N_12817);
nand U18791 (N_18791,N_11344,N_14017);
or U18792 (N_18792,N_12667,N_14102);
xor U18793 (N_18793,N_12921,N_11984);
or U18794 (N_18794,N_12566,N_14436);
xnor U18795 (N_18795,N_11707,N_14467);
and U18796 (N_18796,N_13430,N_12150);
nor U18797 (N_18797,N_13701,N_12168);
nand U18798 (N_18798,N_14158,N_12707);
nand U18799 (N_18799,N_12029,N_14304);
and U18800 (N_18800,N_10343,N_10254);
nor U18801 (N_18801,N_12224,N_12978);
and U18802 (N_18802,N_10374,N_11953);
or U18803 (N_18803,N_11122,N_11988);
nand U18804 (N_18804,N_10723,N_13277);
or U18805 (N_18805,N_12237,N_13463);
xnor U18806 (N_18806,N_12707,N_10526);
nor U18807 (N_18807,N_14719,N_12202);
and U18808 (N_18808,N_11657,N_11468);
nand U18809 (N_18809,N_11036,N_10428);
xnor U18810 (N_18810,N_14845,N_11397);
nand U18811 (N_18811,N_11875,N_10102);
and U18812 (N_18812,N_13745,N_12862);
and U18813 (N_18813,N_13950,N_13464);
nor U18814 (N_18814,N_12607,N_13684);
xor U18815 (N_18815,N_10064,N_14340);
nand U18816 (N_18816,N_13235,N_14405);
xor U18817 (N_18817,N_14606,N_12204);
xnor U18818 (N_18818,N_14746,N_11620);
xor U18819 (N_18819,N_10764,N_14823);
and U18820 (N_18820,N_14262,N_10211);
xnor U18821 (N_18821,N_10952,N_10560);
and U18822 (N_18822,N_14447,N_13714);
or U18823 (N_18823,N_11876,N_11938);
nor U18824 (N_18824,N_13361,N_13562);
and U18825 (N_18825,N_14751,N_11901);
or U18826 (N_18826,N_13303,N_11704);
and U18827 (N_18827,N_13608,N_13373);
or U18828 (N_18828,N_13271,N_14303);
xnor U18829 (N_18829,N_12236,N_10862);
nand U18830 (N_18830,N_10234,N_10902);
nand U18831 (N_18831,N_10658,N_11882);
nand U18832 (N_18832,N_12724,N_14202);
nand U18833 (N_18833,N_13879,N_11795);
xor U18834 (N_18834,N_12457,N_14663);
or U18835 (N_18835,N_11237,N_11343);
nor U18836 (N_18836,N_14325,N_13226);
nand U18837 (N_18837,N_12577,N_14754);
and U18838 (N_18838,N_10698,N_14833);
xnor U18839 (N_18839,N_14491,N_11823);
xor U18840 (N_18840,N_14902,N_11794);
xor U18841 (N_18841,N_10829,N_12672);
and U18842 (N_18842,N_10694,N_12591);
nor U18843 (N_18843,N_12521,N_13555);
xnor U18844 (N_18844,N_10501,N_13110);
and U18845 (N_18845,N_13387,N_13579);
xor U18846 (N_18846,N_11072,N_14748);
nand U18847 (N_18847,N_13098,N_13267);
and U18848 (N_18848,N_14233,N_12702);
or U18849 (N_18849,N_10859,N_12069);
xnor U18850 (N_18850,N_14870,N_10067);
nand U18851 (N_18851,N_14534,N_13208);
nand U18852 (N_18852,N_14768,N_13276);
nand U18853 (N_18853,N_11579,N_11926);
nor U18854 (N_18854,N_11474,N_12380);
and U18855 (N_18855,N_13957,N_10092);
nor U18856 (N_18856,N_12219,N_14200);
xnor U18857 (N_18857,N_13584,N_12805);
nor U18858 (N_18858,N_14786,N_11366);
nand U18859 (N_18859,N_10717,N_13135);
or U18860 (N_18860,N_14790,N_10964);
nor U18861 (N_18861,N_13877,N_11863);
and U18862 (N_18862,N_13767,N_12123);
nand U18863 (N_18863,N_14285,N_14124);
nand U18864 (N_18864,N_10550,N_10191);
xor U18865 (N_18865,N_11001,N_14973);
xor U18866 (N_18866,N_13786,N_10629);
nor U18867 (N_18867,N_11153,N_11098);
or U18868 (N_18868,N_12124,N_11741);
xnor U18869 (N_18869,N_10532,N_14382);
nand U18870 (N_18870,N_13806,N_10509);
xnor U18871 (N_18871,N_11035,N_11550);
nor U18872 (N_18872,N_13416,N_14147);
nand U18873 (N_18873,N_10879,N_14175);
and U18874 (N_18874,N_10495,N_12204);
nand U18875 (N_18875,N_11226,N_12049);
xnor U18876 (N_18876,N_14480,N_11891);
nand U18877 (N_18877,N_12458,N_14327);
xnor U18878 (N_18878,N_10710,N_12562);
and U18879 (N_18879,N_14223,N_10597);
nor U18880 (N_18880,N_14874,N_13761);
nand U18881 (N_18881,N_12869,N_14224);
nor U18882 (N_18882,N_14843,N_10787);
xnor U18883 (N_18883,N_12783,N_12028);
nand U18884 (N_18884,N_13215,N_10807);
nand U18885 (N_18885,N_13968,N_12716);
and U18886 (N_18886,N_12790,N_10882);
and U18887 (N_18887,N_10293,N_13272);
nand U18888 (N_18888,N_13250,N_11895);
nor U18889 (N_18889,N_14297,N_11407);
xnor U18890 (N_18890,N_11929,N_11966);
and U18891 (N_18891,N_13079,N_11928);
nand U18892 (N_18892,N_12213,N_13182);
nor U18893 (N_18893,N_11153,N_12844);
or U18894 (N_18894,N_11018,N_10388);
nand U18895 (N_18895,N_13204,N_10203);
xnor U18896 (N_18896,N_13681,N_10890);
or U18897 (N_18897,N_12292,N_12617);
xnor U18898 (N_18898,N_13678,N_14623);
nor U18899 (N_18899,N_11940,N_13303);
nor U18900 (N_18900,N_14834,N_11877);
and U18901 (N_18901,N_10410,N_11697);
nand U18902 (N_18902,N_11763,N_12434);
or U18903 (N_18903,N_10074,N_14759);
and U18904 (N_18904,N_11316,N_12039);
xnor U18905 (N_18905,N_13324,N_11701);
and U18906 (N_18906,N_13678,N_13683);
nand U18907 (N_18907,N_13786,N_13477);
and U18908 (N_18908,N_11966,N_11931);
xor U18909 (N_18909,N_10856,N_10998);
nand U18910 (N_18910,N_10821,N_13830);
nand U18911 (N_18911,N_12247,N_14670);
nor U18912 (N_18912,N_14223,N_12224);
and U18913 (N_18913,N_10868,N_10853);
and U18914 (N_18914,N_11045,N_10804);
xor U18915 (N_18915,N_10243,N_12521);
xor U18916 (N_18916,N_14967,N_10652);
nor U18917 (N_18917,N_11840,N_13176);
or U18918 (N_18918,N_12791,N_14306);
or U18919 (N_18919,N_13824,N_14219);
nand U18920 (N_18920,N_14195,N_12968);
and U18921 (N_18921,N_11992,N_11368);
or U18922 (N_18922,N_10094,N_10028);
nand U18923 (N_18923,N_11289,N_12746);
xnor U18924 (N_18924,N_12554,N_10257);
nor U18925 (N_18925,N_13683,N_14316);
or U18926 (N_18926,N_12614,N_14726);
and U18927 (N_18927,N_11897,N_12477);
nor U18928 (N_18928,N_12935,N_14161);
and U18929 (N_18929,N_11073,N_10005);
nand U18930 (N_18930,N_10692,N_14666);
and U18931 (N_18931,N_11853,N_10653);
or U18932 (N_18932,N_14166,N_13839);
or U18933 (N_18933,N_12824,N_13427);
and U18934 (N_18934,N_13912,N_10690);
xor U18935 (N_18935,N_11527,N_13598);
nor U18936 (N_18936,N_11291,N_13562);
or U18937 (N_18937,N_13134,N_10986);
and U18938 (N_18938,N_12254,N_12742);
nand U18939 (N_18939,N_12403,N_13650);
or U18940 (N_18940,N_14165,N_13465);
or U18941 (N_18941,N_14892,N_12544);
nor U18942 (N_18942,N_10250,N_11526);
xnor U18943 (N_18943,N_13993,N_13386);
nor U18944 (N_18944,N_12201,N_13890);
xor U18945 (N_18945,N_11928,N_12997);
xor U18946 (N_18946,N_14208,N_12386);
nor U18947 (N_18947,N_10351,N_12469);
nor U18948 (N_18948,N_13902,N_12985);
nand U18949 (N_18949,N_13758,N_14540);
nand U18950 (N_18950,N_12824,N_11387);
xnor U18951 (N_18951,N_14482,N_14194);
xnor U18952 (N_18952,N_11661,N_12417);
or U18953 (N_18953,N_14429,N_14013);
xor U18954 (N_18954,N_14702,N_10036);
and U18955 (N_18955,N_10357,N_10248);
nor U18956 (N_18956,N_10892,N_11508);
nor U18957 (N_18957,N_11371,N_13289);
nor U18958 (N_18958,N_14613,N_13625);
or U18959 (N_18959,N_10170,N_11947);
and U18960 (N_18960,N_14204,N_13449);
or U18961 (N_18961,N_14656,N_14586);
xnor U18962 (N_18962,N_13418,N_11419);
and U18963 (N_18963,N_13985,N_11073);
xnor U18964 (N_18964,N_10415,N_14797);
xnor U18965 (N_18965,N_14439,N_10799);
nand U18966 (N_18966,N_14146,N_13785);
nand U18967 (N_18967,N_10164,N_11576);
or U18968 (N_18968,N_10909,N_10888);
nor U18969 (N_18969,N_11527,N_14033);
xnor U18970 (N_18970,N_12119,N_11304);
xor U18971 (N_18971,N_12609,N_11012);
and U18972 (N_18972,N_14798,N_14861);
xnor U18973 (N_18973,N_12783,N_14022);
and U18974 (N_18974,N_13415,N_14249);
nor U18975 (N_18975,N_11896,N_10799);
and U18976 (N_18976,N_14896,N_13572);
xnor U18977 (N_18977,N_11823,N_13401);
nor U18978 (N_18978,N_10746,N_11568);
xor U18979 (N_18979,N_12054,N_14479);
nand U18980 (N_18980,N_11406,N_13367);
or U18981 (N_18981,N_10448,N_10036);
xnor U18982 (N_18982,N_13082,N_14590);
nand U18983 (N_18983,N_11540,N_14917);
or U18984 (N_18984,N_12527,N_11098);
nand U18985 (N_18985,N_14881,N_12774);
or U18986 (N_18986,N_13319,N_13893);
or U18987 (N_18987,N_13072,N_12313);
xor U18988 (N_18988,N_14726,N_11416);
or U18989 (N_18989,N_11627,N_13469);
and U18990 (N_18990,N_14727,N_10624);
nand U18991 (N_18991,N_14173,N_14933);
nand U18992 (N_18992,N_13800,N_11457);
nor U18993 (N_18993,N_11958,N_11242);
or U18994 (N_18994,N_11317,N_12765);
nand U18995 (N_18995,N_13251,N_13764);
nor U18996 (N_18996,N_10816,N_14590);
nor U18997 (N_18997,N_10317,N_11641);
nor U18998 (N_18998,N_13781,N_14740);
nand U18999 (N_18999,N_11261,N_10095);
and U19000 (N_19000,N_13491,N_13073);
nand U19001 (N_19001,N_14837,N_11162);
or U19002 (N_19002,N_11117,N_14214);
nand U19003 (N_19003,N_11731,N_14234);
or U19004 (N_19004,N_12949,N_14916);
or U19005 (N_19005,N_12523,N_12971);
nor U19006 (N_19006,N_10117,N_14385);
nand U19007 (N_19007,N_14726,N_11043);
and U19008 (N_19008,N_10719,N_12404);
or U19009 (N_19009,N_14967,N_14576);
and U19010 (N_19010,N_14653,N_12274);
xnor U19011 (N_19011,N_11128,N_13097);
or U19012 (N_19012,N_11156,N_14684);
and U19013 (N_19013,N_11198,N_13067);
nand U19014 (N_19014,N_12885,N_12417);
nand U19015 (N_19015,N_10494,N_12079);
and U19016 (N_19016,N_13061,N_13507);
xor U19017 (N_19017,N_13376,N_10748);
and U19018 (N_19018,N_11515,N_13547);
nand U19019 (N_19019,N_14798,N_14744);
and U19020 (N_19020,N_12152,N_14305);
nor U19021 (N_19021,N_13898,N_11527);
and U19022 (N_19022,N_14529,N_10885);
xor U19023 (N_19023,N_11990,N_12565);
xor U19024 (N_19024,N_10557,N_11908);
nor U19025 (N_19025,N_14830,N_11912);
xor U19026 (N_19026,N_13309,N_14959);
or U19027 (N_19027,N_12747,N_12120);
nor U19028 (N_19028,N_14404,N_13443);
or U19029 (N_19029,N_13869,N_10412);
nor U19030 (N_19030,N_12820,N_13158);
nand U19031 (N_19031,N_14953,N_12614);
and U19032 (N_19032,N_12281,N_14739);
or U19033 (N_19033,N_12950,N_12941);
xnor U19034 (N_19034,N_11025,N_13662);
nor U19035 (N_19035,N_12387,N_12814);
or U19036 (N_19036,N_12166,N_10187);
nand U19037 (N_19037,N_11398,N_12409);
nor U19038 (N_19038,N_10686,N_11063);
nand U19039 (N_19039,N_13796,N_11358);
or U19040 (N_19040,N_10145,N_13853);
nand U19041 (N_19041,N_11118,N_11731);
xor U19042 (N_19042,N_12147,N_11407);
and U19043 (N_19043,N_10529,N_13230);
xor U19044 (N_19044,N_14557,N_13962);
and U19045 (N_19045,N_14701,N_10201);
xnor U19046 (N_19046,N_13019,N_14813);
nand U19047 (N_19047,N_14828,N_10845);
xnor U19048 (N_19048,N_14619,N_10295);
or U19049 (N_19049,N_13012,N_10098);
and U19050 (N_19050,N_11560,N_11971);
or U19051 (N_19051,N_13110,N_12319);
and U19052 (N_19052,N_11138,N_10799);
nand U19053 (N_19053,N_14365,N_10759);
nand U19054 (N_19054,N_13626,N_10858);
xnor U19055 (N_19055,N_10544,N_10336);
nor U19056 (N_19056,N_11952,N_11738);
or U19057 (N_19057,N_11833,N_13814);
xnor U19058 (N_19058,N_12627,N_13313);
xnor U19059 (N_19059,N_13134,N_12218);
and U19060 (N_19060,N_14285,N_14147);
nor U19061 (N_19061,N_11423,N_12895);
xnor U19062 (N_19062,N_13506,N_14296);
nand U19063 (N_19063,N_10226,N_10410);
or U19064 (N_19064,N_10662,N_10202);
and U19065 (N_19065,N_12265,N_10933);
nand U19066 (N_19066,N_11384,N_12836);
nor U19067 (N_19067,N_12384,N_10647);
and U19068 (N_19068,N_10883,N_10730);
and U19069 (N_19069,N_11199,N_11316);
and U19070 (N_19070,N_10098,N_13403);
nand U19071 (N_19071,N_10994,N_11853);
xnor U19072 (N_19072,N_11685,N_13406);
or U19073 (N_19073,N_10249,N_12965);
nand U19074 (N_19074,N_10108,N_10021);
xnor U19075 (N_19075,N_12944,N_12669);
nor U19076 (N_19076,N_12464,N_11863);
xnor U19077 (N_19077,N_12072,N_14186);
xnor U19078 (N_19078,N_12422,N_12695);
nor U19079 (N_19079,N_10894,N_12498);
nor U19080 (N_19080,N_11574,N_13151);
nor U19081 (N_19081,N_14394,N_11197);
or U19082 (N_19082,N_10411,N_12246);
xnor U19083 (N_19083,N_14018,N_13565);
xnor U19084 (N_19084,N_13274,N_14046);
xnor U19085 (N_19085,N_11963,N_12610);
xnor U19086 (N_19086,N_13029,N_11702);
and U19087 (N_19087,N_14904,N_14395);
or U19088 (N_19088,N_11583,N_10403);
or U19089 (N_19089,N_11625,N_12326);
or U19090 (N_19090,N_10460,N_12217);
and U19091 (N_19091,N_11689,N_10876);
or U19092 (N_19092,N_13476,N_14259);
and U19093 (N_19093,N_11982,N_11249);
nand U19094 (N_19094,N_13456,N_12671);
nor U19095 (N_19095,N_13863,N_11275);
nand U19096 (N_19096,N_12197,N_11654);
nand U19097 (N_19097,N_11617,N_14220);
or U19098 (N_19098,N_10018,N_13807);
nor U19099 (N_19099,N_13128,N_14798);
or U19100 (N_19100,N_10998,N_14039);
and U19101 (N_19101,N_14478,N_13662);
or U19102 (N_19102,N_13635,N_11843);
and U19103 (N_19103,N_10378,N_12509);
or U19104 (N_19104,N_11515,N_12733);
nand U19105 (N_19105,N_11088,N_10615);
nor U19106 (N_19106,N_13574,N_13686);
and U19107 (N_19107,N_11652,N_11972);
nand U19108 (N_19108,N_14863,N_14927);
and U19109 (N_19109,N_11256,N_13137);
nor U19110 (N_19110,N_13958,N_14689);
and U19111 (N_19111,N_13964,N_11310);
and U19112 (N_19112,N_11329,N_10536);
or U19113 (N_19113,N_11013,N_13357);
and U19114 (N_19114,N_13636,N_13274);
xnor U19115 (N_19115,N_10762,N_10860);
and U19116 (N_19116,N_13555,N_11946);
nand U19117 (N_19117,N_12670,N_14062);
or U19118 (N_19118,N_10704,N_12977);
nand U19119 (N_19119,N_10979,N_10750);
or U19120 (N_19120,N_12893,N_10944);
and U19121 (N_19121,N_12950,N_11825);
or U19122 (N_19122,N_11790,N_11358);
nor U19123 (N_19123,N_11052,N_11973);
xor U19124 (N_19124,N_12133,N_10274);
xor U19125 (N_19125,N_10903,N_12145);
nor U19126 (N_19126,N_14643,N_12281);
and U19127 (N_19127,N_14759,N_13462);
nand U19128 (N_19128,N_12682,N_11156);
nand U19129 (N_19129,N_12351,N_11211);
nand U19130 (N_19130,N_14813,N_13970);
nor U19131 (N_19131,N_14346,N_13029);
xor U19132 (N_19132,N_13467,N_13157);
xor U19133 (N_19133,N_11064,N_13200);
nor U19134 (N_19134,N_10679,N_12369);
nor U19135 (N_19135,N_12942,N_10467);
xor U19136 (N_19136,N_10788,N_12267);
nor U19137 (N_19137,N_14015,N_12824);
or U19138 (N_19138,N_10616,N_10489);
or U19139 (N_19139,N_12891,N_11429);
nand U19140 (N_19140,N_14502,N_12441);
nor U19141 (N_19141,N_10176,N_13819);
nand U19142 (N_19142,N_12716,N_10433);
nor U19143 (N_19143,N_11757,N_12532);
or U19144 (N_19144,N_12759,N_13594);
or U19145 (N_19145,N_12100,N_11975);
nand U19146 (N_19146,N_14384,N_11914);
or U19147 (N_19147,N_14979,N_14349);
nor U19148 (N_19148,N_11396,N_13085);
nand U19149 (N_19149,N_11089,N_14483);
nand U19150 (N_19150,N_10246,N_12060);
xor U19151 (N_19151,N_14552,N_10980);
nand U19152 (N_19152,N_10500,N_10887);
xnor U19153 (N_19153,N_12818,N_12776);
or U19154 (N_19154,N_14070,N_13829);
nor U19155 (N_19155,N_14682,N_13513);
and U19156 (N_19156,N_13086,N_14650);
or U19157 (N_19157,N_10523,N_13901);
nand U19158 (N_19158,N_13707,N_11051);
and U19159 (N_19159,N_10368,N_12657);
and U19160 (N_19160,N_12933,N_11476);
and U19161 (N_19161,N_13462,N_11411);
nand U19162 (N_19162,N_11237,N_11373);
nand U19163 (N_19163,N_12941,N_12238);
nor U19164 (N_19164,N_12013,N_10961);
nor U19165 (N_19165,N_12041,N_13045);
xor U19166 (N_19166,N_14048,N_14122);
and U19167 (N_19167,N_14893,N_13903);
xor U19168 (N_19168,N_14222,N_13739);
and U19169 (N_19169,N_14821,N_12606);
xor U19170 (N_19170,N_12567,N_11113);
xor U19171 (N_19171,N_14351,N_10954);
nor U19172 (N_19172,N_12320,N_11534);
xnor U19173 (N_19173,N_12584,N_10961);
and U19174 (N_19174,N_10674,N_13748);
or U19175 (N_19175,N_11139,N_11369);
xnor U19176 (N_19176,N_14150,N_13129);
or U19177 (N_19177,N_12403,N_10849);
xnor U19178 (N_19178,N_10229,N_14710);
nand U19179 (N_19179,N_11619,N_13826);
nand U19180 (N_19180,N_14765,N_10032);
xnor U19181 (N_19181,N_14376,N_14519);
nor U19182 (N_19182,N_14192,N_10391);
xnor U19183 (N_19183,N_14872,N_14787);
xor U19184 (N_19184,N_10325,N_14356);
nand U19185 (N_19185,N_12705,N_10702);
and U19186 (N_19186,N_13565,N_10829);
nand U19187 (N_19187,N_12748,N_14917);
or U19188 (N_19188,N_14441,N_10601);
and U19189 (N_19189,N_12100,N_13347);
xnor U19190 (N_19190,N_10424,N_13302);
nor U19191 (N_19191,N_14184,N_13526);
or U19192 (N_19192,N_11858,N_11991);
and U19193 (N_19193,N_12777,N_12930);
nor U19194 (N_19194,N_14906,N_11822);
nand U19195 (N_19195,N_11015,N_11252);
nor U19196 (N_19196,N_11516,N_14110);
nand U19197 (N_19197,N_11102,N_10385);
or U19198 (N_19198,N_13859,N_10718);
nor U19199 (N_19199,N_14152,N_10815);
nor U19200 (N_19200,N_14675,N_13558);
or U19201 (N_19201,N_11407,N_10884);
or U19202 (N_19202,N_14669,N_13893);
nor U19203 (N_19203,N_11959,N_12207);
nor U19204 (N_19204,N_14604,N_10800);
or U19205 (N_19205,N_13414,N_14582);
or U19206 (N_19206,N_11274,N_12803);
and U19207 (N_19207,N_13119,N_14487);
or U19208 (N_19208,N_11712,N_14027);
or U19209 (N_19209,N_14829,N_14566);
xor U19210 (N_19210,N_12453,N_11641);
xnor U19211 (N_19211,N_10291,N_13970);
nor U19212 (N_19212,N_10886,N_11883);
or U19213 (N_19213,N_14815,N_11297);
nor U19214 (N_19214,N_12077,N_13283);
or U19215 (N_19215,N_14843,N_10527);
xnor U19216 (N_19216,N_12813,N_14408);
nor U19217 (N_19217,N_13049,N_13126);
or U19218 (N_19218,N_10202,N_13723);
xor U19219 (N_19219,N_13894,N_12652);
nor U19220 (N_19220,N_13643,N_10548);
or U19221 (N_19221,N_11846,N_11948);
or U19222 (N_19222,N_12653,N_14461);
nor U19223 (N_19223,N_13213,N_12976);
or U19224 (N_19224,N_12861,N_10562);
nand U19225 (N_19225,N_13896,N_12021);
nand U19226 (N_19226,N_10928,N_11180);
nor U19227 (N_19227,N_13093,N_11124);
xor U19228 (N_19228,N_13844,N_11505);
and U19229 (N_19229,N_12487,N_13827);
xor U19230 (N_19230,N_14017,N_13005);
nand U19231 (N_19231,N_12549,N_13627);
nand U19232 (N_19232,N_10785,N_10612);
xnor U19233 (N_19233,N_14102,N_12977);
xor U19234 (N_19234,N_11701,N_12428);
xor U19235 (N_19235,N_14333,N_12900);
and U19236 (N_19236,N_10558,N_12823);
and U19237 (N_19237,N_10755,N_13754);
or U19238 (N_19238,N_12873,N_13949);
nand U19239 (N_19239,N_10305,N_13101);
nor U19240 (N_19240,N_13060,N_13243);
and U19241 (N_19241,N_14601,N_10734);
nor U19242 (N_19242,N_11041,N_14816);
or U19243 (N_19243,N_10500,N_14782);
and U19244 (N_19244,N_12302,N_13381);
nor U19245 (N_19245,N_10210,N_13739);
nand U19246 (N_19246,N_11829,N_14187);
xor U19247 (N_19247,N_11556,N_12805);
nor U19248 (N_19248,N_14678,N_11593);
or U19249 (N_19249,N_10883,N_14247);
or U19250 (N_19250,N_11005,N_14368);
nand U19251 (N_19251,N_11001,N_14231);
and U19252 (N_19252,N_14111,N_14670);
xor U19253 (N_19253,N_12750,N_14180);
xor U19254 (N_19254,N_13545,N_11729);
and U19255 (N_19255,N_10079,N_10210);
and U19256 (N_19256,N_10257,N_13709);
or U19257 (N_19257,N_10555,N_10092);
nor U19258 (N_19258,N_10464,N_10291);
and U19259 (N_19259,N_14433,N_12796);
nand U19260 (N_19260,N_11468,N_12824);
and U19261 (N_19261,N_12926,N_14313);
or U19262 (N_19262,N_14317,N_10469);
xnor U19263 (N_19263,N_10177,N_11085);
or U19264 (N_19264,N_13165,N_13524);
nor U19265 (N_19265,N_14713,N_11314);
and U19266 (N_19266,N_12680,N_14523);
or U19267 (N_19267,N_13627,N_10963);
xor U19268 (N_19268,N_14838,N_10524);
and U19269 (N_19269,N_12867,N_10506);
and U19270 (N_19270,N_12819,N_10699);
and U19271 (N_19271,N_11786,N_10332);
or U19272 (N_19272,N_13753,N_10158);
or U19273 (N_19273,N_14624,N_14679);
nor U19274 (N_19274,N_14366,N_13137);
nand U19275 (N_19275,N_14963,N_13252);
nand U19276 (N_19276,N_14200,N_11623);
nand U19277 (N_19277,N_14906,N_13074);
nand U19278 (N_19278,N_12715,N_10714);
xnor U19279 (N_19279,N_12695,N_14710);
nand U19280 (N_19280,N_10393,N_11539);
or U19281 (N_19281,N_14821,N_10379);
and U19282 (N_19282,N_14245,N_10218);
xor U19283 (N_19283,N_13640,N_14786);
xnor U19284 (N_19284,N_12452,N_13916);
or U19285 (N_19285,N_14498,N_14358);
or U19286 (N_19286,N_10395,N_13722);
nor U19287 (N_19287,N_12266,N_11029);
and U19288 (N_19288,N_10633,N_14687);
xnor U19289 (N_19289,N_11059,N_12075);
xnor U19290 (N_19290,N_12331,N_14812);
nor U19291 (N_19291,N_13372,N_10330);
nor U19292 (N_19292,N_13775,N_11821);
nand U19293 (N_19293,N_12347,N_14528);
nand U19294 (N_19294,N_14290,N_12931);
xnor U19295 (N_19295,N_11824,N_10587);
or U19296 (N_19296,N_14024,N_11356);
nand U19297 (N_19297,N_11125,N_11794);
xor U19298 (N_19298,N_10453,N_10148);
nand U19299 (N_19299,N_13472,N_10770);
nor U19300 (N_19300,N_12258,N_11673);
xor U19301 (N_19301,N_11924,N_11548);
and U19302 (N_19302,N_14228,N_14406);
and U19303 (N_19303,N_14535,N_10013);
xnor U19304 (N_19304,N_11458,N_13649);
nand U19305 (N_19305,N_13049,N_12020);
nand U19306 (N_19306,N_13800,N_11731);
or U19307 (N_19307,N_11353,N_10562);
xnor U19308 (N_19308,N_13210,N_14476);
and U19309 (N_19309,N_10221,N_10530);
nor U19310 (N_19310,N_12712,N_12819);
nor U19311 (N_19311,N_10622,N_13424);
xnor U19312 (N_19312,N_14424,N_10439);
and U19313 (N_19313,N_12382,N_13874);
nor U19314 (N_19314,N_14203,N_12197);
nor U19315 (N_19315,N_13086,N_11068);
and U19316 (N_19316,N_14180,N_11071);
xor U19317 (N_19317,N_11121,N_14208);
nor U19318 (N_19318,N_11897,N_11722);
and U19319 (N_19319,N_12068,N_12146);
xor U19320 (N_19320,N_14584,N_11191);
and U19321 (N_19321,N_13460,N_10271);
or U19322 (N_19322,N_13653,N_12139);
and U19323 (N_19323,N_11101,N_11741);
nand U19324 (N_19324,N_12865,N_13162);
nor U19325 (N_19325,N_14603,N_10123);
xor U19326 (N_19326,N_11832,N_13035);
xnor U19327 (N_19327,N_12555,N_10887);
or U19328 (N_19328,N_10474,N_13378);
xnor U19329 (N_19329,N_13140,N_13494);
nand U19330 (N_19330,N_13867,N_10034);
nor U19331 (N_19331,N_14281,N_10027);
nor U19332 (N_19332,N_12599,N_12275);
nor U19333 (N_19333,N_13743,N_11141);
xnor U19334 (N_19334,N_13421,N_13714);
nand U19335 (N_19335,N_11311,N_14142);
or U19336 (N_19336,N_13364,N_14708);
or U19337 (N_19337,N_13472,N_14450);
and U19338 (N_19338,N_10769,N_14308);
nand U19339 (N_19339,N_13972,N_12561);
or U19340 (N_19340,N_11662,N_11908);
xnor U19341 (N_19341,N_11382,N_11669);
xor U19342 (N_19342,N_12198,N_14386);
or U19343 (N_19343,N_11298,N_13568);
and U19344 (N_19344,N_13255,N_12389);
or U19345 (N_19345,N_11961,N_13793);
xor U19346 (N_19346,N_11958,N_14090);
nand U19347 (N_19347,N_12324,N_12076);
or U19348 (N_19348,N_10081,N_10515);
or U19349 (N_19349,N_13217,N_12803);
nor U19350 (N_19350,N_12625,N_11212);
or U19351 (N_19351,N_11937,N_13519);
xnor U19352 (N_19352,N_10797,N_14260);
nand U19353 (N_19353,N_10577,N_11903);
nor U19354 (N_19354,N_14630,N_13608);
xor U19355 (N_19355,N_11882,N_11001);
nor U19356 (N_19356,N_12021,N_11331);
or U19357 (N_19357,N_14940,N_13530);
xor U19358 (N_19358,N_12527,N_11931);
or U19359 (N_19359,N_12044,N_11424);
or U19360 (N_19360,N_13584,N_14512);
nand U19361 (N_19361,N_12293,N_14976);
and U19362 (N_19362,N_10661,N_12609);
or U19363 (N_19363,N_11657,N_10865);
and U19364 (N_19364,N_10149,N_10771);
xnor U19365 (N_19365,N_10759,N_13921);
and U19366 (N_19366,N_13696,N_13376);
nand U19367 (N_19367,N_11764,N_14801);
xnor U19368 (N_19368,N_12376,N_12504);
xor U19369 (N_19369,N_12861,N_13921);
nor U19370 (N_19370,N_10024,N_11911);
nand U19371 (N_19371,N_12259,N_12037);
nor U19372 (N_19372,N_13343,N_13123);
nor U19373 (N_19373,N_12021,N_11586);
nor U19374 (N_19374,N_13642,N_12082);
and U19375 (N_19375,N_12355,N_10155);
nand U19376 (N_19376,N_14871,N_11767);
xor U19377 (N_19377,N_10342,N_12543);
and U19378 (N_19378,N_14868,N_10117);
xor U19379 (N_19379,N_12597,N_11669);
nand U19380 (N_19380,N_10154,N_11023);
or U19381 (N_19381,N_13127,N_13081);
nor U19382 (N_19382,N_10922,N_12370);
xnor U19383 (N_19383,N_12842,N_11034);
and U19384 (N_19384,N_10652,N_12084);
nor U19385 (N_19385,N_14872,N_12207);
nand U19386 (N_19386,N_12061,N_13965);
xnor U19387 (N_19387,N_10168,N_14071);
nor U19388 (N_19388,N_11132,N_12809);
and U19389 (N_19389,N_13597,N_12086);
nand U19390 (N_19390,N_11692,N_10031);
xor U19391 (N_19391,N_13167,N_14438);
nor U19392 (N_19392,N_10042,N_14449);
xor U19393 (N_19393,N_13997,N_11496);
nand U19394 (N_19394,N_10156,N_14748);
nor U19395 (N_19395,N_11987,N_11187);
and U19396 (N_19396,N_10598,N_10366);
xnor U19397 (N_19397,N_11484,N_14185);
and U19398 (N_19398,N_11066,N_12181);
nor U19399 (N_19399,N_10853,N_10332);
xor U19400 (N_19400,N_14756,N_14574);
nand U19401 (N_19401,N_10207,N_13725);
nand U19402 (N_19402,N_11719,N_14578);
xnor U19403 (N_19403,N_14160,N_11653);
and U19404 (N_19404,N_14293,N_10501);
nand U19405 (N_19405,N_11468,N_13772);
or U19406 (N_19406,N_13469,N_10315);
nand U19407 (N_19407,N_14930,N_12463);
and U19408 (N_19408,N_12572,N_10661);
xnor U19409 (N_19409,N_12484,N_11545);
nand U19410 (N_19410,N_11719,N_11011);
nor U19411 (N_19411,N_12622,N_13053);
nand U19412 (N_19412,N_11247,N_13960);
nor U19413 (N_19413,N_13814,N_12547);
or U19414 (N_19414,N_12997,N_13488);
or U19415 (N_19415,N_12521,N_11278);
xor U19416 (N_19416,N_14216,N_10532);
nand U19417 (N_19417,N_13158,N_11741);
or U19418 (N_19418,N_13881,N_14713);
xor U19419 (N_19419,N_12069,N_13944);
nand U19420 (N_19420,N_10415,N_12035);
nand U19421 (N_19421,N_10192,N_14445);
or U19422 (N_19422,N_14863,N_12236);
nor U19423 (N_19423,N_13876,N_13160);
nor U19424 (N_19424,N_10301,N_12125);
or U19425 (N_19425,N_11804,N_11797);
xnor U19426 (N_19426,N_12214,N_10629);
or U19427 (N_19427,N_13802,N_10802);
nand U19428 (N_19428,N_12953,N_12156);
nor U19429 (N_19429,N_12685,N_12156);
and U19430 (N_19430,N_14750,N_10234);
xnor U19431 (N_19431,N_14301,N_13018);
xnor U19432 (N_19432,N_14098,N_12011);
xnor U19433 (N_19433,N_12097,N_14521);
or U19434 (N_19434,N_11794,N_12413);
nor U19435 (N_19435,N_11697,N_14226);
nor U19436 (N_19436,N_13409,N_14819);
or U19437 (N_19437,N_11609,N_12641);
or U19438 (N_19438,N_14801,N_11377);
nand U19439 (N_19439,N_11131,N_11731);
xor U19440 (N_19440,N_12226,N_11675);
or U19441 (N_19441,N_10617,N_14232);
xnor U19442 (N_19442,N_11697,N_12745);
nand U19443 (N_19443,N_12705,N_10114);
xnor U19444 (N_19444,N_12882,N_14105);
nand U19445 (N_19445,N_11711,N_13403);
nand U19446 (N_19446,N_13025,N_14580);
nand U19447 (N_19447,N_11107,N_11611);
and U19448 (N_19448,N_13082,N_13092);
xnor U19449 (N_19449,N_13463,N_13256);
xnor U19450 (N_19450,N_11228,N_10224);
or U19451 (N_19451,N_12823,N_14039);
nor U19452 (N_19452,N_13599,N_10411);
nor U19453 (N_19453,N_13533,N_14413);
or U19454 (N_19454,N_11596,N_11629);
xor U19455 (N_19455,N_10281,N_12940);
xor U19456 (N_19456,N_14957,N_13404);
and U19457 (N_19457,N_11963,N_13775);
nor U19458 (N_19458,N_13258,N_12316);
xor U19459 (N_19459,N_12080,N_10937);
xor U19460 (N_19460,N_14806,N_10951);
nor U19461 (N_19461,N_11541,N_10819);
xnor U19462 (N_19462,N_10214,N_10848);
nor U19463 (N_19463,N_14022,N_11793);
or U19464 (N_19464,N_12264,N_10719);
xor U19465 (N_19465,N_12122,N_14552);
xnor U19466 (N_19466,N_14389,N_13929);
nand U19467 (N_19467,N_10251,N_11757);
nor U19468 (N_19468,N_13593,N_12559);
nor U19469 (N_19469,N_14945,N_12551);
nor U19470 (N_19470,N_12312,N_12635);
and U19471 (N_19471,N_10972,N_12057);
or U19472 (N_19472,N_13075,N_13894);
xnor U19473 (N_19473,N_10482,N_10618);
and U19474 (N_19474,N_11774,N_13711);
nor U19475 (N_19475,N_14747,N_13938);
or U19476 (N_19476,N_14581,N_13515);
and U19477 (N_19477,N_10533,N_10650);
nand U19478 (N_19478,N_11522,N_10658);
nand U19479 (N_19479,N_14199,N_12044);
or U19480 (N_19480,N_11380,N_11652);
xnor U19481 (N_19481,N_14335,N_13153);
xnor U19482 (N_19482,N_14148,N_13923);
nor U19483 (N_19483,N_10305,N_12063);
or U19484 (N_19484,N_14651,N_11532);
and U19485 (N_19485,N_11101,N_12099);
and U19486 (N_19486,N_14731,N_14850);
and U19487 (N_19487,N_10777,N_11259);
xor U19488 (N_19488,N_14233,N_14295);
and U19489 (N_19489,N_13193,N_12781);
or U19490 (N_19490,N_10192,N_11335);
nand U19491 (N_19491,N_10835,N_14047);
nor U19492 (N_19492,N_11904,N_12372);
and U19493 (N_19493,N_14497,N_10617);
or U19494 (N_19494,N_10888,N_10915);
or U19495 (N_19495,N_14549,N_12972);
nor U19496 (N_19496,N_10723,N_13613);
xnor U19497 (N_19497,N_14997,N_13868);
or U19498 (N_19498,N_11628,N_13339);
xor U19499 (N_19499,N_13706,N_10223);
nor U19500 (N_19500,N_14714,N_12381);
xor U19501 (N_19501,N_14301,N_12541);
nor U19502 (N_19502,N_11051,N_12369);
nand U19503 (N_19503,N_10186,N_14869);
nand U19504 (N_19504,N_11977,N_12632);
or U19505 (N_19505,N_13509,N_11169);
or U19506 (N_19506,N_12753,N_14710);
or U19507 (N_19507,N_11749,N_13071);
or U19508 (N_19508,N_12203,N_11304);
and U19509 (N_19509,N_11538,N_10569);
and U19510 (N_19510,N_12028,N_12598);
nand U19511 (N_19511,N_10810,N_11040);
or U19512 (N_19512,N_12388,N_10657);
or U19513 (N_19513,N_14452,N_12524);
and U19514 (N_19514,N_12742,N_10983);
and U19515 (N_19515,N_14975,N_12987);
nand U19516 (N_19516,N_11389,N_13093);
nor U19517 (N_19517,N_11506,N_10089);
nor U19518 (N_19518,N_12014,N_14321);
and U19519 (N_19519,N_14789,N_12293);
and U19520 (N_19520,N_13954,N_13355);
or U19521 (N_19521,N_14034,N_10922);
and U19522 (N_19522,N_10375,N_11968);
xnor U19523 (N_19523,N_11676,N_11542);
nor U19524 (N_19524,N_11460,N_14968);
or U19525 (N_19525,N_10812,N_13902);
xor U19526 (N_19526,N_10787,N_14730);
or U19527 (N_19527,N_10274,N_14204);
nand U19528 (N_19528,N_11731,N_11529);
nor U19529 (N_19529,N_12598,N_11046);
nor U19530 (N_19530,N_10522,N_11736);
or U19531 (N_19531,N_14513,N_12380);
and U19532 (N_19532,N_10643,N_13181);
or U19533 (N_19533,N_10180,N_14100);
or U19534 (N_19534,N_11787,N_10235);
xnor U19535 (N_19535,N_10198,N_14290);
xor U19536 (N_19536,N_10292,N_11533);
nand U19537 (N_19537,N_10384,N_14763);
and U19538 (N_19538,N_13811,N_11899);
nor U19539 (N_19539,N_10103,N_10013);
xnor U19540 (N_19540,N_11334,N_10849);
xnor U19541 (N_19541,N_13568,N_10855);
nand U19542 (N_19542,N_10153,N_10946);
nand U19543 (N_19543,N_13348,N_11776);
nor U19544 (N_19544,N_13133,N_12554);
and U19545 (N_19545,N_14911,N_13768);
and U19546 (N_19546,N_13039,N_11004);
or U19547 (N_19547,N_12679,N_11771);
and U19548 (N_19548,N_14645,N_14686);
nand U19549 (N_19549,N_12459,N_11012);
and U19550 (N_19550,N_13343,N_12738);
xnor U19551 (N_19551,N_12394,N_12475);
nor U19552 (N_19552,N_10806,N_10766);
or U19553 (N_19553,N_10521,N_13943);
nand U19554 (N_19554,N_10938,N_11815);
and U19555 (N_19555,N_11056,N_10308);
nor U19556 (N_19556,N_13941,N_13767);
xnor U19557 (N_19557,N_12426,N_14486);
and U19558 (N_19558,N_12880,N_10161);
and U19559 (N_19559,N_13006,N_10609);
nand U19560 (N_19560,N_13256,N_12802);
nand U19561 (N_19561,N_10981,N_10779);
and U19562 (N_19562,N_10964,N_13324);
xnor U19563 (N_19563,N_14377,N_11606);
or U19564 (N_19564,N_11560,N_14738);
xor U19565 (N_19565,N_12545,N_10664);
and U19566 (N_19566,N_13955,N_10390);
or U19567 (N_19567,N_11845,N_10477);
xor U19568 (N_19568,N_10241,N_12432);
nor U19569 (N_19569,N_10990,N_12534);
nand U19570 (N_19570,N_11534,N_12158);
and U19571 (N_19571,N_13801,N_11296);
and U19572 (N_19572,N_14607,N_11290);
nand U19573 (N_19573,N_14965,N_13996);
xnor U19574 (N_19574,N_14565,N_10990);
nor U19575 (N_19575,N_14900,N_12675);
and U19576 (N_19576,N_10360,N_14801);
or U19577 (N_19577,N_14769,N_12645);
nand U19578 (N_19578,N_11955,N_14615);
and U19579 (N_19579,N_12887,N_10486);
or U19580 (N_19580,N_12523,N_12783);
and U19581 (N_19581,N_14618,N_10506);
or U19582 (N_19582,N_11731,N_11498);
nand U19583 (N_19583,N_13754,N_11498);
xor U19584 (N_19584,N_13970,N_12001);
and U19585 (N_19585,N_10778,N_10049);
and U19586 (N_19586,N_13004,N_12504);
nand U19587 (N_19587,N_11815,N_10976);
or U19588 (N_19588,N_14714,N_10155);
and U19589 (N_19589,N_11558,N_13190);
nor U19590 (N_19590,N_12996,N_13425);
nand U19591 (N_19591,N_14770,N_12765);
nor U19592 (N_19592,N_13384,N_10504);
and U19593 (N_19593,N_13615,N_10249);
and U19594 (N_19594,N_12473,N_10607);
and U19595 (N_19595,N_11958,N_14467);
and U19596 (N_19596,N_11765,N_11713);
and U19597 (N_19597,N_13049,N_12226);
xnor U19598 (N_19598,N_14929,N_11626);
nor U19599 (N_19599,N_10911,N_11111);
and U19600 (N_19600,N_14639,N_13276);
nand U19601 (N_19601,N_13252,N_10143);
nand U19602 (N_19602,N_10122,N_12410);
xnor U19603 (N_19603,N_11539,N_10560);
nor U19604 (N_19604,N_11028,N_14371);
nand U19605 (N_19605,N_14498,N_11089);
xnor U19606 (N_19606,N_12345,N_12930);
and U19607 (N_19607,N_13569,N_12674);
or U19608 (N_19608,N_14357,N_10491);
nand U19609 (N_19609,N_10252,N_10170);
nand U19610 (N_19610,N_14173,N_13803);
xnor U19611 (N_19611,N_13434,N_14412);
nor U19612 (N_19612,N_12365,N_11578);
nor U19613 (N_19613,N_12077,N_13921);
and U19614 (N_19614,N_11425,N_14985);
nand U19615 (N_19615,N_13710,N_11233);
xor U19616 (N_19616,N_14379,N_14792);
and U19617 (N_19617,N_12459,N_13216);
nor U19618 (N_19618,N_12682,N_13138);
or U19619 (N_19619,N_13386,N_13628);
nand U19620 (N_19620,N_14452,N_11803);
xor U19621 (N_19621,N_12291,N_11359);
and U19622 (N_19622,N_14588,N_14498);
nor U19623 (N_19623,N_14557,N_13952);
xor U19624 (N_19624,N_11953,N_12450);
and U19625 (N_19625,N_14468,N_10131);
and U19626 (N_19626,N_12774,N_14420);
or U19627 (N_19627,N_10827,N_14879);
nand U19628 (N_19628,N_12854,N_10846);
or U19629 (N_19629,N_11697,N_14674);
nand U19630 (N_19630,N_13711,N_11532);
or U19631 (N_19631,N_13792,N_10830);
xor U19632 (N_19632,N_11883,N_14647);
xnor U19633 (N_19633,N_10522,N_12381);
and U19634 (N_19634,N_13939,N_13339);
or U19635 (N_19635,N_11631,N_11940);
xnor U19636 (N_19636,N_11797,N_11279);
and U19637 (N_19637,N_12317,N_13771);
and U19638 (N_19638,N_10360,N_10025);
nand U19639 (N_19639,N_10941,N_11377);
and U19640 (N_19640,N_11432,N_14742);
and U19641 (N_19641,N_12548,N_12727);
nand U19642 (N_19642,N_10736,N_14891);
and U19643 (N_19643,N_10797,N_13989);
nand U19644 (N_19644,N_10017,N_13235);
xnor U19645 (N_19645,N_12287,N_13543);
nor U19646 (N_19646,N_11758,N_14213);
nand U19647 (N_19647,N_14567,N_13511);
nor U19648 (N_19648,N_12696,N_14674);
nand U19649 (N_19649,N_10787,N_12599);
nand U19650 (N_19650,N_13281,N_10236);
nand U19651 (N_19651,N_13880,N_11725);
nor U19652 (N_19652,N_11292,N_12758);
and U19653 (N_19653,N_12757,N_11415);
xor U19654 (N_19654,N_11157,N_10291);
or U19655 (N_19655,N_12088,N_12271);
nor U19656 (N_19656,N_10226,N_10111);
xnor U19657 (N_19657,N_13351,N_12032);
nor U19658 (N_19658,N_13264,N_13037);
or U19659 (N_19659,N_13127,N_13004);
xnor U19660 (N_19660,N_10380,N_12271);
nor U19661 (N_19661,N_14234,N_12447);
xnor U19662 (N_19662,N_10327,N_12143);
nand U19663 (N_19663,N_12193,N_14985);
nand U19664 (N_19664,N_13324,N_11449);
nor U19665 (N_19665,N_14192,N_12060);
xor U19666 (N_19666,N_13501,N_13173);
xnor U19667 (N_19667,N_13768,N_14257);
nor U19668 (N_19668,N_14079,N_10861);
nand U19669 (N_19669,N_10821,N_11586);
nand U19670 (N_19670,N_12953,N_10193);
and U19671 (N_19671,N_14034,N_10307);
xnor U19672 (N_19672,N_10594,N_13576);
or U19673 (N_19673,N_10133,N_11042);
nand U19674 (N_19674,N_13020,N_14809);
nor U19675 (N_19675,N_10247,N_10752);
or U19676 (N_19676,N_14721,N_12817);
xnor U19677 (N_19677,N_10992,N_11112);
or U19678 (N_19678,N_13755,N_14367);
and U19679 (N_19679,N_13980,N_12342);
nand U19680 (N_19680,N_14681,N_13180);
xor U19681 (N_19681,N_13177,N_12732);
and U19682 (N_19682,N_13946,N_10376);
xnor U19683 (N_19683,N_10190,N_13620);
xnor U19684 (N_19684,N_11385,N_14340);
xnor U19685 (N_19685,N_13163,N_14184);
nor U19686 (N_19686,N_13029,N_11744);
nor U19687 (N_19687,N_14176,N_12404);
nand U19688 (N_19688,N_13411,N_10985);
nand U19689 (N_19689,N_14267,N_13088);
and U19690 (N_19690,N_14747,N_13455);
nand U19691 (N_19691,N_10222,N_11205);
and U19692 (N_19692,N_10309,N_14743);
nor U19693 (N_19693,N_14117,N_12169);
nand U19694 (N_19694,N_14206,N_13676);
nor U19695 (N_19695,N_14182,N_11869);
and U19696 (N_19696,N_12245,N_13955);
or U19697 (N_19697,N_11637,N_14605);
and U19698 (N_19698,N_11959,N_10784);
and U19699 (N_19699,N_12438,N_12706);
nand U19700 (N_19700,N_10458,N_14474);
and U19701 (N_19701,N_14341,N_10726);
or U19702 (N_19702,N_11938,N_11134);
or U19703 (N_19703,N_14543,N_14528);
and U19704 (N_19704,N_11782,N_11773);
nor U19705 (N_19705,N_12874,N_10963);
and U19706 (N_19706,N_11083,N_12805);
xor U19707 (N_19707,N_13452,N_11192);
nand U19708 (N_19708,N_10475,N_13658);
or U19709 (N_19709,N_10389,N_11311);
nand U19710 (N_19710,N_14320,N_10177);
and U19711 (N_19711,N_10903,N_11795);
nor U19712 (N_19712,N_12426,N_13517);
nor U19713 (N_19713,N_10526,N_10839);
nand U19714 (N_19714,N_14639,N_14196);
or U19715 (N_19715,N_12826,N_12852);
nor U19716 (N_19716,N_13284,N_10520);
xnor U19717 (N_19717,N_12052,N_12938);
and U19718 (N_19718,N_11757,N_12167);
and U19719 (N_19719,N_14666,N_10899);
and U19720 (N_19720,N_14327,N_10515);
nand U19721 (N_19721,N_13002,N_12395);
nand U19722 (N_19722,N_12669,N_11743);
nor U19723 (N_19723,N_12563,N_12559);
xor U19724 (N_19724,N_10293,N_10497);
nor U19725 (N_19725,N_11151,N_12534);
xor U19726 (N_19726,N_13381,N_11516);
nor U19727 (N_19727,N_12631,N_10268);
nand U19728 (N_19728,N_14794,N_14988);
nand U19729 (N_19729,N_13133,N_14600);
xor U19730 (N_19730,N_13552,N_12654);
or U19731 (N_19731,N_10642,N_14926);
and U19732 (N_19732,N_12382,N_13170);
nand U19733 (N_19733,N_10154,N_14721);
or U19734 (N_19734,N_14861,N_13529);
nand U19735 (N_19735,N_13378,N_11301);
or U19736 (N_19736,N_13298,N_13934);
nand U19737 (N_19737,N_12758,N_11058);
and U19738 (N_19738,N_11039,N_10887);
and U19739 (N_19739,N_10836,N_14818);
and U19740 (N_19740,N_11993,N_14751);
nor U19741 (N_19741,N_13994,N_11017);
and U19742 (N_19742,N_11626,N_11425);
and U19743 (N_19743,N_14219,N_12466);
nor U19744 (N_19744,N_13563,N_13365);
or U19745 (N_19745,N_14690,N_14089);
or U19746 (N_19746,N_10510,N_11680);
nand U19747 (N_19747,N_14133,N_10020);
xor U19748 (N_19748,N_14511,N_13666);
nand U19749 (N_19749,N_10348,N_14524);
or U19750 (N_19750,N_10592,N_14224);
nand U19751 (N_19751,N_11645,N_14059);
nand U19752 (N_19752,N_13526,N_12356);
nand U19753 (N_19753,N_14463,N_10289);
xnor U19754 (N_19754,N_13996,N_10101);
nand U19755 (N_19755,N_10835,N_12344);
nand U19756 (N_19756,N_13036,N_13606);
xnor U19757 (N_19757,N_10269,N_11983);
or U19758 (N_19758,N_12567,N_13387);
nor U19759 (N_19759,N_12505,N_12720);
nand U19760 (N_19760,N_13886,N_11099);
and U19761 (N_19761,N_13142,N_12447);
and U19762 (N_19762,N_13309,N_10406);
xor U19763 (N_19763,N_12124,N_14829);
xnor U19764 (N_19764,N_11670,N_12655);
nor U19765 (N_19765,N_14641,N_10844);
nor U19766 (N_19766,N_13550,N_13382);
and U19767 (N_19767,N_10587,N_11250);
and U19768 (N_19768,N_10053,N_13597);
or U19769 (N_19769,N_12426,N_14537);
xnor U19770 (N_19770,N_10543,N_10423);
xnor U19771 (N_19771,N_11479,N_14777);
nand U19772 (N_19772,N_10068,N_14601);
and U19773 (N_19773,N_11753,N_11119);
nand U19774 (N_19774,N_10652,N_10293);
and U19775 (N_19775,N_13336,N_10601);
or U19776 (N_19776,N_14253,N_13488);
and U19777 (N_19777,N_14330,N_13359);
xnor U19778 (N_19778,N_12084,N_13727);
nor U19779 (N_19779,N_10996,N_14521);
xnor U19780 (N_19780,N_12584,N_11172);
nor U19781 (N_19781,N_11998,N_13118);
and U19782 (N_19782,N_13198,N_13987);
and U19783 (N_19783,N_14820,N_12313);
nand U19784 (N_19784,N_13890,N_10297);
or U19785 (N_19785,N_14367,N_12779);
xor U19786 (N_19786,N_12241,N_10979);
nand U19787 (N_19787,N_10745,N_10056);
nor U19788 (N_19788,N_11601,N_14393);
or U19789 (N_19789,N_10296,N_13795);
nor U19790 (N_19790,N_12237,N_11877);
nor U19791 (N_19791,N_10067,N_11570);
nand U19792 (N_19792,N_11642,N_14757);
xor U19793 (N_19793,N_11263,N_12750);
and U19794 (N_19794,N_12356,N_14544);
xor U19795 (N_19795,N_13927,N_13854);
nand U19796 (N_19796,N_14810,N_11577);
xnor U19797 (N_19797,N_12463,N_11129);
nor U19798 (N_19798,N_12048,N_12391);
and U19799 (N_19799,N_14845,N_14657);
nand U19800 (N_19800,N_12725,N_13036);
and U19801 (N_19801,N_11325,N_12213);
or U19802 (N_19802,N_10838,N_12801);
or U19803 (N_19803,N_10617,N_14712);
nor U19804 (N_19804,N_12335,N_11895);
or U19805 (N_19805,N_14382,N_10729);
or U19806 (N_19806,N_12124,N_11907);
or U19807 (N_19807,N_13551,N_12382);
xnor U19808 (N_19808,N_11109,N_14103);
and U19809 (N_19809,N_10185,N_10827);
nand U19810 (N_19810,N_10790,N_12905);
or U19811 (N_19811,N_11462,N_12184);
or U19812 (N_19812,N_13432,N_13501);
or U19813 (N_19813,N_12251,N_14027);
xnor U19814 (N_19814,N_14930,N_13529);
or U19815 (N_19815,N_13586,N_12355);
xor U19816 (N_19816,N_14150,N_12198);
xnor U19817 (N_19817,N_13044,N_13398);
and U19818 (N_19818,N_13019,N_10589);
nand U19819 (N_19819,N_12650,N_12525);
nor U19820 (N_19820,N_11959,N_12360);
xnor U19821 (N_19821,N_11290,N_12448);
xor U19822 (N_19822,N_12731,N_10597);
and U19823 (N_19823,N_12481,N_11038);
or U19824 (N_19824,N_11275,N_10952);
nand U19825 (N_19825,N_11478,N_10092);
and U19826 (N_19826,N_10934,N_10300);
or U19827 (N_19827,N_12691,N_14406);
xor U19828 (N_19828,N_14866,N_10367);
nand U19829 (N_19829,N_14077,N_13385);
and U19830 (N_19830,N_12206,N_10517);
xnor U19831 (N_19831,N_12256,N_14979);
nand U19832 (N_19832,N_13907,N_12373);
nand U19833 (N_19833,N_14641,N_13185);
and U19834 (N_19834,N_14288,N_12891);
xor U19835 (N_19835,N_14710,N_11296);
nand U19836 (N_19836,N_14318,N_10080);
or U19837 (N_19837,N_13448,N_11609);
xnor U19838 (N_19838,N_12923,N_11313);
nand U19839 (N_19839,N_10509,N_13185);
xor U19840 (N_19840,N_13906,N_11767);
nor U19841 (N_19841,N_12107,N_12621);
or U19842 (N_19842,N_14208,N_12128);
nor U19843 (N_19843,N_13532,N_10537);
xor U19844 (N_19844,N_12732,N_14672);
and U19845 (N_19845,N_12782,N_10531);
nand U19846 (N_19846,N_13684,N_12460);
nand U19847 (N_19847,N_14891,N_13841);
nand U19848 (N_19848,N_10273,N_11137);
xnor U19849 (N_19849,N_12086,N_12428);
nor U19850 (N_19850,N_11224,N_13543);
nand U19851 (N_19851,N_14745,N_13895);
or U19852 (N_19852,N_10687,N_10697);
or U19853 (N_19853,N_13123,N_14027);
xnor U19854 (N_19854,N_11778,N_13162);
nor U19855 (N_19855,N_12545,N_11634);
nor U19856 (N_19856,N_10071,N_13511);
nand U19857 (N_19857,N_10128,N_11973);
or U19858 (N_19858,N_13967,N_10201);
nand U19859 (N_19859,N_10662,N_11171);
xnor U19860 (N_19860,N_12563,N_12185);
xor U19861 (N_19861,N_14886,N_13897);
nand U19862 (N_19862,N_11268,N_12977);
xnor U19863 (N_19863,N_12931,N_13045);
xor U19864 (N_19864,N_13368,N_12638);
or U19865 (N_19865,N_10871,N_13040);
xor U19866 (N_19866,N_14437,N_11278);
or U19867 (N_19867,N_13465,N_13282);
nor U19868 (N_19868,N_14358,N_12564);
nor U19869 (N_19869,N_12515,N_10025);
nand U19870 (N_19870,N_13895,N_12319);
nand U19871 (N_19871,N_13739,N_13290);
and U19872 (N_19872,N_12833,N_13025);
or U19873 (N_19873,N_10624,N_12772);
or U19874 (N_19874,N_13068,N_14404);
or U19875 (N_19875,N_11434,N_10529);
xnor U19876 (N_19876,N_14801,N_13173);
and U19877 (N_19877,N_14026,N_14769);
nand U19878 (N_19878,N_12509,N_11328);
and U19879 (N_19879,N_12596,N_10866);
nand U19880 (N_19880,N_13205,N_10140);
or U19881 (N_19881,N_11629,N_13798);
xor U19882 (N_19882,N_12155,N_10750);
or U19883 (N_19883,N_14961,N_13301);
nor U19884 (N_19884,N_14813,N_10012);
and U19885 (N_19885,N_12358,N_11527);
or U19886 (N_19886,N_12243,N_11095);
nand U19887 (N_19887,N_11472,N_13607);
or U19888 (N_19888,N_10313,N_10566);
xnor U19889 (N_19889,N_11366,N_12825);
or U19890 (N_19890,N_12895,N_14974);
xnor U19891 (N_19891,N_10933,N_12800);
and U19892 (N_19892,N_14894,N_13573);
or U19893 (N_19893,N_10736,N_14452);
xnor U19894 (N_19894,N_12316,N_11097);
nand U19895 (N_19895,N_11136,N_14805);
or U19896 (N_19896,N_13378,N_13281);
xnor U19897 (N_19897,N_14876,N_12643);
or U19898 (N_19898,N_12036,N_12600);
or U19899 (N_19899,N_11952,N_12562);
nand U19900 (N_19900,N_12098,N_12379);
nand U19901 (N_19901,N_12048,N_14118);
or U19902 (N_19902,N_14879,N_10669);
and U19903 (N_19903,N_11359,N_10359);
nor U19904 (N_19904,N_10031,N_11901);
xor U19905 (N_19905,N_12742,N_14493);
nor U19906 (N_19906,N_14576,N_14008);
nor U19907 (N_19907,N_11229,N_13559);
and U19908 (N_19908,N_11761,N_14132);
and U19909 (N_19909,N_14180,N_11719);
nand U19910 (N_19910,N_13569,N_12468);
or U19911 (N_19911,N_12335,N_14224);
xnor U19912 (N_19912,N_14479,N_11259);
xor U19913 (N_19913,N_13850,N_13785);
xnor U19914 (N_19914,N_13637,N_13211);
xnor U19915 (N_19915,N_13650,N_11255);
or U19916 (N_19916,N_14387,N_12996);
nand U19917 (N_19917,N_14673,N_14842);
and U19918 (N_19918,N_12050,N_12790);
nand U19919 (N_19919,N_11942,N_10578);
xor U19920 (N_19920,N_11545,N_12751);
and U19921 (N_19921,N_14388,N_13965);
or U19922 (N_19922,N_13753,N_12628);
or U19923 (N_19923,N_13941,N_12463);
or U19924 (N_19924,N_10367,N_13481);
nor U19925 (N_19925,N_14594,N_10091);
and U19926 (N_19926,N_14103,N_10040);
nand U19927 (N_19927,N_12030,N_12897);
nor U19928 (N_19928,N_11102,N_10053);
nor U19929 (N_19929,N_11472,N_10230);
and U19930 (N_19930,N_14610,N_14358);
nand U19931 (N_19931,N_14679,N_10331);
or U19932 (N_19932,N_11016,N_11212);
or U19933 (N_19933,N_10947,N_12645);
xor U19934 (N_19934,N_14970,N_13235);
or U19935 (N_19935,N_14811,N_14560);
and U19936 (N_19936,N_14280,N_10224);
nand U19937 (N_19937,N_12166,N_11935);
nor U19938 (N_19938,N_13636,N_13529);
nor U19939 (N_19939,N_12307,N_11810);
xnor U19940 (N_19940,N_13925,N_12516);
or U19941 (N_19941,N_13221,N_11588);
or U19942 (N_19942,N_14123,N_11003);
nand U19943 (N_19943,N_12576,N_14006);
and U19944 (N_19944,N_10027,N_14327);
xor U19945 (N_19945,N_14400,N_13380);
nand U19946 (N_19946,N_12092,N_10488);
xnor U19947 (N_19947,N_10081,N_10349);
xnor U19948 (N_19948,N_10401,N_12858);
nand U19949 (N_19949,N_10393,N_14254);
xnor U19950 (N_19950,N_11553,N_11537);
xnor U19951 (N_19951,N_14627,N_11703);
nand U19952 (N_19952,N_14953,N_13518);
or U19953 (N_19953,N_12117,N_10793);
and U19954 (N_19954,N_14219,N_13506);
nor U19955 (N_19955,N_12982,N_14270);
and U19956 (N_19956,N_11930,N_14394);
nand U19957 (N_19957,N_14049,N_11696);
nor U19958 (N_19958,N_10904,N_12077);
nor U19959 (N_19959,N_10427,N_12741);
nand U19960 (N_19960,N_13745,N_13486);
xor U19961 (N_19961,N_10109,N_11280);
or U19962 (N_19962,N_11297,N_14551);
nand U19963 (N_19963,N_11796,N_14256);
and U19964 (N_19964,N_12017,N_10259);
nand U19965 (N_19965,N_13631,N_11729);
or U19966 (N_19966,N_12664,N_10486);
or U19967 (N_19967,N_12175,N_10074);
xnor U19968 (N_19968,N_10499,N_13053);
and U19969 (N_19969,N_11129,N_13620);
nand U19970 (N_19970,N_13262,N_10430);
and U19971 (N_19971,N_11419,N_12569);
nand U19972 (N_19972,N_13918,N_11089);
nor U19973 (N_19973,N_14268,N_10512);
nand U19974 (N_19974,N_12664,N_11924);
or U19975 (N_19975,N_13807,N_12666);
nor U19976 (N_19976,N_12956,N_12025);
and U19977 (N_19977,N_13017,N_12693);
nand U19978 (N_19978,N_13402,N_12832);
nor U19979 (N_19979,N_10353,N_11523);
xor U19980 (N_19980,N_11648,N_13270);
nand U19981 (N_19981,N_12592,N_10646);
xnor U19982 (N_19982,N_13942,N_13464);
xnor U19983 (N_19983,N_14540,N_13699);
nand U19984 (N_19984,N_10139,N_12076);
nor U19985 (N_19985,N_13776,N_13112);
xor U19986 (N_19986,N_11524,N_14807);
or U19987 (N_19987,N_13084,N_13965);
and U19988 (N_19988,N_13971,N_14826);
xor U19989 (N_19989,N_13628,N_10018);
nand U19990 (N_19990,N_14474,N_13706);
and U19991 (N_19991,N_10515,N_10750);
xnor U19992 (N_19992,N_11680,N_12655);
nand U19993 (N_19993,N_13021,N_10764);
xor U19994 (N_19994,N_11413,N_12059);
or U19995 (N_19995,N_11557,N_10989);
or U19996 (N_19996,N_10585,N_10074);
nand U19997 (N_19997,N_12464,N_12662);
or U19998 (N_19998,N_11828,N_13647);
nand U19999 (N_19999,N_10790,N_11277);
or UO_0 (O_0,N_15043,N_19871);
xor UO_1 (O_1,N_17823,N_18976);
nor UO_2 (O_2,N_17404,N_15766);
nand UO_3 (O_3,N_17445,N_15324);
and UO_4 (O_4,N_16814,N_18679);
nor UO_5 (O_5,N_16662,N_17938);
nand UO_6 (O_6,N_18838,N_15177);
and UO_7 (O_7,N_18506,N_16382);
and UO_8 (O_8,N_19321,N_18297);
nor UO_9 (O_9,N_16043,N_18373);
nor UO_10 (O_10,N_19065,N_18897);
or UO_11 (O_11,N_17350,N_19406);
and UO_12 (O_12,N_18889,N_15742);
nand UO_13 (O_13,N_19339,N_16848);
and UO_14 (O_14,N_18943,N_16718);
or UO_15 (O_15,N_15107,N_19240);
nor UO_16 (O_16,N_19060,N_19137);
and UO_17 (O_17,N_17164,N_16455);
nor UO_18 (O_18,N_17528,N_19470);
xor UO_19 (O_19,N_16408,N_17692);
or UO_20 (O_20,N_17902,N_16060);
or UO_21 (O_21,N_19216,N_17691);
nor UO_22 (O_22,N_18665,N_16216);
and UO_23 (O_23,N_15501,N_18763);
and UO_24 (O_24,N_16670,N_19664);
nor UO_25 (O_25,N_17503,N_18787);
nand UO_26 (O_26,N_16643,N_18415);
nand UO_27 (O_27,N_18696,N_16011);
xnor UO_28 (O_28,N_16858,N_17578);
or UO_29 (O_29,N_18625,N_17185);
or UO_30 (O_30,N_15607,N_16983);
or UO_31 (O_31,N_17473,N_18132);
xnor UO_32 (O_32,N_15420,N_15235);
nor UO_33 (O_33,N_17270,N_16118);
and UO_34 (O_34,N_17282,N_19688);
xnor UO_35 (O_35,N_18084,N_19064);
or UO_36 (O_36,N_17737,N_16477);
xnor UO_37 (O_37,N_16017,N_16155);
nor UO_38 (O_38,N_19785,N_15091);
or UO_39 (O_39,N_15755,N_18443);
nor UO_40 (O_40,N_15751,N_17640);
and UO_41 (O_41,N_15106,N_17957);
and UO_42 (O_42,N_16990,N_16184);
and UO_43 (O_43,N_18194,N_15659);
and UO_44 (O_44,N_15348,N_19002);
nor UO_45 (O_45,N_15879,N_15977);
xnor UO_46 (O_46,N_19952,N_19887);
nor UO_47 (O_47,N_16215,N_17762);
xor UO_48 (O_48,N_18877,N_19897);
nand UO_49 (O_49,N_15479,N_18395);
xor UO_50 (O_50,N_18796,N_19028);
xor UO_51 (O_51,N_17620,N_19295);
nand UO_52 (O_52,N_18384,N_15374);
and UO_53 (O_53,N_18997,N_16732);
xor UO_54 (O_54,N_19232,N_18706);
or UO_55 (O_55,N_18691,N_15908);
xnor UO_56 (O_56,N_17796,N_16943);
nand UO_57 (O_57,N_19415,N_17644);
nor UO_58 (O_58,N_16225,N_16575);
and UO_59 (O_59,N_19373,N_15567);
nand UO_60 (O_60,N_15138,N_18659);
nand UO_61 (O_61,N_18145,N_17932);
nor UO_62 (O_62,N_18830,N_19241);
or UO_63 (O_63,N_15404,N_16321);
nand UO_64 (O_64,N_15490,N_16931);
or UO_65 (O_65,N_18528,N_19181);
xor UO_66 (O_66,N_15108,N_18870);
and UO_67 (O_67,N_15972,N_18001);
xor UO_68 (O_68,N_16545,N_15475);
and UO_69 (O_69,N_18324,N_19884);
nor UO_70 (O_70,N_18039,N_17713);
or UO_71 (O_71,N_17304,N_18657);
xnor UO_72 (O_72,N_19626,N_15889);
nor UO_73 (O_73,N_15132,N_17968);
nor UO_74 (O_74,N_17712,N_19336);
nor UO_75 (O_75,N_17276,N_17061);
nand UO_76 (O_76,N_19507,N_15485);
and UO_77 (O_77,N_17348,N_15099);
nand UO_78 (O_78,N_16818,N_18173);
or UO_79 (O_79,N_16022,N_17341);
and UO_80 (O_80,N_16507,N_17724);
and UO_81 (O_81,N_18111,N_17857);
nor UO_82 (O_82,N_17098,N_19213);
and UO_83 (O_83,N_18744,N_15805);
and UO_84 (O_84,N_16890,N_15684);
xnor UO_85 (O_85,N_18177,N_18087);
and UO_86 (O_86,N_15537,N_17891);
nor UO_87 (O_87,N_19997,N_17030);
or UO_88 (O_88,N_19631,N_18697);
and UO_89 (O_89,N_19705,N_16597);
nand UO_90 (O_90,N_16768,N_17336);
xnor UO_91 (O_91,N_15649,N_16682);
nand UO_92 (O_92,N_19079,N_17279);
nor UO_93 (O_93,N_15656,N_17116);
or UO_94 (O_94,N_18263,N_19970);
nor UO_95 (O_95,N_15541,N_16266);
or UO_96 (O_96,N_17438,N_19245);
xor UO_97 (O_97,N_18023,N_16885);
and UO_98 (O_98,N_19751,N_16673);
nand UO_99 (O_99,N_18335,N_18982);
nor UO_100 (O_100,N_15858,N_16008);
nor UO_101 (O_101,N_19671,N_18419);
nand UO_102 (O_102,N_16295,N_18839);
nand UO_103 (O_103,N_15340,N_18467);
nand UO_104 (O_104,N_17395,N_17997);
or UO_105 (O_105,N_19004,N_15583);
and UO_106 (O_106,N_17953,N_17267);
and UO_107 (O_107,N_16456,N_19639);
or UO_108 (O_108,N_15346,N_17260);
nand UO_109 (O_109,N_17666,N_19898);
nand UO_110 (O_110,N_18492,N_16121);
or UO_111 (O_111,N_18961,N_17049);
nor UO_112 (O_112,N_17750,N_17172);
nor UO_113 (O_113,N_17794,N_17660);
or UO_114 (O_114,N_19033,N_16632);
nor UO_115 (O_115,N_19836,N_16573);
nand UO_116 (O_116,N_18368,N_15875);
nand UO_117 (O_117,N_16550,N_15354);
xor UO_118 (O_118,N_18267,N_17767);
and UO_119 (O_119,N_15754,N_16301);
xnor UO_120 (O_120,N_18485,N_16766);
nor UO_121 (O_121,N_19266,N_18481);
xor UO_122 (O_122,N_17777,N_18908);
or UO_123 (O_123,N_19961,N_17947);
and UO_124 (O_124,N_19163,N_18050);
nor UO_125 (O_125,N_17568,N_15104);
and UO_126 (O_126,N_15220,N_18955);
nand UO_127 (O_127,N_15591,N_17018);
xor UO_128 (O_128,N_15998,N_17575);
xnor UO_129 (O_129,N_17887,N_17400);
nand UO_130 (O_130,N_15680,N_18228);
xor UO_131 (O_131,N_19642,N_15312);
xor UO_132 (O_132,N_18888,N_19424);
xnor UO_133 (O_133,N_15196,N_16796);
xnor UO_134 (O_134,N_18719,N_16970);
nor UO_135 (O_135,N_18189,N_19650);
nand UO_136 (O_136,N_19867,N_15605);
nand UO_137 (O_137,N_16448,N_18930);
nor UO_138 (O_138,N_15886,N_19636);
xor UO_139 (O_139,N_16792,N_16171);
and UO_140 (O_140,N_17514,N_16316);
xnor UO_141 (O_141,N_17673,N_19349);
xor UO_142 (O_142,N_15559,N_18262);
xor UO_143 (O_143,N_19472,N_16365);
xnor UO_144 (O_144,N_18074,N_15738);
xor UO_145 (O_145,N_18149,N_15009);
nor UO_146 (O_146,N_18826,N_16248);
or UO_147 (O_147,N_17265,N_18722);
xor UO_148 (O_148,N_15226,N_16275);
xnor UO_149 (O_149,N_15601,N_17844);
and UO_150 (O_150,N_19963,N_17342);
and UO_151 (O_151,N_18531,N_15780);
nand UO_152 (O_152,N_17093,N_15744);
nor UO_153 (O_153,N_18604,N_18660);
nor UO_154 (O_154,N_17380,N_18409);
and UO_155 (O_155,N_16744,N_18899);
xnor UO_156 (O_156,N_16499,N_19802);
nand UO_157 (O_157,N_15065,N_17881);
nor UO_158 (O_158,N_17942,N_18669);
xor UO_159 (O_159,N_16734,N_19300);
and UO_160 (O_160,N_16774,N_17023);
nor UO_161 (O_161,N_18049,N_15895);
or UO_162 (O_162,N_18292,N_17833);
xnor UO_163 (O_163,N_17718,N_16871);
xor UO_164 (O_164,N_16019,N_18342);
and UO_165 (O_165,N_18434,N_17719);
nand UO_166 (O_166,N_17923,N_15381);
or UO_167 (O_167,N_17319,N_15116);
and UO_168 (O_168,N_18025,N_19508);
or UO_169 (O_169,N_19347,N_18986);
nor UO_170 (O_170,N_19196,N_19031);
nor UO_171 (O_171,N_16847,N_17301);
or UO_172 (O_172,N_18234,N_18308);
or UO_173 (O_173,N_17624,N_18754);
or UO_174 (O_174,N_15227,N_15838);
nand UO_175 (O_175,N_19673,N_16797);
nor UO_176 (O_176,N_18024,N_16978);
xor UO_177 (O_177,N_19090,N_16218);
or UO_178 (O_178,N_16917,N_19557);
or UO_179 (O_179,N_18595,N_19037);
nand UO_180 (O_180,N_19178,N_19132);
and UO_181 (O_181,N_18314,N_18542);
nor UO_182 (O_182,N_19640,N_17662);
nor UO_183 (O_183,N_15749,N_16405);
nand UO_184 (O_184,N_18242,N_19681);
and UO_185 (O_185,N_19856,N_17109);
nor UO_186 (O_186,N_16254,N_16029);
nand UO_187 (O_187,N_19513,N_15069);
nand UO_188 (O_188,N_16770,N_18143);
xor UO_189 (O_189,N_15014,N_19238);
xnor UO_190 (O_190,N_19246,N_15512);
xnor UO_191 (O_191,N_16046,N_16447);
xnor UO_192 (O_192,N_16803,N_16502);
or UO_193 (O_193,N_17883,N_18104);
or UO_194 (O_194,N_16541,N_19605);
nor UO_195 (O_195,N_16941,N_18885);
nand UO_196 (O_196,N_15549,N_18585);
and UO_197 (O_197,N_19542,N_19994);
xnor UO_198 (O_198,N_17649,N_19713);
nand UO_199 (O_199,N_18654,N_17476);
and UO_200 (O_200,N_18300,N_19381);
xor UO_201 (O_201,N_18476,N_16199);
nand UO_202 (O_202,N_16051,N_15200);
xnor UO_203 (O_203,N_18695,N_19553);
and UO_204 (O_204,N_19382,N_16981);
nor UO_205 (O_205,N_17999,N_19227);
nand UO_206 (O_206,N_17402,N_17466);
xnor UO_207 (O_207,N_16041,N_19692);
nor UO_208 (O_208,N_19676,N_16416);
nor UO_209 (O_209,N_16389,N_19483);
nand UO_210 (O_210,N_18842,N_16355);
and UO_211 (O_211,N_17884,N_17856);
xnor UO_212 (O_212,N_15570,N_15572);
xnor UO_213 (O_213,N_17309,N_19005);
or UO_214 (O_214,N_15251,N_16304);
nand UO_215 (O_215,N_17378,N_18859);
xor UO_216 (O_216,N_17534,N_19129);
nor UO_217 (O_217,N_17687,N_19094);
nand UO_218 (O_218,N_18969,N_15493);
nor UO_219 (O_219,N_15120,N_15987);
or UO_220 (O_220,N_15364,N_15610);
nand UO_221 (O_221,N_17657,N_15525);
xnor UO_222 (O_222,N_17065,N_16690);
and UO_223 (O_223,N_19799,N_18526);
nor UO_224 (O_224,N_19771,N_17496);
nand UO_225 (O_225,N_18362,N_16778);
xor UO_226 (O_226,N_16212,N_19317);
or UO_227 (O_227,N_19123,N_19127);
and UO_228 (O_228,N_19694,N_17631);
and UO_229 (O_229,N_15521,N_17418);
or UO_230 (O_230,N_16129,N_18709);
nor UO_231 (O_231,N_16532,N_15965);
xor UO_232 (O_232,N_15597,N_15462);
nand UO_233 (O_233,N_18014,N_15049);
or UO_234 (O_234,N_15349,N_16214);
xor UO_235 (O_235,N_19807,N_15458);
and UO_236 (O_236,N_18109,N_17286);
nand UO_237 (O_237,N_17074,N_15784);
xor UO_238 (O_238,N_19988,N_16993);
or UO_239 (O_239,N_18320,N_19541);
and UO_240 (O_240,N_19502,N_18602);
nand UO_241 (O_241,N_15699,N_15870);
and UO_242 (O_242,N_15604,N_18344);
nor UO_243 (O_243,N_16854,N_17416);
or UO_244 (O_244,N_16913,N_18636);
nor UO_245 (O_245,N_17746,N_16303);
nor UO_246 (O_246,N_16546,N_18197);
nor UO_247 (O_247,N_16324,N_16982);
xor UO_248 (O_248,N_17625,N_18821);
and UO_249 (O_249,N_16237,N_15830);
or UO_250 (O_250,N_18091,N_16579);
and UO_251 (O_251,N_15953,N_18609);
or UO_252 (O_252,N_18846,N_15012);
and UO_253 (O_253,N_19461,N_16467);
or UO_254 (O_254,N_17616,N_15826);
nand UO_255 (O_255,N_19383,N_18291);
xnor UO_256 (O_256,N_17310,N_18190);
xor UO_257 (O_257,N_17241,N_17629);
and UO_258 (O_258,N_19904,N_15151);
xnor UO_259 (O_259,N_17236,N_19070);
nor UO_260 (O_260,N_15306,N_15565);
nand UO_261 (O_261,N_15590,N_15001);
nor UO_262 (O_262,N_16264,N_19059);
nor UO_263 (O_263,N_15285,N_18425);
or UO_264 (O_264,N_16974,N_17307);
xnor UO_265 (O_265,N_19560,N_18652);
nand UO_266 (O_266,N_16994,N_18963);
nor UO_267 (O_267,N_15487,N_16535);
xor UO_268 (O_268,N_18587,N_15114);
or UO_269 (O_269,N_18393,N_19779);
or UO_270 (O_270,N_17132,N_19394);
nor UO_271 (O_271,N_16916,N_15534);
and UO_272 (O_272,N_15162,N_19501);
or UO_273 (O_273,N_19545,N_18367);
nor UO_274 (O_274,N_16611,N_16517);
nand UO_275 (O_275,N_17009,N_16182);
nor UO_276 (O_276,N_18203,N_16220);
and UO_277 (O_277,N_19801,N_16281);
nand UO_278 (O_278,N_19220,N_19716);
nor UO_279 (O_279,N_16010,N_19708);
or UO_280 (O_280,N_19253,N_16428);
nor UO_281 (O_281,N_17564,N_16378);
xnor UO_282 (O_282,N_19555,N_15956);
nand UO_283 (O_283,N_16126,N_16213);
xor UO_284 (O_284,N_18155,N_16508);
nand UO_285 (O_285,N_16044,N_18260);
nor UO_286 (O_286,N_15642,N_19320);
nand UO_287 (O_287,N_17269,N_15882);
or UO_288 (O_288,N_19599,N_15667);
xor UO_289 (O_289,N_18707,N_15428);
or UO_290 (O_290,N_19831,N_16644);
nand UO_291 (O_291,N_16671,N_19808);
and UO_292 (O_292,N_18097,N_18243);
xor UO_293 (O_293,N_18977,N_15693);
nand UO_294 (O_294,N_15124,N_19385);
nor UO_295 (O_295,N_18357,N_19927);
nand UO_296 (O_296,N_18293,N_19554);
nor UO_297 (O_297,N_19047,N_19454);
nand UO_298 (O_298,N_17806,N_18555);
xnor UO_299 (O_299,N_15332,N_17707);
and UO_300 (O_300,N_15973,N_17663);
xnor UO_301 (O_301,N_17256,N_15763);
nand UO_302 (O_302,N_17860,N_17144);
and UO_303 (O_303,N_16329,N_18900);
nor UO_304 (O_304,N_19832,N_15382);
and UO_305 (O_305,N_15623,N_19119);
nand UO_306 (O_306,N_15816,N_16158);
nand UO_307 (O_307,N_17391,N_18122);
xor UO_308 (O_308,N_16584,N_15960);
nor UO_309 (O_309,N_17982,N_19355);
or UO_310 (O_310,N_18017,N_17372);
nand UO_311 (O_311,N_17607,N_15403);
or UO_312 (O_312,N_17513,N_17003);
nand UO_313 (O_313,N_17218,N_15711);
nor UO_314 (O_314,N_18804,N_16676);
nor UO_315 (O_315,N_19893,N_19899);
nor UO_316 (O_316,N_19298,N_19931);
and UO_317 (O_317,N_15032,N_18359);
or UO_318 (O_318,N_17990,N_15622);
nand UO_319 (O_319,N_17775,N_19409);
nand UO_320 (O_320,N_18926,N_18829);
xnor UO_321 (O_321,N_16352,N_16819);
nand UO_322 (O_322,N_17863,N_15421);
xor UO_323 (O_323,N_15581,N_19484);
and UO_324 (O_324,N_17216,N_19390);
nor UO_325 (O_325,N_17509,N_17075);
nand UO_326 (O_326,N_18865,N_16484);
or UO_327 (O_327,N_15730,N_19029);
and UO_328 (O_328,N_15773,N_17318);
xnor UO_329 (O_329,N_18245,N_19559);
nor UO_330 (O_330,N_15267,N_19476);
xnor UO_331 (O_331,N_18273,N_16927);
nor UO_332 (O_332,N_15466,N_18752);
or UO_333 (O_333,N_18762,N_17339);
or UO_334 (O_334,N_15734,N_15918);
or UO_335 (O_335,N_19941,N_16536);
nor UO_336 (O_336,N_18034,N_15233);
nand UO_337 (O_337,N_19010,N_19395);
nand UO_338 (O_338,N_17701,N_18910);
nand UO_339 (O_339,N_18389,N_18869);
nand UO_340 (O_340,N_16771,N_18330);
nand UO_341 (O_341,N_19161,N_17014);
or UO_342 (O_342,N_16386,N_16585);
xor UO_343 (O_343,N_18271,N_15914);
nor UO_344 (O_344,N_18855,N_16646);
nand UO_345 (O_345,N_15405,N_16483);
and UO_346 (O_346,N_17428,N_18945);
nor UO_347 (O_347,N_15058,N_17917);
or UO_348 (O_348,N_19932,N_16678);
nand UO_349 (O_349,N_16150,N_16837);
nand UO_350 (O_350,N_19616,N_18550);
xor UO_351 (O_351,N_18252,N_17951);
nand UO_352 (O_352,N_19365,N_17151);
xnor UO_353 (O_353,N_18250,N_18802);
nor UO_354 (O_354,N_18033,N_17804);
nor UO_355 (O_355,N_16251,N_16345);
and UO_356 (O_356,N_16178,N_19099);
nand UO_357 (O_357,N_15414,N_16106);
nand UO_358 (O_358,N_15672,N_16552);
xnor UO_359 (O_359,N_17035,N_19564);
and UO_360 (O_360,N_16967,N_18824);
nand UO_361 (O_361,N_19593,N_19793);
nand UO_362 (O_362,N_18350,N_15216);
xor UO_363 (O_363,N_18503,N_19125);
nor UO_364 (O_364,N_17095,N_17756);
nand UO_365 (O_365,N_18729,N_19619);
xor UO_366 (O_366,N_18529,N_18360);
nor UO_367 (O_367,N_17403,N_18840);
and UO_368 (O_368,N_15315,N_16265);
or UO_369 (O_369,N_16901,N_19297);
nand UO_370 (O_370,N_16424,N_15606);
and UO_371 (O_371,N_16804,N_19140);
nor UO_372 (O_372,N_15673,N_16557);
nand UO_373 (O_373,N_15319,N_19500);
xor UO_374 (O_374,N_16161,N_18572);
or UO_375 (O_375,N_15686,N_18134);
or UO_376 (O_376,N_15300,N_15630);
xor UO_377 (O_377,N_16025,N_17056);
nand UO_378 (O_378,N_18499,N_16465);
or UO_379 (O_379,N_18483,N_16101);
nor UO_380 (O_380,N_17683,N_16273);
and UO_381 (O_381,N_17134,N_16039);
xnor UO_382 (O_382,N_17532,N_16960);
nand UO_383 (O_383,N_17731,N_19209);
xor UO_384 (O_384,N_18430,N_18215);
and UO_385 (O_385,N_16038,N_16294);
and UO_386 (O_386,N_19819,N_18131);
xor UO_387 (O_387,N_18002,N_17803);
nor UO_388 (O_388,N_18450,N_15687);
or UO_389 (O_389,N_17545,N_17419);
nand UO_390 (O_390,N_16874,N_18639);
or UO_391 (O_391,N_19653,N_16357);
xnor UO_392 (O_392,N_19647,N_17600);
nand UO_393 (O_393,N_18785,N_19052);
nor UO_394 (O_394,N_16454,N_19598);
or UO_395 (O_395,N_19886,N_18406);
xor UO_396 (O_396,N_19685,N_17436);
or UO_397 (O_397,N_15080,N_15411);
or UO_398 (O_398,N_18876,N_17453);
nand UO_399 (O_399,N_19767,N_15040);
and UO_400 (O_400,N_18372,N_18800);
nand UO_401 (O_401,N_16433,N_19156);
nand UO_402 (O_402,N_17246,N_19485);
and UO_403 (O_403,N_15310,N_19736);
xnor UO_404 (O_404,N_19435,N_15234);
or UO_405 (O_405,N_18890,N_18480);
or UO_406 (O_406,N_19743,N_17755);
nand UO_407 (O_407,N_17627,N_16256);
nor UO_408 (O_408,N_15096,N_16627);
or UO_409 (O_409,N_16807,N_15427);
nor UO_410 (O_410,N_16107,N_15905);
nor UO_411 (O_411,N_16347,N_16714);
or UO_412 (O_412,N_18628,N_17203);
or UO_413 (O_413,N_15585,N_16005);
and UO_414 (O_414,N_18692,N_19265);
nand UO_415 (O_415,N_18274,N_17650);
nand UO_416 (O_416,N_17455,N_16775);
xnor UO_417 (O_417,N_17481,N_17300);
and UO_418 (O_418,N_15229,N_19782);
nor UO_419 (O_419,N_16228,N_19166);
and UO_420 (O_420,N_15539,N_15843);
or UO_421 (O_421,N_17551,N_18083);
and UO_422 (O_422,N_17001,N_18683);
xor UO_423 (O_423,N_19345,N_19878);
nor UO_424 (O_424,N_17868,N_16612);
or UO_425 (O_425,N_17434,N_18934);
and UO_426 (O_426,N_15863,N_19548);
or UO_427 (O_427,N_17250,N_19849);
or UO_428 (O_428,N_17059,N_15327);
nand UO_429 (O_429,N_18886,N_18037);
xor UO_430 (O_430,N_18183,N_18036);
or UO_431 (O_431,N_17055,N_18730);
xnor UO_432 (O_432,N_16896,N_15061);
xnor UO_433 (O_433,N_15392,N_17682);
xnor UO_434 (O_434,N_15287,N_17334);
and UO_435 (O_435,N_15631,N_19362);
xor UO_436 (O_436,N_17748,N_15517);
xnor UO_437 (O_437,N_16193,N_15048);
and UO_438 (O_438,N_15413,N_19506);
xnor UO_439 (O_439,N_16271,N_19134);
nor UO_440 (O_440,N_16889,N_19902);
and UO_441 (O_441,N_18449,N_17373);
xnor UO_442 (O_442,N_15011,N_15646);
xor UO_443 (O_443,N_19654,N_16131);
or UO_444 (O_444,N_18244,N_17569);
nor UO_445 (O_445,N_16151,N_18540);
nand UO_446 (O_446,N_19913,N_19596);
and UO_447 (O_447,N_19344,N_15620);
nand UO_448 (O_448,N_19221,N_18556);
or UO_449 (O_449,N_16886,N_16030);
and UO_450 (O_450,N_17326,N_18216);
xor UO_451 (O_451,N_17901,N_17052);
and UO_452 (O_452,N_18196,N_17321);
nor UO_453 (O_453,N_19306,N_18516);
xor UO_454 (O_454,N_15239,N_18217);
or UO_455 (O_455,N_16162,N_18786);
or UO_456 (O_456,N_15185,N_16134);
or UO_457 (O_457,N_16729,N_15067);
nor UO_458 (O_458,N_15855,N_17119);
nor UO_459 (O_459,N_15967,N_17138);
nor UO_460 (O_460,N_18805,N_19858);
or UO_461 (O_461,N_16244,N_15593);
or UO_462 (O_462,N_19313,N_19342);
or UO_463 (O_463,N_19526,N_16918);
xor UO_464 (O_464,N_16229,N_18779);
nand UO_465 (O_465,N_17141,N_16144);
xor UO_466 (O_466,N_15308,N_18282);
and UO_467 (O_467,N_17798,N_17854);
xnor UO_468 (O_468,N_15975,N_18959);
nor UO_469 (O_469,N_17542,N_18536);
nor UO_470 (O_470,N_16239,N_17556);
and UO_471 (O_471,N_15957,N_16786);
nor UO_472 (O_472,N_19837,N_17169);
nor UO_473 (O_473,N_17610,N_16168);
nand UO_474 (O_474,N_15166,N_16474);
nor UO_475 (O_475,N_15868,N_18159);
nor UO_476 (O_476,N_17944,N_16739);
and UO_477 (O_477,N_16139,N_17802);
nand UO_478 (O_478,N_15560,N_16683);
or UO_479 (O_479,N_17898,N_17050);
xnor UO_480 (O_480,N_19724,N_19758);
nand UO_481 (O_481,N_16476,N_17952);
xnor UO_482 (O_482,N_15901,N_19568);
nand UO_483 (O_483,N_19975,N_17442);
xnor UO_484 (O_484,N_19003,N_19086);
nor UO_485 (O_485,N_19728,N_17886);
or UO_486 (O_486,N_17920,N_17308);
nor UO_487 (O_487,N_16551,N_17103);
xnor UO_488 (O_488,N_15980,N_15491);
nand UO_489 (O_489,N_18346,N_18079);
xnor UO_490 (O_490,N_15561,N_19592);
xnor UO_491 (O_491,N_19393,N_19648);
or UO_492 (O_492,N_15708,N_15510);
or UO_493 (O_493,N_16834,N_17477);
or UO_494 (O_494,N_17160,N_18422);
xor UO_495 (O_495,N_15976,N_17457);
nor UO_496 (O_496,N_15296,N_17278);
xnor UO_497 (O_497,N_17928,N_17826);
and UO_498 (O_498,N_19124,N_17129);
nor UO_499 (O_499,N_17435,N_19268);
and UO_500 (O_500,N_16120,N_15007);
or UO_501 (O_501,N_18644,N_15823);
nor UO_502 (O_502,N_15542,N_15825);
and UO_503 (O_503,N_17684,N_18073);
nor UO_504 (O_504,N_18509,N_16638);
or UO_505 (O_505,N_17225,N_15347);
nor UO_506 (O_506,N_15402,N_17567);
and UO_507 (O_507,N_18154,N_15183);
nor UO_508 (O_508,N_15934,N_18579);
xnor UO_509 (O_509,N_16130,N_18276);
nor UO_510 (O_510,N_18676,N_18921);
nor UO_511 (O_511,N_15194,N_17432);
xor UO_512 (O_512,N_19080,N_16759);
nand UO_513 (O_513,N_19023,N_15996);
or UO_514 (O_514,N_15515,N_17839);
and UO_515 (O_515,N_15232,N_19580);
xnor UO_516 (O_516,N_18851,N_18093);
nor UO_517 (O_517,N_16501,N_15596);
or UO_518 (O_518,N_19388,N_19701);
nor UO_519 (O_519,N_16925,N_16122);
and UO_520 (O_520,N_18407,N_15768);
nand UO_521 (O_521,N_19536,N_16629);
and UO_522 (O_522,N_15357,N_18428);
and UO_523 (O_523,N_17446,N_17029);
and UO_524 (O_524,N_17175,N_17694);
xnor UO_525 (O_525,N_19201,N_18984);
nor UO_526 (O_526,N_17740,N_18849);
or UO_527 (O_527,N_15051,N_19702);
and UO_528 (O_528,N_16663,N_18788);
nor UO_529 (O_529,N_18218,N_18936);
xor UO_530 (O_530,N_18720,N_19738);
nor UO_531 (O_531,N_18753,N_15213);
xnor UO_532 (O_532,N_19438,N_15318);
and UO_533 (O_533,N_17087,N_19992);
and UO_534 (O_534,N_19584,N_19916);
nand UO_535 (O_535,N_16102,N_19632);
and UO_536 (O_536,N_19749,N_18402);
xnor UO_537 (O_537,N_16831,N_18819);
or UO_538 (O_538,N_19637,N_17572);
nor UO_539 (O_539,N_15822,N_19044);
and UO_540 (O_540,N_17044,N_15279);
nor UO_541 (O_541,N_15530,N_17742);
or UO_542 (O_542,N_19069,N_15925);
nor UO_543 (O_543,N_17805,N_19281);
xnor UO_544 (O_544,N_18975,N_16317);
or UO_545 (O_545,N_15781,N_16364);
and UO_546 (O_546,N_19457,N_18311);
or UO_547 (O_547,N_17911,N_15988);
xnor UO_548 (O_548,N_17693,N_17817);
nand UO_549 (O_549,N_19873,N_15481);
and UO_550 (O_550,N_19575,N_15679);
or UO_551 (O_551,N_19911,N_16018);
or UO_552 (O_552,N_19260,N_17288);
or UO_553 (O_553,N_18632,N_17706);
nand UO_554 (O_554,N_16906,N_15283);
xnor UO_555 (O_555,N_15893,N_17851);
nand UO_556 (O_556,N_16381,N_19440);
nand UO_557 (O_557,N_15142,N_17343);
nand UO_558 (O_558,N_16701,N_15911);
and UO_559 (O_559,N_16711,N_17240);
or UO_560 (O_560,N_16955,N_17589);
nand UO_561 (O_561,N_15180,N_18988);
nor UO_562 (O_562,N_17197,N_18880);
nand UO_563 (O_563,N_18455,N_18207);
or UO_564 (O_564,N_17900,N_19815);
or UO_565 (O_565,N_15497,N_16080);
xor UO_566 (O_566,N_19680,N_15304);
nand UO_567 (O_567,N_18400,N_17739);
nand UO_568 (O_568,N_17668,N_18634);
nor UO_569 (O_569,N_19458,N_19489);
nand UO_570 (O_570,N_19257,N_19428);
nor UO_571 (O_571,N_19030,N_17573);
xnor UO_572 (O_572,N_18166,N_19309);
xnor UO_573 (O_573,N_19739,N_18633);
xor UO_574 (O_574,N_17214,N_15650);
xor UO_575 (O_575,N_16688,N_18004);
nor UO_576 (O_576,N_15335,N_16063);
nand UO_577 (O_577,N_15328,N_16642);
xnor UO_578 (O_578,N_18418,N_17778);
nor UO_579 (O_579,N_16191,N_16135);
xnor UO_580 (O_580,N_15297,N_19248);
nand UO_581 (O_581,N_16109,N_17226);
and UO_582 (O_582,N_16396,N_18170);
or UO_583 (O_583,N_15223,N_15127);
or UO_584 (O_584,N_18351,N_15066);
and UO_585 (O_585,N_15619,N_19914);
xnor UO_586 (O_586,N_16968,N_18120);
or UO_587 (O_587,N_18474,N_19491);
and UO_588 (O_588,N_19089,N_15792);
and UO_589 (O_589,N_19964,N_18462);
xnor UO_590 (O_590,N_15859,N_15073);
or UO_591 (O_591,N_17787,N_16249);
xnor UO_592 (O_592,N_16547,N_15674);
or UO_593 (O_593,N_15459,N_18844);
and UO_594 (O_594,N_18179,N_15746);
or UO_595 (O_595,N_15872,N_17885);
nand UO_596 (O_596,N_19912,N_19503);
or UO_597 (O_597,N_19375,N_16272);
nor UO_598 (O_598,N_15368,N_17948);
xor UO_599 (O_599,N_17338,N_18337);
nor UO_600 (O_600,N_15092,N_16375);
nand UO_601 (O_601,N_19106,N_15303);
and UO_602 (O_602,N_18992,N_16315);
xnor UO_603 (O_603,N_15117,N_17845);
xor UO_604 (O_604,N_19670,N_19254);
xor UO_605 (O_605,N_15636,N_16064);
xor UO_606 (O_606,N_16680,N_16061);
or UO_607 (O_607,N_15322,N_18205);
nand UO_608 (O_608,N_17120,N_19517);
xnor UO_609 (O_609,N_19130,N_15024);
and UO_610 (O_610,N_16194,N_15696);
nand UO_611 (O_611,N_17769,N_17560);
nor UO_612 (O_612,N_18363,N_18285);
and UO_613 (O_613,N_18775,N_19550);
xor UO_614 (O_614,N_16677,N_16924);
nor UO_615 (O_615,N_16594,N_19303);
and UO_616 (O_616,N_16331,N_17824);
and UO_617 (O_617,N_18045,N_18011);
and UO_618 (O_618,N_19971,N_19293);
xor UO_619 (O_619,N_17306,N_16875);
or UO_620 (O_620,N_16056,N_15782);
and UO_621 (O_621,N_15513,N_16042);
xor UO_622 (O_622,N_17108,N_16421);
nor UO_623 (O_623,N_15774,N_18171);
or UO_624 (O_624,N_16843,N_18508);
and UO_625 (O_625,N_18774,N_16009);
xor UO_626 (O_626,N_16861,N_16669);
nand UO_627 (O_627,N_17007,N_15111);
xnor UO_628 (O_628,N_17905,N_18251);
or UO_629 (O_629,N_19566,N_16031);
and UO_630 (O_630,N_19841,N_19944);
nor UO_631 (O_631,N_19544,N_16791);
nor UO_632 (O_632,N_16348,N_18141);
nor UO_633 (O_633,N_19719,N_16828);
xnor UO_634 (O_634,N_16092,N_19982);
or UO_635 (O_635,N_16188,N_16311);
nor UO_636 (O_636,N_17180,N_17797);
and UO_637 (O_637,N_16404,N_19759);
nand UO_638 (O_638,N_15770,N_15499);
xor UO_639 (O_639,N_15209,N_18670);
and UO_640 (O_640,N_18912,N_17426);
or UO_641 (O_641,N_17679,N_17959);
xor UO_642 (O_642,N_19630,N_17506);
xor UO_643 (O_643,N_19062,N_19532);
or UO_644 (O_644,N_19258,N_17490);
xnor UO_645 (O_645,N_15920,N_17484);
or UO_646 (O_646,N_16761,N_17500);
nor UO_647 (O_647,N_18358,N_16402);
and UO_648 (O_648,N_15750,N_17872);
or UO_649 (O_649,N_17234,N_17954);
nor UO_650 (O_650,N_19668,N_19663);
or UO_651 (O_651,N_15641,N_15006);
and UO_652 (O_652,N_18184,N_15355);
nand UO_653 (O_653,N_17471,N_16338);
and UO_654 (O_654,N_18128,N_18502);
and UO_655 (O_655,N_17618,N_18593);
xnor UO_656 (O_656,N_19624,N_17450);
nor UO_657 (O_657,N_17315,N_19894);
or UO_658 (O_658,N_17958,N_16684);
and UO_659 (O_659,N_17222,N_19479);
or UO_660 (O_660,N_17264,N_15070);
or UO_661 (O_661,N_19081,N_15506);
and UO_662 (O_662,N_18758,N_18144);
nor UO_663 (O_663,N_16040,N_18615);
and UO_664 (O_664,N_15836,N_15828);
nor UO_665 (O_665,N_17126,N_17934);
xor UO_666 (O_666,N_15556,N_18578);
xnor UO_667 (O_667,N_15424,N_16442);
nor UO_668 (O_668,N_19327,N_19876);
or UO_669 (O_669,N_19466,N_18392);
or UO_670 (O_670,N_18915,N_18681);
and UO_671 (O_671,N_19756,N_15632);
xnor UO_672 (O_672,N_18309,N_16608);
nand UO_673 (O_673,N_19136,N_16556);
nand UO_674 (O_674,N_18442,N_15121);
and UO_675 (O_675,N_18115,N_16749);
or UO_676 (O_676,N_18622,N_17971);
nand UO_677 (O_677,N_16743,N_15113);
and UO_678 (O_678,N_19237,N_16072);
xnor UO_679 (O_679,N_15529,N_16084);
and UO_680 (O_680,N_16868,N_19905);
nand UO_681 (O_681,N_15383,N_16650);
nor UO_682 (O_682,N_16259,N_18557);
or UO_683 (O_683,N_16817,N_19984);
and UO_684 (O_684,N_16258,N_16667);
xor UO_685 (O_685,N_17873,N_16180);
or UO_686 (O_686,N_16850,N_18248);
xnor UO_687 (O_687,N_17879,N_15874);
nand UO_688 (O_688,N_17281,N_16359);
xor UO_689 (O_689,N_19061,N_17782);
and UO_690 (O_690,N_15846,N_17669);
nand UO_691 (O_691,N_16179,N_17448);
or UO_692 (O_692,N_15993,N_19294);
xnor UO_693 (O_693,N_17993,N_19173);
xnor UO_694 (O_694,N_18361,N_17910);
or UO_695 (O_695,N_18699,N_15720);
xor UO_696 (O_696,N_17051,N_16777);
xnor UO_697 (O_697,N_17521,N_17972);
xnor UO_698 (O_698,N_15902,N_19111);
or UO_699 (O_699,N_16310,N_18871);
nor UO_700 (O_700,N_16123,N_16879);
and UO_701 (O_701,N_18057,N_18672);
nor UO_702 (O_702,N_19307,N_18687);
or UO_703 (O_703,N_15437,N_19212);
xor UO_704 (O_704,N_19186,N_18607);
xnor UO_705 (O_705,N_18006,N_16789);
or UO_706 (O_706,N_16565,N_19107);
or UO_707 (O_707,N_16075,N_17285);
nand UO_708 (O_708,N_17427,N_18062);
or UO_709 (O_709,N_15765,N_16712);
nand UO_710 (O_710,N_16856,N_19430);
nand UO_711 (O_711,N_17058,N_18716);
and UO_712 (O_712,N_19820,N_15256);
nand UO_713 (O_713,N_19959,N_19380);
nand UO_714 (O_714,N_16607,N_16289);
and UO_715 (O_715,N_15473,N_17594);
nand UO_716 (O_716,N_19574,N_18047);
nor UO_717 (O_717,N_16738,N_16422);
xor UO_718 (O_718,N_19888,N_19270);
xor UO_719 (O_719,N_18044,N_19549);
nor UO_720 (O_720,N_17102,N_17096);
or UO_721 (O_721,N_18811,N_18405);
xor UO_722 (O_722,N_18790,N_15602);
nand UO_723 (O_723,N_19925,N_19026);
and UO_724 (O_724,N_16672,N_16829);
and UO_725 (O_725,N_15756,N_19486);
nor UO_726 (O_726,N_18641,N_15927);
nor UO_727 (O_727,N_17495,N_19754);
nor UO_728 (O_728,N_15309,N_19601);
xor UO_729 (O_729,N_17228,N_17414);
and UO_730 (O_730,N_19278,N_16521);
and UO_731 (O_731,N_15455,N_19956);
xnor UO_732 (O_732,N_16649,N_15795);
and UO_733 (O_733,N_16520,N_16154);
or UO_734 (O_734,N_17728,N_17005);
nor UO_735 (O_735,N_17818,N_15373);
or UO_736 (O_736,N_19825,N_19460);
nand UO_737 (O_737,N_15369,N_17766);
and UO_738 (O_738,N_16809,N_18086);
xnor UO_739 (O_739,N_15955,N_15495);
and UO_740 (O_740,N_17410,N_15027);
and UO_741 (O_741,N_18452,N_15119);
nand UO_742 (O_742,N_19796,N_18764);
nor UO_743 (O_743,N_18290,N_17838);
and UO_744 (O_744,N_16923,N_17801);
nand UO_745 (O_745,N_18065,N_18032);
nor UO_746 (O_746,N_17345,N_15841);
xnor UO_747 (O_747,N_19623,N_19529);
or UO_748 (O_748,N_16252,N_16760);
nand UO_749 (O_749,N_15395,N_15728);
xnor UO_750 (O_750,N_16755,N_15496);
or UO_751 (O_751,N_18605,N_15710);
xnor UO_752 (O_752,N_16332,N_19826);
and UO_753 (O_753,N_15468,N_15257);
nor UO_754 (O_754,N_19847,N_19978);
and UO_755 (O_755,N_15130,N_19729);
xor UO_756 (O_756,N_17715,N_15055);
and UO_757 (O_757,N_19153,N_19478);
xnor UO_758 (O_758,N_17783,N_17221);
nor UO_759 (O_759,N_18674,N_15566);
xor UO_760 (O_760,N_17809,N_17415);
nor UO_761 (O_761,N_17157,N_19284);
xor UO_762 (O_762,N_17671,N_17057);
or UO_763 (O_763,N_17217,N_19290);
nand UO_764 (O_764,N_15299,N_15550);
nor UO_765 (O_765,N_15818,N_19881);
nor UO_766 (O_766,N_15432,N_19223);
xnor UO_767 (O_767,N_17195,N_15637);
xor UO_768 (O_768,N_16383,N_17136);
nor UO_769 (O_769,N_17361,N_18493);
and UO_770 (O_770,N_15187,N_15563);
and UO_771 (O_771,N_18640,N_17760);
xnor UO_772 (O_772,N_19588,N_15807);
nand UO_773 (O_773,N_15618,N_15676);
and UO_774 (O_774,N_17362,N_19571);
and UO_775 (O_775,N_19603,N_19050);
and UO_776 (O_776,N_18322,N_18600);
or UO_777 (O_777,N_15528,N_15292);
and UO_778 (O_778,N_19158,N_16325);
and UO_779 (O_779,N_18257,N_17700);
xnor UO_780 (O_780,N_16783,N_19049);
xnor UO_781 (O_781,N_15430,N_18884);
nor UO_782 (O_782,N_19301,N_15158);
nor UO_783 (O_783,N_15337,N_15938);
nand UO_784 (O_784,N_18808,N_18951);
or UO_785 (O_785,N_15931,N_18993);
nor UO_786 (O_786,N_15277,N_17199);
nand UO_787 (O_787,N_16052,N_19991);
or UO_788 (O_788,N_17698,N_16920);
or UO_789 (O_789,N_17581,N_15269);
xnor UO_790 (O_790,N_15943,N_16371);
or UO_791 (O_791,N_19823,N_18519);
or UO_792 (O_792,N_19896,N_18340);
and UO_793 (O_793,N_16954,N_16992);
and UO_794 (O_794,N_15429,N_15189);
nor UO_795 (O_795,N_18451,N_18211);
or UO_796 (O_796,N_18301,N_18414);
xor UO_797 (O_797,N_15727,N_19402);
nand UO_798 (O_798,N_15122,N_16720);
nor UO_799 (O_799,N_17193,N_18410);
xor UO_800 (O_800,N_18355,N_15071);
nand UO_801 (O_801,N_19750,N_15492);
and UO_802 (O_802,N_16140,N_17356);
and UO_803 (O_803,N_17425,N_17976);
and UO_804 (O_804,N_15666,N_19733);
and UO_805 (O_805,N_15115,N_15097);
nor UO_806 (O_806,N_17579,N_17523);
xnor UO_807 (O_807,N_15477,N_18092);
nand UO_808 (O_808,N_16950,N_19475);
nor UO_809 (O_809,N_18204,N_15665);
nor UO_810 (O_810,N_16503,N_15910);
nand UO_811 (O_811,N_16240,N_17271);
xnor UO_812 (O_812,N_16339,N_18028);
or UO_813 (O_813,N_19146,N_18942);
xnor UO_814 (O_814,N_18546,N_16219);
nor UO_815 (O_815,N_17440,N_17557);
nand UO_816 (O_816,N_15400,N_15041);
nor UO_817 (O_817,N_15135,N_16204);
nand UO_818 (O_818,N_19611,N_15712);
xnor UO_819 (O_819,N_16045,N_15022);
nand UO_820 (O_820,N_16958,N_16351);
nor UO_821 (O_821,N_18755,N_15467);
nand UO_822 (O_822,N_19938,N_18598);
and UO_823 (O_823,N_15817,N_16784);
nand UO_824 (O_824,N_19943,N_19492);
and UO_825 (O_825,N_18306,N_18341);
xnor UO_826 (O_826,N_17480,N_16431);
and UO_827 (O_827,N_18326,N_16984);
nand UO_828 (O_828,N_17695,N_18460);
xnor UO_829 (O_829,N_16839,N_16057);
nor UO_830 (O_830,N_17303,N_18559);
nor UO_831 (O_831,N_16991,N_16822);
or UO_832 (O_832,N_15023,N_15313);
and UO_833 (O_833,N_17131,N_17654);
or UO_834 (O_834,N_17370,N_18863);
nor UO_835 (O_835,N_19131,N_15867);
or UO_836 (O_836,N_17086,N_18745);
xnor UO_837 (O_837,N_15586,N_17325);
nor UO_838 (O_838,N_15835,N_16141);
nor UO_839 (O_839,N_19405,N_18532);
nor UO_840 (O_840,N_19731,N_16074);
nor UO_841 (O_841,N_17411,N_18937);
nor UO_842 (O_842,N_19045,N_19473);
or UO_843 (O_843,N_16243,N_16933);
xnor UO_844 (O_844,N_15700,N_18354);
or UO_845 (O_845,N_16037,N_18931);
xor UO_846 (O_846,N_16633,N_17962);
nor UO_847 (O_847,N_18048,N_17609);
nand UO_848 (O_848,N_16636,N_15434);
and UO_849 (O_849,N_16985,N_19228);
nor UO_850 (O_850,N_17045,N_19780);
or UO_851 (O_851,N_19909,N_16965);
and UO_852 (O_852,N_19949,N_15638);
nor UO_853 (O_853,N_19835,N_18663);
nor UO_854 (O_854,N_15695,N_19703);
xnor UO_855 (O_855,N_16276,N_18894);
nand UO_856 (O_856,N_15716,N_18454);
nand UO_857 (O_857,N_19748,N_17123);
and UO_858 (O_858,N_19868,N_18560);
and UO_859 (O_859,N_16342,N_19874);
nor UO_860 (O_860,N_18478,N_16392);
nor UO_861 (O_861,N_16125,N_18015);
nand UO_862 (O_862,N_15359,N_15569);
nand UO_863 (O_863,N_16723,N_19795);
nor UO_864 (O_864,N_16293,N_17576);
nor UO_865 (O_865,N_16190,N_18489);
nor UO_866 (O_866,N_16232,N_17016);
and UO_867 (O_867,N_16537,N_16027);
and UO_868 (O_868,N_19935,N_18971);
and UO_869 (O_869,N_15932,N_19352);
nor UO_870 (O_870,N_16951,N_15675);
nand UO_871 (O_871,N_17531,N_19195);
or UO_872 (O_872,N_19776,N_16234);
and UO_873 (O_873,N_16334,N_15971);
xor UO_874 (O_874,N_16915,N_16469);
xor UO_875 (O_875,N_15726,N_17355);
and UO_876 (O_876,N_16936,N_19691);
and UO_877 (O_877,N_19364,N_17674);
or UO_878 (O_878,N_17996,N_19885);
nand UO_879 (O_879,N_19224,N_15025);
nor UO_880 (O_880,N_16117,N_19730);
xnor UO_881 (O_881,N_18694,N_17211);
and UO_882 (O_882,N_19817,N_16088);
or UO_883 (O_883,N_17588,N_15547);
xnor UO_884 (O_884,N_18387,N_16956);
nand UO_885 (O_885,N_16937,N_16250);
nand UO_886 (O_886,N_17143,N_16087);
xnor UO_887 (O_887,N_18726,N_19523);
or UO_888 (O_888,N_19429,N_15325);
or UO_889 (O_889,N_17258,N_15747);
nor UO_890 (O_890,N_15398,N_19085);
and UO_891 (O_891,N_16262,N_17210);
xor UO_892 (O_892,N_17470,N_15105);
or UO_893 (O_893,N_19323,N_15005);
xnor UO_894 (O_894,N_16769,N_19547);
or UO_895 (O_895,N_15019,N_15237);
nand UO_896 (O_896,N_18857,N_17789);
or UO_897 (O_897,N_16236,N_19824);
xnor UO_898 (O_898,N_15573,N_15984);
nand UO_899 (O_899,N_16269,N_16222);
nand UO_900 (O_900,N_19155,N_18229);
xor UO_901 (O_901,N_15899,N_17903);
xor UO_902 (O_902,N_18794,N_19614);
or UO_903 (O_903,N_17111,N_19590);
nor UO_904 (O_904,N_15509,N_16763);
or UO_905 (O_905,N_15154,N_16715);
and UO_906 (O_906,N_16808,N_15311);
nand UO_907 (O_907,N_18020,N_17612);
nand UO_908 (O_908,N_16619,N_16479);
or UO_909 (O_909,N_18981,N_15851);
nor UO_910 (O_910,N_19410,N_16833);
or UO_911 (O_911,N_16196,N_16198);
nand UO_912 (O_912,N_18682,N_19903);
or UO_913 (O_913,N_16224,N_16802);
and UO_914 (O_914,N_19877,N_19147);
and UO_915 (O_915,N_18631,N_16372);
and UO_916 (O_916,N_16013,N_18135);
or UO_917 (O_917,N_16944,N_19942);
nor UO_918 (O_918,N_18140,N_19890);
xnor UO_919 (O_919,N_16905,N_15683);
nand UO_920 (O_920,N_15133,N_18703);
nand UO_921 (O_921,N_16436,N_16746);
nand UO_922 (O_922,N_19222,N_19019);
or UO_923 (O_923,N_18280,N_19427);
and UO_924 (O_924,N_16754,N_15589);
xor UO_925 (O_925,N_19034,N_19296);
and UO_926 (O_926,N_15293,N_16606);
and UO_927 (O_927,N_18439,N_16429);
xnor UO_928 (O_928,N_19162,N_19291);
xnor UO_929 (O_929,N_19813,N_16085);
nor UO_930 (O_930,N_17741,N_16113);
nor UO_931 (O_931,N_18860,N_16466);
or UO_932 (O_932,N_18099,N_16696);
xor UO_933 (O_933,N_18138,N_16624);
and UO_934 (O_934,N_17155,N_18394);
nor UO_935 (O_935,N_17461,N_16497);
and UO_936 (O_936,N_17807,N_17002);
and UO_937 (O_937,N_16510,N_15016);
or UO_938 (O_938,N_17178,N_16288);
and UO_939 (O_939,N_19009,N_19842);
nor UO_940 (O_940,N_19610,N_15447);
nand UO_941 (O_941,N_17605,N_17812);
nor UO_942 (O_942,N_17209,N_18723);
nor UO_943 (O_943,N_17125,N_19789);
or UO_944 (O_944,N_18510,N_16296);
nor UO_945 (O_945,N_16910,N_19948);
nor UO_946 (O_946,N_16679,N_17753);
xor UO_947 (O_947,N_17574,N_18650);
nand UO_948 (O_948,N_17925,N_17070);
xnor UO_949 (O_949,N_18381,N_16059);
nor UO_950 (O_950,N_15345,N_16437);
xnor UO_951 (O_951,N_15840,N_17031);
and UO_952 (O_952,N_17849,N_18077);
and UO_953 (O_953,N_19058,N_17312);
nand UO_954 (O_954,N_16108,N_19036);
nand UO_955 (O_955,N_15562,N_19976);
xor UO_956 (O_956,N_15059,N_19012);
xor UO_957 (O_957,N_15249,N_15323);
and UO_958 (O_958,N_18371,N_18737);
or UO_959 (O_959,N_19833,N_17295);
and UO_960 (O_960,N_16529,N_15038);
or UO_961 (O_961,N_18739,N_15376);
xor UO_962 (O_962,N_19379,N_18743);
or UO_963 (O_963,N_19643,N_18272);
nand UO_964 (O_964,N_18470,N_19338);
xor UO_965 (O_965,N_17156,N_18873);
nor UO_966 (O_966,N_18702,N_18258);
nor UO_967 (O_967,N_18264,N_16656);
and UO_968 (O_968,N_19582,N_17703);
and UO_969 (O_969,N_15543,N_15204);
nor UO_970 (O_970,N_16793,N_18379);
nor UO_971 (O_971,N_18746,N_18875);
nand UO_972 (O_972,N_16959,N_18479);
xnor UO_973 (O_973,N_17861,N_18881);
xnor UO_974 (O_974,N_16757,N_18107);
xnor UO_975 (O_975,N_16119,N_17493);
nor UO_976 (O_976,N_16911,N_17565);
xnor UO_977 (O_977,N_19777,N_15892);
nand UO_978 (O_978,N_18448,N_19524);
and UO_979 (O_979,N_15640,N_16995);
and UO_980 (O_980,N_16050,N_17313);
nor UO_981 (O_981,N_17048,N_16620);
xnor UO_982 (O_982,N_19883,N_19120);
nor UO_983 (O_983,N_18181,N_16898);
nor UO_984 (O_984,N_15915,N_16735);
and UO_985 (O_985,N_18469,N_17522);
nor UO_986 (O_986,N_15331,N_18396);
xor UO_987 (O_987,N_17145,N_16756);
nor UO_988 (O_988,N_15168,N_16090);
or UO_989 (O_989,N_15554,N_15344);
or UO_990 (O_990,N_15176,N_19164);
nand UO_991 (O_991,N_17946,N_18377);
xnor UO_992 (O_992,N_15579,N_18728);
or UO_993 (O_993,N_18918,N_17864);
and UO_994 (O_994,N_17316,N_18386);
and UO_995 (O_995,N_16036,N_18468);
xor UO_996 (O_996,N_16894,N_18566);
nor UO_997 (O_997,N_19378,N_16023);
and UO_998 (O_998,N_15243,N_15503);
or UO_999 (O_999,N_17469,N_18698);
nor UO_1000 (O_1000,N_18398,N_17168);
and UO_1001 (O_1001,N_19741,N_18933);
and UO_1002 (O_1002,N_17516,N_17212);
nand UO_1003 (O_1003,N_18535,N_19669);
xnor UO_1004 (O_1004,N_17463,N_18247);
or UO_1005 (O_1005,N_19512,N_15440);
xnor UO_1006 (O_1006,N_18760,N_15544);
xnor UO_1007 (O_1007,N_16639,N_18343);
or UO_1008 (O_1008,N_15100,N_16245);
nor UO_1009 (O_1009,N_16674,N_15246);
nor UO_1010 (O_1010,N_17555,N_15824);
and UO_1011 (O_1011,N_19910,N_18312);
or UO_1012 (O_1012,N_18375,N_17732);
or UO_1013 (O_1013,N_17158,N_16574);
xnor UO_1014 (O_1014,N_17915,N_15118);
nand UO_1015 (O_1015,N_16363,N_16571);
or UO_1016 (O_1016,N_19744,N_16519);
nor UO_1017 (O_1017,N_17254,N_19818);
or UO_1018 (O_1018,N_18968,N_15961);
and UO_1019 (O_1019,N_18225,N_16586);
xor UO_1020 (O_1020,N_18334,N_19051);
nor UO_1021 (O_1021,N_19139,N_15564);
nor UO_1022 (O_1022,N_16452,N_19450);
xnor UO_1023 (O_1023,N_18887,N_19214);
and UO_1024 (O_1024,N_19117,N_15945);
and UO_1025 (O_1025,N_19615,N_19445);
and UO_1026 (O_1026,N_17585,N_19606);
nand UO_1027 (O_1027,N_15849,N_16138);
nor UO_1028 (O_1028,N_19589,N_17389);
xnor UO_1029 (O_1029,N_15076,N_16689);
or UO_1030 (O_1030,N_15657,N_16790);
and UO_1031 (O_1031,N_15265,N_16747);
xor UO_1032 (O_1032,N_15426,N_15060);
nor UO_1033 (O_1033,N_17379,N_19299);
or UO_1034 (O_1034,N_18701,N_17930);
xnor UO_1035 (O_1035,N_16488,N_17115);
xnor UO_1036 (O_1036,N_16086,N_19190);
xnor UO_1037 (O_1037,N_17037,N_18680);
nor UO_1038 (O_1038,N_18941,N_19459);
or UO_1039 (O_1039,N_18953,N_15808);
and UO_1040 (O_1040,N_16173,N_18630);
nand UO_1041 (O_1041,N_17940,N_19543);
and UO_1042 (O_1042,N_15811,N_17980);
and UO_1043 (O_1043,N_19455,N_15207);
or UO_1044 (O_1044,N_17985,N_18978);
nand UO_1045 (O_1045,N_16658,N_16935);
and UO_1046 (O_1046,N_16257,N_15030);
nand UO_1047 (O_1047,N_18972,N_15390);
xor UO_1048 (O_1048,N_19498,N_18562);
nor UO_1049 (O_1049,N_15692,N_18112);
xor UO_1050 (O_1050,N_18323,N_18150);
or UO_1051 (O_1051,N_19628,N_16544);
or UO_1052 (O_1052,N_19011,N_18275);
or UO_1053 (O_1053,N_16492,N_15125);
xor UO_1054 (O_1054,N_17974,N_17866);
and UO_1055 (O_1055,N_16369,N_16704);
or UO_1056 (O_1056,N_17711,N_16811);
or UO_1057 (O_1057,N_17914,N_19556);
and UO_1058 (O_1058,N_16975,N_17754);
xnor UO_1059 (O_1059,N_18068,N_17710);
nand UO_1060 (O_1060,N_16780,N_18734);
xor UO_1061 (O_1061,N_18954,N_18119);
nand UO_1062 (O_1062,N_15668,N_17603);
nor UO_1063 (O_1063,N_19854,N_17422);
nor UO_1064 (O_1064,N_18721,N_15690);
nand UO_1065 (O_1065,N_18030,N_18995);
nand UO_1066 (O_1066,N_16393,N_18440);
or UO_1067 (O_1067,N_17725,N_15877);
and UO_1068 (O_1068,N_19985,N_18580);
and UO_1069 (O_1069,N_18944,N_17262);
nand UO_1070 (O_1070,N_17895,N_18055);
or UO_1071 (O_1071,N_19329,N_16340);
nand UO_1072 (O_1072,N_18441,N_17998);
nor UO_1073 (O_1073,N_18799,N_18391);
nor UO_1074 (O_1074,N_15317,N_18237);
or UO_1075 (O_1075,N_18445,N_17830);
nor UO_1076 (O_1076,N_18980,N_17284);
or UO_1077 (O_1077,N_15629,N_15363);
nand UO_1078 (O_1078,N_17268,N_18612);
xor UO_1079 (O_1079,N_15046,N_18298);
nand UO_1080 (O_1080,N_18102,N_17505);
xnor UO_1081 (O_1081,N_19784,N_19958);
and UO_1082 (O_1082,N_16261,N_19184);
nor UO_1083 (O_1083,N_19850,N_15688);
and UO_1084 (O_1084,N_16246,N_15441);
or UO_1085 (O_1085,N_19569,N_17472);
nand UO_1086 (O_1086,N_18761,N_15507);
nor UO_1087 (O_1087,N_16548,N_16934);
and UO_1088 (O_1088,N_17239,N_18651);
nor UO_1089 (O_1089,N_16200,N_15463);
xor UO_1090 (O_1090,N_16862,N_16657);
and UO_1091 (O_1091,N_19351,N_15647);
nor UO_1092 (O_1092,N_17459,N_15361);
xnor UO_1093 (O_1093,N_18152,N_19401);
xnor UO_1094 (O_1094,N_15288,N_15989);
or UO_1095 (O_1095,N_16026,N_17613);
or UO_1096 (O_1096,N_16827,N_15682);
nand UO_1097 (O_1097,N_15906,N_16360);
xor UO_1098 (O_1098,N_18836,N_17877);
xnor UO_1099 (O_1099,N_19658,N_15709);
nor UO_1100 (O_1100,N_15587,N_19966);
and UO_1101 (O_1101,N_19250,N_17405);
and UO_1102 (O_1102,N_19576,N_18113);
and UO_1103 (O_1103,N_15008,N_18365);
or UO_1104 (O_1104,N_19625,N_15054);
nand UO_1105 (O_1105,N_17648,N_19561);
or UO_1106 (O_1106,N_17596,N_16313);
nand UO_1107 (O_1107,N_16260,N_17277);
nor UO_1108 (O_1108,N_17837,N_19534);
nor UO_1109 (O_1109,N_19451,N_19141);
nor UO_1110 (O_1110,N_15449,N_19604);
or UO_1111 (O_1111,N_15802,N_15442);
nand UO_1112 (O_1112,N_18438,N_18175);
nor UO_1113 (O_1113,N_15655,N_16590);
or UO_1114 (O_1114,N_17869,N_18567);
xnor UO_1115 (O_1115,N_15801,N_15850);
nand UO_1116 (O_1116,N_19940,N_17015);
xor UO_1117 (O_1117,N_16116,N_15790);
or UO_1118 (O_1118,N_19318,N_16932);
nand UO_1119 (O_1119,N_15134,N_15422);
nor UO_1120 (O_1120,N_19742,N_17943);
or UO_1121 (O_1121,N_19493,N_17774);
or UO_1122 (O_1122,N_18085,N_18019);
and UO_1123 (O_1123,N_18231,N_15820);
xnor UO_1124 (O_1124,N_19068,N_16434);
or UO_1125 (O_1125,N_19247,N_19804);
nand UO_1126 (O_1126,N_19449,N_16238);
xnor UO_1127 (O_1127,N_16758,N_19638);
nand UO_1128 (O_1128,N_17069,N_19252);
and UO_1129 (O_1129,N_18339,N_15064);
nand UO_1130 (O_1130,N_15997,N_15913);
or UO_1131 (O_1131,N_16820,N_19115);
nand UO_1132 (O_1132,N_15338,N_17949);
nand UO_1133 (O_1133,N_15540,N_17681);
or UO_1134 (O_1134,N_16857,N_19311);
nor UO_1135 (O_1135,N_17580,N_16397);
or UO_1136 (O_1136,N_17488,N_17353);
and UO_1137 (O_1137,N_17977,N_16569);
xor UO_1138 (O_1138,N_16561,N_17518);
xnor UO_1139 (O_1139,N_17337,N_18296);
nor UO_1140 (O_1140,N_15789,N_16538);
nor UO_1141 (O_1141,N_15236,N_17670);
nor UO_1142 (O_1142,N_17332,N_16686);
nor UO_1143 (O_1143,N_15377,N_15149);
nand UO_1144 (O_1144,N_18026,N_18747);
or UO_1145 (O_1145,N_17191,N_16945);
xnor UO_1146 (O_1146,N_19407,N_15372);
nor UO_1147 (O_1147,N_17150,N_17152);
or UO_1148 (O_1148,N_16438,N_15000);
or UO_1149 (O_1149,N_18907,N_15842);
and UO_1150 (O_1150,N_16491,N_15399);
nor UO_1151 (O_1151,N_18427,N_15757);
or UO_1152 (O_1152,N_17963,N_15284);
and UO_1153 (O_1153,N_15110,N_19712);
nand UO_1154 (O_1154,N_17960,N_16922);
nor UO_1155 (O_1155,N_15651,N_18219);
or UO_1156 (O_1156,N_15713,N_17779);
and UO_1157 (O_1157,N_15329,N_18964);
or UO_1158 (O_1158,N_17298,N_17068);
and UO_1159 (O_1159,N_15128,N_18929);
xnor UO_1160 (O_1160,N_15478,N_17936);
nor UO_1161 (O_1161,N_16414,N_17975);
or UO_1162 (O_1162,N_15511,N_17196);
nand UO_1163 (O_1163,N_17969,N_15929);
nor UO_1164 (O_1164,N_17768,N_15922);
or UO_1165 (O_1165,N_18447,N_19934);
xor UO_1166 (O_1166,N_16413,N_19171);
and UO_1167 (O_1167,N_15574,N_19737);
or UO_1168 (O_1168,N_15815,N_15378);
and UO_1169 (O_1169,N_18283,N_18845);
nor UO_1170 (O_1170,N_17984,N_18129);
nand UO_1171 (O_1171,N_18611,N_19447);
nor UO_1172 (O_1172,N_19919,N_16724);
or UO_1173 (O_1173,N_15471,N_17458);
xnor UO_1174 (O_1174,N_19126,N_15252);
xnor UO_1175 (O_1175,N_17582,N_16900);
or UO_1176 (O_1176,N_17060,N_15238);
and UO_1177 (O_1177,N_19482,N_15089);
or UO_1178 (O_1178,N_19008,N_15225);
nand UO_1179 (O_1179,N_17853,N_15873);
nand UO_1180 (O_1180,N_17081,N_17659);
and UO_1181 (O_1181,N_18347,N_15393);
xnor UO_1182 (O_1182,N_19678,N_19261);
and UO_1183 (O_1183,N_17918,N_18331);
nor UO_1184 (O_1184,N_16821,N_17836);
nor UO_1185 (O_1185,N_19955,N_18035);
nor UO_1186 (O_1186,N_17223,N_19612);
and UO_1187 (O_1187,N_18182,N_17063);
nor UO_1188 (O_1188,N_16267,N_15148);
and UO_1189 (O_1189,N_17382,N_15753);
xnor UO_1190 (O_1190,N_15614,N_18417);
and UO_1191 (O_1191,N_15776,N_16952);
and UO_1192 (O_1192,N_17922,N_17867);
xnor UO_1193 (O_1193,N_19682,N_16341);
nand UO_1194 (O_1194,N_16601,N_18617);
or UO_1195 (O_1195,N_19839,N_18178);
xnor UO_1196 (O_1196,N_19113,N_17813);
or UO_1197 (O_1197,N_18459,N_18538);
nand UO_1198 (O_1198,N_15217,N_19552);
or UO_1199 (O_1199,N_16432,N_15926);
xor UO_1200 (O_1200,N_19993,N_19343);
nor UO_1201 (O_1201,N_19255,N_16600);
or UO_1202 (O_1202,N_18317,N_15643);
xor UO_1203 (O_1203,N_16417,N_17590);
xnor UO_1204 (O_1204,N_18594,N_15508);
xor UO_1205 (O_1205,N_19463,N_18563);
xnor UO_1206 (O_1206,N_16490,N_15379);
or UO_1207 (O_1207,N_19696,N_18623);
nand UO_1208 (O_1208,N_15033,N_15532);
and UO_1209 (O_1209,N_16515,N_19276);
or UO_1210 (O_1210,N_17046,N_19684);
or UO_1211 (O_1211,N_16016,N_19828);
and UO_1212 (O_1212,N_17413,N_15339);
xor UO_1213 (O_1213,N_15350,N_19467);
xor UO_1214 (O_1214,N_18319,N_17179);
or UO_1215 (O_1215,N_15169,N_19416);
nor UO_1216 (O_1216,N_17452,N_17716);
xor UO_1217 (O_1217,N_16307,N_16427);
or UO_1218 (O_1218,N_15192,N_19076);
nor UO_1219 (O_1219,N_19434,N_17167);
or UO_1220 (O_1220,N_16282,N_16695);
nor UO_1221 (O_1221,N_16914,N_19150);
xor UO_1222 (O_1222,N_18029,N_17987);
or UO_1223 (O_1223,N_15280,N_17465);
and UO_1224 (O_1224,N_17110,N_15112);
xor UO_1225 (O_1225,N_19656,N_17735);
xnor UO_1226 (O_1226,N_17010,N_17913);
and UO_1227 (O_1227,N_18710,N_18072);
nand UO_1228 (O_1228,N_17956,N_16707);
or UO_1229 (O_1229,N_16172,N_15191);
or UO_1230 (O_1230,N_17727,N_19860);
and UO_1231 (O_1231,N_18399,N_16708);
nand UO_1232 (O_1232,N_15454,N_19262);
and UO_1233 (O_1233,N_17107,N_19135);
nand UO_1234 (O_1234,N_17791,N_19007);
xnor UO_1235 (O_1235,N_16591,N_19322);
xnor UO_1236 (O_1236,N_17346,N_16810);
xor UO_1237 (O_1237,N_19188,N_18847);
xnor UO_1238 (O_1238,N_18643,N_15334);
nand UO_1239 (O_1239,N_17738,N_19510);
nand UO_1240 (O_1240,N_15685,N_17908);
xor UO_1241 (O_1241,N_18596,N_17548);
xor UO_1242 (O_1242,N_15968,N_18277);
nor UO_1243 (O_1243,N_19310,N_17344);
or UO_1244 (O_1244,N_16592,N_16844);
nor UO_1245 (O_1245,N_16980,N_18565);
nor UO_1246 (O_1246,N_17188,N_17561);
and UO_1247 (O_1247,N_17617,N_17501);
and UO_1248 (O_1248,N_18577,N_18648);
and UO_1249 (O_1249,N_17311,N_18833);
nand UO_1250 (O_1250,N_17577,N_16553);
and UO_1251 (O_1251,N_15274,N_16263);
nand UO_1252 (O_1252,N_19361,N_17255);
xor UO_1253 (O_1253,N_16385,N_19481);
xnor UO_1254 (O_1254,N_15366,N_18713);
xnor UO_1255 (O_1255,N_15952,N_16845);
or UO_1256 (O_1256,N_18076,N_16506);
xor UO_1257 (O_1257,N_15470,N_15273);
xor UO_1258 (O_1258,N_17970,N_19709);
nand UO_1259 (O_1259,N_17008,N_16685);
nand UO_1260 (O_1260,N_16157,N_18018);
nor UO_1261 (O_1261,N_17352,N_17517);
nand UO_1262 (O_1262,N_16851,N_18791);
and UO_1263 (O_1263,N_19229,N_16380);
xnor UO_1264 (O_1264,N_19219,N_16001);
and UO_1265 (O_1265,N_17757,N_16189);
nand UO_1266 (O_1266,N_18704,N_17137);
nor UO_1267 (O_1267,N_18742,N_17717);
nand UO_1268 (O_1268,N_19422,N_16480);
xor UO_1269 (O_1269,N_18420,N_16566);
nand UO_1270 (O_1270,N_16904,N_18548);
or UO_1271 (O_1271,N_19686,N_16727);
nand UO_1272 (O_1272,N_19289,N_18939);
nand UO_1273 (O_1273,N_19128,N_15951);
nand UO_1274 (O_1274,N_15336,N_15087);
nand UO_1275 (O_1275,N_18732,N_17347);
nand UO_1276 (O_1276,N_15681,N_15890);
or UO_1277 (O_1277,N_19488,N_19073);
nand UO_1278 (O_1278,N_17630,N_19022);
nor UO_1279 (O_1279,N_17478,N_15375);
and UO_1280 (O_1280,N_15155,N_17552);
xor UO_1281 (O_1281,N_19998,N_18962);
nor UO_1282 (O_1282,N_17835,N_18172);
xor UO_1283 (O_1283,N_15242,N_15365);
nor UO_1284 (O_1284,N_19439,N_19540);
or UO_1285 (O_1285,N_19231,N_15775);
or UO_1286 (O_1286,N_17104,N_17554);
nor UO_1287 (O_1287,N_15264,N_17101);
xnor UO_1288 (O_1288,N_16379,N_19720);
xnor UO_1289 (O_1289,N_15992,N_18070);
or UO_1290 (O_1290,N_19471,N_15645);
or UO_1291 (O_1291,N_19732,N_16703);
and UO_1292 (O_1292,N_16753,N_16887);
nor UO_1293 (O_1293,N_19769,N_17821);
or UO_1294 (O_1294,N_19244,N_17076);
or UO_1295 (O_1295,N_17351,N_15184);
nand UO_1296 (O_1296,N_19305,N_16622);
nor UO_1297 (O_1297,N_19551,N_18989);
and UO_1298 (O_1298,N_15260,N_16864);
or UO_1299 (O_1299,N_16444,N_19622);
or UO_1300 (O_1300,N_16079,N_16094);
nand UO_1301 (O_1301,N_19468,N_16077);
or UO_1302 (O_1302,N_19400,N_18541);
xnor UO_1303 (O_1303,N_19657,N_16800);
and UO_1304 (O_1304,N_15615,N_15178);
nand UO_1305 (O_1305,N_19271,N_15153);
or UO_1306 (O_1306,N_15995,N_15444);
nand UO_1307 (O_1307,N_17032,N_15415);
nor UO_1308 (O_1308,N_17696,N_16826);
and UO_1309 (O_1309,N_18431,N_17317);
xnor UO_1310 (O_1310,N_16000,N_17992);
nand UO_1311 (O_1311,N_17636,N_19861);
or UO_1312 (O_1312,N_18458,N_15484);
and UO_1313 (O_1313,N_16181,N_15519);
nand UO_1314 (O_1314,N_15211,N_17685);
xor UO_1315 (O_1315,N_16300,N_19063);
xor UO_1316 (O_1316,N_15536,N_15599);
nor UO_1317 (O_1317,N_19048,N_15717);
and UO_1318 (O_1318,N_17004,N_15963);
and UO_1319 (O_1319,N_15809,N_16899);
xor UO_1320 (O_1320,N_15034,N_16426);
or UO_1321 (O_1321,N_17252,N_17406);
nand UO_1322 (O_1322,N_18088,N_19859);
or UO_1323 (O_1323,N_18518,N_18013);
and UO_1324 (O_1324,N_18552,N_15488);
and UO_1325 (O_1325,N_15621,N_15276);
nor UO_1326 (O_1326,N_17606,N_17187);
nand UO_1327 (O_1327,N_19889,N_18882);
nand UO_1328 (O_1328,N_16722,N_16459);
and UO_1329 (O_1329,N_19537,N_15199);
or UO_1330 (O_1330,N_15804,N_19921);
xnor UO_1331 (O_1331,N_17651,N_18278);
nor UO_1332 (O_1332,N_17906,N_15909);
nand UO_1333 (O_1333,N_17536,N_18996);
and UO_1334 (O_1334,N_17595,N_16235);
nor UO_1335 (O_1335,N_16461,N_17122);
nand UO_1336 (O_1336,N_18991,N_15248);
nor UO_1337 (O_1337,N_15436,N_16370);
xnor UO_1338 (O_1338,N_18376,N_17912);
or UO_1339 (O_1339,N_19565,N_17251);
or UO_1340 (O_1340,N_19448,N_19396);
or UO_1341 (O_1341,N_18685,N_16152);
nor UO_1342 (O_1342,N_15289,N_17224);
or UO_1343 (O_1343,N_17634,N_17843);
and UO_1344 (O_1344,N_15609,N_18922);
and UO_1345 (O_1345,N_16354,N_16972);
and UO_1346 (O_1346,N_15095,N_15464);
and UO_1347 (O_1347,N_16750,N_15786);
or UO_1348 (O_1348,N_16435,N_17828);
nand UO_1349 (O_1349,N_19497,N_15291);
nand UO_1350 (O_1350,N_16083,N_17034);
nor UO_1351 (O_1351,N_19509,N_17890);
xnor UO_1352 (O_1352,N_19722,N_16588);
and UO_1353 (O_1353,N_16798,N_17375);
or UO_1354 (O_1354,N_15966,N_17937);
xor UO_1355 (O_1355,N_15778,N_19496);
nor UO_1356 (O_1356,N_19211,N_16645);
xnor UO_1357 (O_1357,N_16147,N_18125);
and UO_1358 (O_1358,N_15797,N_15748);
xnor UO_1359 (O_1359,N_15555,N_16058);
nand UO_1360 (O_1360,N_16336,N_15788);
nand UO_1361 (O_1361,N_16388,N_16988);
or UO_1362 (O_1362,N_19444,N_16660);
or UO_1363 (O_1363,N_17464,N_16762);
or UO_1364 (O_1364,N_16095,N_17437);
nor UO_1365 (O_1365,N_18806,N_16568);
nor UO_1366 (O_1366,N_17291,N_18570);
nand UO_1367 (O_1367,N_18883,N_17926);
or UO_1368 (O_1368,N_15050,N_15779);
and UO_1369 (O_1369,N_17097,N_16986);
nor UO_1370 (O_1370,N_16795,N_16966);
nand UO_1371 (O_1371,N_16962,N_15482);
xnor UO_1372 (O_1372,N_15819,N_19499);
nand UO_1373 (O_1373,N_17995,N_15974);
nor UO_1374 (O_1374,N_15270,N_18561);
and UO_1375 (O_1375,N_15101,N_17206);
nand UO_1376 (O_1376,N_15448,N_17124);
nor UO_1377 (O_1377,N_19791,N_18898);
and UO_1378 (O_1378,N_19707,N_18187);
and UO_1379 (O_1379,N_16053,N_15903);
or UO_1380 (O_1380,N_19760,N_18928);
or UO_1381 (O_1381,N_16020,N_18232);
or UO_1382 (O_1382,N_19335,N_15878);
nor UO_1383 (O_1383,N_18527,N_18642);
or UO_1384 (O_1384,N_17680,N_16505);
nand UO_1385 (O_1385,N_15986,N_16033);
nand UO_1386 (O_1386,N_18046,N_19734);
and UO_1387 (O_1387,N_17449,N_15764);
nand UO_1388 (O_1388,N_19084,N_19230);
nor UO_1389 (O_1389,N_17273,N_19790);
and UO_1390 (O_1390,N_16206,N_19233);
and UO_1391 (O_1391,N_19096,N_17924);
xor UO_1392 (O_1392,N_18169,N_18054);
xnor UO_1393 (O_1393,N_17899,N_19172);
or UO_1394 (O_1394,N_19617,N_17667);
xnor UO_1395 (O_1395,N_17686,N_16473);
nand UO_1396 (O_1396,N_16587,N_18413);
xnor UO_1397 (O_1397,N_17744,N_16268);
or UO_1398 (O_1398,N_16593,N_18490);
xor UO_1399 (O_1399,N_17520,N_19377);
nor UO_1400 (O_1400,N_15333,N_16500);
or UO_1401 (O_1401,N_17689,N_19359);
nor UO_1402 (O_1402,N_18364,N_17017);
nor UO_1403 (O_1403,N_16343,N_15088);
nand UO_1404 (O_1404,N_15465,N_16909);
nor UO_1405 (O_1405,N_17672,N_18576);
and UO_1406 (O_1406,N_15702,N_15266);
or UO_1407 (O_1407,N_18151,N_19078);
xnor UO_1408 (O_1408,N_17665,N_16964);
or UO_1409 (O_1409,N_15962,N_16443);
xor UO_1410 (O_1410,N_16785,N_15660);
and UO_1411 (O_1411,N_17889,N_16938);
nor UO_1412 (O_1412,N_17772,N_17090);
nor UO_1413 (O_1413,N_19234,N_18059);
nand UO_1414 (O_1414,N_16840,N_17888);
and UO_1415 (O_1415,N_19046,N_18163);
nand UO_1416 (O_1416,N_19778,N_17305);
or UO_1417 (O_1417,N_17053,N_15167);
and UO_1418 (O_1418,N_18090,N_18667);
xor UO_1419 (O_1419,N_15351,N_18772);
or UO_1420 (O_1420,N_15412,N_16699);
or UO_1421 (O_1421,N_17429,N_18513);
xnor UO_1422 (O_1422,N_19880,N_15062);
nand UO_1423 (O_1423,N_15635,N_19723);
and UO_1424 (O_1424,N_19765,N_15739);
nand UO_1425 (O_1425,N_16623,N_18637);
nand UO_1426 (O_1426,N_17261,N_18206);
or UO_1427 (O_1427,N_18751,N_19142);
nand UO_1428 (O_1428,N_16855,N_16615);
and UO_1429 (O_1429,N_16625,N_17628);
nor UO_1430 (O_1430,N_17702,N_16721);
and UO_1431 (O_1431,N_19367,N_15571);
or UO_1432 (O_1432,N_16021,N_16283);
xor UO_1433 (O_1433,N_19088,N_16208);
nand UO_1434 (O_1434,N_18482,N_18464);
and UO_1435 (O_1435,N_18858,N_18571);
nand UO_1436 (O_1436,N_15664,N_17991);
nand UO_1437 (O_1437,N_19714,N_15255);
nor UO_1438 (O_1438,N_16787,N_18353);
nand UO_1439 (O_1439,N_15950,N_18210);
nor UO_1440 (O_1440,N_16716,N_18378);
nor UO_1441 (O_1441,N_19337,N_18835);
nand UO_1442 (O_1442,N_15860,N_16048);
and UO_1443 (O_1443,N_19170,N_16504);
nand UO_1444 (O_1444,N_16939,N_17024);
or UO_1445 (O_1445,N_19761,N_18673);
xnor UO_1446 (O_1446,N_16888,N_15078);
xor UO_1447 (O_1447,N_18069,N_19855);
xnor UO_1448 (O_1448,N_15714,N_16457);
nor UO_1449 (O_1449,N_19399,N_18127);
and UO_1450 (O_1450,N_16323,N_15253);
and UO_1451 (O_1451,N_15472,N_15281);
or UO_1452 (O_1452,N_18136,N_17562);
and UO_1453 (O_1453,N_16211,N_15758);
xor UO_1454 (O_1454,N_17130,N_17099);
nor UO_1455 (O_1455,N_15182,N_17335);
nor UO_1456 (O_1456,N_16709,N_15548);
nor UO_1457 (O_1457,N_15939,N_17697);
or UO_1458 (O_1458,N_15093,N_18313);
nand UO_1459 (O_1459,N_19504,N_19764);
nand UO_1460 (O_1460,N_16533,N_16049);
and UO_1461 (O_1461,N_17088,N_15810);
nand UO_1462 (O_1462,N_18003,N_17543);
nor UO_1463 (O_1463,N_16835,N_18522);
and UO_1464 (O_1464,N_15186,N_18999);
or UO_1465 (O_1465,N_17771,N_16280);
xnor UO_1466 (O_1466,N_16713,N_15588);
xor UO_1467 (O_1467,N_16940,N_15603);
xnor UO_1468 (O_1468,N_17213,N_15558);
or UO_1469 (O_1469,N_18891,N_18213);
xor UO_1470 (O_1470,N_16513,N_15037);
or UO_1471 (O_1471,N_18736,N_15718);
or UO_1472 (O_1472,N_17831,N_15912);
and UO_1473 (O_1473,N_18212,N_17705);
or UO_1474 (O_1474,N_19689,N_19302);
nor UO_1475 (O_1475,N_16979,N_16805);
nand UO_1476 (O_1476,N_19494,N_16387);
nand UO_1477 (O_1477,N_17202,N_17244);
nand UO_1478 (O_1478,N_19644,N_16014);
nor UO_1479 (O_1479,N_17423,N_19814);
and UO_1480 (O_1480,N_17366,N_19387);
nand UO_1481 (O_1481,N_16641,N_18987);
nor UO_1482 (O_1482,N_16973,N_15535);
or UO_1483 (O_1483,N_19041,N_19110);
nand UO_1484 (O_1484,N_15074,N_18383);
nand UO_1485 (O_1485,N_18101,N_15457);
nor UO_1486 (O_1486,N_15385,N_19869);
nand UO_1487 (O_1487,N_16209,N_18336);
or UO_1488 (O_1488,N_18671,N_19116);
or UO_1489 (O_1489,N_19711,N_18328);
nand UO_1490 (O_1490,N_18318,N_19174);
nand UO_1491 (O_1491,N_15848,N_16253);
nor UO_1492 (O_1492,N_19528,N_17570);
or UO_1493 (O_1493,N_17189,N_17085);
or UO_1494 (O_1494,N_16175,N_17331);
and UO_1495 (O_1495,N_15813,N_19772);
nand UO_1496 (O_1496,N_16919,N_17792);
nand UO_1497 (O_1497,N_19651,N_18725);
xnor UO_1498 (O_1498,N_19585,N_17112);
or UO_1499 (O_1499,N_16160,N_15947);
nand UO_1500 (O_1500,N_17927,N_16788);
xnor UO_1501 (O_1501,N_18583,N_17825);
xnor UO_1502 (O_1502,N_15887,N_17814);
or UO_1503 (O_1503,N_17967,N_17474);
nand UO_1504 (O_1504,N_15812,N_18437);
and UO_1505 (O_1505,N_17293,N_18892);
xnor UO_1506 (O_1506,N_16736,N_17243);
xor UO_1507 (O_1507,N_18708,N_15407);
nor UO_1508 (O_1508,N_15362,N_16302);
nand UO_1509 (O_1509,N_18965,N_16971);
nand UO_1510 (O_1510,N_15671,N_17508);
nand UO_1511 (O_1511,N_16164,N_18629);
or UO_1512 (O_1512,N_18426,N_19586);
xor UO_1513 (O_1513,N_19757,N_15272);
nor UO_1514 (O_1514,N_18056,N_15469);
xor UO_1515 (O_1515,N_15940,N_18832);
nor UO_1516 (O_1516,N_15904,N_18770);
xor UO_1517 (O_1517,N_15982,N_17456);
nand UO_1518 (O_1518,N_18031,N_16554);
and UO_1519 (O_1519,N_16782,N_16328);
and UO_1520 (O_1520,N_15608,N_19892);
nand UO_1521 (O_1521,N_18823,N_19346);
nor UO_1522 (O_1522,N_16346,N_15769);
xnor UO_1523 (O_1523,N_15326,N_17173);
nand UO_1524 (O_1524,N_19634,N_19787);
nor UO_1525 (O_1525,N_18192,N_16285);
xor UO_1526 (O_1526,N_18432,N_17929);
and UO_1527 (O_1527,N_16779,N_19602);
and UO_1528 (O_1528,N_17941,N_16306);
nand UO_1529 (O_1529,N_19200,N_19515);
xor UO_1530 (O_1530,N_16893,N_17743);
nand UO_1531 (O_1531,N_15082,N_19020);
xnor UO_1532 (O_1532,N_18818,N_16176);
and UO_1533 (O_1533,N_19098,N_15553);
and UO_1534 (O_1534,N_16635,N_19986);
or UO_1535 (O_1535,N_17314,N_16953);
nor UO_1536 (O_1536,N_18348,N_18621);
nand UO_1537 (O_1537,N_15979,N_18186);
nor UO_1538 (O_1538,N_16054,N_18958);
nor UO_1539 (O_1539,N_19519,N_15538);
and UO_1540 (O_1540,N_16441,N_19840);
nand UO_1541 (O_1541,N_19154,N_15862);
nor UO_1542 (O_1542,N_19418,N_19423);
nor UO_1543 (O_1543,N_19879,N_18960);
or UO_1544 (O_1544,N_19706,N_19675);
or UO_1545 (O_1545,N_18496,N_17387);
xnor UO_1546 (O_1546,N_17511,N_19017);
nor UO_1547 (O_1547,N_16853,N_16327);
nand UO_1548 (O_1548,N_19421,N_17394);
or UO_1549 (O_1549,N_17637,N_16812);
nor UO_1550 (O_1550,N_15991,N_16308);
or UO_1551 (O_1551,N_15648,N_16589);
nand UO_1552 (O_1552,N_18022,N_16740);
nor UO_1553 (O_1553,N_18530,N_19189);
xor UO_1554 (O_1554,N_16481,N_18599);
nand UO_1555 (O_1555,N_18534,N_19929);
and UO_1556 (O_1556,N_19700,N_18864);
or UO_1557 (O_1557,N_16602,N_17064);
and UO_1558 (O_1558,N_16948,N_15384);
or UO_1559 (O_1559,N_18435,N_18773);
and UO_1560 (O_1560,N_19431,N_18613);
and UO_1561 (O_1561,N_19205,N_15985);
and UO_1562 (O_1562,N_17302,N_17047);
nor UO_1563 (O_1563,N_19595,N_19937);
nand UO_1564 (O_1564,N_16912,N_17994);
nor UO_1565 (O_1565,N_18553,N_16872);
and UO_1566 (O_1566,N_16297,N_17248);
xor UO_1567 (O_1567,N_19727,N_16528);
nor UO_1568 (O_1568,N_18116,N_16210);
or UO_1569 (O_1569,N_16299,N_15195);
and UO_1570 (O_1570,N_17294,N_16136);
or UO_1571 (O_1571,N_17829,N_18117);
or UO_1572 (O_1572,N_18684,N_18647);
or UO_1573 (O_1573,N_19000,N_19521);
nand UO_1574 (O_1574,N_19620,N_19288);
and UO_1575 (O_1575,N_19267,N_16815);
or UO_1576 (O_1576,N_17799,N_18544);
and UO_1577 (O_1577,N_19752,N_17894);
or UO_1578 (O_1578,N_18558,N_16486);
or UO_1579 (O_1579,N_19864,N_16002);
nor UO_1580 (O_1580,N_15634,N_19165);
or UO_1581 (O_1581,N_16949,N_17215);
nor UO_1582 (O_1582,N_19043,N_16773);
xnor UO_1583 (O_1583,N_15936,N_19928);
or UO_1584 (O_1584,N_18689,N_19208);
nor UO_1585 (O_1585,N_15644,N_17524);
nand UO_1586 (O_1586,N_17541,N_15438);
nand UO_1587 (O_1587,N_16485,N_15081);
xor UO_1588 (O_1588,N_16572,N_15202);
nor UO_1589 (O_1589,N_17733,N_16977);
nand UO_1590 (O_1590,N_18893,N_15489);
nand UO_1591 (O_1591,N_17547,N_17444);
nor UO_1592 (O_1592,N_18500,N_17190);
xor UO_1593 (O_1593,N_15741,N_19570);
or UO_1594 (O_1594,N_18484,N_17079);
xnor UO_1595 (O_1595,N_19573,N_19082);
nand UO_1596 (O_1596,N_19204,N_15231);
xor UO_1597 (O_1597,N_17498,N_15829);
nor UO_1598 (O_1598,N_17810,N_18848);
or UO_1599 (O_1599,N_16527,N_18905);
and UO_1600 (O_1600,N_19875,N_17852);
and UO_1601 (O_1601,N_19001,N_18731);
nand UO_1602 (O_1602,N_15021,N_16618);
nand UO_1603 (O_1603,N_16751,N_17329);
xor UO_1604 (O_1604,N_17559,N_16374);
nand UO_1605 (O_1605,N_16668,N_18227);
nor UO_1606 (O_1606,N_18446,N_16412);
and UO_1607 (O_1607,N_18162,N_19446);
nand UO_1608 (O_1608,N_16478,N_18066);
nand UO_1609 (O_1609,N_18008,N_15262);
or UO_1610 (O_1610,N_18471,N_15450);
or UO_1611 (O_1611,N_15219,N_15139);
xor UO_1612 (O_1612,N_18224,N_19594);
or UO_1613 (O_1613,N_19918,N_15268);
xnor UO_1614 (O_1614,N_19957,N_17722);
nand UO_1615 (O_1615,N_19319,N_19806);
or UO_1616 (O_1616,N_18043,N_15174);
or UO_1617 (O_1617,N_19792,N_17154);
xnor UO_1618 (O_1618,N_15370,N_15942);
xnor UO_1619 (O_1619,N_18573,N_17354);
and UO_1620 (O_1620,N_16034,N_16640);
or UO_1621 (O_1621,N_16445,N_16838);
and UO_1622 (O_1622,N_19376,N_18901);
nand UO_1623 (O_1623,N_15394,N_19316);
xor UO_1624 (O_1624,N_15990,N_16167);
nand UO_1625 (O_1625,N_19242,N_15150);
xor UO_1626 (O_1626,N_15389,N_19464);
xor UO_1627 (O_1627,N_17658,N_18501);
and UO_1628 (O_1628,N_17368,N_19693);
nor UO_1629 (O_1629,N_17420,N_18872);
and UO_1630 (O_1630,N_17790,N_19075);
or UO_1631 (O_1631,N_15600,N_18397);
and UO_1632 (O_1632,N_18266,N_18512);
nor UO_1633 (O_1633,N_16185,N_16832);
and UO_1634 (O_1634,N_19432,N_16356);
nand UO_1635 (O_1635,N_18158,N_17263);
or UO_1636 (O_1636,N_17106,N_18866);
or UO_1637 (O_1637,N_15752,N_19794);
nor UO_1638 (O_1638,N_15129,N_16705);
nand UO_1639 (O_1639,N_18494,N_19505);
and UO_1640 (O_1640,N_18757,N_15627);
or UO_1641 (O_1641,N_18103,N_15245);
or UO_1642 (O_1642,N_15179,N_15885);
xor UO_1643 (O_1643,N_15689,N_17083);
and UO_1644 (O_1644,N_19384,N_19053);
nand UO_1645 (O_1645,N_17289,N_18735);
and UO_1646 (O_1646,N_16376,N_19597);
nand UO_1647 (O_1647,N_16733,N_15367);
xnor UO_1648 (O_1648,N_15522,N_17847);
or UO_1649 (O_1649,N_15896,N_16111);
and UO_1650 (O_1650,N_17723,N_19933);
xnor UO_1651 (O_1651,N_18236,N_19236);
nand UO_1652 (O_1652,N_18195,N_18403);
xor UO_1653 (O_1653,N_17067,N_19811);
xor UO_1654 (O_1654,N_16286,N_16115);
nor UO_1655 (O_1655,N_15224,N_15864);
or UO_1656 (O_1656,N_18477,N_17066);
and UO_1657 (O_1657,N_18075,N_19627);
xor UO_1658 (O_1658,N_15137,N_15446);
nand UO_1659 (O_1659,N_17133,N_17489);
and UO_1660 (O_1660,N_19256,N_18913);
nand UO_1661 (O_1661,N_17431,N_19923);
or UO_1662 (O_1662,N_17412,N_18920);
or UO_1663 (O_1663,N_17082,N_19287);
nor UO_1664 (O_1664,N_17208,N_15723);
nand UO_1665 (O_1665,N_17253,N_16987);
xor UO_1666 (O_1666,N_19969,N_19101);
or UO_1667 (O_1667,N_17274,N_17597);
or UO_1668 (O_1668,N_18656,N_15247);
and UO_1669 (O_1669,N_17483,N_16860);
and UO_1670 (O_1670,N_17388,N_16741);
xor UO_1671 (O_1671,N_16869,N_19122);
and UO_1672 (O_1672,N_18188,N_18012);
nand UO_1673 (O_1673,N_15210,N_18983);
xnor UO_1674 (O_1674,N_17897,N_19087);
nor UO_1675 (O_1675,N_18620,N_16032);
or UO_1676 (O_1676,N_16367,N_16725);
and UO_1677 (O_1677,N_15978,N_19618);
xnor UO_1678 (O_1678,N_19945,N_16186);
nand UO_1679 (O_1679,N_18058,N_15391);
nand UO_1680 (O_1680,N_16524,N_15443);
nand UO_1681 (O_1681,N_17989,N_18862);
or UO_1682 (O_1682,N_15144,N_15188);
xnor UO_1683 (O_1683,N_19054,N_17033);
xnor UO_1684 (O_1684,N_17249,N_18903);
nor UO_1685 (O_1685,N_19193,N_15856);
xnor UO_1686 (O_1686,N_17655,N_17978);
nor UO_1687 (O_1687,N_19326,N_16873);
nor UO_1688 (O_1688,N_19652,N_18064);
or UO_1689 (O_1689,N_17736,N_16693);
nand UO_1690 (O_1690,N_17113,N_17409);
nor UO_1691 (O_1691,N_18366,N_19016);
nor UO_1692 (O_1692,N_18575,N_16202);
and UO_1693 (O_1693,N_15894,N_17275);
and UO_1694 (O_1694,N_17527,N_19695);
or UO_1695 (O_1695,N_16358,N_17664);
or UO_1696 (O_1696,N_19420,N_17299);
or UO_1697 (O_1697,N_16287,N_15715);
xor UO_1698 (O_1698,N_15639,N_16398);
or UO_1699 (O_1699,N_19870,N_18453);
nand UO_1700 (O_1700,N_19411,N_19717);
nor UO_1701 (O_1701,N_18220,N_15928);
and UO_1702 (O_1702,N_19800,N_16647);
or UO_1703 (O_1703,N_15145,N_17194);
and UO_1704 (O_1704,N_17358,N_15171);
and UO_1705 (O_1705,N_17676,N_15937);
xor UO_1706 (O_1706,N_16201,N_19645);
and UO_1707 (O_1707,N_18798,N_15881);
xor UO_1708 (O_1708,N_16963,N_18769);
or UO_1709 (O_1709,N_16284,N_18302);
or UO_1710 (O_1710,N_19272,N_15159);
or UO_1711 (O_1711,N_18815,N_16003);
or UO_1712 (O_1712,N_15584,N_18653);
xor UO_1713 (O_1713,N_18914,N_19203);
nor UO_1714 (O_1714,N_16697,N_18543);
and UO_1715 (O_1715,N_18919,N_19152);
or UO_1716 (O_1716,N_15771,N_18896);
nor UO_1717 (O_1717,N_15921,N_16067);
nor UO_1718 (O_1718,N_15451,N_18294);
or UO_1719 (O_1719,N_19097,N_19967);
nand UO_1720 (O_1720,N_19829,N_17371);
xnor UO_1721 (O_1721,N_19226,N_15729);
and UO_1722 (O_1722,N_16495,N_18021);
or UO_1723 (O_1723,N_18511,N_16071);
nor UO_1724 (O_1724,N_15502,N_17198);
and UO_1725 (O_1725,N_17128,N_18265);
and UO_1726 (O_1726,N_15056,N_18316);
nor UO_1727 (O_1727,N_15847,N_18094);
nand UO_1728 (O_1728,N_17955,N_15888);
nand UO_1729 (O_1729,N_19655,N_18797);
xnor UO_1730 (O_1730,N_16419,N_16100);
nand UO_1731 (O_1731,N_16255,N_18661);
nand UO_1732 (O_1732,N_16460,N_17546);
xor UO_1733 (O_1733,N_19844,N_16322);
and UO_1734 (O_1734,N_16626,N_15028);
or UO_1735 (O_1735,N_16446,N_15261);
and UO_1736 (O_1736,N_18504,N_18949);
xor UO_1737 (O_1737,N_17583,N_16468);
or UO_1738 (O_1738,N_19514,N_16366);
or UO_1739 (O_1739,N_15698,N_16004);
or UO_1740 (O_1740,N_15218,N_16458);
xor UO_1741 (O_1741,N_16555,N_19533);
nor UO_1742 (O_1742,N_15052,N_16163);
nand UO_1743 (O_1743,N_15516,N_19275);
xnor UO_1744 (O_1744,N_19102,N_18382);
and UO_1745 (O_1745,N_15290,N_17357);
nor UO_1746 (O_1746,N_15035,N_18998);
xor UO_1747 (O_1747,N_18408,N_16531);
and UO_1748 (O_1748,N_19018,N_18780);
nor UO_1749 (O_1749,N_15136,N_16470);
nor UO_1750 (O_1750,N_16799,N_16187);
or UO_1751 (O_1751,N_15109,N_19834);
xnor UO_1752 (O_1752,N_15205,N_19013);
and UO_1753 (O_1753,N_18924,N_19522);
nor UO_1754 (O_1754,N_19108,N_19951);
or UO_1755 (O_1755,N_18837,N_19149);
nand UO_1756 (O_1756,N_17247,N_16534);
xnor UO_1757 (O_1757,N_19915,N_15839);
nor UO_1758 (O_1758,N_16425,N_19114);
nor UO_1759 (O_1759,N_18457,N_16599);
nand UO_1760 (O_1760,N_17451,N_18201);
or UO_1761 (O_1761,N_15161,N_19456);
and UO_1762 (O_1762,N_16247,N_18436);
and UO_1763 (O_1763,N_17142,N_15514);
or UO_1764 (O_1764,N_18081,N_18935);
nor UO_1765 (O_1765,N_17376,N_15633);
xor UO_1766 (O_1766,N_19292,N_19562);
xnor UO_1767 (O_1767,N_18895,N_15316);
xor UO_1768 (O_1768,N_16737,N_17374);
nand UO_1769 (O_1769,N_17604,N_18861);
nand UO_1770 (O_1770,N_18515,N_17858);
nand UO_1771 (O_1771,N_17013,N_18352);
xnor UO_1772 (O_1772,N_16183,N_18466);
nand UO_1773 (O_1773,N_18927,N_17092);
or UO_1774 (O_1774,N_15557,N_19179);
xor UO_1775 (O_1775,N_19922,N_16564);
nor UO_1776 (O_1776,N_17238,N_17148);
and UO_1777 (O_1777,N_16603,N_15500);
xor UO_1778 (O_1778,N_15342,N_16169);
or UO_1779 (O_1779,N_18198,N_16598);
or UO_1780 (O_1780,N_16407,N_19525);
or UO_1781 (O_1781,N_17749,N_19286);
nor UO_1782 (O_1782,N_18126,N_18979);
xor UO_1783 (O_1783,N_19040,N_19198);
and UO_1784 (O_1784,N_18717,N_18776);
nor UO_1785 (O_1785,N_15474,N_18060);
and UO_1786 (O_1786,N_18238,N_19157);
nor UO_1787 (O_1787,N_17730,N_15418);
or UO_1788 (O_1788,N_16883,N_15068);
nor UO_1789 (O_1789,N_16558,N_19015);
xor UO_1790 (O_1790,N_17181,N_16511);
nor UO_1791 (O_1791,N_16530,N_18700);
and UO_1792 (O_1792,N_18137,N_19683);
nand UO_1793 (O_1793,N_19755,N_17192);
and UO_1794 (O_1794,N_17492,N_17091);
xnor UO_1795 (O_1795,N_16292,N_15143);
xor UO_1796 (O_1796,N_16226,N_19983);
xor UO_1797 (O_1797,N_18778,N_17751);
nor UO_1798 (O_1798,N_19210,N_19197);
xnor UO_1799 (O_1799,N_17633,N_17973);
xor UO_1800 (O_1800,N_16902,N_15397);
nor UO_1801 (O_1801,N_17041,N_17363);
and UO_1802 (O_1802,N_16015,N_17486);
nor UO_1803 (O_1803,N_15330,N_17526);
and UO_1804 (O_1804,N_16634,N_19414);
and UO_1805 (O_1805,N_17333,N_18200);
xnor UO_1806 (O_1806,N_15003,N_15767);
and UO_1807 (O_1807,N_16170,N_16706);
nand UO_1808 (O_1808,N_17407,N_16884);
nor UO_1809 (O_1809,N_19697,N_18000);
nor UO_1810 (O_1810,N_16137,N_17227);
or UO_1811 (O_1811,N_16562,N_19477);
nand UO_1812 (O_1812,N_15173,N_17369);
and UO_1813 (O_1813,N_17328,N_19662);
nand UO_1814 (O_1814,N_19145,N_17950);
and UO_1815 (O_1815,N_15244,N_15653);
or UO_1816 (O_1816,N_16394,N_15026);
and UO_1817 (O_1817,N_17734,N_17170);
or UO_1818 (O_1818,N_16661,N_16596);
and UO_1819 (O_1819,N_18784,N_19403);
nor UO_1820 (O_1820,N_18488,N_16637);
nand UO_1821 (O_1821,N_17062,N_19104);
nand UO_1822 (O_1822,N_18582,N_18767);
nor UO_1823 (O_1823,N_15258,N_18733);
xnor UO_1824 (O_1824,N_18281,N_17025);
xnor UO_1825 (O_1825,N_18686,N_19953);
nor UO_1826 (O_1826,N_17688,N_17162);
nor UO_1827 (O_1827,N_18675,N_17840);
nand UO_1828 (O_1828,N_19148,N_19038);
xor UO_1829 (O_1829,N_17811,N_15386);
nor UO_1830 (O_1830,N_18825,N_17297);
nand UO_1831 (O_1831,N_17071,N_19629);
or UO_1832 (O_1832,N_16159,N_18646);
and UO_1833 (O_1833,N_17089,N_19783);
nand UO_1834 (O_1834,N_19437,N_15983);
nor UO_1835 (O_1835,N_16876,N_15919);
xor UO_1836 (O_1836,N_19774,N_18329);
or UO_1837 (O_1837,N_19735,N_15612);
xnor UO_1838 (O_1838,N_16207,N_17022);
or UO_1839 (O_1839,N_19981,N_18027);
nor UO_1840 (O_1840,N_15520,N_18157);
xnor UO_1841 (O_1841,N_18241,N_19443);
or UO_1842 (O_1842,N_15408,N_17397);
nand UO_1843 (O_1843,N_16091,N_15031);
or UO_1844 (O_1844,N_16082,N_15737);
or UO_1845 (O_1845,N_19398,N_17646);
or UO_1846 (O_1846,N_16745,N_19579);
nand UO_1847 (O_1847,N_16112,N_17964);
or UO_1848 (O_1848,N_16291,N_15141);
xor UO_1849 (O_1849,N_16055,N_16717);
or UO_1850 (O_1850,N_17704,N_17121);
and UO_1851 (O_1851,N_17072,N_17842);
or UO_1852 (O_1852,N_18638,N_19646);
xnor UO_1853 (O_1853,N_15798,N_19331);
and UO_1854 (O_1854,N_19987,N_15837);
nor UO_1855 (O_1855,N_15131,N_18904);
xor UO_1856 (O_1856,N_15356,N_18591);
nand UO_1857 (O_1857,N_17981,N_15735);
nand UO_1858 (O_1858,N_19067,N_15410);
nor UO_1859 (O_1859,N_17266,N_18771);
xor UO_1860 (O_1860,N_16007,N_18433);
and UO_1861 (O_1861,N_19325,N_16024);
or UO_1862 (O_1862,N_17820,N_19539);
xor UO_1863 (O_1863,N_15799,N_17678);
xnor UO_1864 (O_1864,N_19370,N_17324);
nand UO_1865 (O_1865,N_16989,N_16525);
nor UO_1866 (O_1866,N_19773,N_17012);
or UO_1867 (O_1867,N_17904,N_15286);
and UO_1868 (O_1868,N_18917,N_18038);
and UO_1869 (O_1869,N_18130,N_19371);
nor UO_1870 (O_1870,N_18486,N_19666);
xnor UO_1871 (O_1871,N_15958,N_19810);
nor UO_1872 (O_1872,N_17862,N_18678);
or UO_1873 (O_1873,N_19660,N_15360);
nand UO_1874 (O_1874,N_16451,N_17795);
nor UO_1875 (O_1875,N_18524,N_15880);
xnor UO_1876 (O_1876,N_17094,N_17149);
and UO_1877 (O_1877,N_19330,N_15933);
nor UO_1878 (O_1878,N_18016,N_16197);
nor UO_1879 (O_1879,N_16415,N_18310);
or UO_1880 (O_1880,N_15897,N_16496);
nand UO_1881 (O_1881,N_16344,N_17468);
or UO_1882 (O_1882,N_16559,N_18586);
xnor UO_1883 (O_1883,N_15733,N_19360);
nand UO_1884 (O_1884,N_16752,N_18095);
nor UO_1885 (O_1885,N_17874,N_19581);
or UO_1886 (O_1886,N_15582,N_18517);
or UO_1887 (O_1887,N_16692,N_16440);
nor UO_1888 (O_1888,N_18666,N_15228);
or UO_1889 (O_1889,N_17776,N_18783);
or UO_1890 (O_1890,N_17430,N_15094);
nand UO_1891 (O_1891,N_17871,N_15341);
nand UO_1892 (O_1892,N_19851,N_15575);
nand UO_1893 (O_1893,N_19358,N_16305);
and UO_1894 (O_1894,N_16870,N_17159);
xnor UO_1895 (O_1895,N_17327,N_18114);
xor UO_1896 (O_1896,N_17726,N_17643);
nand UO_1897 (O_1897,N_16767,N_18042);
nor UO_1898 (O_1898,N_15772,N_19857);
nor UO_1899 (O_1899,N_18946,N_16377);
or UO_1900 (O_1900,N_19350,N_17174);
or UO_1901 (O_1901,N_15221,N_19563);
nor UO_1902 (O_1902,N_16320,N_18249);
xnor UO_1903 (O_1903,N_15701,N_18167);
nand UO_1904 (O_1904,N_18662,N_15175);
nor UO_1905 (O_1905,N_19822,N_16996);
xnor UO_1906 (O_1906,N_16373,N_18940);
nor UO_1907 (O_1907,N_16846,N_16104);
nand UO_1908 (O_1908,N_19357,N_15964);
nand UO_1909 (O_1909,N_19917,N_18473);
nand UO_1910 (O_1910,N_16217,N_17283);
nand UO_1911 (O_1911,N_18180,N_17078);
and UO_1912 (O_1912,N_17758,N_16464);
nand UO_1913 (O_1913,N_16089,N_19530);
xnor UO_1914 (O_1914,N_17598,N_19462);
or UO_1915 (O_1915,N_15423,N_18803);
xor UO_1916 (O_1916,N_16816,N_15123);
nor UO_1917 (O_1917,N_15431,N_15759);
or UO_1918 (O_1918,N_16062,N_18521);
xnor UO_1919 (O_1919,N_18879,N_17399);
or UO_1920 (O_1920,N_18253,N_16514);
xnor UO_1921 (O_1921,N_15865,N_15827);
nand UO_1922 (O_1922,N_18168,N_17280);
and UO_1923 (O_1923,N_19243,N_16403);
nand UO_1924 (O_1924,N_16411,N_18749);
nand UO_1925 (O_1925,N_15930,N_19391);
xnor UO_1926 (O_1926,N_17601,N_17635);
or UO_1927 (O_1927,N_16681,N_18052);
nand UO_1928 (O_1928,N_19194,N_15456);
or UO_1929 (O_1929,N_16223,N_15970);
or UO_1930 (O_1930,N_18831,N_17677);
nand UO_1931 (O_1931,N_19511,N_15580);
nor UO_1932 (O_1932,N_16409,N_18284);
nand UO_1933 (O_1933,N_15800,N_17393);
nor UO_1934 (O_1934,N_15527,N_17235);
xnor UO_1935 (O_1935,N_19469,N_19746);
and UO_1936 (O_1936,N_15072,N_18750);
xor UO_1937 (O_1937,N_16391,N_15891);
nor UO_1938 (O_1938,N_15871,N_15063);
nor UO_1939 (O_1939,N_18235,N_16903);
xnor UO_1940 (O_1940,N_16930,N_18792);
nand UO_1941 (O_1941,N_18209,N_15240);
nand UO_1942 (O_1942,N_17232,N_15613);
nand UO_1943 (O_1943,N_17893,N_15883);
nor UO_1944 (O_1944,N_18147,N_18814);
or UO_1945 (O_1945,N_17602,N_16278);
or UO_1946 (O_1946,N_19133,N_17652);
nor UO_1947 (O_1947,N_15545,N_18768);
nor UO_1948 (O_1948,N_19972,N_16006);
nor UO_1949 (O_1949,N_19635,N_15498);
or UO_1950 (O_1950,N_15017,N_15703);
nand UO_1951 (O_1951,N_18349,N_18507);
or UO_1952 (O_1952,N_17621,N_17512);
or UO_1953 (O_1953,N_17614,N_17819);
xnor UO_1954 (O_1954,N_17039,N_17808);
or UO_1955 (O_1955,N_19715,N_15916);
and UO_1956 (O_1956,N_16070,N_16772);
and UO_1957 (O_1957,N_19710,N_18106);
xor UO_1958 (O_1958,N_15616,N_15406);
nand UO_1959 (O_1959,N_17011,N_19853);
xor UO_1960 (O_1960,N_15505,N_16842);
or UO_1961 (O_1961,N_19665,N_16277);
and UO_1962 (O_1962,N_17979,N_18853);
nor UO_1963 (O_1963,N_19263,N_17623);
or UO_1964 (O_1964,N_19389,N_15039);
nand UO_1965 (O_1965,N_18156,N_19249);
nand UO_1966 (O_1966,N_17816,N_18208);
or UO_1967 (O_1967,N_15740,N_18909);
nor UO_1968 (O_1968,N_18423,N_18185);
and UO_1969 (O_1969,N_18759,N_19621);
and UO_1970 (O_1970,N_19679,N_16836);
or UO_1971 (O_1971,N_18793,N_17882);
or UO_1972 (O_1972,N_17784,N_18089);
or UO_1973 (O_1973,N_18288,N_15380);
xnor UO_1974 (O_1974,N_18240,N_18874);
or UO_1975 (O_1975,N_16270,N_15935);
nand UO_1976 (O_1976,N_17105,N_17966);
or UO_1977 (O_1977,N_19354,N_16395);
nor UO_1978 (O_1978,N_17245,N_18925);
xor UO_1979 (O_1979,N_15624,N_19333);
or UO_1980 (O_1980,N_19520,N_17036);
xor UO_1981 (O_1981,N_18966,N_17530);
nand UO_1982 (O_1982,N_15250,N_17454);
and UO_1983 (O_1983,N_15083,N_17146);
or UO_1984 (O_1984,N_16567,N_17896);
and UO_1985 (O_1985,N_18369,N_16309);
nand UO_1986 (O_1986,N_17257,N_19979);
nor UO_1987 (O_1987,N_16648,N_19990);
and UO_1988 (O_1988,N_18110,N_19718);
nand UO_1989 (O_1989,N_18304,N_18063);
xor UO_1990 (O_1990,N_15416,N_19118);
xor UO_1991 (O_1991,N_18388,N_17499);
xor UO_1992 (O_1992,N_16542,N_17040);
or UO_1993 (O_1993,N_16509,N_15098);
nor UO_1994 (O_1994,N_17139,N_18421);
and UO_1995 (O_1995,N_19487,N_16823);
or UO_1996 (O_1996,N_16659,N_15844);
or UO_1997 (O_1997,N_17533,N_17729);
or UO_1998 (O_1998,N_18627,N_19027);
and UO_1999 (O_1999,N_18202,N_17848);
xnor UO_2000 (O_2000,N_15163,N_19225);
xnor UO_2001 (O_2001,N_19891,N_16849);
or UO_2002 (O_2002,N_18813,N_15198);
nor UO_2003 (O_2003,N_15724,N_15010);
nand UO_2004 (O_2004,N_16652,N_18338);
or UO_2005 (O_2005,N_15959,N_18568);
and UO_2006 (O_2006,N_17421,N_15241);
nor UO_2007 (O_2007,N_15057,N_19846);
or UO_2008 (O_2008,N_19538,N_15853);
or UO_2009 (O_2009,N_19687,N_17491);
nand UO_2010 (O_2010,N_15147,N_18624);
xnor UO_2011 (O_2011,N_17584,N_15015);
xor UO_2012 (O_2012,N_19474,N_17641);
or UO_2013 (O_2013,N_15625,N_16578);
nand UO_2014 (O_2014,N_18142,N_19324);
xnor UO_2015 (O_2015,N_16143,N_19277);
and UO_2016 (O_2016,N_18239,N_17916);
nand UO_2017 (O_2017,N_16882,N_19613);
or UO_2018 (O_2018,N_17608,N_15900);
nor UO_2019 (O_2019,N_18165,N_17043);
and UO_2020 (O_2020,N_18974,N_15814);
or UO_2021 (O_2021,N_18153,N_17708);
or UO_2022 (O_2022,N_17487,N_19908);
or UO_2023 (O_2023,N_18714,N_15628);
and UO_2024 (O_2024,N_17638,N_19274);
xnor UO_2025 (O_2025,N_18461,N_19865);
xnor UO_2026 (O_2026,N_19768,N_16581);
nand UO_2027 (O_2027,N_17204,N_19169);
or UO_2028 (O_2028,N_19103,N_18222);
nand UO_2029 (O_2029,N_19182,N_19954);
nor UO_2030 (O_2030,N_19453,N_17909);
or UO_2031 (O_2031,N_18080,N_19112);
xnor UO_2032 (O_2032,N_19386,N_18380);
or UO_2033 (O_2033,N_17907,N_17519);
nand UO_2034 (O_2034,N_16946,N_17865);
or UO_2035 (O_2035,N_17653,N_19930);
and UO_2036 (O_2036,N_19280,N_16726);
nor UO_2037 (O_2037,N_19308,N_16880);
nand UO_2038 (O_2038,N_16730,N_15796);
nor UO_2039 (O_2039,N_15876,N_15794);
nor UO_2040 (O_2040,N_16406,N_16824);
nand UO_2041 (O_2041,N_17390,N_19490);
and UO_2042 (O_2042,N_16595,N_16867);
xor UO_2043 (O_2043,N_15954,N_15944);
nor UO_2044 (O_2044,N_19057,N_18299);
nand UO_2045 (O_2045,N_18938,N_17140);
and UO_2046 (O_2046,N_16813,N_19105);
xnor UO_2047 (O_2047,N_16976,N_17721);
or UO_2048 (O_2048,N_16012,N_15721);
nor UO_2049 (O_2049,N_15999,N_17166);
nor UO_2050 (O_2050,N_16852,N_17100);
nand UO_2051 (O_2051,N_18256,N_17720);
nand UO_2052 (O_2052,N_17675,N_19374);
xor UO_2053 (O_2053,N_15206,N_15760);
xor UO_2054 (O_2054,N_17587,N_18867);
xnor UO_2055 (O_2055,N_17292,N_16047);
nor UO_2056 (O_2056,N_19803,N_16231);
xor UO_2057 (O_2057,N_16098,N_15949);
xnor UO_2058 (O_2058,N_17510,N_15917);
nor UO_2059 (O_2059,N_15857,N_16400);
nand UO_2060 (O_2060,N_17592,N_17381);
xor UO_2061 (O_2061,N_15670,N_19168);
nand UO_2062 (O_2062,N_16881,N_17622);
nor UO_2063 (O_2063,N_17349,N_17165);
xnor UO_2064 (O_2064,N_19920,N_17880);
and UO_2065 (O_2065,N_17359,N_16765);
and UO_2066 (O_2066,N_15743,N_19901);
or UO_2067 (O_2067,N_19202,N_19797);
nand UO_2068 (O_2068,N_15568,N_19066);
xnor UO_2069 (O_2069,N_16361,N_17764);
or UO_2070 (O_2070,N_18828,N_19980);
nor UO_2071 (O_2071,N_18100,N_17841);
and UO_2072 (O_2072,N_19138,N_16349);
xor UO_2073 (O_2073,N_17021,N_15791);
nor UO_2074 (O_2074,N_15783,N_16399);
and UO_2075 (O_2075,N_15578,N_18990);
nand UO_2076 (O_2076,N_18315,N_16418);
xnor UO_2077 (O_2077,N_17118,N_17323);
nand UO_2078 (O_2078,N_19798,N_15663);
xnor UO_2079 (O_2079,N_15103,N_17540);
xor UO_2080 (O_2080,N_16096,N_16700);
or UO_2081 (O_2081,N_18411,N_16430);
xnor UO_2082 (O_2082,N_16631,N_19852);
nand UO_2083 (O_2083,N_19368,N_15387);
and UO_2084 (O_2084,N_15453,N_15480);
or UO_2085 (O_2085,N_19583,N_19071);
xnor UO_2086 (O_2086,N_17834,N_18610);
xor UO_2087 (O_2087,N_16475,N_17377);
xor UO_2088 (O_2088,N_18807,N_18947);
nor UO_2089 (O_2089,N_15518,N_17876);
and UO_2090 (O_2090,N_19143,N_15806);
nand UO_2091 (O_2091,N_19452,N_15282);
nand UO_2092 (O_2092,N_19535,N_17320);
or UO_2093 (O_2093,N_15576,N_18010);
and UO_2094 (O_2094,N_17586,N_17553);
and UO_2095 (O_2095,N_16675,N_16613);
or UO_2096 (O_2096,N_15314,N_19279);
or UO_2097 (O_2097,N_18614,N_16866);
nand UO_2098 (O_2098,N_18385,N_15706);
nand UO_2099 (O_2099,N_16494,N_19095);
or UO_2100 (O_2100,N_15592,N_18789);
xor UO_2101 (O_2101,N_15761,N_18325);
xor UO_2102 (O_2102,N_16651,N_18261);
xnor UO_2103 (O_2103,N_18289,N_15941);
nor UO_2104 (O_2104,N_18677,N_17038);
or UO_2105 (O_2105,N_15156,N_18616);
nand UO_2106 (O_2106,N_15821,N_17117);
nand UO_2107 (O_2107,N_15476,N_19527);
and UO_2108 (O_2108,N_19843,N_18495);
nand UO_2109 (O_2109,N_16908,N_16863);
nor UO_2110 (O_2110,N_16576,N_19531);
xnor UO_2111 (O_2111,N_18096,N_15719);
nand UO_2112 (O_2112,N_19264,N_15524);
nand UO_2113 (O_2113,N_19328,N_16073);
nand UO_2114 (O_2114,N_19092,N_15546);
nand UO_2115 (O_2115,N_17642,N_15832);
nand UO_2116 (O_2116,N_16764,N_15494);
or UO_2117 (O_2117,N_19425,N_18523);
or UO_2118 (O_2118,N_15212,N_16099);
xnor UO_2119 (O_2119,N_16142,N_15298);
and UO_2120 (O_2120,N_16153,N_19285);
xor UO_2121 (O_2121,N_15170,N_18118);
nand UO_2122 (O_2122,N_17846,N_17827);
nand UO_2123 (O_2123,N_16097,N_15626);
nand UO_2124 (O_2124,N_15018,N_16687);
or UO_2125 (O_2125,N_18305,N_15924);
or UO_2126 (O_2126,N_19906,N_16279);
nand UO_2127 (O_2127,N_17793,N_19356);
and UO_2128 (O_2128,N_17529,N_17988);
or UO_2129 (O_2129,N_15181,N_18668);
nand UO_2130 (O_2130,N_15090,N_18268);
nand UO_2131 (O_2131,N_18345,N_19740);
and UO_2132 (O_2132,N_16897,N_18718);
nor UO_2133 (O_2133,N_17447,N_19218);
nand UO_2134 (O_2134,N_18878,N_16621);
xnor UO_2135 (O_2135,N_16891,N_18810);
nor UO_2136 (O_2136,N_15352,N_19426);
nor UO_2137 (O_2137,N_15594,N_19021);
or UO_2138 (O_2138,N_16895,N_16233);
nor UO_2139 (O_2139,N_17745,N_15736);
or UO_2140 (O_2140,N_18456,N_18705);
or UO_2141 (O_2141,N_17287,N_17182);
or UO_2142 (O_2142,N_16516,N_17781);
or UO_2143 (O_2143,N_18664,N_19947);
xor UO_2144 (O_2144,N_17537,N_17026);
nand UO_2145 (O_2145,N_15321,N_18333);
and UO_2146 (O_2146,N_16498,N_18332);
and UO_2147 (O_2147,N_16698,N_17259);
nand UO_2148 (O_2148,N_16570,N_18618);
or UO_2149 (O_2149,N_15222,N_18191);
xnor UO_2150 (O_2150,N_16942,N_15214);
nand UO_2151 (O_2151,N_19907,N_19014);
xor UO_2152 (O_2152,N_15707,N_19340);
xnor UO_2153 (O_2153,N_19442,N_18279);
or UO_2154 (O_2154,N_17785,N_16128);
or UO_2155 (O_2155,N_19838,N_18295);
and UO_2156 (O_2156,N_15085,N_19055);
or UO_2157 (O_2157,N_18841,N_18581);
or UO_2158 (O_2158,N_19926,N_18230);
or UO_2159 (O_2159,N_19006,N_19465);
nor UO_2160 (O_2160,N_15948,N_17201);
and UO_2161 (O_2161,N_15803,N_16035);
and UO_2162 (O_2162,N_15731,N_15611);
nor UO_2163 (O_2163,N_19762,N_19866);
nand UO_2164 (O_2164,N_19674,N_16410);
nor UO_2165 (O_2165,N_18148,N_17933);
or UO_2166 (O_2166,N_18554,N_15531);
and UO_2167 (O_2167,N_17639,N_19753);
and UO_2168 (O_2168,N_15793,N_18606);
xor UO_2169 (O_2169,N_19372,N_15845);
or UO_2170 (O_2170,N_17815,N_19996);
or UO_2171 (O_2171,N_19770,N_17006);
or UO_2172 (O_2172,N_16312,N_19518);
or UO_2173 (O_2173,N_18416,N_19609);
and UO_2174 (O_2174,N_17752,N_19180);
or UO_2175 (O_2175,N_18463,N_16384);
or UO_2176 (O_2176,N_16961,N_15732);
nand UO_2177 (O_2177,N_15146,N_18412);
xor UO_2178 (O_2178,N_16710,N_16654);
and UO_2179 (O_2179,N_16605,N_15526);
nor UO_2180 (O_2180,N_19187,N_18923);
xnor UO_2181 (O_2181,N_17443,N_17441);
or UO_2182 (O_2182,N_15677,N_18727);
nand UO_2183 (O_2183,N_19845,N_18254);
nor UO_2184 (O_2184,N_19167,N_18834);
nand UO_2185 (O_2185,N_18950,N_15691);
nand UO_2186 (O_2186,N_18608,N_18584);
and UO_2187 (O_2187,N_15425,N_17921);
nand UO_2188 (O_2188,N_16337,N_15230);
and UO_2189 (O_2189,N_16742,N_16702);
or UO_2190 (O_2190,N_16560,N_19973);
or UO_2191 (O_2191,N_17535,N_16290);
xor UO_2192 (O_2192,N_17544,N_17147);
or UO_2193 (O_2193,N_15044,N_19144);
or UO_2194 (O_2194,N_18592,N_15271);
and UO_2195 (O_2195,N_17384,N_17296);
and UO_2196 (O_2196,N_18121,N_16523);
and UO_2197 (O_2197,N_16078,N_15215);
and UO_2198 (O_2198,N_16543,N_18041);
and UO_2199 (O_2199,N_17396,N_15047);
nand UO_2200 (O_2200,N_18124,N_19348);
and UO_2201 (O_2201,N_19315,N_15157);
nor UO_2202 (O_2202,N_18589,N_18424);
or UO_2203 (O_2203,N_18067,N_18619);
and UO_2204 (O_2204,N_19025,N_19939);
and UO_2205 (O_2205,N_16540,N_17135);
nor UO_2206 (O_2206,N_17392,N_18514);
nor UO_2207 (O_2207,N_19962,N_16069);
nor UO_2208 (O_2208,N_17028,N_15452);
and UO_2209 (O_2209,N_16362,N_18645);
and UO_2210 (O_2210,N_18199,N_15777);
xor UO_2211 (O_2211,N_19672,N_15320);
nand UO_2212 (O_2212,N_15533,N_17385);
or UO_2213 (O_2213,N_15053,N_17205);
nand UO_2214 (O_2214,N_17822,N_17965);
nand UO_2215 (O_2215,N_16563,N_18161);
xnor UO_2216 (O_2216,N_15042,N_18255);
and UO_2217 (O_2217,N_19726,N_15307);
nand UO_2218 (O_2218,N_15898,N_15275);
nand UO_2219 (O_2219,N_15029,N_19369);
or UO_2220 (O_2220,N_19353,N_18108);
nand UO_2221 (O_2221,N_17919,N_18711);
and UO_2222 (O_2222,N_19608,N_16653);
nor UO_2223 (O_2223,N_17765,N_15697);
or UO_2224 (O_2224,N_18816,N_19239);
nand UO_2225 (O_2225,N_15396,N_17763);
or UO_2226 (O_2226,N_16664,N_15102);
or UO_2227 (O_2227,N_19649,N_19441);
xor UO_2228 (O_2228,N_19334,N_19725);
and UO_2229 (O_2229,N_15045,N_16114);
xnor UO_2230 (O_2230,N_17207,N_17507);
nor UO_2231 (O_2231,N_16628,N_18868);
xnor UO_2232 (O_2232,N_16892,N_19032);
nor UO_2233 (O_2233,N_16582,N_17042);
or UO_2234 (O_2234,N_16549,N_18635);
or UO_2235 (O_2235,N_15020,N_15140);
or UO_2236 (O_2236,N_18801,N_18827);
and UO_2237 (O_2237,N_15694,N_16165);
xnor UO_2238 (O_2238,N_16830,N_17272);
nor UO_2239 (O_2239,N_18658,N_16242);
nor UO_2240 (O_2240,N_19558,N_15002);
nand UO_2241 (O_2241,N_15152,N_16333);
nor UO_2242 (O_2242,N_18176,N_17773);
and UO_2243 (O_2243,N_15301,N_15523);
or UO_2244 (O_2244,N_19788,N_17550);
and UO_2245 (O_2245,N_19304,N_19436);
nand UO_2246 (O_2246,N_17184,N_17761);
or UO_2247 (O_2247,N_16794,N_16825);
nor UO_2248 (O_2248,N_17233,N_19312);
and UO_2249 (O_2249,N_19251,N_19786);
nand UO_2250 (O_2250,N_19314,N_18146);
or UO_2251 (O_2251,N_16145,N_16728);
or UO_2252 (O_2252,N_18009,N_19206);
nor UO_2253 (O_2253,N_15704,N_15409);
xor UO_2254 (O_2254,N_17077,N_18078);
or UO_2255 (O_2255,N_16462,N_15165);
and UO_2256 (O_2256,N_17229,N_16630);
or UO_2257 (O_2257,N_18952,N_17433);
and UO_2258 (O_2258,N_18603,N_17367);
nor UO_2259 (O_2259,N_18916,N_18133);
or UO_2260 (O_2260,N_18321,N_19924);
nor UO_2261 (O_2261,N_16694,N_18626);
nor UO_2262 (O_2262,N_19812,N_15833);
and UO_2263 (O_2263,N_15662,N_16450);
and UO_2264 (O_2264,N_18465,N_16105);
xor UO_2265 (O_2265,N_16878,N_19872);
or UO_2266 (O_2266,N_18472,N_19747);
nor UO_2267 (O_2267,N_15371,N_19809);
or UO_2268 (O_2268,N_18948,N_16124);
nand UO_2269 (O_2269,N_16929,N_16691);
or UO_2270 (O_2270,N_17591,N_15084);
nor UO_2271 (O_2271,N_15595,N_19900);
nor UO_2272 (O_2272,N_19587,N_17619);
xnor UO_2273 (O_2273,N_18533,N_17566);
nand UO_2274 (O_2274,N_15077,N_18525);
nor UO_2275 (O_2275,N_18547,N_19577);
xnor UO_2276 (O_2276,N_17171,N_17709);
and UO_2277 (O_2277,N_18214,N_18551);
or UO_2278 (O_2278,N_19100,N_16205);
or UO_2279 (O_2279,N_17424,N_17626);
nand UO_2280 (O_2280,N_17850,N_16617);
xor UO_2281 (O_2281,N_18356,N_17364);
nor UO_2282 (O_2282,N_19816,N_19159);
or UO_2283 (O_2283,N_16997,N_18588);
or UO_2284 (O_2284,N_17462,N_19273);
nand UO_2285 (O_2285,N_19408,N_18973);
or UO_2286 (O_2286,N_18537,N_16298);
and UO_2287 (O_2287,N_16103,N_15203);
and UO_2288 (O_2288,N_19936,N_17647);
xnor UO_2289 (O_2289,N_15417,N_19217);
and UO_2290 (O_2290,N_17231,N_16156);
or UO_2291 (O_2291,N_19366,N_16132);
nor UO_2292 (O_2292,N_18590,N_19392);
nor UO_2293 (O_2293,N_18985,N_18545);
nor UO_2294 (O_2294,N_15669,N_15126);
and UO_2295 (O_2295,N_17599,N_18287);
nor UO_2296 (O_2296,N_17322,N_16274);
or UO_2297 (O_2297,N_17504,N_16420);
and UO_2298 (O_2298,N_16453,N_19805);
or UO_2299 (O_2299,N_17593,N_19121);
or UO_2300 (O_2300,N_17127,N_15433);
xor UO_2301 (O_2301,N_19419,N_18007);
and UO_2302 (O_2302,N_18649,N_15079);
or UO_2303 (O_2303,N_16471,N_18098);
and UO_2304 (O_2304,N_18856,N_16614);
and UO_2305 (O_2305,N_16065,N_15661);
nor UO_2306 (O_2306,N_19341,N_19035);
or UO_2307 (O_2307,N_15598,N_16390);
nor UO_2308 (O_2308,N_19667,N_17479);
xor UO_2309 (O_2309,N_16776,N_19591);
xnor UO_2310 (O_2310,N_15834,N_18655);
nand UO_2311 (O_2311,N_16423,N_18429);
nand UO_2312 (O_2312,N_15787,N_19704);
or UO_2313 (O_2313,N_16127,N_15086);
nor UO_2314 (O_2314,N_16221,N_17983);
and UO_2315 (O_2315,N_17460,N_19109);
or UO_2316 (O_2316,N_17176,N_18401);
or UO_2317 (O_2317,N_15164,N_19968);
nor UO_2318 (O_2318,N_16314,N_17114);
or UO_2319 (O_2319,N_17656,N_18902);
or UO_2320 (O_2320,N_16449,N_17759);
or UO_2321 (O_2321,N_18498,N_16577);
nand UO_2322 (O_2322,N_17401,N_16928);
and UO_2323 (O_2323,N_18817,N_17661);
and UO_2324 (O_2324,N_19781,N_18777);
nand UO_2325 (O_2325,N_15762,N_15435);
and UO_2326 (O_2326,N_16580,N_19546);
nor UO_2327 (O_2327,N_19151,N_16068);
nor UO_2328 (O_2328,N_15254,N_15994);
or UO_2329 (O_2329,N_18574,N_16177);
and UO_2330 (O_2330,N_18259,N_17645);
nor UO_2331 (O_2331,N_18782,N_19677);
nor UO_2332 (O_2332,N_18160,N_17161);
nor UO_2333 (O_2333,N_19191,N_15884);
or UO_2334 (O_2334,N_16066,N_15852);
nand UO_2335 (O_2335,N_15652,N_18852);
nor UO_2336 (O_2336,N_17386,N_16609);
nor UO_2337 (O_2337,N_17417,N_18809);
nand UO_2338 (O_2338,N_19480,N_16166);
and UO_2339 (O_2339,N_18444,N_15678);
and UO_2340 (O_2340,N_18994,N_17242);
or UO_2341 (O_2341,N_19965,N_16148);
xnor UO_2342 (O_2342,N_19215,N_17408);
xnor UO_2343 (O_2343,N_16610,N_15486);
nor UO_2344 (O_2344,N_19074,N_16877);
nand UO_2345 (O_2345,N_15259,N_17237);
nand UO_2346 (O_2346,N_18123,N_19775);
nor UO_2347 (O_2347,N_18040,N_17747);
and UO_2348 (O_2348,N_18967,N_17870);
xor UO_2349 (O_2349,N_17330,N_17054);
nor UO_2350 (O_2350,N_16227,N_15193);
or UO_2351 (O_2351,N_15172,N_16192);
and UO_2352 (O_2352,N_16604,N_16522);
nor UO_2353 (O_2353,N_19093,N_17571);
xnor UO_2354 (O_2354,N_16655,N_19659);
and UO_2355 (O_2355,N_18226,N_15302);
nand UO_2356 (O_2356,N_19862,N_15013);
and UO_2357 (O_2357,N_19042,N_18906);
and UO_2358 (O_2358,N_19989,N_18843);
and UO_2359 (O_2359,N_16719,N_15388);
or UO_2360 (O_2360,N_16368,N_18370);
nand UO_2361 (O_2361,N_17073,N_19661);
nor UO_2362 (O_2362,N_17153,N_15869);
xor UO_2363 (O_2363,N_15461,N_15923);
xnor UO_2364 (O_2364,N_19821,N_18850);
or UO_2365 (O_2365,N_17563,N_18193);
nor UO_2366 (O_2366,N_18307,N_18475);
xnor UO_2367 (O_2367,N_18956,N_15866);
and UO_2368 (O_2368,N_16133,N_16512);
nand UO_2369 (O_2369,N_18854,N_18795);
or UO_2370 (O_2370,N_19699,N_19607);
nand UO_2371 (O_2371,N_17439,N_16146);
or UO_2372 (O_2372,N_18564,N_16335);
or UO_2373 (O_2373,N_15295,N_17186);
xor UO_2374 (O_2374,N_18139,N_19056);
xnor UO_2375 (O_2375,N_17027,N_17177);
nand UO_2376 (O_2376,N_19995,N_15552);
nor UO_2377 (O_2377,N_15722,N_16731);
nand UO_2378 (O_2378,N_17230,N_17800);
or UO_2379 (O_2379,N_18270,N_16489);
or UO_2380 (O_2380,N_16318,N_17220);
nor UO_2381 (O_2381,N_15705,N_17360);
and UO_2382 (O_2382,N_17878,N_16076);
and UO_2383 (O_2383,N_19766,N_16801);
nand UO_2384 (O_2384,N_16859,N_19641);
nor UO_2385 (O_2385,N_15504,N_16028);
or UO_2386 (O_2386,N_19745,N_16806);
xor UO_2387 (O_2387,N_19633,N_18724);
nand UO_2388 (O_2388,N_18911,N_16947);
or UO_2389 (O_2389,N_17020,N_16149);
nand UO_2390 (O_2390,N_15969,N_15419);
and UO_2391 (O_2391,N_19863,N_16539);
nor UO_2392 (O_2392,N_19183,N_16781);
and UO_2393 (O_2393,N_16241,N_18246);
xor UO_2394 (O_2394,N_15190,N_17611);
nor UO_2395 (O_2395,N_19192,N_18970);
nor UO_2396 (O_2396,N_19077,N_17494);
and UO_2397 (O_2397,N_15305,N_17632);
nand UO_2398 (O_2398,N_18715,N_17945);
xnor UO_2399 (O_2399,N_15004,N_15460);
xnor UO_2400 (O_2400,N_17690,N_16439);
xor UO_2401 (O_2401,N_17714,N_17200);
and UO_2402 (O_2402,N_17788,N_17770);
nor UO_2403 (O_2403,N_15854,N_16482);
and UO_2404 (O_2404,N_17000,N_17080);
nor UO_2405 (O_2405,N_18756,N_18223);
nor UO_2406 (O_2406,N_18497,N_16472);
and UO_2407 (O_2407,N_15483,N_18822);
or UO_2408 (O_2408,N_18327,N_17892);
and UO_2409 (O_2409,N_18741,N_19417);
nor UO_2410 (O_2410,N_17163,N_19516);
or UO_2411 (O_2411,N_16493,N_19690);
xor UO_2412 (O_2412,N_16081,N_17515);
nor UO_2413 (O_2413,N_17855,N_17986);
and UO_2414 (O_2414,N_18051,N_17485);
xnor UO_2415 (O_2415,N_16865,N_17497);
nand UO_2416 (O_2416,N_17859,N_19413);
nor UO_2417 (O_2417,N_19763,N_18491);
or UO_2418 (O_2418,N_17780,N_17935);
nor UO_2419 (O_2419,N_16841,N_15907);
nand UO_2420 (O_2420,N_19572,N_17558);
and UO_2421 (O_2421,N_18569,N_18390);
xor UO_2422 (O_2422,N_19495,N_16230);
nor UO_2423 (O_2423,N_16969,N_18303);
and UO_2424 (O_2424,N_19363,N_18105);
xnor UO_2425 (O_2425,N_18748,N_18597);
or UO_2426 (O_2426,N_18932,N_16666);
nand UO_2427 (O_2427,N_19950,N_17961);
or UO_2428 (O_2428,N_18082,N_19397);
nand UO_2429 (O_2429,N_16616,N_16921);
and UO_2430 (O_2430,N_18740,N_16174);
nand UO_2431 (O_2431,N_18765,N_15353);
nand UO_2432 (O_2432,N_18053,N_19977);
or UO_2433 (O_2433,N_18269,N_19024);
nor UO_2434 (O_2434,N_16093,N_19177);
nand UO_2435 (O_2435,N_16999,N_17549);
xor UO_2436 (O_2436,N_15278,N_15745);
or UO_2437 (O_2437,N_18781,N_15343);
xnor UO_2438 (O_2438,N_19974,N_16319);
nand UO_2439 (O_2439,N_16665,N_18071);
xnor UO_2440 (O_2440,N_18766,N_16487);
and UO_2441 (O_2441,N_17538,N_16957);
nand UO_2442 (O_2442,N_19039,N_15075);
or UO_2443 (O_2443,N_18812,N_19176);
nor UO_2444 (O_2444,N_19175,N_15785);
and UO_2445 (O_2445,N_15160,N_15617);
nand UO_2446 (O_2446,N_18005,N_18690);
nor UO_2447 (O_2447,N_15358,N_17939);
xnor UO_2448 (O_2448,N_16748,N_19721);
xnor UO_2449 (O_2449,N_18539,N_15725);
and UO_2450 (O_2450,N_19404,N_19578);
xor UO_2451 (O_2451,N_18738,N_16518);
and UO_2452 (O_2452,N_19160,N_18820);
xnor UO_2453 (O_2453,N_15658,N_16110);
and UO_2454 (O_2454,N_17786,N_19895);
and UO_2455 (O_2455,N_19960,N_16326);
nand UO_2456 (O_2456,N_19567,N_17525);
nor UO_2457 (O_2457,N_17502,N_17475);
and UO_2458 (O_2458,N_18164,N_16583);
or UO_2459 (O_2459,N_19083,N_15036);
nand UO_2460 (O_2460,N_18221,N_19433);
or UO_2461 (O_2461,N_19207,N_17365);
and UO_2462 (O_2462,N_19848,N_15201);
or UO_2463 (O_2463,N_17290,N_18487);
nand UO_2464 (O_2464,N_15654,N_18233);
and UO_2465 (O_2465,N_19600,N_19698);
nor UO_2466 (O_2466,N_18404,N_18601);
or UO_2467 (O_2467,N_16330,N_15946);
or UO_2468 (O_2468,N_19072,N_18505);
xor UO_2469 (O_2469,N_19259,N_18286);
or UO_2470 (O_2470,N_19235,N_16926);
nor UO_2471 (O_2471,N_16195,N_16353);
xor UO_2472 (O_2472,N_17699,N_19282);
nor UO_2473 (O_2473,N_19091,N_18712);
and UO_2474 (O_2474,N_17019,N_15861);
nand UO_2475 (O_2475,N_19283,N_16463);
xnor UO_2476 (O_2476,N_16401,N_17482);
and UO_2477 (O_2477,N_18061,N_16526);
xnor UO_2478 (O_2478,N_17467,N_15981);
and UO_2479 (O_2479,N_17183,N_19882);
nand UO_2480 (O_2480,N_15401,N_18693);
nor UO_2481 (O_2481,N_16998,N_17931);
nand UO_2482 (O_2482,N_15263,N_17539);
nand UO_2483 (O_2483,N_19199,N_19332);
xnor UO_2484 (O_2484,N_19830,N_17383);
nor UO_2485 (O_2485,N_18374,N_15197);
nand UO_2486 (O_2486,N_16907,N_15294);
or UO_2487 (O_2487,N_17832,N_18174);
nor UO_2488 (O_2488,N_15551,N_17340);
nor UO_2489 (O_2489,N_19269,N_18520);
nor UO_2490 (O_2490,N_19946,N_15831);
or UO_2491 (O_2491,N_19185,N_15439);
xor UO_2492 (O_2492,N_17875,N_15445);
xor UO_2493 (O_2493,N_16203,N_19999);
xor UO_2494 (O_2494,N_18549,N_16350);
or UO_2495 (O_2495,N_17084,N_18688);
xor UO_2496 (O_2496,N_19412,N_17219);
xor UO_2497 (O_2497,N_15208,N_19827);
nor UO_2498 (O_2498,N_17398,N_17615);
nand UO_2499 (O_2499,N_18957,N_15577);
endmodule