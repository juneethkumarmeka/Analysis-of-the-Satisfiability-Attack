module basic_2500_25000_3000_5_levels_10xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
xor U0 (N_0,In_175,In_2339);
or U1 (N_1,In_1555,In_178);
and U2 (N_2,In_94,In_214);
xor U3 (N_3,In_2172,In_2365);
nor U4 (N_4,In_1965,In_2465);
and U5 (N_5,In_1041,In_1142);
or U6 (N_6,In_2231,In_1359);
and U7 (N_7,In_409,In_1714);
nand U8 (N_8,In_1260,In_2075);
xor U9 (N_9,In_2089,In_814);
nand U10 (N_10,In_341,In_1466);
and U11 (N_11,In_1299,In_40);
nand U12 (N_12,In_1331,In_1872);
xnor U13 (N_13,In_1831,In_1945);
or U14 (N_14,In_799,In_538);
xor U15 (N_15,In_2326,In_1074);
xor U16 (N_16,In_141,In_2021);
and U17 (N_17,In_46,In_1650);
nor U18 (N_18,In_1881,In_1743);
nand U19 (N_19,In_1439,In_2472);
and U20 (N_20,In_1649,In_1647);
nor U21 (N_21,In_897,In_669);
and U22 (N_22,In_2155,In_391);
xor U23 (N_23,In_2253,In_734);
or U24 (N_24,In_593,In_497);
nor U25 (N_25,In_2257,In_840);
nand U26 (N_26,In_563,In_1869);
nand U27 (N_27,In_235,In_1504);
or U28 (N_28,In_1636,In_394);
and U29 (N_29,In_348,In_584);
nand U30 (N_30,In_284,In_2066);
nor U31 (N_31,In_393,In_537);
xor U32 (N_32,In_1007,In_1775);
nor U33 (N_33,In_1762,In_1612);
nand U34 (N_34,In_1129,In_250);
nand U35 (N_35,In_2245,In_826);
xor U36 (N_36,In_1680,In_1319);
and U37 (N_37,In_323,In_1237);
or U38 (N_38,In_660,In_665);
or U39 (N_39,In_189,In_1428);
nand U40 (N_40,In_1002,In_659);
nand U41 (N_41,In_1355,In_1336);
xnor U42 (N_42,In_157,In_859);
nor U43 (N_43,In_1099,In_601);
xnor U44 (N_44,In_392,In_783);
and U45 (N_45,In_645,In_1370);
or U46 (N_46,In_219,In_1772);
nor U47 (N_47,In_2251,In_6);
or U48 (N_48,In_2111,In_1597);
xnor U49 (N_49,In_1075,In_1445);
xnor U50 (N_50,In_371,In_778);
nor U51 (N_51,In_1654,In_1613);
xor U52 (N_52,In_1685,In_1242);
xor U53 (N_53,In_2278,In_1713);
nand U54 (N_54,In_1012,In_692);
or U55 (N_55,In_1978,In_332);
nor U56 (N_56,In_953,In_1987);
and U57 (N_57,In_1692,In_180);
nor U58 (N_58,In_2003,In_354);
nand U59 (N_59,In_123,In_905);
or U60 (N_60,In_898,In_2043);
xor U61 (N_61,In_926,In_2330);
xor U62 (N_62,In_1936,In_66);
and U63 (N_63,In_700,In_1641);
nand U64 (N_64,In_122,In_23);
nand U65 (N_65,In_79,In_2364);
xor U66 (N_66,In_518,In_532);
nand U67 (N_67,In_662,In_1186);
xor U68 (N_68,In_213,In_2080);
and U69 (N_69,In_2417,In_2007);
xnor U70 (N_70,In_689,In_1414);
xor U71 (N_71,In_1939,In_291);
or U72 (N_72,In_2203,In_2039);
or U73 (N_73,In_390,In_2427);
or U74 (N_74,In_386,In_970);
nand U75 (N_75,In_282,In_1499);
nor U76 (N_76,In_2463,In_2232);
nor U77 (N_77,In_1658,In_2275);
or U78 (N_78,In_1410,In_1113);
nor U79 (N_79,In_204,In_1590);
nand U80 (N_80,In_998,In_1290);
xnor U81 (N_81,In_84,In_2009);
nand U82 (N_82,In_1033,In_1868);
or U83 (N_83,In_649,In_1028);
and U84 (N_84,In_1853,In_2138);
and U85 (N_85,In_242,In_2149);
nand U86 (N_86,In_479,In_2217);
and U87 (N_87,In_565,In_2185);
and U88 (N_88,In_1747,In_854);
xor U89 (N_89,In_1737,In_2421);
and U90 (N_90,In_476,In_1917);
or U91 (N_91,In_958,In_548);
xor U92 (N_92,In_2143,In_1357);
nand U93 (N_93,In_71,In_1746);
or U94 (N_94,In_1158,In_1572);
or U95 (N_95,In_1801,In_2261);
xor U96 (N_96,In_786,In_980);
xor U97 (N_97,In_224,In_1494);
and U98 (N_98,In_531,In_1855);
nand U99 (N_99,In_1971,In_2166);
and U100 (N_100,In_2206,In_1530);
nor U101 (N_101,In_1477,In_2052);
nand U102 (N_102,In_1206,In_668);
nand U103 (N_103,In_2340,In_2436);
or U104 (N_104,In_2101,In_2086);
and U105 (N_105,In_1856,In_2491);
and U106 (N_106,In_1284,In_251);
xor U107 (N_107,In_1994,In_930);
xor U108 (N_108,In_1546,In_2177);
nand U109 (N_109,In_2268,In_1644);
nand U110 (N_110,In_1066,In_1585);
or U111 (N_111,In_1086,In_1578);
nand U112 (N_112,In_1688,In_1553);
or U113 (N_113,In_1098,In_1887);
nand U114 (N_114,In_2032,In_1449);
nor U115 (N_115,In_1134,In_1305);
nor U116 (N_116,In_128,In_1720);
or U117 (N_117,In_300,In_368);
and U118 (N_118,In_1764,In_1678);
or U119 (N_119,In_871,In_1210);
and U120 (N_120,In_858,In_2377);
nor U121 (N_121,In_2316,In_1037);
xnor U122 (N_122,In_100,In_232);
nor U123 (N_123,In_505,In_1042);
nor U124 (N_124,In_776,In_794);
and U125 (N_125,In_1224,In_82);
and U126 (N_126,In_2460,In_1929);
xor U127 (N_127,In_329,In_1227);
nor U128 (N_128,In_2334,In_1958);
xnor U129 (N_129,In_975,In_252);
nor U130 (N_130,In_2422,In_95);
nor U131 (N_131,In_1493,In_1806);
nor U132 (N_132,In_2034,In_1683);
xnor U133 (N_133,In_1922,In_749);
nor U134 (N_134,In_891,In_363);
or U135 (N_135,In_1396,In_1263);
and U136 (N_136,In_194,In_1267);
and U137 (N_137,In_719,In_850);
xor U138 (N_138,In_1778,In_429);
nor U139 (N_139,In_2338,In_2384);
or U140 (N_140,In_1233,In_1600);
or U141 (N_141,In_328,In_2132);
xor U142 (N_142,In_2309,In_1670);
nor U143 (N_143,In_295,In_1858);
nand U144 (N_144,In_1123,In_1541);
nand U145 (N_145,In_864,In_248);
nor U146 (N_146,In_1666,In_2022);
and U147 (N_147,In_2091,In_2467);
nor U148 (N_148,In_583,In_913);
and U149 (N_149,In_31,In_2108);
xor U150 (N_150,In_158,In_1973);
and U151 (N_151,In_809,In_1053);
and U152 (N_152,In_2296,In_1866);
xnor U153 (N_153,In_1560,In_174);
xnor U154 (N_154,In_1380,In_925);
nand U155 (N_155,In_257,In_651);
and U156 (N_156,In_424,In_1852);
and U157 (N_157,In_1561,In_991);
nand U158 (N_158,In_1417,In_427);
and U159 (N_159,In_1722,In_202);
nand U160 (N_160,In_1470,In_2103);
xor U161 (N_161,In_2264,In_1223);
or U162 (N_162,In_1820,In_489);
and U163 (N_163,In_2133,In_109);
nand U164 (N_164,In_1972,In_2337);
or U165 (N_165,In_698,In_824);
and U166 (N_166,In_2462,In_1140);
nor U167 (N_167,In_347,In_2490);
nor U168 (N_168,In_261,In_615);
and U169 (N_169,In_1937,In_1532);
and U170 (N_170,In_2321,In_2492);
xnor U171 (N_171,In_2119,In_1838);
and U172 (N_172,In_724,In_1427);
nor U173 (N_173,In_682,In_2451);
and U174 (N_174,In_1418,In_1802);
nor U175 (N_175,In_1489,In_2450);
nor U176 (N_176,In_894,In_1593);
nand U177 (N_177,In_748,In_1615);
nor U178 (N_178,In_238,In_24);
or U179 (N_179,In_1162,In_1859);
or U180 (N_180,In_1784,In_1245);
xor U181 (N_181,In_661,In_993);
nor U182 (N_182,In_632,In_1501);
nand U183 (N_183,In_1883,In_83);
nand U184 (N_184,In_359,In_737);
or U185 (N_185,In_2051,In_1356);
or U186 (N_186,In_1787,In_863);
nor U187 (N_187,In_1222,In_1566);
or U188 (N_188,In_1824,In_713);
and U189 (N_189,In_350,In_2409);
nand U190 (N_190,In_977,In_1576);
nor U191 (N_191,In_417,In_2239);
nand U192 (N_192,In_1551,In_1239);
xnor U193 (N_193,In_1926,In_2248);
or U194 (N_194,In_412,In_800);
nor U195 (N_195,In_852,In_278);
or U196 (N_196,In_228,In_2184);
nand U197 (N_197,In_104,In_1264);
nand U198 (N_198,In_1165,In_12);
and U199 (N_199,In_1034,In_1554);
nand U200 (N_200,In_236,In_1520);
and U201 (N_201,In_145,In_1949);
nand U202 (N_202,In_2214,In_1312);
and U203 (N_203,In_1379,In_2348);
nor U204 (N_204,In_1163,In_1334);
nor U205 (N_205,In_1719,In_2197);
or U206 (N_206,In_265,In_2288);
or U207 (N_207,In_326,In_389);
nor U208 (N_208,In_316,In_1464);
and U209 (N_209,In_751,In_990);
nor U210 (N_210,In_2298,In_136);
xnor U211 (N_211,In_179,In_1731);
xnor U212 (N_212,In_1730,In_263);
or U213 (N_213,In_514,In_42);
nand U214 (N_214,In_1988,In_2096);
or U215 (N_215,In_1300,In_2192);
nand U216 (N_216,In_432,In_156);
nand U217 (N_217,In_1810,In_1019);
or U218 (N_218,In_1207,In_1347);
xnor U219 (N_219,In_483,In_801);
nor U220 (N_220,In_1628,In_1216);
or U221 (N_221,In_1540,In_846);
nor U222 (N_222,In_1502,In_2160);
nand U223 (N_223,In_2107,In_663);
or U224 (N_224,In_1055,In_1202);
and U225 (N_225,In_1897,In_591);
and U226 (N_226,In_922,In_1339);
or U227 (N_227,In_1458,In_1382);
xor U228 (N_228,In_149,In_673);
nor U229 (N_229,In_2434,In_1841);
nor U230 (N_230,In_470,In_444);
or U231 (N_231,In_415,In_2292);
xor U232 (N_232,In_804,In_2148);
and U233 (N_233,In_2265,In_2050);
nor U234 (N_234,In_2225,In_1921);
or U235 (N_235,In_1294,In_1911);
nand U236 (N_236,In_866,In_1960);
or U237 (N_237,In_511,In_2286);
or U238 (N_238,In_954,In_186);
nor U239 (N_239,In_1441,In_2006);
xor U240 (N_240,In_1259,In_1729);
nand U241 (N_241,In_899,In_1409);
nor U242 (N_242,In_1558,In_2152);
and U243 (N_243,In_1387,In_2224);
and U244 (N_244,In_699,In_227);
nand U245 (N_245,In_1057,In_2415);
nor U246 (N_246,In_1862,In_694);
xnor U247 (N_247,In_1545,In_2025);
xor U248 (N_248,In_159,In_225);
and U249 (N_249,In_2129,In_75);
and U250 (N_250,In_312,In_572);
or U251 (N_251,In_2341,In_2024);
nand U252 (N_252,In_1811,In_1669);
xor U253 (N_253,In_1990,In_657);
nor U254 (N_254,In_64,In_2084);
and U255 (N_255,In_1742,In_672);
xor U256 (N_256,In_1372,In_683);
xor U257 (N_257,In_705,In_2379);
xnor U258 (N_258,In_2213,In_318);
xnor U259 (N_259,In_1150,In_1715);
and U260 (N_260,In_861,In_1350);
nand U261 (N_261,In_1953,In_2473);
xnor U262 (N_262,In_299,In_2060);
or U263 (N_263,In_1465,In_540);
or U264 (N_264,In_1082,In_857);
xnor U265 (N_265,In_289,In_2351);
xnor U266 (N_266,In_1705,In_2123);
xnor U267 (N_267,In_249,In_357);
xor U268 (N_268,In_568,In_1984);
nand U269 (N_269,In_1995,In_2163);
xor U270 (N_270,In_1352,In_845);
xnor U271 (N_271,In_1480,In_2355);
nand U272 (N_272,In_50,In_810);
and U273 (N_273,In_1825,In_1663);
or U274 (N_274,In_1420,In_1419);
and U275 (N_275,In_2033,In_1138);
and U276 (N_276,In_60,In_573);
and U277 (N_277,In_2469,In_791);
or U278 (N_278,In_86,In_2190);
and U279 (N_279,In_1254,In_892);
nand U280 (N_280,In_723,In_637);
nand U281 (N_281,In_653,In_1518);
and U282 (N_282,In_2497,In_1905);
nand U283 (N_283,In_1635,In_2130);
and U284 (N_284,In_982,In_2036);
or U285 (N_285,In_1864,In_87);
nand U286 (N_286,In_634,In_113);
and U287 (N_287,In_1890,In_2414);
nand U288 (N_288,In_851,In_221);
nand U289 (N_289,In_2346,In_1845);
xor U290 (N_290,In_1891,In_1633);
nor U291 (N_291,In_667,In_121);
nand U292 (N_292,In_1107,In_274);
nand U293 (N_293,In_731,In_464);
and U294 (N_294,In_1416,In_1812);
nand U295 (N_295,In_703,In_22);
nor U296 (N_296,In_853,In_743);
nand U297 (N_297,In_1095,In_870);
nand U298 (N_298,In_495,In_1269);
nor U299 (N_299,In_675,In_1790);
nor U300 (N_300,In_2136,In_1592);
xnor U301 (N_301,In_1084,In_865);
and U302 (N_302,In_552,In_450);
nand U303 (N_303,In_1009,In_1094);
or U304 (N_304,In_1457,In_2029);
xnor U305 (N_305,In_2229,In_1923);
nor U306 (N_306,In_1059,In_191);
nand U307 (N_307,In_607,In_217);
nor U308 (N_308,In_2402,In_2280);
nand U309 (N_309,In_349,In_519);
xor U310 (N_310,In_1423,In_2423);
or U311 (N_311,In_162,In_2097);
nor U312 (N_312,In_1006,In_2470);
nand U313 (N_313,In_1570,In_2484);
nor U314 (N_314,In_1961,In_2183);
nor U315 (N_315,In_2110,In_346);
and U316 (N_316,In_331,In_276);
nor U317 (N_317,In_2223,In_395);
xor U318 (N_318,In_912,In_333);
or U319 (N_319,In_493,In_1884);
nand U320 (N_320,In_1744,In_2358);
xor U321 (N_321,In_596,In_1101);
nor U322 (N_322,In_2131,In_51);
nand U323 (N_323,In_1383,In_55);
xnor U324 (N_324,In_603,In_1789);
nor U325 (N_325,In_1488,In_119);
or U326 (N_326,In_1511,In_681);
nor U327 (N_327,In_1909,In_1882);
and U328 (N_328,In_307,In_1193);
nand U329 (N_329,In_2076,In_1924);
nor U330 (N_330,In_2437,In_197);
nand U331 (N_331,In_463,In_1433);
nand U332 (N_332,In_2312,In_860);
and U333 (N_333,In_481,In_674);
nor U334 (N_334,In_847,In_1854);
nor U335 (N_335,In_1345,In_2287);
or U336 (N_336,In_901,In_1467);
or U337 (N_337,In_1885,In_397);
xor U338 (N_338,In_304,In_1384);
nor U339 (N_339,In_1249,In_1371);
nand U340 (N_340,In_2063,In_2283);
or U341 (N_341,In_2461,In_2078);
nor U342 (N_342,In_617,In_1351);
or U343 (N_343,In_137,In_2241);
or U344 (N_344,In_226,In_15);
xor U345 (N_345,In_484,In_1303);
nor U346 (N_346,In_380,In_1252);
nand U347 (N_347,In_1673,In_2387);
and U348 (N_348,In_2015,In_1124);
nor U349 (N_349,In_269,In_2452);
or U350 (N_350,In_153,In_2204);
or U351 (N_351,In_618,In_20);
or U352 (N_352,In_2082,In_775);
and U353 (N_353,In_1954,In_1940);
nor U354 (N_354,In_1127,In_2226);
and U355 (N_355,In_1759,In_1393);
and U356 (N_356,In_869,In_1308);
and U357 (N_357,In_728,In_1927);
nand U358 (N_358,In_2019,In_1521);
nand U359 (N_359,In_1310,In_2016);
or U360 (N_360,In_570,In_2094);
xor U361 (N_361,In_1736,In_478);
nor U362 (N_362,In_1378,In_1172);
nor U363 (N_363,In_1894,In_73);
nor U364 (N_364,In_1577,In_1694);
nor U365 (N_365,In_406,In_1657);
nand U366 (N_366,In_1281,In_2295);
or U367 (N_367,In_446,In_1221);
and U368 (N_368,In_1725,In_1873);
nor U369 (N_369,In_556,In_1998);
xor U370 (N_370,In_1429,In_862);
and U371 (N_371,In_1947,In_272);
and U372 (N_372,In_696,In_2055);
nor U373 (N_373,In_1071,In_240);
nand U374 (N_374,In_971,In_1340);
xnor U375 (N_375,In_1146,In_1563);
xor U376 (N_376,In_770,In_2318);
and U377 (N_377,In_258,In_2040);
nand U378 (N_378,In_34,In_99);
and U379 (N_379,In_1933,In_678);
or U380 (N_380,In_2013,In_2366);
xnor U381 (N_381,In_53,In_77);
xnor U382 (N_382,In_989,In_2099);
nand U383 (N_383,In_2297,In_528);
and U384 (N_384,In_1443,In_27);
xor U385 (N_385,In_1161,In_2109);
or U386 (N_386,In_1748,In_2401);
xor U387 (N_387,In_2201,In_1803);
or U388 (N_388,In_2256,In_788);
xor U389 (N_389,In_1826,In_697);
nor U390 (N_390,In_513,In_222);
nor U391 (N_391,In_233,In_932);
xor U392 (N_392,In_2398,In_1605);
nand U393 (N_393,In_1286,In_1079);
nor U394 (N_394,In_500,In_1951);
and U395 (N_395,In_1377,In_1814);
and U396 (N_396,In_1614,In_1788);
and U397 (N_397,In_1693,In_1178);
nor U398 (N_398,In_2262,In_1438);
nand U399 (N_399,In_590,In_542);
nor U400 (N_400,In_1471,In_592);
or U401 (N_401,In_340,In_1609);
xor U402 (N_402,In_437,In_1255);
or U403 (N_403,In_773,In_283);
or U404 (N_404,In_1106,In_2125);
nor U405 (N_405,In_1681,In_1332);
xor U406 (N_406,In_576,In_2393);
nor U407 (N_407,In_1726,In_554);
xor U408 (N_408,In_1874,In_942);
xnor U409 (N_409,In_2236,In_1840);
nand U410 (N_410,In_1950,In_1968);
xnor U411 (N_411,In_402,In_420);
or U412 (N_412,In_887,In_2390);
or U413 (N_413,In_729,In_2215);
or U414 (N_414,In_2211,In_1587);
xor U415 (N_415,In_268,In_578);
nand U416 (N_416,In_294,In_1050);
nor U417 (N_417,In_1112,In_598);
nand U418 (N_418,In_886,In_296);
xnor U419 (N_419,In_2005,In_1205);
and U420 (N_420,In_353,In_834);
or U421 (N_421,In_647,In_2322);
and U422 (N_422,In_582,In_2222);
nor U423 (N_423,In_1583,In_223);
and U424 (N_424,In_1358,In_676);
or U425 (N_425,In_762,In_802);
or U426 (N_426,In_1794,In_2046);
nor U427 (N_427,In_1584,In_1979);
and U428 (N_428,In_1608,In_1529);
nand U429 (N_429,In_408,In_680);
or U430 (N_430,In_1157,In_1324);
nand U431 (N_431,In_650,In_1996);
nor U432 (N_432,In_1816,In_2323);
or U433 (N_433,In_1181,In_1413);
xnor U434 (N_434,In_445,In_37);
and U435 (N_435,In_44,In_237);
xnor U436 (N_436,In_1238,In_1989);
nand U437 (N_437,In_1738,In_716);
or U438 (N_438,In_461,In_2361);
nor U439 (N_439,In_1089,In_1456);
or U440 (N_440,In_1510,In_2475);
or U441 (N_441,In_2030,In_654);
nand U442 (N_442,In_1625,In_1620);
and U443 (N_443,In_2416,In_2430);
nor U444 (N_444,In_301,In_2244);
nand U445 (N_445,In_1860,In_1580);
nor U446 (N_446,In_943,In_494);
or U447 (N_447,In_1035,In_1970);
or U448 (N_448,In_1513,In_198);
or U449 (N_449,In_411,In_1315);
nor U450 (N_450,In_2140,In_1646);
nand U451 (N_451,In_11,In_47);
nand U452 (N_452,In_1011,In_963);
and U453 (N_453,In_396,In_74);
nor U454 (N_454,In_2081,In_695);
nor U455 (N_455,In_1388,In_2333);
and U456 (N_456,In_1629,In_1373);
nor U457 (N_457,In_453,In_2207);
xor U458 (N_458,In_1671,In_1436);
or U459 (N_459,In_1039,In_1808);
nand U460 (N_460,In_14,In_1791);
nand U461 (N_461,In_1783,In_112);
and U462 (N_462,In_2221,In_606);
or U463 (N_463,In_485,In_1696);
and U464 (N_464,In_1473,In_374);
xnor U465 (N_465,In_419,In_1000);
xor U466 (N_466,In_2282,In_1076);
nand U467 (N_467,In_1195,In_1807);
nand U468 (N_468,In_1607,In_2435);
or U469 (N_469,In_725,In_1991);
nand U470 (N_470,In_1268,In_588);
xor U471 (N_471,In_325,In_959);
or U472 (N_472,In_594,In_1068);
nor U473 (N_473,In_45,In_836);
and U474 (N_474,In_1048,In_973);
or U475 (N_475,In_1631,In_1301);
nand U476 (N_476,In_155,In_566);
xor U477 (N_477,In_164,In_712);
nor U478 (N_478,In_992,In_1490);
or U479 (N_479,In_766,In_828);
and U480 (N_480,In_2153,In_343);
or U481 (N_481,In_848,In_2271);
nand U482 (N_482,In_130,In_986);
and U483 (N_483,In_1918,In_1621);
xnor U484 (N_484,In_984,In_2182);
nor U485 (N_485,In_1200,In_1478);
and U486 (N_486,In_1411,In_1166);
or U487 (N_487,In_1786,In_1323);
and U488 (N_488,In_1500,In_1226);
nand U489 (N_489,In_1728,In_2202);
nor U490 (N_490,In_101,In_297);
and U491 (N_491,In_1344,In_2315);
nand U492 (N_492,In_2456,In_1754);
xor U493 (N_493,In_614,In_2342);
and U494 (N_494,In_527,In_2112);
xnor U495 (N_495,In_143,In_739);
or U496 (N_496,In_338,In_2233);
nand U497 (N_497,In_193,In_2382);
xnor U498 (N_498,In_2480,In_2065);
and U499 (N_499,In_1486,In_1652);
or U500 (N_500,In_62,In_260);
nand U501 (N_501,In_2299,In_1088);
nor U502 (N_502,In_835,In_273);
xnor U503 (N_503,In_2105,In_1491);
nand U504 (N_504,In_2289,In_337);
or U505 (N_505,In_2234,In_2372);
and U506 (N_506,In_1931,In_1538);
or U507 (N_507,In_1509,In_1562);
and U508 (N_508,In_808,In_2062);
and U509 (N_509,In_413,In_935);
xnor U510 (N_510,In_1220,In_2068);
and U511 (N_511,In_76,In_327);
or U512 (N_512,In_2162,In_2117);
xnor U513 (N_513,In_133,In_706);
nand U514 (N_514,In_29,In_581);
or U515 (N_515,In_2499,In_523);
and U516 (N_516,In_1718,In_927);
or U517 (N_517,In_1367,In_1219);
xnor U518 (N_518,In_1120,In_670);
nand U519 (N_519,In_2432,In_2073);
xnor U520 (N_520,In_1262,In_638);
xnor U521 (N_521,In_308,In_267);
and U522 (N_522,In_543,In_1974);
xnor U523 (N_523,In_1516,In_2157);
nand U524 (N_524,In_1253,In_1777);
nand U525 (N_525,In_1780,In_1225);
xor U526 (N_526,In_1201,In_401);
and U527 (N_527,In_2407,In_1935);
nand U528 (N_528,In_2165,In_1288);
xor U529 (N_529,In_1667,In_1505);
and U530 (N_530,In_1295,In_375);
xnor U531 (N_531,In_2147,In_792);
xnor U532 (N_532,In_2468,In_2164);
xor U533 (N_533,In_1865,In_2260);
and U534 (N_534,In_1391,In_812);
nor U535 (N_535,In_1879,In_968);
and U536 (N_536,In_431,In_1248);
and U537 (N_537,In_1085,In_1064);
or U538 (N_538,In_2494,In_1363);
nor U539 (N_539,In_2293,In_207);
and U540 (N_540,In_1495,In_2189);
nand U541 (N_541,In_2385,In_2057);
nand U542 (N_542,In_934,In_1559);
nor U543 (N_543,In_1153,In_933);
nand U544 (N_544,In_1627,In_1228);
or U545 (N_545,In_2240,In_1311);
and U546 (N_546,In_2424,In_1376);
nor U547 (N_547,In_192,In_946);
or U548 (N_548,In_896,In_1077);
and U549 (N_549,In_883,In_1131);
or U550 (N_550,In_589,In_2325);
xnor U551 (N_551,In_972,In_701);
and U552 (N_552,In_1708,In_486);
or U553 (N_553,In_1136,In_522);
nand U554 (N_554,In_919,In_8);
and U555 (N_555,In_741,In_1648);
xnor U556 (N_556,In_1765,In_1460);
nor U557 (N_557,In_69,In_1533);
or U558 (N_558,In_182,In_1156);
nor U559 (N_559,In_2156,In_1687);
nand U560 (N_560,In_1761,In_208);
nand U561 (N_561,In_2174,In_1374);
or U562 (N_562,In_414,In_502);
nand U563 (N_563,In_163,In_2227);
and U564 (N_564,In_1348,In_1755);
and U565 (N_565,In_714,In_2270);
and U566 (N_566,In_416,In_1063);
nor U567 (N_567,In_1451,In_790);
and U568 (N_568,In_1707,In_2028);
or U569 (N_569,In_1622,In_831);
nor U570 (N_570,In_2400,In_533);
nand U571 (N_571,In_1274,In_462);
and U572 (N_572,In_421,In_2018);
and U573 (N_573,In_1481,In_2403);
or U574 (N_574,In_2263,In_2235);
and U575 (N_575,In_1103,In_314);
and U576 (N_576,In_1325,In_165);
xnor U577 (N_577,In_880,In_586);
and U578 (N_578,In_1168,In_203);
nor U579 (N_579,In_1361,In_1750);
xor U580 (N_580,In_1208,In_1758);
or U581 (N_581,In_287,In_436);
nor U582 (N_582,In_2284,In_1589);
or U583 (N_583,In_1606,In_2049);
nor U584 (N_584,In_1946,In_2059);
nor U585 (N_585,In_423,In_1769);
nor U586 (N_586,In_1187,In_2048);
nand U587 (N_587,In_1174,In_1976);
nor U588 (N_588,In_2104,In_1137);
and U589 (N_589,In_367,In_184);
nor U590 (N_590,In_1781,In_2085);
or U591 (N_591,In_1752,In_907);
or U592 (N_592,In_1699,In_994);
nand U593 (N_593,In_784,In_1243);
or U594 (N_594,In_1828,In_1712);
nor U595 (N_595,In_2158,In_1536);
xor U596 (N_596,In_715,In_21);
nor U597 (N_597,In_2308,In_2114);
nand U598 (N_598,In_2126,In_30);
nor U599 (N_599,In_422,In_736);
xnor U600 (N_600,In_2406,In_856);
and U601 (N_601,In_452,In_1934);
or U602 (N_602,In_2479,In_1360);
nand U603 (N_603,In_1525,In_906);
and U604 (N_604,In_448,In_2483);
or U605 (N_605,In_2383,In_2276);
and U606 (N_606,In_147,In_1637);
nand U607 (N_607,In_1964,In_2319);
nand U608 (N_608,In_1013,In_2336);
nor U609 (N_609,In_1512,In_759);
or U610 (N_610,In_1674,In_1655);
nor U611 (N_611,In_735,In_1318);
nor U612 (N_612,In_1899,In_1848);
or U613 (N_613,In_1321,In_434);
xor U614 (N_614,In_1517,In_878);
or U615 (N_615,In_2307,In_2173);
nand U616 (N_616,In_376,In_1676);
or U617 (N_617,In_1240,In_1804);
and U618 (N_618,In_825,In_438);
xnor U619 (N_619,In_2272,In_286);
and U620 (N_620,In_1293,In_1903);
nor U621 (N_621,In_777,In_983);
nor U622 (N_622,In_2311,In_2420);
nand U623 (N_623,In_822,In_1723);
xor U624 (N_624,In_1975,In_17);
and U625 (N_625,In_1322,In_1930);
nand U626 (N_626,In_2357,In_1073);
or U627 (N_627,In_32,In_319);
nor U628 (N_628,In_1767,In_1645);
and U629 (N_629,In_711,In_1703);
nor U630 (N_630,In_629,In_2150);
xor U631 (N_631,In_628,In_957);
and U632 (N_632,In_255,In_433);
nor U633 (N_633,In_303,In_2464);
or U634 (N_634,In_1506,In_1544);
and U635 (N_635,In_160,In_2195);
and U636 (N_636,In_2412,In_2250);
nand U637 (N_637,In_89,In_873);
and U638 (N_638,In_2041,In_524);
nand U639 (N_639,In_1537,In_2302);
and U640 (N_640,In_458,In_1170);
nor U641 (N_641,In_456,In_1959);
xor U642 (N_642,In_335,In_909);
nand U643 (N_643,In_1381,In_798);
xor U644 (N_644,In_931,In_2077);
nor U645 (N_645,In_345,In_510);
or U646 (N_646,In_2061,In_1406);
xnor U647 (N_647,In_1045,In_1183);
and U648 (N_648,In_1199,In_2376);
nor U649 (N_649,In_466,In_1425);
or U650 (N_650,In_1401,In_379);
and U651 (N_651,In_787,In_1582);
and U652 (N_652,In_460,In_1919);
nand U653 (N_653,In_562,In_1198);
nor U654 (N_654,In_1479,In_1328);
xor U655 (N_655,In_652,In_1022);
and U656 (N_656,In_63,In_111);
xnor U657 (N_657,In_138,In_655);
xnor U658 (N_658,In_2363,In_19);
nor U659 (N_659,In_764,In_1815);
and U660 (N_660,In_1813,In_1152);
nor U661 (N_661,In_1482,In_1404);
or U662 (N_662,In_1304,In_1796);
or U663 (N_663,In_1141,In_620);
nand U664 (N_664,In_923,In_311);
or U665 (N_665,In_1462,In_1003);
xor U666 (N_666,In_781,In_1330);
nor U667 (N_667,In_1682,In_1450);
or U668 (N_668,In_1739,In_1756);
and U669 (N_669,In_1285,In_893);
and U670 (N_670,In_1817,In_1782);
xnor U671 (N_671,In_2127,In_220);
or U672 (N_672,In_1836,In_1702);
nand U673 (N_673,In_85,In_2139);
or U674 (N_674,In_1125,In_135);
nand U675 (N_675,In_2145,In_530);
xor U676 (N_676,In_844,In_2178);
or U677 (N_677,In_2443,In_2482);
or U678 (N_678,In_1966,In_888);
and U679 (N_679,In_1044,In_471);
or U680 (N_680,In_1070,In_440);
xor U681 (N_681,In_1118,In_2359);
nor U682 (N_682,In_1058,In_1706);
or U683 (N_683,In_1008,In_910);
nand U684 (N_684,In_200,In_969);
nand U685 (N_685,In_362,In_558);
nand U686 (N_686,In_546,In_721);
or U687 (N_687,In_2026,In_1832);
nand U688 (N_688,In_1915,In_785);
nand U689 (N_689,In_360,In_1397);
nor U690 (N_690,In_2255,In_1122);
nor U691 (N_691,In_1876,In_1271);
or U692 (N_692,In_955,In_1032);
or U693 (N_693,In_351,In_1167);
nor U694 (N_694,In_921,In_266);
and U695 (N_695,In_1052,In_1639);
nand U696 (N_696,In_1487,In_152);
and U697 (N_697,In_939,In_1709);
nor U698 (N_698,In_988,In_57);
and U699 (N_699,In_817,In_68);
or U700 (N_700,In_1054,In_1661);
nor U701 (N_701,In_2273,In_1539);
or U702 (N_702,In_823,In_2433);
nor U703 (N_703,In_1036,In_517);
and U704 (N_704,In_974,In_754);
xnor U705 (N_705,In_229,In_1797);
nand U706 (N_706,In_1920,In_383);
nor U707 (N_707,In_795,In_96);
and U708 (N_708,In_25,In_1507);
nand U709 (N_709,In_507,In_467);
nor U710 (N_710,In_2106,In_172);
or U711 (N_711,In_1999,In_356);
nand U712 (N_712,In_755,In_1851);
nor U713 (N_713,In_146,In_1251);
nand U714 (N_714,In_1638,In_1145);
nand U715 (N_715,In_843,In_1306);
xor U716 (N_716,In_410,In_1944);
and U717 (N_717,In_1565,In_1912);
or U718 (N_718,In_2368,In_1618);
or U719 (N_719,In_539,In_1132);
and U720 (N_720,In_2476,In_1721);
nor U721 (N_721,In_911,In_428);
xor U722 (N_722,In_1474,In_43);
and U723 (N_723,In_39,In_1176);
and U724 (N_724,In_2493,In_1);
nor U725 (N_725,In_443,In_2489);
nand U726 (N_726,In_1065,In_313);
or U727 (N_727,In_90,In_2014);
or U728 (N_728,In_2053,In_439);
xnor U729 (N_729,In_206,In_1829);
and U730 (N_730,In_1030,In_187);
nor U731 (N_731,In_545,In_398);
nor U732 (N_732,In_28,In_551);
xnor U733 (N_733,In_960,In_1871);
xnor U734 (N_734,In_2444,In_2237);
nor U735 (N_735,In_1010,In_1117);
xnor U736 (N_736,In_664,In_2254);
xnor U737 (N_737,In_1595,In_1431);
and U738 (N_738,In_474,In_310);
or U739 (N_739,In_1932,In_2481);
and U740 (N_740,In_451,In_298);
nor U741 (N_741,In_855,In_2056);
xnor U742 (N_742,In_2012,In_1368);
or U743 (N_743,In_499,In_1476);
or U744 (N_744,In_1837,In_2392);
nand U745 (N_745,In_1795,In_1497);
or U746 (N_746,In_1320,In_169);
or U747 (N_747,In_35,In_595);
and U748 (N_748,In_1619,In_1596);
xnor U749 (N_749,In_976,In_2004);
nand U750 (N_750,In_1038,In_2266);
xor U751 (N_751,In_1437,In_1446);
nor U752 (N_752,In_1880,In_10);
nor U753 (N_753,In_2335,In_2405);
or U754 (N_754,In_1611,In_1185);
and U755 (N_755,In_702,In_521);
nand U756 (N_756,In_1403,In_129);
or U757 (N_757,In_612,In_937);
or U758 (N_758,In_1492,In_2252);
xnor U759 (N_759,In_239,In_2378);
xor U760 (N_760,In_2281,In_837);
or U761 (N_761,In_677,In_2176);
or U762 (N_762,In_5,In_2304);
nand U763 (N_763,In_1567,In_496);
nand U764 (N_764,In_1955,In_1434);
nand U765 (N_765,In_315,In_1190);
nand U766 (N_766,In_1689,In_2001);
xor U767 (N_767,In_106,In_2124);
or U768 (N_768,In_1234,In_830);
nor U769 (N_769,In_161,In_950);
xnor U770 (N_770,In_1277,In_916);
xor U771 (N_771,In_48,In_279);
or U772 (N_772,In_358,In_1067);
nand U773 (N_773,In_631,In_2445);
and U774 (N_774,In_1400,In_1213);
xor U775 (N_775,In_730,In_1901);
or U776 (N_776,In_2303,In_704);
xor U777 (N_777,In_2179,In_1716);
nor U778 (N_778,In_752,In_1483);
xor U779 (N_779,In_2210,In_1279);
and U780 (N_780,In_181,In_780);
xnor U781 (N_781,In_388,In_2045);
nand U782 (N_782,In_281,In_407);
nand U783 (N_783,In_2453,In_2181);
and U784 (N_784,In_920,In_482);
nand U785 (N_785,In_903,In_718);
or U786 (N_786,In_1115,In_2426);
xor U787 (N_787,In_2277,In_1272);
xnor U788 (N_788,In_512,In_515);
nor U789 (N_789,In_579,In_1229);
nand U790 (N_790,In_967,In_1405);
nand U791 (N_791,In_120,In_807);
nand U792 (N_792,In_1847,In_1329);
nand U793 (N_793,In_154,In_1734);
xor U794 (N_794,In_945,In_1514);
nand U795 (N_795,In_234,In_2243);
xor U796 (N_796,In_833,In_806);
xor U797 (N_797,In_1992,In_1651);
nand U798 (N_798,In_150,In_2353);
nand U799 (N_799,In_1604,In_321);
nand U800 (N_800,In_2171,In_1977);
nor U801 (N_801,In_1818,In_874);
or U802 (N_802,In_342,In_372);
nand U803 (N_803,In_365,In_2449);
xnor U804 (N_804,In_2356,In_382);
or U805 (N_805,In_1610,In_1745);
and U806 (N_806,In_2259,In_1155);
nand U807 (N_807,In_442,In_738);
nor U808 (N_808,In_38,In_1395);
or U809 (N_809,In_1078,In_1522);
nand U810 (N_810,In_1362,In_1527);
and U811 (N_811,In_2498,In_369);
and U812 (N_812,In_52,In_1475);
or U813 (N_813,In_2209,In_740);
and U814 (N_814,In_1016,In_480);
or U815 (N_815,In_1046,In_2345);
xnor U816 (N_816,In_1913,In_2399);
and U817 (N_817,In_642,In_2120);
xor U818 (N_818,In_81,In_1843);
and U819 (N_819,In_477,In_2344);
nor U820 (N_820,In_330,In_2332);
xnor U821 (N_821,In_838,In_475);
xor U822 (N_822,In_640,In_1800);
xnor U823 (N_823,In_2100,In_671);
and U824 (N_824,In_387,In_1834);
nand U825 (N_825,In_167,In_1724);
nand U826 (N_826,In_132,In_2440);
xor U827 (N_827,In_1004,In_1697);
xnor U828 (N_828,In_1983,In_1957);
nor U829 (N_829,In_1878,In_684);
and U830 (N_830,In_97,In_2069);
nand U831 (N_831,In_339,In_2064);
nand U832 (N_832,In_549,In_107);
nor U833 (N_833,In_1849,In_185);
xor U834 (N_834,In_564,In_2098);
nor U835 (N_835,In_2305,In_1907);
xor U836 (N_836,In_127,In_33);
nor U837 (N_837,In_2074,In_449);
nor U838 (N_838,In_2418,In_41);
xnor U839 (N_839,In_2429,In_915);
xnor U840 (N_840,In_2457,In_2455);
or U841 (N_841,In_218,In_1598);
xor U842 (N_842,In_1399,In_1571);
nor U843 (N_843,In_2389,In_1139);
nand U844 (N_844,In_2218,In_1341);
nand U845 (N_845,In_1569,In_473);
or U846 (N_846,In_1291,In_1447);
nand U847 (N_847,In_1215,In_80);
nand U848 (N_848,In_666,In_1160);
or U849 (N_849,In_140,In_1247);
nor U850 (N_850,In_173,In_979);
xor U851 (N_851,In_2198,In_2313);
or U852 (N_852,In_245,In_78);
and U853 (N_853,In_1133,In_625);
or U854 (N_854,In_1298,In_426);
or U855 (N_855,In_2391,In_1444);
xnor U856 (N_856,In_2238,In_627);
or U857 (N_857,In_285,In_1792);
nand U858 (N_858,In_1735,In_488);
xnor U859 (N_859,In_796,In_938);
nand U860 (N_860,In_2485,In_613);
or U861 (N_861,In_2347,In_1938);
or U862 (N_862,In_733,In_717);
and U863 (N_863,In_211,In_2290);
or U864 (N_864,In_88,In_636);
nor U865 (N_865,In_557,In_633);
xor U866 (N_866,In_457,In_1154);
xnor U867 (N_867,In_535,In_575);
xor U868 (N_868,In_1867,In_956);
nand U869 (N_869,In_2141,In_2300);
or U870 (N_870,In_117,In_805);
nand U871 (N_871,In_447,In_1793);
xnor U872 (N_872,In_768,In_1993);
and U873 (N_873,In_1111,In_1798);
xnor U874 (N_874,In_1586,In_720);
xnor U875 (N_875,In_277,In_567);
xnor U876 (N_876,In_1943,In_1753);
xnor U877 (N_877,In_621,In_908);
xor U878 (N_878,In_1180,In_487);
nand U879 (N_879,In_1617,In_2031);
or U880 (N_880,In_1727,In_2187);
nand U881 (N_881,In_658,In_441);
or U882 (N_882,In_1177,In_1896);
xnor U883 (N_883,In_418,In_2072);
nand U884 (N_884,In_364,In_550);
or U885 (N_885,In_2396,In_1029);
or U886 (N_886,In_1025,In_803);
nor U887 (N_887,In_914,In_879);
nand U888 (N_888,In_2327,In_2137);
and U889 (N_889,In_1556,In_771);
nor U890 (N_890,In_1656,In_1257);
nand U891 (N_891,In_2386,In_622);
nor U892 (N_892,In_1543,In_2011);
nand U893 (N_893,In_1732,In_262);
or U894 (N_894,In_1952,In_2488);
and U895 (N_895,In_679,In_1452);
nor U896 (N_896,In_1942,In_18);
xor U897 (N_897,In_1194,In_1421);
xor U898 (N_898,In_199,In_1928);
nor U899 (N_899,In_1270,In_608);
nand U900 (N_900,In_2458,In_2228);
nor U901 (N_901,In_1981,In_2135);
and U902 (N_902,In_691,In_985);
and U903 (N_903,In_1515,In_2010);
nor U904 (N_904,In_384,In_1179);
or U905 (N_905,In_2431,In_2329);
or U906 (N_906,In_490,In_1785);
nand U907 (N_907,In_1455,In_1542);
nor U908 (N_908,In_2194,In_832);
nor U909 (N_909,In_793,In_758);
or U910 (N_910,In_246,In_195);
nor U911 (N_911,In_1534,In_1547);
or U912 (N_912,In_1159,In_67);
xor U913 (N_913,In_305,In_2274);
and U914 (N_914,In_2380,In_1895);
nor U915 (N_915,In_2425,In_2291);
or U916 (N_916,In_2167,In_2186);
nand U917 (N_917,In_1484,In_1307);
xor U918 (N_918,In_2373,In_114);
nor U919 (N_919,In_2478,In_105);
or U920 (N_920,In_400,In_1774);
nand U921 (N_921,In_306,In_2267);
or U922 (N_922,In_1969,In_49);
and U923 (N_923,In_115,In_816);
xnor U924 (N_924,In_827,In_302);
nand U925 (N_925,In_623,In_1292);
nand U926 (N_926,In_1760,In_2144);
or U927 (N_927,In_1925,In_1302);
nor U928 (N_928,In_2246,In_2193);
nand U929 (N_929,In_102,In_2044);
nand U930 (N_930,In_2219,In_2087);
and U931 (N_931,In_1276,In_1863);
nand U932 (N_932,In_1664,In_209);
nor U933 (N_933,In_580,In_2037);
and U934 (N_934,In_829,In_526);
nor U935 (N_935,In_1018,In_1844);
nand U936 (N_936,In_1910,In_2369);
or U937 (N_937,In_952,In_2367);
or U938 (N_938,In_587,In_1642);
nor U939 (N_939,In_710,In_1005);
nand U940 (N_940,In_1900,In_760);
nor U941 (N_941,In_1105,In_91);
nor U942 (N_942,In_2331,In_1001);
and U943 (N_943,In_1850,In_1232);
nand U944 (N_944,In_243,In_889);
and U945 (N_945,In_611,In_1568);
nand U946 (N_946,In_216,In_2038);
xnor U947 (N_947,In_961,In_1822);
xnor U948 (N_948,In_688,In_1698);
xor U949 (N_949,In_544,In_1857);
and U950 (N_950,In_686,In_1346);
nor U951 (N_951,In_1870,In_1888);
nand U952 (N_952,In_585,In_1408);
or U953 (N_953,In_813,In_1072);
or U954 (N_954,In_468,In_244);
nor U955 (N_955,In_1135,In_1564);
or U956 (N_956,In_2095,In_1779);
or U957 (N_957,In_1763,In_2180);
and U958 (N_958,In_644,In_2362);
or U959 (N_959,In_270,In_2374);
xor U960 (N_960,In_188,In_108);
and U961 (N_961,In_72,In_2306);
nor U962 (N_962,In_600,In_604);
xnor U963 (N_963,In_1591,In_1246);
nor U964 (N_964,In_1496,In_2205);
or U965 (N_965,In_2446,In_819);
and U966 (N_966,In_275,In_708);
and U967 (N_967,In_2230,In_2151);
nor U968 (N_968,In_797,In_1442);
and U969 (N_969,In_1861,In_964);
or U970 (N_970,In_520,In_1632);
xnor U971 (N_971,In_2191,In_336);
nor U972 (N_972,In_1024,In_491);
nand U973 (N_973,In_1963,In_2413);
xor U974 (N_974,In_1327,In_2419);
nand U975 (N_975,In_2301,In_54);
xor U976 (N_976,In_1773,In_2454);
and U977 (N_977,In_1169,In_1503);
nor U978 (N_978,In_936,In_2188);
or U979 (N_979,In_1126,In_2121);
and U980 (N_980,In_2212,In_509);
or U981 (N_981,In_882,In_2200);
nor U982 (N_982,In_171,In_405);
nor U983 (N_983,In_196,In_254);
and U984 (N_984,In_2067,In_536);
or U985 (N_985,In_1061,In_148);
xnor U986 (N_986,In_1402,In_1108);
or U987 (N_987,In_1144,In_648);
xor U988 (N_988,In_1212,In_1967);
and U989 (N_989,In_2071,In_190);
nor U990 (N_990,In_2447,In_1508);
nand U991 (N_991,In_1192,In_504);
nand U992 (N_992,In_1261,In_2128);
or U993 (N_993,In_2175,In_290);
nor U994 (N_994,In_746,In_1892);
nor U995 (N_995,In_1015,In_2352);
nand U996 (N_996,In_1768,In_1603);
and U997 (N_997,In_2058,In_98);
or U998 (N_998,In_1275,In_508);
and U999 (N_999,In_1426,In_1757);
and U1000 (N_1000,In_247,In_2441);
nand U1001 (N_1001,In_1230,In_2208);
or U1002 (N_1002,In_2442,In_2242);
xnor U1003 (N_1003,In_58,In_872);
nand U1004 (N_1004,In_1588,In_610);
xor U1005 (N_1005,In_693,In_1717);
xnor U1006 (N_1006,In_1695,In_1342);
and U1007 (N_1007,In_643,In_1119);
and U1008 (N_1008,In_1904,In_1415);
or U1009 (N_1009,In_1104,In_1700);
nand U1010 (N_1010,In_656,In_868);
xnor U1011 (N_1011,In_1081,In_1463);
or U1012 (N_1012,In_516,In_1557);
nand U1013 (N_1013,In_1313,In_1102);
or U1014 (N_1014,In_7,In_1948);
or U1015 (N_1015,In_1660,In_574);
nor U1016 (N_1016,In_2381,In_1594);
or U1017 (N_1017,In_1616,In_2);
xor U1018 (N_1018,In_1833,In_1021);
xor U1019 (N_1019,In_947,In_2349);
or U1020 (N_1020,In_2083,In_134);
nand U1021 (N_1021,In_1733,In_1549);
nand U1022 (N_1022,In_26,In_320);
nor U1023 (N_1023,In_1805,In_1175);
nand U1024 (N_1024,In_1665,In_1100);
nor U1025 (N_1025,In_1147,In_212);
nand U1026 (N_1026,In_1244,In_1908);
and U1027 (N_1027,In_1017,In_110);
nor U1028 (N_1028,In_1114,In_1148);
and U1029 (N_1029,In_2027,In_1333);
or U1030 (N_1030,In_1266,In_1751);
nor U1031 (N_1031,In_378,In_1711);
nand U1032 (N_1032,In_547,In_732);
and U1033 (N_1033,In_1353,In_1093);
or U1034 (N_1034,In_2146,In_2168);
and U1035 (N_1035,In_1386,In_1398);
or U1036 (N_1036,In_1060,In_1314);
nor U1037 (N_1037,In_1191,In_769);
or U1038 (N_1038,In_1839,In_2486);
nor U1039 (N_1039,In_2496,In_1083);
nand U1040 (N_1040,In_1485,In_2047);
nand U1041 (N_1041,In_1893,In_1809);
nand U1042 (N_1042,In_177,In_722);
nor U1043 (N_1043,In_1047,In_503);
xnor U1044 (N_1044,In_2017,In_1027);
nand U1045 (N_1045,In_292,In_2404);
and U1046 (N_1046,In_498,In_818);
or U1047 (N_1047,In_753,In_1823);
nor U1048 (N_1048,In_1273,In_2448);
nor U1049 (N_1049,In_1898,In_765);
nor U1050 (N_1050,In_116,In_687);
nor U1051 (N_1051,In_929,In_1283);
and U1052 (N_1052,In_1776,In_1548);
nand U1053 (N_1053,In_2216,In_1623);
nand U1054 (N_1054,In_560,In_1846);
nand U1055 (N_1055,In_1258,In_1519);
xnor U1056 (N_1056,In_501,In_1550);
or U1057 (N_1057,In_2495,In_205);
nor U1058 (N_1058,In_1096,In_309);
nand U1059 (N_1059,In_1602,In_1278);
nand U1060 (N_1060,In_1256,In_529);
xor U1061 (N_1061,In_2279,In_890);
nand U1062 (N_1062,In_1526,In_215);
nand U1063 (N_1063,In_1296,In_1316);
or U1064 (N_1064,In_2079,In_506);
xor U1065 (N_1065,In_690,In_944);
xnor U1066 (N_1066,In_355,In_767);
nand U1067 (N_1067,In_940,In_2070);
xnor U1068 (N_1068,In_324,In_1343);
and U1069 (N_1069,In_1469,In_1235);
nand U1070 (N_1070,In_1842,In_1188);
xor U1071 (N_1071,In_981,In_377);
or U1072 (N_1072,In_877,In_124);
xnor U1073 (N_1073,In_231,In_264);
or U1074 (N_1074,In_1090,In_472);
xnor U1075 (N_1075,In_1349,In_1231);
xor U1076 (N_1076,In_1454,In_92);
nand U1077 (N_1077,In_1309,In_201);
nand U1078 (N_1078,In_1461,In_492);
and U1079 (N_1079,In_334,In_756);
nand U1080 (N_1080,In_2090,In_900);
and U1081 (N_1081,In_0,In_2020);
or U1082 (N_1082,In_1440,In_1217);
nand U1083 (N_1083,In_1448,In_1407);
nor U1084 (N_1084,In_1830,In_1128);
nor U1085 (N_1085,In_1412,In_1980);
or U1086 (N_1086,In_2142,In_2360);
nor U1087 (N_1087,In_1143,In_1690);
and U1088 (N_1088,In_1280,In_1424);
and U1089 (N_1089,In_1121,In_13);
and U1090 (N_1090,In_1189,In_65);
nor U1091 (N_1091,In_2487,In_1203);
and U1092 (N_1092,In_820,In_1528);
nor U1093 (N_1093,In_36,In_2159);
nor U1094 (N_1094,In_1749,In_1710);
and U1095 (N_1095,In_2042,In_2343);
nor U1096 (N_1096,In_1640,In_1827);
and U1097 (N_1097,In_2118,In_941);
nand U1098 (N_1098,In_2054,In_256);
nand U1099 (N_1099,In_435,In_2471);
nand U1100 (N_1100,In_1164,In_2269);
nand U1101 (N_1101,In_1265,In_1741);
nor U1102 (N_1102,In_381,In_1365);
or U1103 (N_1103,In_996,In_1366);
and U1104 (N_1104,In_3,In_93);
and U1105 (N_1105,In_895,In_1109);
or U1106 (N_1106,In_1043,In_1821);
xor U1107 (N_1107,In_561,In_2035);
xnor U1108 (N_1108,In_1552,In_1581);
or U1109 (N_1109,In_1422,In_9);
nor U1110 (N_1110,In_1287,In_2161);
nand U1111 (N_1111,In_747,In_962);
nor U1112 (N_1112,In_1182,In_2102);
nand U1113 (N_1113,In_1902,In_842);
or U1114 (N_1114,In_2394,In_789);
xnor U1115 (N_1115,In_2196,In_1056);
xor U1116 (N_1116,In_1364,In_1337);
or U1117 (N_1117,In_2371,In_949);
or U1118 (N_1118,In_841,In_1875);
or U1119 (N_1119,In_2438,In_1338);
xor U1120 (N_1120,In_1601,In_126);
nor U1121 (N_1121,In_183,In_1432);
nand U1122 (N_1122,In_1886,In_1662);
xnor U1123 (N_1123,In_1531,In_641);
nor U1124 (N_1124,In_259,In_125);
nand U1125 (N_1125,In_1130,In_280);
and U1126 (N_1126,In_2466,In_1092);
xor U1127 (N_1127,In_1297,In_1317);
or U1128 (N_1128,In_1385,In_2285);
xnor U1129 (N_1129,In_995,In_139);
nand U1130 (N_1130,In_1236,In_1659);
nor U1131 (N_1131,In_399,In_230);
xor U1132 (N_1132,In_1799,In_1173);
and U1133 (N_1133,In_1023,In_541);
and U1134 (N_1134,In_2314,In_709);
and U1135 (N_1135,In_1634,In_727);
nor U1136 (N_1136,In_2169,In_2354);
nand U1137 (N_1137,In_1250,In_1062);
nand U1138 (N_1138,In_1459,In_2324);
nor U1139 (N_1139,In_2122,In_902);
nand U1140 (N_1140,In_1677,In_1031);
and U1141 (N_1141,In_1472,In_525);
or U1142 (N_1142,In_271,In_553);
or U1143 (N_1143,In_1579,In_559);
xnor U1144 (N_1144,In_2395,In_965);
or U1145 (N_1145,In_815,In_875);
nor U1146 (N_1146,In_2477,In_2000);
nand U1147 (N_1147,In_1986,In_430);
xnor U1148 (N_1148,In_571,In_2474);
xnor U1149 (N_1149,In_1211,In_811);
and U1150 (N_1150,In_881,In_2170);
xnor U1151 (N_1151,In_2093,In_924);
and U1152 (N_1152,In_1906,In_1498);
xnor U1153 (N_1153,In_997,In_948);
xor U1154 (N_1154,In_602,In_2397);
nor U1155 (N_1155,In_344,In_1209);
or U1156 (N_1156,In_1672,In_569);
nand U1157 (N_1157,In_2320,In_779);
and U1158 (N_1158,In_999,In_454);
nand U1159 (N_1159,In_1691,In_1204);
or U1160 (N_1160,In_1770,In_366);
xor U1161 (N_1161,In_763,In_1997);
or U1162 (N_1162,In_2317,In_1675);
xnor U1163 (N_1163,In_1624,In_1282);
nand U1164 (N_1164,In_1375,In_626);
and U1165 (N_1165,In_1653,In_1049);
or U1166 (N_1166,In_1051,In_176);
nor U1167 (N_1167,In_2370,In_742);
or U1168 (N_1168,In_1116,In_577);
or U1169 (N_1169,In_821,In_774);
and U1170 (N_1170,In_884,In_951);
and U1171 (N_1171,In_761,In_555);
xor U1172 (N_1172,In_1435,In_1394);
nor U1173 (N_1173,In_459,In_2258);
nor U1174 (N_1174,In_385,In_639);
nor U1175 (N_1175,In_1626,In_2002);
xnor U1176 (N_1176,In_151,In_170);
or U1177 (N_1177,In_1184,In_118);
or U1178 (N_1178,In_2088,In_4);
and U1179 (N_1179,In_2116,In_1686);
or U1180 (N_1180,In_361,In_726);
and U1181 (N_1181,In_61,In_772);
xor U1182 (N_1182,In_1241,In_635);
or U1183 (N_1183,In_253,In_1985);
nand U1184 (N_1184,In_1668,In_2310);
or U1185 (N_1185,In_646,In_839);
nand U1186 (N_1186,In_928,In_1171);
nand U1187 (N_1187,In_1819,In_917);
nor U1188 (N_1188,In_744,In_597);
xnor U1189 (N_1189,In_144,In_1956);
or U1190 (N_1190,In_2408,In_745);
or U1191 (N_1191,In_56,In_2199);
or U1192 (N_1192,In_978,In_1040);
and U1193 (N_1193,In_876,In_1684);
nor U1194 (N_1194,In_2113,In_1289);
nor U1195 (N_1195,In_1069,In_624);
and U1196 (N_1196,In_1941,In_619);
or U1197 (N_1197,In_2092,In_1766);
nor U1198 (N_1198,In_849,In_1889);
nor U1199 (N_1199,In_1468,In_685);
and U1200 (N_1200,In_1430,In_1630);
and U1201 (N_1201,In_469,In_352);
and U1202 (N_1202,In_1740,In_1962);
and U1203 (N_1203,In_288,In_1643);
xor U1204 (N_1204,In_1877,In_142);
and U1205 (N_1205,In_1087,In_293);
or U1206 (N_1206,In_59,In_2459);
nor U1207 (N_1207,In_1679,In_1392);
and U1208 (N_1208,In_465,In_987);
nor U1209 (N_1209,In_1214,In_317);
nand U1210 (N_1210,In_2375,In_373);
and U1211 (N_1211,In_1390,In_707);
or U1212 (N_1212,In_2008,In_2439);
or U1213 (N_1213,In_131,In_1196);
and U1214 (N_1214,In_1091,In_605);
xnor U1215 (N_1215,In_1701,In_370);
nand U1216 (N_1216,In_616,In_609);
xnor U1217 (N_1217,In_1110,In_2388);
xor U1218 (N_1218,In_1535,In_2428);
or U1219 (N_1219,In_966,In_1026);
nor U1220 (N_1220,In_210,In_1335);
or U1221 (N_1221,In_1835,In_168);
or U1222 (N_1222,In_757,In_1524);
nor U1223 (N_1223,In_1771,In_918);
or U1224 (N_1224,In_2247,In_1453);
or U1225 (N_1225,In_2134,In_455);
nand U1226 (N_1226,In_2328,In_1575);
nand U1227 (N_1227,In_1574,In_534);
or U1228 (N_1228,In_1218,In_1916);
or U1229 (N_1229,In_599,In_1599);
nand U1230 (N_1230,In_1197,In_403);
nand U1231 (N_1231,In_1097,In_16);
nor U1232 (N_1232,In_904,In_2154);
nor U1233 (N_1233,In_1523,In_2115);
nor U1234 (N_1234,In_1704,In_885);
nand U1235 (N_1235,In_2220,In_1014);
nor U1236 (N_1236,In_1982,In_404);
nor U1237 (N_1237,In_630,In_2023);
and U1238 (N_1238,In_1389,In_1080);
nand U1239 (N_1239,In_70,In_322);
nand U1240 (N_1240,In_1369,In_782);
and U1241 (N_1241,In_867,In_1354);
nor U1242 (N_1242,In_103,In_2410);
nand U1243 (N_1243,In_1151,In_1149);
xnor U1244 (N_1244,In_1326,In_2411);
nor U1245 (N_1245,In_1020,In_1914);
xnor U1246 (N_1246,In_2350,In_1573);
nand U1247 (N_1247,In_166,In_750);
nor U1248 (N_1248,In_241,In_2294);
xor U1249 (N_1249,In_425,In_2249);
nand U1250 (N_1250,In_927,In_89);
or U1251 (N_1251,In_464,In_935);
nand U1252 (N_1252,In_2062,In_749);
or U1253 (N_1253,In_1923,In_877);
nand U1254 (N_1254,In_1988,In_1140);
and U1255 (N_1255,In_257,In_479);
and U1256 (N_1256,In_1215,In_1468);
nor U1257 (N_1257,In_1735,In_480);
and U1258 (N_1258,In_1450,In_56);
nor U1259 (N_1259,In_367,In_2130);
nor U1260 (N_1260,In_405,In_211);
xor U1261 (N_1261,In_1496,In_17);
nor U1262 (N_1262,In_1921,In_898);
xnor U1263 (N_1263,In_1384,In_1133);
nand U1264 (N_1264,In_2226,In_1832);
xnor U1265 (N_1265,In_1947,In_1304);
nor U1266 (N_1266,In_2461,In_813);
xnor U1267 (N_1267,In_1719,In_496);
nor U1268 (N_1268,In_438,In_1746);
nor U1269 (N_1269,In_2225,In_1943);
or U1270 (N_1270,In_2230,In_3);
nor U1271 (N_1271,In_1544,In_549);
xor U1272 (N_1272,In_260,In_424);
nor U1273 (N_1273,In_2462,In_871);
or U1274 (N_1274,In_1030,In_1454);
and U1275 (N_1275,In_2474,In_1709);
nor U1276 (N_1276,In_1504,In_1711);
and U1277 (N_1277,In_1674,In_930);
nand U1278 (N_1278,In_336,In_76);
and U1279 (N_1279,In_1860,In_1822);
nand U1280 (N_1280,In_1248,In_820);
xnor U1281 (N_1281,In_582,In_1472);
nor U1282 (N_1282,In_1309,In_1520);
nor U1283 (N_1283,In_437,In_198);
or U1284 (N_1284,In_2002,In_2228);
nand U1285 (N_1285,In_2411,In_1593);
nand U1286 (N_1286,In_1040,In_1404);
nor U1287 (N_1287,In_1447,In_2376);
nor U1288 (N_1288,In_1184,In_628);
or U1289 (N_1289,In_428,In_404);
nor U1290 (N_1290,In_2399,In_1053);
xnor U1291 (N_1291,In_1658,In_635);
nor U1292 (N_1292,In_1343,In_1146);
and U1293 (N_1293,In_2102,In_2379);
nor U1294 (N_1294,In_1051,In_2146);
or U1295 (N_1295,In_646,In_771);
nand U1296 (N_1296,In_1169,In_2240);
xnor U1297 (N_1297,In_673,In_2306);
nand U1298 (N_1298,In_974,In_535);
nor U1299 (N_1299,In_1366,In_2482);
and U1300 (N_1300,In_332,In_2290);
or U1301 (N_1301,In_2062,In_2484);
nor U1302 (N_1302,In_1187,In_2370);
and U1303 (N_1303,In_371,In_78);
or U1304 (N_1304,In_1774,In_1702);
nand U1305 (N_1305,In_200,In_213);
nand U1306 (N_1306,In_2056,In_2153);
xor U1307 (N_1307,In_767,In_2275);
or U1308 (N_1308,In_1752,In_1811);
xor U1309 (N_1309,In_1150,In_2109);
nor U1310 (N_1310,In_2109,In_308);
nand U1311 (N_1311,In_2269,In_1082);
nor U1312 (N_1312,In_1344,In_1218);
or U1313 (N_1313,In_1111,In_1781);
xor U1314 (N_1314,In_646,In_1695);
nor U1315 (N_1315,In_541,In_325);
or U1316 (N_1316,In_613,In_238);
nand U1317 (N_1317,In_2155,In_1944);
or U1318 (N_1318,In_561,In_83);
nor U1319 (N_1319,In_695,In_411);
nand U1320 (N_1320,In_1053,In_1895);
xor U1321 (N_1321,In_2246,In_68);
xnor U1322 (N_1322,In_1628,In_1305);
nor U1323 (N_1323,In_1656,In_1753);
or U1324 (N_1324,In_154,In_2130);
and U1325 (N_1325,In_821,In_1765);
nor U1326 (N_1326,In_1524,In_1122);
xor U1327 (N_1327,In_2387,In_1031);
or U1328 (N_1328,In_301,In_387);
nor U1329 (N_1329,In_2092,In_970);
or U1330 (N_1330,In_1651,In_1697);
and U1331 (N_1331,In_1434,In_499);
nand U1332 (N_1332,In_330,In_1227);
xnor U1333 (N_1333,In_1428,In_1543);
nand U1334 (N_1334,In_983,In_78);
xnor U1335 (N_1335,In_584,In_1456);
nand U1336 (N_1336,In_1861,In_524);
nor U1337 (N_1337,In_1427,In_2455);
nand U1338 (N_1338,In_459,In_1036);
and U1339 (N_1339,In_817,In_2462);
nand U1340 (N_1340,In_627,In_650);
and U1341 (N_1341,In_2192,In_2417);
xnor U1342 (N_1342,In_146,In_79);
or U1343 (N_1343,In_666,In_2050);
nand U1344 (N_1344,In_175,In_2266);
nand U1345 (N_1345,In_1593,In_851);
nand U1346 (N_1346,In_2018,In_1826);
nor U1347 (N_1347,In_1145,In_69);
nor U1348 (N_1348,In_1747,In_419);
and U1349 (N_1349,In_467,In_697);
or U1350 (N_1350,In_1811,In_1694);
and U1351 (N_1351,In_1326,In_2032);
xnor U1352 (N_1352,In_2179,In_485);
nand U1353 (N_1353,In_151,In_561);
and U1354 (N_1354,In_824,In_2301);
and U1355 (N_1355,In_250,In_465);
nor U1356 (N_1356,In_1995,In_984);
and U1357 (N_1357,In_648,In_1220);
xnor U1358 (N_1358,In_47,In_2274);
or U1359 (N_1359,In_1226,In_1291);
or U1360 (N_1360,In_2446,In_1760);
and U1361 (N_1361,In_2100,In_1894);
nor U1362 (N_1362,In_1475,In_2454);
or U1363 (N_1363,In_1455,In_2007);
nor U1364 (N_1364,In_873,In_622);
xnor U1365 (N_1365,In_306,In_2251);
xor U1366 (N_1366,In_644,In_1695);
xnor U1367 (N_1367,In_1682,In_1763);
and U1368 (N_1368,In_1205,In_1452);
and U1369 (N_1369,In_1185,In_838);
or U1370 (N_1370,In_1553,In_217);
nand U1371 (N_1371,In_1922,In_1307);
nand U1372 (N_1372,In_2027,In_1127);
xnor U1373 (N_1373,In_2496,In_2342);
nand U1374 (N_1374,In_786,In_1086);
nand U1375 (N_1375,In_1737,In_2130);
or U1376 (N_1376,In_2093,In_2074);
xor U1377 (N_1377,In_1862,In_661);
nor U1378 (N_1378,In_1141,In_1417);
or U1379 (N_1379,In_1780,In_1865);
and U1380 (N_1380,In_777,In_786);
xor U1381 (N_1381,In_1676,In_57);
or U1382 (N_1382,In_990,In_2398);
nand U1383 (N_1383,In_1753,In_2320);
and U1384 (N_1384,In_479,In_2214);
or U1385 (N_1385,In_520,In_1295);
nor U1386 (N_1386,In_512,In_1534);
and U1387 (N_1387,In_665,In_0);
nand U1388 (N_1388,In_1871,In_77);
or U1389 (N_1389,In_2310,In_2392);
and U1390 (N_1390,In_1388,In_2086);
nor U1391 (N_1391,In_1333,In_539);
or U1392 (N_1392,In_1120,In_2174);
and U1393 (N_1393,In_2368,In_527);
and U1394 (N_1394,In_1145,In_1057);
or U1395 (N_1395,In_1606,In_1403);
nand U1396 (N_1396,In_1366,In_942);
nor U1397 (N_1397,In_278,In_1666);
xnor U1398 (N_1398,In_16,In_2080);
nor U1399 (N_1399,In_1717,In_431);
or U1400 (N_1400,In_1885,In_600);
xor U1401 (N_1401,In_1015,In_1271);
xor U1402 (N_1402,In_1161,In_1767);
and U1403 (N_1403,In_895,In_2313);
nor U1404 (N_1404,In_660,In_1100);
nand U1405 (N_1405,In_778,In_1229);
or U1406 (N_1406,In_467,In_28);
or U1407 (N_1407,In_645,In_2032);
or U1408 (N_1408,In_674,In_151);
xnor U1409 (N_1409,In_1616,In_2149);
and U1410 (N_1410,In_90,In_575);
or U1411 (N_1411,In_1300,In_1244);
or U1412 (N_1412,In_1227,In_2349);
xnor U1413 (N_1413,In_909,In_1747);
and U1414 (N_1414,In_1336,In_608);
and U1415 (N_1415,In_1715,In_2302);
xor U1416 (N_1416,In_1562,In_579);
nand U1417 (N_1417,In_1014,In_400);
nor U1418 (N_1418,In_922,In_977);
nand U1419 (N_1419,In_703,In_1154);
or U1420 (N_1420,In_1473,In_2312);
xnor U1421 (N_1421,In_1590,In_1267);
nor U1422 (N_1422,In_402,In_1097);
and U1423 (N_1423,In_2144,In_1857);
nor U1424 (N_1424,In_1724,In_1945);
xor U1425 (N_1425,In_560,In_1924);
nor U1426 (N_1426,In_236,In_284);
xnor U1427 (N_1427,In_1991,In_2498);
nor U1428 (N_1428,In_2290,In_1686);
nor U1429 (N_1429,In_1518,In_422);
or U1430 (N_1430,In_205,In_2313);
nor U1431 (N_1431,In_2391,In_2358);
nor U1432 (N_1432,In_2357,In_821);
nor U1433 (N_1433,In_1504,In_1849);
nand U1434 (N_1434,In_1809,In_1320);
and U1435 (N_1435,In_182,In_1246);
xor U1436 (N_1436,In_1092,In_2272);
xnor U1437 (N_1437,In_2304,In_108);
nor U1438 (N_1438,In_1103,In_1343);
xor U1439 (N_1439,In_10,In_1936);
nor U1440 (N_1440,In_451,In_332);
nor U1441 (N_1441,In_402,In_255);
and U1442 (N_1442,In_747,In_2073);
or U1443 (N_1443,In_1568,In_1810);
and U1444 (N_1444,In_2231,In_384);
nor U1445 (N_1445,In_242,In_1297);
and U1446 (N_1446,In_91,In_608);
and U1447 (N_1447,In_2248,In_1548);
or U1448 (N_1448,In_1139,In_603);
nand U1449 (N_1449,In_2439,In_55);
nand U1450 (N_1450,In_1504,In_545);
and U1451 (N_1451,In_610,In_1256);
nand U1452 (N_1452,In_1199,In_2042);
nor U1453 (N_1453,In_1950,In_2389);
xor U1454 (N_1454,In_2078,In_576);
and U1455 (N_1455,In_1372,In_1300);
nor U1456 (N_1456,In_2443,In_1137);
and U1457 (N_1457,In_57,In_204);
nor U1458 (N_1458,In_2254,In_1230);
nor U1459 (N_1459,In_681,In_260);
or U1460 (N_1460,In_2018,In_1884);
or U1461 (N_1461,In_1081,In_1144);
xnor U1462 (N_1462,In_750,In_2413);
nand U1463 (N_1463,In_1505,In_2377);
xnor U1464 (N_1464,In_484,In_1544);
and U1465 (N_1465,In_344,In_1215);
xor U1466 (N_1466,In_405,In_2455);
and U1467 (N_1467,In_222,In_2435);
nand U1468 (N_1468,In_1401,In_782);
or U1469 (N_1469,In_312,In_489);
nand U1470 (N_1470,In_1792,In_1186);
nor U1471 (N_1471,In_171,In_1301);
nor U1472 (N_1472,In_1773,In_131);
nor U1473 (N_1473,In_2030,In_529);
nor U1474 (N_1474,In_1847,In_1646);
nor U1475 (N_1475,In_1106,In_232);
or U1476 (N_1476,In_398,In_355);
nor U1477 (N_1477,In_410,In_51);
and U1478 (N_1478,In_1718,In_882);
nor U1479 (N_1479,In_1271,In_666);
or U1480 (N_1480,In_1725,In_1203);
nor U1481 (N_1481,In_1721,In_185);
nor U1482 (N_1482,In_1748,In_474);
nand U1483 (N_1483,In_1650,In_1996);
xor U1484 (N_1484,In_2186,In_1295);
nand U1485 (N_1485,In_555,In_36);
nand U1486 (N_1486,In_1309,In_2456);
and U1487 (N_1487,In_143,In_1774);
nor U1488 (N_1488,In_355,In_505);
and U1489 (N_1489,In_1028,In_2345);
nor U1490 (N_1490,In_1190,In_1153);
and U1491 (N_1491,In_1416,In_1823);
xnor U1492 (N_1492,In_1194,In_1994);
nand U1493 (N_1493,In_488,In_602);
nand U1494 (N_1494,In_2383,In_240);
and U1495 (N_1495,In_396,In_1314);
and U1496 (N_1496,In_262,In_1842);
xnor U1497 (N_1497,In_485,In_1161);
or U1498 (N_1498,In_427,In_89);
nand U1499 (N_1499,In_524,In_2016);
or U1500 (N_1500,In_2061,In_1989);
nor U1501 (N_1501,In_1624,In_1113);
xnor U1502 (N_1502,In_1359,In_1540);
xor U1503 (N_1503,In_2104,In_490);
xor U1504 (N_1504,In_2058,In_1336);
xnor U1505 (N_1505,In_1954,In_678);
nor U1506 (N_1506,In_1184,In_1933);
xor U1507 (N_1507,In_2424,In_446);
nand U1508 (N_1508,In_1227,In_125);
xnor U1509 (N_1509,In_1615,In_1239);
nand U1510 (N_1510,In_1064,In_282);
nor U1511 (N_1511,In_1528,In_2334);
nand U1512 (N_1512,In_2028,In_1409);
and U1513 (N_1513,In_2438,In_1838);
nand U1514 (N_1514,In_2049,In_1216);
xor U1515 (N_1515,In_1506,In_576);
and U1516 (N_1516,In_1851,In_1976);
nand U1517 (N_1517,In_846,In_1040);
nand U1518 (N_1518,In_103,In_933);
nand U1519 (N_1519,In_1449,In_1240);
nor U1520 (N_1520,In_2127,In_705);
and U1521 (N_1521,In_989,In_987);
and U1522 (N_1522,In_1473,In_1588);
nor U1523 (N_1523,In_1778,In_545);
or U1524 (N_1524,In_762,In_2468);
nand U1525 (N_1525,In_1490,In_818);
or U1526 (N_1526,In_429,In_151);
and U1527 (N_1527,In_1049,In_1093);
nand U1528 (N_1528,In_1986,In_806);
and U1529 (N_1529,In_28,In_1781);
or U1530 (N_1530,In_2372,In_1667);
or U1531 (N_1531,In_1667,In_2421);
nand U1532 (N_1532,In_1640,In_1620);
nor U1533 (N_1533,In_74,In_2311);
nand U1534 (N_1534,In_2481,In_1789);
or U1535 (N_1535,In_43,In_435);
nand U1536 (N_1536,In_99,In_1450);
or U1537 (N_1537,In_1154,In_708);
nand U1538 (N_1538,In_1269,In_2052);
xnor U1539 (N_1539,In_703,In_2232);
and U1540 (N_1540,In_2162,In_1556);
and U1541 (N_1541,In_1563,In_1824);
nand U1542 (N_1542,In_466,In_1564);
or U1543 (N_1543,In_1267,In_318);
and U1544 (N_1544,In_2398,In_126);
nand U1545 (N_1545,In_2455,In_817);
nand U1546 (N_1546,In_2430,In_2392);
or U1547 (N_1547,In_2182,In_901);
xnor U1548 (N_1548,In_277,In_1167);
nand U1549 (N_1549,In_1123,In_946);
or U1550 (N_1550,In_2184,In_2462);
and U1551 (N_1551,In_1740,In_2164);
xnor U1552 (N_1552,In_1316,In_584);
or U1553 (N_1553,In_425,In_322);
and U1554 (N_1554,In_1726,In_1385);
and U1555 (N_1555,In_2193,In_256);
or U1556 (N_1556,In_916,In_703);
and U1557 (N_1557,In_1947,In_1770);
nand U1558 (N_1558,In_741,In_1490);
xnor U1559 (N_1559,In_2298,In_1386);
nor U1560 (N_1560,In_865,In_2242);
xnor U1561 (N_1561,In_917,In_364);
xor U1562 (N_1562,In_1463,In_1664);
and U1563 (N_1563,In_988,In_1062);
nor U1564 (N_1564,In_247,In_2210);
xor U1565 (N_1565,In_444,In_595);
nand U1566 (N_1566,In_873,In_848);
xnor U1567 (N_1567,In_1596,In_767);
and U1568 (N_1568,In_2298,In_1760);
nand U1569 (N_1569,In_1294,In_68);
nor U1570 (N_1570,In_2492,In_2160);
and U1571 (N_1571,In_2304,In_291);
or U1572 (N_1572,In_348,In_831);
nand U1573 (N_1573,In_2,In_2332);
and U1574 (N_1574,In_1714,In_1244);
and U1575 (N_1575,In_109,In_1504);
nor U1576 (N_1576,In_1723,In_2129);
nand U1577 (N_1577,In_24,In_1426);
xor U1578 (N_1578,In_764,In_1019);
xnor U1579 (N_1579,In_2372,In_558);
xor U1580 (N_1580,In_1408,In_148);
xnor U1581 (N_1581,In_2290,In_1965);
nand U1582 (N_1582,In_1771,In_900);
and U1583 (N_1583,In_821,In_660);
xnor U1584 (N_1584,In_1396,In_1264);
nor U1585 (N_1585,In_699,In_1322);
nor U1586 (N_1586,In_118,In_1339);
or U1587 (N_1587,In_1099,In_2319);
and U1588 (N_1588,In_1956,In_2285);
nor U1589 (N_1589,In_1170,In_238);
xor U1590 (N_1590,In_346,In_531);
and U1591 (N_1591,In_1341,In_1442);
and U1592 (N_1592,In_1324,In_1087);
and U1593 (N_1593,In_1054,In_1329);
and U1594 (N_1594,In_1043,In_715);
nor U1595 (N_1595,In_1310,In_2290);
and U1596 (N_1596,In_2179,In_1001);
and U1597 (N_1597,In_961,In_2050);
and U1598 (N_1598,In_1320,In_892);
xor U1599 (N_1599,In_1083,In_1226);
xnor U1600 (N_1600,In_1484,In_772);
or U1601 (N_1601,In_1497,In_1074);
and U1602 (N_1602,In_384,In_726);
or U1603 (N_1603,In_948,In_2404);
nand U1604 (N_1604,In_1393,In_696);
nand U1605 (N_1605,In_1985,In_154);
or U1606 (N_1606,In_1741,In_1935);
nor U1607 (N_1607,In_1245,In_690);
and U1608 (N_1608,In_1858,In_337);
and U1609 (N_1609,In_419,In_2124);
or U1610 (N_1610,In_1083,In_2074);
or U1611 (N_1611,In_1898,In_440);
xnor U1612 (N_1612,In_2458,In_1724);
xor U1613 (N_1613,In_107,In_267);
nor U1614 (N_1614,In_1424,In_2199);
nor U1615 (N_1615,In_2246,In_747);
or U1616 (N_1616,In_153,In_1556);
or U1617 (N_1617,In_2333,In_1953);
or U1618 (N_1618,In_987,In_2134);
xnor U1619 (N_1619,In_1129,In_2285);
nand U1620 (N_1620,In_102,In_2364);
and U1621 (N_1621,In_1234,In_1953);
xnor U1622 (N_1622,In_349,In_313);
and U1623 (N_1623,In_1880,In_1245);
and U1624 (N_1624,In_820,In_190);
and U1625 (N_1625,In_2430,In_938);
nor U1626 (N_1626,In_1719,In_497);
or U1627 (N_1627,In_885,In_321);
and U1628 (N_1628,In_2048,In_1538);
nand U1629 (N_1629,In_580,In_1234);
and U1630 (N_1630,In_1866,In_1631);
and U1631 (N_1631,In_1450,In_1635);
xnor U1632 (N_1632,In_2130,In_1853);
nand U1633 (N_1633,In_76,In_1334);
and U1634 (N_1634,In_1964,In_1768);
nor U1635 (N_1635,In_665,In_920);
or U1636 (N_1636,In_214,In_1242);
nand U1637 (N_1637,In_554,In_1584);
nor U1638 (N_1638,In_2018,In_1229);
nand U1639 (N_1639,In_248,In_1102);
and U1640 (N_1640,In_822,In_1371);
or U1641 (N_1641,In_2298,In_2305);
or U1642 (N_1642,In_735,In_2300);
xor U1643 (N_1643,In_1739,In_964);
nand U1644 (N_1644,In_554,In_2438);
or U1645 (N_1645,In_9,In_959);
nand U1646 (N_1646,In_782,In_65);
and U1647 (N_1647,In_1993,In_2406);
and U1648 (N_1648,In_1196,In_2283);
or U1649 (N_1649,In_1891,In_1942);
xnor U1650 (N_1650,In_408,In_268);
nand U1651 (N_1651,In_2130,In_71);
xnor U1652 (N_1652,In_471,In_858);
nand U1653 (N_1653,In_2174,In_232);
xnor U1654 (N_1654,In_542,In_1342);
and U1655 (N_1655,In_2173,In_1637);
xnor U1656 (N_1656,In_728,In_155);
and U1657 (N_1657,In_1402,In_2465);
nand U1658 (N_1658,In_1545,In_1687);
and U1659 (N_1659,In_2489,In_827);
nand U1660 (N_1660,In_583,In_366);
xnor U1661 (N_1661,In_1620,In_1529);
nor U1662 (N_1662,In_1784,In_723);
nand U1663 (N_1663,In_849,In_1571);
nor U1664 (N_1664,In_11,In_29);
and U1665 (N_1665,In_1127,In_1410);
nand U1666 (N_1666,In_317,In_815);
xnor U1667 (N_1667,In_1612,In_186);
nand U1668 (N_1668,In_219,In_2359);
and U1669 (N_1669,In_839,In_1353);
xor U1670 (N_1670,In_2185,In_381);
and U1671 (N_1671,In_771,In_2431);
nor U1672 (N_1672,In_1554,In_495);
nand U1673 (N_1673,In_788,In_41);
xor U1674 (N_1674,In_2482,In_2470);
or U1675 (N_1675,In_1207,In_2109);
nand U1676 (N_1676,In_1154,In_152);
or U1677 (N_1677,In_44,In_2483);
nor U1678 (N_1678,In_953,In_525);
or U1679 (N_1679,In_936,In_2117);
nand U1680 (N_1680,In_1588,In_1431);
nand U1681 (N_1681,In_742,In_1862);
nor U1682 (N_1682,In_2088,In_166);
nand U1683 (N_1683,In_2248,In_1611);
xor U1684 (N_1684,In_2431,In_1514);
and U1685 (N_1685,In_718,In_2295);
nand U1686 (N_1686,In_908,In_567);
nand U1687 (N_1687,In_1314,In_627);
nand U1688 (N_1688,In_2178,In_64);
nor U1689 (N_1689,In_219,In_2164);
and U1690 (N_1690,In_2213,In_2393);
nand U1691 (N_1691,In_404,In_1511);
nor U1692 (N_1692,In_2271,In_670);
and U1693 (N_1693,In_1198,In_2171);
nand U1694 (N_1694,In_1902,In_1184);
nand U1695 (N_1695,In_250,In_245);
nand U1696 (N_1696,In_2200,In_600);
nand U1697 (N_1697,In_2323,In_914);
nor U1698 (N_1698,In_1274,In_1801);
or U1699 (N_1699,In_2456,In_2309);
or U1700 (N_1700,In_2005,In_1976);
or U1701 (N_1701,In_1429,In_498);
nand U1702 (N_1702,In_1201,In_221);
and U1703 (N_1703,In_1678,In_1350);
nand U1704 (N_1704,In_2100,In_1829);
or U1705 (N_1705,In_575,In_597);
xnor U1706 (N_1706,In_1457,In_2461);
nand U1707 (N_1707,In_1405,In_678);
xor U1708 (N_1708,In_614,In_470);
nand U1709 (N_1709,In_414,In_2499);
nor U1710 (N_1710,In_26,In_2390);
or U1711 (N_1711,In_1842,In_2145);
or U1712 (N_1712,In_2202,In_1016);
nor U1713 (N_1713,In_80,In_191);
xnor U1714 (N_1714,In_22,In_1635);
nand U1715 (N_1715,In_633,In_1010);
xnor U1716 (N_1716,In_809,In_2172);
or U1717 (N_1717,In_1169,In_1867);
xor U1718 (N_1718,In_662,In_1277);
and U1719 (N_1719,In_1736,In_219);
or U1720 (N_1720,In_1427,In_1291);
nand U1721 (N_1721,In_259,In_2115);
nor U1722 (N_1722,In_2455,In_1747);
nand U1723 (N_1723,In_664,In_161);
nand U1724 (N_1724,In_1338,In_2271);
xnor U1725 (N_1725,In_1464,In_2309);
nor U1726 (N_1726,In_1947,In_734);
nand U1727 (N_1727,In_212,In_859);
and U1728 (N_1728,In_1800,In_57);
xor U1729 (N_1729,In_1576,In_1525);
and U1730 (N_1730,In_1977,In_1020);
xor U1731 (N_1731,In_1922,In_909);
or U1732 (N_1732,In_2423,In_1328);
nand U1733 (N_1733,In_2032,In_184);
xor U1734 (N_1734,In_105,In_119);
nand U1735 (N_1735,In_788,In_2386);
nor U1736 (N_1736,In_2133,In_1866);
nand U1737 (N_1737,In_488,In_1075);
nand U1738 (N_1738,In_795,In_111);
xnor U1739 (N_1739,In_2390,In_1361);
nor U1740 (N_1740,In_771,In_1235);
and U1741 (N_1741,In_237,In_189);
xnor U1742 (N_1742,In_1299,In_910);
and U1743 (N_1743,In_2345,In_1426);
or U1744 (N_1744,In_1414,In_2392);
nor U1745 (N_1745,In_2458,In_1057);
or U1746 (N_1746,In_724,In_2429);
xnor U1747 (N_1747,In_867,In_1569);
or U1748 (N_1748,In_468,In_1722);
or U1749 (N_1749,In_1579,In_1274);
nor U1750 (N_1750,In_2090,In_842);
or U1751 (N_1751,In_443,In_1757);
and U1752 (N_1752,In_1573,In_558);
and U1753 (N_1753,In_1215,In_205);
nor U1754 (N_1754,In_2326,In_1178);
xor U1755 (N_1755,In_2195,In_300);
or U1756 (N_1756,In_2100,In_1280);
and U1757 (N_1757,In_1112,In_1965);
or U1758 (N_1758,In_1350,In_2432);
or U1759 (N_1759,In_2307,In_986);
and U1760 (N_1760,In_1226,In_1172);
xnor U1761 (N_1761,In_2249,In_787);
or U1762 (N_1762,In_442,In_1701);
nor U1763 (N_1763,In_706,In_1203);
xnor U1764 (N_1764,In_996,In_1404);
xor U1765 (N_1765,In_1268,In_1773);
nand U1766 (N_1766,In_2395,In_1246);
nor U1767 (N_1767,In_293,In_67);
nand U1768 (N_1768,In_1810,In_1518);
nand U1769 (N_1769,In_457,In_2494);
or U1770 (N_1770,In_1492,In_1893);
xor U1771 (N_1771,In_2469,In_2247);
xnor U1772 (N_1772,In_1417,In_104);
or U1773 (N_1773,In_1822,In_1043);
or U1774 (N_1774,In_1945,In_1482);
xor U1775 (N_1775,In_271,In_16);
and U1776 (N_1776,In_916,In_805);
xnor U1777 (N_1777,In_562,In_908);
nand U1778 (N_1778,In_860,In_686);
nand U1779 (N_1779,In_1841,In_426);
xnor U1780 (N_1780,In_1160,In_542);
xor U1781 (N_1781,In_424,In_92);
nand U1782 (N_1782,In_128,In_2293);
and U1783 (N_1783,In_1601,In_1804);
or U1784 (N_1784,In_1252,In_2252);
and U1785 (N_1785,In_2300,In_1019);
or U1786 (N_1786,In_1416,In_991);
xnor U1787 (N_1787,In_1747,In_636);
xor U1788 (N_1788,In_1095,In_2363);
nor U1789 (N_1789,In_1417,In_164);
and U1790 (N_1790,In_649,In_1318);
nand U1791 (N_1791,In_2203,In_1579);
xor U1792 (N_1792,In_905,In_2007);
nand U1793 (N_1793,In_1062,In_28);
and U1794 (N_1794,In_1158,In_492);
nor U1795 (N_1795,In_319,In_1799);
or U1796 (N_1796,In_775,In_1089);
or U1797 (N_1797,In_33,In_854);
xor U1798 (N_1798,In_486,In_2346);
nand U1799 (N_1799,In_807,In_2338);
nand U1800 (N_1800,In_413,In_134);
and U1801 (N_1801,In_783,In_321);
xor U1802 (N_1802,In_2314,In_1729);
xnor U1803 (N_1803,In_1198,In_337);
or U1804 (N_1804,In_1007,In_1057);
or U1805 (N_1805,In_1013,In_801);
or U1806 (N_1806,In_63,In_142);
or U1807 (N_1807,In_2473,In_2424);
nor U1808 (N_1808,In_1618,In_1706);
nor U1809 (N_1809,In_1864,In_1022);
and U1810 (N_1810,In_267,In_2462);
or U1811 (N_1811,In_2462,In_1856);
and U1812 (N_1812,In_1891,In_2256);
xor U1813 (N_1813,In_619,In_1212);
nor U1814 (N_1814,In_298,In_200);
xnor U1815 (N_1815,In_1161,In_2077);
and U1816 (N_1816,In_1302,In_1690);
nand U1817 (N_1817,In_972,In_1075);
xor U1818 (N_1818,In_2217,In_2267);
or U1819 (N_1819,In_1740,In_273);
nor U1820 (N_1820,In_743,In_352);
or U1821 (N_1821,In_1296,In_1607);
nor U1822 (N_1822,In_1237,In_616);
and U1823 (N_1823,In_1322,In_1175);
or U1824 (N_1824,In_325,In_460);
xnor U1825 (N_1825,In_551,In_2073);
xor U1826 (N_1826,In_2147,In_233);
or U1827 (N_1827,In_596,In_1631);
xor U1828 (N_1828,In_2074,In_1581);
or U1829 (N_1829,In_508,In_199);
nor U1830 (N_1830,In_1477,In_705);
or U1831 (N_1831,In_1869,In_1879);
or U1832 (N_1832,In_965,In_109);
nor U1833 (N_1833,In_100,In_2331);
or U1834 (N_1834,In_1823,In_142);
xnor U1835 (N_1835,In_2114,In_60);
or U1836 (N_1836,In_502,In_2089);
nand U1837 (N_1837,In_2465,In_1444);
or U1838 (N_1838,In_726,In_717);
xnor U1839 (N_1839,In_571,In_1931);
nor U1840 (N_1840,In_839,In_1139);
nor U1841 (N_1841,In_525,In_1367);
nor U1842 (N_1842,In_2193,In_1526);
xor U1843 (N_1843,In_1881,In_1753);
nand U1844 (N_1844,In_153,In_406);
nor U1845 (N_1845,In_567,In_417);
nor U1846 (N_1846,In_2068,In_1303);
or U1847 (N_1847,In_2251,In_2240);
nand U1848 (N_1848,In_451,In_1528);
xor U1849 (N_1849,In_247,In_2389);
or U1850 (N_1850,In_240,In_1484);
or U1851 (N_1851,In_1565,In_1626);
nand U1852 (N_1852,In_1159,In_1826);
nand U1853 (N_1853,In_2398,In_2247);
xor U1854 (N_1854,In_86,In_196);
xor U1855 (N_1855,In_1092,In_948);
nor U1856 (N_1856,In_2474,In_530);
nand U1857 (N_1857,In_1862,In_2040);
and U1858 (N_1858,In_271,In_1391);
and U1859 (N_1859,In_1377,In_1515);
and U1860 (N_1860,In_2461,In_442);
nor U1861 (N_1861,In_853,In_244);
nand U1862 (N_1862,In_1554,In_320);
nand U1863 (N_1863,In_718,In_2215);
nand U1864 (N_1864,In_765,In_515);
xnor U1865 (N_1865,In_1717,In_616);
xor U1866 (N_1866,In_302,In_2091);
nor U1867 (N_1867,In_606,In_593);
xnor U1868 (N_1868,In_848,In_2120);
nand U1869 (N_1869,In_298,In_2083);
or U1870 (N_1870,In_1531,In_1828);
nor U1871 (N_1871,In_1264,In_1016);
nand U1872 (N_1872,In_1483,In_1688);
nand U1873 (N_1873,In_1034,In_2159);
nand U1874 (N_1874,In_922,In_1656);
or U1875 (N_1875,In_459,In_1466);
or U1876 (N_1876,In_1156,In_2475);
and U1877 (N_1877,In_1126,In_271);
xnor U1878 (N_1878,In_2463,In_1795);
nand U1879 (N_1879,In_1455,In_1918);
nor U1880 (N_1880,In_731,In_512);
and U1881 (N_1881,In_38,In_2278);
or U1882 (N_1882,In_261,In_104);
nand U1883 (N_1883,In_1639,In_1085);
xor U1884 (N_1884,In_2267,In_395);
or U1885 (N_1885,In_513,In_1787);
nand U1886 (N_1886,In_1721,In_2029);
xor U1887 (N_1887,In_2411,In_1287);
xor U1888 (N_1888,In_2049,In_1938);
and U1889 (N_1889,In_1111,In_2173);
and U1890 (N_1890,In_446,In_17);
and U1891 (N_1891,In_613,In_486);
nand U1892 (N_1892,In_1503,In_897);
nand U1893 (N_1893,In_1869,In_2133);
nor U1894 (N_1894,In_1415,In_1300);
and U1895 (N_1895,In_1997,In_1506);
and U1896 (N_1896,In_816,In_1150);
xnor U1897 (N_1897,In_1430,In_2072);
xor U1898 (N_1898,In_530,In_794);
or U1899 (N_1899,In_900,In_1192);
and U1900 (N_1900,In_723,In_2430);
or U1901 (N_1901,In_78,In_1036);
and U1902 (N_1902,In_2180,In_1539);
and U1903 (N_1903,In_902,In_2134);
and U1904 (N_1904,In_1930,In_1823);
nand U1905 (N_1905,In_1882,In_1133);
nand U1906 (N_1906,In_1956,In_1531);
and U1907 (N_1907,In_2411,In_2378);
xnor U1908 (N_1908,In_2195,In_385);
and U1909 (N_1909,In_1294,In_1346);
and U1910 (N_1910,In_1481,In_443);
xor U1911 (N_1911,In_1916,In_498);
and U1912 (N_1912,In_1181,In_433);
and U1913 (N_1913,In_1007,In_517);
or U1914 (N_1914,In_1592,In_2148);
xor U1915 (N_1915,In_2360,In_2413);
nand U1916 (N_1916,In_616,In_1572);
or U1917 (N_1917,In_180,In_1080);
or U1918 (N_1918,In_86,In_1339);
nand U1919 (N_1919,In_1533,In_455);
xor U1920 (N_1920,In_1467,In_136);
or U1921 (N_1921,In_1259,In_298);
and U1922 (N_1922,In_515,In_382);
and U1923 (N_1923,In_1103,In_2293);
or U1924 (N_1924,In_1636,In_1669);
and U1925 (N_1925,In_2172,In_1446);
xor U1926 (N_1926,In_1715,In_802);
nor U1927 (N_1927,In_6,In_1252);
nand U1928 (N_1928,In_784,In_697);
or U1929 (N_1929,In_1636,In_2087);
xnor U1930 (N_1930,In_1104,In_100);
and U1931 (N_1931,In_28,In_2287);
and U1932 (N_1932,In_2396,In_692);
nor U1933 (N_1933,In_100,In_949);
nor U1934 (N_1934,In_482,In_325);
and U1935 (N_1935,In_774,In_285);
and U1936 (N_1936,In_2413,In_915);
nor U1937 (N_1937,In_503,In_324);
nor U1938 (N_1938,In_1708,In_889);
or U1939 (N_1939,In_1890,In_2029);
and U1940 (N_1940,In_2413,In_2027);
nor U1941 (N_1941,In_881,In_42);
and U1942 (N_1942,In_1265,In_743);
or U1943 (N_1943,In_234,In_1385);
nor U1944 (N_1944,In_2185,In_558);
xnor U1945 (N_1945,In_751,In_2276);
or U1946 (N_1946,In_2281,In_2222);
and U1947 (N_1947,In_2124,In_497);
xnor U1948 (N_1948,In_2354,In_1143);
nor U1949 (N_1949,In_169,In_321);
or U1950 (N_1950,In_321,In_2457);
nor U1951 (N_1951,In_1242,In_207);
nor U1952 (N_1952,In_1961,In_2070);
nand U1953 (N_1953,In_1623,In_665);
nand U1954 (N_1954,In_1017,In_318);
nand U1955 (N_1955,In_1532,In_1384);
xnor U1956 (N_1956,In_1908,In_2117);
nor U1957 (N_1957,In_776,In_670);
nand U1958 (N_1958,In_1225,In_843);
nor U1959 (N_1959,In_709,In_827);
or U1960 (N_1960,In_374,In_2403);
nor U1961 (N_1961,In_493,In_741);
or U1962 (N_1962,In_1817,In_729);
xor U1963 (N_1963,In_326,In_1180);
or U1964 (N_1964,In_411,In_2457);
nand U1965 (N_1965,In_667,In_520);
or U1966 (N_1966,In_1146,In_848);
or U1967 (N_1967,In_139,In_2245);
nor U1968 (N_1968,In_1577,In_1803);
or U1969 (N_1969,In_1452,In_1047);
or U1970 (N_1970,In_2435,In_239);
xor U1971 (N_1971,In_264,In_586);
and U1972 (N_1972,In_2442,In_752);
nor U1973 (N_1973,In_867,In_2288);
nor U1974 (N_1974,In_1162,In_184);
and U1975 (N_1975,In_1291,In_1530);
nor U1976 (N_1976,In_849,In_444);
xnor U1977 (N_1977,In_1575,In_965);
or U1978 (N_1978,In_1350,In_2027);
nor U1979 (N_1979,In_1140,In_1945);
and U1980 (N_1980,In_252,In_686);
or U1981 (N_1981,In_636,In_2091);
and U1982 (N_1982,In_421,In_2294);
or U1983 (N_1983,In_409,In_13);
and U1984 (N_1984,In_1684,In_430);
or U1985 (N_1985,In_1897,In_2126);
or U1986 (N_1986,In_2101,In_2256);
nand U1987 (N_1987,In_1626,In_2028);
xnor U1988 (N_1988,In_2439,In_86);
nor U1989 (N_1989,In_2188,In_1533);
and U1990 (N_1990,In_773,In_379);
xnor U1991 (N_1991,In_452,In_1968);
nand U1992 (N_1992,In_1714,In_2100);
and U1993 (N_1993,In_81,In_2102);
xor U1994 (N_1994,In_45,In_1286);
xnor U1995 (N_1995,In_872,In_273);
nand U1996 (N_1996,In_638,In_2023);
and U1997 (N_1997,In_383,In_2013);
nor U1998 (N_1998,In_2368,In_1265);
nand U1999 (N_1999,In_713,In_773);
xor U2000 (N_2000,In_568,In_361);
and U2001 (N_2001,In_1977,In_1681);
xnor U2002 (N_2002,In_1221,In_2252);
xnor U2003 (N_2003,In_761,In_437);
nand U2004 (N_2004,In_1476,In_2262);
or U2005 (N_2005,In_1835,In_2365);
xnor U2006 (N_2006,In_1237,In_1562);
nor U2007 (N_2007,In_1543,In_201);
or U2008 (N_2008,In_1773,In_1728);
nand U2009 (N_2009,In_827,In_212);
and U2010 (N_2010,In_13,In_1886);
nor U2011 (N_2011,In_1455,In_1744);
nor U2012 (N_2012,In_1858,In_990);
xor U2013 (N_2013,In_1928,In_1100);
nor U2014 (N_2014,In_1377,In_1479);
nor U2015 (N_2015,In_1518,In_794);
nor U2016 (N_2016,In_1703,In_1831);
nand U2017 (N_2017,In_940,In_853);
xor U2018 (N_2018,In_74,In_665);
or U2019 (N_2019,In_1878,In_822);
xor U2020 (N_2020,In_747,In_1306);
or U2021 (N_2021,In_302,In_684);
or U2022 (N_2022,In_2179,In_591);
or U2023 (N_2023,In_20,In_2491);
xnor U2024 (N_2024,In_999,In_709);
nand U2025 (N_2025,In_107,In_1444);
or U2026 (N_2026,In_1070,In_973);
xor U2027 (N_2027,In_1729,In_1827);
nand U2028 (N_2028,In_20,In_1375);
and U2029 (N_2029,In_1255,In_575);
nor U2030 (N_2030,In_122,In_737);
or U2031 (N_2031,In_33,In_13);
xor U2032 (N_2032,In_644,In_2318);
and U2033 (N_2033,In_797,In_1862);
xor U2034 (N_2034,In_1900,In_2148);
nand U2035 (N_2035,In_1379,In_985);
and U2036 (N_2036,In_1165,In_2399);
nor U2037 (N_2037,In_2282,In_1729);
or U2038 (N_2038,In_1625,In_988);
or U2039 (N_2039,In_290,In_873);
nor U2040 (N_2040,In_1417,In_955);
and U2041 (N_2041,In_1991,In_2077);
xnor U2042 (N_2042,In_777,In_820);
nor U2043 (N_2043,In_2337,In_523);
and U2044 (N_2044,In_2403,In_521);
nor U2045 (N_2045,In_1061,In_618);
nor U2046 (N_2046,In_1642,In_750);
or U2047 (N_2047,In_48,In_1508);
or U2048 (N_2048,In_147,In_1387);
xnor U2049 (N_2049,In_2193,In_800);
xnor U2050 (N_2050,In_668,In_263);
and U2051 (N_2051,In_1552,In_1755);
and U2052 (N_2052,In_503,In_465);
nor U2053 (N_2053,In_577,In_717);
nand U2054 (N_2054,In_2314,In_248);
or U2055 (N_2055,In_116,In_207);
nand U2056 (N_2056,In_842,In_1893);
nand U2057 (N_2057,In_1672,In_23);
nand U2058 (N_2058,In_710,In_1030);
nand U2059 (N_2059,In_340,In_264);
nor U2060 (N_2060,In_1829,In_1250);
xnor U2061 (N_2061,In_1123,In_363);
xnor U2062 (N_2062,In_1558,In_1821);
nor U2063 (N_2063,In_970,In_1004);
nor U2064 (N_2064,In_1667,In_1265);
xor U2065 (N_2065,In_1277,In_684);
or U2066 (N_2066,In_649,In_1907);
and U2067 (N_2067,In_1340,In_515);
and U2068 (N_2068,In_73,In_1467);
or U2069 (N_2069,In_2445,In_443);
or U2070 (N_2070,In_585,In_2395);
xor U2071 (N_2071,In_1388,In_171);
or U2072 (N_2072,In_1077,In_1400);
and U2073 (N_2073,In_2468,In_2217);
nand U2074 (N_2074,In_311,In_353);
nand U2075 (N_2075,In_717,In_522);
or U2076 (N_2076,In_920,In_1485);
nand U2077 (N_2077,In_2115,In_1599);
nand U2078 (N_2078,In_1099,In_1715);
nor U2079 (N_2079,In_1813,In_250);
and U2080 (N_2080,In_2268,In_1487);
nand U2081 (N_2081,In_1494,In_659);
or U2082 (N_2082,In_211,In_373);
nor U2083 (N_2083,In_531,In_2388);
or U2084 (N_2084,In_2212,In_2095);
nor U2085 (N_2085,In_1959,In_1652);
xor U2086 (N_2086,In_2226,In_2044);
and U2087 (N_2087,In_830,In_339);
nor U2088 (N_2088,In_998,In_377);
nor U2089 (N_2089,In_1588,In_507);
and U2090 (N_2090,In_657,In_2356);
xnor U2091 (N_2091,In_463,In_443);
or U2092 (N_2092,In_1845,In_795);
and U2093 (N_2093,In_1132,In_446);
or U2094 (N_2094,In_1634,In_2027);
nand U2095 (N_2095,In_3,In_2337);
and U2096 (N_2096,In_1547,In_2429);
or U2097 (N_2097,In_2300,In_1609);
nor U2098 (N_2098,In_1036,In_1850);
nand U2099 (N_2099,In_1182,In_1369);
xnor U2100 (N_2100,In_265,In_1763);
or U2101 (N_2101,In_1854,In_391);
nor U2102 (N_2102,In_1761,In_701);
or U2103 (N_2103,In_1859,In_34);
or U2104 (N_2104,In_1581,In_1896);
or U2105 (N_2105,In_1055,In_1513);
nor U2106 (N_2106,In_648,In_1554);
or U2107 (N_2107,In_291,In_1576);
and U2108 (N_2108,In_1410,In_1163);
nand U2109 (N_2109,In_1541,In_1159);
xnor U2110 (N_2110,In_2461,In_511);
nand U2111 (N_2111,In_853,In_1969);
or U2112 (N_2112,In_1563,In_1409);
xor U2113 (N_2113,In_1805,In_1609);
or U2114 (N_2114,In_222,In_347);
xnor U2115 (N_2115,In_2132,In_977);
or U2116 (N_2116,In_1888,In_1706);
xor U2117 (N_2117,In_1362,In_1572);
nand U2118 (N_2118,In_2067,In_726);
nor U2119 (N_2119,In_318,In_638);
or U2120 (N_2120,In_2490,In_521);
nor U2121 (N_2121,In_1721,In_1762);
xnor U2122 (N_2122,In_1488,In_673);
xnor U2123 (N_2123,In_1540,In_1312);
or U2124 (N_2124,In_559,In_1399);
and U2125 (N_2125,In_1662,In_530);
nor U2126 (N_2126,In_2029,In_1360);
nand U2127 (N_2127,In_1882,In_1235);
or U2128 (N_2128,In_693,In_2260);
nor U2129 (N_2129,In_712,In_2431);
xnor U2130 (N_2130,In_475,In_385);
nor U2131 (N_2131,In_719,In_1632);
xor U2132 (N_2132,In_1324,In_2329);
nor U2133 (N_2133,In_298,In_837);
nand U2134 (N_2134,In_1435,In_520);
nand U2135 (N_2135,In_180,In_378);
or U2136 (N_2136,In_964,In_737);
xor U2137 (N_2137,In_765,In_1978);
nor U2138 (N_2138,In_1263,In_1427);
or U2139 (N_2139,In_1260,In_303);
xnor U2140 (N_2140,In_306,In_1705);
and U2141 (N_2141,In_2418,In_735);
or U2142 (N_2142,In_106,In_1086);
nand U2143 (N_2143,In_2411,In_1754);
and U2144 (N_2144,In_1060,In_1147);
xnor U2145 (N_2145,In_248,In_2219);
and U2146 (N_2146,In_1546,In_1913);
nor U2147 (N_2147,In_1698,In_95);
or U2148 (N_2148,In_1588,In_397);
nand U2149 (N_2149,In_139,In_111);
xor U2150 (N_2150,In_1296,In_824);
or U2151 (N_2151,In_1282,In_1935);
nor U2152 (N_2152,In_897,In_1181);
xnor U2153 (N_2153,In_665,In_329);
and U2154 (N_2154,In_874,In_973);
and U2155 (N_2155,In_1676,In_461);
and U2156 (N_2156,In_2363,In_1223);
and U2157 (N_2157,In_125,In_1947);
nor U2158 (N_2158,In_1471,In_753);
or U2159 (N_2159,In_593,In_812);
xnor U2160 (N_2160,In_1251,In_372);
nor U2161 (N_2161,In_934,In_1346);
nand U2162 (N_2162,In_232,In_2423);
xnor U2163 (N_2163,In_2357,In_1765);
and U2164 (N_2164,In_1574,In_548);
or U2165 (N_2165,In_372,In_604);
nand U2166 (N_2166,In_1235,In_1713);
nand U2167 (N_2167,In_734,In_1284);
nand U2168 (N_2168,In_1562,In_1528);
nor U2169 (N_2169,In_408,In_1103);
and U2170 (N_2170,In_585,In_1699);
xor U2171 (N_2171,In_766,In_2377);
and U2172 (N_2172,In_2395,In_1170);
xnor U2173 (N_2173,In_2274,In_2232);
or U2174 (N_2174,In_2372,In_465);
or U2175 (N_2175,In_2280,In_803);
nor U2176 (N_2176,In_2404,In_1581);
nor U2177 (N_2177,In_1387,In_1803);
nor U2178 (N_2178,In_2061,In_927);
and U2179 (N_2179,In_2327,In_1909);
nand U2180 (N_2180,In_1608,In_626);
or U2181 (N_2181,In_545,In_262);
nand U2182 (N_2182,In_1576,In_2490);
or U2183 (N_2183,In_1345,In_209);
and U2184 (N_2184,In_181,In_2115);
and U2185 (N_2185,In_257,In_834);
and U2186 (N_2186,In_676,In_461);
nor U2187 (N_2187,In_260,In_651);
xor U2188 (N_2188,In_1613,In_2128);
xor U2189 (N_2189,In_1607,In_114);
nand U2190 (N_2190,In_233,In_2329);
xor U2191 (N_2191,In_2446,In_1695);
or U2192 (N_2192,In_934,In_391);
or U2193 (N_2193,In_7,In_302);
nand U2194 (N_2194,In_209,In_1633);
nor U2195 (N_2195,In_2026,In_2133);
xnor U2196 (N_2196,In_762,In_307);
nor U2197 (N_2197,In_113,In_196);
nand U2198 (N_2198,In_332,In_195);
xnor U2199 (N_2199,In_1076,In_2477);
nor U2200 (N_2200,In_1976,In_2080);
nand U2201 (N_2201,In_1039,In_2104);
and U2202 (N_2202,In_659,In_2001);
and U2203 (N_2203,In_306,In_292);
nand U2204 (N_2204,In_968,In_1986);
and U2205 (N_2205,In_1354,In_842);
xnor U2206 (N_2206,In_110,In_795);
nand U2207 (N_2207,In_2343,In_1771);
nand U2208 (N_2208,In_2248,In_2096);
nor U2209 (N_2209,In_853,In_954);
or U2210 (N_2210,In_1380,In_1034);
or U2211 (N_2211,In_1054,In_1101);
and U2212 (N_2212,In_378,In_1541);
and U2213 (N_2213,In_595,In_2347);
and U2214 (N_2214,In_169,In_1857);
or U2215 (N_2215,In_2184,In_423);
and U2216 (N_2216,In_866,In_2470);
or U2217 (N_2217,In_289,In_1577);
or U2218 (N_2218,In_51,In_423);
xnor U2219 (N_2219,In_1528,In_2320);
and U2220 (N_2220,In_1860,In_151);
or U2221 (N_2221,In_2130,In_1297);
nand U2222 (N_2222,In_932,In_587);
or U2223 (N_2223,In_411,In_316);
xnor U2224 (N_2224,In_1693,In_1978);
nor U2225 (N_2225,In_790,In_327);
nand U2226 (N_2226,In_653,In_2128);
xor U2227 (N_2227,In_1522,In_1390);
nor U2228 (N_2228,In_118,In_1196);
and U2229 (N_2229,In_2294,In_63);
nand U2230 (N_2230,In_1741,In_2202);
xor U2231 (N_2231,In_2474,In_1717);
nand U2232 (N_2232,In_730,In_193);
xnor U2233 (N_2233,In_78,In_2380);
xor U2234 (N_2234,In_291,In_2378);
nor U2235 (N_2235,In_1359,In_1749);
xnor U2236 (N_2236,In_941,In_117);
or U2237 (N_2237,In_2264,In_1686);
and U2238 (N_2238,In_1451,In_2361);
nor U2239 (N_2239,In_772,In_596);
nand U2240 (N_2240,In_1736,In_1478);
nor U2241 (N_2241,In_1682,In_213);
xor U2242 (N_2242,In_69,In_2124);
nor U2243 (N_2243,In_514,In_1025);
nand U2244 (N_2244,In_1586,In_1552);
nor U2245 (N_2245,In_2104,In_922);
nand U2246 (N_2246,In_1162,In_951);
xor U2247 (N_2247,In_1587,In_1816);
or U2248 (N_2248,In_2339,In_169);
nor U2249 (N_2249,In_546,In_57);
xnor U2250 (N_2250,In_2306,In_76);
or U2251 (N_2251,In_1835,In_1060);
or U2252 (N_2252,In_1796,In_2417);
or U2253 (N_2253,In_2319,In_2085);
xor U2254 (N_2254,In_1037,In_331);
nand U2255 (N_2255,In_968,In_55);
xnor U2256 (N_2256,In_173,In_1769);
xnor U2257 (N_2257,In_36,In_1609);
nand U2258 (N_2258,In_2431,In_2227);
or U2259 (N_2259,In_1587,In_2351);
and U2260 (N_2260,In_1048,In_657);
xnor U2261 (N_2261,In_146,In_1502);
nor U2262 (N_2262,In_1019,In_143);
nor U2263 (N_2263,In_95,In_1696);
and U2264 (N_2264,In_128,In_2287);
and U2265 (N_2265,In_1609,In_1771);
or U2266 (N_2266,In_1151,In_1715);
or U2267 (N_2267,In_2047,In_60);
nand U2268 (N_2268,In_1804,In_2277);
xnor U2269 (N_2269,In_17,In_1002);
nand U2270 (N_2270,In_283,In_738);
or U2271 (N_2271,In_2321,In_2365);
or U2272 (N_2272,In_252,In_338);
nor U2273 (N_2273,In_2060,In_826);
and U2274 (N_2274,In_2360,In_2087);
or U2275 (N_2275,In_2003,In_938);
nand U2276 (N_2276,In_2217,In_1703);
nor U2277 (N_2277,In_965,In_1596);
and U2278 (N_2278,In_1741,In_790);
xnor U2279 (N_2279,In_1946,In_321);
or U2280 (N_2280,In_842,In_583);
nor U2281 (N_2281,In_20,In_2303);
nor U2282 (N_2282,In_517,In_1316);
nand U2283 (N_2283,In_367,In_381);
xnor U2284 (N_2284,In_2141,In_1173);
nand U2285 (N_2285,In_492,In_1966);
and U2286 (N_2286,In_1104,In_1725);
and U2287 (N_2287,In_122,In_1204);
and U2288 (N_2288,In_1462,In_300);
nor U2289 (N_2289,In_2228,In_1913);
nand U2290 (N_2290,In_1319,In_163);
and U2291 (N_2291,In_1232,In_2413);
and U2292 (N_2292,In_556,In_1264);
or U2293 (N_2293,In_2045,In_2161);
nor U2294 (N_2294,In_2493,In_1721);
nor U2295 (N_2295,In_1995,In_804);
and U2296 (N_2296,In_673,In_908);
xnor U2297 (N_2297,In_813,In_1870);
nor U2298 (N_2298,In_234,In_607);
or U2299 (N_2299,In_2116,In_2449);
nand U2300 (N_2300,In_480,In_619);
nor U2301 (N_2301,In_1722,In_2270);
or U2302 (N_2302,In_2250,In_528);
xnor U2303 (N_2303,In_314,In_1299);
or U2304 (N_2304,In_1630,In_1520);
or U2305 (N_2305,In_879,In_2004);
nand U2306 (N_2306,In_727,In_223);
or U2307 (N_2307,In_1099,In_1014);
nand U2308 (N_2308,In_613,In_43);
nor U2309 (N_2309,In_1060,In_1994);
nand U2310 (N_2310,In_1552,In_2114);
and U2311 (N_2311,In_1649,In_99);
nor U2312 (N_2312,In_1832,In_2102);
xnor U2313 (N_2313,In_1235,In_5);
nand U2314 (N_2314,In_191,In_2411);
and U2315 (N_2315,In_1735,In_1095);
xor U2316 (N_2316,In_2351,In_1537);
nor U2317 (N_2317,In_894,In_1988);
nor U2318 (N_2318,In_1691,In_1157);
xnor U2319 (N_2319,In_146,In_1523);
or U2320 (N_2320,In_1722,In_783);
nor U2321 (N_2321,In_2208,In_313);
or U2322 (N_2322,In_2306,In_2080);
nor U2323 (N_2323,In_2119,In_929);
or U2324 (N_2324,In_683,In_1170);
nor U2325 (N_2325,In_1588,In_1099);
nor U2326 (N_2326,In_2069,In_7);
xnor U2327 (N_2327,In_2178,In_1174);
and U2328 (N_2328,In_341,In_223);
nand U2329 (N_2329,In_2472,In_873);
nand U2330 (N_2330,In_1449,In_2333);
and U2331 (N_2331,In_1773,In_464);
xnor U2332 (N_2332,In_1377,In_1438);
nor U2333 (N_2333,In_1870,In_1937);
or U2334 (N_2334,In_1381,In_643);
or U2335 (N_2335,In_74,In_1913);
nand U2336 (N_2336,In_574,In_1055);
nor U2337 (N_2337,In_1227,In_1217);
nor U2338 (N_2338,In_408,In_250);
or U2339 (N_2339,In_2261,In_1092);
nor U2340 (N_2340,In_803,In_1889);
or U2341 (N_2341,In_2304,In_1304);
or U2342 (N_2342,In_1337,In_1280);
and U2343 (N_2343,In_814,In_1535);
and U2344 (N_2344,In_1250,In_876);
xor U2345 (N_2345,In_161,In_1463);
nand U2346 (N_2346,In_463,In_1508);
xor U2347 (N_2347,In_1067,In_2279);
or U2348 (N_2348,In_1020,In_433);
and U2349 (N_2349,In_1765,In_1202);
or U2350 (N_2350,In_1311,In_1956);
xnor U2351 (N_2351,In_1581,In_1477);
or U2352 (N_2352,In_2142,In_7);
or U2353 (N_2353,In_1579,In_1749);
nand U2354 (N_2354,In_1230,In_1732);
and U2355 (N_2355,In_1206,In_938);
nor U2356 (N_2356,In_318,In_501);
nor U2357 (N_2357,In_2364,In_1963);
nor U2358 (N_2358,In_295,In_98);
xor U2359 (N_2359,In_1251,In_89);
nand U2360 (N_2360,In_1790,In_493);
nand U2361 (N_2361,In_996,In_2069);
nand U2362 (N_2362,In_608,In_2383);
and U2363 (N_2363,In_2357,In_1633);
and U2364 (N_2364,In_2072,In_1909);
nor U2365 (N_2365,In_1392,In_1076);
or U2366 (N_2366,In_803,In_364);
nor U2367 (N_2367,In_2283,In_207);
and U2368 (N_2368,In_672,In_2282);
nand U2369 (N_2369,In_2296,In_356);
nand U2370 (N_2370,In_1648,In_2352);
or U2371 (N_2371,In_2158,In_2217);
xor U2372 (N_2372,In_165,In_1679);
xnor U2373 (N_2373,In_2075,In_83);
xor U2374 (N_2374,In_2303,In_1361);
nand U2375 (N_2375,In_1431,In_1272);
or U2376 (N_2376,In_1257,In_1992);
or U2377 (N_2377,In_2148,In_976);
nor U2378 (N_2378,In_366,In_648);
nor U2379 (N_2379,In_1888,In_1649);
or U2380 (N_2380,In_29,In_988);
nand U2381 (N_2381,In_1695,In_1272);
or U2382 (N_2382,In_951,In_320);
nor U2383 (N_2383,In_2214,In_1133);
and U2384 (N_2384,In_283,In_1442);
or U2385 (N_2385,In_1221,In_1922);
or U2386 (N_2386,In_769,In_1137);
xor U2387 (N_2387,In_2027,In_1760);
xnor U2388 (N_2388,In_486,In_1258);
xor U2389 (N_2389,In_46,In_1546);
and U2390 (N_2390,In_2083,In_442);
or U2391 (N_2391,In_175,In_1168);
nand U2392 (N_2392,In_823,In_2288);
nand U2393 (N_2393,In_238,In_527);
and U2394 (N_2394,In_1923,In_634);
and U2395 (N_2395,In_485,In_1984);
and U2396 (N_2396,In_156,In_1977);
xor U2397 (N_2397,In_415,In_2364);
xor U2398 (N_2398,In_1473,In_47);
nand U2399 (N_2399,In_76,In_1557);
and U2400 (N_2400,In_1492,In_2213);
nor U2401 (N_2401,In_1315,In_1953);
and U2402 (N_2402,In_2495,In_1826);
and U2403 (N_2403,In_574,In_2318);
or U2404 (N_2404,In_2491,In_2125);
and U2405 (N_2405,In_1644,In_2207);
or U2406 (N_2406,In_1891,In_765);
and U2407 (N_2407,In_243,In_2240);
xnor U2408 (N_2408,In_235,In_2466);
nor U2409 (N_2409,In_997,In_1392);
nand U2410 (N_2410,In_65,In_1698);
xor U2411 (N_2411,In_2116,In_1683);
or U2412 (N_2412,In_2175,In_2452);
nand U2413 (N_2413,In_2480,In_1974);
nor U2414 (N_2414,In_854,In_2272);
and U2415 (N_2415,In_2191,In_1308);
nand U2416 (N_2416,In_2246,In_831);
or U2417 (N_2417,In_200,In_627);
nor U2418 (N_2418,In_1661,In_1690);
nor U2419 (N_2419,In_77,In_714);
or U2420 (N_2420,In_983,In_2053);
xnor U2421 (N_2421,In_1376,In_1821);
nor U2422 (N_2422,In_2192,In_914);
nand U2423 (N_2423,In_2458,In_8);
xnor U2424 (N_2424,In_428,In_2338);
nand U2425 (N_2425,In_2246,In_343);
and U2426 (N_2426,In_37,In_287);
or U2427 (N_2427,In_238,In_1665);
nor U2428 (N_2428,In_2251,In_2215);
or U2429 (N_2429,In_2205,In_1430);
nor U2430 (N_2430,In_186,In_532);
nor U2431 (N_2431,In_201,In_1151);
nor U2432 (N_2432,In_171,In_2013);
xor U2433 (N_2433,In_1994,In_551);
xnor U2434 (N_2434,In_233,In_993);
and U2435 (N_2435,In_1900,In_847);
nor U2436 (N_2436,In_480,In_1310);
and U2437 (N_2437,In_814,In_1599);
and U2438 (N_2438,In_1135,In_511);
xor U2439 (N_2439,In_2480,In_1148);
xor U2440 (N_2440,In_2155,In_504);
nor U2441 (N_2441,In_770,In_1351);
xor U2442 (N_2442,In_1196,In_367);
and U2443 (N_2443,In_1590,In_1187);
nor U2444 (N_2444,In_2189,In_1773);
nand U2445 (N_2445,In_1538,In_1734);
nand U2446 (N_2446,In_84,In_795);
and U2447 (N_2447,In_1229,In_799);
nor U2448 (N_2448,In_1959,In_700);
nand U2449 (N_2449,In_363,In_2362);
and U2450 (N_2450,In_251,In_885);
or U2451 (N_2451,In_1150,In_980);
xnor U2452 (N_2452,In_1696,In_1095);
nand U2453 (N_2453,In_829,In_213);
or U2454 (N_2454,In_1466,In_1301);
or U2455 (N_2455,In_859,In_2165);
and U2456 (N_2456,In_1184,In_555);
xor U2457 (N_2457,In_774,In_425);
or U2458 (N_2458,In_943,In_883);
xor U2459 (N_2459,In_1794,In_453);
nor U2460 (N_2460,In_1963,In_632);
nand U2461 (N_2461,In_1133,In_2351);
and U2462 (N_2462,In_326,In_1084);
or U2463 (N_2463,In_1664,In_623);
nand U2464 (N_2464,In_291,In_578);
xnor U2465 (N_2465,In_1403,In_656);
and U2466 (N_2466,In_2088,In_1290);
xor U2467 (N_2467,In_2232,In_1721);
or U2468 (N_2468,In_578,In_172);
and U2469 (N_2469,In_331,In_1895);
and U2470 (N_2470,In_1990,In_557);
nand U2471 (N_2471,In_1789,In_751);
nand U2472 (N_2472,In_670,In_2495);
nor U2473 (N_2473,In_2438,In_2275);
nand U2474 (N_2474,In_2497,In_1465);
nor U2475 (N_2475,In_813,In_667);
and U2476 (N_2476,In_358,In_559);
nand U2477 (N_2477,In_780,In_1333);
or U2478 (N_2478,In_1338,In_1625);
nor U2479 (N_2479,In_977,In_803);
or U2480 (N_2480,In_830,In_84);
and U2481 (N_2481,In_42,In_1448);
nor U2482 (N_2482,In_382,In_1204);
nand U2483 (N_2483,In_2415,In_476);
and U2484 (N_2484,In_2492,In_145);
or U2485 (N_2485,In_1175,In_685);
nand U2486 (N_2486,In_2466,In_42);
xor U2487 (N_2487,In_578,In_1870);
or U2488 (N_2488,In_51,In_2457);
xnor U2489 (N_2489,In_306,In_1526);
nand U2490 (N_2490,In_394,In_2424);
xor U2491 (N_2491,In_1762,In_2403);
and U2492 (N_2492,In_1096,In_907);
nand U2493 (N_2493,In_896,In_254);
xor U2494 (N_2494,In_849,In_1223);
or U2495 (N_2495,In_1434,In_2118);
nand U2496 (N_2496,In_2024,In_2487);
xor U2497 (N_2497,In_1483,In_669);
xor U2498 (N_2498,In_1370,In_2217);
or U2499 (N_2499,In_1436,In_551);
and U2500 (N_2500,In_1453,In_894);
nand U2501 (N_2501,In_1068,In_2274);
xor U2502 (N_2502,In_1850,In_2285);
and U2503 (N_2503,In_310,In_566);
or U2504 (N_2504,In_1184,In_2066);
xnor U2505 (N_2505,In_2362,In_2254);
nand U2506 (N_2506,In_634,In_1920);
nor U2507 (N_2507,In_2277,In_1343);
nor U2508 (N_2508,In_2263,In_1675);
nand U2509 (N_2509,In_215,In_961);
nand U2510 (N_2510,In_2207,In_952);
xnor U2511 (N_2511,In_11,In_1376);
nand U2512 (N_2512,In_2215,In_2107);
xor U2513 (N_2513,In_1389,In_1831);
xnor U2514 (N_2514,In_567,In_2246);
or U2515 (N_2515,In_709,In_937);
xor U2516 (N_2516,In_849,In_1208);
or U2517 (N_2517,In_756,In_1974);
or U2518 (N_2518,In_2211,In_1797);
or U2519 (N_2519,In_2129,In_1986);
or U2520 (N_2520,In_2142,In_48);
nor U2521 (N_2521,In_1384,In_2432);
or U2522 (N_2522,In_1045,In_847);
or U2523 (N_2523,In_434,In_435);
and U2524 (N_2524,In_2295,In_1033);
nand U2525 (N_2525,In_184,In_667);
nand U2526 (N_2526,In_2033,In_68);
xor U2527 (N_2527,In_624,In_571);
nor U2528 (N_2528,In_1086,In_2153);
nor U2529 (N_2529,In_1086,In_48);
nor U2530 (N_2530,In_978,In_1892);
nor U2531 (N_2531,In_169,In_705);
nand U2532 (N_2532,In_810,In_651);
or U2533 (N_2533,In_1378,In_849);
nor U2534 (N_2534,In_1491,In_965);
nor U2535 (N_2535,In_98,In_1438);
and U2536 (N_2536,In_231,In_201);
nor U2537 (N_2537,In_254,In_1873);
and U2538 (N_2538,In_1070,In_1092);
xor U2539 (N_2539,In_2142,In_1665);
nand U2540 (N_2540,In_2141,In_2271);
nor U2541 (N_2541,In_1747,In_2073);
nor U2542 (N_2542,In_1688,In_451);
nand U2543 (N_2543,In_607,In_1131);
and U2544 (N_2544,In_521,In_92);
and U2545 (N_2545,In_669,In_892);
nor U2546 (N_2546,In_1131,In_1758);
nand U2547 (N_2547,In_77,In_842);
nand U2548 (N_2548,In_2421,In_2043);
nor U2549 (N_2549,In_1488,In_1962);
xnor U2550 (N_2550,In_769,In_1150);
nor U2551 (N_2551,In_1515,In_372);
nand U2552 (N_2552,In_1923,In_2093);
nor U2553 (N_2553,In_38,In_1892);
nor U2554 (N_2554,In_2378,In_2141);
or U2555 (N_2555,In_1837,In_1173);
nor U2556 (N_2556,In_1563,In_744);
or U2557 (N_2557,In_431,In_2100);
and U2558 (N_2558,In_835,In_684);
xor U2559 (N_2559,In_1322,In_2225);
xnor U2560 (N_2560,In_393,In_1326);
or U2561 (N_2561,In_490,In_1695);
xnor U2562 (N_2562,In_1771,In_137);
nor U2563 (N_2563,In_270,In_140);
xnor U2564 (N_2564,In_1300,In_67);
nand U2565 (N_2565,In_1881,In_733);
or U2566 (N_2566,In_541,In_2495);
and U2567 (N_2567,In_1102,In_1011);
nand U2568 (N_2568,In_2295,In_67);
or U2569 (N_2569,In_551,In_2385);
or U2570 (N_2570,In_2349,In_1403);
and U2571 (N_2571,In_1387,In_1579);
and U2572 (N_2572,In_1381,In_1848);
and U2573 (N_2573,In_2380,In_1778);
nand U2574 (N_2574,In_593,In_1556);
or U2575 (N_2575,In_1139,In_437);
nand U2576 (N_2576,In_1894,In_1583);
or U2577 (N_2577,In_130,In_2414);
or U2578 (N_2578,In_530,In_67);
nand U2579 (N_2579,In_630,In_1837);
and U2580 (N_2580,In_1324,In_18);
or U2581 (N_2581,In_2000,In_1939);
nand U2582 (N_2582,In_410,In_1591);
nor U2583 (N_2583,In_1711,In_2236);
and U2584 (N_2584,In_2453,In_1992);
or U2585 (N_2585,In_1144,In_2121);
and U2586 (N_2586,In_145,In_1268);
and U2587 (N_2587,In_498,In_178);
and U2588 (N_2588,In_1675,In_2348);
nor U2589 (N_2589,In_1765,In_2268);
nor U2590 (N_2590,In_1188,In_799);
nor U2591 (N_2591,In_1522,In_1241);
nand U2592 (N_2592,In_1914,In_1536);
nand U2593 (N_2593,In_331,In_2273);
nand U2594 (N_2594,In_1973,In_1887);
nor U2595 (N_2595,In_1959,In_1638);
nor U2596 (N_2596,In_1916,In_2475);
and U2597 (N_2597,In_1942,In_1358);
nand U2598 (N_2598,In_110,In_1563);
xnor U2599 (N_2599,In_2304,In_118);
and U2600 (N_2600,In_2487,In_1949);
nand U2601 (N_2601,In_1652,In_564);
xnor U2602 (N_2602,In_218,In_735);
nand U2603 (N_2603,In_1148,In_983);
or U2604 (N_2604,In_1349,In_2405);
or U2605 (N_2605,In_1745,In_151);
or U2606 (N_2606,In_290,In_2148);
xnor U2607 (N_2607,In_24,In_502);
nor U2608 (N_2608,In_1216,In_485);
xnor U2609 (N_2609,In_2217,In_1674);
and U2610 (N_2610,In_111,In_1732);
nand U2611 (N_2611,In_759,In_373);
xor U2612 (N_2612,In_2322,In_481);
nor U2613 (N_2613,In_218,In_724);
or U2614 (N_2614,In_1843,In_1553);
or U2615 (N_2615,In_1981,In_460);
xnor U2616 (N_2616,In_661,In_1039);
nor U2617 (N_2617,In_1340,In_1947);
xnor U2618 (N_2618,In_375,In_1756);
xnor U2619 (N_2619,In_2079,In_138);
nand U2620 (N_2620,In_1318,In_1418);
or U2621 (N_2621,In_214,In_1465);
nor U2622 (N_2622,In_1888,In_2065);
xor U2623 (N_2623,In_976,In_1190);
nor U2624 (N_2624,In_1355,In_516);
nor U2625 (N_2625,In_2032,In_413);
xnor U2626 (N_2626,In_1562,In_1801);
nand U2627 (N_2627,In_2430,In_173);
xnor U2628 (N_2628,In_2325,In_1106);
and U2629 (N_2629,In_252,In_2041);
xor U2630 (N_2630,In_2223,In_842);
and U2631 (N_2631,In_1568,In_1667);
nor U2632 (N_2632,In_2409,In_1975);
or U2633 (N_2633,In_2160,In_489);
or U2634 (N_2634,In_278,In_979);
and U2635 (N_2635,In_1630,In_1969);
or U2636 (N_2636,In_815,In_1457);
or U2637 (N_2637,In_1813,In_2190);
and U2638 (N_2638,In_1462,In_617);
nand U2639 (N_2639,In_1263,In_503);
xor U2640 (N_2640,In_834,In_315);
nand U2641 (N_2641,In_42,In_1793);
or U2642 (N_2642,In_1968,In_92);
and U2643 (N_2643,In_1547,In_2448);
nand U2644 (N_2644,In_2215,In_2371);
and U2645 (N_2645,In_1591,In_1830);
nor U2646 (N_2646,In_73,In_2058);
nor U2647 (N_2647,In_736,In_417);
xnor U2648 (N_2648,In_2030,In_1124);
or U2649 (N_2649,In_372,In_1761);
nand U2650 (N_2650,In_1340,In_2285);
nor U2651 (N_2651,In_598,In_1883);
nand U2652 (N_2652,In_2150,In_1285);
nand U2653 (N_2653,In_1833,In_142);
nand U2654 (N_2654,In_521,In_274);
and U2655 (N_2655,In_2182,In_1171);
or U2656 (N_2656,In_1305,In_587);
nand U2657 (N_2657,In_2129,In_2128);
nor U2658 (N_2658,In_1630,In_2439);
and U2659 (N_2659,In_2250,In_2355);
nor U2660 (N_2660,In_877,In_412);
nor U2661 (N_2661,In_1520,In_760);
nand U2662 (N_2662,In_540,In_2365);
xnor U2663 (N_2663,In_235,In_1438);
or U2664 (N_2664,In_2459,In_810);
or U2665 (N_2665,In_630,In_2389);
and U2666 (N_2666,In_1973,In_2239);
or U2667 (N_2667,In_2073,In_783);
nand U2668 (N_2668,In_341,In_451);
nand U2669 (N_2669,In_314,In_1581);
or U2670 (N_2670,In_1986,In_1718);
nand U2671 (N_2671,In_952,In_982);
or U2672 (N_2672,In_2298,In_2409);
xor U2673 (N_2673,In_1957,In_1157);
nand U2674 (N_2674,In_643,In_2029);
and U2675 (N_2675,In_200,In_2332);
nand U2676 (N_2676,In_2105,In_2349);
or U2677 (N_2677,In_2174,In_1546);
nand U2678 (N_2678,In_1463,In_1754);
or U2679 (N_2679,In_2279,In_731);
nand U2680 (N_2680,In_43,In_1552);
nand U2681 (N_2681,In_1071,In_956);
xor U2682 (N_2682,In_2128,In_1615);
xor U2683 (N_2683,In_1238,In_1110);
and U2684 (N_2684,In_833,In_914);
nor U2685 (N_2685,In_789,In_480);
or U2686 (N_2686,In_1151,In_1815);
nand U2687 (N_2687,In_2014,In_896);
nand U2688 (N_2688,In_1406,In_950);
and U2689 (N_2689,In_1148,In_2375);
xnor U2690 (N_2690,In_2427,In_508);
nand U2691 (N_2691,In_666,In_2322);
nor U2692 (N_2692,In_1004,In_893);
nand U2693 (N_2693,In_1961,In_34);
or U2694 (N_2694,In_837,In_829);
xor U2695 (N_2695,In_304,In_1120);
nor U2696 (N_2696,In_69,In_180);
nor U2697 (N_2697,In_56,In_438);
xnor U2698 (N_2698,In_2237,In_1358);
and U2699 (N_2699,In_2032,In_1311);
and U2700 (N_2700,In_218,In_1392);
nor U2701 (N_2701,In_2072,In_113);
and U2702 (N_2702,In_2315,In_2016);
nand U2703 (N_2703,In_2101,In_2131);
and U2704 (N_2704,In_2260,In_2378);
or U2705 (N_2705,In_2014,In_1852);
and U2706 (N_2706,In_994,In_113);
nor U2707 (N_2707,In_1258,In_1130);
nor U2708 (N_2708,In_1329,In_762);
xnor U2709 (N_2709,In_538,In_397);
and U2710 (N_2710,In_1657,In_779);
nand U2711 (N_2711,In_1064,In_1464);
or U2712 (N_2712,In_1911,In_944);
nand U2713 (N_2713,In_1023,In_1897);
or U2714 (N_2714,In_2471,In_1165);
or U2715 (N_2715,In_2308,In_1691);
xor U2716 (N_2716,In_2036,In_1358);
or U2717 (N_2717,In_2275,In_265);
nor U2718 (N_2718,In_585,In_760);
and U2719 (N_2719,In_316,In_847);
nand U2720 (N_2720,In_305,In_2165);
or U2721 (N_2721,In_247,In_422);
nand U2722 (N_2722,In_1752,In_1093);
xor U2723 (N_2723,In_2253,In_51);
and U2724 (N_2724,In_1106,In_1809);
or U2725 (N_2725,In_1171,In_2146);
xor U2726 (N_2726,In_501,In_665);
and U2727 (N_2727,In_1295,In_1901);
xor U2728 (N_2728,In_356,In_253);
nor U2729 (N_2729,In_248,In_2498);
xnor U2730 (N_2730,In_861,In_188);
xor U2731 (N_2731,In_1238,In_2003);
and U2732 (N_2732,In_9,In_1758);
and U2733 (N_2733,In_1035,In_1807);
nand U2734 (N_2734,In_146,In_2449);
and U2735 (N_2735,In_1273,In_1736);
and U2736 (N_2736,In_989,In_1578);
xnor U2737 (N_2737,In_1206,In_1294);
xor U2738 (N_2738,In_2437,In_1880);
xnor U2739 (N_2739,In_504,In_1497);
or U2740 (N_2740,In_1910,In_333);
nor U2741 (N_2741,In_1776,In_2211);
and U2742 (N_2742,In_473,In_2303);
or U2743 (N_2743,In_380,In_2279);
or U2744 (N_2744,In_118,In_2032);
xnor U2745 (N_2745,In_271,In_1416);
and U2746 (N_2746,In_1988,In_1092);
or U2747 (N_2747,In_736,In_339);
xnor U2748 (N_2748,In_1850,In_1616);
or U2749 (N_2749,In_1916,In_766);
xor U2750 (N_2750,In_606,In_1731);
nor U2751 (N_2751,In_1745,In_2392);
nor U2752 (N_2752,In_2164,In_650);
and U2753 (N_2753,In_282,In_93);
and U2754 (N_2754,In_738,In_1135);
and U2755 (N_2755,In_753,In_996);
and U2756 (N_2756,In_953,In_183);
nor U2757 (N_2757,In_188,In_566);
nor U2758 (N_2758,In_97,In_1126);
xnor U2759 (N_2759,In_123,In_1166);
nor U2760 (N_2760,In_1041,In_2006);
nand U2761 (N_2761,In_1668,In_2375);
nand U2762 (N_2762,In_1852,In_968);
or U2763 (N_2763,In_1723,In_1493);
nor U2764 (N_2764,In_15,In_1915);
nand U2765 (N_2765,In_2362,In_370);
nor U2766 (N_2766,In_932,In_1019);
xor U2767 (N_2767,In_133,In_2233);
or U2768 (N_2768,In_672,In_2118);
xor U2769 (N_2769,In_2357,In_1428);
or U2770 (N_2770,In_402,In_1837);
and U2771 (N_2771,In_1889,In_739);
nor U2772 (N_2772,In_666,In_1502);
xor U2773 (N_2773,In_2223,In_11);
or U2774 (N_2774,In_222,In_1273);
nand U2775 (N_2775,In_2403,In_2118);
and U2776 (N_2776,In_1074,In_2098);
or U2777 (N_2777,In_583,In_1704);
or U2778 (N_2778,In_114,In_1069);
xnor U2779 (N_2779,In_143,In_458);
nand U2780 (N_2780,In_2059,In_690);
xor U2781 (N_2781,In_2269,In_381);
and U2782 (N_2782,In_970,In_1836);
xor U2783 (N_2783,In_1386,In_534);
nor U2784 (N_2784,In_1093,In_1254);
and U2785 (N_2785,In_408,In_523);
nand U2786 (N_2786,In_1740,In_1878);
nand U2787 (N_2787,In_56,In_2434);
nor U2788 (N_2788,In_172,In_1664);
nand U2789 (N_2789,In_1201,In_245);
or U2790 (N_2790,In_2148,In_709);
xnor U2791 (N_2791,In_1854,In_2082);
nand U2792 (N_2792,In_545,In_799);
nand U2793 (N_2793,In_1572,In_1393);
nor U2794 (N_2794,In_246,In_1196);
and U2795 (N_2795,In_762,In_1183);
and U2796 (N_2796,In_843,In_1603);
nand U2797 (N_2797,In_1125,In_369);
or U2798 (N_2798,In_2282,In_1987);
xor U2799 (N_2799,In_330,In_1999);
and U2800 (N_2800,In_2193,In_68);
nand U2801 (N_2801,In_898,In_1533);
and U2802 (N_2802,In_311,In_1470);
and U2803 (N_2803,In_716,In_363);
xor U2804 (N_2804,In_890,In_1386);
xnor U2805 (N_2805,In_1233,In_2479);
and U2806 (N_2806,In_2238,In_2159);
nand U2807 (N_2807,In_1252,In_1313);
nor U2808 (N_2808,In_1852,In_83);
nand U2809 (N_2809,In_1041,In_2259);
and U2810 (N_2810,In_1287,In_62);
or U2811 (N_2811,In_2166,In_1757);
nand U2812 (N_2812,In_55,In_1750);
and U2813 (N_2813,In_458,In_2066);
nand U2814 (N_2814,In_255,In_324);
or U2815 (N_2815,In_999,In_1150);
xnor U2816 (N_2816,In_1153,In_11);
nand U2817 (N_2817,In_2053,In_1419);
or U2818 (N_2818,In_563,In_1617);
nor U2819 (N_2819,In_538,In_109);
nand U2820 (N_2820,In_351,In_2266);
or U2821 (N_2821,In_1294,In_1585);
nand U2822 (N_2822,In_396,In_770);
xor U2823 (N_2823,In_1182,In_1797);
xnor U2824 (N_2824,In_841,In_2189);
nor U2825 (N_2825,In_2031,In_298);
or U2826 (N_2826,In_302,In_1745);
and U2827 (N_2827,In_260,In_1675);
nand U2828 (N_2828,In_1808,In_2207);
nand U2829 (N_2829,In_1211,In_2353);
nand U2830 (N_2830,In_1770,In_776);
nor U2831 (N_2831,In_1936,In_1602);
nand U2832 (N_2832,In_1672,In_503);
nor U2833 (N_2833,In_2141,In_2086);
nand U2834 (N_2834,In_2416,In_1235);
nor U2835 (N_2835,In_783,In_84);
and U2836 (N_2836,In_172,In_801);
xnor U2837 (N_2837,In_1579,In_2268);
xor U2838 (N_2838,In_756,In_762);
nand U2839 (N_2839,In_2312,In_1609);
or U2840 (N_2840,In_484,In_1290);
nand U2841 (N_2841,In_1064,In_2423);
nand U2842 (N_2842,In_2091,In_2473);
or U2843 (N_2843,In_1833,In_467);
nor U2844 (N_2844,In_1248,In_1805);
or U2845 (N_2845,In_1957,In_1954);
nor U2846 (N_2846,In_45,In_2318);
nand U2847 (N_2847,In_2012,In_1191);
xnor U2848 (N_2848,In_120,In_85);
and U2849 (N_2849,In_641,In_504);
nor U2850 (N_2850,In_2263,In_2236);
or U2851 (N_2851,In_801,In_1867);
and U2852 (N_2852,In_1318,In_2058);
and U2853 (N_2853,In_1601,In_1741);
nand U2854 (N_2854,In_813,In_2191);
xnor U2855 (N_2855,In_834,In_2492);
xor U2856 (N_2856,In_1650,In_319);
xor U2857 (N_2857,In_1223,In_655);
and U2858 (N_2858,In_2314,In_2057);
nor U2859 (N_2859,In_2268,In_292);
xor U2860 (N_2860,In_1898,In_550);
nor U2861 (N_2861,In_39,In_2382);
and U2862 (N_2862,In_1913,In_1033);
and U2863 (N_2863,In_2277,In_1021);
nor U2864 (N_2864,In_1152,In_2307);
xnor U2865 (N_2865,In_1354,In_351);
and U2866 (N_2866,In_608,In_208);
or U2867 (N_2867,In_1774,In_858);
and U2868 (N_2868,In_584,In_1929);
or U2869 (N_2869,In_2490,In_1628);
xor U2870 (N_2870,In_634,In_1004);
xnor U2871 (N_2871,In_1653,In_1503);
xnor U2872 (N_2872,In_2296,In_2490);
nor U2873 (N_2873,In_1617,In_1373);
and U2874 (N_2874,In_400,In_2484);
and U2875 (N_2875,In_1328,In_1752);
xor U2876 (N_2876,In_159,In_1228);
nor U2877 (N_2877,In_2499,In_2030);
or U2878 (N_2878,In_1218,In_2247);
or U2879 (N_2879,In_2398,In_1513);
xnor U2880 (N_2880,In_2345,In_408);
nand U2881 (N_2881,In_1048,In_989);
or U2882 (N_2882,In_1734,In_2266);
and U2883 (N_2883,In_1767,In_101);
and U2884 (N_2884,In_2498,In_1828);
or U2885 (N_2885,In_1305,In_167);
or U2886 (N_2886,In_2155,In_2322);
nand U2887 (N_2887,In_2120,In_2229);
xor U2888 (N_2888,In_1015,In_711);
and U2889 (N_2889,In_1838,In_1506);
and U2890 (N_2890,In_734,In_1779);
nand U2891 (N_2891,In_1596,In_123);
nand U2892 (N_2892,In_2233,In_2435);
or U2893 (N_2893,In_1805,In_548);
nor U2894 (N_2894,In_1389,In_1553);
and U2895 (N_2895,In_1359,In_1687);
nand U2896 (N_2896,In_2319,In_291);
xor U2897 (N_2897,In_1998,In_2412);
nor U2898 (N_2898,In_762,In_1423);
nand U2899 (N_2899,In_2444,In_790);
and U2900 (N_2900,In_2181,In_562);
and U2901 (N_2901,In_2453,In_1093);
nor U2902 (N_2902,In_278,In_1497);
nor U2903 (N_2903,In_312,In_265);
nor U2904 (N_2904,In_736,In_926);
and U2905 (N_2905,In_2446,In_1722);
and U2906 (N_2906,In_348,In_2243);
nand U2907 (N_2907,In_2266,In_1050);
nor U2908 (N_2908,In_884,In_1404);
nand U2909 (N_2909,In_2428,In_521);
nand U2910 (N_2910,In_1951,In_1136);
and U2911 (N_2911,In_1533,In_2341);
xor U2912 (N_2912,In_180,In_1813);
nand U2913 (N_2913,In_811,In_1151);
xnor U2914 (N_2914,In_1855,In_1403);
xor U2915 (N_2915,In_583,In_1008);
xor U2916 (N_2916,In_202,In_2007);
xor U2917 (N_2917,In_1800,In_603);
and U2918 (N_2918,In_1457,In_2047);
and U2919 (N_2919,In_725,In_1327);
nand U2920 (N_2920,In_476,In_1235);
nor U2921 (N_2921,In_2050,In_947);
and U2922 (N_2922,In_1021,In_873);
nor U2923 (N_2923,In_2146,In_1294);
xor U2924 (N_2924,In_900,In_2238);
nand U2925 (N_2925,In_43,In_1978);
nand U2926 (N_2926,In_1463,In_106);
xnor U2927 (N_2927,In_1388,In_1275);
nor U2928 (N_2928,In_614,In_1184);
nor U2929 (N_2929,In_1467,In_2332);
and U2930 (N_2930,In_1886,In_2398);
and U2931 (N_2931,In_257,In_2416);
and U2932 (N_2932,In_352,In_1293);
nand U2933 (N_2933,In_90,In_1538);
and U2934 (N_2934,In_1284,In_1357);
nand U2935 (N_2935,In_1257,In_1599);
nand U2936 (N_2936,In_1894,In_878);
and U2937 (N_2937,In_1649,In_313);
nor U2938 (N_2938,In_2487,In_2171);
nand U2939 (N_2939,In_798,In_324);
xor U2940 (N_2940,In_2176,In_388);
xnor U2941 (N_2941,In_208,In_2197);
nand U2942 (N_2942,In_544,In_1865);
and U2943 (N_2943,In_1148,In_1280);
xor U2944 (N_2944,In_396,In_422);
or U2945 (N_2945,In_1073,In_1637);
or U2946 (N_2946,In_295,In_1638);
or U2947 (N_2947,In_199,In_1350);
and U2948 (N_2948,In_1029,In_878);
nor U2949 (N_2949,In_1849,In_432);
xor U2950 (N_2950,In_2384,In_1279);
nor U2951 (N_2951,In_1264,In_439);
nand U2952 (N_2952,In_684,In_1276);
nand U2953 (N_2953,In_903,In_1582);
nor U2954 (N_2954,In_230,In_1534);
and U2955 (N_2955,In_1790,In_182);
or U2956 (N_2956,In_186,In_775);
or U2957 (N_2957,In_2464,In_2429);
nand U2958 (N_2958,In_1442,In_1429);
and U2959 (N_2959,In_834,In_356);
nand U2960 (N_2960,In_132,In_1214);
nand U2961 (N_2961,In_1291,In_1880);
and U2962 (N_2962,In_2438,In_582);
or U2963 (N_2963,In_1253,In_1002);
nor U2964 (N_2964,In_1214,In_1704);
or U2965 (N_2965,In_2022,In_47);
and U2966 (N_2966,In_697,In_2128);
or U2967 (N_2967,In_2441,In_287);
nand U2968 (N_2968,In_1698,In_261);
or U2969 (N_2969,In_1938,In_339);
nor U2970 (N_2970,In_2035,In_598);
nand U2971 (N_2971,In_257,In_1133);
and U2972 (N_2972,In_474,In_1991);
nor U2973 (N_2973,In_209,In_438);
and U2974 (N_2974,In_2463,In_1344);
or U2975 (N_2975,In_1099,In_87);
nor U2976 (N_2976,In_1683,In_144);
nor U2977 (N_2977,In_1323,In_1410);
nand U2978 (N_2978,In_1167,In_319);
xnor U2979 (N_2979,In_682,In_198);
nor U2980 (N_2980,In_1978,In_385);
nor U2981 (N_2981,In_945,In_1196);
and U2982 (N_2982,In_1368,In_180);
and U2983 (N_2983,In_346,In_50);
xor U2984 (N_2984,In_1259,In_272);
and U2985 (N_2985,In_1314,In_399);
or U2986 (N_2986,In_662,In_196);
nor U2987 (N_2987,In_508,In_1291);
or U2988 (N_2988,In_1174,In_2072);
and U2989 (N_2989,In_2091,In_127);
and U2990 (N_2990,In_1110,In_728);
xnor U2991 (N_2991,In_1711,In_802);
and U2992 (N_2992,In_600,In_1781);
and U2993 (N_2993,In_1539,In_846);
or U2994 (N_2994,In_2065,In_960);
and U2995 (N_2995,In_10,In_162);
and U2996 (N_2996,In_560,In_1637);
nor U2997 (N_2997,In_2357,In_954);
and U2998 (N_2998,In_2178,In_1123);
nand U2999 (N_2999,In_1271,In_1003);
nor U3000 (N_3000,In_2075,In_140);
or U3001 (N_3001,In_1263,In_2288);
or U3002 (N_3002,In_37,In_2473);
nand U3003 (N_3003,In_1623,In_1598);
xnor U3004 (N_3004,In_1902,In_1009);
and U3005 (N_3005,In_703,In_2136);
nand U3006 (N_3006,In_1627,In_1211);
nor U3007 (N_3007,In_1559,In_1117);
nor U3008 (N_3008,In_2366,In_635);
nand U3009 (N_3009,In_1371,In_776);
nand U3010 (N_3010,In_602,In_2305);
nand U3011 (N_3011,In_497,In_439);
nor U3012 (N_3012,In_858,In_35);
or U3013 (N_3013,In_1656,In_106);
nor U3014 (N_3014,In_1337,In_278);
nand U3015 (N_3015,In_125,In_253);
nand U3016 (N_3016,In_1560,In_170);
nand U3017 (N_3017,In_1109,In_1756);
or U3018 (N_3018,In_204,In_2240);
xnor U3019 (N_3019,In_164,In_2484);
nand U3020 (N_3020,In_26,In_912);
nor U3021 (N_3021,In_223,In_1767);
nor U3022 (N_3022,In_608,In_1372);
or U3023 (N_3023,In_948,In_2360);
nor U3024 (N_3024,In_938,In_642);
xnor U3025 (N_3025,In_128,In_865);
nand U3026 (N_3026,In_2416,In_658);
nor U3027 (N_3027,In_1229,In_1359);
nor U3028 (N_3028,In_1692,In_2201);
and U3029 (N_3029,In_186,In_1507);
or U3030 (N_3030,In_593,In_2006);
or U3031 (N_3031,In_688,In_2424);
xnor U3032 (N_3032,In_197,In_660);
or U3033 (N_3033,In_1196,In_624);
xnor U3034 (N_3034,In_388,In_133);
nand U3035 (N_3035,In_1820,In_2169);
or U3036 (N_3036,In_836,In_977);
nor U3037 (N_3037,In_746,In_650);
nand U3038 (N_3038,In_647,In_241);
xnor U3039 (N_3039,In_1654,In_34);
and U3040 (N_3040,In_525,In_1535);
nor U3041 (N_3041,In_1761,In_603);
or U3042 (N_3042,In_556,In_1530);
and U3043 (N_3043,In_555,In_1505);
xnor U3044 (N_3044,In_1200,In_1409);
xor U3045 (N_3045,In_753,In_1311);
xnor U3046 (N_3046,In_1451,In_1156);
and U3047 (N_3047,In_73,In_381);
or U3048 (N_3048,In_1058,In_964);
and U3049 (N_3049,In_1831,In_1297);
or U3050 (N_3050,In_492,In_2337);
or U3051 (N_3051,In_1008,In_970);
nor U3052 (N_3052,In_2298,In_1658);
or U3053 (N_3053,In_1244,In_440);
nor U3054 (N_3054,In_251,In_1997);
xor U3055 (N_3055,In_1007,In_1995);
xnor U3056 (N_3056,In_2475,In_1556);
and U3057 (N_3057,In_442,In_635);
and U3058 (N_3058,In_1113,In_455);
xnor U3059 (N_3059,In_1198,In_1813);
xnor U3060 (N_3060,In_2262,In_649);
nor U3061 (N_3061,In_1815,In_199);
nor U3062 (N_3062,In_1619,In_2095);
or U3063 (N_3063,In_2005,In_1322);
nor U3064 (N_3064,In_2109,In_1135);
and U3065 (N_3065,In_823,In_64);
and U3066 (N_3066,In_1134,In_2419);
nand U3067 (N_3067,In_1328,In_2367);
xnor U3068 (N_3068,In_729,In_584);
nor U3069 (N_3069,In_447,In_1277);
xor U3070 (N_3070,In_897,In_1436);
xor U3071 (N_3071,In_2469,In_559);
and U3072 (N_3072,In_2390,In_1151);
xor U3073 (N_3073,In_35,In_302);
nor U3074 (N_3074,In_2482,In_895);
nand U3075 (N_3075,In_519,In_673);
nor U3076 (N_3076,In_647,In_921);
or U3077 (N_3077,In_2076,In_886);
xnor U3078 (N_3078,In_465,In_2460);
and U3079 (N_3079,In_1885,In_2231);
and U3080 (N_3080,In_734,In_2333);
and U3081 (N_3081,In_1763,In_2479);
nor U3082 (N_3082,In_1589,In_2122);
and U3083 (N_3083,In_726,In_1835);
and U3084 (N_3084,In_2365,In_1580);
nor U3085 (N_3085,In_1950,In_905);
and U3086 (N_3086,In_1211,In_754);
nor U3087 (N_3087,In_1931,In_938);
or U3088 (N_3088,In_11,In_109);
or U3089 (N_3089,In_2355,In_626);
and U3090 (N_3090,In_479,In_1551);
or U3091 (N_3091,In_1555,In_609);
and U3092 (N_3092,In_1857,In_239);
or U3093 (N_3093,In_1996,In_1731);
nand U3094 (N_3094,In_844,In_1207);
or U3095 (N_3095,In_1804,In_2017);
xnor U3096 (N_3096,In_615,In_1238);
nand U3097 (N_3097,In_1876,In_1628);
nand U3098 (N_3098,In_69,In_796);
xnor U3099 (N_3099,In_733,In_2419);
nor U3100 (N_3100,In_1251,In_1465);
or U3101 (N_3101,In_2407,In_2170);
nand U3102 (N_3102,In_1888,In_940);
nand U3103 (N_3103,In_2348,In_581);
xor U3104 (N_3104,In_2367,In_1350);
nand U3105 (N_3105,In_1857,In_1570);
xor U3106 (N_3106,In_2063,In_1144);
and U3107 (N_3107,In_1017,In_1611);
or U3108 (N_3108,In_1171,In_298);
nor U3109 (N_3109,In_2447,In_910);
nor U3110 (N_3110,In_1621,In_1978);
nand U3111 (N_3111,In_1162,In_521);
xnor U3112 (N_3112,In_1642,In_2314);
xnor U3113 (N_3113,In_921,In_1753);
nand U3114 (N_3114,In_2199,In_868);
xor U3115 (N_3115,In_1971,In_2254);
nor U3116 (N_3116,In_847,In_2467);
and U3117 (N_3117,In_1027,In_1643);
xor U3118 (N_3118,In_1256,In_2475);
or U3119 (N_3119,In_72,In_1485);
and U3120 (N_3120,In_2157,In_28);
and U3121 (N_3121,In_1100,In_1695);
xnor U3122 (N_3122,In_1833,In_1147);
xor U3123 (N_3123,In_1887,In_1624);
xor U3124 (N_3124,In_401,In_827);
or U3125 (N_3125,In_2250,In_1498);
and U3126 (N_3126,In_1232,In_1599);
nor U3127 (N_3127,In_1444,In_2037);
nand U3128 (N_3128,In_2363,In_2213);
nor U3129 (N_3129,In_197,In_1188);
and U3130 (N_3130,In_511,In_942);
and U3131 (N_3131,In_2053,In_222);
nand U3132 (N_3132,In_1576,In_2156);
nor U3133 (N_3133,In_1347,In_1442);
xor U3134 (N_3134,In_253,In_71);
and U3135 (N_3135,In_915,In_521);
or U3136 (N_3136,In_2316,In_1456);
and U3137 (N_3137,In_524,In_2484);
nand U3138 (N_3138,In_533,In_142);
nor U3139 (N_3139,In_2462,In_617);
nor U3140 (N_3140,In_847,In_642);
nor U3141 (N_3141,In_881,In_1316);
xnor U3142 (N_3142,In_1952,In_511);
xor U3143 (N_3143,In_1520,In_1103);
xor U3144 (N_3144,In_603,In_2496);
nand U3145 (N_3145,In_1265,In_304);
or U3146 (N_3146,In_1247,In_745);
nand U3147 (N_3147,In_1373,In_1780);
nand U3148 (N_3148,In_2153,In_2054);
nor U3149 (N_3149,In_1693,In_1382);
or U3150 (N_3150,In_576,In_2472);
and U3151 (N_3151,In_1141,In_33);
and U3152 (N_3152,In_1649,In_934);
nand U3153 (N_3153,In_2217,In_1305);
nand U3154 (N_3154,In_1160,In_1937);
or U3155 (N_3155,In_76,In_42);
xnor U3156 (N_3156,In_1793,In_962);
nand U3157 (N_3157,In_856,In_211);
nor U3158 (N_3158,In_1091,In_1845);
nor U3159 (N_3159,In_471,In_1150);
xor U3160 (N_3160,In_77,In_1842);
nand U3161 (N_3161,In_2334,In_636);
and U3162 (N_3162,In_1884,In_285);
xor U3163 (N_3163,In_510,In_77);
nor U3164 (N_3164,In_773,In_1194);
and U3165 (N_3165,In_1092,In_1516);
nor U3166 (N_3166,In_1130,In_134);
and U3167 (N_3167,In_1706,In_702);
nand U3168 (N_3168,In_2344,In_474);
or U3169 (N_3169,In_450,In_715);
nor U3170 (N_3170,In_1945,In_1134);
or U3171 (N_3171,In_1894,In_2255);
or U3172 (N_3172,In_1381,In_1880);
nand U3173 (N_3173,In_457,In_1077);
or U3174 (N_3174,In_639,In_2147);
and U3175 (N_3175,In_2225,In_1295);
nand U3176 (N_3176,In_803,In_2290);
xor U3177 (N_3177,In_101,In_1714);
xor U3178 (N_3178,In_779,In_869);
xnor U3179 (N_3179,In_1688,In_153);
nor U3180 (N_3180,In_850,In_2145);
or U3181 (N_3181,In_76,In_25);
or U3182 (N_3182,In_504,In_2012);
and U3183 (N_3183,In_1336,In_1662);
xnor U3184 (N_3184,In_1355,In_1213);
or U3185 (N_3185,In_2260,In_1787);
or U3186 (N_3186,In_1691,In_429);
xor U3187 (N_3187,In_777,In_2021);
or U3188 (N_3188,In_1527,In_1125);
nor U3189 (N_3189,In_1852,In_2315);
xor U3190 (N_3190,In_2106,In_1744);
nor U3191 (N_3191,In_278,In_473);
and U3192 (N_3192,In_1592,In_1291);
or U3193 (N_3193,In_544,In_1673);
nor U3194 (N_3194,In_140,In_2031);
nand U3195 (N_3195,In_2283,In_1311);
nor U3196 (N_3196,In_174,In_638);
nand U3197 (N_3197,In_1328,In_1072);
nor U3198 (N_3198,In_1670,In_252);
nor U3199 (N_3199,In_1467,In_2247);
nand U3200 (N_3200,In_1975,In_2076);
xnor U3201 (N_3201,In_398,In_2294);
or U3202 (N_3202,In_2327,In_597);
nand U3203 (N_3203,In_1839,In_1349);
nand U3204 (N_3204,In_1126,In_409);
xor U3205 (N_3205,In_114,In_2132);
xnor U3206 (N_3206,In_703,In_1639);
or U3207 (N_3207,In_1652,In_1939);
xor U3208 (N_3208,In_704,In_1181);
xor U3209 (N_3209,In_1273,In_2018);
or U3210 (N_3210,In_2395,In_2312);
or U3211 (N_3211,In_1055,In_1057);
nor U3212 (N_3212,In_1980,In_962);
nor U3213 (N_3213,In_1880,In_1247);
and U3214 (N_3214,In_1704,In_1517);
and U3215 (N_3215,In_2295,In_1419);
nor U3216 (N_3216,In_2048,In_250);
xor U3217 (N_3217,In_672,In_1340);
nand U3218 (N_3218,In_2298,In_1103);
xnor U3219 (N_3219,In_173,In_2411);
xnor U3220 (N_3220,In_645,In_1384);
xnor U3221 (N_3221,In_2153,In_1070);
xor U3222 (N_3222,In_1210,In_1342);
and U3223 (N_3223,In_600,In_1113);
nor U3224 (N_3224,In_634,In_1095);
nor U3225 (N_3225,In_732,In_1331);
and U3226 (N_3226,In_2424,In_1613);
nand U3227 (N_3227,In_1768,In_2286);
nor U3228 (N_3228,In_773,In_1812);
nand U3229 (N_3229,In_794,In_72);
or U3230 (N_3230,In_1516,In_409);
nand U3231 (N_3231,In_58,In_1019);
and U3232 (N_3232,In_1344,In_948);
nand U3233 (N_3233,In_1531,In_1066);
nor U3234 (N_3234,In_317,In_221);
or U3235 (N_3235,In_1999,In_2482);
and U3236 (N_3236,In_1706,In_2211);
nand U3237 (N_3237,In_1613,In_369);
nor U3238 (N_3238,In_1622,In_901);
nor U3239 (N_3239,In_2377,In_896);
xor U3240 (N_3240,In_2213,In_2408);
xnor U3241 (N_3241,In_2164,In_252);
and U3242 (N_3242,In_2258,In_1324);
and U3243 (N_3243,In_1300,In_632);
or U3244 (N_3244,In_2217,In_2333);
and U3245 (N_3245,In_593,In_2479);
nor U3246 (N_3246,In_864,In_1839);
and U3247 (N_3247,In_658,In_1100);
and U3248 (N_3248,In_1354,In_2478);
or U3249 (N_3249,In_2221,In_1928);
xor U3250 (N_3250,In_936,In_9);
or U3251 (N_3251,In_1094,In_251);
and U3252 (N_3252,In_758,In_2048);
nor U3253 (N_3253,In_1212,In_870);
and U3254 (N_3254,In_1760,In_2443);
and U3255 (N_3255,In_1556,In_1937);
xor U3256 (N_3256,In_782,In_1585);
and U3257 (N_3257,In_809,In_2318);
or U3258 (N_3258,In_2110,In_1712);
nor U3259 (N_3259,In_1653,In_864);
and U3260 (N_3260,In_1529,In_25);
nor U3261 (N_3261,In_1498,In_1064);
xnor U3262 (N_3262,In_760,In_2055);
and U3263 (N_3263,In_650,In_747);
xor U3264 (N_3264,In_1531,In_1546);
nand U3265 (N_3265,In_52,In_1408);
or U3266 (N_3266,In_768,In_1603);
xnor U3267 (N_3267,In_1590,In_2108);
xor U3268 (N_3268,In_1851,In_506);
nand U3269 (N_3269,In_1804,In_987);
nand U3270 (N_3270,In_725,In_362);
xnor U3271 (N_3271,In_2081,In_321);
nand U3272 (N_3272,In_2238,In_263);
and U3273 (N_3273,In_1458,In_1023);
nor U3274 (N_3274,In_1877,In_1290);
nor U3275 (N_3275,In_134,In_1168);
or U3276 (N_3276,In_956,In_2473);
or U3277 (N_3277,In_1505,In_902);
nand U3278 (N_3278,In_1908,In_2385);
nor U3279 (N_3279,In_398,In_57);
xor U3280 (N_3280,In_457,In_146);
nor U3281 (N_3281,In_763,In_1406);
nor U3282 (N_3282,In_1698,In_2190);
nand U3283 (N_3283,In_1873,In_1366);
and U3284 (N_3284,In_1050,In_904);
nand U3285 (N_3285,In_687,In_1765);
nor U3286 (N_3286,In_1543,In_1411);
nand U3287 (N_3287,In_1631,In_88);
nor U3288 (N_3288,In_1288,In_2136);
and U3289 (N_3289,In_2168,In_872);
or U3290 (N_3290,In_218,In_2081);
or U3291 (N_3291,In_1042,In_30);
nor U3292 (N_3292,In_820,In_65);
xnor U3293 (N_3293,In_2466,In_1510);
xnor U3294 (N_3294,In_408,In_728);
nor U3295 (N_3295,In_510,In_2400);
or U3296 (N_3296,In_955,In_1427);
or U3297 (N_3297,In_1937,In_909);
and U3298 (N_3298,In_1781,In_2131);
or U3299 (N_3299,In_2132,In_387);
nor U3300 (N_3300,In_1144,In_1435);
or U3301 (N_3301,In_1341,In_1257);
xnor U3302 (N_3302,In_2116,In_354);
nand U3303 (N_3303,In_1600,In_1996);
xor U3304 (N_3304,In_1335,In_894);
nor U3305 (N_3305,In_2408,In_495);
xor U3306 (N_3306,In_1512,In_1770);
and U3307 (N_3307,In_109,In_2182);
or U3308 (N_3308,In_228,In_997);
or U3309 (N_3309,In_1424,In_99);
nor U3310 (N_3310,In_2292,In_1070);
and U3311 (N_3311,In_2236,In_681);
nand U3312 (N_3312,In_1018,In_586);
or U3313 (N_3313,In_1479,In_577);
nor U3314 (N_3314,In_1881,In_791);
nand U3315 (N_3315,In_1697,In_19);
nand U3316 (N_3316,In_128,In_2286);
or U3317 (N_3317,In_2405,In_2432);
nand U3318 (N_3318,In_2164,In_2075);
nand U3319 (N_3319,In_528,In_1772);
and U3320 (N_3320,In_411,In_2058);
xnor U3321 (N_3321,In_485,In_1903);
or U3322 (N_3322,In_677,In_1950);
nor U3323 (N_3323,In_1213,In_788);
or U3324 (N_3324,In_166,In_1714);
nor U3325 (N_3325,In_2278,In_507);
and U3326 (N_3326,In_1969,In_753);
and U3327 (N_3327,In_699,In_1803);
xnor U3328 (N_3328,In_411,In_395);
xor U3329 (N_3329,In_810,In_2002);
nor U3330 (N_3330,In_1025,In_1338);
nand U3331 (N_3331,In_2172,In_2160);
and U3332 (N_3332,In_265,In_142);
and U3333 (N_3333,In_237,In_2365);
and U3334 (N_3334,In_1811,In_816);
nand U3335 (N_3335,In_368,In_1362);
and U3336 (N_3336,In_2239,In_1512);
nand U3337 (N_3337,In_973,In_2473);
nand U3338 (N_3338,In_1668,In_25);
xnor U3339 (N_3339,In_1190,In_2273);
nand U3340 (N_3340,In_1680,In_687);
and U3341 (N_3341,In_875,In_1822);
nand U3342 (N_3342,In_648,In_1052);
nand U3343 (N_3343,In_305,In_2426);
or U3344 (N_3344,In_326,In_762);
or U3345 (N_3345,In_667,In_1372);
nand U3346 (N_3346,In_1435,In_1933);
nor U3347 (N_3347,In_1258,In_2189);
and U3348 (N_3348,In_2266,In_804);
nand U3349 (N_3349,In_115,In_1155);
nor U3350 (N_3350,In_1202,In_1912);
or U3351 (N_3351,In_288,In_2458);
and U3352 (N_3352,In_2324,In_2494);
nor U3353 (N_3353,In_1998,In_1473);
or U3354 (N_3354,In_1297,In_1303);
or U3355 (N_3355,In_1827,In_1367);
nand U3356 (N_3356,In_332,In_1178);
nand U3357 (N_3357,In_1442,In_1315);
or U3358 (N_3358,In_2044,In_1155);
or U3359 (N_3359,In_778,In_1721);
or U3360 (N_3360,In_2287,In_1828);
or U3361 (N_3361,In_278,In_405);
nand U3362 (N_3362,In_1185,In_768);
and U3363 (N_3363,In_1335,In_233);
xnor U3364 (N_3364,In_164,In_16);
xor U3365 (N_3365,In_1174,In_202);
or U3366 (N_3366,In_475,In_1556);
or U3367 (N_3367,In_1755,In_1401);
and U3368 (N_3368,In_279,In_2193);
and U3369 (N_3369,In_748,In_1849);
or U3370 (N_3370,In_993,In_1598);
nor U3371 (N_3371,In_509,In_2488);
nor U3372 (N_3372,In_64,In_836);
nor U3373 (N_3373,In_1975,In_731);
xor U3374 (N_3374,In_2482,In_257);
nand U3375 (N_3375,In_1851,In_1885);
nor U3376 (N_3376,In_473,In_2114);
nand U3377 (N_3377,In_1763,In_604);
nand U3378 (N_3378,In_645,In_2253);
nor U3379 (N_3379,In_2404,In_684);
xor U3380 (N_3380,In_1797,In_1476);
nor U3381 (N_3381,In_93,In_889);
nand U3382 (N_3382,In_2256,In_141);
nor U3383 (N_3383,In_1186,In_2410);
nand U3384 (N_3384,In_1593,In_2313);
or U3385 (N_3385,In_659,In_8);
or U3386 (N_3386,In_2323,In_692);
or U3387 (N_3387,In_700,In_1422);
xnor U3388 (N_3388,In_728,In_589);
nand U3389 (N_3389,In_512,In_2252);
nor U3390 (N_3390,In_334,In_83);
nand U3391 (N_3391,In_1443,In_170);
and U3392 (N_3392,In_2455,In_2413);
nor U3393 (N_3393,In_1582,In_1554);
and U3394 (N_3394,In_1155,In_1070);
and U3395 (N_3395,In_1939,In_1625);
or U3396 (N_3396,In_1109,In_324);
or U3397 (N_3397,In_391,In_704);
nand U3398 (N_3398,In_1416,In_827);
nor U3399 (N_3399,In_136,In_1121);
xor U3400 (N_3400,In_1751,In_525);
xor U3401 (N_3401,In_462,In_1164);
nor U3402 (N_3402,In_1784,In_2299);
or U3403 (N_3403,In_2000,In_1437);
nor U3404 (N_3404,In_557,In_1467);
nor U3405 (N_3405,In_587,In_2311);
xor U3406 (N_3406,In_276,In_1394);
nand U3407 (N_3407,In_2358,In_1855);
nand U3408 (N_3408,In_550,In_1817);
xnor U3409 (N_3409,In_67,In_1066);
nor U3410 (N_3410,In_62,In_1231);
or U3411 (N_3411,In_2448,In_163);
or U3412 (N_3412,In_1013,In_595);
xor U3413 (N_3413,In_2263,In_2104);
nand U3414 (N_3414,In_284,In_2170);
xnor U3415 (N_3415,In_1154,In_915);
xnor U3416 (N_3416,In_568,In_2228);
nand U3417 (N_3417,In_960,In_1113);
or U3418 (N_3418,In_375,In_1226);
or U3419 (N_3419,In_2043,In_735);
xnor U3420 (N_3420,In_928,In_2225);
nor U3421 (N_3421,In_1254,In_1765);
nand U3422 (N_3422,In_160,In_1566);
nand U3423 (N_3423,In_495,In_1001);
nand U3424 (N_3424,In_1827,In_127);
nand U3425 (N_3425,In_2304,In_599);
and U3426 (N_3426,In_620,In_10);
nor U3427 (N_3427,In_91,In_2059);
nand U3428 (N_3428,In_1607,In_1856);
or U3429 (N_3429,In_2166,In_454);
nor U3430 (N_3430,In_894,In_593);
xor U3431 (N_3431,In_70,In_1500);
nor U3432 (N_3432,In_2351,In_2412);
nor U3433 (N_3433,In_331,In_1875);
xor U3434 (N_3434,In_1022,In_345);
xor U3435 (N_3435,In_239,In_1944);
nand U3436 (N_3436,In_2124,In_940);
and U3437 (N_3437,In_1256,In_560);
and U3438 (N_3438,In_638,In_1061);
nand U3439 (N_3439,In_947,In_57);
xor U3440 (N_3440,In_830,In_1210);
and U3441 (N_3441,In_1336,In_299);
xnor U3442 (N_3442,In_894,In_35);
or U3443 (N_3443,In_947,In_2267);
xor U3444 (N_3444,In_65,In_1039);
nor U3445 (N_3445,In_795,In_1710);
nand U3446 (N_3446,In_1845,In_1954);
xnor U3447 (N_3447,In_2308,In_371);
and U3448 (N_3448,In_80,In_1077);
xor U3449 (N_3449,In_699,In_1701);
xnor U3450 (N_3450,In_1303,In_1708);
or U3451 (N_3451,In_1595,In_2419);
or U3452 (N_3452,In_1688,In_202);
nand U3453 (N_3453,In_1671,In_429);
nor U3454 (N_3454,In_1270,In_2127);
xor U3455 (N_3455,In_597,In_1028);
and U3456 (N_3456,In_169,In_756);
nor U3457 (N_3457,In_2320,In_1712);
and U3458 (N_3458,In_874,In_1711);
nand U3459 (N_3459,In_149,In_164);
nor U3460 (N_3460,In_913,In_769);
xor U3461 (N_3461,In_1115,In_228);
or U3462 (N_3462,In_712,In_597);
and U3463 (N_3463,In_2234,In_2485);
xnor U3464 (N_3464,In_1209,In_1085);
nor U3465 (N_3465,In_742,In_2437);
nor U3466 (N_3466,In_2431,In_272);
and U3467 (N_3467,In_2344,In_697);
nor U3468 (N_3468,In_146,In_2435);
nand U3469 (N_3469,In_833,In_2033);
or U3470 (N_3470,In_463,In_302);
or U3471 (N_3471,In_591,In_2092);
nand U3472 (N_3472,In_2387,In_1330);
nand U3473 (N_3473,In_416,In_165);
or U3474 (N_3474,In_1960,In_2430);
or U3475 (N_3475,In_2016,In_548);
or U3476 (N_3476,In_300,In_495);
and U3477 (N_3477,In_2292,In_89);
nor U3478 (N_3478,In_2338,In_2006);
or U3479 (N_3479,In_1255,In_1758);
xor U3480 (N_3480,In_844,In_1819);
nand U3481 (N_3481,In_1617,In_7);
nand U3482 (N_3482,In_1067,In_1889);
nand U3483 (N_3483,In_62,In_1904);
nor U3484 (N_3484,In_1,In_1635);
xnor U3485 (N_3485,In_2443,In_1295);
or U3486 (N_3486,In_580,In_2185);
xor U3487 (N_3487,In_558,In_2156);
and U3488 (N_3488,In_2174,In_1550);
and U3489 (N_3489,In_1691,In_1707);
xnor U3490 (N_3490,In_1452,In_1505);
nor U3491 (N_3491,In_2484,In_1129);
or U3492 (N_3492,In_564,In_2005);
xor U3493 (N_3493,In_1863,In_1013);
and U3494 (N_3494,In_2487,In_1055);
and U3495 (N_3495,In_1260,In_1290);
or U3496 (N_3496,In_177,In_500);
and U3497 (N_3497,In_1930,In_1446);
xnor U3498 (N_3498,In_1938,In_1803);
nor U3499 (N_3499,In_1790,In_1286);
and U3500 (N_3500,In_384,In_1621);
or U3501 (N_3501,In_154,In_1988);
or U3502 (N_3502,In_814,In_484);
nor U3503 (N_3503,In_1648,In_2085);
and U3504 (N_3504,In_2310,In_1777);
nor U3505 (N_3505,In_1404,In_578);
nand U3506 (N_3506,In_203,In_2053);
or U3507 (N_3507,In_862,In_1647);
nand U3508 (N_3508,In_1568,In_2426);
nor U3509 (N_3509,In_1209,In_2437);
nor U3510 (N_3510,In_1497,In_828);
xnor U3511 (N_3511,In_1159,In_1446);
and U3512 (N_3512,In_377,In_1709);
or U3513 (N_3513,In_1898,In_686);
xor U3514 (N_3514,In_2303,In_1355);
and U3515 (N_3515,In_2001,In_1256);
xor U3516 (N_3516,In_379,In_2188);
xnor U3517 (N_3517,In_552,In_255);
xnor U3518 (N_3518,In_85,In_2422);
nand U3519 (N_3519,In_800,In_1985);
xnor U3520 (N_3520,In_913,In_680);
xnor U3521 (N_3521,In_19,In_2368);
nor U3522 (N_3522,In_2100,In_1801);
xnor U3523 (N_3523,In_1067,In_157);
xor U3524 (N_3524,In_919,In_2089);
xor U3525 (N_3525,In_113,In_333);
nand U3526 (N_3526,In_422,In_839);
xnor U3527 (N_3527,In_1140,In_336);
nand U3528 (N_3528,In_1124,In_374);
nand U3529 (N_3529,In_279,In_1020);
nand U3530 (N_3530,In_1305,In_302);
nand U3531 (N_3531,In_2205,In_208);
or U3532 (N_3532,In_950,In_1533);
xor U3533 (N_3533,In_907,In_1509);
or U3534 (N_3534,In_1692,In_1201);
nand U3535 (N_3535,In_2189,In_681);
xor U3536 (N_3536,In_870,In_1411);
nor U3537 (N_3537,In_204,In_1171);
nor U3538 (N_3538,In_1253,In_1360);
nand U3539 (N_3539,In_1052,In_1552);
nand U3540 (N_3540,In_949,In_2365);
nor U3541 (N_3541,In_354,In_397);
xnor U3542 (N_3542,In_1336,In_1847);
and U3543 (N_3543,In_1174,In_818);
nand U3544 (N_3544,In_512,In_1952);
or U3545 (N_3545,In_90,In_411);
nand U3546 (N_3546,In_1331,In_254);
nor U3547 (N_3547,In_1550,In_409);
nor U3548 (N_3548,In_834,In_2045);
or U3549 (N_3549,In_824,In_2287);
and U3550 (N_3550,In_1159,In_1370);
nor U3551 (N_3551,In_259,In_151);
xnor U3552 (N_3552,In_1402,In_1773);
or U3553 (N_3553,In_1840,In_312);
xnor U3554 (N_3554,In_1073,In_1409);
nor U3555 (N_3555,In_461,In_688);
xnor U3556 (N_3556,In_460,In_1233);
and U3557 (N_3557,In_758,In_1932);
and U3558 (N_3558,In_1273,In_333);
nor U3559 (N_3559,In_1474,In_2362);
and U3560 (N_3560,In_910,In_2337);
nand U3561 (N_3561,In_1699,In_1875);
nor U3562 (N_3562,In_672,In_1139);
nor U3563 (N_3563,In_1503,In_1152);
or U3564 (N_3564,In_574,In_378);
nand U3565 (N_3565,In_873,In_2299);
nand U3566 (N_3566,In_2021,In_1486);
nand U3567 (N_3567,In_185,In_1971);
xor U3568 (N_3568,In_2128,In_67);
xnor U3569 (N_3569,In_261,In_608);
and U3570 (N_3570,In_263,In_615);
xnor U3571 (N_3571,In_1339,In_2352);
nand U3572 (N_3572,In_147,In_509);
nand U3573 (N_3573,In_465,In_810);
or U3574 (N_3574,In_629,In_556);
or U3575 (N_3575,In_1894,In_800);
and U3576 (N_3576,In_510,In_1346);
xor U3577 (N_3577,In_1171,In_614);
and U3578 (N_3578,In_1305,In_1150);
and U3579 (N_3579,In_2315,In_882);
nand U3580 (N_3580,In_534,In_150);
or U3581 (N_3581,In_2474,In_2316);
nor U3582 (N_3582,In_46,In_475);
nor U3583 (N_3583,In_1367,In_2164);
and U3584 (N_3584,In_211,In_1803);
nand U3585 (N_3585,In_476,In_495);
and U3586 (N_3586,In_343,In_2341);
nor U3587 (N_3587,In_2058,In_1442);
or U3588 (N_3588,In_218,In_2418);
nand U3589 (N_3589,In_93,In_1300);
or U3590 (N_3590,In_138,In_1985);
nor U3591 (N_3591,In_307,In_139);
or U3592 (N_3592,In_2237,In_1218);
nand U3593 (N_3593,In_1633,In_1697);
xnor U3594 (N_3594,In_1917,In_83);
and U3595 (N_3595,In_1790,In_2380);
or U3596 (N_3596,In_1690,In_1972);
and U3597 (N_3597,In_442,In_1161);
and U3598 (N_3598,In_1084,In_915);
or U3599 (N_3599,In_843,In_207);
nand U3600 (N_3600,In_1400,In_1965);
and U3601 (N_3601,In_1867,In_996);
xnor U3602 (N_3602,In_1941,In_492);
and U3603 (N_3603,In_1743,In_37);
xor U3604 (N_3604,In_261,In_2204);
and U3605 (N_3605,In_225,In_1810);
xor U3606 (N_3606,In_1096,In_1093);
and U3607 (N_3607,In_815,In_839);
or U3608 (N_3608,In_2454,In_2319);
nand U3609 (N_3609,In_2178,In_1177);
xnor U3610 (N_3610,In_1251,In_623);
nor U3611 (N_3611,In_1207,In_1308);
nand U3612 (N_3612,In_1881,In_639);
or U3613 (N_3613,In_879,In_695);
or U3614 (N_3614,In_369,In_1531);
nand U3615 (N_3615,In_2217,In_2492);
xnor U3616 (N_3616,In_146,In_971);
and U3617 (N_3617,In_1121,In_114);
nand U3618 (N_3618,In_1354,In_1957);
nand U3619 (N_3619,In_1778,In_428);
nand U3620 (N_3620,In_407,In_726);
or U3621 (N_3621,In_2087,In_818);
xor U3622 (N_3622,In_1325,In_1161);
or U3623 (N_3623,In_1701,In_2132);
nand U3624 (N_3624,In_136,In_157);
xnor U3625 (N_3625,In_1459,In_1487);
or U3626 (N_3626,In_157,In_273);
and U3627 (N_3627,In_2162,In_128);
xnor U3628 (N_3628,In_1501,In_1585);
nor U3629 (N_3629,In_418,In_1077);
nand U3630 (N_3630,In_513,In_666);
nand U3631 (N_3631,In_816,In_470);
xnor U3632 (N_3632,In_8,In_704);
nand U3633 (N_3633,In_2431,In_848);
nor U3634 (N_3634,In_1759,In_86);
xnor U3635 (N_3635,In_1248,In_2101);
or U3636 (N_3636,In_396,In_496);
or U3637 (N_3637,In_1479,In_1828);
nor U3638 (N_3638,In_2192,In_545);
or U3639 (N_3639,In_485,In_1090);
or U3640 (N_3640,In_602,In_2267);
or U3641 (N_3641,In_2242,In_1282);
or U3642 (N_3642,In_1980,In_1891);
xnor U3643 (N_3643,In_1014,In_2387);
and U3644 (N_3644,In_1430,In_430);
or U3645 (N_3645,In_1744,In_1935);
or U3646 (N_3646,In_979,In_2116);
or U3647 (N_3647,In_2461,In_1639);
and U3648 (N_3648,In_82,In_2336);
xnor U3649 (N_3649,In_1772,In_1614);
nand U3650 (N_3650,In_1302,In_280);
nand U3651 (N_3651,In_99,In_1608);
or U3652 (N_3652,In_2205,In_2272);
nand U3653 (N_3653,In_1578,In_1975);
nand U3654 (N_3654,In_961,In_340);
nor U3655 (N_3655,In_2271,In_1942);
nor U3656 (N_3656,In_1625,In_1437);
or U3657 (N_3657,In_1893,In_1940);
xnor U3658 (N_3658,In_1488,In_1199);
and U3659 (N_3659,In_280,In_2081);
and U3660 (N_3660,In_1387,In_1643);
nor U3661 (N_3661,In_48,In_619);
nand U3662 (N_3662,In_1190,In_1281);
and U3663 (N_3663,In_936,In_1420);
nor U3664 (N_3664,In_2300,In_902);
nor U3665 (N_3665,In_375,In_510);
xor U3666 (N_3666,In_2177,In_390);
xor U3667 (N_3667,In_317,In_1543);
nand U3668 (N_3668,In_1836,In_2345);
or U3669 (N_3669,In_1634,In_171);
xor U3670 (N_3670,In_1716,In_625);
nor U3671 (N_3671,In_1930,In_175);
nor U3672 (N_3672,In_2064,In_1650);
nor U3673 (N_3673,In_2240,In_1576);
nand U3674 (N_3674,In_214,In_1773);
nand U3675 (N_3675,In_2468,In_1374);
or U3676 (N_3676,In_536,In_1247);
nor U3677 (N_3677,In_1168,In_1629);
xnor U3678 (N_3678,In_1902,In_1186);
xor U3679 (N_3679,In_2047,In_827);
nor U3680 (N_3680,In_1244,In_637);
or U3681 (N_3681,In_2093,In_630);
nand U3682 (N_3682,In_971,In_1737);
nor U3683 (N_3683,In_1726,In_2360);
and U3684 (N_3684,In_2473,In_2440);
and U3685 (N_3685,In_12,In_1140);
nand U3686 (N_3686,In_298,In_423);
or U3687 (N_3687,In_934,In_18);
and U3688 (N_3688,In_1516,In_1310);
xor U3689 (N_3689,In_715,In_2428);
nor U3690 (N_3690,In_594,In_1010);
nor U3691 (N_3691,In_778,In_2216);
or U3692 (N_3692,In_1375,In_1227);
xor U3693 (N_3693,In_1287,In_2182);
xor U3694 (N_3694,In_875,In_2282);
nand U3695 (N_3695,In_147,In_724);
xnor U3696 (N_3696,In_2238,In_1269);
nor U3697 (N_3697,In_789,In_62);
xnor U3698 (N_3698,In_2282,In_308);
nand U3699 (N_3699,In_60,In_446);
xnor U3700 (N_3700,In_297,In_2255);
and U3701 (N_3701,In_2114,In_2489);
or U3702 (N_3702,In_239,In_140);
or U3703 (N_3703,In_938,In_2080);
nand U3704 (N_3704,In_1116,In_787);
xor U3705 (N_3705,In_1340,In_2243);
xor U3706 (N_3706,In_2014,In_1950);
nor U3707 (N_3707,In_625,In_1320);
and U3708 (N_3708,In_284,In_1071);
nand U3709 (N_3709,In_1279,In_417);
nor U3710 (N_3710,In_2415,In_1171);
nor U3711 (N_3711,In_402,In_2384);
nand U3712 (N_3712,In_500,In_636);
or U3713 (N_3713,In_478,In_761);
nand U3714 (N_3714,In_2261,In_2429);
or U3715 (N_3715,In_1353,In_1813);
and U3716 (N_3716,In_840,In_1882);
and U3717 (N_3717,In_2452,In_1586);
or U3718 (N_3718,In_564,In_1883);
or U3719 (N_3719,In_1403,In_1545);
and U3720 (N_3720,In_1054,In_541);
and U3721 (N_3721,In_2011,In_599);
xor U3722 (N_3722,In_328,In_2445);
nor U3723 (N_3723,In_2461,In_1151);
and U3724 (N_3724,In_159,In_1146);
nor U3725 (N_3725,In_301,In_2012);
nor U3726 (N_3726,In_474,In_2055);
and U3727 (N_3727,In_2348,In_1416);
nor U3728 (N_3728,In_167,In_694);
nor U3729 (N_3729,In_720,In_773);
nand U3730 (N_3730,In_920,In_613);
nand U3731 (N_3731,In_1465,In_1680);
xor U3732 (N_3732,In_1477,In_1623);
xor U3733 (N_3733,In_843,In_1709);
nand U3734 (N_3734,In_2144,In_1480);
nor U3735 (N_3735,In_655,In_801);
xnor U3736 (N_3736,In_1038,In_905);
or U3737 (N_3737,In_719,In_871);
or U3738 (N_3738,In_2070,In_1639);
nand U3739 (N_3739,In_1466,In_494);
or U3740 (N_3740,In_1217,In_1058);
nand U3741 (N_3741,In_1373,In_1967);
xnor U3742 (N_3742,In_1107,In_743);
nand U3743 (N_3743,In_1979,In_2104);
nor U3744 (N_3744,In_2084,In_2);
nor U3745 (N_3745,In_1928,In_2020);
nand U3746 (N_3746,In_2332,In_2452);
xor U3747 (N_3747,In_2436,In_2479);
nor U3748 (N_3748,In_248,In_1909);
and U3749 (N_3749,In_338,In_1280);
xnor U3750 (N_3750,In_1828,In_1552);
xor U3751 (N_3751,In_1981,In_500);
and U3752 (N_3752,In_1859,In_2149);
nor U3753 (N_3753,In_1223,In_1674);
xor U3754 (N_3754,In_1674,In_778);
and U3755 (N_3755,In_837,In_1112);
nand U3756 (N_3756,In_844,In_1425);
and U3757 (N_3757,In_1341,In_1657);
or U3758 (N_3758,In_2120,In_2391);
or U3759 (N_3759,In_2013,In_1738);
and U3760 (N_3760,In_787,In_810);
xnor U3761 (N_3761,In_906,In_475);
or U3762 (N_3762,In_1043,In_0);
and U3763 (N_3763,In_1795,In_528);
and U3764 (N_3764,In_2193,In_1789);
xor U3765 (N_3765,In_614,In_38);
or U3766 (N_3766,In_2047,In_584);
nor U3767 (N_3767,In_1215,In_996);
xnor U3768 (N_3768,In_1904,In_251);
or U3769 (N_3769,In_1531,In_117);
nand U3770 (N_3770,In_2341,In_504);
nor U3771 (N_3771,In_1175,In_862);
nor U3772 (N_3772,In_965,In_1053);
xor U3773 (N_3773,In_1548,In_2152);
nor U3774 (N_3774,In_681,In_1848);
xor U3775 (N_3775,In_1582,In_1333);
nand U3776 (N_3776,In_60,In_1996);
nor U3777 (N_3777,In_1820,In_1495);
or U3778 (N_3778,In_1910,In_2493);
or U3779 (N_3779,In_404,In_2312);
nand U3780 (N_3780,In_70,In_1317);
nor U3781 (N_3781,In_1780,In_973);
nor U3782 (N_3782,In_2155,In_827);
xor U3783 (N_3783,In_529,In_384);
and U3784 (N_3784,In_794,In_321);
and U3785 (N_3785,In_1,In_1201);
nor U3786 (N_3786,In_623,In_1109);
nand U3787 (N_3787,In_1199,In_1096);
and U3788 (N_3788,In_358,In_2149);
and U3789 (N_3789,In_2394,In_1125);
nand U3790 (N_3790,In_1279,In_1400);
nor U3791 (N_3791,In_33,In_1355);
nand U3792 (N_3792,In_659,In_1876);
or U3793 (N_3793,In_2,In_1353);
xor U3794 (N_3794,In_2434,In_245);
nand U3795 (N_3795,In_1644,In_1543);
xor U3796 (N_3796,In_2036,In_2442);
nand U3797 (N_3797,In_252,In_2134);
or U3798 (N_3798,In_1101,In_2134);
xor U3799 (N_3799,In_2061,In_402);
xnor U3800 (N_3800,In_780,In_1885);
nor U3801 (N_3801,In_41,In_966);
xnor U3802 (N_3802,In_1077,In_1815);
nand U3803 (N_3803,In_2177,In_2400);
or U3804 (N_3804,In_1110,In_2327);
nor U3805 (N_3805,In_784,In_1591);
or U3806 (N_3806,In_1131,In_1969);
or U3807 (N_3807,In_481,In_1865);
xnor U3808 (N_3808,In_1507,In_94);
or U3809 (N_3809,In_576,In_2058);
xnor U3810 (N_3810,In_1006,In_2220);
or U3811 (N_3811,In_2304,In_249);
or U3812 (N_3812,In_947,In_697);
xnor U3813 (N_3813,In_1923,In_1445);
xnor U3814 (N_3814,In_2347,In_298);
xor U3815 (N_3815,In_1916,In_1169);
nand U3816 (N_3816,In_932,In_1648);
xor U3817 (N_3817,In_1049,In_2248);
or U3818 (N_3818,In_1406,In_185);
or U3819 (N_3819,In_1343,In_582);
xnor U3820 (N_3820,In_2496,In_2203);
xor U3821 (N_3821,In_957,In_1442);
or U3822 (N_3822,In_1818,In_1007);
xnor U3823 (N_3823,In_1798,In_231);
nand U3824 (N_3824,In_1542,In_2005);
xnor U3825 (N_3825,In_10,In_1768);
xor U3826 (N_3826,In_2478,In_328);
nand U3827 (N_3827,In_1757,In_2054);
nand U3828 (N_3828,In_2131,In_1525);
nand U3829 (N_3829,In_948,In_1600);
nor U3830 (N_3830,In_1739,In_1545);
xnor U3831 (N_3831,In_93,In_667);
nand U3832 (N_3832,In_1382,In_445);
and U3833 (N_3833,In_2382,In_1085);
xnor U3834 (N_3834,In_1350,In_2433);
nor U3835 (N_3835,In_1005,In_2128);
and U3836 (N_3836,In_396,In_1412);
xnor U3837 (N_3837,In_2183,In_1580);
xnor U3838 (N_3838,In_439,In_208);
nor U3839 (N_3839,In_2331,In_2307);
xnor U3840 (N_3840,In_1891,In_2082);
and U3841 (N_3841,In_832,In_2190);
and U3842 (N_3842,In_2313,In_279);
nor U3843 (N_3843,In_691,In_166);
nor U3844 (N_3844,In_117,In_1436);
and U3845 (N_3845,In_1068,In_503);
or U3846 (N_3846,In_1122,In_2458);
nor U3847 (N_3847,In_1640,In_1705);
nand U3848 (N_3848,In_165,In_329);
or U3849 (N_3849,In_2253,In_1643);
nor U3850 (N_3850,In_663,In_812);
xnor U3851 (N_3851,In_1369,In_563);
or U3852 (N_3852,In_1817,In_2234);
xor U3853 (N_3853,In_2132,In_2189);
nand U3854 (N_3854,In_513,In_418);
or U3855 (N_3855,In_1606,In_658);
nand U3856 (N_3856,In_1,In_2339);
and U3857 (N_3857,In_133,In_1338);
xnor U3858 (N_3858,In_95,In_234);
nor U3859 (N_3859,In_2287,In_865);
nand U3860 (N_3860,In_395,In_1657);
or U3861 (N_3861,In_1627,In_538);
nand U3862 (N_3862,In_14,In_2210);
nand U3863 (N_3863,In_1352,In_1935);
nand U3864 (N_3864,In_740,In_626);
nand U3865 (N_3865,In_1429,In_1541);
and U3866 (N_3866,In_1275,In_1987);
nor U3867 (N_3867,In_2279,In_264);
nand U3868 (N_3868,In_2255,In_618);
nand U3869 (N_3869,In_994,In_1719);
nand U3870 (N_3870,In_1317,In_1074);
nand U3871 (N_3871,In_212,In_766);
nor U3872 (N_3872,In_444,In_510);
xor U3873 (N_3873,In_1809,In_1298);
nor U3874 (N_3874,In_2387,In_796);
nor U3875 (N_3875,In_638,In_702);
xor U3876 (N_3876,In_138,In_1016);
and U3877 (N_3877,In_339,In_298);
nor U3878 (N_3878,In_1326,In_58);
nand U3879 (N_3879,In_458,In_1830);
xnor U3880 (N_3880,In_1292,In_2402);
xor U3881 (N_3881,In_387,In_19);
or U3882 (N_3882,In_2441,In_2285);
or U3883 (N_3883,In_1328,In_2363);
nor U3884 (N_3884,In_653,In_406);
nor U3885 (N_3885,In_172,In_2010);
nand U3886 (N_3886,In_751,In_2170);
and U3887 (N_3887,In_1522,In_1195);
or U3888 (N_3888,In_841,In_2240);
nor U3889 (N_3889,In_1213,In_1502);
nand U3890 (N_3890,In_2296,In_1606);
nor U3891 (N_3891,In_2127,In_2425);
nor U3892 (N_3892,In_312,In_1843);
or U3893 (N_3893,In_849,In_1712);
or U3894 (N_3894,In_958,In_2259);
nor U3895 (N_3895,In_1490,In_1861);
and U3896 (N_3896,In_2149,In_2265);
or U3897 (N_3897,In_2185,In_289);
nor U3898 (N_3898,In_1386,In_899);
and U3899 (N_3899,In_1187,In_603);
nor U3900 (N_3900,In_361,In_2496);
nor U3901 (N_3901,In_2149,In_1589);
xor U3902 (N_3902,In_1273,In_637);
or U3903 (N_3903,In_2483,In_2437);
nor U3904 (N_3904,In_1132,In_1405);
and U3905 (N_3905,In_984,In_525);
nor U3906 (N_3906,In_165,In_1373);
nand U3907 (N_3907,In_1213,In_1085);
nor U3908 (N_3908,In_1428,In_1750);
xor U3909 (N_3909,In_249,In_37);
nand U3910 (N_3910,In_2279,In_1668);
nand U3911 (N_3911,In_307,In_1688);
nor U3912 (N_3912,In_1929,In_1726);
and U3913 (N_3913,In_1247,In_1297);
nand U3914 (N_3914,In_650,In_2119);
and U3915 (N_3915,In_213,In_945);
and U3916 (N_3916,In_1733,In_2130);
and U3917 (N_3917,In_943,In_908);
nand U3918 (N_3918,In_708,In_1286);
nor U3919 (N_3919,In_360,In_1752);
or U3920 (N_3920,In_1128,In_202);
or U3921 (N_3921,In_915,In_92);
or U3922 (N_3922,In_1198,In_1022);
xnor U3923 (N_3923,In_2191,In_756);
nor U3924 (N_3924,In_941,In_1692);
nand U3925 (N_3925,In_2445,In_846);
or U3926 (N_3926,In_2214,In_189);
or U3927 (N_3927,In_1175,In_1079);
nand U3928 (N_3928,In_700,In_1210);
nand U3929 (N_3929,In_1203,In_770);
or U3930 (N_3930,In_1640,In_1367);
xnor U3931 (N_3931,In_1800,In_741);
nand U3932 (N_3932,In_2198,In_2234);
nand U3933 (N_3933,In_707,In_1332);
and U3934 (N_3934,In_1840,In_967);
or U3935 (N_3935,In_118,In_985);
or U3936 (N_3936,In_598,In_1518);
xnor U3937 (N_3937,In_1399,In_407);
nor U3938 (N_3938,In_978,In_1282);
nand U3939 (N_3939,In_1848,In_1604);
nand U3940 (N_3940,In_1548,In_1003);
xnor U3941 (N_3941,In_1837,In_1379);
and U3942 (N_3942,In_746,In_2151);
and U3943 (N_3943,In_655,In_1098);
xor U3944 (N_3944,In_2334,In_1446);
xor U3945 (N_3945,In_1982,In_1267);
nand U3946 (N_3946,In_2156,In_770);
and U3947 (N_3947,In_405,In_103);
xor U3948 (N_3948,In_838,In_2144);
or U3949 (N_3949,In_836,In_1753);
or U3950 (N_3950,In_36,In_792);
nand U3951 (N_3951,In_2125,In_276);
or U3952 (N_3952,In_2047,In_866);
and U3953 (N_3953,In_1031,In_1719);
nand U3954 (N_3954,In_1976,In_2189);
nand U3955 (N_3955,In_1543,In_337);
or U3956 (N_3956,In_831,In_1745);
or U3957 (N_3957,In_1328,In_1058);
nand U3958 (N_3958,In_2003,In_2225);
or U3959 (N_3959,In_1908,In_145);
and U3960 (N_3960,In_948,In_573);
or U3961 (N_3961,In_2467,In_1692);
nand U3962 (N_3962,In_2278,In_717);
nand U3963 (N_3963,In_344,In_754);
xnor U3964 (N_3964,In_1073,In_1680);
or U3965 (N_3965,In_2195,In_869);
nand U3966 (N_3966,In_2255,In_393);
and U3967 (N_3967,In_833,In_1413);
or U3968 (N_3968,In_75,In_1354);
or U3969 (N_3969,In_1806,In_1249);
or U3970 (N_3970,In_2168,In_1498);
nor U3971 (N_3971,In_2008,In_1556);
xnor U3972 (N_3972,In_563,In_577);
nor U3973 (N_3973,In_699,In_1582);
nand U3974 (N_3974,In_2117,In_1470);
nor U3975 (N_3975,In_1403,In_855);
xor U3976 (N_3976,In_248,In_458);
and U3977 (N_3977,In_1276,In_1767);
xnor U3978 (N_3978,In_89,In_1479);
and U3979 (N_3979,In_486,In_931);
xor U3980 (N_3980,In_943,In_550);
xor U3981 (N_3981,In_777,In_361);
or U3982 (N_3982,In_510,In_1484);
and U3983 (N_3983,In_2329,In_663);
or U3984 (N_3984,In_441,In_1137);
or U3985 (N_3985,In_1167,In_208);
nor U3986 (N_3986,In_1243,In_2388);
and U3987 (N_3987,In_1175,In_1214);
nor U3988 (N_3988,In_974,In_1853);
and U3989 (N_3989,In_444,In_1937);
nor U3990 (N_3990,In_1352,In_881);
nor U3991 (N_3991,In_2385,In_1094);
nand U3992 (N_3992,In_378,In_1607);
xor U3993 (N_3993,In_1725,In_237);
and U3994 (N_3994,In_35,In_2296);
xor U3995 (N_3995,In_344,In_2258);
nand U3996 (N_3996,In_370,In_1635);
or U3997 (N_3997,In_145,In_1423);
and U3998 (N_3998,In_209,In_1687);
nor U3999 (N_3999,In_2136,In_487);
xnor U4000 (N_4000,In_2123,In_588);
xnor U4001 (N_4001,In_130,In_867);
xor U4002 (N_4002,In_1159,In_2106);
xnor U4003 (N_4003,In_1489,In_590);
nor U4004 (N_4004,In_500,In_2250);
or U4005 (N_4005,In_453,In_581);
or U4006 (N_4006,In_1219,In_166);
nor U4007 (N_4007,In_2496,In_1918);
or U4008 (N_4008,In_301,In_1454);
and U4009 (N_4009,In_2291,In_1311);
or U4010 (N_4010,In_788,In_2480);
or U4011 (N_4011,In_1013,In_2438);
and U4012 (N_4012,In_942,In_2423);
or U4013 (N_4013,In_233,In_1913);
and U4014 (N_4014,In_1961,In_1378);
and U4015 (N_4015,In_547,In_2188);
and U4016 (N_4016,In_2404,In_152);
or U4017 (N_4017,In_1142,In_457);
nor U4018 (N_4018,In_915,In_1542);
xor U4019 (N_4019,In_541,In_1773);
and U4020 (N_4020,In_501,In_2295);
or U4021 (N_4021,In_51,In_1870);
nor U4022 (N_4022,In_1260,In_2089);
nand U4023 (N_4023,In_86,In_781);
nor U4024 (N_4024,In_525,In_1955);
nand U4025 (N_4025,In_1298,In_962);
and U4026 (N_4026,In_1876,In_187);
xor U4027 (N_4027,In_396,In_2360);
or U4028 (N_4028,In_1255,In_2471);
or U4029 (N_4029,In_1006,In_905);
nand U4030 (N_4030,In_719,In_384);
xnor U4031 (N_4031,In_321,In_2089);
xor U4032 (N_4032,In_734,In_2283);
nand U4033 (N_4033,In_334,In_2397);
xor U4034 (N_4034,In_518,In_2466);
and U4035 (N_4035,In_192,In_798);
xor U4036 (N_4036,In_1179,In_494);
or U4037 (N_4037,In_2006,In_1499);
or U4038 (N_4038,In_1110,In_1568);
xor U4039 (N_4039,In_2280,In_556);
nor U4040 (N_4040,In_1936,In_568);
nand U4041 (N_4041,In_1860,In_2287);
nand U4042 (N_4042,In_1995,In_2165);
nand U4043 (N_4043,In_1518,In_669);
xor U4044 (N_4044,In_585,In_1825);
or U4045 (N_4045,In_2172,In_649);
and U4046 (N_4046,In_110,In_539);
nand U4047 (N_4047,In_1961,In_1272);
and U4048 (N_4048,In_1249,In_2356);
and U4049 (N_4049,In_1679,In_1486);
and U4050 (N_4050,In_1607,In_230);
nand U4051 (N_4051,In_1419,In_961);
xor U4052 (N_4052,In_128,In_71);
xnor U4053 (N_4053,In_1535,In_806);
xnor U4054 (N_4054,In_256,In_1666);
nand U4055 (N_4055,In_1499,In_1444);
xnor U4056 (N_4056,In_154,In_2402);
xor U4057 (N_4057,In_1555,In_458);
and U4058 (N_4058,In_767,In_2408);
nand U4059 (N_4059,In_159,In_2482);
or U4060 (N_4060,In_1777,In_872);
nand U4061 (N_4061,In_159,In_2400);
or U4062 (N_4062,In_1637,In_2205);
xnor U4063 (N_4063,In_331,In_1995);
and U4064 (N_4064,In_2259,In_1084);
nand U4065 (N_4065,In_830,In_1051);
xnor U4066 (N_4066,In_1909,In_1445);
or U4067 (N_4067,In_1660,In_1438);
and U4068 (N_4068,In_2128,In_2035);
xor U4069 (N_4069,In_68,In_1267);
and U4070 (N_4070,In_1265,In_213);
nand U4071 (N_4071,In_2198,In_920);
xnor U4072 (N_4072,In_2242,In_1116);
or U4073 (N_4073,In_43,In_2141);
nor U4074 (N_4074,In_1422,In_1284);
nand U4075 (N_4075,In_1035,In_252);
nand U4076 (N_4076,In_349,In_2079);
nor U4077 (N_4077,In_2145,In_1730);
nand U4078 (N_4078,In_842,In_1648);
xor U4079 (N_4079,In_1087,In_2242);
nand U4080 (N_4080,In_208,In_948);
nand U4081 (N_4081,In_1135,In_1380);
nand U4082 (N_4082,In_2499,In_1501);
nand U4083 (N_4083,In_1945,In_1759);
or U4084 (N_4084,In_741,In_329);
or U4085 (N_4085,In_2096,In_1880);
nor U4086 (N_4086,In_1943,In_1664);
and U4087 (N_4087,In_919,In_1275);
and U4088 (N_4088,In_275,In_440);
or U4089 (N_4089,In_1085,In_213);
or U4090 (N_4090,In_393,In_2286);
and U4091 (N_4091,In_94,In_1696);
xor U4092 (N_4092,In_2383,In_123);
nor U4093 (N_4093,In_1951,In_1295);
and U4094 (N_4094,In_59,In_2443);
nand U4095 (N_4095,In_1726,In_1284);
nor U4096 (N_4096,In_755,In_2006);
xor U4097 (N_4097,In_481,In_181);
or U4098 (N_4098,In_1700,In_1059);
and U4099 (N_4099,In_1961,In_83);
xnor U4100 (N_4100,In_2134,In_2449);
nand U4101 (N_4101,In_912,In_1117);
xor U4102 (N_4102,In_342,In_2275);
or U4103 (N_4103,In_660,In_387);
nand U4104 (N_4104,In_473,In_1720);
xnor U4105 (N_4105,In_801,In_1018);
and U4106 (N_4106,In_1683,In_91);
and U4107 (N_4107,In_906,In_678);
nand U4108 (N_4108,In_2389,In_2473);
xor U4109 (N_4109,In_1629,In_522);
nand U4110 (N_4110,In_885,In_2079);
and U4111 (N_4111,In_1825,In_186);
and U4112 (N_4112,In_642,In_1810);
or U4113 (N_4113,In_718,In_1088);
nor U4114 (N_4114,In_734,In_1116);
xnor U4115 (N_4115,In_815,In_1518);
nand U4116 (N_4116,In_1468,In_1889);
and U4117 (N_4117,In_655,In_1632);
nand U4118 (N_4118,In_1448,In_1748);
nand U4119 (N_4119,In_815,In_1215);
nand U4120 (N_4120,In_106,In_906);
nand U4121 (N_4121,In_1702,In_1535);
and U4122 (N_4122,In_2378,In_1566);
or U4123 (N_4123,In_1211,In_1169);
nor U4124 (N_4124,In_2437,In_2051);
or U4125 (N_4125,In_604,In_2345);
or U4126 (N_4126,In_1468,In_639);
or U4127 (N_4127,In_1801,In_2024);
or U4128 (N_4128,In_301,In_131);
nor U4129 (N_4129,In_1317,In_547);
nand U4130 (N_4130,In_1848,In_341);
and U4131 (N_4131,In_2361,In_1819);
xor U4132 (N_4132,In_2271,In_2119);
or U4133 (N_4133,In_702,In_1559);
xor U4134 (N_4134,In_822,In_301);
and U4135 (N_4135,In_1313,In_418);
nor U4136 (N_4136,In_1095,In_236);
nand U4137 (N_4137,In_1363,In_4);
nor U4138 (N_4138,In_479,In_745);
nand U4139 (N_4139,In_764,In_373);
nand U4140 (N_4140,In_1864,In_216);
xor U4141 (N_4141,In_2320,In_1329);
and U4142 (N_4142,In_1917,In_2360);
and U4143 (N_4143,In_2321,In_966);
or U4144 (N_4144,In_2090,In_1287);
and U4145 (N_4145,In_2077,In_1348);
xor U4146 (N_4146,In_1746,In_94);
xnor U4147 (N_4147,In_306,In_93);
nor U4148 (N_4148,In_1373,In_4);
xnor U4149 (N_4149,In_477,In_2067);
or U4150 (N_4150,In_1506,In_1255);
or U4151 (N_4151,In_1940,In_983);
xor U4152 (N_4152,In_233,In_44);
nor U4153 (N_4153,In_1902,In_66);
xnor U4154 (N_4154,In_1378,In_908);
nor U4155 (N_4155,In_2022,In_1988);
and U4156 (N_4156,In_2474,In_1265);
xnor U4157 (N_4157,In_2356,In_1742);
nand U4158 (N_4158,In_637,In_1056);
and U4159 (N_4159,In_1896,In_1826);
nand U4160 (N_4160,In_778,In_1511);
or U4161 (N_4161,In_1562,In_2443);
and U4162 (N_4162,In_2449,In_870);
or U4163 (N_4163,In_204,In_1820);
xor U4164 (N_4164,In_1816,In_2481);
xnor U4165 (N_4165,In_1064,In_337);
nor U4166 (N_4166,In_2165,In_647);
nor U4167 (N_4167,In_1668,In_1172);
or U4168 (N_4168,In_2243,In_1380);
or U4169 (N_4169,In_2385,In_604);
xnor U4170 (N_4170,In_766,In_879);
xnor U4171 (N_4171,In_2195,In_1925);
or U4172 (N_4172,In_651,In_2045);
nand U4173 (N_4173,In_827,In_1873);
nor U4174 (N_4174,In_25,In_463);
or U4175 (N_4175,In_835,In_620);
xor U4176 (N_4176,In_695,In_843);
or U4177 (N_4177,In_533,In_2420);
xor U4178 (N_4178,In_286,In_1410);
xor U4179 (N_4179,In_1599,In_1821);
or U4180 (N_4180,In_2418,In_2076);
or U4181 (N_4181,In_810,In_1921);
and U4182 (N_4182,In_287,In_671);
or U4183 (N_4183,In_758,In_1915);
xnor U4184 (N_4184,In_1006,In_2273);
and U4185 (N_4185,In_937,In_1336);
and U4186 (N_4186,In_401,In_924);
and U4187 (N_4187,In_2261,In_553);
xor U4188 (N_4188,In_1626,In_1322);
and U4189 (N_4189,In_1405,In_590);
xnor U4190 (N_4190,In_1315,In_68);
xnor U4191 (N_4191,In_334,In_2242);
nor U4192 (N_4192,In_2156,In_931);
nor U4193 (N_4193,In_821,In_2060);
nand U4194 (N_4194,In_1177,In_2374);
xor U4195 (N_4195,In_455,In_1435);
or U4196 (N_4196,In_1269,In_2251);
nand U4197 (N_4197,In_2199,In_336);
xor U4198 (N_4198,In_1242,In_2397);
and U4199 (N_4199,In_1974,In_2381);
and U4200 (N_4200,In_2016,In_1071);
xor U4201 (N_4201,In_1590,In_565);
or U4202 (N_4202,In_641,In_2456);
nor U4203 (N_4203,In_1204,In_1355);
xnor U4204 (N_4204,In_517,In_1964);
or U4205 (N_4205,In_1320,In_412);
or U4206 (N_4206,In_1612,In_468);
or U4207 (N_4207,In_1576,In_1660);
and U4208 (N_4208,In_1328,In_490);
and U4209 (N_4209,In_1557,In_1718);
nand U4210 (N_4210,In_1595,In_1364);
or U4211 (N_4211,In_2408,In_2125);
xnor U4212 (N_4212,In_1221,In_1422);
and U4213 (N_4213,In_2164,In_185);
nand U4214 (N_4214,In_2098,In_1012);
nand U4215 (N_4215,In_1544,In_420);
xor U4216 (N_4216,In_613,In_2112);
nor U4217 (N_4217,In_759,In_2215);
or U4218 (N_4218,In_1909,In_2264);
nand U4219 (N_4219,In_1391,In_2128);
or U4220 (N_4220,In_2308,In_426);
nor U4221 (N_4221,In_2083,In_390);
or U4222 (N_4222,In_1440,In_2061);
xnor U4223 (N_4223,In_2245,In_159);
xor U4224 (N_4224,In_1618,In_2270);
and U4225 (N_4225,In_1153,In_1941);
xor U4226 (N_4226,In_664,In_1444);
xor U4227 (N_4227,In_1883,In_2225);
and U4228 (N_4228,In_329,In_160);
xor U4229 (N_4229,In_2027,In_483);
xnor U4230 (N_4230,In_1278,In_321);
or U4231 (N_4231,In_2430,In_1804);
and U4232 (N_4232,In_943,In_384);
nor U4233 (N_4233,In_309,In_1208);
or U4234 (N_4234,In_1059,In_2407);
xor U4235 (N_4235,In_2395,In_262);
xnor U4236 (N_4236,In_1848,In_1724);
nand U4237 (N_4237,In_267,In_2116);
and U4238 (N_4238,In_1491,In_2195);
and U4239 (N_4239,In_1886,In_240);
and U4240 (N_4240,In_1284,In_1094);
xor U4241 (N_4241,In_1940,In_188);
nand U4242 (N_4242,In_2445,In_2040);
and U4243 (N_4243,In_867,In_2301);
or U4244 (N_4244,In_1122,In_1851);
and U4245 (N_4245,In_60,In_1649);
xnor U4246 (N_4246,In_1277,In_1344);
nor U4247 (N_4247,In_2188,In_77);
nor U4248 (N_4248,In_1543,In_388);
or U4249 (N_4249,In_1294,In_1017);
xor U4250 (N_4250,In_845,In_1584);
nor U4251 (N_4251,In_420,In_242);
xor U4252 (N_4252,In_986,In_1154);
nand U4253 (N_4253,In_1291,In_2408);
xor U4254 (N_4254,In_430,In_9);
xor U4255 (N_4255,In_1591,In_1335);
nor U4256 (N_4256,In_607,In_664);
nand U4257 (N_4257,In_63,In_120);
nand U4258 (N_4258,In_977,In_292);
nand U4259 (N_4259,In_670,In_2210);
or U4260 (N_4260,In_1667,In_1127);
and U4261 (N_4261,In_1869,In_1688);
or U4262 (N_4262,In_325,In_506);
nor U4263 (N_4263,In_343,In_1506);
nand U4264 (N_4264,In_1629,In_87);
xnor U4265 (N_4265,In_2218,In_974);
nor U4266 (N_4266,In_453,In_422);
nand U4267 (N_4267,In_1556,In_2226);
or U4268 (N_4268,In_1293,In_1843);
xor U4269 (N_4269,In_447,In_2402);
nand U4270 (N_4270,In_147,In_2217);
nand U4271 (N_4271,In_1527,In_1006);
or U4272 (N_4272,In_904,In_511);
or U4273 (N_4273,In_558,In_282);
or U4274 (N_4274,In_1073,In_1495);
nor U4275 (N_4275,In_1221,In_2128);
or U4276 (N_4276,In_58,In_273);
and U4277 (N_4277,In_2236,In_1203);
nor U4278 (N_4278,In_2195,In_2015);
xnor U4279 (N_4279,In_691,In_1799);
or U4280 (N_4280,In_1943,In_810);
xnor U4281 (N_4281,In_708,In_1423);
or U4282 (N_4282,In_1348,In_30);
or U4283 (N_4283,In_809,In_1337);
xor U4284 (N_4284,In_1235,In_2300);
nand U4285 (N_4285,In_1083,In_2424);
nor U4286 (N_4286,In_1833,In_1905);
xor U4287 (N_4287,In_1880,In_1573);
xnor U4288 (N_4288,In_279,In_296);
and U4289 (N_4289,In_1724,In_625);
nor U4290 (N_4290,In_2268,In_262);
nand U4291 (N_4291,In_1109,In_689);
xor U4292 (N_4292,In_25,In_2354);
or U4293 (N_4293,In_809,In_2221);
nand U4294 (N_4294,In_2054,In_2229);
and U4295 (N_4295,In_984,In_1636);
nor U4296 (N_4296,In_2169,In_2497);
and U4297 (N_4297,In_965,In_1830);
or U4298 (N_4298,In_744,In_2283);
and U4299 (N_4299,In_1435,In_611);
nor U4300 (N_4300,In_57,In_1336);
xnor U4301 (N_4301,In_321,In_1021);
nor U4302 (N_4302,In_2489,In_2129);
and U4303 (N_4303,In_44,In_931);
or U4304 (N_4304,In_1069,In_1637);
nand U4305 (N_4305,In_567,In_1609);
and U4306 (N_4306,In_1739,In_2150);
nand U4307 (N_4307,In_2423,In_435);
and U4308 (N_4308,In_1732,In_539);
xor U4309 (N_4309,In_2432,In_1572);
xnor U4310 (N_4310,In_821,In_1584);
nor U4311 (N_4311,In_1824,In_519);
xor U4312 (N_4312,In_1920,In_1351);
nand U4313 (N_4313,In_1389,In_1265);
nand U4314 (N_4314,In_2305,In_1498);
and U4315 (N_4315,In_152,In_2230);
or U4316 (N_4316,In_655,In_2439);
or U4317 (N_4317,In_2126,In_645);
nand U4318 (N_4318,In_490,In_2369);
nor U4319 (N_4319,In_1983,In_347);
nor U4320 (N_4320,In_371,In_351);
nor U4321 (N_4321,In_133,In_2159);
nor U4322 (N_4322,In_1274,In_1161);
or U4323 (N_4323,In_1753,In_692);
or U4324 (N_4324,In_1057,In_941);
nand U4325 (N_4325,In_1479,In_2401);
nor U4326 (N_4326,In_1993,In_1154);
nor U4327 (N_4327,In_1182,In_1214);
nor U4328 (N_4328,In_543,In_2444);
xor U4329 (N_4329,In_729,In_175);
nand U4330 (N_4330,In_54,In_241);
or U4331 (N_4331,In_467,In_844);
nor U4332 (N_4332,In_308,In_318);
nand U4333 (N_4333,In_506,In_1646);
nor U4334 (N_4334,In_720,In_77);
nor U4335 (N_4335,In_1378,In_163);
nor U4336 (N_4336,In_2227,In_1516);
or U4337 (N_4337,In_1988,In_1125);
nor U4338 (N_4338,In_330,In_1958);
nor U4339 (N_4339,In_554,In_1565);
or U4340 (N_4340,In_2092,In_1102);
or U4341 (N_4341,In_816,In_1540);
nor U4342 (N_4342,In_243,In_2028);
or U4343 (N_4343,In_37,In_1313);
nor U4344 (N_4344,In_2025,In_111);
nand U4345 (N_4345,In_2385,In_1461);
or U4346 (N_4346,In_2494,In_471);
xnor U4347 (N_4347,In_106,In_1800);
xnor U4348 (N_4348,In_1597,In_812);
and U4349 (N_4349,In_941,In_2436);
and U4350 (N_4350,In_373,In_1484);
and U4351 (N_4351,In_2234,In_991);
nor U4352 (N_4352,In_2383,In_328);
or U4353 (N_4353,In_870,In_431);
xnor U4354 (N_4354,In_2357,In_89);
or U4355 (N_4355,In_2354,In_1586);
nand U4356 (N_4356,In_2017,In_1025);
xnor U4357 (N_4357,In_1894,In_839);
nand U4358 (N_4358,In_1710,In_2060);
and U4359 (N_4359,In_536,In_1688);
xnor U4360 (N_4360,In_84,In_284);
and U4361 (N_4361,In_2184,In_1547);
and U4362 (N_4362,In_2480,In_188);
nand U4363 (N_4363,In_1557,In_2106);
and U4364 (N_4364,In_726,In_1272);
or U4365 (N_4365,In_566,In_2447);
or U4366 (N_4366,In_1941,In_289);
or U4367 (N_4367,In_1082,In_711);
nand U4368 (N_4368,In_1704,In_169);
or U4369 (N_4369,In_2050,In_570);
or U4370 (N_4370,In_1630,In_2167);
xnor U4371 (N_4371,In_1822,In_475);
nor U4372 (N_4372,In_750,In_863);
and U4373 (N_4373,In_1931,In_264);
and U4374 (N_4374,In_1438,In_2229);
nand U4375 (N_4375,In_860,In_2318);
and U4376 (N_4376,In_1082,In_1211);
nand U4377 (N_4377,In_1856,In_2368);
nor U4378 (N_4378,In_1818,In_1032);
nand U4379 (N_4379,In_784,In_2402);
nor U4380 (N_4380,In_761,In_1396);
xnor U4381 (N_4381,In_236,In_1272);
nor U4382 (N_4382,In_321,In_437);
xor U4383 (N_4383,In_1429,In_1690);
and U4384 (N_4384,In_58,In_243);
or U4385 (N_4385,In_2003,In_72);
xnor U4386 (N_4386,In_1433,In_273);
or U4387 (N_4387,In_1376,In_111);
xor U4388 (N_4388,In_2309,In_2358);
xor U4389 (N_4389,In_2147,In_1809);
or U4390 (N_4390,In_1615,In_696);
xor U4391 (N_4391,In_296,In_477);
nand U4392 (N_4392,In_1346,In_847);
nor U4393 (N_4393,In_307,In_1985);
and U4394 (N_4394,In_445,In_704);
and U4395 (N_4395,In_1568,In_2455);
or U4396 (N_4396,In_588,In_1215);
xnor U4397 (N_4397,In_1477,In_2029);
nor U4398 (N_4398,In_1724,In_336);
and U4399 (N_4399,In_318,In_1539);
nor U4400 (N_4400,In_228,In_1844);
xor U4401 (N_4401,In_663,In_387);
and U4402 (N_4402,In_2408,In_1362);
nor U4403 (N_4403,In_91,In_89);
and U4404 (N_4404,In_886,In_295);
nand U4405 (N_4405,In_371,In_2177);
nor U4406 (N_4406,In_1223,In_815);
nor U4407 (N_4407,In_1603,In_1025);
nor U4408 (N_4408,In_1277,In_531);
xnor U4409 (N_4409,In_1842,In_295);
nor U4410 (N_4410,In_672,In_2190);
xor U4411 (N_4411,In_124,In_881);
nand U4412 (N_4412,In_1634,In_1042);
xor U4413 (N_4413,In_706,In_653);
and U4414 (N_4414,In_397,In_2429);
nor U4415 (N_4415,In_1827,In_1246);
or U4416 (N_4416,In_458,In_342);
and U4417 (N_4417,In_37,In_1783);
nand U4418 (N_4418,In_233,In_200);
xor U4419 (N_4419,In_220,In_834);
xnor U4420 (N_4420,In_2112,In_2303);
nand U4421 (N_4421,In_825,In_2444);
nand U4422 (N_4422,In_1011,In_45);
or U4423 (N_4423,In_1583,In_2350);
nor U4424 (N_4424,In_2150,In_888);
or U4425 (N_4425,In_1306,In_1318);
or U4426 (N_4426,In_264,In_2238);
and U4427 (N_4427,In_2050,In_1778);
and U4428 (N_4428,In_517,In_494);
or U4429 (N_4429,In_1096,In_1537);
xnor U4430 (N_4430,In_332,In_65);
nand U4431 (N_4431,In_1443,In_982);
xnor U4432 (N_4432,In_2492,In_1066);
nand U4433 (N_4433,In_1396,In_23);
xor U4434 (N_4434,In_245,In_2498);
nor U4435 (N_4435,In_2046,In_873);
xnor U4436 (N_4436,In_1859,In_737);
xnor U4437 (N_4437,In_733,In_2288);
and U4438 (N_4438,In_860,In_908);
nor U4439 (N_4439,In_1370,In_1779);
xor U4440 (N_4440,In_276,In_2285);
and U4441 (N_4441,In_1685,In_133);
or U4442 (N_4442,In_2219,In_1880);
or U4443 (N_4443,In_694,In_2172);
nand U4444 (N_4444,In_688,In_2324);
nand U4445 (N_4445,In_2342,In_848);
nand U4446 (N_4446,In_1677,In_1497);
xnor U4447 (N_4447,In_294,In_524);
xnor U4448 (N_4448,In_712,In_2462);
nand U4449 (N_4449,In_2276,In_1170);
or U4450 (N_4450,In_1287,In_2425);
nand U4451 (N_4451,In_1629,In_1935);
nor U4452 (N_4452,In_999,In_933);
nor U4453 (N_4453,In_885,In_775);
and U4454 (N_4454,In_2376,In_1937);
nor U4455 (N_4455,In_2175,In_1144);
nand U4456 (N_4456,In_449,In_1515);
nand U4457 (N_4457,In_1682,In_991);
and U4458 (N_4458,In_1610,In_2233);
nand U4459 (N_4459,In_875,In_746);
nand U4460 (N_4460,In_1407,In_26);
xor U4461 (N_4461,In_954,In_1403);
or U4462 (N_4462,In_2283,In_1999);
nand U4463 (N_4463,In_19,In_1098);
xnor U4464 (N_4464,In_1889,In_1947);
nand U4465 (N_4465,In_1349,In_2375);
and U4466 (N_4466,In_693,In_2371);
nand U4467 (N_4467,In_846,In_1001);
and U4468 (N_4468,In_2476,In_83);
nor U4469 (N_4469,In_1069,In_464);
and U4470 (N_4470,In_2431,In_81);
and U4471 (N_4471,In_1945,In_489);
nor U4472 (N_4472,In_243,In_1381);
and U4473 (N_4473,In_415,In_1112);
xnor U4474 (N_4474,In_1519,In_110);
xor U4475 (N_4475,In_2106,In_720);
nand U4476 (N_4476,In_2173,In_1822);
and U4477 (N_4477,In_1792,In_562);
nor U4478 (N_4478,In_1172,In_2124);
and U4479 (N_4479,In_2044,In_590);
and U4480 (N_4480,In_86,In_293);
nand U4481 (N_4481,In_684,In_1589);
nand U4482 (N_4482,In_58,In_2142);
or U4483 (N_4483,In_838,In_1363);
and U4484 (N_4484,In_430,In_205);
or U4485 (N_4485,In_2329,In_2268);
xor U4486 (N_4486,In_274,In_1096);
and U4487 (N_4487,In_2041,In_2446);
xor U4488 (N_4488,In_710,In_2065);
nor U4489 (N_4489,In_2022,In_1078);
and U4490 (N_4490,In_1812,In_1806);
and U4491 (N_4491,In_2278,In_1348);
and U4492 (N_4492,In_746,In_296);
and U4493 (N_4493,In_1438,In_774);
nand U4494 (N_4494,In_268,In_1679);
nand U4495 (N_4495,In_941,In_711);
nand U4496 (N_4496,In_1222,In_1412);
nand U4497 (N_4497,In_1690,In_1459);
nand U4498 (N_4498,In_2274,In_2277);
xor U4499 (N_4499,In_2043,In_1378);
or U4500 (N_4500,In_511,In_2205);
xor U4501 (N_4501,In_1997,In_2024);
and U4502 (N_4502,In_2476,In_2484);
or U4503 (N_4503,In_1066,In_527);
or U4504 (N_4504,In_2170,In_239);
and U4505 (N_4505,In_936,In_691);
and U4506 (N_4506,In_713,In_1014);
nand U4507 (N_4507,In_370,In_1278);
or U4508 (N_4508,In_2441,In_2035);
nor U4509 (N_4509,In_944,In_262);
or U4510 (N_4510,In_2495,In_524);
and U4511 (N_4511,In_2172,In_124);
nor U4512 (N_4512,In_183,In_1195);
nor U4513 (N_4513,In_1352,In_1051);
or U4514 (N_4514,In_1923,In_804);
and U4515 (N_4515,In_283,In_1520);
nand U4516 (N_4516,In_2404,In_864);
nand U4517 (N_4517,In_40,In_947);
nand U4518 (N_4518,In_2336,In_1383);
and U4519 (N_4519,In_1223,In_547);
or U4520 (N_4520,In_1997,In_2156);
nand U4521 (N_4521,In_2433,In_69);
or U4522 (N_4522,In_2460,In_730);
or U4523 (N_4523,In_724,In_1722);
xnor U4524 (N_4524,In_804,In_2280);
or U4525 (N_4525,In_922,In_1073);
xnor U4526 (N_4526,In_1276,In_1082);
and U4527 (N_4527,In_1926,In_1050);
nand U4528 (N_4528,In_893,In_2153);
xor U4529 (N_4529,In_1705,In_1507);
and U4530 (N_4530,In_855,In_2376);
xor U4531 (N_4531,In_486,In_2378);
xor U4532 (N_4532,In_2387,In_1199);
nand U4533 (N_4533,In_1132,In_314);
nand U4534 (N_4534,In_2360,In_1035);
nor U4535 (N_4535,In_496,In_491);
nor U4536 (N_4536,In_1999,In_233);
and U4537 (N_4537,In_365,In_1686);
nor U4538 (N_4538,In_29,In_274);
xnor U4539 (N_4539,In_1570,In_314);
nand U4540 (N_4540,In_631,In_2213);
and U4541 (N_4541,In_886,In_1065);
or U4542 (N_4542,In_715,In_1098);
nor U4543 (N_4543,In_552,In_2182);
nor U4544 (N_4544,In_741,In_991);
or U4545 (N_4545,In_1674,In_243);
or U4546 (N_4546,In_1964,In_1330);
and U4547 (N_4547,In_872,In_1555);
or U4548 (N_4548,In_1727,In_230);
nand U4549 (N_4549,In_495,In_2257);
nand U4550 (N_4550,In_1339,In_2023);
nor U4551 (N_4551,In_1991,In_619);
or U4552 (N_4552,In_570,In_1489);
nand U4553 (N_4553,In_565,In_1217);
and U4554 (N_4554,In_1720,In_504);
nand U4555 (N_4555,In_2243,In_1855);
or U4556 (N_4556,In_1291,In_124);
and U4557 (N_4557,In_1609,In_882);
xor U4558 (N_4558,In_798,In_1354);
and U4559 (N_4559,In_1126,In_580);
or U4560 (N_4560,In_1313,In_1579);
xnor U4561 (N_4561,In_2228,In_354);
nand U4562 (N_4562,In_1561,In_1801);
nand U4563 (N_4563,In_797,In_116);
and U4564 (N_4564,In_1037,In_1346);
and U4565 (N_4565,In_215,In_2379);
xor U4566 (N_4566,In_2046,In_474);
nor U4567 (N_4567,In_462,In_1384);
xnor U4568 (N_4568,In_1602,In_2194);
and U4569 (N_4569,In_2108,In_2025);
nand U4570 (N_4570,In_497,In_834);
and U4571 (N_4571,In_224,In_652);
xnor U4572 (N_4572,In_2029,In_1349);
and U4573 (N_4573,In_1472,In_2299);
nand U4574 (N_4574,In_1486,In_1015);
xor U4575 (N_4575,In_719,In_2151);
nor U4576 (N_4576,In_885,In_1371);
and U4577 (N_4577,In_1838,In_1293);
nand U4578 (N_4578,In_1825,In_2046);
nand U4579 (N_4579,In_1097,In_661);
and U4580 (N_4580,In_1987,In_454);
and U4581 (N_4581,In_539,In_909);
or U4582 (N_4582,In_85,In_1345);
and U4583 (N_4583,In_2134,In_1909);
or U4584 (N_4584,In_461,In_151);
nand U4585 (N_4585,In_2442,In_826);
xnor U4586 (N_4586,In_2233,In_2012);
or U4587 (N_4587,In_23,In_1207);
nand U4588 (N_4588,In_1603,In_813);
xnor U4589 (N_4589,In_582,In_395);
nor U4590 (N_4590,In_1075,In_1576);
or U4591 (N_4591,In_2455,In_823);
and U4592 (N_4592,In_106,In_224);
nand U4593 (N_4593,In_524,In_1373);
xor U4594 (N_4594,In_2341,In_762);
or U4595 (N_4595,In_1863,In_1120);
and U4596 (N_4596,In_437,In_2063);
and U4597 (N_4597,In_1833,In_1636);
nand U4598 (N_4598,In_1816,In_1118);
nand U4599 (N_4599,In_1115,In_1590);
nand U4600 (N_4600,In_621,In_1655);
xor U4601 (N_4601,In_1920,In_1617);
or U4602 (N_4602,In_578,In_1207);
nand U4603 (N_4603,In_1154,In_1755);
nor U4604 (N_4604,In_13,In_67);
or U4605 (N_4605,In_818,In_458);
nand U4606 (N_4606,In_482,In_391);
xnor U4607 (N_4607,In_1022,In_1093);
xnor U4608 (N_4608,In_965,In_110);
xor U4609 (N_4609,In_967,In_1816);
or U4610 (N_4610,In_1078,In_271);
nor U4611 (N_4611,In_84,In_343);
and U4612 (N_4612,In_1479,In_968);
nor U4613 (N_4613,In_2426,In_249);
nor U4614 (N_4614,In_508,In_1438);
xnor U4615 (N_4615,In_411,In_2011);
xnor U4616 (N_4616,In_1629,In_370);
and U4617 (N_4617,In_688,In_1907);
or U4618 (N_4618,In_1080,In_921);
or U4619 (N_4619,In_647,In_2368);
and U4620 (N_4620,In_1603,In_678);
xor U4621 (N_4621,In_1117,In_691);
nand U4622 (N_4622,In_448,In_507);
nand U4623 (N_4623,In_1700,In_880);
and U4624 (N_4624,In_1803,In_37);
and U4625 (N_4625,In_615,In_491);
nand U4626 (N_4626,In_1053,In_398);
xor U4627 (N_4627,In_333,In_2285);
nor U4628 (N_4628,In_1419,In_233);
or U4629 (N_4629,In_559,In_130);
or U4630 (N_4630,In_589,In_1928);
or U4631 (N_4631,In_1228,In_2312);
nor U4632 (N_4632,In_1236,In_1060);
xor U4633 (N_4633,In_684,In_1493);
or U4634 (N_4634,In_360,In_2078);
and U4635 (N_4635,In_1810,In_1189);
or U4636 (N_4636,In_1112,In_821);
nand U4637 (N_4637,In_2315,In_263);
or U4638 (N_4638,In_1586,In_658);
and U4639 (N_4639,In_1826,In_1555);
xnor U4640 (N_4640,In_1690,In_1251);
nand U4641 (N_4641,In_754,In_1282);
xor U4642 (N_4642,In_1849,In_1511);
nor U4643 (N_4643,In_2392,In_2329);
xnor U4644 (N_4644,In_939,In_2078);
nand U4645 (N_4645,In_1174,In_1133);
and U4646 (N_4646,In_557,In_1076);
nand U4647 (N_4647,In_1396,In_1952);
or U4648 (N_4648,In_682,In_258);
or U4649 (N_4649,In_890,In_221);
nor U4650 (N_4650,In_1597,In_1116);
nand U4651 (N_4651,In_2433,In_2454);
or U4652 (N_4652,In_159,In_1382);
xnor U4653 (N_4653,In_231,In_1729);
nand U4654 (N_4654,In_1266,In_2453);
nand U4655 (N_4655,In_1667,In_1952);
nand U4656 (N_4656,In_1700,In_179);
or U4657 (N_4657,In_2238,In_655);
or U4658 (N_4658,In_556,In_1101);
xor U4659 (N_4659,In_1444,In_1120);
nor U4660 (N_4660,In_1421,In_1919);
xnor U4661 (N_4661,In_805,In_669);
and U4662 (N_4662,In_1724,In_1928);
nor U4663 (N_4663,In_1579,In_2008);
or U4664 (N_4664,In_631,In_739);
nand U4665 (N_4665,In_257,In_242);
and U4666 (N_4666,In_1313,In_2160);
or U4667 (N_4667,In_1109,In_2353);
or U4668 (N_4668,In_2141,In_395);
and U4669 (N_4669,In_2433,In_349);
xnor U4670 (N_4670,In_1886,In_115);
and U4671 (N_4671,In_2424,In_454);
xor U4672 (N_4672,In_1344,In_852);
xor U4673 (N_4673,In_2445,In_1541);
and U4674 (N_4674,In_2017,In_1632);
or U4675 (N_4675,In_166,In_1617);
xnor U4676 (N_4676,In_918,In_1799);
or U4677 (N_4677,In_2257,In_1779);
or U4678 (N_4678,In_2113,In_501);
or U4679 (N_4679,In_1110,In_641);
or U4680 (N_4680,In_1575,In_1097);
or U4681 (N_4681,In_474,In_1086);
nand U4682 (N_4682,In_2044,In_501);
or U4683 (N_4683,In_1684,In_1559);
and U4684 (N_4684,In_1172,In_1576);
and U4685 (N_4685,In_536,In_814);
nor U4686 (N_4686,In_2492,In_1746);
nand U4687 (N_4687,In_988,In_103);
nand U4688 (N_4688,In_307,In_2306);
nor U4689 (N_4689,In_755,In_1016);
or U4690 (N_4690,In_1040,In_663);
nor U4691 (N_4691,In_1948,In_110);
and U4692 (N_4692,In_208,In_748);
and U4693 (N_4693,In_940,In_1944);
and U4694 (N_4694,In_1982,In_390);
nand U4695 (N_4695,In_1789,In_1062);
nor U4696 (N_4696,In_29,In_191);
xor U4697 (N_4697,In_39,In_513);
or U4698 (N_4698,In_135,In_1578);
nor U4699 (N_4699,In_216,In_2397);
nand U4700 (N_4700,In_960,In_805);
nand U4701 (N_4701,In_1961,In_497);
or U4702 (N_4702,In_1596,In_114);
and U4703 (N_4703,In_1891,In_2486);
nand U4704 (N_4704,In_901,In_1478);
or U4705 (N_4705,In_1045,In_621);
and U4706 (N_4706,In_1426,In_1548);
nand U4707 (N_4707,In_1993,In_354);
and U4708 (N_4708,In_1845,In_436);
nor U4709 (N_4709,In_2102,In_1434);
or U4710 (N_4710,In_1191,In_1051);
and U4711 (N_4711,In_1302,In_1649);
or U4712 (N_4712,In_1186,In_1336);
and U4713 (N_4713,In_1134,In_2241);
xnor U4714 (N_4714,In_1821,In_1335);
xnor U4715 (N_4715,In_1199,In_1371);
or U4716 (N_4716,In_1134,In_1066);
nor U4717 (N_4717,In_1130,In_1368);
and U4718 (N_4718,In_2008,In_1601);
or U4719 (N_4719,In_167,In_753);
nor U4720 (N_4720,In_714,In_1353);
nor U4721 (N_4721,In_449,In_969);
xnor U4722 (N_4722,In_1942,In_614);
or U4723 (N_4723,In_611,In_253);
or U4724 (N_4724,In_2169,In_1597);
nor U4725 (N_4725,In_2217,In_1032);
or U4726 (N_4726,In_2195,In_817);
xor U4727 (N_4727,In_1510,In_521);
nor U4728 (N_4728,In_1382,In_1622);
xor U4729 (N_4729,In_1872,In_2126);
xnor U4730 (N_4730,In_1099,In_578);
and U4731 (N_4731,In_275,In_1303);
nor U4732 (N_4732,In_2162,In_2227);
nor U4733 (N_4733,In_2364,In_2021);
nor U4734 (N_4734,In_1890,In_2014);
or U4735 (N_4735,In_547,In_325);
nor U4736 (N_4736,In_2094,In_257);
xnor U4737 (N_4737,In_327,In_1117);
and U4738 (N_4738,In_546,In_2268);
xnor U4739 (N_4739,In_2429,In_937);
xnor U4740 (N_4740,In_2140,In_423);
xnor U4741 (N_4741,In_308,In_1455);
nor U4742 (N_4742,In_2499,In_866);
or U4743 (N_4743,In_52,In_370);
xor U4744 (N_4744,In_2324,In_597);
and U4745 (N_4745,In_1860,In_1459);
xnor U4746 (N_4746,In_165,In_2435);
or U4747 (N_4747,In_2063,In_1859);
nand U4748 (N_4748,In_1810,In_250);
nor U4749 (N_4749,In_1867,In_864);
nand U4750 (N_4750,In_2222,In_1069);
nand U4751 (N_4751,In_1778,In_2318);
xor U4752 (N_4752,In_2143,In_696);
nand U4753 (N_4753,In_866,In_2384);
nor U4754 (N_4754,In_272,In_1265);
or U4755 (N_4755,In_378,In_1398);
nor U4756 (N_4756,In_792,In_2227);
and U4757 (N_4757,In_753,In_1481);
nand U4758 (N_4758,In_790,In_2042);
xnor U4759 (N_4759,In_2296,In_1918);
or U4760 (N_4760,In_2092,In_1357);
nor U4761 (N_4761,In_165,In_1088);
nand U4762 (N_4762,In_2225,In_1713);
or U4763 (N_4763,In_389,In_1878);
xnor U4764 (N_4764,In_1413,In_49);
and U4765 (N_4765,In_1670,In_173);
and U4766 (N_4766,In_1621,In_1593);
xor U4767 (N_4767,In_1810,In_1496);
and U4768 (N_4768,In_17,In_7);
or U4769 (N_4769,In_783,In_1605);
nand U4770 (N_4770,In_2174,In_2490);
nand U4771 (N_4771,In_1130,In_1945);
nand U4772 (N_4772,In_107,In_1645);
nor U4773 (N_4773,In_1863,In_1289);
nand U4774 (N_4774,In_95,In_1422);
nor U4775 (N_4775,In_605,In_2189);
nor U4776 (N_4776,In_2017,In_118);
and U4777 (N_4777,In_387,In_2488);
and U4778 (N_4778,In_695,In_1460);
nor U4779 (N_4779,In_1788,In_1037);
and U4780 (N_4780,In_1869,In_65);
nor U4781 (N_4781,In_1437,In_1894);
or U4782 (N_4782,In_1452,In_1134);
nand U4783 (N_4783,In_352,In_1950);
and U4784 (N_4784,In_29,In_1178);
nor U4785 (N_4785,In_599,In_83);
or U4786 (N_4786,In_839,In_2212);
nand U4787 (N_4787,In_859,In_68);
nand U4788 (N_4788,In_2016,In_26);
or U4789 (N_4789,In_1400,In_633);
xor U4790 (N_4790,In_560,In_801);
or U4791 (N_4791,In_2035,In_432);
nor U4792 (N_4792,In_875,In_1183);
nor U4793 (N_4793,In_1267,In_2133);
nand U4794 (N_4794,In_1587,In_314);
xnor U4795 (N_4795,In_466,In_132);
nor U4796 (N_4796,In_827,In_596);
and U4797 (N_4797,In_1773,In_1893);
nor U4798 (N_4798,In_1319,In_730);
nand U4799 (N_4799,In_2351,In_2435);
xor U4800 (N_4800,In_1713,In_1898);
nand U4801 (N_4801,In_2118,In_1475);
and U4802 (N_4802,In_1757,In_885);
nand U4803 (N_4803,In_1497,In_1768);
or U4804 (N_4804,In_1133,In_1462);
and U4805 (N_4805,In_2216,In_2234);
nand U4806 (N_4806,In_1189,In_879);
xnor U4807 (N_4807,In_351,In_879);
nand U4808 (N_4808,In_1819,In_1524);
and U4809 (N_4809,In_997,In_35);
and U4810 (N_4810,In_536,In_1256);
or U4811 (N_4811,In_1499,In_1240);
nand U4812 (N_4812,In_426,In_154);
nor U4813 (N_4813,In_876,In_549);
and U4814 (N_4814,In_313,In_842);
or U4815 (N_4815,In_1010,In_2014);
or U4816 (N_4816,In_606,In_2003);
xnor U4817 (N_4817,In_486,In_1386);
nand U4818 (N_4818,In_228,In_448);
and U4819 (N_4819,In_869,In_1457);
nand U4820 (N_4820,In_1130,In_869);
xor U4821 (N_4821,In_1638,In_1941);
nor U4822 (N_4822,In_97,In_2116);
nand U4823 (N_4823,In_1884,In_1590);
xor U4824 (N_4824,In_2125,In_1214);
nor U4825 (N_4825,In_107,In_2000);
and U4826 (N_4826,In_2208,In_774);
xnor U4827 (N_4827,In_48,In_1727);
nor U4828 (N_4828,In_1659,In_135);
and U4829 (N_4829,In_966,In_2302);
nor U4830 (N_4830,In_711,In_930);
and U4831 (N_4831,In_350,In_2260);
nand U4832 (N_4832,In_586,In_1575);
and U4833 (N_4833,In_1255,In_140);
xnor U4834 (N_4834,In_2267,In_250);
or U4835 (N_4835,In_115,In_699);
or U4836 (N_4836,In_1107,In_1981);
and U4837 (N_4837,In_1476,In_1661);
nor U4838 (N_4838,In_1030,In_334);
and U4839 (N_4839,In_1652,In_1971);
and U4840 (N_4840,In_2028,In_75);
or U4841 (N_4841,In_963,In_1051);
xor U4842 (N_4842,In_1615,In_958);
nand U4843 (N_4843,In_366,In_2428);
nand U4844 (N_4844,In_1611,In_1724);
nand U4845 (N_4845,In_149,In_2073);
nand U4846 (N_4846,In_1529,In_1299);
nand U4847 (N_4847,In_15,In_502);
or U4848 (N_4848,In_1756,In_919);
or U4849 (N_4849,In_349,In_606);
nor U4850 (N_4850,In_1879,In_747);
xnor U4851 (N_4851,In_2261,In_1717);
or U4852 (N_4852,In_520,In_1908);
nor U4853 (N_4853,In_1743,In_2004);
nor U4854 (N_4854,In_525,In_329);
xnor U4855 (N_4855,In_45,In_2333);
xnor U4856 (N_4856,In_2478,In_4);
and U4857 (N_4857,In_776,In_1634);
and U4858 (N_4858,In_2101,In_1087);
nor U4859 (N_4859,In_1651,In_1480);
xnor U4860 (N_4860,In_562,In_2446);
and U4861 (N_4861,In_1340,In_453);
xor U4862 (N_4862,In_1538,In_809);
and U4863 (N_4863,In_1071,In_1358);
nor U4864 (N_4864,In_1680,In_315);
and U4865 (N_4865,In_1842,In_1148);
nor U4866 (N_4866,In_813,In_17);
and U4867 (N_4867,In_291,In_1359);
nand U4868 (N_4868,In_130,In_488);
nand U4869 (N_4869,In_84,In_1824);
nor U4870 (N_4870,In_1717,In_2378);
nor U4871 (N_4871,In_1617,In_2010);
nor U4872 (N_4872,In_1201,In_848);
or U4873 (N_4873,In_352,In_558);
xnor U4874 (N_4874,In_419,In_420);
nand U4875 (N_4875,In_2273,In_2329);
and U4876 (N_4876,In_1857,In_1472);
xnor U4877 (N_4877,In_1625,In_1911);
or U4878 (N_4878,In_1801,In_1581);
and U4879 (N_4879,In_676,In_1795);
nand U4880 (N_4880,In_1182,In_1209);
nor U4881 (N_4881,In_2410,In_1325);
xor U4882 (N_4882,In_1471,In_264);
or U4883 (N_4883,In_244,In_909);
or U4884 (N_4884,In_2439,In_345);
or U4885 (N_4885,In_594,In_1705);
and U4886 (N_4886,In_903,In_1870);
nand U4887 (N_4887,In_567,In_1607);
nor U4888 (N_4888,In_1129,In_1092);
xor U4889 (N_4889,In_1483,In_459);
nand U4890 (N_4890,In_1668,In_2189);
or U4891 (N_4891,In_2126,In_876);
and U4892 (N_4892,In_3,In_1431);
or U4893 (N_4893,In_2092,In_2253);
xnor U4894 (N_4894,In_1151,In_1583);
and U4895 (N_4895,In_2173,In_2207);
or U4896 (N_4896,In_1752,In_347);
and U4897 (N_4897,In_2004,In_326);
xor U4898 (N_4898,In_764,In_894);
and U4899 (N_4899,In_658,In_2140);
nor U4900 (N_4900,In_1554,In_340);
xnor U4901 (N_4901,In_1701,In_1994);
nand U4902 (N_4902,In_1949,In_576);
xor U4903 (N_4903,In_671,In_1060);
nand U4904 (N_4904,In_56,In_968);
nand U4905 (N_4905,In_2447,In_298);
nand U4906 (N_4906,In_1150,In_389);
xor U4907 (N_4907,In_1852,In_931);
xnor U4908 (N_4908,In_2124,In_1398);
nor U4909 (N_4909,In_708,In_81);
or U4910 (N_4910,In_335,In_459);
nand U4911 (N_4911,In_1259,In_1081);
xor U4912 (N_4912,In_1126,In_2391);
nor U4913 (N_4913,In_2071,In_370);
and U4914 (N_4914,In_2072,In_1088);
nor U4915 (N_4915,In_65,In_1509);
xor U4916 (N_4916,In_211,In_21);
and U4917 (N_4917,In_297,In_2047);
xnor U4918 (N_4918,In_1367,In_394);
nor U4919 (N_4919,In_769,In_1338);
xnor U4920 (N_4920,In_1200,In_1766);
nor U4921 (N_4921,In_698,In_265);
or U4922 (N_4922,In_686,In_444);
or U4923 (N_4923,In_1443,In_2256);
nor U4924 (N_4924,In_2172,In_1865);
nand U4925 (N_4925,In_1570,In_427);
nand U4926 (N_4926,In_2337,In_817);
or U4927 (N_4927,In_1878,In_1869);
and U4928 (N_4928,In_12,In_1347);
nor U4929 (N_4929,In_1109,In_1865);
and U4930 (N_4930,In_1754,In_1037);
nand U4931 (N_4931,In_1867,In_1320);
xor U4932 (N_4932,In_977,In_2372);
nand U4933 (N_4933,In_220,In_1394);
or U4934 (N_4934,In_339,In_1946);
nor U4935 (N_4935,In_799,In_930);
nor U4936 (N_4936,In_267,In_1852);
nand U4937 (N_4937,In_2272,In_1855);
or U4938 (N_4938,In_2136,In_496);
or U4939 (N_4939,In_1113,In_767);
xor U4940 (N_4940,In_944,In_1049);
xor U4941 (N_4941,In_582,In_2234);
nand U4942 (N_4942,In_2379,In_150);
nor U4943 (N_4943,In_207,In_176);
or U4944 (N_4944,In_1014,In_1111);
nand U4945 (N_4945,In_704,In_1973);
or U4946 (N_4946,In_1604,In_237);
nor U4947 (N_4947,In_59,In_876);
xnor U4948 (N_4948,In_1868,In_1129);
xor U4949 (N_4949,In_716,In_1984);
nor U4950 (N_4950,In_2226,In_159);
or U4951 (N_4951,In_1298,In_1421);
nand U4952 (N_4952,In_1969,In_1737);
and U4953 (N_4953,In_536,In_1041);
and U4954 (N_4954,In_812,In_1793);
nor U4955 (N_4955,In_271,In_567);
xor U4956 (N_4956,In_1175,In_1880);
xnor U4957 (N_4957,In_2365,In_2316);
and U4958 (N_4958,In_960,In_2403);
or U4959 (N_4959,In_1611,In_2465);
xnor U4960 (N_4960,In_183,In_1852);
xnor U4961 (N_4961,In_107,In_1526);
nor U4962 (N_4962,In_50,In_1734);
nor U4963 (N_4963,In_2425,In_853);
nor U4964 (N_4964,In_1232,In_585);
or U4965 (N_4965,In_2288,In_1995);
xnor U4966 (N_4966,In_1226,In_1174);
nor U4967 (N_4967,In_195,In_631);
nand U4968 (N_4968,In_1420,In_2306);
or U4969 (N_4969,In_1479,In_1193);
nor U4970 (N_4970,In_1829,In_2054);
and U4971 (N_4971,In_1762,In_324);
xor U4972 (N_4972,In_1996,In_1680);
and U4973 (N_4973,In_153,In_38);
and U4974 (N_4974,In_649,In_1610);
and U4975 (N_4975,In_1510,In_1350);
xnor U4976 (N_4976,In_2118,In_1917);
nand U4977 (N_4977,In_1564,In_1781);
or U4978 (N_4978,In_1735,In_1852);
xor U4979 (N_4979,In_371,In_1042);
or U4980 (N_4980,In_233,In_2425);
xor U4981 (N_4981,In_672,In_2012);
or U4982 (N_4982,In_1478,In_364);
and U4983 (N_4983,In_541,In_1829);
xor U4984 (N_4984,In_413,In_1104);
xor U4985 (N_4985,In_1936,In_2032);
or U4986 (N_4986,In_2221,In_573);
xor U4987 (N_4987,In_1409,In_283);
xor U4988 (N_4988,In_2363,In_1641);
and U4989 (N_4989,In_855,In_634);
nand U4990 (N_4990,In_1103,In_1731);
xor U4991 (N_4991,In_1392,In_2468);
or U4992 (N_4992,In_1211,In_292);
nor U4993 (N_4993,In_1087,In_557);
xor U4994 (N_4994,In_1513,In_1811);
xnor U4995 (N_4995,In_175,In_1325);
and U4996 (N_4996,In_307,In_450);
nand U4997 (N_4997,In_1846,In_2134);
nor U4998 (N_4998,In_1108,In_2040);
nor U4999 (N_4999,In_2395,In_100);
xor U5000 (N_5000,N_3069,N_444);
xor U5001 (N_5001,N_4870,N_3520);
xor U5002 (N_5002,N_4951,N_2765);
or U5003 (N_5003,N_2267,N_4592);
xnor U5004 (N_5004,N_4890,N_2252);
and U5005 (N_5005,N_3212,N_2319);
and U5006 (N_5006,N_2174,N_2997);
xnor U5007 (N_5007,N_1007,N_461);
and U5008 (N_5008,N_4352,N_616);
xor U5009 (N_5009,N_349,N_4880);
nand U5010 (N_5010,N_1244,N_1422);
nand U5011 (N_5011,N_2354,N_4500);
xor U5012 (N_5012,N_669,N_4257);
and U5013 (N_5013,N_3716,N_2138);
nand U5014 (N_5014,N_582,N_2981);
nor U5015 (N_5015,N_1955,N_243);
and U5016 (N_5016,N_3454,N_1188);
xor U5017 (N_5017,N_3615,N_591);
xor U5018 (N_5018,N_1600,N_3917);
nand U5019 (N_5019,N_1277,N_4550);
xnor U5020 (N_5020,N_1642,N_3558);
nand U5021 (N_5021,N_318,N_3116);
and U5022 (N_5022,N_4864,N_4410);
xnor U5023 (N_5023,N_3852,N_4699);
and U5024 (N_5024,N_739,N_834);
nand U5025 (N_5025,N_3792,N_3576);
and U5026 (N_5026,N_4935,N_681);
nand U5027 (N_5027,N_4976,N_1827);
nand U5028 (N_5028,N_2651,N_4373);
and U5029 (N_5029,N_2240,N_965);
and U5030 (N_5030,N_76,N_4248);
nand U5031 (N_5031,N_1843,N_1591);
nand U5032 (N_5032,N_4797,N_813);
xnor U5033 (N_5033,N_1928,N_709);
xnor U5034 (N_5034,N_937,N_3431);
and U5035 (N_5035,N_3152,N_3952);
xnor U5036 (N_5036,N_915,N_2444);
nand U5037 (N_5037,N_4524,N_4288);
or U5038 (N_5038,N_116,N_4220);
and U5039 (N_5039,N_3401,N_3727);
nor U5040 (N_5040,N_4484,N_3875);
nor U5041 (N_5041,N_3166,N_209);
or U5042 (N_5042,N_1117,N_960);
nand U5043 (N_5043,N_377,N_245);
nand U5044 (N_5044,N_2735,N_2431);
nand U5045 (N_5045,N_3637,N_1572);
nand U5046 (N_5046,N_3430,N_3246);
xor U5047 (N_5047,N_3196,N_3713);
xnor U5048 (N_5048,N_3273,N_1593);
xnor U5049 (N_5049,N_4551,N_3377);
xnor U5050 (N_5050,N_2649,N_4185);
nor U5051 (N_5051,N_3386,N_2385);
and U5052 (N_5052,N_372,N_455);
nand U5053 (N_5053,N_3658,N_3493);
xnor U5054 (N_5054,N_2601,N_3410);
nor U5055 (N_5055,N_2030,N_3910);
and U5056 (N_5056,N_2464,N_1754);
or U5057 (N_5057,N_4121,N_1597);
and U5058 (N_5058,N_1525,N_1198);
and U5059 (N_5059,N_3075,N_1959);
nand U5060 (N_5060,N_1370,N_4584);
xnor U5061 (N_5061,N_430,N_495);
and U5062 (N_5062,N_2116,N_3800);
and U5063 (N_5063,N_2533,N_2375);
nor U5064 (N_5064,N_3328,N_4214);
and U5065 (N_5065,N_2245,N_376);
xor U5066 (N_5066,N_354,N_1087);
or U5067 (N_5067,N_4440,N_1866);
and U5068 (N_5068,N_358,N_4806);
nor U5069 (N_5069,N_4009,N_127);
and U5070 (N_5070,N_1564,N_3711);
nand U5071 (N_5071,N_4044,N_3770);
or U5072 (N_5072,N_605,N_1851);
nand U5073 (N_5073,N_2335,N_3543);
nand U5074 (N_5074,N_4741,N_3657);
nand U5075 (N_5075,N_744,N_2494);
or U5076 (N_5076,N_458,N_1510);
nand U5077 (N_5077,N_4777,N_1646);
nor U5078 (N_5078,N_440,N_4049);
nand U5079 (N_5079,N_2034,N_1448);
xor U5080 (N_5080,N_4832,N_687);
nand U5081 (N_5081,N_2092,N_1474);
xor U5082 (N_5082,N_4636,N_2785);
or U5083 (N_5083,N_1963,N_2280);
nor U5084 (N_5084,N_3214,N_2923);
nor U5085 (N_5085,N_1753,N_2455);
or U5086 (N_5086,N_1814,N_4126);
or U5087 (N_5087,N_1392,N_469);
xnor U5088 (N_5088,N_2855,N_4368);
xnor U5089 (N_5089,N_4385,N_2946);
or U5090 (N_5090,N_4293,N_3099);
or U5091 (N_5091,N_2578,N_4828);
nor U5092 (N_5092,N_2163,N_4161);
xnor U5093 (N_5093,N_2373,N_4125);
nand U5094 (N_5094,N_1307,N_147);
nor U5095 (N_5095,N_3754,N_2344);
or U5096 (N_5096,N_1423,N_1469);
xor U5097 (N_5097,N_3361,N_2986);
xnor U5098 (N_5098,N_713,N_4349);
nor U5099 (N_5099,N_1019,N_3913);
and U5100 (N_5100,N_2766,N_3843);
xnor U5101 (N_5101,N_2207,N_568);
nand U5102 (N_5102,N_4568,N_895);
and U5103 (N_5103,N_19,N_98);
xnor U5104 (N_5104,N_1042,N_53);
and U5105 (N_5105,N_1463,N_1693);
or U5106 (N_5106,N_4108,N_77);
xor U5107 (N_5107,N_660,N_2057);
nand U5108 (N_5108,N_3550,N_894);
or U5109 (N_5109,N_1943,N_4278);
nor U5110 (N_5110,N_4065,N_1082);
or U5111 (N_5111,N_3083,N_3086);
xnor U5112 (N_5112,N_1156,N_4781);
or U5113 (N_5113,N_909,N_1755);
and U5114 (N_5114,N_3975,N_722);
nor U5115 (N_5115,N_4234,N_2282);
and U5116 (N_5116,N_727,N_889);
nand U5117 (N_5117,N_4541,N_486);
or U5118 (N_5118,N_769,N_235);
nor U5119 (N_5119,N_317,N_1275);
nand U5120 (N_5120,N_2067,N_2586);
and U5121 (N_5121,N_3644,N_122);
or U5122 (N_5122,N_4256,N_3584);
nor U5123 (N_5123,N_143,N_899);
nand U5124 (N_5124,N_624,N_282);
xor U5125 (N_5125,N_4029,N_1992);
or U5126 (N_5126,N_1706,N_857);
and U5127 (N_5127,N_2691,N_1503);
nor U5128 (N_5128,N_2883,N_3502);
or U5129 (N_5129,N_2203,N_1450);
xor U5130 (N_5130,N_3516,N_2301);
nor U5131 (N_5131,N_4767,N_1142);
xnor U5132 (N_5132,N_1954,N_729);
and U5133 (N_5133,N_4355,N_4305);
or U5134 (N_5134,N_1923,N_389);
and U5135 (N_5135,N_4894,N_241);
and U5136 (N_5136,N_3753,N_3318);
xnor U5137 (N_5137,N_75,N_770);
or U5138 (N_5138,N_1530,N_2599);
nand U5139 (N_5139,N_916,N_2332);
or U5140 (N_5140,N_1739,N_2417);
or U5141 (N_5141,N_347,N_1934);
and U5142 (N_5142,N_1173,N_2291);
nand U5143 (N_5143,N_1653,N_580);
nor U5144 (N_5144,N_1080,N_386);
and U5145 (N_5145,N_18,N_2108);
or U5146 (N_5146,N_535,N_4237);
or U5147 (N_5147,N_2930,N_3158);
nor U5148 (N_5148,N_2739,N_184);
xor U5149 (N_5149,N_2210,N_2374);
xor U5150 (N_5150,N_4513,N_938);
and U5151 (N_5151,N_4332,N_3106);
xor U5152 (N_5152,N_4926,N_2906);
and U5153 (N_5153,N_180,N_1926);
and U5154 (N_5154,N_1489,N_82);
nor U5155 (N_5155,N_2638,N_3265);
nand U5156 (N_5156,N_4084,N_1581);
or U5157 (N_5157,N_1844,N_964);
nand U5158 (N_5158,N_2017,N_68);
xor U5159 (N_5159,N_3162,N_1339);
or U5160 (N_5160,N_3860,N_401);
nor U5161 (N_5161,N_974,N_3779);
nor U5162 (N_5162,N_485,N_4239);
nand U5163 (N_5163,N_3109,N_2672);
nand U5164 (N_5164,N_3927,N_1266);
nor U5165 (N_5165,N_3877,N_2758);
and U5166 (N_5166,N_4061,N_2061);
and U5167 (N_5167,N_3302,N_3521);
nor U5168 (N_5168,N_308,N_4936);
and U5169 (N_5169,N_1621,N_2682);
or U5170 (N_5170,N_3536,N_3900);
nor U5171 (N_5171,N_778,N_4981);
nor U5172 (N_5172,N_1768,N_2401);
nor U5173 (N_5173,N_92,N_1774);
and U5174 (N_5174,N_38,N_1598);
xnor U5175 (N_5175,N_2224,N_1273);
xnor U5176 (N_5176,N_3087,N_1004);
or U5177 (N_5177,N_4578,N_2933);
or U5178 (N_5178,N_1748,N_3908);
nand U5179 (N_5179,N_2737,N_2580);
or U5180 (N_5180,N_3478,N_784);
xor U5181 (N_5181,N_2802,N_3856);
or U5182 (N_5182,N_3971,N_4365);
or U5183 (N_5183,N_2716,N_3367);
nand U5184 (N_5184,N_4342,N_103);
and U5185 (N_5185,N_3280,N_3271);
and U5186 (N_5186,N_1967,N_1281);
xor U5187 (N_5187,N_357,N_2503);
nor U5188 (N_5188,N_4983,N_906);
nand U5189 (N_5189,N_3305,N_4988);
and U5190 (N_5190,N_3651,N_2629);
xor U5191 (N_5191,N_2306,N_4246);
and U5192 (N_5192,N_2890,N_4261);
nand U5193 (N_5193,N_8,N_4768);
or U5194 (N_5194,N_2979,N_2489);
and U5195 (N_5195,N_764,N_2775);
and U5196 (N_5196,N_2180,N_598);
xor U5197 (N_5197,N_1770,N_3032);
xor U5198 (N_5198,N_2162,N_3320);
and U5199 (N_5199,N_2956,N_3479);
nor U5200 (N_5200,N_866,N_3412);
or U5201 (N_5201,N_4778,N_1543);
or U5202 (N_5202,N_3055,N_4684);
nor U5203 (N_5203,N_2197,N_2110);
and U5204 (N_5204,N_2149,N_674);
nor U5205 (N_5205,N_572,N_2078);
and U5206 (N_5206,N_797,N_3031);
nand U5207 (N_5207,N_1038,N_2697);
nand U5208 (N_5208,N_396,N_206);
or U5209 (N_5209,N_4226,N_4640);
nand U5210 (N_5210,N_2005,N_99);
and U5211 (N_5211,N_3591,N_1028);
xnor U5212 (N_5212,N_3895,N_3552);
nand U5213 (N_5213,N_3326,N_1170);
nor U5214 (N_5214,N_4760,N_848);
nor U5215 (N_5215,N_4001,N_4526);
nor U5216 (N_5216,N_309,N_2103);
or U5217 (N_5217,N_11,N_3380);
xnor U5218 (N_5218,N_4804,N_3013);
or U5219 (N_5219,N_2394,N_904);
nand U5220 (N_5220,N_2941,N_635);
and U5221 (N_5221,N_721,N_2873);
or U5222 (N_5222,N_3924,N_2704);
nand U5223 (N_5223,N_2606,N_3732);
nor U5224 (N_5224,N_4851,N_699);
and U5225 (N_5225,N_749,N_4364);
nand U5226 (N_5226,N_2454,N_119);
nand U5227 (N_5227,N_10,N_1366);
or U5228 (N_5228,N_1268,N_1141);
or U5229 (N_5229,N_2463,N_4201);
xnor U5230 (N_5230,N_3681,N_1711);
xor U5231 (N_5231,N_1363,N_4522);
nand U5232 (N_5232,N_2475,N_1084);
and U5233 (N_5233,N_4409,N_4715);
nand U5234 (N_5234,N_4947,N_2688);
or U5235 (N_5235,N_4092,N_2683);
and U5236 (N_5236,N_4294,N_4112);
nor U5237 (N_5237,N_3,N_4518);
xnor U5238 (N_5238,N_1482,N_1295);
or U5239 (N_5239,N_205,N_1861);
or U5240 (N_5240,N_4077,N_4634);
xnor U5241 (N_5241,N_2963,N_1115);
or U5242 (N_5242,N_724,N_3472);
or U5243 (N_5243,N_4,N_972);
or U5244 (N_5244,N_384,N_3095);
xnor U5245 (N_5245,N_3457,N_4591);
xnor U5246 (N_5246,N_1476,N_4380);
xnor U5247 (N_5247,N_1394,N_4067);
and U5248 (N_5248,N_939,N_3553);
xnor U5249 (N_5249,N_753,N_4948);
and U5250 (N_5250,N_2769,N_4900);
xnor U5251 (N_5251,N_2850,N_4348);
and U5252 (N_5252,N_913,N_1574);
nand U5253 (N_5253,N_1998,N_2040);
or U5254 (N_5254,N_4339,N_1888);
nand U5255 (N_5255,N_1949,N_4235);
nand U5256 (N_5256,N_4224,N_4959);
nor U5257 (N_5257,N_2190,N_4018);
nand U5258 (N_5258,N_4456,N_1538);
nor U5259 (N_5259,N_4771,N_1267);
and U5260 (N_5260,N_168,N_3025);
nand U5261 (N_5261,N_4367,N_2857);
or U5262 (N_5262,N_3567,N_1900);
nor U5263 (N_5263,N_2294,N_824);
nand U5264 (N_5264,N_1415,N_3476);
nand U5265 (N_5265,N_1015,N_4765);
and U5266 (N_5266,N_1067,N_2339);
xor U5267 (N_5267,N_1622,N_2141);
nand U5268 (N_5268,N_2099,N_923);
or U5269 (N_5269,N_4898,N_3504);
nand U5270 (N_5270,N_4286,N_200);
xor U5271 (N_5271,N_3663,N_4530);
nor U5272 (N_5272,N_3486,N_1553);
nand U5273 (N_5273,N_3330,N_517);
nand U5274 (N_5274,N_4124,N_1668);
or U5275 (N_5275,N_167,N_3883);
nor U5276 (N_5276,N_3635,N_1131);
nor U5277 (N_5277,N_2673,N_2208);
or U5278 (N_5278,N_695,N_524);
and U5279 (N_5279,N_719,N_4712);
or U5280 (N_5280,N_299,N_2556);
xor U5281 (N_5281,N_1279,N_4128);
or U5282 (N_5282,N_3389,N_410);
nand U5283 (N_5283,N_422,N_4897);
nor U5284 (N_5284,N_3204,N_434);
and U5285 (N_5285,N_4709,N_2473);
xnor U5286 (N_5286,N_4388,N_2388);
nor U5287 (N_5287,N_3098,N_3861);
nor U5288 (N_5288,N_3721,N_3627);
or U5289 (N_5289,N_1696,N_1618);
and U5290 (N_5290,N_52,N_4917);
and U5291 (N_5291,N_2815,N_2939);
xor U5292 (N_5292,N_2699,N_3787);
nor U5293 (N_5293,N_4993,N_4282);
or U5294 (N_5294,N_4735,N_1335);
or U5295 (N_5295,N_2434,N_558);
nand U5296 (N_5296,N_3668,N_2485);
xnor U5297 (N_5297,N_4151,N_2701);
xor U5298 (N_5298,N_2383,N_3451);
xnor U5299 (N_5299,N_2367,N_3511);
nand U5300 (N_5300,N_1094,N_163);
nand U5301 (N_5301,N_13,N_4639);
nand U5302 (N_5302,N_2389,N_1807);
xnor U5303 (N_5303,N_4102,N_230);
nand U5304 (N_5304,N_1810,N_2700);
and U5305 (N_5305,N_1070,N_141);
and U5306 (N_5306,N_2405,N_2353);
nand U5307 (N_5307,N_3124,N_4865);
xnor U5308 (N_5308,N_651,N_1933);
or U5309 (N_5309,N_518,N_4701);
xnor U5310 (N_5310,N_1406,N_2725);
or U5311 (N_5311,N_4691,N_4274);
or U5312 (N_5312,N_946,N_1701);
nand U5313 (N_5313,N_4271,N_1132);
and U5314 (N_5314,N_2520,N_1662);
or U5315 (N_5315,N_1982,N_3400);
xnor U5316 (N_5316,N_4031,N_819);
nand U5317 (N_5317,N_686,N_1232);
xnor U5318 (N_5318,N_3030,N_584);
nor U5319 (N_5319,N_2171,N_1166);
nand U5320 (N_5320,N_2443,N_3755);
and U5321 (N_5321,N_3278,N_2396);
or U5322 (N_5322,N_2891,N_1317);
nand U5323 (N_5323,N_1932,N_4082);
and U5324 (N_5324,N_1672,N_144);
or U5325 (N_5325,N_4042,N_4775);
xor U5326 (N_5326,N_1913,N_1740);
or U5327 (N_5327,N_4310,N_4321);
and U5328 (N_5328,N_1439,N_4955);
nor U5329 (N_5329,N_66,N_818);
or U5330 (N_5330,N_601,N_777);
nor U5331 (N_5331,N_453,N_2729);
and U5332 (N_5332,N_1983,N_2973);
nand U5333 (N_5333,N_1729,N_3979);
xor U5334 (N_5334,N_4844,N_3091);
nor U5335 (N_5335,N_4670,N_706);
nand U5336 (N_5336,N_3348,N_1535);
and U5337 (N_5337,N_438,N_314);
or U5338 (N_5338,N_992,N_94);
nor U5339 (N_5339,N_1200,N_2772);
or U5340 (N_5340,N_3648,N_3827);
nor U5341 (N_5341,N_14,N_4437);
xnor U5342 (N_5342,N_3944,N_4602);
nand U5343 (N_5343,N_1342,N_1570);
nand U5344 (N_5344,N_1319,N_1425);
or U5345 (N_5345,N_4340,N_4991);
xnor U5346 (N_5346,N_4974,N_1429);
xnor U5347 (N_5347,N_3425,N_3596);
and U5348 (N_5348,N_4298,N_2472);
nor U5349 (N_5349,N_2880,N_4595);
and U5350 (N_5350,N_1210,N_4643);
or U5351 (N_5351,N_4879,N_3043);
nand U5352 (N_5352,N_383,N_1705);
or U5353 (N_5353,N_2840,N_711);
nand U5354 (N_5354,N_1234,N_4301);
nor U5355 (N_5355,N_647,N_1507);
nand U5356 (N_5356,N_4142,N_645);
xnor U5357 (N_5357,N_3948,N_3725);
xor U5358 (N_5358,N_489,N_4451);
nor U5359 (N_5359,N_3974,N_3394);
xor U5360 (N_5360,N_3081,N_158);
nor U5361 (N_5361,N_1956,N_2131);
nand U5362 (N_5362,N_9,N_3830);
nor U5363 (N_5363,N_61,N_3918);
or U5364 (N_5364,N_3020,N_2045);
and U5365 (N_5365,N_4876,N_2970);
and U5366 (N_5366,N_4064,N_3440);
and U5367 (N_5367,N_4626,N_3199);
nor U5368 (N_5368,N_771,N_216);
nand U5369 (N_5369,N_4136,N_126);
nor U5370 (N_5370,N_1731,N_828);
and U5371 (N_5371,N_4134,N_1787);
nand U5372 (N_5372,N_4496,N_4867);
nand U5373 (N_5373,N_4786,N_1346);
and U5374 (N_5374,N_2976,N_4040);
nor U5375 (N_5375,N_3808,N_407);
nor U5376 (N_5376,N_2242,N_233);
and U5377 (N_5377,N_4997,N_809);
nand U5378 (N_5378,N_213,N_1571);
or U5379 (N_5379,N_4381,N_2243);
nand U5380 (N_5380,N_302,N_931);
nand U5381 (N_5381,N_3832,N_3359);
nand U5382 (N_5382,N_4269,N_1251);
and U5383 (N_5383,N_2847,N_2988);
xnor U5384 (N_5384,N_4962,N_4430);
or U5385 (N_5385,N_2510,N_1182);
nand U5386 (N_5386,N_2290,N_3899);
nand U5387 (N_5387,N_1097,N_1874);
or U5388 (N_5388,N_653,N_3107);
xnor U5389 (N_5389,N_3463,N_2736);
or U5390 (N_5390,N_4180,N_3512);
or U5391 (N_5391,N_2093,N_2265);
xor U5392 (N_5392,N_4860,N_4395);
and U5393 (N_5393,N_4093,N_2286);
nor U5394 (N_5394,N_301,N_3513);
nor U5395 (N_5395,N_2756,N_28);
or U5396 (N_5396,N_297,N_2778);
or U5397 (N_5397,N_3064,N_4443);
and U5398 (N_5398,N_867,N_4869);
nor U5399 (N_5399,N_3569,N_4647);
nor U5400 (N_5400,N_2753,N_4529);
or U5401 (N_5401,N_187,N_173);
and U5402 (N_5402,N_3159,N_3173);
xnor U5403 (N_5403,N_3989,N_3560);
nor U5404 (N_5404,N_4507,N_732);
xnor U5405 (N_5405,N_4359,N_671);
and U5406 (N_5406,N_1402,N_3764);
nor U5407 (N_5407,N_2415,N_4555);
nand U5408 (N_5408,N_1821,N_3722);
and U5409 (N_5409,N_924,N_1472);
xor U5410 (N_5410,N_3052,N_63);
nand U5411 (N_5411,N_2300,N_3597);
xor U5412 (N_5412,N_3884,N_878);
xor U5413 (N_5413,N_3988,N_4280);
or U5414 (N_5414,N_1936,N_3660);
xor U5415 (N_5415,N_880,N_1792);
xnor U5416 (N_5416,N_312,N_3607);
and U5417 (N_5417,N_631,N_3531);
nand U5418 (N_5418,N_31,N_2898);
xor U5419 (N_5419,N_3855,N_123);
xor U5420 (N_5420,N_4710,N_1501);
xnor U5421 (N_5421,N_2193,N_1579);
nand U5422 (N_5422,N_4553,N_50);
and U5423 (N_5423,N_851,N_155);
xor U5424 (N_5424,N_4621,N_1318);
and U5425 (N_5425,N_1767,N_3969);
or U5426 (N_5426,N_1605,N_1678);
xnor U5427 (N_5427,N_519,N_3643);
or U5428 (N_5428,N_4776,N_4546);
nand U5429 (N_5429,N_1987,N_4004);
and U5430 (N_5430,N_1578,N_538);
and U5431 (N_5431,N_2878,N_4232);
nand U5432 (N_5432,N_1824,N_4360);
xnor U5433 (N_5433,N_3471,N_4027);
or U5434 (N_5434,N_3369,N_2184);
and U5435 (N_5435,N_4785,N_1111);
nor U5436 (N_5436,N_4115,N_4953);
or U5437 (N_5437,N_1663,N_4987);
and U5438 (N_5438,N_1059,N_1322);
nor U5439 (N_5439,N_2414,N_2044);
nor U5440 (N_5440,N_1609,N_3775);
and U5441 (N_5441,N_1099,N_2077);
xnor U5442 (N_5442,N_2094,N_1011);
or U5443 (N_5443,N_1620,N_4356);
or U5444 (N_5444,N_339,N_840);
nor U5445 (N_5445,N_1684,N_1452);
nand U5446 (N_5446,N_2271,N_1973);
xnor U5447 (N_5447,N_3114,N_3997);
nor U5448 (N_5448,N_2577,N_2948);
or U5449 (N_5449,N_3784,N_2176);
or U5450 (N_5450,N_788,N_4852);
and U5451 (N_5451,N_3903,N_3857);
xnor U5452 (N_5452,N_4399,N_1256);
or U5453 (N_5453,N_3227,N_2752);
or U5454 (N_5454,N_4230,N_1565);
nor U5455 (N_5455,N_4048,N_185);
nand U5456 (N_5456,N_883,N_190);
and U5457 (N_5457,N_2554,N_4449);
xor U5458 (N_5458,N_2380,N_3245);
or U5459 (N_5459,N_3379,N_3327);
and U5460 (N_5460,N_1387,N_2142);
nor U5461 (N_5461,N_3015,N_1758);
or U5462 (N_5462,N_1907,N_4014);
or U5463 (N_5463,N_1494,N_1459);
xnor U5464 (N_5464,N_2714,N_2655);
xor U5465 (N_5465,N_468,N_4868);
xnor U5466 (N_5466,N_4374,N_4651);
and U5467 (N_5467,N_4527,N_3845);
xor U5468 (N_5468,N_4160,N_4980);
xnor U5469 (N_5469,N_4941,N_4608);
nand U5470 (N_5470,N_2025,N_2812);
xnor U5471 (N_5471,N_1925,N_2555);
xnor U5472 (N_5472,N_569,N_553);
or U5473 (N_5473,N_3492,N_2524);
nor U5474 (N_5474,N_3272,N_1168);
nand U5475 (N_5475,N_4264,N_1610);
xor U5476 (N_5476,N_3695,N_1481);
xor U5477 (N_5477,N_3561,N_4107);
xor U5478 (N_5478,N_1927,N_2495);
and U5479 (N_5479,N_3949,N_3774);
and U5480 (N_5480,N_1899,N_661);
xor U5481 (N_5481,N_3276,N_2338);
nor U5482 (N_5482,N_1677,N_2079);
and U5483 (N_5483,N_1613,N_2476);
nand U5484 (N_5484,N_2258,N_3200);
or U5485 (N_5485,N_3940,N_2450);
xor U5486 (N_5486,N_4570,N_4521);
and U5487 (N_5487,N_4075,N_4925);
xnor U5488 (N_5488,N_2810,N_2813);
or U5489 (N_5489,N_702,N_4095);
and U5490 (N_5490,N_3142,N_390);
nand U5491 (N_5491,N_4087,N_4931);
nand U5492 (N_5492,N_2310,N_2945);
nand U5493 (N_5493,N_694,N_2496);
and U5494 (N_5494,N_1424,N_1098);
nor U5495 (N_5495,N_1833,N_1855);
xnor U5496 (N_5496,N_1180,N_4476);
and U5497 (N_5497,N_3128,N_836);
or U5498 (N_5498,N_27,N_1977);
xor U5499 (N_5499,N_1534,N_1588);
nor U5500 (N_5500,N_4158,N_2439);
xor U5501 (N_5501,N_1438,N_3983);
or U5502 (N_5502,N_991,N_2727);
and U5503 (N_5503,N_3718,N_3680);
nor U5504 (N_5504,N_2196,N_293);
nand U5505 (N_5505,N_3088,N_1981);
and U5506 (N_5506,N_4317,N_1941);
nand U5507 (N_5507,N_630,N_1030);
nor U5508 (N_5508,N_1154,N_3281);
nand U5509 (N_5509,N_1468,N_1327);
xnor U5510 (N_5510,N_3606,N_947);
nor U5511 (N_5511,N_4617,N_4453);
nand U5512 (N_5512,N_3218,N_2230);
nor U5513 (N_5513,N_2852,N_3191);
nor U5514 (N_5514,N_1831,N_2133);
xor U5515 (N_5515,N_3009,N_2333);
nor U5516 (N_5516,N_3869,N_846);
xor U5517 (N_5517,N_835,N_1779);
xnor U5518 (N_5518,N_4303,N_4861);
nand U5519 (N_5519,N_1435,N_2573);
and U5520 (N_5520,N_2486,N_3092);
nor U5521 (N_5521,N_4628,N_4078);
or U5522 (N_5522,N_211,N_2220);
nor U5523 (N_5523,N_4752,N_1694);
nor U5524 (N_5524,N_2340,N_1138);
nor U5525 (N_5525,N_2720,N_4164);
xnor U5526 (N_5526,N_4243,N_832);
nand U5527 (N_5527,N_1047,N_4069);
nor U5528 (N_5528,N_1911,N_1569);
and U5529 (N_5529,N_456,N_3448);
nor U5530 (N_5530,N_4604,N_4299);
nor U5531 (N_5531,N_3790,N_3223);
xor U5532 (N_5532,N_1576,N_2685);
nand U5533 (N_5533,N_3066,N_1383);
xor U5534 (N_5534,N_3057,N_3825);
nor U5535 (N_5535,N_4780,N_4163);
xor U5536 (N_5536,N_201,N_1430);
or U5537 (N_5537,N_648,N_839);
and U5538 (N_5538,N_531,N_3118);
and U5539 (N_5539,N_1276,N_1040);
and U5540 (N_5540,N_1842,N_3554);
or U5541 (N_5541,N_3794,N_513);
nand U5542 (N_5542,N_1355,N_4404);
and U5543 (N_5543,N_984,N_4319);
and U5544 (N_5544,N_3195,N_3548);
and U5545 (N_5545,N_969,N_1968);
and U5546 (N_5546,N_1944,N_4464);
or U5547 (N_5547,N_1718,N_3700);
nor U5548 (N_5548,N_3639,N_4450);
xor U5549 (N_5549,N_4896,N_1069);
nand U5550 (N_5550,N_2407,N_1896);
or U5551 (N_5551,N_4086,N_3368);
or U5552 (N_5552,N_3203,N_4291);
and U5553 (N_5553,N_3583,N_4229);
and U5554 (N_5554,N_2001,N_525);
xnor U5555 (N_5555,N_2867,N_1114);
xor U5556 (N_5556,N_1398,N_1749);
and U5557 (N_5557,N_505,N_1879);
nor U5558 (N_5558,N_161,N_504);
nand U5559 (N_5559,N_3004,N_2920);
or U5560 (N_5560,N_4267,N_4135);
nand U5561 (N_5561,N_798,N_2853);
or U5562 (N_5562,N_1024,N_3491);
and U5563 (N_5563,N_2304,N_3252);
xnor U5564 (N_5564,N_3450,N_2546);
or U5565 (N_5565,N_4739,N_2166);
nor U5566 (N_5566,N_1730,N_3117);
and U5567 (N_5567,N_4207,N_1895);
xnor U5568 (N_5568,N_2349,N_4596);
nor U5569 (N_5569,N_2119,N_1940);
nor U5570 (N_5570,N_2014,N_4292);
xnor U5571 (N_5571,N_4169,N_2442);
nand U5572 (N_5572,N_1785,N_3810);
nor U5573 (N_5573,N_789,N_4520);
or U5574 (N_5574,N_2154,N_1136);
xor U5575 (N_5575,N_3964,N_3547);
xnor U5576 (N_5576,N_4782,N_3858);
nand U5577 (N_5577,N_2378,N_641);
xnor U5578 (N_5578,N_4788,N_313);
nand U5579 (N_5579,N_4968,N_1736);
or U5580 (N_5580,N_2026,N_2734);
or U5581 (N_5581,N_4079,N_2188);
xnor U5582 (N_5582,N_1492,N_4688);
xnor U5583 (N_5583,N_1630,N_4800);
xnor U5584 (N_5584,N_4627,N_2278);
xnor U5585 (N_5585,N_4912,N_2363);
and U5586 (N_5586,N_2113,N_714);
nand U5587 (N_5587,N_2132,N_1191);
and U5588 (N_5588,N_608,N_2090);
or U5589 (N_5589,N_487,N_2185);
nor U5590 (N_5590,N_2816,N_81);
xnor U5591 (N_5591,N_1344,N_3846);
nor U5592 (N_5592,N_2515,N_1560);
nand U5593 (N_5593,N_2246,N_1629);
or U5594 (N_5594,N_4732,N_4964);
and U5595 (N_5595,N_3357,N_3709);
xor U5596 (N_5596,N_1129,N_4052);
or U5597 (N_5597,N_4714,N_4693);
nor U5598 (N_5598,N_4311,N_2052);
or U5599 (N_5599,N_3160,N_2901);
and U5600 (N_5600,N_2613,N_327);
nand U5601 (N_5601,N_1829,N_4244);
nand U5602 (N_5602,N_4790,N_4652);
or U5603 (N_5603,N_4233,N_2312);
or U5604 (N_5604,N_4891,N_3115);
xor U5605 (N_5605,N_3541,N_994);
nor U5606 (N_5606,N_2957,N_1032);
or U5607 (N_5607,N_4548,N_2070);
nor U5608 (N_5608,N_676,N_4645);
nor U5609 (N_5609,N_3164,N_3889);
xor U5610 (N_5610,N_655,N_4028);
or U5611 (N_5611,N_397,N_4393);
nor U5612 (N_5612,N_640,N_4287);
and U5613 (N_5613,N_3529,N_3815);
or U5614 (N_5614,N_3094,N_1382);
or U5615 (N_5615,N_290,N_2865);
or U5616 (N_5616,N_4966,N_4493);
nor U5617 (N_5617,N_3838,N_737);
xor U5618 (N_5618,N_1633,N_1409);
and U5619 (N_5619,N_3482,N_2732);
xnor U5620 (N_5620,N_4644,N_4460);
xnor U5621 (N_5621,N_3300,N_2616);
and U5622 (N_5622,N_820,N_1471);
and U5623 (N_5623,N_3676,N_1635);
nor U5624 (N_5624,N_4198,N_3498);
nand U5625 (N_5625,N_2307,N_421);
xor U5626 (N_5626,N_2547,N_196);
or U5627 (N_5627,N_1513,N_3414);
and U5628 (N_5628,N_2708,N_3866);
xor U5629 (N_5629,N_898,N_3747);
xnor U5630 (N_5630,N_4885,N_4187);
and U5631 (N_5631,N_2391,N_507);
and U5632 (N_5632,N_3277,N_2531);
or U5633 (N_5633,N_4620,N_1852);
nand U5634 (N_5634,N_4759,N_137);
or U5635 (N_5635,N_3586,N_466);
and U5636 (N_5636,N_445,N_223);
nand U5637 (N_5637,N_4692,N_2421);
and U5638 (N_5638,N_3003,N_106);
and U5639 (N_5639,N_4698,N_3629);
xnor U5640 (N_5640,N_166,N_2127);
xor U5641 (N_5641,N_1286,N_1083);
nand U5642 (N_5642,N_4315,N_1766);
and U5643 (N_5643,N_1615,N_716);
and U5644 (N_5644,N_4727,N_2798);
nand U5645 (N_5645,N_3082,N_1808);
or U5646 (N_5646,N_1385,N_2565);
xor U5647 (N_5647,N_1876,N_3694);
nor U5648 (N_5648,N_1163,N_4725);
nor U5649 (N_5649,N_4354,N_2365);
nand U5650 (N_5650,N_2501,N_45);
and U5651 (N_5651,N_1143,N_4300);
xor U5652 (N_5652,N_4946,N_2861);
nor U5653 (N_5653,N_2399,N_928);
nand U5654 (N_5654,N_1433,N_2347);
or U5655 (N_5655,N_4819,N_2804);
or U5656 (N_5656,N_4401,N_1947);
nand U5657 (N_5657,N_2549,N_4706);
xor U5658 (N_5658,N_462,N_3210);
nand U5659 (N_5659,N_3955,N_3939);
and U5660 (N_5660,N_412,N_2967);
nand U5661 (N_5661,N_4007,N_1826);
nand U5662 (N_5662,N_2172,N_3021);
nor U5663 (N_5663,N_4313,N_2006);
nor U5664 (N_5664,N_1887,N_2669);
nand U5665 (N_5665,N_3331,N_1797);
nand U5666 (N_5666,N_807,N_2075);
or U5667 (N_5667,N_4749,N_2771);
nor U5668 (N_5668,N_3972,N_32);
nand U5669 (N_5669,N_3444,N_2257);
and U5670 (N_5670,N_1676,N_2530);
or U5671 (N_5671,N_3911,N_2218);
nor U5672 (N_5672,N_2974,N_1348);
or U5673 (N_5673,N_224,N_3748);
or U5674 (N_5674,N_1147,N_4182);
nor U5675 (N_5675,N_4433,N_4967);
or U5676 (N_5676,N_1857,N_4024);
nand U5677 (N_5677,N_3434,N_2938);
xnor U5678 (N_5678,N_2059,N_4942);
and U5679 (N_5679,N_1195,N_436);
nor U5680 (N_5680,N_217,N_3008);
or U5681 (N_5681,N_3060,N_1938);
and U5682 (N_5682,N_3294,N_2671);
or U5683 (N_5683,N_882,N_4754);
xnor U5684 (N_5684,N_2478,N_3891);
xor U5685 (N_5685,N_2591,N_1413);
nor U5686 (N_5686,N_4502,N_2317);
nor U5687 (N_5687,N_665,N_4116);
nor U5688 (N_5688,N_2567,N_348);
or U5689 (N_5689,N_3175,N_408);
and U5690 (N_5690,N_1243,N_3984);
nand U5691 (N_5691,N_2177,N_4787);
and U5692 (N_5692,N_3198,N_2437);
and U5693 (N_5693,N_1049,N_1648);
nor U5694 (N_5694,N_3180,N_4255);
and U5695 (N_5695,N_2991,N_4051);
or U5696 (N_5696,N_4632,N_1839);
and U5697 (N_5697,N_1838,N_1643);
or U5698 (N_5698,N_4272,N_2398);
and U5699 (N_5699,N_890,N_2235);
or U5700 (N_5700,N_1884,N_4369);
nand U5701 (N_5701,N_403,N_1009);
and U5702 (N_5702,N_2821,N_945);
and U5703 (N_5703,N_494,N_4718);
or U5704 (N_5704,N_3590,N_343);
and U5705 (N_5705,N_2703,N_4970);
or U5706 (N_5706,N_4724,N_2889);
nor U5707 (N_5707,N_2448,N_2803);
nand U5708 (N_5708,N_1966,N_1850);
nor U5709 (N_5709,N_3915,N_2035);
or U5710 (N_5710,N_3679,N_4677);
nor U5711 (N_5711,N_1972,N_1551);
xnor U5712 (N_5712,N_4571,N_4002);
nor U5713 (N_5713,N_2912,N_2227);
or U5714 (N_5714,N_2424,N_1502);
xnor U5715 (N_5715,N_4512,N_973);
xor U5716 (N_5716,N_1769,N_3634);
or U5717 (N_5717,N_4683,N_1377);
nor U5718 (N_5718,N_3496,N_3682);
nand U5719 (N_5719,N_43,N_2273);
xnor U5720 (N_5720,N_3638,N_4515);
xor U5721 (N_5721,N_2940,N_340);
or U5722 (N_5722,N_4445,N_2170);
and U5723 (N_5723,N_3065,N_3363);
or U5724 (N_5724,N_4238,N_4899);
nand U5725 (N_5725,N_578,N_884);
nand U5726 (N_5726,N_4793,N_2470);
nor U5727 (N_5727,N_4217,N_4689);
nor U5728 (N_5728,N_464,N_160);
and U5729 (N_5729,N_1149,N_1284);
xor U5730 (N_5730,N_1061,N_4285);
and U5731 (N_5731,N_1695,N_892);
xor U5732 (N_5732,N_1003,N_3112);
nor U5733 (N_5733,N_3799,N_1691);
or U5734 (N_5734,N_656,N_179);
and U5735 (N_5735,N_4610,N_2153);
xor U5736 (N_5736,N_2611,N_1403);
and U5737 (N_5737,N_2666,N_298);
nor U5738 (N_5738,N_3288,N_474);
xor U5739 (N_5739,N_4707,N_3620);
or U5740 (N_5740,N_3452,N_3295);
or U5741 (N_5741,N_988,N_3260);
nand U5742 (N_5742,N_1703,N_3206);
nand U5743 (N_5743,N_4114,N_1760);
nand U5744 (N_5744,N_4019,N_4603);
xor U5745 (N_5745,N_2283,N_1257);
or U5746 (N_5746,N_467,N_4810);
nand U5747 (N_5747,N_4492,N_3613);
or U5748 (N_5748,N_514,N_277);
and U5749 (N_5749,N_3585,N_3514);
nand U5750 (N_5750,N_1179,N_1153);
nand U5751 (N_5751,N_3556,N_2481);
nand U5752 (N_5752,N_2817,N_3678);
xnor U5753 (N_5753,N_1443,N_952);
and U5754 (N_5754,N_2334,N_1063);
xnor U5755 (N_5755,N_2647,N_1637);
nand U5756 (N_5756,N_1208,N_2710);
xnor U5757 (N_5757,N_4196,N_4184);
or U5758 (N_5758,N_4062,N_515);
nand U5759 (N_5759,N_1465,N_4432);
or U5760 (N_5760,N_4744,N_93);
nand U5761 (N_5761,N_691,N_3104);
nand U5762 (N_5762,N_599,N_2028);
and U5763 (N_5763,N_1230,N_252);
xnor U5764 (N_5764,N_3821,N_3959);
nand U5765 (N_5765,N_3742,N_4103);
or U5766 (N_5766,N_3795,N_3659);
and U5767 (N_5767,N_2728,N_955);
xnor U5768 (N_5768,N_3738,N_3089);
nor U5769 (N_5769,N_1835,N_1121);
xnor U5770 (N_5770,N_1066,N_3938);
nand U5771 (N_5771,N_1556,N_2897);
and U5772 (N_5772,N_322,N_618);
xnor U5773 (N_5773,N_4309,N_3691);
xor U5774 (N_5774,N_1848,N_3572);
or U5775 (N_5775,N_2293,N_2095);
nand U5776 (N_5776,N_3618,N_879);
nand U5777 (N_5777,N_2509,N_4909);
nand U5778 (N_5778,N_2882,N_3143);
nand U5779 (N_5779,N_2147,N_419);
and U5780 (N_5780,N_1796,N_1008);
xnor U5781 (N_5781,N_4989,N_1428);
and U5782 (N_5782,N_560,N_1898);
or U5783 (N_5783,N_3985,N_3667);
and U5784 (N_5784,N_2858,N_833);
nor U5785 (N_5785,N_4576,N_3608);
nor U5786 (N_5786,N_2302,N_2659);
and U5787 (N_5787,N_1240,N_2091);
nand U5788 (N_5788,N_3370,N_547);
or U5789 (N_5789,N_3720,N_1367);
or U5790 (N_5790,N_286,N_3423);
xnor U5791 (N_5791,N_415,N_4215);
or U5792 (N_5792,N_2796,N_956);
nand U5793 (N_5793,N_2837,N_452);
or U5794 (N_5794,N_1986,N_1112);
or U5795 (N_5795,N_1636,N_842);
xor U5796 (N_5796,N_3517,N_2750);
nor U5797 (N_5797,N_776,N_3796);
nor U5798 (N_5798,N_2461,N_3238);
or U5799 (N_5799,N_4803,N_1820);
nor U5800 (N_5800,N_3253,N_3282);
nand U5801 (N_5801,N_420,N_3188);
nand U5802 (N_5802,N_2051,N_1738);
nor U5803 (N_5803,N_1679,N_1397);
xnor U5804 (N_5804,N_4347,N_2919);
and U5805 (N_5805,N_90,N_2870);
nand U5806 (N_5806,N_2745,N_2325);
nand U5807 (N_5807,N_484,N_2042);
nor U5808 (N_5808,N_3483,N_743);
or U5809 (N_5809,N_2994,N_1667);
xor U5810 (N_5810,N_3982,N_295);
nand U5811 (N_5811,N_250,N_424);
and U5812 (N_5812,N_4660,N_926);
and U5813 (N_5813,N_1227,N_1076);
xor U5814 (N_5814,N_2839,N_3500);
and U5815 (N_5815,N_4036,N_4045);
nor U5816 (N_5816,N_74,N_404);
nand U5817 (N_5817,N_3374,N_2846);
and U5818 (N_5818,N_23,N_2887);
nand U5819 (N_5819,N_1700,N_47);
nand U5820 (N_5820,N_3242,N_2978);
nor U5821 (N_5821,N_4442,N_1717);
or U5822 (N_5822,N_2996,N_2575);
and U5823 (N_5823,N_3063,N_1119);
nand U5824 (N_5824,N_1483,N_237);
xor U5825 (N_5825,N_3497,N_2689);
or U5826 (N_5826,N_1144,N_1157);
nor U5827 (N_5827,N_3565,N_3693);
xnor U5828 (N_5828,N_4081,N_2326);
or U5829 (N_5829,N_682,N_948);
or U5830 (N_5830,N_765,N_1336);
nor U5831 (N_5831,N_2198,N_2249);
or U5832 (N_5832,N_670,N_1549);
and U5833 (N_5833,N_2781,N_3197);
nand U5834 (N_5834,N_521,N_3044);
or U5835 (N_5835,N_4037,N_2977);
nor U5836 (N_5836,N_3465,N_814);
nand U5837 (N_5837,N_4862,N_3862);
nor U5838 (N_5838,N_4809,N_2292);
xor U5839 (N_5839,N_5,N_2763);
nand U5840 (N_5840,N_3446,N_1477);
and U5841 (N_5841,N_4454,N_3714);
xor U5842 (N_5842,N_289,N_3251);
or U5843 (N_5843,N_379,N_957);
or U5844 (N_5844,N_1939,N_2041);
and U5845 (N_5845,N_1690,N_3907);
or U5846 (N_5846,N_3781,N_3669);
or U5847 (N_5847,N_3387,N_1640);
xor U5848 (N_5848,N_845,N_2024);
or U5849 (N_5849,N_3022,N_4503);
xnor U5850 (N_5850,N_4886,N_4874);
xor U5851 (N_5851,N_1021,N_4770);
nand U5852 (N_5852,N_374,N_3067);
nor U5853 (N_5853,N_2592,N_3602);
xnor U5854 (N_5854,N_557,N_4648);
xnor U5855 (N_5855,N_72,N_3731);
nor U5856 (N_5856,N_4999,N_4969);
or U5857 (N_5857,N_306,N_326);
or U5858 (N_5858,N_4200,N_3710);
nor U5859 (N_5859,N_1488,N_4438);
and U5860 (N_5860,N_2420,N_275);
xor U5861 (N_5861,N_971,N_3892);
and U5862 (N_5862,N_3261,N_287);
xor U5863 (N_5863,N_1892,N_3257);
xnor U5864 (N_5864,N_1665,N_181);
nor U5865 (N_5865,N_3090,N_4954);
nor U5866 (N_5866,N_2086,N_1071);
nand U5867 (N_5867,N_612,N_4297);
nand U5868 (N_5868,N_4562,N_2126);
nor U5869 (N_5869,N_78,N_1715);
xnor U5870 (N_5870,N_3728,N_4758);
and U5871 (N_5871,N_4854,N_3371);
nand U5872 (N_5872,N_3375,N_1133);
and U5873 (N_5873,N_4378,N_271);
xor U5874 (N_5874,N_4537,N_2003);
xnor U5875 (N_5875,N_3923,N_270);
and U5876 (N_5876,N_4016,N_1937);
nor U5877 (N_5877,N_4730,N_4420);
xnor U5878 (N_5878,N_2779,N_3051);
and U5879 (N_5879,N_2289,N_3244);
nand U5880 (N_5880,N_4212,N_3134);
nand U5881 (N_5881,N_1041,N_2260);
or U5882 (N_5882,N_2854,N_3666);
nand U5883 (N_5883,N_869,N_4318);
and U5884 (N_5884,N_1490,N_3580);
and U5885 (N_5885,N_3555,N_3987);
or U5886 (N_5886,N_4379,N_983);
or U5887 (N_5887,N_2106,N_3791);
and U5888 (N_5888,N_1611,N_332);
and U5889 (N_5889,N_4875,N_2268);
nand U5890 (N_5890,N_1803,N_4605);
nand U5891 (N_5891,N_2377,N_1374);
nor U5892 (N_5892,N_4871,N_400);
or U5893 (N_5893,N_2859,N_4769);
or U5894 (N_5894,N_3937,N_3168);
and U5895 (N_5895,N_2557,N_442);
nand U5896 (N_5896,N_1199,N_981);
xnor U5897 (N_5897,N_2722,N_1645);
or U5898 (N_5898,N_1673,N_3100);
xnor U5899 (N_5899,N_431,N_1316);
or U5900 (N_5900,N_3193,N_1401);
nand U5901 (N_5901,N_3393,N_3750);
nand U5902 (N_5902,N_2010,N_1224);
nand U5903 (N_5903,N_1301,N_805);
nor U5904 (N_5904,N_280,N_2830);
nor U5905 (N_5905,N_2724,N_4325);
or U5906 (N_5906,N_901,N_3865);
or U5907 (N_5907,N_549,N_1324);
nor U5908 (N_5908,N_2004,N_4704);
nor U5909 (N_5909,N_3213,N_1356);
or U5910 (N_5910,N_4441,N_2950);
or U5911 (N_5911,N_1096,N_1751);
nor U5912 (N_5912,N_4855,N_662);
nor U5913 (N_5913,N_3935,N_790);
nor U5914 (N_5914,N_1546,N_3932);
nand U5915 (N_5915,N_4446,N_1444);
nor U5916 (N_5916,N_4462,N_3705);
nor U5917 (N_5917,N_3594,N_920);
nor U5918 (N_5918,N_4511,N_4371);
or U5919 (N_5919,N_4162,N_3167);
and U5920 (N_5920,N_2021,N_174);
nand U5921 (N_5921,N_2213,N_980);
or U5922 (N_5922,N_1997,N_3157);
nor U5923 (N_5923,N_3980,N_1446);
and U5924 (N_5924,N_506,N_1177);
xor U5925 (N_5925,N_1809,N_896);
or U5926 (N_5926,N_1592,N_4783);
nor U5927 (N_5927,N_1437,N_2605);
xnor U5928 (N_5928,N_718,N_2983);
nand U5929 (N_5929,N_4129,N_2872);
and U5930 (N_5930,N_1235,N_2844);
and U5931 (N_5931,N_266,N_2820);
and U5932 (N_5932,N_4375,N_592);
or U5933 (N_5933,N_265,N_4296);
xor U5934 (N_5934,N_4856,N_646);
xor U5935 (N_5935,N_3391,N_2355);
nor U5936 (N_5936,N_847,N_4487);
and U5937 (N_5937,N_2914,N_875);
nand U5938 (N_5938,N_4060,N_1293);
and U5939 (N_5939,N_2000,N_567);
nand U5940 (N_5940,N_496,N_720);
and U5941 (N_5941,N_3546,N_1719);
nor U5942 (N_5942,N_2916,N_4322);
and U5943 (N_5943,N_540,N_4950);
nor U5944 (N_5944,N_4973,N_2838);
or U5945 (N_5945,N_3998,N_80);
or U5946 (N_5946,N_2343,N_3187);
nand U5947 (N_5947,N_2358,N_2877);
xnor U5948 (N_5948,N_588,N_2780);
or U5949 (N_5949,N_3631,N_316);
xor U5950 (N_5950,N_1453,N_1311);
xnor U5951 (N_5951,N_1671,N_4582);
or U5952 (N_5952,N_2899,N_4618);
or U5953 (N_5953,N_2248,N_4463);
nor U5954 (N_5954,N_3462,N_2845);
nand U5955 (N_5955,N_3352,N_2369);
xor U5956 (N_5956,N_4335,N_1455);
and U5957 (N_5957,N_1819,N_1847);
xnor U5958 (N_5958,N_949,N_2783);
and U5959 (N_5959,N_4559,N_2526);
nor U5960 (N_5960,N_4117,N_4831);
and U5961 (N_5961,N_1350,N_3426);
and U5962 (N_5962,N_2490,N_2428);
and U5963 (N_5963,N_2123,N_2137);
or U5964 (N_5964,N_2504,N_4405);
nand U5965 (N_5965,N_3963,N_2308);
nor U5966 (N_5966,N_2905,N_2359);
nor U5967 (N_5967,N_1707,N_1205);
xor U5968 (N_5968,N_4205,N_3871);
or U5969 (N_5969,N_3147,N_3490);
and U5970 (N_5970,N_1890,N_863);
nor U5971 (N_5971,N_1487,N_4022);
nand U5972 (N_5972,N_4138,N_3687);
and U5973 (N_5973,N_1903,N_1841);
or U5974 (N_5974,N_4774,N_2516);
nand U5975 (N_5975,N_860,N_4560);
xor U5976 (N_5976,N_4005,N_4473);
xor U5977 (N_5977,N_3074,N_2623);
nand U5978 (N_5978,N_1650,N_378);
or U5979 (N_5979,N_4904,N_2048);
xnor U5980 (N_5980,N_689,N_3205);
and U5981 (N_5981,N_1536,N_3045);
or U5982 (N_5982,N_263,N_1791);
nor U5983 (N_5983,N_2517,N_3418);
nand U5984 (N_5984,N_2453,N_4025);
and U5985 (N_5985,N_4872,N_3145);
nand U5986 (N_5986,N_3535,N_940);
and U5987 (N_5987,N_2219,N_2071);
or U5988 (N_5988,N_2645,N_1440);
nand U5989 (N_5989,N_652,N_954);
nor U5990 (N_5990,N_3007,N_79);
or U5991 (N_5991,N_3316,N_4431);
xor U5992 (N_5992,N_3925,N_3306);
or U5993 (N_5993,N_3507,N_4304);
or U5994 (N_5994,N_725,N_222);
and U5995 (N_5995,N_3729,N_4594);
xnor U5996 (N_5996,N_338,N_2811);
nor U5997 (N_5997,N_1562,N_446);
xnor U5998 (N_5998,N_4960,N_4480);
nor U5999 (N_5999,N_2896,N_4895);
or U6000 (N_6000,N_4572,N_406);
or U6001 (N_6001,N_4396,N_2926);
and U6002 (N_6002,N_2955,N_1405);
and U6003 (N_6003,N_3802,N_2707);
or U6004 (N_6004,N_3208,N_4588);
or U6005 (N_6005,N_2712,N_510);
or U6006 (N_6006,N_324,N_2426);
nor U6007 (N_6007,N_1822,N_865);
xnor U6008 (N_6008,N_4144,N_4873);
xnor U6009 (N_6009,N_3125,N_2563);
and U6010 (N_6010,N_1916,N_571);
nor U6011 (N_6011,N_1805,N_3103);
xor U6012 (N_6012,N_3445,N_1798);
nand U6013 (N_6013,N_1126,N_1457);
or U6014 (N_6014,N_2085,N_2346);
or U6015 (N_6015,N_3850,N_3309);
and U6016 (N_6016,N_2545,N_4376);
and U6017 (N_6017,N_2871,N_2357);
and U6018 (N_6018,N_3751,N_3934);
or U6019 (N_6019,N_3050,N_191);
or U6020 (N_6020,N_3803,N_199);
nor U6021 (N_6021,N_4035,N_2161);
nand U6022 (N_6022,N_4893,N_3464);
nor U6023 (N_6023,N_276,N_2733);
xnor U6024 (N_6024,N_1416,N_2929);
or U6025 (N_6025,N_4932,N_3780);
nand U6026 (N_6026,N_1589,N_4833);
or U6027 (N_6027,N_4362,N_1155);
nor U6028 (N_6028,N_26,N_2255);
nand U6029 (N_6029,N_1960,N_2937);
nor U6030 (N_6030,N_334,N_2382);
or U6031 (N_6031,N_2337,N_4384);
nand U6032 (N_6032,N_543,N_1325);
or U6033 (N_6033,N_49,N_2522);
xnor U6034 (N_6034,N_4653,N_4343);
nor U6035 (N_6035,N_3035,N_2596);
or U6036 (N_6036,N_3181,N_3275);
xor U6037 (N_6037,N_4242,N_3723);
and U6038 (N_6038,N_1520,N_856);
or U6039 (N_6039,N_2951,N_1456);
nor U6040 (N_6040,N_4723,N_3477);
or U6041 (N_6041,N_2570,N_4137);
xnor U6042 (N_6042,N_249,N_2323);
nand U6043 (N_6043,N_2222,N_528);
and U6044 (N_6044,N_4930,N_3042);
and U6045 (N_6045,N_470,N_2251);
nand U6046 (N_6046,N_4150,N_1220);
xor U6047 (N_6047,N_1984,N_2425);
xnor U6048 (N_6048,N_3028,N_4083);
and U6049 (N_6049,N_1441,N_811);
or U6050 (N_6050,N_4649,N_808);
or U6051 (N_6051,N_4377,N_156);
xor U6052 (N_6052,N_1818,N_1419);
nand U6053 (N_6053,N_4063,N_3698);
or U6054 (N_6054,N_2462,N_600);
or U6055 (N_6055,N_335,N_1005);
and U6056 (N_6056,N_4351,N_876);
xnor U6057 (N_6057,N_3149,N_4549);
nor U6058 (N_6058,N_3376,N_4837);
nand U6059 (N_6059,N_3353,N_195);
xnor U6060 (N_6060,N_4817,N_333);
nand U6061 (N_6061,N_2656,N_2422);
nor U6062 (N_6062,N_2773,N_1287);
nand U6063 (N_6063,N_3820,N_2427);
and U6064 (N_6064,N_1832,N_4091);
or U6065 (N_6065,N_291,N_1623);
xor U6066 (N_6066,N_2642,N_636);
nand U6067 (N_6067,N_3922,N_2836);
nand U6068 (N_6068,N_1054,N_188);
and U6069 (N_6069,N_2612,N_3532);
nor U6070 (N_6070,N_2824,N_2136);
nand U6071 (N_6071,N_1122,N_583);
or U6072 (N_6072,N_2403,N_3217);
or U6073 (N_6073,N_4099,N_3140);
xor U6074 (N_6074,N_3837,N_17);
xnor U6075 (N_6075,N_4581,N_1603);
nand U6076 (N_6076,N_4331,N_1023);
or U6077 (N_6077,N_2316,N_3416);
nand U6078 (N_6078,N_4307,N_3809);
nand U6079 (N_6079,N_1343,N_1055);
xnor U6080 (N_6080,N_473,N_1771);
xor U6081 (N_6081,N_607,N_3381);
or U6082 (N_6082,N_2990,N_2789);
nor U6083 (N_6083,N_2759,N_4849);
and U6084 (N_6084,N_3262,N_1442);
and U6085 (N_6085,N_288,N_2564);
nor U6086 (N_6086,N_4662,N_2762);
or U6087 (N_6087,N_2390,N_1599);
nor U6088 (N_6088,N_2541,N_1371);
nor U6089 (N_6089,N_1511,N_3818);
nand U6090 (N_6090,N_4853,N_703);
or U6091 (N_6091,N_4505,N_488);
xnor U6092 (N_6092,N_2600,N_4003);
nor U6093 (N_6093,N_4514,N_2921);
and U6094 (N_6094,N_104,N_4344);
xnor U6095 (N_6095,N_2191,N_2971);
and U6096 (N_6096,N_3957,N_4398);
nand U6097 (N_6097,N_4746,N_2114);
nand U6098 (N_6098,N_2639,N_3105);
and U6099 (N_6099,N_3902,N_2418);
nand U6100 (N_6100,N_2211,N_3898);
nor U6101 (N_6101,N_2791,N_2801);
xnor U6102 (N_6102,N_4789,N_1309);
nor U6103 (N_6103,N_548,N_4017);
xnor U6104 (N_6104,N_4944,N_966);
nor U6105 (N_6105,N_4488,N_56);
xor U6106 (N_6106,N_1113,N_4266);
nand U6107 (N_6107,N_3916,N_4361);
nor U6108 (N_6108,N_1320,N_3851);
nor U6109 (N_6109,N_2740,N_1331);
nand U6110 (N_6110,N_4422,N_4104);
and U6111 (N_6111,N_4753,N_1207);
nor U6112 (N_6112,N_481,N_3575);
nor U6113 (N_6113,N_2199,N_4073);
and U6114 (N_6114,N_3812,N_4907);
xor U6115 (N_6115,N_4848,N_3926);
xnor U6116 (N_6116,N_150,N_4834);
xor U6117 (N_6117,N_110,N_341);
nor U6118 (N_6118,N_782,N_4556);
nor U6119 (N_6119,N_1995,N_95);
nand U6120 (N_6120,N_4720,N_602);
nand U6121 (N_6121,N_1078,N_1657);
or U6122 (N_6122,N_4929,N_3170);
nor U6123 (N_6123,N_3358,N_4391);
or U6124 (N_6124,N_3836,N_3111);
nor U6125 (N_6125,N_2835,N_3593);
xor U6126 (N_6126,N_1685,N_172);
or U6127 (N_6127,N_4485,N_728);
and U6128 (N_6128,N_4807,N_3909);
or U6129 (N_6129,N_1952,N_4577);
or U6130 (N_6130,N_12,N_626);
nor U6131 (N_6131,N_1586,N_4106);
or U6132 (N_6132,N_1854,N_1612);
and U6133 (N_6133,N_4181,N_3285);
or U6134 (N_6134,N_1245,N_1988);
and U6135 (N_6135,N_3699,N_1270);
or U6136 (N_6136,N_3616,N_3308);
nand U6137 (N_6137,N_4251,N_139);
and U6138 (N_6138,N_4076,N_1447);
or U6139 (N_6139,N_1379,N_4690);
nor U6140 (N_6140,N_457,N_4253);
xnor U6141 (N_6141,N_4327,N_3945);
nand U6142 (N_6142,N_177,N_1171);
or U6143 (N_6143,N_958,N_69);
nor U6144 (N_6144,N_1773,N_3329);
nand U6145 (N_6145,N_4761,N_3826);
and U6146 (N_6146,N_2483,N_414);
nand U6147 (N_6147,N_2869,N_3258);
nand U6148 (N_6148,N_450,N_576);
xor U6149 (N_6149,N_781,N_3570);
and U6150 (N_6150,N_1389,N_1658);
and U6151 (N_6151,N_1150,N_1587);
or U6152 (N_6152,N_4543,N_2330);
and U6153 (N_6153,N_2843,N_2571);
nand U6154 (N_6154,N_2924,N_2748);
xnor U6155 (N_6155,N_1048,N_3919);
nor U6156 (N_6156,N_615,N_4146);
or U6157 (N_6157,N_4262,N_356);
or U6158 (N_6158,N_2535,N_1102);
and U6159 (N_6159,N_4447,N_3612);
or U6160 (N_6160,N_3757,N_370);
and U6161 (N_6161,N_2430,N_4695);
nand U6162 (N_6162,N_2022,N_2074);
xor U6163 (N_6163,N_4270,N_3346);
nor U6164 (N_6164,N_1644,N_1302);
nand U6165 (N_6165,N_796,N_871);
nor U6166 (N_6166,N_409,N_633);
and U6167 (N_6167,N_3068,N_2731);
nand U6168 (N_6168,N_4557,N_3345);
xor U6169 (N_6169,N_3744,N_2104);
or U6170 (N_6170,N_3942,N_3409);
and U6171 (N_6171,N_3653,N_1255);
nor U6172 (N_6172,N_2525,N_1338);
nand U6173 (N_6173,N_1604,N_1865);
nand U6174 (N_6174,N_4459,N_231);
and U6175 (N_6175,N_759,N_3342);
and U6176 (N_6176,N_1873,N_3039);
and U6177 (N_6177,N_1479,N_3283);
or U6178 (N_6178,N_220,N_4583);
xnor U6179 (N_6179,N_6,N_1500);
nor U6180 (N_6180,N_2863,N_1186);
or U6181 (N_6181,N_3905,N_1278);
nor U6182 (N_6182,N_274,N_823);
and U6183 (N_6183,N_751,N_3343);
and U6184 (N_6184,N_989,N_3943);
xor U6185 (N_6185,N_1541,N_1178);
nor U6186 (N_6186,N_3274,N_4483);
or U6187 (N_6187,N_4863,N_3058);
nand U6188 (N_6188,N_2918,N_3783);
nor U6189 (N_6189,N_4402,N_259);
nor U6190 (N_6190,N_2054,N_1567);
and U6191 (N_6191,N_3417,N_726);
xor U6192 (N_6192,N_2542,N_2356);
and U6193 (N_6193,N_3527,N_4664);
or U6194 (N_6194,N_4259,N_4471);
nor U6195 (N_6195,N_2787,N_3515);
nand U6196 (N_6196,N_2674,N_4961);
nor U6197 (N_6197,N_3192,N_3292);
or U6198 (N_6198,N_4222,N_1010);
or U6199 (N_6199,N_3470,N_2506);
and U6200 (N_6200,N_3130,N_307);
xor U6201 (N_6201,N_4672,N_1092);
nor U6202 (N_6202,N_2667,N_2187);
and U6203 (N_6203,N_1306,N_360);
and U6204 (N_6204,N_1237,N_1929);
xor U6205 (N_6205,N_1139,N_4629);
nand U6206 (N_6206,N_4721,N_2743);
and U6207 (N_6207,N_1869,N_4545);
nor U6208 (N_6208,N_135,N_2618);
nor U6209 (N_6209,N_2709,N_791);
and U6210 (N_6210,N_169,N_2107);
nor U6211 (N_6211,N_131,N_3150);
and U6212 (N_6212,N_2631,N_736);
and U6213 (N_6213,N_2993,N_587);
or U6214 (N_6214,N_4254,N_806);
and U6215 (N_6215,N_2457,N_3973);
and U6216 (N_6216,N_794,N_900);
nand U6217 (N_6217,N_1332,N_3562);
or U6218 (N_6218,N_2913,N_111);
xnor U6219 (N_6219,N_3351,N_3756);
nand U6220 (N_6220,N_1480,N_1493);
nand U6221 (N_6221,N_1022,N_2284);
and U6222 (N_6222,N_3993,N_1212);
or U6223 (N_6223,N_362,N_731);
xnor U6224 (N_6224,N_3798,N_912);
nand U6225 (N_6225,N_3689,N_3805);
and U6226 (N_6226,N_1313,N_2760);
xnor U6227 (N_6227,N_258,N_4892);
xor U6228 (N_6228,N_4435,N_1550);
nor U6229 (N_6229,N_746,N_283);
nor U6230 (N_6230,N_1475,N_4346);
nand U6231 (N_6231,N_1522,N_1451);
or U6232 (N_6232,N_2195,N_1090);
nor U6233 (N_6233,N_1634,N_3835);
nand U6234 (N_6234,N_1863,N_500);
nand U6235 (N_6235,N_3743,N_1145);
and U6236 (N_6236,N_4990,N_4928);
nor U6237 (N_6237,N_3823,N_4623);
xor U6238 (N_6238,N_3788,N_4687);
and U6239 (N_6239,N_3786,N_1811);
nor U6240 (N_6240,N_3041,N_2287);
and U6241 (N_6241,N_742,N_1976);
nand U6242 (N_6242,N_1682,N_1689);
nand U6243 (N_6243,N_1248,N_1464);
and U6244 (N_6244,N_4428,N_454);
nor U6245 (N_6245,N_3958,N_1434);
and U6246 (N_6246,N_2653,N_433);
nor U6247 (N_6247,N_838,N_3564);
xnor U6248 (N_6248,N_1031,N_3853);
or U6249 (N_6249,N_4178,N_1542);
and U6250 (N_6250,N_903,N_1528);
nand U6251 (N_6251,N_639,N_1260);
nor U6252 (N_6252,N_2569,N_673);
xnor U6253 (N_6253,N_2237,N_492);
and U6254 (N_6254,N_2492,N_3221);
or U6255 (N_6255,N_539,N_593);
nand U6256 (N_6256,N_2379,N_919);
nor U6257 (N_6257,N_1582,N_4210);
or U6258 (N_6258,N_3768,N_3876);
nand U6259 (N_6259,N_417,N_4268);
xor U6260 (N_6260,N_4053,N_2833);
xor U6261 (N_6261,N_1123,N_3340);
or U6262 (N_6262,N_1957,N_1563);
xnor U6263 (N_6263,N_3268,N_2036);
nand U6264 (N_6264,N_46,N_4824);
or U6265 (N_6265,N_2037,N_2135);
nor U6266 (N_6266,N_4419,N_1213);
or U6267 (N_6267,N_1904,N_125);
nor U6268 (N_6268,N_555,N_4998);
nor U6269 (N_6269,N_472,N_3225);
xor U6270 (N_6270,N_1226,N_1310);
or U6271 (N_6271,N_4155,N_2751);
or U6272 (N_6272,N_927,N_922);
or U6273 (N_6273,N_2007,N_221);
or U6274 (N_6274,N_3697,N_2893);
nand U6275 (N_6275,N_907,N_4606);
xor U6276 (N_6276,N_1039,N_3034);
nor U6277 (N_6277,N_1962,N_107);
xnor U6278 (N_6278,N_1652,N_3420);
and U6279 (N_6279,N_4252,N_3333);
nor U6280 (N_6280,N_1872,N_885);
or U6281 (N_6281,N_4328,N_1264);
nor U6282 (N_6282,N_3286,N_942);
xor U6283 (N_6283,N_3266,N_304);
nand U6284 (N_6284,N_4829,N_2934);
and U6285 (N_6285,N_330,N_29);
xnor U6286 (N_6286,N_2665,N_775);
xor U6287 (N_6287,N_3991,N_4614);
nand U6288 (N_6288,N_2372,N_2635);
and U6289 (N_6289,N_3215,N_761);
and U6290 (N_6290,N_3458,N_2892);
or U6291 (N_6291,N_2164,N_1218);
nand U6292 (N_6292,N_1189,N_2644);
nand U6293 (N_6293,N_3293,N_2256);
and U6294 (N_6294,N_3759,N_3270);
nor U6295 (N_6295,N_4835,N_1670);
nor U6296 (N_6296,N_2179,N_1360);
or U6297 (N_6297,N_1252,N_2276);
nand U6298 (N_6298,N_210,N_87);
xor U6299 (N_6299,N_3339,N_4836);
and U6300 (N_6300,N_3953,N_4726);
nor U6301 (N_6301,N_3313,N_4247);
xnor U6302 (N_6302,N_4772,N_4685);
nor U6303 (N_6303,N_2232,N_3814);
nand U6304 (N_6304,N_3734,N_512);
nor U6305 (N_6305,N_4902,N_3936);
or U6306 (N_6306,N_1985,N_1384);
or U6307 (N_6307,N_3772,N_189);
nor U6308 (N_6308,N_242,N_2234);
nor U6309 (N_6309,N_2792,N_1614);
or U6310 (N_6310,N_3929,N_715);
nand U6311 (N_6311,N_1886,N_365);
nand U6312 (N_6312,N_4345,N_1206);
nor U6313 (N_6313,N_2794,N_1420);
nand U6314 (N_6314,N_3234,N_4611);
nand U6315 (N_6315,N_1628,N_692);
nor U6316 (N_6316,N_1783,N_2205);
and U6317 (N_6317,N_2062,N_3867);
and U6318 (N_6318,N_2746,N_1261);
xor U6319 (N_6319,N_1027,N_1880);
or U6320 (N_6320,N_1996,N_2617);
nor U6321 (N_6321,N_33,N_2822);
nor U6322 (N_6322,N_2143,N_1073);
and U6323 (N_6323,N_1341,N_2774);
nand U6324 (N_6324,N_4679,N_1664);
or U6325 (N_6325,N_2966,N_562);
xor U6326 (N_6326,N_145,N_2636);
and U6327 (N_6327,N_351,N_4673);
or U6328 (N_6328,N_917,N_2630);
nand U6329 (N_6329,N_3211,N_2992);
or U6330 (N_6330,N_2932,N_3816);
or U6331 (N_6331,N_2266,N_701);
or U6332 (N_6332,N_3354,N_888);
nand U6333 (N_6333,N_4566,N_2272);
and U6334 (N_6334,N_373,N_886);
xor U6335 (N_6335,N_1735,N_3186);
xnor U6336 (N_6336,N_4219,N_465);
or U6337 (N_6337,N_843,N_284);
and U6338 (N_6338,N_4908,N_3778);
or U6339 (N_6339,N_2786,N_3849);
xor U6340 (N_6340,N_3765,N_2681);
nor U6341 (N_6341,N_183,N_4825);
xnor U6342 (N_6342,N_4532,N_2129);
and U6343 (N_6343,N_4619,N_2058);
and U6344 (N_6344,N_4826,N_2507);
and U6345 (N_6345,N_1823,N_3789);
or U6346 (N_6346,N_4382,N_4302);
nor U6347 (N_6347,N_554,N_4696);
nand U6348 (N_6348,N_2884,N_511);
nand U6349 (N_6349,N_1750,N_34);
nand U6350 (N_6350,N_1782,N_3661);
or U6351 (N_6351,N_4674,N_1704);
and U6352 (N_6352,N_4708,N_1353);
nor U6353 (N_6353,N_1323,N_4276);
and U6354 (N_6354,N_4199,N_1858);
and U6355 (N_6355,N_4153,N_4579);
xnor U6356 (N_6356,N_2900,N_238);
and U6357 (N_6357,N_2904,N_1734);
xnor U6358 (N_6358,N_1408,N_1151);
or U6359 (N_6359,N_480,N_392);
nor U6360 (N_6360,N_4784,N_4072);
xnor U6361 (N_6361,N_3842,N_2019);
or U6362 (N_6362,N_1146,N_369);
xor U6363 (N_6363,N_604,N_4694);
or U6364 (N_6364,N_1741,N_986);
or U6365 (N_6365,N_3621,N_1368);
and U6366 (N_6366,N_2650,N_118);
nand U6367 (N_6367,N_3161,N_1661);
nand U6368 (N_6368,N_4963,N_2262);
xnor U6369 (N_6369,N_4387,N_3344);
or U6370 (N_6370,N_1778,N_448);
or U6371 (N_6371,N_359,N_3110);
or U6372 (N_6372,N_4039,N_2156);
nor U6373 (N_6373,N_734,N_2500);
nand U6374 (N_6374,N_4448,N_2788);
and U6375 (N_6375,N_4279,N_3712);
nor U6376 (N_6376,N_2809,N_1641);
nor U6377 (N_6377,N_1091,N_215);
xnor U6378 (N_6378,N_2576,N_193);
or U6379 (N_6379,N_4597,N_2660);
nand U6380 (N_6380,N_3752,N_3421);
nor U6381 (N_6381,N_1372,N_4911);
xnor U6382 (N_6382,N_859,N_2008);
xor U6383 (N_6383,N_4805,N_1499);
or U6384 (N_6384,N_874,N_1484);
nand U6385 (N_6385,N_375,N_2528);
nor U6386 (N_6386,N_4228,N_1436);
and U6387 (N_6387,N_1724,N_4197);
and U6388 (N_6388,N_566,N_649);
nand U6389 (N_6389,N_4417,N_2879);
and U6390 (N_6390,N_1196,N_2466);
and U6391 (N_6391,N_697,N_1894);
and U6392 (N_6392,N_2693,N_632);
nor U6393 (N_6393,N_3219,N_3263);
nand U6394 (N_6394,N_3382,N_523);
and U6395 (N_6395,N_165,N_3538);
nor U6396 (N_6396,N_254,N_4468);
and U6397 (N_6397,N_1878,N_3811);
nor U6398 (N_6398,N_4046,N_672);
and U6399 (N_6399,N_3897,N_617);
xor U6400 (N_6400,N_2806,N_2318);
or U6401 (N_6401,N_1557,N_108);
nand U6402 (N_6402,N_4038,N_3422);
and U6403 (N_6403,N_3595,N_3549);
xnor U6404 (N_6404,N_4519,N_305);
or U6405 (N_6405,N_4157,N_2253);
or U6406 (N_6406,N_3012,N_3120);
nand U6407 (N_6407,N_3247,N_1174);
xor U6408 (N_6408,N_4717,N_693);
nand U6409 (N_6409,N_2795,N_1203);
nand U6410 (N_6410,N_3970,N_2279);
or U6411 (N_6411,N_773,N_2800);
nand U6412 (N_6412,N_1001,N_1655);
and U6413 (N_6413,N_2063,N_4389);
nor U6414 (N_6414,N_3151,N_3672);
or U6415 (N_6415,N_1806,N_3807);
xnor U6416 (N_6416,N_3207,N_366);
nand U6417 (N_6417,N_1241,N_65);
nor U6418 (N_6418,N_2909,N_2588);
nand U6419 (N_6419,N_1964,N_2834);
and U6420 (N_6420,N_628,N_4156);
and U6421 (N_6421,N_3947,N_4383);
nor U6422 (N_6422,N_2767,N_696);
xnor U6423 (N_6423,N_987,N_747);
and U6424 (N_6424,N_1193,N_772);
xnor U6425 (N_6425,N_3236,N_2532);
nor U6426 (N_6426,N_2480,N_3882);
or U6427 (N_6427,N_3623,N_3847);
xnor U6428 (N_6428,N_774,N_3441);
nor U6429 (N_6429,N_463,N_2247);
nand U6430 (N_6430,N_101,N_91);
and U6431 (N_6431,N_4655,N_4494);
and U6432 (N_6432,N_976,N_3165);
and U6433 (N_6433,N_4218,N_1035);
or U6434 (N_6434,N_96,N_2226);
nor U6435 (N_6435,N_998,N_2080);
nor U6436 (N_6436,N_3533,N_2598);
and U6437 (N_6437,N_2423,N_2314);
or U6438 (N_6438,N_4444,N_678);
xnor U6439 (N_6439,N_2468,N_1033);
nand U6440 (N_6440,N_4958,N_498);
or U6441 (N_6441,N_285,N_1804);
nand U6442 (N_6442,N_1060,N_1108);
nand U6443 (N_6443,N_2519,N_4498);
and U6444 (N_6444,N_3745,N_1400);
and U6445 (N_6445,N_70,N_3048);
nor U6446 (N_6446,N_1545,N_921);
xor U6447 (N_6447,N_4213,N_2098);
or U6448 (N_6448,N_4635,N_1577);
xnor U6449 (N_6449,N_4478,N_2238);
and U6450 (N_6450,N_3216,N_1608);
nor U6451 (N_6451,N_4338,N_2015);
xnor U6452 (N_6452,N_2178,N_2209);
nand U6453 (N_6453,N_88,N_710);
or U6454 (N_6454,N_4815,N_2676);
nor U6455 (N_6455,N_2275,N_1445);
and U6456 (N_6456,N_4646,N_3996);
or U6457 (N_6457,N_1491,N_2818);
nor U6458 (N_6458,N_2917,N_1176);
nand U6459 (N_6459,N_3990,N_2866);
nor U6460 (N_6460,N_3981,N_2173);
and U6461 (N_6461,N_793,N_3874);
or U6462 (N_6462,N_3194,N_785);
and U6463 (N_6463,N_3906,N_2055);
nor U6464 (N_6464,N_182,N_911);
nor U6465 (N_6465,N_2624,N_837);
nor U6466 (N_6466,N_3655,N_4467);
nor U6467 (N_6467,N_4090,N_4206);
nand U6468 (N_6468,N_3383,N_2634);
nand U6469 (N_6469,N_4472,N_534);
and U6470 (N_6470,N_416,N_3468);
or U6471 (N_6471,N_2411,N_1347);
xor U6472 (N_6472,N_1759,N_1882);
and U6473 (N_6473,N_3459,N_4407);
xnor U6474 (N_6474,N_3588,N_1737);
and U6475 (N_6475,N_4728,N_3696);
or U6476 (N_6476,N_1853,N_2023);
nor U6477 (N_6477,N_2115,N_1815);
xnor U6478 (N_6478,N_3864,N_2206);
or U6479 (N_6479,N_3427,N_792);
nand U6480 (N_6480,N_644,N_3267);
and U6481 (N_6481,N_1052,N_3665);
nand U6482 (N_6482,N_675,N_3762);
nand U6483 (N_6483,N_740,N_2633);
nand U6484 (N_6484,N_4563,N_4475);
nor U6485 (N_6485,N_4411,N_4426);
xor U6486 (N_6486,N_3311,N_1217);
nand U6487 (N_6487,N_2350,N_1742);
xor U6488 (N_6488,N_3887,N_2670);
nor U6489 (N_6489,N_2742,N_1290);
or U6490 (N_6490,N_186,N_428);
or U6491 (N_6491,N_3447,N_1294);
nor U6492 (N_6492,N_3179,N_522);
or U6493 (N_6493,N_2718,N_4111);
nand U6494 (N_6494,N_4757,N_4877);
or U6495 (N_6495,N_2607,N_868);
or U6496 (N_6496,N_3888,N_3226);
nand U6497 (N_6497,N_3467,N_4424);
and U6498 (N_6498,N_1308,N_611);
nand U6499 (N_6499,N_4984,N_1524);
nand U6500 (N_6500,N_1390,N_1547);
nand U6501 (N_6501,N_342,N_1710);
xor U6502 (N_6502,N_1135,N_2089);
or U6503 (N_6503,N_4032,N_1757);
nand U6504 (N_6504,N_4638,N_4023);
or U6505 (N_6505,N_2121,N_667);
or U6506 (N_6506,N_3360,N_2295);
nor U6507 (N_6507,N_4663,N_4751);
nor U6508 (N_6508,N_1775,N_2646);
nand U6509 (N_6509,N_2831,N_2160);
nor U6510 (N_6510,N_3670,N_1721);
nor U6511 (N_6511,N_586,N_950);
nand U6512 (N_6512,N_1817,N_877);
xnor U6513 (N_6513,N_37,N_501);
and U6514 (N_6514,N_3397,N_129);
and U6515 (N_6515,N_3704,N_4273);
nor U6516 (N_6516,N_3291,N_2229);
and U6517 (N_6517,N_4667,N_1512);
xor U6518 (N_6518,N_2827,N_816);
nor U6519 (N_6519,N_2911,N_2033);
or U6520 (N_6520,N_3763,N_3230);
nor U6521 (N_6521,N_3001,N_2602);
xnor U6522 (N_6522,N_2433,N_1432);
nor U6523 (N_6523,N_2947,N_4455);
and U6524 (N_6524,N_1051,N_352);
nor U6525 (N_6525,N_1167,N_668);
nor U6526 (N_6526,N_105,N_1376);
or U6527 (N_6527,N_4666,N_382);
nand U6528 (N_6528,N_2723,N_2679);
and U6529 (N_6529,N_2925,N_3622);
and U6530 (N_6530,N_3844,N_4650);
nand U6531 (N_6531,N_2680,N_1265);
nor U6532 (N_6532,N_449,N_1391);
and U6533 (N_6533,N_1340,N_3407);
nand U6534 (N_6534,N_4847,N_2620);
and U6535 (N_6535,N_1109,N_1127);
or U6536 (N_6536,N_4510,N_4949);
nand U6537 (N_6537,N_3854,N_4586);
xnor U6538 (N_6538,N_4295,N_1726);
nor U6539 (N_6539,N_723,N_1950);
nor U6540 (N_6540,N_3571,N_1762);
nor U6541 (N_6541,N_1269,N_577);
nand U6542 (N_6542,N_575,N_4697);
and U6543 (N_6543,N_2790,N_3994);
nor U6544 (N_6544,N_2982,N_2675);
or U6545 (N_6545,N_4109,N_4122);
xnor U6546 (N_6546,N_4020,N_1025);
nand U6547 (N_6547,N_1093,N_1920);
nor U6548 (N_6548,N_2551,N_3038);
nor U6549 (N_6549,N_4814,N_1118);
nand U6550 (N_6550,N_2661,N_3928);
xnor U6551 (N_6551,N_1994,N_3950);
nor U6552 (N_6552,N_1781,N_3040);
nor U6553 (N_6553,N_3080,N_212);
xnor U6554 (N_6554,N_2259,N_4734);
nor U6555 (N_6555,N_2313,N_3097);
nor U6556 (N_6556,N_1000,N_1583);
xnor U6557 (N_6557,N_3954,N_3868);
or U6558 (N_6558,N_4743,N_1859);
xor U6559 (N_6559,N_2216,N_4971);
nand U6560 (N_6560,N_2684,N_2274);
nor U6561 (N_6561,N_346,N_1062);
or U6562 (N_6562,N_2819,N_2362);
nand U6563 (N_6563,N_3960,N_563);
nor U6564 (N_6564,N_2327,N_3702);
nor U6565 (N_6565,N_67,N_802);
xnor U6566 (N_6566,N_4881,N_750);
nand U6567 (N_6567,N_581,N_368);
or U6568 (N_6568,N_2105,N_1239);
or U6569 (N_6569,N_3078,N_2529);
nand U6570 (N_6570,N_1496,N_1526);
nor U6571 (N_6571,N_1194,N_3172);
or U6572 (N_6572,N_3396,N_4132);
and U6573 (N_6573,N_685,N_849);
xnor U6574 (N_6574,N_1192,N_2826);
and U6575 (N_6575,N_1991,N_3102);
xor U6576 (N_6576,N_4940,N_2324);
or U6577 (N_6577,N_2508,N_411);
nand U6578 (N_6578,N_0,N_4762);
nand U6579 (N_6579,N_4972,N_1566);
nand U6580 (N_6580,N_1617,N_1250);
or U6581 (N_6581,N_4154,N_1698);
xnor U6582 (N_6582,N_3626,N_1527);
xnor U6583 (N_6583,N_4284,N_2544);
and U6584 (N_6584,N_3250,N_2706);
xnor U6585 (N_6585,N_3129,N_3364);
or U6586 (N_6586,N_1315,N_4353);
or U6587 (N_6587,N_4008,N_3388);
nand U6588 (N_6588,N_3435,N_2368);
or U6589 (N_6589,N_4306,N_1172);
or U6590 (N_6590,N_3505,N_2640);
nor U6591 (N_6591,N_2895,N_2828);
or U6592 (N_6592,N_3096,N_1974);
nor U6593 (N_6593,N_4066,N_597);
or U6594 (N_6594,N_3540,N_4508);
xor U6595 (N_6595,N_1509,N_4277);
or U6596 (N_6596,N_2764,N_3077);
or U6597 (N_6597,N_1431,N_4558);
xor U6598 (N_6598,N_1263,N_4952);
nor U6599 (N_6599,N_2715,N_478);
xor U6600 (N_6600,N_1531,N_3056);
nor U6601 (N_6601,N_4565,N_2169);
xnor U6602 (N_6602,N_1312,N_830);
nor U6603 (N_6603,N_4043,N_3314);
nand U6604 (N_6604,N_1352,N_2029);
or U6605 (N_6605,N_2603,N_4764);
or U6606 (N_6606,N_4054,N_2574);
nor U6607 (N_6607,N_2296,N_893);
xnor U6608 (N_6608,N_2122,N_2768);
nor U6609 (N_6609,N_2972,N_2046);
nor U6610 (N_6610,N_4542,N_3131);
xor U6611 (N_6611,N_570,N_596);
and U6612 (N_6612,N_872,N_2221);
xor U6613 (N_6613,N_64,N_2663);
nand U6614 (N_6614,N_1058,N_2011);
and U6615 (N_6615,N_3817,N_4615);
xor U6616 (N_6616,N_1813,N_3222);
xor U6617 (N_6617,N_228,N_1945);
nor U6618 (N_6618,N_3019,N_3355);
or U6619 (N_6619,N_754,N_2687);
nand U6620 (N_6620,N_395,N_1860);
xor U6621 (N_6621,N_855,N_2713);
and U6622 (N_6622,N_1358,N_1922);
and U6623 (N_6623,N_3813,N_2168);
nor U6624 (N_6624,N_4682,N_1359);
xor U6625 (N_6625,N_3461,N_1271);
nand U6626 (N_6626,N_3495,N_2231);
xor U6627 (N_6627,N_918,N_130);
nor U6628 (N_6628,N_1029,N_2587);
nor U6629 (N_6629,N_745,N_544);
and U6630 (N_6630,N_3785,N_1845);
xnor U6631 (N_6631,N_1037,N_3760);
nand U6632 (N_6632,N_2610,N_4208);
and U6633 (N_6633,N_2328,N_3133);
xnor U6634 (N_6634,N_1961,N_1931);
xnor U6635 (N_6635,N_85,N_4167);
or U6636 (N_6636,N_364,N_2484);
and U6637 (N_6637,N_4601,N_4481);
and U6638 (N_6638,N_2416,N_4585);
nand U6639 (N_6639,N_4625,N_3885);
nor U6640 (N_6640,N_4517,N_2505);
or U6641 (N_6641,N_4263,N_1140);
and U6642 (N_6642,N_1231,N_2548);
and U6643 (N_6643,N_154,N_2654);
xor U6644 (N_6644,N_1214,N_4202);
nand U6645 (N_6645,N_2285,N_1328);
nor U6646 (N_6646,N_2069,N_1561);
and U6647 (N_6647,N_707,N_4098);
xor U6648 (N_6648,N_4842,N_623);
nor U6649 (N_6649,N_2128,N_2590);
nor U6650 (N_6650,N_4681,N_3921);
nand U6651 (N_6651,N_822,N_1793);
nor U6652 (N_6652,N_766,N_3872);
xor U6653 (N_6653,N_3633,N_4733);
or U6654 (N_6654,N_3373,N_4439);
nor U6655 (N_6655,N_1053,N_460);
and U6656 (N_6656,N_2412,N_2888);
nor U6657 (N_6657,N_3733,N_4700);
nor U6658 (N_6658,N_4813,N_3356);
or U6659 (N_6659,N_2083,N_2413);
nor U6660 (N_6660,N_2406,N_861);
nor U6661 (N_6661,N_4535,N_1953);
nor U6662 (N_6662,N_3024,N_3804);
xnor U6663 (N_6663,N_3411,N_3671);
nand U6664 (N_6664,N_4839,N_4236);
and U6665 (N_6665,N_1259,N_479);
nand U6666 (N_6666,N_3599,N_2695);
xnor U6667 (N_6667,N_3901,N_3726);
xnor U6668 (N_6668,N_1999,N_2118);
nand U6669 (N_6669,N_1647,N_4329);
nor U6670 (N_6670,N_204,N_1161);
or U6671 (N_6671,N_3338,N_1812);
xor U6672 (N_6672,N_3894,N_654);
and U6673 (N_6673,N_2047,N_97);
nand U6674 (N_6674,N_2698,N_260);
xor U6675 (N_6675,N_4992,N_4400);
and U6676 (N_6676,N_3473,N_4554);
xnor U6677 (N_6677,N_4386,N_1552);
xnor U6678 (N_6678,N_2881,N_1202);
xor U6679 (N_6679,N_4889,N_4821);
nor U6680 (N_6680,N_4920,N_4798);
or U6681 (N_6681,N_2499,N_2641);
nand U6682 (N_6682,N_100,N_3146);
and U6683 (N_6683,N_4888,N_4841);
nor U6684 (N_6684,N_3766,N_4736);
or U6685 (N_6685,N_73,N_4194);
xnor U6686 (N_6686,N_2183,N_1978);
nand U6687 (N_6687,N_4659,N_2523);
nand U6688 (N_6688,N_1699,N_3026);
xor U6689 (N_6689,N_953,N_2965);
xor U6690 (N_6690,N_1897,N_717);
and U6691 (N_6691,N_2568,N_3645);
xnor U6692 (N_6692,N_2139,N_4506);
or U6693 (N_6693,N_4056,N_4680);
and U6694 (N_6694,N_1333,N_748);
xnor U6695 (N_6695,N_4996,N_3303);
and U6696 (N_6696,N_4249,N_2250);
and U6697 (N_6697,N_267,N_2954);
xnor U6698 (N_6698,N_113,N_2125);
nand U6699 (N_6699,N_371,N_594);
nor U6700 (N_6700,N_3310,N_1877);
and U6701 (N_6701,N_1686,N_3741);
nor U6702 (N_6702,N_4538,N_198);
nand U6703 (N_6703,N_2452,N_2961);
and U6704 (N_6704,N_253,N_1130);
and U6705 (N_6705,N_3132,N_2239);
nor U6706 (N_6706,N_2770,N_136);
nor U6707 (N_6707,N_590,N_3499);
and U6708 (N_6708,N_300,N_1505);
or U6709 (N_6709,N_4216,N_2053);
or U6710 (N_6710,N_1466,N_3053);
and U6711 (N_6711,N_2559,N_1651);
or U6712 (N_6712,N_3235,N_3962);
and U6713 (N_6713,N_4882,N_2482);
or U6714 (N_6714,N_367,N_2908);
and U6715 (N_6715,N_4580,N_1074);
xor U6716 (N_6716,N_3474,N_4574);
and U6717 (N_6717,N_2165,N_690);
xor U6718 (N_6718,N_207,N_3385);
or U6719 (N_6719,N_4812,N_3703);
or U6720 (N_6720,N_4427,N_1746);
nand U6721 (N_6721,N_3941,N_3240);
and U6722 (N_6722,N_2849,N_1606);
nand U6723 (N_6723,N_4918,N_4033);
and U6724 (N_6724,N_4074,N_194);
or U6725 (N_6725,N_311,N_2158);
or U6726 (N_6726,N_3735,N_4152);
nor U6727 (N_6727,N_3614,N_3717);
or U6728 (N_6728,N_2860,N_520);
or U6729 (N_6729,N_2064,N_2471);
or U6730 (N_6730,N_529,N_1764);
or U6731 (N_6731,N_2404,N_3404);
and U6732 (N_6732,N_2236,N_1930);
nand U6733 (N_6733,N_426,N_4906);
nand U6734 (N_6734,N_1846,N_1233);
nand U6735 (N_6735,N_1849,N_1124);
xor U6736 (N_6736,N_3737,N_292);
xnor U6737 (N_6737,N_1575,N_128);
xor U6738 (N_6738,N_4026,N_1584);
and U6739 (N_6739,N_83,N_4085);
xor U6740 (N_6740,N_2432,N_4609);
xnor U6741 (N_6741,N_1619,N_2980);
nor U6742 (N_6742,N_2182,N_559);
and U6743 (N_6743,N_3119,N_4742);
nor U6744 (N_6744,N_4330,N_1816);
nand U6745 (N_6745,N_4477,N_1134);
or U6746 (N_6746,N_733,N_2270);
or U6747 (N_6747,N_1056,N_4006);
and U6748 (N_6748,N_4846,N_1772);
xnor U6749 (N_6749,N_4922,N_4552);
and U6750 (N_6750,N_2479,N_4452);
or U6751 (N_6751,N_2371,N_3609);
and U6752 (N_6752,N_3284,N_2622);
and U6753 (N_6753,N_757,N_4924);
nor U6754 (N_6754,N_1917,N_2381);
xor U6755 (N_6755,N_2894,N_3719);
nor U6756 (N_6756,N_4225,N_783);
xnor U6757 (N_6757,N_2782,N_4170);
nand U6758 (N_6758,N_2619,N_3185);
xor U6759 (N_6759,N_561,N_1159);
nor U6760 (N_6760,N_2664,N_2215);
or U6761 (N_6761,N_1558,N_4589);
nor U6762 (N_6762,N_680,N_149);
xnor U6763 (N_6763,N_2298,N_2387);
or U6764 (N_6764,N_4575,N_4536);
and U6765 (N_6765,N_2625,N_4533);
xnor U6766 (N_6766,N_2020,N_1540);
nor U6767 (N_6767,N_3189,N_1881);
xnor U6768 (N_6768,N_2658,N_4250);
and U6769 (N_6769,N_1639,N_2608);
nand U6770 (N_6770,N_4240,N_2543);
nor U6771 (N_6771,N_2875,N_3600);
and U6772 (N_6772,N_2777,N_4458);
and U6773 (N_6773,N_2081,N_3177);
and U6774 (N_6774,N_1375,N_4569);
xor U6775 (N_6775,N_850,N_4531);
nand U6776 (N_6776,N_3248,N_3834);
nor U6777 (N_6777,N_4705,N_2150);
or U6778 (N_6778,N_1288,N_3736);
nand U6779 (N_6779,N_1165,N_2458);
xor U6780 (N_6780,N_3965,N_4094);
or U6781 (N_6781,N_1902,N_3337);
or U6782 (N_6782,N_1152,N_3136);
xor U6783 (N_6783,N_1386,N_1258);
nand U6784 (N_6784,N_1296,N_3652);
and U6785 (N_6785,N_278,N_1602);
and U6786 (N_6786,N_3439,N_4057);
nand U6787 (N_6787,N_1914,N_3350);
and U6788 (N_6788,N_482,N_2534);
xor U6789 (N_6789,N_2013,N_659);
or U6790 (N_6790,N_4737,N_1979);
nor U6791 (N_6791,N_1185,N_2793);
xor U6792 (N_6792,N_3209,N_429);
nand U6793 (N_6793,N_4165,N_4425);
nand U6794 (N_6794,N_873,N_565);
xnor U6795 (N_6795,N_2145,N_1514);
nand U6796 (N_6796,N_2518,N_516);
and U6797 (N_6797,N_1870,N_4713);
xnor U6798 (N_6798,N_2200,N_4956);
or U6799 (N_6799,N_810,N_936);
nor U6800 (N_6800,N_1364,N_2593);
nand U6801 (N_6801,N_2151,N_1362);
xnor U6802 (N_6802,N_3646,N_393);
nor U6803 (N_6803,N_4119,N_1529);
nor U6804 (N_6804,N_109,N_256);
and U6805 (N_6805,N_1725,N_1181);
nand U6806 (N_6806,N_1225,N_16);
or U6807 (N_6807,N_3568,N_35);
nand U6808 (N_6808,N_2615,N_3047);
xor U6809 (N_6809,N_3372,N_2336);
or U6810 (N_6810,N_2705,N_2456);
nand U6811 (N_6811,N_2066,N_4499);
nand U6812 (N_6812,N_4366,N_1148);
nor U6813 (N_6813,N_1107,N_3630);
nand U6814 (N_6814,N_248,N_1160);
or U6815 (N_6815,N_870,N_4965);
or U6816 (N_6816,N_2562,N_3437);
nand U6817 (N_6817,N_2886,N_3154);
xnor U6818 (N_6818,N_142,N_4884);
nor U6819 (N_6819,N_4979,N_153);
or U6820 (N_6820,N_3603,N_2537);
or U6821 (N_6821,N_1989,N_273);
and U6822 (N_6822,N_3690,N_4408);
xor U6823 (N_6823,N_175,N_4593);
nor U6824 (N_6824,N_4985,N_4995);
and U6825 (N_6825,N_3341,N_2446);
nand U6826 (N_6826,N_363,N_2395);
nand U6827 (N_6827,N_2181,N_3793);
and U6828 (N_6828,N_133,N_2513);
nor U6829 (N_6829,N_3135,N_1554);
nor U6830 (N_6830,N_4791,N_320);
nand U6831 (N_6831,N_4975,N_3184);
nor U6832 (N_6832,N_841,N_756);
or U6833 (N_6833,N_3522,N_627);
xor U6834 (N_6834,N_4350,N_666);
nor U6835 (N_6835,N_57,N_197);
xor U6836 (N_6836,N_1580,N_3619);
xor U6837 (N_6837,N_4838,N_3501);
and U6838 (N_6838,N_3494,N_996);
nand U6839 (N_6839,N_443,N_3485);
and U6840 (N_6840,N_1473,N_1871);
nor U6841 (N_6841,N_3601,N_1539);
nand U6842 (N_6842,N_1204,N_236);
nand U6843 (N_6843,N_3890,N_1125);
nor U6844 (N_6844,N_1085,N_3956);
nand U6845 (N_6845,N_1795,N_218);
or U6846 (N_6846,N_361,N_4118);
nor U6847 (N_6847,N_4795,N_3579);
nor U6848 (N_6848,N_2386,N_634);
and U6849 (N_6849,N_4491,N_3611);
nor U6850 (N_6850,N_3347,N_3625);
and U6851 (N_6851,N_2233,N_2799);
xnor U6852 (N_6852,N_4921,N_152);
or U6853 (N_6853,N_4050,N_3828);
xnor U6854 (N_6854,N_4275,N_3455);
xnor U6855 (N_6855,N_1215,N_1101);
or U6856 (N_6856,N_1649,N_925);
nand U6857 (N_6857,N_3046,N_20);
nand U6858 (N_6858,N_536,N_1801);
nand U6859 (N_6859,N_1828,N_1596);
xnor U6860 (N_6860,N_4333,N_4245);
and U6861 (N_6861,N_2397,N_1559);
xor U6862 (N_6862,N_3829,N_3006);
xnor U6863 (N_6863,N_3487,N_1089);
and U6864 (N_6864,N_683,N_1292);
xor U6865 (N_6865,N_2566,N_650);
or U6866 (N_6866,N_2558,N_1924);
xor U6867 (N_6867,N_579,N_799);
or U6868 (N_6868,N_4479,N_684);
or U6869 (N_6869,N_4703,N_2540);
or U6870 (N_6870,N_3914,N_3229);
or U6871 (N_6871,N_910,N_1627);
nand U6872 (N_6872,N_1544,N_1064);
xor U6873 (N_6873,N_2189,N_4738);
nand U6874 (N_6874,N_3724,N_3831);
nand U6875 (N_6875,N_2419,N_3178);
and U6876 (N_6876,N_1418,N_3144);
xnor U6877 (N_6877,N_2370,N_1272);
or U6878 (N_6878,N_4792,N_2112);
and U6879 (N_6879,N_3449,N_2073);
and U6880 (N_6880,N_4041,N_1274);
and U6881 (N_6881,N_1247,N_3442);
nor U6882 (N_6882,N_541,N_4489);
and U6883 (N_6883,N_4957,N_3893);
nand U6884 (N_6884,N_1631,N_2754);
nor U6885 (N_6885,N_2212,N_244);
or U6886 (N_6886,N_138,N_2776);
nor U6887 (N_6887,N_423,N_3534);
and U6888 (N_6888,N_4159,N_2964);
xnor U6889 (N_6889,N_1045,N_2995);
and U6890 (N_6890,N_4172,N_4096);
nand U6891 (N_6891,N_303,N_3773);
nand U6892 (N_6892,N_3297,N_2341);
or U6893 (N_6893,N_4977,N_610);
and U6894 (N_6894,N_3526,N_4173);
xor U6895 (N_6895,N_2146,N_2902);
nor U6896 (N_6896,N_1788,N_1357);
xnor U6897 (N_6897,N_42,N_767);
nor U6898 (N_6898,N_1369,N_4641);
or U6899 (N_6899,N_3489,N_2686);
nand U6900 (N_6900,N_4612,N_2192);
or U6901 (N_6901,N_1993,N_1669);
and U6902 (N_6902,N_1980,N_2797);
nor U6903 (N_6903,N_975,N_2056);
nand U6904 (N_6904,N_2244,N_1100);
nor U6905 (N_6905,N_1585,N_3758);
or U6906 (N_6906,N_2467,N_4722);
or U6907 (N_6907,N_89,N_4097);
nand U6908 (N_6908,N_3254,N_3577);
or U6909 (N_6909,N_4631,N_4203);
or U6910 (N_6910,N_1918,N_1901);
nand U6911 (N_6911,N_2435,N_102);
and U6912 (N_6912,N_2761,N_232);
xor U6913 (N_6913,N_2572,N_2497);
nand U6914 (N_6914,N_2204,N_1088);
and U6915 (N_6915,N_959,N_4336);
nor U6916 (N_6916,N_3662,N_3336);
nor U6917 (N_6917,N_3141,N_542);
nor U6918 (N_6918,N_1460,N_815);
and U6919 (N_6919,N_3930,N_929);
nand U6920 (N_6920,N_3650,N_1043);
and U6921 (N_6921,N_944,N_4177);
and U6922 (N_6922,N_967,N_157);
nand U6923 (N_6923,N_2084,N_3169);
nor U6924 (N_6924,N_3684,N_2459);
nor U6925 (N_6925,N_779,N_1399);
or U6926 (N_6926,N_4188,N_2155);
nand U6927 (N_6927,N_4661,N_4939);
and U6928 (N_6928,N_3683,N_1478);
nor U6929 (N_6929,N_934,N_1184);
and U6930 (N_6930,N_3509,N_3362);
and U6931 (N_6931,N_2721,N_688);
nand U6932 (N_6932,N_2254,N_1105);
nand U6933 (N_6933,N_4675,N_1723);
nand U6934 (N_6934,N_1727,N_2281);
nor U6935 (N_6935,N_3392,N_3138);
xor U6936 (N_6936,N_4801,N_4818);
or U6937 (N_6937,N_323,N_4916);
xor U6938 (N_6938,N_995,N_1013);
nor U6939 (N_6939,N_336,N_2807);
xnor U6940 (N_6940,N_997,N_3933);
nand U6941 (N_6941,N_4600,N_1830);
nand U6942 (N_6942,N_1885,N_4630);
and U6943 (N_6943,N_1304,N_2082);
xor U6944 (N_6944,N_2393,N_3563);
nor U6945 (N_6945,N_1002,N_2140);
xnor U6946 (N_6946,N_4779,N_435);
xnor U6947 (N_6947,N_3239,N_3740);
nand U6948 (N_6948,N_762,N_2038);
nand U6949 (N_6949,N_4539,N_970);
or U6950 (N_6950,N_3503,N_4820);
xnor U6951 (N_6951,N_475,N_497);
nand U6952 (N_6952,N_3967,N_2584);
and U6953 (N_6953,N_4141,N_905);
xnor U6954 (N_6954,N_2621,N_441);
or U6955 (N_6955,N_3992,N_4000);
or U6956 (N_6956,N_3518,N_4994);
nand U6957 (N_6957,N_2087,N_1495);
xnor U6958 (N_6958,N_4080,N_4143);
and U6959 (N_6959,N_3307,N_804);
or U6960 (N_6960,N_3428,N_3137);
nor U6961 (N_6961,N_1393,N_1378);
nor U6962 (N_6962,N_768,N_1254);
nand U6963 (N_6963,N_3279,N_3079);
or U6964 (N_6964,N_4573,N_642);
and U6965 (N_6965,N_812,N_350);
nand U6966 (N_6966,N_609,N_3589);
and U6967 (N_6967,N_527,N_345);
xor U6968 (N_6968,N_3624,N_2445);
and U6969 (N_6969,N_533,N_1674);
or U6970 (N_6970,N_1201,N_3061);
nand U6971 (N_6971,N_41,N_4766);
nor U6972 (N_6972,N_1345,N_2594);
and U6973 (N_6973,N_3528,N_4857);
or U6974 (N_6974,N_3201,N_1868);
nor U6975 (N_6975,N_3977,N_171);
or U6976 (N_6976,N_2202,N_4633);
and U6977 (N_6977,N_537,N_315);
xnor U6978 (N_6978,N_4883,N_3378);
or U6979 (N_6979,N_1632,N_1103);
nor U6980 (N_6980,N_4176,N_2690);
or U6981 (N_6981,N_385,N_2952);
nand U6982 (N_6982,N_643,N_620);
xor U6983 (N_6983,N_4516,N_1262);
or U6984 (N_6984,N_1380,N_1761);
xnor U6985 (N_6985,N_854,N_3123);
or U6986 (N_6986,N_3062,N_4799);
xnor U6987 (N_6987,N_1410,N_891);
nand U6988 (N_6988,N_380,N_2049);
and U6989 (N_6989,N_3881,N_3259);
and U6990 (N_6990,N_3415,N_3848);
and U6991 (N_6991,N_4211,N_4745);
or U6992 (N_6992,N_2264,N_585);
or U6993 (N_6993,N_490,N_2514);
xor U6994 (N_6994,N_1012,N_427);
and U6995 (N_6995,N_4403,N_381);
or U6996 (N_6996,N_2449,N_170);
nand U6997 (N_6997,N_4166,N_4669);
or U6998 (N_6998,N_255,N_2862);
and U6999 (N_6999,N_4740,N_4413);
and U7000 (N_7000,N_328,N_3545);
nor U7001 (N_7001,N_2214,N_3870);
nand U7002 (N_7002,N_1034,N_3460);
nand U7003 (N_7003,N_2152,N_3365);
xnor U7004 (N_7004,N_1228,N_3647);
or U7005 (N_7005,N_2009,N_1426);
xnor U7006 (N_7006,N_2469,N_3771);
xor U7007 (N_7007,N_1519,N_4058);
nor U7008 (N_7008,N_3156,N_3398);
nand U7009 (N_7009,N_1548,N_48);
nand U7010 (N_7010,N_4341,N_4131);
and U7011 (N_7011,N_1506,N_589);
nor U7012 (N_7012,N_4127,N_3113);
nand U7013 (N_7013,N_4731,N_388);
or U7014 (N_7014,N_1799,N_4642);
and U7015 (N_7015,N_698,N_1745);
nand U7016 (N_7016,N_2876,N_1675);
nand U7017 (N_7017,N_603,N_2345);
xor U7018 (N_7018,N_1517,N_4465);
or U7019 (N_7019,N_114,N_1975);
nor U7020 (N_7020,N_730,N_2582);
or U7021 (N_7021,N_405,N_712);
xnor U7022 (N_7022,N_22,N_3126);
and U7023 (N_7023,N_1238,N_3999);
and U7024 (N_7024,N_2175,N_1601);
xor U7025 (N_7025,N_219,N_261);
or U7026 (N_7026,N_4191,N_4823);
nand U7027 (N_7027,N_3488,N_1836);
xnor U7028 (N_7028,N_7,N_4747);
xor U7029 (N_7029,N_124,N_4145);
nor U7030 (N_7030,N_2757,N_4822);
nand U7031 (N_7031,N_3121,N_62);
nor U7032 (N_7032,N_3321,N_3027);
or U7033 (N_7033,N_4668,N_1388);
xor U7034 (N_7034,N_4657,N_1862);
or U7035 (N_7035,N_1411,N_3966);
and U7036 (N_7036,N_1518,N_4802);
nand U7037 (N_7037,N_3701,N_961);
or U7038 (N_7038,N_3233,N_4676);
nand U7039 (N_7039,N_3951,N_2315);
nor U7040 (N_7040,N_1086,N_2441);
nand U7041 (N_7041,N_1289,N_4209);
nand U7042 (N_7042,N_2829,N_3475);
nor U7043 (N_7043,N_54,N_1044);
or U7044 (N_7044,N_3264,N_2730);
nand U7045 (N_7045,N_2969,N_281);
nand U7046 (N_7046,N_117,N_1104);
and U7047 (N_7047,N_3654,N_2277);
nor U7048 (N_7048,N_1187,N_3819);
xor U7049 (N_7049,N_25,N_3641);
or U7050 (N_7050,N_4059,N_1334);
nor U7051 (N_7051,N_355,N_294);
and U7052 (N_7052,N_3715,N_2402);
nor U7053 (N_7053,N_1747,N_3249);
nand U7054 (N_7054,N_1743,N_3174);
nor U7055 (N_7055,N_887,N_787);
xnor U7056 (N_7056,N_3005,N_3673);
xnor U7057 (N_7057,N_1072,N_176);
and U7058 (N_7058,N_1427,N_3801);
nand U7059 (N_7059,N_2628,N_4756);
or U7060 (N_7060,N_4190,N_3183);
xor U7061 (N_7061,N_4656,N_4528);
nor U7062 (N_7062,N_2561,N_4123);
nor U7063 (N_7063,N_4139,N_1291);
or U7064 (N_7064,N_3824,N_4934);
nor U7065 (N_7065,N_3101,N_3968);
xnor U7066 (N_7066,N_1702,N_1776);
nand U7067 (N_7067,N_1190,N_4015);
xnor U7068 (N_7068,N_3334,N_2856);
xor U7069 (N_7069,N_2627,N_451);
xnor U7070 (N_7070,N_1222,N_3986);
xor U7071 (N_7071,N_1789,N_3566);
xor U7072 (N_7072,N_1298,N_800);
or U7073 (N_7073,N_4101,N_4490);
or U7074 (N_7074,N_1486,N_437);
and U7075 (N_7075,N_2088,N_638);
nor U7076 (N_7076,N_4241,N_2512);
or U7077 (N_7077,N_2157,N_3405);
and U7078 (N_7078,N_2329,N_2749);
or U7079 (N_7079,N_3163,N_2583);
nor U7080 (N_7080,N_398,N_4482);
and U7081 (N_7081,N_3269,N_2351);
nand U7082 (N_7082,N_545,N_3016);
or U7083 (N_7083,N_2228,N_3686);
and U7084 (N_7084,N_3544,N_1856);
xnor U7085 (N_7085,N_3746,N_3324);
nand U7086 (N_7086,N_2117,N_148);
nor U7087 (N_7087,N_2303,N_3822);
or U7088 (N_7088,N_1867,N_621);
nor U7089 (N_7089,N_3036,N_2842);
or U7090 (N_7090,N_1708,N_999);
or U7091 (N_7091,N_2560,N_862);
nand U7092 (N_7092,N_2536,N_4567);
nor U7093 (N_7093,N_2487,N_1625);
xnor U7094 (N_7094,N_930,N_4525);
and U7095 (N_7095,N_4149,N_162);
xnor U7096 (N_7096,N_4320,N_908);
or U7097 (N_7097,N_3232,N_1236);
xor U7098 (N_7098,N_705,N_3610);
nand U7099 (N_7099,N_2805,N_4982);
nand U7100 (N_7100,N_2120,N_1253);
xor U7101 (N_7101,N_36,N_3224);
nand U7102 (N_7102,N_3122,N_3978);
xor U7103 (N_7103,N_4416,N_4504);
nor U7104 (N_7104,N_483,N_864);
nand U7105 (N_7105,N_4423,N_2440);
and U7106 (N_7106,N_2999,N_3739);
and U7107 (N_7107,N_2614,N_4397);
xnor U7108 (N_7108,N_4923,N_1523);
nor U7109 (N_7109,N_3298,N_4827);
xnor U7110 (N_7110,N_239,N_2968);
and U7111 (N_7111,N_1018,N_629);
nor U7112 (N_7112,N_4509,N_3349);
xnor U7113 (N_7113,N_1714,N_817);
nor U7114 (N_7114,N_2702,N_4316);
xnor U7115 (N_7115,N_1942,N_3776);
xor U7116 (N_7116,N_532,N_2552);
and U7117 (N_7117,N_2477,N_990);
and U7118 (N_7118,N_4068,N_2100);
xnor U7119 (N_7119,N_1361,N_4055);
nand U7120 (N_7120,N_1249,N_1020);
and U7121 (N_7121,N_493,N_2521);
and U7122 (N_7122,N_4223,N_3961);
nor U7123 (N_7123,N_3029,N_4773);
nor U7124 (N_7124,N_3605,N_619);
and U7125 (N_7125,N_178,N_2928);
nand U7126 (N_7126,N_1395,N_1744);
and U7127 (N_7127,N_2039,N_331);
nand U7128 (N_7128,N_2408,N_2585);
nand U7129 (N_7129,N_1242,N_4808);
and U7130 (N_7130,N_1508,N_3931);
nand U7131 (N_7131,N_476,N_2016);
or U7132 (N_7132,N_509,N_3582);
and U7133 (N_7133,N_941,N_1219);
nor U7134 (N_7134,N_2944,N_477);
nand U7135 (N_7135,N_4088,N_1516);
nor U7136 (N_7136,N_402,N_2808);
nor U7137 (N_7137,N_1656,N_353);
xor U7138 (N_7138,N_2493,N_3017);
and U7139 (N_7139,N_1282,N_2159);
xnor U7140 (N_7140,N_4678,N_3551);
and U7141 (N_7141,N_1790,N_2632);
xnor U7142 (N_7142,N_4174,N_2960);
and U7143 (N_7143,N_3912,N_3202);
nor U7144 (N_7144,N_2696,N_1624);
xor U7145 (N_7145,N_1970,N_4326);
and U7146 (N_7146,N_3070,N_4394);
xor U7147 (N_7147,N_4011,N_225);
nand U7148 (N_7148,N_795,N_4421);
xnor U7149 (N_7149,N_4021,N_439);
nand U7150 (N_7150,N_1763,N_1414);
xor U7151 (N_7151,N_951,N_2962);
xnor U7152 (N_7152,N_3508,N_4357);
xnor U7153 (N_7153,N_4258,N_4755);
and U7154 (N_7154,N_2553,N_935);
nor U7155 (N_7155,N_2392,N_844);
or U7156 (N_7156,N_1381,N_3155);
nor U7157 (N_7157,N_3480,N_3797);
nand U7158 (N_7158,N_3408,N_1990);
or U7159 (N_7159,N_3685,N_963);
and U7160 (N_7160,N_3530,N_2018);
nand U7161 (N_7161,N_4811,N_3059);
and U7162 (N_7162,N_3904,N_663);
nor U7163 (N_7163,N_2922,N_3241);
nor U7164 (N_7164,N_1638,N_3806);
or U7165 (N_7165,N_1912,N_2311);
nor U7166 (N_7166,N_2915,N_4587);
or U7167 (N_7167,N_932,N_4616);
nor U7168 (N_7168,N_399,N_1305);
nand U7169 (N_7169,N_4547,N_3581);
nand U7170 (N_7170,N_2885,N_4564);
and U7171 (N_7171,N_3010,N_4937);
and U7172 (N_7172,N_574,N_2784);
and U7173 (N_7173,N_2903,N_1681);
xnor U7174 (N_7174,N_4260,N_2447);
or U7175 (N_7175,N_262,N_2366);
or U7176 (N_7176,N_2511,N_4013);
nor U7177 (N_7177,N_786,N_1321);
nor U7178 (N_7178,N_977,N_3037);
or U7179 (N_7179,N_2299,N_4501);
and U7180 (N_7180,N_4598,N_394);
and U7181 (N_7181,N_1014,N_4434);
or U7182 (N_7182,N_4665,N_978);
nor U7183 (N_7183,N_4845,N_3220);
xor U7184 (N_7184,N_3287,N_1280);
or U7185 (N_7185,N_1485,N_3525);
or U7186 (N_7186,N_2111,N_4816);
or U7187 (N_7187,N_2101,N_2959);
or U7188 (N_7188,N_2677,N_1948);
xor U7189 (N_7189,N_132,N_2352);
xor U7190 (N_7190,N_2297,N_1720);
nor U7191 (N_7191,N_4100,N_1687);
nor U7192 (N_7192,N_3880,N_1595);
and U7193 (N_7193,N_2747,N_2);
and U7194 (N_7194,N_3664,N_3127);
and U7195 (N_7195,N_1351,N_1326);
nor U7196 (N_7196,N_1568,N_3322);
and U7197 (N_7197,N_226,N_3002);
or U7198 (N_7198,N_2662,N_491);
or U7199 (N_7199,N_3243,N_268);
nand U7200 (N_7200,N_4281,N_3636);
xor U7201 (N_7201,N_1909,N_530);
and U7202 (N_7202,N_1314,N_2348);
or U7203 (N_7203,N_3730,N_4978);
or U7204 (N_7204,N_1590,N_831);
and U7205 (N_7205,N_1893,N_3255);
xor U7206 (N_7206,N_827,N_4599);
and U7207 (N_7207,N_3335,N_246);
nand U7208 (N_7208,N_1079,N_3598);
xor U7209 (N_7209,N_1461,N_760);
xor U7210 (N_7210,N_3390,N_2953);
and U7211 (N_7211,N_1713,N_257);
nor U7212 (N_7212,N_203,N_310);
nand U7213 (N_7213,N_3231,N_755);
xnor U7214 (N_7214,N_1965,N_1883);
nand U7215 (N_7215,N_2360,N_4193);
xnor U7216 (N_7216,N_4671,N_1889);
nand U7217 (N_7217,N_821,N_44);
nand U7218 (N_7218,N_1454,N_3481);
nor U7219 (N_7219,N_2609,N_1354);
or U7220 (N_7220,N_4750,N_4544);
and U7221 (N_7221,N_2527,N_425);
and U7222 (N_7222,N_1158,N_3000);
xnor U7223 (N_7223,N_3419,N_4859);
nand U7224 (N_7224,N_4047,N_3332);
and U7225 (N_7225,N_1330,N_858);
and U7226 (N_7226,N_4719,N_84);
and U7227 (N_7227,N_3076,N_2539);
xnor U7228 (N_7228,N_825,N_2692);
or U7229 (N_7229,N_3617,N_3014);
nor U7230 (N_7230,N_2288,N_4089);
xor U7231 (N_7231,N_4372,N_1910);
xnor U7232 (N_7232,N_700,N_3878);
nand U7233 (N_7233,N_1211,N_3384);
and U7234 (N_7234,N_914,N_546);
or U7235 (N_7235,N_4231,N_4622);
xor U7236 (N_7236,N_3976,N_3573);
or U7237 (N_7237,N_1283,N_159);
and U7238 (N_7238,N_2027,N_4071);
xor U7239 (N_7239,N_4186,N_4283);
xor U7240 (N_7240,N_552,N_2958);
nor U7241 (N_7241,N_1680,N_2851);
or U7242 (N_7242,N_459,N_1209);
nand U7243 (N_7243,N_2987,N_1825);
or U7244 (N_7244,N_3592,N_21);
nor U7245 (N_7245,N_3688,N_3443);
or U7246 (N_7246,N_2321,N_39);
and U7247 (N_7247,N_4120,N_3054);
xnor U7248 (N_7248,N_3537,N_2134);
nor U7249 (N_7249,N_4133,N_3587);
or U7250 (N_7250,N_2096,N_1915);
and U7251 (N_7251,N_3406,N_2050);
nor U7252 (N_7252,N_2648,N_269);
nor U7253 (N_7253,N_3749,N_3523);
or U7254 (N_7254,N_418,N_4457);
nand U7255 (N_7255,N_1626,N_4637);
xor U7256 (N_7256,N_3171,N_4540);
nor U7257 (N_7257,N_503,N_4903);
xor U7258 (N_7258,N_1533,N_344);
nor U7259 (N_7259,N_853,N_1329);
nand U7260 (N_7260,N_1412,N_1110);
or U7261 (N_7261,N_1017,N_3506);
and U7262 (N_7262,N_2726,N_550);
nand U7263 (N_7263,N_3484,N_3782);
and U7264 (N_7264,N_3767,N_4878);
nor U7265 (N_7265,N_595,N_852);
and U7266 (N_7266,N_1246,N_2538);
xor U7267 (N_7267,N_3841,N_2031);
xor U7268 (N_7268,N_1285,N_943);
nand U7269 (N_7269,N_4221,N_3071);
nand U7270 (N_7270,N_1777,N_40);
xor U7271 (N_7271,N_2002,N_140);
nand U7272 (N_7272,N_3896,N_1837);
and U7273 (N_7273,N_2738,N_3413);
xor U7274 (N_7274,N_202,N_4392);
nand U7275 (N_7275,N_3429,N_3085);
and U7276 (N_7276,N_2410,N_3304);
nand U7277 (N_7277,N_1404,N_3677);
nand U7278 (N_7278,N_337,N_2931);
nand U7279 (N_7279,N_4414,N_664);
xor U7280 (N_7280,N_3708,N_2076);
xnor U7281 (N_7281,N_4070,N_3299);
and U7282 (N_7282,N_3946,N_1906);
or U7283 (N_7283,N_4030,N_432);
nand U7284 (N_7284,N_1462,N_4796);
or U7285 (N_7285,N_55,N_2429);
nor U7286 (N_7286,N_2984,N_1688);
xnor U7287 (N_7287,N_4470,N_319);
and U7288 (N_7288,N_962,N_1716);
and U7289 (N_7289,N_1521,N_2498);
xor U7290 (N_7290,N_3542,N_4843);
nand U7291 (N_7291,N_1594,N_3539);
or U7292 (N_7292,N_758,N_4938);
nor U7293 (N_7293,N_1935,N_1128);
or U7294 (N_7294,N_4919,N_1183);
xor U7295 (N_7295,N_3438,N_2376);
or U7296 (N_7296,N_164,N_1421);
or U7297 (N_7297,N_2223,N_3628);
nor U7298 (N_7298,N_2148,N_4105);
nand U7299 (N_7299,N_502,N_4390);
nor U7300 (N_7300,N_3033,N_2261);
and U7301 (N_7301,N_4012,N_4850);
and U7302 (N_7302,N_2097,N_564);
and U7303 (N_7303,N_272,N_2225);
nand U7304 (N_7304,N_4415,N_2269);
or U7305 (N_7305,N_4474,N_4436);
or U7306 (N_7306,N_4034,N_3325);
nor U7307 (N_7307,N_30,N_2942);
nand U7308 (N_7308,N_4986,N_3706);
or U7309 (N_7309,N_4148,N_4914);
xnor U7310 (N_7310,N_1026,N_279);
nor U7311 (N_7311,N_1709,N_1555);
nor U7312 (N_7312,N_803,N_471);
nor U7313 (N_7313,N_4711,N_3301);
nand U7314 (N_7314,N_4561,N_3073);
or U7315 (N_7315,N_2460,N_4945);
or U7316 (N_7316,N_2331,N_4324);
nand U7317 (N_7317,N_4658,N_1068);
nor U7318 (N_7318,N_2814,N_1050);
nor U7319 (N_7319,N_3524,N_4915);
nand U7320 (N_7320,N_704,N_4523);
nand U7321 (N_7321,N_1458,N_3632);
xor U7322 (N_7322,N_3402,N_556);
xor U7323 (N_7323,N_2102,N_3153);
nand U7324 (N_7324,N_1951,N_4130);
nor U7325 (N_7325,N_2322,N_3018);
or U7326 (N_7326,N_2384,N_60);
and U7327 (N_7327,N_4227,N_2409);
nor U7328 (N_7328,N_613,N_902);
xnor U7329 (N_7329,N_2201,N_2678);
nand U7330 (N_7330,N_933,N_985);
or U7331 (N_7331,N_741,N_2320);
nand U7332 (N_7332,N_2465,N_3578);
or U7333 (N_7333,N_387,N_763);
and U7334 (N_7334,N_3424,N_1006);
or U7335 (N_7335,N_120,N_4140);
nor U7336 (N_7336,N_1106,N_2012);
nor U7337 (N_7337,N_2719,N_573);
and U7338 (N_7338,N_15,N_780);
or U7339 (N_7339,N_2400,N_1802);
xor U7340 (N_7340,N_2124,N_4901);
nand U7341 (N_7341,N_4858,N_115);
xnor U7342 (N_7342,N_3692,N_826);
nand U7343 (N_7343,N_2581,N_4183);
and U7344 (N_7344,N_2502,N_625);
nand U7345 (N_7345,N_3833,N_2823);
nand U7346 (N_7346,N_1969,N_4175);
nand U7347 (N_7347,N_1697,N_229);
nand U7348 (N_7348,N_3237,N_1300);
nand U7349 (N_7349,N_1197,N_4334);
nand U7350 (N_7350,N_1840,N_2989);
nand U7351 (N_7351,N_2597,N_1057);
nand U7352 (N_7352,N_2438,N_325);
or U7353 (N_7353,N_3296,N_2668);
xnor U7354 (N_7354,N_499,N_4314);
or U7355 (N_7355,N_1299,N_614);
nor U7356 (N_7356,N_4308,N_1116);
nor U7357 (N_7357,N_4406,N_146);
nand U7358 (N_7358,N_2711,N_1654);
or U7359 (N_7359,N_3108,N_4265);
xnor U7360 (N_7360,N_1666,N_3289);
and U7361 (N_7361,N_4469,N_968);
and U7362 (N_7362,N_247,N_24);
xor U7363 (N_7363,N_4358,N_1532);
nand U7364 (N_7364,N_234,N_4461);
and U7365 (N_7365,N_3675,N_4590);
nand U7366 (N_7366,N_4290,N_1065);
xnor U7367 (N_7367,N_3656,N_4113);
or U7368 (N_7368,N_3084,N_4716);
nand U7369 (N_7369,N_3366,N_829);
and U7370 (N_7370,N_151,N_2626);
xor U7371 (N_7371,N_3642,N_3072);
xnor U7372 (N_7372,N_3466,N_2841);
nor U7373 (N_7373,N_1373,N_2985);
and U7374 (N_7374,N_1081,N_214);
nand U7375 (N_7375,N_227,N_4905);
or U7376 (N_7376,N_2657,N_1958);
or U7377 (N_7377,N_2936,N_2717);
and U7378 (N_7378,N_3519,N_2998);
nor U7379 (N_7379,N_447,N_321);
xor U7380 (N_7380,N_3256,N_3228);
nand U7381 (N_7381,N_2032,N_2868);
or U7382 (N_7382,N_251,N_2263);
nor U7383 (N_7383,N_526,N_3453);
xnor U7384 (N_7384,N_3863,N_391);
nand U7385 (N_7385,N_1470,N_1095);
and U7386 (N_7386,N_4189,N_657);
or U7387 (N_7387,N_3176,N_1407);
or U7388 (N_7388,N_1875,N_1786);
and U7389 (N_7389,N_3840,N_3319);
or U7390 (N_7390,N_1365,N_2043);
nor U7391 (N_7391,N_1728,N_4748);
nand U7392 (N_7392,N_1498,N_3395);
nor U7393 (N_7393,N_2491,N_3777);
xnor U7394 (N_7394,N_2144,N_2652);
nor U7395 (N_7395,N_4913,N_1046);
nor U7396 (N_7396,N_4412,N_2825);
or U7397 (N_7397,N_1467,N_3290);
nor U7398 (N_7398,N_3469,N_4168);
or U7399 (N_7399,N_3323,N_4729);
nand U7400 (N_7400,N_4933,N_1732);
nor U7401 (N_7401,N_735,N_3674);
nor U7402 (N_7402,N_2604,N_3182);
nand U7403 (N_7403,N_1784,N_3920);
xor U7404 (N_7404,N_1,N_4607);
and U7405 (N_7405,N_3859,N_3399);
and U7406 (N_7406,N_752,N_1515);
nor U7407 (N_7407,N_4866,N_3557);
or U7408 (N_7408,N_264,N_1765);
nor U7409 (N_7409,N_2305,N_1175);
and U7410 (N_7410,N_3312,N_3769);
and U7411 (N_7411,N_4624,N_1573);
and U7412 (N_7412,N_4497,N_3707);
or U7413 (N_7413,N_1077,N_3456);
and U7414 (N_7414,N_1834,N_4179);
or U7415 (N_7415,N_2451,N_2364);
or U7416 (N_7416,N_2975,N_4840);
xor U7417 (N_7417,N_1752,N_2309);
nor U7418 (N_7418,N_2474,N_2241);
or U7419 (N_7419,N_1349,N_508);
nor U7420 (N_7420,N_2217,N_1905);
nand U7421 (N_7421,N_1120,N_2864);
and U7422 (N_7422,N_1497,N_329);
nand U7423 (N_7423,N_2361,N_4195);
or U7424 (N_7424,N_1449,N_3649);
xnor U7425 (N_7425,N_4363,N_1137);
nor U7426 (N_7426,N_3436,N_2167);
and U7427 (N_7427,N_1016,N_4486);
nand U7428 (N_7428,N_3093,N_551);
nand U7429 (N_7429,N_4686,N_1908);
or U7430 (N_7430,N_1036,N_606);
nor U7431 (N_7431,N_2910,N_1712);
and U7432 (N_7432,N_4927,N_679);
and U7433 (N_7433,N_86,N_4943);
and U7434 (N_7434,N_112,N_1971);
or U7435 (N_7435,N_4110,N_2755);
nand U7436 (N_7436,N_1169,N_2643);
nor U7437 (N_7437,N_1221,N_1756);
nand U7438 (N_7438,N_4887,N_59);
nor U7439 (N_7439,N_4192,N_1075);
nor U7440 (N_7440,N_2694,N_1659);
nand U7441 (N_7441,N_413,N_1164);
xor U7442 (N_7442,N_801,N_3886);
or U7443 (N_7443,N_993,N_2436);
and U7444 (N_7444,N_2935,N_4171);
or U7445 (N_7445,N_1864,N_1607);
and U7446 (N_7446,N_3640,N_3148);
and U7447 (N_7447,N_2848,N_3315);
nand U7448 (N_7448,N_4654,N_2907);
and U7449 (N_7449,N_1229,N_677);
xor U7450 (N_7450,N_2186,N_881);
nor U7451 (N_7451,N_2488,N_192);
xor U7452 (N_7452,N_1303,N_3190);
and U7453 (N_7453,N_1921,N_2741);
xnor U7454 (N_7454,N_2589,N_240);
nor U7455 (N_7455,N_3604,N_1800);
nor U7456 (N_7456,N_2065,N_3023);
and U7457 (N_7457,N_1216,N_1683);
nand U7458 (N_7458,N_637,N_2874);
or U7459 (N_7459,N_2342,N_1504);
or U7460 (N_7460,N_3761,N_2832);
nand U7461 (N_7461,N_2637,N_2550);
xor U7462 (N_7462,N_4429,N_3510);
nand U7463 (N_7463,N_4312,N_1537);
nand U7464 (N_7464,N_3049,N_658);
xnor U7465 (N_7465,N_3433,N_738);
xnor U7466 (N_7466,N_1616,N_4418);
and U7467 (N_7467,N_2579,N_3139);
xor U7468 (N_7468,N_121,N_4204);
or U7469 (N_7469,N_1891,N_208);
or U7470 (N_7470,N_4534,N_4910);
xnor U7471 (N_7471,N_4830,N_979);
or U7472 (N_7472,N_1162,N_1794);
nor U7473 (N_7473,N_2130,N_2595);
nand U7474 (N_7474,N_622,N_71);
xor U7475 (N_7475,N_3432,N_296);
xnor U7476 (N_7476,N_4495,N_1223);
xor U7477 (N_7477,N_4794,N_4466);
nand U7478 (N_7478,N_1946,N_3317);
nor U7479 (N_7479,N_1780,N_3873);
xnor U7480 (N_7480,N_4613,N_2949);
or U7481 (N_7481,N_708,N_3995);
nor U7482 (N_7482,N_4763,N_4010);
nand U7483 (N_7483,N_1417,N_1396);
or U7484 (N_7484,N_1297,N_134);
xor U7485 (N_7485,N_2943,N_4337);
xnor U7486 (N_7486,N_2927,N_2194);
nor U7487 (N_7487,N_3879,N_2068);
or U7488 (N_7488,N_1337,N_4370);
and U7489 (N_7489,N_2109,N_1919);
or U7490 (N_7490,N_1660,N_3574);
nor U7491 (N_7491,N_1692,N_1733);
nor U7492 (N_7492,N_3011,N_3559);
nand U7493 (N_7493,N_2744,N_3403);
xor U7494 (N_7494,N_1722,N_4289);
nand U7495 (N_7495,N_982,N_58);
or U7496 (N_7496,N_4323,N_2072);
nand U7497 (N_7497,N_897,N_2060);
nand U7498 (N_7498,N_3839,N_51);
xor U7499 (N_7499,N_4702,N_4147);
nand U7500 (N_7500,N_1561,N_1543);
nand U7501 (N_7501,N_22,N_2417);
or U7502 (N_7502,N_365,N_3984);
nand U7503 (N_7503,N_2991,N_1460);
xor U7504 (N_7504,N_2497,N_85);
and U7505 (N_7505,N_2836,N_2800);
xor U7506 (N_7506,N_4145,N_4373);
and U7507 (N_7507,N_2789,N_4751);
nand U7508 (N_7508,N_820,N_4365);
or U7509 (N_7509,N_536,N_183);
nor U7510 (N_7510,N_198,N_2731);
nor U7511 (N_7511,N_2580,N_3895);
xor U7512 (N_7512,N_422,N_3737);
nand U7513 (N_7513,N_909,N_4957);
or U7514 (N_7514,N_2036,N_1389);
or U7515 (N_7515,N_4125,N_204);
or U7516 (N_7516,N_1133,N_4890);
nand U7517 (N_7517,N_4659,N_823);
nand U7518 (N_7518,N_396,N_3333);
nand U7519 (N_7519,N_2939,N_1886);
or U7520 (N_7520,N_688,N_982);
nor U7521 (N_7521,N_3949,N_2211);
nor U7522 (N_7522,N_4334,N_4202);
xor U7523 (N_7523,N_4701,N_1080);
nor U7524 (N_7524,N_1249,N_2813);
nor U7525 (N_7525,N_4446,N_3663);
nor U7526 (N_7526,N_2854,N_4388);
nor U7527 (N_7527,N_73,N_2664);
xor U7528 (N_7528,N_2341,N_4460);
or U7529 (N_7529,N_1812,N_1434);
and U7530 (N_7530,N_2222,N_102);
or U7531 (N_7531,N_431,N_3749);
xor U7532 (N_7532,N_3913,N_4539);
or U7533 (N_7533,N_915,N_2905);
xnor U7534 (N_7534,N_303,N_4774);
nand U7535 (N_7535,N_4785,N_572);
xor U7536 (N_7536,N_2085,N_1939);
and U7537 (N_7537,N_2932,N_504);
nand U7538 (N_7538,N_1371,N_2086);
or U7539 (N_7539,N_1436,N_186);
nor U7540 (N_7540,N_4815,N_3288);
nor U7541 (N_7541,N_4599,N_1302);
xnor U7542 (N_7542,N_394,N_486);
and U7543 (N_7543,N_2469,N_2384);
xnor U7544 (N_7544,N_3421,N_398);
or U7545 (N_7545,N_949,N_192);
or U7546 (N_7546,N_1691,N_1746);
nor U7547 (N_7547,N_894,N_2839);
nand U7548 (N_7548,N_2299,N_3475);
xor U7549 (N_7549,N_3149,N_3241);
and U7550 (N_7550,N_1263,N_431);
and U7551 (N_7551,N_98,N_3750);
or U7552 (N_7552,N_4665,N_4587);
nand U7553 (N_7553,N_4048,N_3411);
nor U7554 (N_7554,N_3356,N_4567);
and U7555 (N_7555,N_3806,N_3937);
nand U7556 (N_7556,N_1428,N_1800);
or U7557 (N_7557,N_109,N_1975);
nand U7558 (N_7558,N_4879,N_115);
xor U7559 (N_7559,N_2815,N_2319);
and U7560 (N_7560,N_1504,N_1676);
xnor U7561 (N_7561,N_3837,N_426);
xor U7562 (N_7562,N_3524,N_1499);
and U7563 (N_7563,N_787,N_2906);
nor U7564 (N_7564,N_297,N_1586);
or U7565 (N_7565,N_2593,N_42);
or U7566 (N_7566,N_4080,N_2309);
or U7567 (N_7567,N_2569,N_1976);
nand U7568 (N_7568,N_529,N_3767);
or U7569 (N_7569,N_1648,N_4600);
nand U7570 (N_7570,N_810,N_3193);
nor U7571 (N_7571,N_3527,N_4954);
nor U7572 (N_7572,N_3677,N_4316);
nor U7573 (N_7573,N_988,N_3168);
and U7574 (N_7574,N_599,N_1535);
or U7575 (N_7575,N_2401,N_3138);
xnor U7576 (N_7576,N_3159,N_1181);
and U7577 (N_7577,N_1544,N_1486);
nand U7578 (N_7578,N_2792,N_178);
or U7579 (N_7579,N_3607,N_3000);
and U7580 (N_7580,N_3623,N_4543);
or U7581 (N_7581,N_4699,N_2184);
and U7582 (N_7582,N_3110,N_4854);
or U7583 (N_7583,N_2997,N_2810);
xnor U7584 (N_7584,N_2030,N_2112);
and U7585 (N_7585,N_4536,N_1053);
xnor U7586 (N_7586,N_4632,N_3119);
nor U7587 (N_7587,N_2164,N_1761);
and U7588 (N_7588,N_1982,N_1600);
nand U7589 (N_7589,N_3599,N_3059);
nand U7590 (N_7590,N_2428,N_164);
and U7591 (N_7591,N_1226,N_2314);
xor U7592 (N_7592,N_3274,N_3752);
nor U7593 (N_7593,N_3201,N_641);
nand U7594 (N_7594,N_1334,N_4083);
or U7595 (N_7595,N_1188,N_1046);
nand U7596 (N_7596,N_834,N_811);
xor U7597 (N_7597,N_1185,N_288);
nand U7598 (N_7598,N_736,N_4456);
or U7599 (N_7599,N_1640,N_3799);
xor U7600 (N_7600,N_1957,N_1323);
xnor U7601 (N_7601,N_2507,N_1168);
xor U7602 (N_7602,N_2004,N_4886);
or U7603 (N_7603,N_958,N_3426);
xor U7604 (N_7604,N_3772,N_1587);
and U7605 (N_7605,N_3133,N_3440);
or U7606 (N_7606,N_695,N_967);
nand U7607 (N_7607,N_1476,N_3581);
or U7608 (N_7608,N_2889,N_522);
nand U7609 (N_7609,N_1217,N_111);
or U7610 (N_7610,N_649,N_2785);
xnor U7611 (N_7611,N_302,N_2901);
nor U7612 (N_7612,N_1677,N_3989);
or U7613 (N_7613,N_3758,N_1915);
nor U7614 (N_7614,N_2368,N_2480);
nand U7615 (N_7615,N_2128,N_1328);
or U7616 (N_7616,N_4519,N_4974);
nand U7617 (N_7617,N_4664,N_3135);
and U7618 (N_7618,N_2934,N_4627);
nor U7619 (N_7619,N_1518,N_1420);
or U7620 (N_7620,N_3136,N_2725);
xnor U7621 (N_7621,N_3365,N_2096);
nor U7622 (N_7622,N_1332,N_3767);
or U7623 (N_7623,N_2927,N_1277);
nor U7624 (N_7624,N_4928,N_3641);
nand U7625 (N_7625,N_1739,N_19);
or U7626 (N_7626,N_3048,N_3882);
nand U7627 (N_7627,N_2717,N_484);
or U7628 (N_7628,N_743,N_3311);
and U7629 (N_7629,N_1351,N_3137);
xor U7630 (N_7630,N_2294,N_2482);
or U7631 (N_7631,N_2692,N_595);
xor U7632 (N_7632,N_3856,N_1232);
xor U7633 (N_7633,N_2581,N_4896);
or U7634 (N_7634,N_4035,N_3769);
and U7635 (N_7635,N_4340,N_3627);
and U7636 (N_7636,N_3917,N_2819);
xor U7637 (N_7637,N_2386,N_3669);
xor U7638 (N_7638,N_2970,N_821);
nor U7639 (N_7639,N_4749,N_3984);
xnor U7640 (N_7640,N_4194,N_172);
nor U7641 (N_7641,N_785,N_3449);
nor U7642 (N_7642,N_4577,N_4923);
nand U7643 (N_7643,N_2265,N_474);
nor U7644 (N_7644,N_2592,N_4092);
xor U7645 (N_7645,N_1511,N_4075);
xor U7646 (N_7646,N_2824,N_4009);
or U7647 (N_7647,N_4395,N_3050);
and U7648 (N_7648,N_3730,N_4352);
xor U7649 (N_7649,N_1685,N_1838);
nand U7650 (N_7650,N_1567,N_3443);
and U7651 (N_7651,N_2314,N_1441);
xor U7652 (N_7652,N_1802,N_738);
and U7653 (N_7653,N_4833,N_3343);
or U7654 (N_7654,N_2962,N_4541);
nand U7655 (N_7655,N_3502,N_117);
nand U7656 (N_7656,N_2781,N_1123);
or U7657 (N_7657,N_4736,N_1000);
and U7658 (N_7658,N_4276,N_3342);
or U7659 (N_7659,N_2368,N_3785);
or U7660 (N_7660,N_1245,N_4141);
nand U7661 (N_7661,N_1812,N_1767);
nor U7662 (N_7662,N_3018,N_678);
and U7663 (N_7663,N_1023,N_4606);
nor U7664 (N_7664,N_3871,N_1965);
nor U7665 (N_7665,N_4727,N_1498);
xnor U7666 (N_7666,N_2940,N_3317);
nor U7667 (N_7667,N_2688,N_1618);
nand U7668 (N_7668,N_2086,N_1976);
and U7669 (N_7669,N_578,N_1089);
nor U7670 (N_7670,N_350,N_2603);
xor U7671 (N_7671,N_836,N_1955);
xor U7672 (N_7672,N_157,N_2061);
and U7673 (N_7673,N_301,N_162);
or U7674 (N_7674,N_4312,N_2193);
or U7675 (N_7675,N_4558,N_3788);
or U7676 (N_7676,N_424,N_3756);
nand U7677 (N_7677,N_1469,N_4765);
and U7678 (N_7678,N_461,N_3626);
xor U7679 (N_7679,N_1486,N_4749);
nand U7680 (N_7680,N_1415,N_3084);
or U7681 (N_7681,N_2551,N_4844);
nor U7682 (N_7682,N_3722,N_3289);
nand U7683 (N_7683,N_2847,N_3018);
xor U7684 (N_7684,N_1231,N_1027);
nor U7685 (N_7685,N_2465,N_2883);
nor U7686 (N_7686,N_2032,N_4291);
xor U7687 (N_7687,N_1147,N_3355);
and U7688 (N_7688,N_243,N_1586);
nand U7689 (N_7689,N_2398,N_1212);
and U7690 (N_7690,N_81,N_3713);
and U7691 (N_7691,N_3252,N_4449);
xnor U7692 (N_7692,N_3592,N_2137);
or U7693 (N_7693,N_4263,N_2610);
xnor U7694 (N_7694,N_992,N_955);
nand U7695 (N_7695,N_2388,N_31);
xor U7696 (N_7696,N_4311,N_1518);
nor U7697 (N_7697,N_4346,N_1008);
nand U7698 (N_7698,N_3215,N_4458);
or U7699 (N_7699,N_4318,N_1532);
xor U7700 (N_7700,N_4154,N_105);
xnor U7701 (N_7701,N_343,N_4091);
nor U7702 (N_7702,N_686,N_279);
nand U7703 (N_7703,N_471,N_543);
nor U7704 (N_7704,N_1133,N_1602);
or U7705 (N_7705,N_3289,N_556);
xor U7706 (N_7706,N_3843,N_1527);
xor U7707 (N_7707,N_2295,N_240);
or U7708 (N_7708,N_1341,N_4307);
nand U7709 (N_7709,N_1987,N_3394);
nor U7710 (N_7710,N_2180,N_3519);
and U7711 (N_7711,N_3252,N_1858);
xnor U7712 (N_7712,N_3801,N_425);
xor U7713 (N_7713,N_3818,N_4749);
nor U7714 (N_7714,N_4227,N_2108);
or U7715 (N_7715,N_4050,N_2602);
nor U7716 (N_7716,N_442,N_2646);
or U7717 (N_7717,N_1600,N_2582);
or U7718 (N_7718,N_1108,N_4227);
or U7719 (N_7719,N_4873,N_1647);
nand U7720 (N_7720,N_3097,N_2521);
and U7721 (N_7721,N_2233,N_3833);
and U7722 (N_7722,N_276,N_2135);
nor U7723 (N_7723,N_4859,N_2906);
or U7724 (N_7724,N_3021,N_3343);
xnor U7725 (N_7725,N_984,N_3773);
xnor U7726 (N_7726,N_217,N_4138);
or U7727 (N_7727,N_1683,N_535);
nor U7728 (N_7728,N_4876,N_911);
nand U7729 (N_7729,N_3246,N_184);
and U7730 (N_7730,N_1458,N_4484);
or U7731 (N_7731,N_869,N_307);
nor U7732 (N_7732,N_2290,N_2751);
nor U7733 (N_7733,N_4008,N_4655);
and U7734 (N_7734,N_2642,N_2120);
and U7735 (N_7735,N_3571,N_2188);
xor U7736 (N_7736,N_4314,N_3404);
xnor U7737 (N_7737,N_4964,N_1270);
and U7738 (N_7738,N_2168,N_1416);
xor U7739 (N_7739,N_1802,N_1729);
xor U7740 (N_7740,N_253,N_645);
xor U7741 (N_7741,N_1377,N_2764);
or U7742 (N_7742,N_2356,N_1360);
nand U7743 (N_7743,N_1482,N_1971);
nand U7744 (N_7744,N_4032,N_63);
nor U7745 (N_7745,N_1459,N_156);
xor U7746 (N_7746,N_3721,N_4593);
nor U7747 (N_7747,N_2741,N_3322);
or U7748 (N_7748,N_1014,N_4780);
nand U7749 (N_7749,N_1113,N_3453);
nor U7750 (N_7750,N_2541,N_1840);
and U7751 (N_7751,N_3396,N_4266);
and U7752 (N_7752,N_4519,N_2676);
and U7753 (N_7753,N_710,N_3831);
nor U7754 (N_7754,N_4523,N_3581);
nor U7755 (N_7755,N_743,N_2997);
nand U7756 (N_7756,N_1011,N_2757);
nand U7757 (N_7757,N_4446,N_3874);
or U7758 (N_7758,N_685,N_2669);
xnor U7759 (N_7759,N_4115,N_3503);
nand U7760 (N_7760,N_4844,N_2028);
and U7761 (N_7761,N_3277,N_2611);
and U7762 (N_7762,N_1576,N_3312);
nand U7763 (N_7763,N_788,N_1669);
xor U7764 (N_7764,N_702,N_2729);
or U7765 (N_7765,N_395,N_4291);
nand U7766 (N_7766,N_849,N_1674);
xnor U7767 (N_7767,N_3038,N_2189);
or U7768 (N_7768,N_1174,N_3528);
nor U7769 (N_7769,N_4777,N_2794);
nand U7770 (N_7770,N_1313,N_1677);
or U7771 (N_7771,N_420,N_4600);
or U7772 (N_7772,N_1278,N_4139);
and U7773 (N_7773,N_4488,N_3742);
nand U7774 (N_7774,N_4756,N_994);
and U7775 (N_7775,N_1107,N_2319);
or U7776 (N_7776,N_1508,N_3930);
nor U7777 (N_7777,N_4293,N_763);
or U7778 (N_7778,N_2366,N_4173);
xor U7779 (N_7779,N_637,N_3335);
nand U7780 (N_7780,N_246,N_1804);
nand U7781 (N_7781,N_4068,N_2270);
xor U7782 (N_7782,N_2272,N_1162);
nand U7783 (N_7783,N_2979,N_4691);
nand U7784 (N_7784,N_682,N_1300);
and U7785 (N_7785,N_4603,N_3154);
nand U7786 (N_7786,N_448,N_2501);
and U7787 (N_7787,N_4178,N_460);
nor U7788 (N_7788,N_2883,N_569);
xor U7789 (N_7789,N_3363,N_1796);
nor U7790 (N_7790,N_1253,N_2473);
or U7791 (N_7791,N_1684,N_2448);
nor U7792 (N_7792,N_3968,N_2105);
or U7793 (N_7793,N_2835,N_4234);
nand U7794 (N_7794,N_1968,N_2485);
or U7795 (N_7795,N_902,N_2316);
and U7796 (N_7796,N_2001,N_750);
nand U7797 (N_7797,N_4859,N_2152);
nor U7798 (N_7798,N_181,N_4611);
nand U7799 (N_7799,N_1928,N_1562);
nand U7800 (N_7800,N_4375,N_3369);
and U7801 (N_7801,N_1078,N_4147);
or U7802 (N_7802,N_3726,N_1307);
nand U7803 (N_7803,N_3706,N_4436);
nand U7804 (N_7804,N_202,N_4032);
xor U7805 (N_7805,N_1067,N_1810);
nor U7806 (N_7806,N_4721,N_283);
and U7807 (N_7807,N_4194,N_3908);
nor U7808 (N_7808,N_739,N_15);
or U7809 (N_7809,N_2330,N_3288);
or U7810 (N_7810,N_2834,N_4430);
nor U7811 (N_7811,N_4468,N_4332);
nor U7812 (N_7812,N_1880,N_634);
nand U7813 (N_7813,N_3957,N_2948);
nand U7814 (N_7814,N_180,N_218);
xor U7815 (N_7815,N_2471,N_2410);
or U7816 (N_7816,N_3586,N_3423);
nor U7817 (N_7817,N_1092,N_1659);
and U7818 (N_7818,N_3001,N_4297);
nor U7819 (N_7819,N_853,N_707);
or U7820 (N_7820,N_2944,N_1902);
nor U7821 (N_7821,N_3801,N_4779);
nor U7822 (N_7822,N_65,N_1990);
or U7823 (N_7823,N_4144,N_2385);
and U7824 (N_7824,N_4200,N_2836);
nand U7825 (N_7825,N_4357,N_146);
and U7826 (N_7826,N_3215,N_316);
nor U7827 (N_7827,N_416,N_4297);
xnor U7828 (N_7828,N_2441,N_659);
xor U7829 (N_7829,N_3,N_1041);
and U7830 (N_7830,N_283,N_1868);
nor U7831 (N_7831,N_4630,N_4277);
or U7832 (N_7832,N_4178,N_4691);
or U7833 (N_7833,N_4022,N_3925);
or U7834 (N_7834,N_3490,N_475);
nand U7835 (N_7835,N_1713,N_1747);
nand U7836 (N_7836,N_2787,N_2251);
or U7837 (N_7837,N_3671,N_3545);
nand U7838 (N_7838,N_1657,N_4566);
nand U7839 (N_7839,N_473,N_3887);
nand U7840 (N_7840,N_770,N_417);
or U7841 (N_7841,N_1450,N_3676);
xnor U7842 (N_7842,N_3715,N_2673);
xor U7843 (N_7843,N_2052,N_2109);
xnor U7844 (N_7844,N_4860,N_1415);
xnor U7845 (N_7845,N_4033,N_3765);
and U7846 (N_7846,N_2520,N_2131);
nand U7847 (N_7847,N_2487,N_3000);
or U7848 (N_7848,N_1182,N_4547);
nor U7849 (N_7849,N_4337,N_377);
and U7850 (N_7850,N_905,N_462);
nand U7851 (N_7851,N_4138,N_3390);
xor U7852 (N_7852,N_1481,N_3769);
nand U7853 (N_7853,N_4131,N_1793);
xnor U7854 (N_7854,N_789,N_1693);
nand U7855 (N_7855,N_3615,N_1391);
nand U7856 (N_7856,N_789,N_1190);
nor U7857 (N_7857,N_128,N_567);
nand U7858 (N_7858,N_394,N_2478);
xor U7859 (N_7859,N_773,N_263);
or U7860 (N_7860,N_1427,N_2232);
and U7861 (N_7861,N_1572,N_2183);
nand U7862 (N_7862,N_4228,N_414);
or U7863 (N_7863,N_3718,N_2893);
xor U7864 (N_7864,N_907,N_4029);
xnor U7865 (N_7865,N_130,N_2954);
nand U7866 (N_7866,N_346,N_4903);
xnor U7867 (N_7867,N_2174,N_4229);
xor U7868 (N_7868,N_365,N_4604);
nand U7869 (N_7869,N_3061,N_1613);
or U7870 (N_7870,N_986,N_81);
nand U7871 (N_7871,N_383,N_2030);
xor U7872 (N_7872,N_1814,N_2633);
nand U7873 (N_7873,N_4943,N_3380);
and U7874 (N_7874,N_4079,N_4121);
or U7875 (N_7875,N_1457,N_4031);
nand U7876 (N_7876,N_170,N_2859);
and U7877 (N_7877,N_1988,N_4903);
and U7878 (N_7878,N_193,N_470);
nand U7879 (N_7879,N_680,N_3301);
and U7880 (N_7880,N_2611,N_3207);
nor U7881 (N_7881,N_3297,N_1866);
xor U7882 (N_7882,N_2526,N_322);
or U7883 (N_7883,N_766,N_1934);
and U7884 (N_7884,N_1072,N_908);
xnor U7885 (N_7885,N_3548,N_709);
xor U7886 (N_7886,N_4697,N_4165);
xor U7887 (N_7887,N_4096,N_3771);
xnor U7888 (N_7888,N_2160,N_4377);
xnor U7889 (N_7889,N_1880,N_357);
or U7890 (N_7890,N_277,N_4457);
nand U7891 (N_7891,N_3465,N_1152);
nor U7892 (N_7892,N_3250,N_3083);
or U7893 (N_7893,N_3901,N_1088);
and U7894 (N_7894,N_3116,N_3312);
and U7895 (N_7895,N_550,N_2074);
nand U7896 (N_7896,N_3755,N_1535);
or U7897 (N_7897,N_3828,N_1322);
or U7898 (N_7898,N_363,N_4396);
xnor U7899 (N_7899,N_3309,N_2295);
or U7900 (N_7900,N_3376,N_2275);
nand U7901 (N_7901,N_3525,N_3386);
nand U7902 (N_7902,N_4004,N_1775);
xor U7903 (N_7903,N_793,N_3110);
nand U7904 (N_7904,N_282,N_2334);
and U7905 (N_7905,N_3259,N_2891);
nand U7906 (N_7906,N_4017,N_2765);
or U7907 (N_7907,N_2444,N_1812);
nor U7908 (N_7908,N_1212,N_2848);
and U7909 (N_7909,N_2253,N_2118);
xnor U7910 (N_7910,N_2302,N_4580);
xor U7911 (N_7911,N_1837,N_4432);
nor U7912 (N_7912,N_875,N_627);
and U7913 (N_7913,N_3304,N_2124);
and U7914 (N_7914,N_2952,N_2874);
or U7915 (N_7915,N_2649,N_2931);
xnor U7916 (N_7916,N_600,N_3565);
xnor U7917 (N_7917,N_227,N_1726);
or U7918 (N_7918,N_4520,N_2805);
and U7919 (N_7919,N_2282,N_21);
or U7920 (N_7920,N_4477,N_129);
nand U7921 (N_7921,N_1716,N_2138);
and U7922 (N_7922,N_3612,N_3539);
xnor U7923 (N_7923,N_802,N_3144);
and U7924 (N_7924,N_3430,N_1968);
nor U7925 (N_7925,N_3032,N_2439);
or U7926 (N_7926,N_2200,N_2672);
or U7927 (N_7927,N_2596,N_4129);
xor U7928 (N_7928,N_4882,N_129);
nand U7929 (N_7929,N_3472,N_2436);
and U7930 (N_7930,N_831,N_2399);
xor U7931 (N_7931,N_1906,N_3757);
and U7932 (N_7932,N_1710,N_3674);
xor U7933 (N_7933,N_812,N_1992);
or U7934 (N_7934,N_3164,N_4795);
or U7935 (N_7935,N_4498,N_200);
or U7936 (N_7936,N_3645,N_4656);
and U7937 (N_7937,N_1788,N_4533);
xor U7938 (N_7938,N_2757,N_1122);
xor U7939 (N_7939,N_825,N_605);
or U7940 (N_7940,N_4384,N_3553);
nand U7941 (N_7941,N_1794,N_287);
or U7942 (N_7942,N_3783,N_1658);
xnor U7943 (N_7943,N_1985,N_4347);
and U7944 (N_7944,N_4942,N_2645);
nor U7945 (N_7945,N_95,N_4757);
and U7946 (N_7946,N_3150,N_3267);
xnor U7947 (N_7947,N_2816,N_1162);
xor U7948 (N_7948,N_878,N_2596);
xor U7949 (N_7949,N_4825,N_4369);
nand U7950 (N_7950,N_4147,N_3745);
or U7951 (N_7951,N_4092,N_2560);
xor U7952 (N_7952,N_1217,N_3630);
nor U7953 (N_7953,N_114,N_1266);
nor U7954 (N_7954,N_2665,N_2649);
nand U7955 (N_7955,N_3858,N_4456);
nand U7956 (N_7956,N_4263,N_4057);
xor U7957 (N_7957,N_4507,N_580);
and U7958 (N_7958,N_1990,N_4392);
or U7959 (N_7959,N_1579,N_3221);
or U7960 (N_7960,N_1876,N_330);
and U7961 (N_7961,N_2961,N_1711);
and U7962 (N_7962,N_3286,N_3542);
nor U7963 (N_7963,N_3641,N_406);
xor U7964 (N_7964,N_1438,N_629);
and U7965 (N_7965,N_3585,N_1825);
and U7966 (N_7966,N_1474,N_269);
nand U7967 (N_7967,N_1840,N_4146);
or U7968 (N_7968,N_3109,N_3803);
nor U7969 (N_7969,N_1465,N_4906);
or U7970 (N_7970,N_726,N_1048);
and U7971 (N_7971,N_439,N_2064);
xnor U7972 (N_7972,N_2719,N_1395);
or U7973 (N_7973,N_1139,N_4034);
nor U7974 (N_7974,N_1670,N_229);
or U7975 (N_7975,N_3516,N_459);
nor U7976 (N_7976,N_1081,N_4068);
and U7977 (N_7977,N_4771,N_4084);
or U7978 (N_7978,N_4867,N_2469);
and U7979 (N_7979,N_3335,N_2056);
and U7980 (N_7980,N_2181,N_3366);
and U7981 (N_7981,N_3065,N_2459);
nand U7982 (N_7982,N_4935,N_3213);
and U7983 (N_7983,N_987,N_3466);
or U7984 (N_7984,N_1882,N_3017);
and U7985 (N_7985,N_1157,N_4864);
nand U7986 (N_7986,N_4377,N_2156);
xnor U7987 (N_7987,N_1089,N_1228);
nand U7988 (N_7988,N_4306,N_528);
and U7989 (N_7989,N_4458,N_2327);
nor U7990 (N_7990,N_2342,N_3037);
or U7991 (N_7991,N_1493,N_2902);
xor U7992 (N_7992,N_3026,N_4383);
xor U7993 (N_7993,N_4916,N_3094);
xnor U7994 (N_7994,N_445,N_1700);
or U7995 (N_7995,N_1288,N_3354);
nand U7996 (N_7996,N_925,N_1343);
and U7997 (N_7997,N_2256,N_3886);
nand U7998 (N_7998,N_3780,N_1362);
nor U7999 (N_7999,N_3848,N_1660);
nand U8000 (N_8000,N_963,N_395);
and U8001 (N_8001,N_4991,N_3336);
and U8002 (N_8002,N_4405,N_155);
nor U8003 (N_8003,N_3881,N_2344);
or U8004 (N_8004,N_4497,N_601);
nand U8005 (N_8005,N_4309,N_2478);
or U8006 (N_8006,N_1459,N_3724);
or U8007 (N_8007,N_494,N_2843);
and U8008 (N_8008,N_1559,N_1378);
and U8009 (N_8009,N_3522,N_1518);
and U8010 (N_8010,N_1198,N_2583);
nor U8011 (N_8011,N_3316,N_1751);
and U8012 (N_8012,N_308,N_4789);
xor U8013 (N_8013,N_4092,N_3969);
nor U8014 (N_8014,N_4906,N_1912);
nor U8015 (N_8015,N_4793,N_4677);
and U8016 (N_8016,N_3955,N_3184);
nor U8017 (N_8017,N_3468,N_4114);
nor U8018 (N_8018,N_2375,N_973);
nor U8019 (N_8019,N_868,N_444);
nand U8020 (N_8020,N_4359,N_2044);
and U8021 (N_8021,N_2524,N_1795);
xnor U8022 (N_8022,N_957,N_512);
xor U8023 (N_8023,N_1650,N_4260);
nand U8024 (N_8024,N_448,N_1287);
or U8025 (N_8025,N_4930,N_2135);
nor U8026 (N_8026,N_3951,N_1039);
nand U8027 (N_8027,N_3500,N_2006);
nor U8028 (N_8028,N_3567,N_1833);
nor U8029 (N_8029,N_3076,N_4891);
or U8030 (N_8030,N_100,N_2588);
xnor U8031 (N_8031,N_2688,N_1938);
nand U8032 (N_8032,N_2396,N_4514);
nor U8033 (N_8033,N_1341,N_1374);
nand U8034 (N_8034,N_316,N_4140);
and U8035 (N_8035,N_4378,N_4468);
nand U8036 (N_8036,N_2718,N_4830);
nand U8037 (N_8037,N_3172,N_1792);
xor U8038 (N_8038,N_4317,N_1521);
nor U8039 (N_8039,N_2673,N_2260);
xnor U8040 (N_8040,N_3743,N_1134);
xnor U8041 (N_8041,N_3536,N_1382);
nand U8042 (N_8042,N_1688,N_2125);
nor U8043 (N_8043,N_3751,N_4149);
nor U8044 (N_8044,N_4400,N_1627);
xnor U8045 (N_8045,N_4243,N_4482);
xor U8046 (N_8046,N_64,N_4122);
or U8047 (N_8047,N_1121,N_3521);
or U8048 (N_8048,N_1123,N_2559);
xor U8049 (N_8049,N_4705,N_2642);
and U8050 (N_8050,N_86,N_1448);
nor U8051 (N_8051,N_120,N_1066);
xnor U8052 (N_8052,N_328,N_2260);
xnor U8053 (N_8053,N_2611,N_3484);
and U8054 (N_8054,N_4302,N_871);
nor U8055 (N_8055,N_1384,N_3891);
or U8056 (N_8056,N_4526,N_4645);
nor U8057 (N_8057,N_342,N_1312);
and U8058 (N_8058,N_3232,N_4894);
and U8059 (N_8059,N_2336,N_1734);
and U8060 (N_8060,N_648,N_88);
nand U8061 (N_8061,N_4131,N_3191);
and U8062 (N_8062,N_2907,N_4084);
nor U8063 (N_8063,N_4295,N_3220);
and U8064 (N_8064,N_4307,N_1406);
or U8065 (N_8065,N_1174,N_3580);
nand U8066 (N_8066,N_2132,N_2806);
or U8067 (N_8067,N_3638,N_3916);
and U8068 (N_8068,N_2353,N_3001);
or U8069 (N_8069,N_3651,N_945);
xnor U8070 (N_8070,N_3890,N_3579);
nor U8071 (N_8071,N_1886,N_4122);
or U8072 (N_8072,N_3726,N_1463);
or U8073 (N_8073,N_398,N_130);
and U8074 (N_8074,N_2877,N_4536);
or U8075 (N_8075,N_3802,N_4332);
xnor U8076 (N_8076,N_1664,N_2609);
nand U8077 (N_8077,N_2459,N_1370);
nor U8078 (N_8078,N_321,N_1402);
nor U8079 (N_8079,N_69,N_904);
and U8080 (N_8080,N_167,N_1270);
or U8081 (N_8081,N_2946,N_969);
or U8082 (N_8082,N_4130,N_2801);
nor U8083 (N_8083,N_3623,N_4093);
nand U8084 (N_8084,N_1268,N_1850);
nand U8085 (N_8085,N_3776,N_3036);
and U8086 (N_8086,N_2287,N_4525);
xor U8087 (N_8087,N_644,N_2879);
nor U8088 (N_8088,N_2342,N_3101);
or U8089 (N_8089,N_838,N_620);
nand U8090 (N_8090,N_519,N_2132);
nor U8091 (N_8091,N_4333,N_2864);
xor U8092 (N_8092,N_1017,N_874);
nand U8093 (N_8093,N_3811,N_2720);
nand U8094 (N_8094,N_3888,N_743);
xnor U8095 (N_8095,N_3484,N_1755);
or U8096 (N_8096,N_1978,N_520);
xor U8097 (N_8097,N_495,N_1809);
nor U8098 (N_8098,N_4746,N_4672);
or U8099 (N_8099,N_4708,N_1117);
nand U8100 (N_8100,N_1467,N_2986);
nor U8101 (N_8101,N_2133,N_624);
xnor U8102 (N_8102,N_804,N_1953);
and U8103 (N_8103,N_2013,N_3471);
and U8104 (N_8104,N_3710,N_2334);
xnor U8105 (N_8105,N_3386,N_4292);
xor U8106 (N_8106,N_2634,N_2243);
or U8107 (N_8107,N_2376,N_3105);
or U8108 (N_8108,N_4689,N_1084);
nor U8109 (N_8109,N_173,N_1051);
or U8110 (N_8110,N_286,N_2567);
nand U8111 (N_8111,N_4130,N_3351);
and U8112 (N_8112,N_1108,N_4316);
or U8113 (N_8113,N_1340,N_1456);
or U8114 (N_8114,N_474,N_3718);
xnor U8115 (N_8115,N_4045,N_3848);
and U8116 (N_8116,N_1487,N_2677);
and U8117 (N_8117,N_4418,N_3161);
or U8118 (N_8118,N_3628,N_4587);
and U8119 (N_8119,N_3108,N_4036);
and U8120 (N_8120,N_2088,N_4240);
xor U8121 (N_8121,N_3317,N_3351);
nor U8122 (N_8122,N_4010,N_4720);
xor U8123 (N_8123,N_2073,N_2029);
or U8124 (N_8124,N_1584,N_3299);
nand U8125 (N_8125,N_632,N_4675);
or U8126 (N_8126,N_4336,N_3451);
xor U8127 (N_8127,N_4118,N_3418);
and U8128 (N_8128,N_2572,N_1882);
nor U8129 (N_8129,N_4660,N_2109);
or U8130 (N_8130,N_2886,N_1195);
or U8131 (N_8131,N_1071,N_4962);
xor U8132 (N_8132,N_3453,N_3688);
xnor U8133 (N_8133,N_3378,N_3044);
or U8134 (N_8134,N_1872,N_4245);
nor U8135 (N_8135,N_1251,N_764);
nor U8136 (N_8136,N_4057,N_2184);
xnor U8137 (N_8137,N_775,N_4267);
or U8138 (N_8138,N_1888,N_1913);
xor U8139 (N_8139,N_3147,N_3160);
or U8140 (N_8140,N_2441,N_1254);
nor U8141 (N_8141,N_3601,N_1407);
nand U8142 (N_8142,N_630,N_2109);
xnor U8143 (N_8143,N_4037,N_1818);
or U8144 (N_8144,N_2129,N_300);
or U8145 (N_8145,N_1330,N_3323);
nand U8146 (N_8146,N_3757,N_704);
nor U8147 (N_8147,N_4321,N_3193);
nand U8148 (N_8148,N_2827,N_2366);
nand U8149 (N_8149,N_545,N_344);
and U8150 (N_8150,N_3607,N_1065);
nand U8151 (N_8151,N_898,N_1361);
or U8152 (N_8152,N_3834,N_719);
nand U8153 (N_8153,N_2014,N_3254);
nand U8154 (N_8154,N_447,N_4620);
or U8155 (N_8155,N_3534,N_960);
nand U8156 (N_8156,N_99,N_2884);
nor U8157 (N_8157,N_2189,N_3264);
and U8158 (N_8158,N_3857,N_599);
nand U8159 (N_8159,N_2777,N_3854);
and U8160 (N_8160,N_1227,N_2551);
nor U8161 (N_8161,N_4918,N_3370);
or U8162 (N_8162,N_1778,N_1384);
nor U8163 (N_8163,N_1088,N_2378);
nor U8164 (N_8164,N_75,N_4359);
nor U8165 (N_8165,N_1031,N_2512);
xor U8166 (N_8166,N_2,N_524);
nand U8167 (N_8167,N_1945,N_1379);
nand U8168 (N_8168,N_4363,N_3556);
xor U8169 (N_8169,N_1315,N_2363);
or U8170 (N_8170,N_2156,N_2928);
or U8171 (N_8171,N_4813,N_3281);
and U8172 (N_8172,N_2917,N_2143);
nand U8173 (N_8173,N_538,N_1620);
nor U8174 (N_8174,N_621,N_2880);
nor U8175 (N_8175,N_684,N_3886);
nor U8176 (N_8176,N_2989,N_3363);
nand U8177 (N_8177,N_4288,N_656);
nor U8178 (N_8178,N_3159,N_4941);
nand U8179 (N_8179,N_933,N_3672);
xor U8180 (N_8180,N_523,N_1777);
nand U8181 (N_8181,N_3248,N_1991);
or U8182 (N_8182,N_3261,N_1476);
or U8183 (N_8183,N_768,N_988);
nand U8184 (N_8184,N_3567,N_3147);
nor U8185 (N_8185,N_2305,N_894);
nor U8186 (N_8186,N_4332,N_2273);
and U8187 (N_8187,N_431,N_4181);
or U8188 (N_8188,N_2079,N_2537);
nand U8189 (N_8189,N_2183,N_1078);
and U8190 (N_8190,N_3780,N_2607);
nand U8191 (N_8191,N_4878,N_1918);
or U8192 (N_8192,N_3991,N_1319);
nand U8193 (N_8193,N_3688,N_1562);
nand U8194 (N_8194,N_1506,N_190);
and U8195 (N_8195,N_3249,N_4459);
xnor U8196 (N_8196,N_1459,N_1889);
nor U8197 (N_8197,N_1579,N_3551);
nand U8198 (N_8198,N_4799,N_1324);
nand U8199 (N_8199,N_3923,N_2781);
nor U8200 (N_8200,N_1378,N_3165);
or U8201 (N_8201,N_2374,N_713);
nor U8202 (N_8202,N_3667,N_4714);
nor U8203 (N_8203,N_2716,N_3857);
or U8204 (N_8204,N_1625,N_1005);
and U8205 (N_8205,N_653,N_4936);
nand U8206 (N_8206,N_3990,N_4136);
nor U8207 (N_8207,N_3668,N_2213);
xor U8208 (N_8208,N_2118,N_3762);
or U8209 (N_8209,N_1107,N_1362);
nor U8210 (N_8210,N_1369,N_1663);
nand U8211 (N_8211,N_1922,N_2272);
and U8212 (N_8212,N_1447,N_196);
xnor U8213 (N_8213,N_2301,N_4595);
nor U8214 (N_8214,N_2781,N_1488);
nand U8215 (N_8215,N_2359,N_4753);
and U8216 (N_8216,N_1019,N_214);
xor U8217 (N_8217,N_2950,N_1459);
or U8218 (N_8218,N_2665,N_2499);
or U8219 (N_8219,N_3709,N_3318);
nand U8220 (N_8220,N_3195,N_2487);
nand U8221 (N_8221,N_3630,N_4776);
and U8222 (N_8222,N_1307,N_559);
nor U8223 (N_8223,N_152,N_2467);
nand U8224 (N_8224,N_1830,N_4242);
and U8225 (N_8225,N_4090,N_3680);
and U8226 (N_8226,N_4274,N_1565);
and U8227 (N_8227,N_3623,N_4529);
nand U8228 (N_8228,N_4259,N_2557);
nand U8229 (N_8229,N_3808,N_795);
and U8230 (N_8230,N_442,N_4826);
nand U8231 (N_8231,N_252,N_3276);
nand U8232 (N_8232,N_1264,N_4602);
or U8233 (N_8233,N_2579,N_1978);
xor U8234 (N_8234,N_2495,N_2233);
or U8235 (N_8235,N_1409,N_498);
and U8236 (N_8236,N_3431,N_414);
nand U8237 (N_8237,N_3366,N_3508);
and U8238 (N_8238,N_4874,N_4626);
nand U8239 (N_8239,N_3258,N_3685);
nor U8240 (N_8240,N_3110,N_2718);
or U8241 (N_8241,N_3078,N_3688);
or U8242 (N_8242,N_4942,N_1114);
nand U8243 (N_8243,N_756,N_3327);
and U8244 (N_8244,N_2441,N_1394);
and U8245 (N_8245,N_4803,N_552);
nand U8246 (N_8246,N_3231,N_2328);
xor U8247 (N_8247,N_4688,N_2420);
and U8248 (N_8248,N_1085,N_1699);
nor U8249 (N_8249,N_94,N_677);
xnor U8250 (N_8250,N_4660,N_1964);
xnor U8251 (N_8251,N_4527,N_323);
nand U8252 (N_8252,N_1067,N_4264);
and U8253 (N_8253,N_1165,N_2935);
or U8254 (N_8254,N_3212,N_3842);
or U8255 (N_8255,N_669,N_736);
or U8256 (N_8256,N_3912,N_4721);
nor U8257 (N_8257,N_3365,N_3311);
nand U8258 (N_8258,N_484,N_4277);
and U8259 (N_8259,N_1496,N_2191);
and U8260 (N_8260,N_2862,N_253);
and U8261 (N_8261,N_3271,N_32);
and U8262 (N_8262,N_2763,N_1419);
and U8263 (N_8263,N_1592,N_4706);
xnor U8264 (N_8264,N_3886,N_4922);
or U8265 (N_8265,N_2870,N_476);
nand U8266 (N_8266,N_4289,N_4434);
or U8267 (N_8267,N_2262,N_4139);
xnor U8268 (N_8268,N_2086,N_1834);
or U8269 (N_8269,N_3785,N_470);
or U8270 (N_8270,N_396,N_3441);
and U8271 (N_8271,N_1359,N_4270);
nand U8272 (N_8272,N_4591,N_1477);
or U8273 (N_8273,N_1903,N_4568);
nand U8274 (N_8274,N_3817,N_3665);
and U8275 (N_8275,N_3159,N_4172);
or U8276 (N_8276,N_2013,N_2348);
nand U8277 (N_8277,N_1533,N_1891);
xor U8278 (N_8278,N_2627,N_1757);
or U8279 (N_8279,N_3648,N_4258);
and U8280 (N_8280,N_285,N_3765);
nand U8281 (N_8281,N_2036,N_1766);
and U8282 (N_8282,N_4150,N_699);
or U8283 (N_8283,N_1603,N_4821);
nand U8284 (N_8284,N_4629,N_4027);
nand U8285 (N_8285,N_3524,N_1839);
or U8286 (N_8286,N_820,N_2846);
nor U8287 (N_8287,N_828,N_2551);
nand U8288 (N_8288,N_3778,N_2129);
nand U8289 (N_8289,N_3198,N_351);
or U8290 (N_8290,N_4855,N_3094);
xnor U8291 (N_8291,N_2329,N_2327);
and U8292 (N_8292,N_1201,N_4270);
and U8293 (N_8293,N_1449,N_4499);
or U8294 (N_8294,N_10,N_4225);
xor U8295 (N_8295,N_788,N_4509);
xnor U8296 (N_8296,N_4502,N_3703);
nor U8297 (N_8297,N_4340,N_4575);
nand U8298 (N_8298,N_3868,N_2974);
and U8299 (N_8299,N_3130,N_2110);
nor U8300 (N_8300,N_1456,N_4222);
and U8301 (N_8301,N_614,N_1088);
xor U8302 (N_8302,N_2804,N_2735);
nand U8303 (N_8303,N_4548,N_4331);
or U8304 (N_8304,N_4165,N_3161);
or U8305 (N_8305,N_1606,N_3993);
and U8306 (N_8306,N_1708,N_1631);
or U8307 (N_8307,N_781,N_2605);
or U8308 (N_8308,N_1383,N_4804);
nor U8309 (N_8309,N_2120,N_4928);
or U8310 (N_8310,N_3065,N_2984);
nor U8311 (N_8311,N_109,N_2277);
nor U8312 (N_8312,N_2956,N_1596);
and U8313 (N_8313,N_1390,N_3035);
or U8314 (N_8314,N_3470,N_1554);
nor U8315 (N_8315,N_1135,N_165);
xnor U8316 (N_8316,N_2901,N_1115);
nor U8317 (N_8317,N_4933,N_2710);
nand U8318 (N_8318,N_1045,N_4223);
nand U8319 (N_8319,N_1996,N_3619);
and U8320 (N_8320,N_3075,N_4627);
or U8321 (N_8321,N_1419,N_1841);
and U8322 (N_8322,N_2426,N_4980);
and U8323 (N_8323,N_4984,N_2280);
nand U8324 (N_8324,N_4160,N_49);
xnor U8325 (N_8325,N_4888,N_2131);
or U8326 (N_8326,N_845,N_3847);
nor U8327 (N_8327,N_1353,N_1661);
nor U8328 (N_8328,N_4934,N_2526);
xnor U8329 (N_8329,N_4301,N_893);
and U8330 (N_8330,N_3969,N_4635);
xor U8331 (N_8331,N_942,N_4858);
nor U8332 (N_8332,N_2773,N_1556);
nand U8333 (N_8333,N_4411,N_504);
nor U8334 (N_8334,N_1134,N_4497);
xnor U8335 (N_8335,N_2192,N_4500);
and U8336 (N_8336,N_2090,N_3547);
nor U8337 (N_8337,N_1474,N_3570);
and U8338 (N_8338,N_3323,N_3964);
or U8339 (N_8339,N_2361,N_2773);
nand U8340 (N_8340,N_1803,N_4983);
or U8341 (N_8341,N_4026,N_4911);
and U8342 (N_8342,N_4213,N_4872);
nand U8343 (N_8343,N_2173,N_1352);
xnor U8344 (N_8344,N_1491,N_658);
xnor U8345 (N_8345,N_511,N_1492);
xor U8346 (N_8346,N_2282,N_4191);
nor U8347 (N_8347,N_3017,N_458);
nand U8348 (N_8348,N_1466,N_4458);
xor U8349 (N_8349,N_1485,N_852);
or U8350 (N_8350,N_1002,N_453);
or U8351 (N_8351,N_1915,N_1357);
and U8352 (N_8352,N_2497,N_2377);
and U8353 (N_8353,N_442,N_4186);
and U8354 (N_8354,N_1171,N_368);
or U8355 (N_8355,N_4749,N_1700);
and U8356 (N_8356,N_4849,N_688);
and U8357 (N_8357,N_392,N_803);
xor U8358 (N_8358,N_4306,N_558);
or U8359 (N_8359,N_4705,N_2525);
nand U8360 (N_8360,N_3246,N_2016);
nor U8361 (N_8361,N_3369,N_368);
nand U8362 (N_8362,N_3127,N_2189);
nand U8363 (N_8363,N_3197,N_2661);
and U8364 (N_8364,N_2307,N_3504);
xnor U8365 (N_8365,N_2672,N_1968);
xnor U8366 (N_8366,N_540,N_365);
xor U8367 (N_8367,N_3796,N_4320);
or U8368 (N_8368,N_2304,N_1484);
nor U8369 (N_8369,N_2335,N_2543);
xnor U8370 (N_8370,N_4479,N_3932);
nor U8371 (N_8371,N_216,N_1312);
xnor U8372 (N_8372,N_1359,N_504);
or U8373 (N_8373,N_3417,N_2729);
or U8374 (N_8374,N_90,N_1573);
nor U8375 (N_8375,N_2795,N_2215);
nand U8376 (N_8376,N_1140,N_16);
xor U8377 (N_8377,N_966,N_2020);
nand U8378 (N_8378,N_1534,N_4484);
nand U8379 (N_8379,N_2011,N_2370);
nand U8380 (N_8380,N_3531,N_2736);
nand U8381 (N_8381,N_4123,N_4925);
and U8382 (N_8382,N_1039,N_1967);
or U8383 (N_8383,N_2517,N_4243);
nand U8384 (N_8384,N_2636,N_4026);
and U8385 (N_8385,N_4001,N_106);
nor U8386 (N_8386,N_1997,N_3968);
or U8387 (N_8387,N_293,N_1924);
or U8388 (N_8388,N_9,N_3502);
or U8389 (N_8389,N_3465,N_1402);
and U8390 (N_8390,N_4395,N_3318);
nand U8391 (N_8391,N_4744,N_4814);
and U8392 (N_8392,N_4023,N_4809);
nor U8393 (N_8393,N_470,N_940);
xnor U8394 (N_8394,N_2110,N_2304);
or U8395 (N_8395,N_57,N_576);
nand U8396 (N_8396,N_3291,N_195);
or U8397 (N_8397,N_4696,N_3243);
or U8398 (N_8398,N_4350,N_369);
or U8399 (N_8399,N_3416,N_1961);
xor U8400 (N_8400,N_3801,N_405);
nor U8401 (N_8401,N_2550,N_3878);
and U8402 (N_8402,N_4271,N_4425);
nand U8403 (N_8403,N_4238,N_2509);
nand U8404 (N_8404,N_4269,N_4190);
nand U8405 (N_8405,N_2688,N_4356);
nand U8406 (N_8406,N_711,N_1396);
nor U8407 (N_8407,N_3487,N_1775);
or U8408 (N_8408,N_10,N_3002);
or U8409 (N_8409,N_2159,N_2121);
or U8410 (N_8410,N_2155,N_2060);
nor U8411 (N_8411,N_3901,N_2633);
and U8412 (N_8412,N_3483,N_4307);
nor U8413 (N_8413,N_2105,N_833);
nand U8414 (N_8414,N_1015,N_3421);
and U8415 (N_8415,N_3319,N_3291);
and U8416 (N_8416,N_3243,N_4141);
nor U8417 (N_8417,N_2998,N_143);
xor U8418 (N_8418,N_4794,N_3558);
nand U8419 (N_8419,N_3528,N_72);
or U8420 (N_8420,N_2877,N_3337);
xnor U8421 (N_8421,N_2926,N_4386);
nor U8422 (N_8422,N_4569,N_4970);
and U8423 (N_8423,N_2204,N_2853);
nand U8424 (N_8424,N_1857,N_4253);
or U8425 (N_8425,N_1062,N_4818);
xnor U8426 (N_8426,N_1512,N_937);
and U8427 (N_8427,N_1938,N_4690);
and U8428 (N_8428,N_4647,N_4498);
xor U8429 (N_8429,N_4302,N_2206);
xor U8430 (N_8430,N_2819,N_1444);
xnor U8431 (N_8431,N_3524,N_2343);
xor U8432 (N_8432,N_3001,N_3314);
or U8433 (N_8433,N_4159,N_395);
nor U8434 (N_8434,N_2694,N_2459);
nand U8435 (N_8435,N_3598,N_4190);
nor U8436 (N_8436,N_3757,N_3248);
and U8437 (N_8437,N_3086,N_1090);
xnor U8438 (N_8438,N_1994,N_1206);
or U8439 (N_8439,N_3411,N_4651);
xor U8440 (N_8440,N_3625,N_1281);
and U8441 (N_8441,N_1084,N_3136);
or U8442 (N_8442,N_860,N_1998);
nor U8443 (N_8443,N_552,N_2113);
or U8444 (N_8444,N_2929,N_1022);
xnor U8445 (N_8445,N_4367,N_2675);
and U8446 (N_8446,N_4245,N_1888);
nor U8447 (N_8447,N_3195,N_3656);
nor U8448 (N_8448,N_4315,N_530);
or U8449 (N_8449,N_4321,N_590);
nor U8450 (N_8450,N_3794,N_759);
nand U8451 (N_8451,N_2008,N_4775);
and U8452 (N_8452,N_4166,N_2746);
nand U8453 (N_8453,N_4601,N_402);
and U8454 (N_8454,N_2741,N_3999);
and U8455 (N_8455,N_4255,N_3095);
or U8456 (N_8456,N_4982,N_4334);
nor U8457 (N_8457,N_3961,N_1383);
nor U8458 (N_8458,N_4935,N_1835);
nand U8459 (N_8459,N_4765,N_571);
nand U8460 (N_8460,N_1835,N_486);
or U8461 (N_8461,N_2153,N_626);
and U8462 (N_8462,N_1972,N_3825);
and U8463 (N_8463,N_601,N_2902);
or U8464 (N_8464,N_330,N_4729);
nor U8465 (N_8465,N_3756,N_2691);
and U8466 (N_8466,N_397,N_3032);
nand U8467 (N_8467,N_3908,N_463);
nor U8468 (N_8468,N_2329,N_42);
xnor U8469 (N_8469,N_2855,N_3974);
xnor U8470 (N_8470,N_4103,N_1308);
or U8471 (N_8471,N_2851,N_2476);
nor U8472 (N_8472,N_4201,N_1167);
nand U8473 (N_8473,N_3813,N_4533);
or U8474 (N_8474,N_4060,N_3711);
nor U8475 (N_8475,N_1739,N_3275);
and U8476 (N_8476,N_3185,N_4277);
nor U8477 (N_8477,N_3435,N_3873);
and U8478 (N_8478,N_873,N_1138);
nand U8479 (N_8479,N_671,N_2097);
nor U8480 (N_8480,N_3262,N_2726);
or U8481 (N_8481,N_3333,N_1319);
or U8482 (N_8482,N_806,N_1933);
and U8483 (N_8483,N_955,N_4324);
nand U8484 (N_8484,N_4279,N_1589);
or U8485 (N_8485,N_995,N_3682);
or U8486 (N_8486,N_1911,N_3071);
nor U8487 (N_8487,N_3468,N_706);
nand U8488 (N_8488,N_2761,N_861);
nor U8489 (N_8489,N_858,N_4946);
nand U8490 (N_8490,N_4506,N_2911);
xnor U8491 (N_8491,N_4322,N_2607);
nand U8492 (N_8492,N_4948,N_1621);
nor U8493 (N_8493,N_1423,N_4719);
nor U8494 (N_8494,N_4859,N_4025);
nand U8495 (N_8495,N_4902,N_1072);
and U8496 (N_8496,N_2258,N_1863);
and U8497 (N_8497,N_1429,N_163);
xnor U8498 (N_8498,N_2634,N_4435);
nand U8499 (N_8499,N_1658,N_613);
or U8500 (N_8500,N_3096,N_797);
xor U8501 (N_8501,N_1203,N_1066);
nand U8502 (N_8502,N_4064,N_3573);
nand U8503 (N_8503,N_4308,N_1589);
nor U8504 (N_8504,N_3551,N_118);
or U8505 (N_8505,N_912,N_3941);
xnor U8506 (N_8506,N_927,N_1996);
xnor U8507 (N_8507,N_4350,N_1009);
nor U8508 (N_8508,N_2015,N_989);
or U8509 (N_8509,N_4221,N_1358);
or U8510 (N_8510,N_1438,N_4427);
nor U8511 (N_8511,N_4817,N_4099);
nand U8512 (N_8512,N_1519,N_1682);
nor U8513 (N_8513,N_3787,N_3125);
xor U8514 (N_8514,N_2100,N_2046);
xor U8515 (N_8515,N_4516,N_4787);
nand U8516 (N_8516,N_516,N_1396);
or U8517 (N_8517,N_1695,N_3211);
and U8518 (N_8518,N_270,N_4393);
nor U8519 (N_8519,N_3536,N_1295);
nand U8520 (N_8520,N_1866,N_1734);
nand U8521 (N_8521,N_2574,N_2796);
or U8522 (N_8522,N_3567,N_1170);
or U8523 (N_8523,N_4708,N_271);
or U8524 (N_8524,N_3917,N_4706);
xor U8525 (N_8525,N_177,N_828);
and U8526 (N_8526,N_4339,N_708);
or U8527 (N_8527,N_4492,N_17);
or U8528 (N_8528,N_130,N_4245);
nand U8529 (N_8529,N_2349,N_2331);
nor U8530 (N_8530,N_2914,N_3874);
nor U8531 (N_8531,N_318,N_2995);
or U8532 (N_8532,N_52,N_4642);
nand U8533 (N_8533,N_3717,N_3032);
or U8534 (N_8534,N_554,N_2387);
or U8535 (N_8535,N_2268,N_2367);
nand U8536 (N_8536,N_1946,N_1923);
and U8537 (N_8537,N_1604,N_1722);
xnor U8538 (N_8538,N_4565,N_4033);
nor U8539 (N_8539,N_3087,N_2765);
nor U8540 (N_8540,N_1471,N_4629);
nand U8541 (N_8541,N_4664,N_3831);
and U8542 (N_8542,N_3478,N_3263);
or U8543 (N_8543,N_1573,N_4898);
nand U8544 (N_8544,N_4641,N_504);
nand U8545 (N_8545,N_1822,N_3656);
nand U8546 (N_8546,N_1406,N_629);
and U8547 (N_8547,N_2234,N_3132);
nand U8548 (N_8548,N_3002,N_1409);
nand U8549 (N_8549,N_1266,N_3977);
nand U8550 (N_8550,N_1053,N_3702);
xnor U8551 (N_8551,N_3143,N_3662);
xor U8552 (N_8552,N_4484,N_3175);
xnor U8553 (N_8553,N_1705,N_305);
and U8554 (N_8554,N_0,N_1519);
or U8555 (N_8555,N_3889,N_4477);
or U8556 (N_8556,N_2388,N_2242);
nand U8557 (N_8557,N_2472,N_4540);
nand U8558 (N_8558,N_1108,N_4466);
xnor U8559 (N_8559,N_4174,N_2512);
and U8560 (N_8560,N_77,N_30);
xor U8561 (N_8561,N_458,N_4387);
nand U8562 (N_8562,N_4156,N_1294);
nor U8563 (N_8563,N_2964,N_4203);
xor U8564 (N_8564,N_260,N_2571);
and U8565 (N_8565,N_4070,N_911);
nand U8566 (N_8566,N_2541,N_4290);
or U8567 (N_8567,N_1737,N_3087);
nor U8568 (N_8568,N_3631,N_4763);
or U8569 (N_8569,N_1295,N_2825);
xor U8570 (N_8570,N_4268,N_3469);
nor U8571 (N_8571,N_1806,N_3753);
or U8572 (N_8572,N_1404,N_3267);
or U8573 (N_8573,N_1734,N_2517);
nand U8574 (N_8574,N_67,N_4612);
nand U8575 (N_8575,N_2932,N_1679);
or U8576 (N_8576,N_1436,N_4371);
and U8577 (N_8577,N_4116,N_2273);
or U8578 (N_8578,N_1620,N_3528);
or U8579 (N_8579,N_105,N_4834);
or U8580 (N_8580,N_3203,N_4554);
and U8581 (N_8581,N_1477,N_3874);
xnor U8582 (N_8582,N_1171,N_3711);
nand U8583 (N_8583,N_1645,N_229);
nor U8584 (N_8584,N_3553,N_4437);
nand U8585 (N_8585,N_1767,N_3842);
nor U8586 (N_8586,N_3274,N_1875);
nor U8587 (N_8587,N_35,N_531);
nor U8588 (N_8588,N_2922,N_1533);
nor U8589 (N_8589,N_1538,N_2683);
or U8590 (N_8590,N_2074,N_3826);
nor U8591 (N_8591,N_4384,N_950);
and U8592 (N_8592,N_1673,N_1534);
or U8593 (N_8593,N_2831,N_2165);
and U8594 (N_8594,N_3416,N_510);
nand U8595 (N_8595,N_3696,N_2643);
nand U8596 (N_8596,N_3378,N_168);
xor U8597 (N_8597,N_1166,N_3009);
or U8598 (N_8598,N_3850,N_1193);
xor U8599 (N_8599,N_2585,N_2092);
or U8600 (N_8600,N_3664,N_442);
nor U8601 (N_8601,N_1308,N_4029);
or U8602 (N_8602,N_1423,N_2883);
or U8603 (N_8603,N_1748,N_3789);
xnor U8604 (N_8604,N_4622,N_3987);
xor U8605 (N_8605,N_2005,N_4657);
xor U8606 (N_8606,N_2911,N_688);
and U8607 (N_8607,N_561,N_3012);
xor U8608 (N_8608,N_1288,N_2051);
nand U8609 (N_8609,N_2153,N_4495);
nand U8610 (N_8610,N_3585,N_4076);
xnor U8611 (N_8611,N_1040,N_4798);
xor U8612 (N_8612,N_3012,N_3819);
nor U8613 (N_8613,N_2363,N_4876);
nor U8614 (N_8614,N_1890,N_3600);
and U8615 (N_8615,N_2343,N_314);
nor U8616 (N_8616,N_3001,N_1696);
xnor U8617 (N_8617,N_645,N_4149);
xnor U8618 (N_8618,N_1576,N_611);
or U8619 (N_8619,N_3934,N_1397);
nor U8620 (N_8620,N_4790,N_1098);
or U8621 (N_8621,N_1388,N_1226);
or U8622 (N_8622,N_3862,N_2659);
nor U8623 (N_8623,N_3360,N_1303);
nor U8624 (N_8624,N_3207,N_930);
nor U8625 (N_8625,N_3684,N_561);
xnor U8626 (N_8626,N_4320,N_41);
or U8627 (N_8627,N_782,N_3938);
nor U8628 (N_8628,N_664,N_3564);
nor U8629 (N_8629,N_163,N_4556);
xor U8630 (N_8630,N_3434,N_3385);
nor U8631 (N_8631,N_545,N_3127);
or U8632 (N_8632,N_4181,N_3845);
and U8633 (N_8633,N_4585,N_3475);
xnor U8634 (N_8634,N_2804,N_2482);
and U8635 (N_8635,N_3654,N_2496);
and U8636 (N_8636,N_1991,N_4625);
and U8637 (N_8637,N_2634,N_2240);
xor U8638 (N_8638,N_4509,N_2115);
or U8639 (N_8639,N_1295,N_1149);
or U8640 (N_8640,N_4170,N_112);
xor U8641 (N_8641,N_857,N_3689);
xnor U8642 (N_8642,N_1115,N_4228);
nor U8643 (N_8643,N_2771,N_1751);
nor U8644 (N_8644,N_4365,N_3957);
nor U8645 (N_8645,N_2500,N_4212);
nand U8646 (N_8646,N_221,N_2453);
xnor U8647 (N_8647,N_2239,N_1958);
xnor U8648 (N_8648,N_2876,N_3078);
xnor U8649 (N_8649,N_4497,N_4648);
nand U8650 (N_8650,N_4079,N_4127);
xor U8651 (N_8651,N_3381,N_123);
nand U8652 (N_8652,N_4713,N_4448);
or U8653 (N_8653,N_1896,N_3287);
and U8654 (N_8654,N_3290,N_69);
and U8655 (N_8655,N_1695,N_3488);
nand U8656 (N_8656,N_4941,N_2861);
and U8657 (N_8657,N_3202,N_4056);
nand U8658 (N_8658,N_815,N_4180);
xnor U8659 (N_8659,N_4359,N_4738);
nor U8660 (N_8660,N_2849,N_3562);
nor U8661 (N_8661,N_524,N_561);
and U8662 (N_8662,N_819,N_3300);
and U8663 (N_8663,N_3414,N_3335);
xnor U8664 (N_8664,N_3268,N_1671);
nand U8665 (N_8665,N_3936,N_4739);
nor U8666 (N_8666,N_676,N_3081);
xnor U8667 (N_8667,N_3072,N_3478);
or U8668 (N_8668,N_3939,N_2813);
and U8669 (N_8669,N_2997,N_1451);
nor U8670 (N_8670,N_2020,N_2821);
nor U8671 (N_8671,N_3400,N_1572);
and U8672 (N_8672,N_4062,N_2146);
nand U8673 (N_8673,N_3538,N_234);
or U8674 (N_8674,N_395,N_3685);
xnor U8675 (N_8675,N_3339,N_3093);
nor U8676 (N_8676,N_3776,N_4921);
xnor U8677 (N_8677,N_3130,N_4465);
nor U8678 (N_8678,N_4133,N_4308);
or U8679 (N_8679,N_161,N_1748);
nand U8680 (N_8680,N_2402,N_4356);
nand U8681 (N_8681,N_2866,N_3948);
nor U8682 (N_8682,N_1595,N_271);
or U8683 (N_8683,N_4357,N_1391);
or U8684 (N_8684,N_2259,N_2732);
or U8685 (N_8685,N_775,N_3393);
xnor U8686 (N_8686,N_1536,N_2452);
or U8687 (N_8687,N_780,N_1744);
nor U8688 (N_8688,N_4909,N_3246);
nand U8689 (N_8689,N_2595,N_2006);
and U8690 (N_8690,N_3875,N_1561);
and U8691 (N_8691,N_3401,N_1215);
or U8692 (N_8692,N_42,N_2160);
and U8693 (N_8693,N_4560,N_3033);
nand U8694 (N_8694,N_268,N_763);
and U8695 (N_8695,N_4450,N_2142);
nor U8696 (N_8696,N_1772,N_1700);
nor U8697 (N_8697,N_460,N_1486);
and U8698 (N_8698,N_4514,N_3499);
xnor U8699 (N_8699,N_4329,N_3496);
and U8700 (N_8700,N_3241,N_1680);
nand U8701 (N_8701,N_4790,N_2855);
xnor U8702 (N_8702,N_2565,N_2302);
and U8703 (N_8703,N_1331,N_3719);
or U8704 (N_8704,N_2148,N_293);
nand U8705 (N_8705,N_1700,N_1055);
or U8706 (N_8706,N_2864,N_4883);
and U8707 (N_8707,N_1611,N_3332);
and U8708 (N_8708,N_494,N_3729);
nand U8709 (N_8709,N_2957,N_1565);
xnor U8710 (N_8710,N_1475,N_1527);
xnor U8711 (N_8711,N_3832,N_4822);
nand U8712 (N_8712,N_3376,N_3507);
nand U8713 (N_8713,N_997,N_847);
nand U8714 (N_8714,N_4410,N_2565);
and U8715 (N_8715,N_2471,N_2623);
xnor U8716 (N_8716,N_384,N_2523);
xor U8717 (N_8717,N_1748,N_484);
or U8718 (N_8718,N_4767,N_3173);
and U8719 (N_8719,N_1466,N_290);
xnor U8720 (N_8720,N_3506,N_4981);
and U8721 (N_8721,N_1355,N_4919);
nor U8722 (N_8722,N_2949,N_1945);
xnor U8723 (N_8723,N_1244,N_1006);
xor U8724 (N_8724,N_1525,N_796);
and U8725 (N_8725,N_4597,N_1773);
nor U8726 (N_8726,N_3103,N_2548);
nand U8727 (N_8727,N_3520,N_3003);
xor U8728 (N_8728,N_1522,N_11);
nor U8729 (N_8729,N_4478,N_923);
xor U8730 (N_8730,N_1123,N_1523);
nand U8731 (N_8731,N_2871,N_1516);
and U8732 (N_8732,N_3237,N_1681);
nor U8733 (N_8733,N_4776,N_4365);
nor U8734 (N_8734,N_3098,N_637);
or U8735 (N_8735,N_2511,N_231);
and U8736 (N_8736,N_4808,N_3535);
nand U8737 (N_8737,N_1252,N_479);
nand U8738 (N_8738,N_434,N_4178);
and U8739 (N_8739,N_1819,N_971);
nand U8740 (N_8740,N_2719,N_3516);
or U8741 (N_8741,N_1634,N_3300);
nand U8742 (N_8742,N_262,N_7);
and U8743 (N_8743,N_1750,N_4520);
and U8744 (N_8744,N_4366,N_901);
and U8745 (N_8745,N_4161,N_3364);
nand U8746 (N_8746,N_4995,N_1786);
or U8747 (N_8747,N_3545,N_2828);
and U8748 (N_8748,N_3817,N_2539);
xor U8749 (N_8749,N_1261,N_3117);
nand U8750 (N_8750,N_4920,N_1499);
nand U8751 (N_8751,N_1239,N_4010);
xnor U8752 (N_8752,N_735,N_3339);
and U8753 (N_8753,N_4823,N_3735);
nand U8754 (N_8754,N_537,N_1993);
and U8755 (N_8755,N_2246,N_4570);
nand U8756 (N_8756,N_3071,N_4785);
or U8757 (N_8757,N_2178,N_3289);
or U8758 (N_8758,N_3962,N_4888);
nor U8759 (N_8759,N_2061,N_1097);
or U8760 (N_8760,N_4986,N_320);
and U8761 (N_8761,N_2072,N_2760);
nor U8762 (N_8762,N_2831,N_4859);
or U8763 (N_8763,N_88,N_2041);
nor U8764 (N_8764,N_1450,N_3049);
nand U8765 (N_8765,N_1414,N_56);
and U8766 (N_8766,N_3290,N_2817);
nand U8767 (N_8767,N_4695,N_2434);
xnor U8768 (N_8768,N_1604,N_888);
or U8769 (N_8769,N_3527,N_1645);
xor U8770 (N_8770,N_4392,N_2804);
and U8771 (N_8771,N_848,N_550);
and U8772 (N_8772,N_3021,N_3869);
or U8773 (N_8773,N_4862,N_3481);
xor U8774 (N_8774,N_2900,N_749);
xor U8775 (N_8775,N_3241,N_3960);
and U8776 (N_8776,N_69,N_3308);
or U8777 (N_8777,N_2055,N_709);
nor U8778 (N_8778,N_1288,N_3667);
nand U8779 (N_8779,N_3179,N_3202);
or U8780 (N_8780,N_576,N_3850);
nor U8781 (N_8781,N_4962,N_2886);
or U8782 (N_8782,N_748,N_177);
xor U8783 (N_8783,N_1883,N_2745);
nand U8784 (N_8784,N_2806,N_3570);
or U8785 (N_8785,N_2525,N_2138);
nand U8786 (N_8786,N_4839,N_4943);
nor U8787 (N_8787,N_2938,N_611);
or U8788 (N_8788,N_3261,N_4028);
nor U8789 (N_8789,N_3005,N_2000);
and U8790 (N_8790,N_2354,N_1578);
xor U8791 (N_8791,N_166,N_1395);
xor U8792 (N_8792,N_4576,N_994);
nand U8793 (N_8793,N_118,N_962);
nand U8794 (N_8794,N_76,N_3131);
xnor U8795 (N_8795,N_2359,N_4363);
xor U8796 (N_8796,N_1015,N_2636);
or U8797 (N_8797,N_846,N_4953);
nor U8798 (N_8798,N_1801,N_2368);
and U8799 (N_8799,N_1785,N_2146);
xnor U8800 (N_8800,N_4271,N_3046);
nor U8801 (N_8801,N_2495,N_1749);
nand U8802 (N_8802,N_3842,N_1410);
nor U8803 (N_8803,N_584,N_347);
or U8804 (N_8804,N_3959,N_1953);
nand U8805 (N_8805,N_3096,N_4090);
xor U8806 (N_8806,N_3002,N_4150);
xor U8807 (N_8807,N_384,N_2595);
nor U8808 (N_8808,N_3647,N_3183);
and U8809 (N_8809,N_647,N_2404);
and U8810 (N_8810,N_456,N_2820);
xnor U8811 (N_8811,N_3753,N_1089);
xor U8812 (N_8812,N_976,N_1478);
nand U8813 (N_8813,N_838,N_539);
nor U8814 (N_8814,N_3345,N_4587);
or U8815 (N_8815,N_3675,N_3159);
nor U8816 (N_8816,N_4202,N_2828);
xnor U8817 (N_8817,N_245,N_2081);
or U8818 (N_8818,N_4775,N_2241);
and U8819 (N_8819,N_3261,N_33);
nor U8820 (N_8820,N_759,N_560);
or U8821 (N_8821,N_4168,N_1974);
or U8822 (N_8822,N_4646,N_4895);
xnor U8823 (N_8823,N_597,N_416);
and U8824 (N_8824,N_3250,N_4021);
nor U8825 (N_8825,N_2110,N_300);
xor U8826 (N_8826,N_2195,N_2027);
and U8827 (N_8827,N_3023,N_1428);
or U8828 (N_8828,N_4586,N_4127);
or U8829 (N_8829,N_3181,N_1422);
nor U8830 (N_8830,N_536,N_3292);
nand U8831 (N_8831,N_1667,N_4501);
and U8832 (N_8832,N_4956,N_4793);
nand U8833 (N_8833,N_4753,N_3704);
nor U8834 (N_8834,N_2675,N_3675);
and U8835 (N_8835,N_2315,N_2903);
and U8836 (N_8836,N_947,N_2510);
or U8837 (N_8837,N_1853,N_2247);
nand U8838 (N_8838,N_3892,N_3841);
or U8839 (N_8839,N_1556,N_992);
nand U8840 (N_8840,N_2909,N_1598);
nand U8841 (N_8841,N_858,N_41);
or U8842 (N_8842,N_2606,N_3054);
nand U8843 (N_8843,N_1893,N_3825);
and U8844 (N_8844,N_2126,N_3872);
nor U8845 (N_8845,N_1766,N_2961);
or U8846 (N_8846,N_810,N_4347);
or U8847 (N_8847,N_1382,N_2477);
nand U8848 (N_8848,N_3871,N_980);
xor U8849 (N_8849,N_640,N_2970);
or U8850 (N_8850,N_3661,N_4025);
and U8851 (N_8851,N_3387,N_4188);
nand U8852 (N_8852,N_4343,N_2825);
nand U8853 (N_8853,N_244,N_4009);
xnor U8854 (N_8854,N_4091,N_361);
and U8855 (N_8855,N_1199,N_731);
xnor U8856 (N_8856,N_3384,N_669);
and U8857 (N_8857,N_4319,N_3488);
or U8858 (N_8858,N_3768,N_1599);
and U8859 (N_8859,N_368,N_2968);
nor U8860 (N_8860,N_3959,N_3385);
xnor U8861 (N_8861,N_4295,N_3269);
and U8862 (N_8862,N_304,N_1621);
and U8863 (N_8863,N_3781,N_1325);
nor U8864 (N_8864,N_2108,N_1998);
nand U8865 (N_8865,N_725,N_1994);
nand U8866 (N_8866,N_2561,N_1495);
nor U8867 (N_8867,N_442,N_1658);
and U8868 (N_8868,N_4946,N_1642);
and U8869 (N_8869,N_2731,N_1363);
xnor U8870 (N_8870,N_3802,N_653);
or U8871 (N_8871,N_485,N_3492);
nand U8872 (N_8872,N_2483,N_1590);
or U8873 (N_8873,N_2427,N_2803);
nand U8874 (N_8874,N_3612,N_3388);
nand U8875 (N_8875,N_900,N_1160);
and U8876 (N_8876,N_3429,N_4672);
nor U8877 (N_8877,N_2822,N_4541);
and U8878 (N_8878,N_4137,N_2900);
nand U8879 (N_8879,N_865,N_155);
and U8880 (N_8880,N_3182,N_4109);
nor U8881 (N_8881,N_1054,N_2106);
and U8882 (N_8882,N_2001,N_921);
or U8883 (N_8883,N_4139,N_1149);
nor U8884 (N_8884,N_4226,N_752);
and U8885 (N_8885,N_4067,N_2624);
nor U8886 (N_8886,N_2076,N_2116);
nand U8887 (N_8887,N_3704,N_3799);
nand U8888 (N_8888,N_4456,N_229);
or U8889 (N_8889,N_154,N_1192);
or U8890 (N_8890,N_3790,N_3916);
or U8891 (N_8891,N_2195,N_715);
xor U8892 (N_8892,N_3029,N_1289);
nand U8893 (N_8893,N_758,N_4621);
and U8894 (N_8894,N_3246,N_4420);
xor U8895 (N_8895,N_2556,N_276);
nor U8896 (N_8896,N_264,N_2324);
or U8897 (N_8897,N_614,N_1114);
nand U8898 (N_8898,N_3433,N_1675);
or U8899 (N_8899,N_1282,N_2667);
and U8900 (N_8900,N_1312,N_1088);
or U8901 (N_8901,N_155,N_4312);
nand U8902 (N_8902,N_344,N_616);
nand U8903 (N_8903,N_3123,N_1416);
nor U8904 (N_8904,N_1818,N_859);
or U8905 (N_8905,N_1871,N_3786);
xnor U8906 (N_8906,N_1018,N_540);
or U8907 (N_8907,N_4276,N_95);
and U8908 (N_8908,N_3726,N_2464);
and U8909 (N_8909,N_4588,N_2046);
nor U8910 (N_8910,N_3786,N_2817);
and U8911 (N_8911,N_1404,N_3540);
and U8912 (N_8912,N_1682,N_4076);
xor U8913 (N_8913,N_3513,N_1737);
nor U8914 (N_8914,N_1653,N_1553);
and U8915 (N_8915,N_1862,N_452);
nand U8916 (N_8916,N_4035,N_521);
or U8917 (N_8917,N_1778,N_2728);
nor U8918 (N_8918,N_3545,N_1455);
and U8919 (N_8919,N_4442,N_4111);
and U8920 (N_8920,N_2603,N_1225);
and U8921 (N_8921,N_1877,N_4859);
and U8922 (N_8922,N_2736,N_3415);
or U8923 (N_8923,N_1496,N_4817);
or U8924 (N_8924,N_4161,N_1490);
or U8925 (N_8925,N_1829,N_3009);
or U8926 (N_8926,N_832,N_3382);
or U8927 (N_8927,N_2734,N_3674);
and U8928 (N_8928,N_701,N_4852);
or U8929 (N_8929,N_3305,N_625);
xnor U8930 (N_8930,N_1073,N_1793);
and U8931 (N_8931,N_4483,N_739);
xnor U8932 (N_8932,N_1705,N_839);
xor U8933 (N_8933,N_4768,N_748);
or U8934 (N_8934,N_4446,N_2513);
or U8935 (N_8935,N_2821,N_1527);
or U8936 (N_8936,N_1241,N_3011);
or U8937 (N_8937,N_1773,N_1408);
nor U8938 (N_8938,N_4774,N_4788);
nand U8939 (N_8939,N_4985,N_3980);
nand U8940 (N_8940,N_4717,N_498);
or U8941 (N_8941,N_1618,N_825);
nand U8942 (N_8942,N_624,N_2922);
or U8943 (N_8943,N_79,N_4296);
xnor U8944 (N_8944,N_3643,N_3723);
xor U8945 (N_8945,N_2222,N_4073);
nor U8946 (N_8946,N_3737,N_4811);
or U8947 (N_8947,N_3688,N_4188);
nor U8948 (N_8948,N_1437,N_179);
or U8949 (N_8949,N_1013,N_1208);
nand U8950 (N_8950,N_1962,N_510);
and U8951 (N_8951,N_2578,N_4727);
or U8952 (N_8952,N_952,N_2952);
xnor U8953 (N_8953,N_1737,N_4695);
nor U8954 (N_8954,N_1761,N_3527);
nor U8955 (N_8955,N_957,N_3010);
and U8956 (N_8956,N_2643,N_4280);
nand U8957 (N_8957,N_1002,N_1021);
nand U8958 (N_8958,N_1618,N_3564);
xnor U8959 (N_8959,N_244,N_1616);
and U8960 (N_8960,N_4705,N_1706);
nand U8961 (N_8961,N_1674,N_2404);
nand U8962 (N_8962,N_2683,N_1717);
xnor U8963 (N_8963,N_4751,N_4425);
and U8964 (N_8964,N_3965,N_3852);
and U8965 (N_8965,N_2627,N_2934);
or U8966 (N_8966,N_3892,N_968);
nor U8967 (N_8967,N_671,N_4372);
xor U8968 (N_8968,N_4182,N_607);
xor U8969 (N_8969,N_3965,N_320);
xnor U8970 (N_8970,N_1493,N_126);
nand U8971 (N_8971,N_1826,N_1275);
or U8972 (N_8972,N_1680,N_624);
nor U8973 (N_8973,N_2426,N_719);
nor U8974 (N_8974,N_1811,N_1143);
xnor U8975 (N_8975,N_3671,N_1398);
nor U8976 (N_8976,N_332,N_2730);
nand U8977 (N_8977,N_1641,N_951);
or U8978 (N_8978,N_3358,N_175);
and U8979 (N_8979,N_1928,N_3857);
nand U8980 (N_8980,N_4528,N_1080);
xnor U8981 (N_8981,N_3690,N_4140);
nor U8982 (N_8982,N_3384,N_11);
or U8983 (N_8983,N_897,N_4495);
nand U8984 (N_8984,N_553,N_2953);
and U8985 (N_8985,N_4313,N_2447);
nor U8986 (N_8986,N_881,N_4087);
nor U8987 (N_8987,N_4898,N_3450);
nor U8988 (N_8988,N_4733,N_1474);
xnor U8989 (N_8989,N_576,N_1794);
nor U8990 (N_8990,N_3409,N_1685);
nand U8991 (N_8991,N_3166,N_2812);
nand U8992 (N_8992,N_2132,N_3737);
or U8993 (N_8993,N_764,N_2940);
or U8994 (N_8994,N_1273,N_1804);
or U8995 (N_8995,N_3264,N_2510);
nand U8996 (N_8996,N_2058,N_4872);
and U8997 (N_8997,N_1401,N_1654);
xor U8998 (N_8998,N_4250,N_1161);
and U8999 (N_8999,N_3904,N_2267);
nor U9000 (N_9000,N_2459,N_1568);
nand U9001 (N_9001,N_3659,N_597);
nand U9002 (N_9002,N_1962,N_4023);
nor U9003 (N_9003,N_189,N_371);
nor U9004 (N_9004,N_4109,N_1171);
xor U9005 (N_9005,N_4279,N_2942);
xor U9006 (N_9006,N_4599,N_2357);
nand U9007 (N_9007,N_1625,N_2724);
and U9008 (N_9008,N_96,N_1670);
or U9009 (N_9009,N_3643,N_2770);
nor U9010 (N_9010,N_3176,N_3119);
nor U9011 (N_9011,N_1515,N_1956);
nor U9012 (N_9012,N_2334,N_2196);
xor U9013 (N_9013,N_1328,N_514);
and U9014 (N_9014,N_4623,N_3803);
and U9015 (N_9015,N_4289,N_2290);
or U9016 (N_9016,N_1109,N_1114);
nand U9017 (N_9017,N_14,N_225);
or U9018 (N_9018,N_1467,N_253);
xnor U9019 (N_9019,N_739,N_4812);
nor U9020 (N_9020,N_2696,N_4131);
or U9021 (N_9021,N_491,N_2159);
nor U9022 (N_9022,N_4316,N_4399);
or U9023 (N_9023,N_1781,N_1002);
xnor U9024 (N_9024,N_898,N_392);
xnor U9025 (N_9025,N_1470,N_1377);
nand U9026 (N_9026,N_2939,N_2155);
or U9027 (N_9027,N_284,N_4153);
nor U9028 (N_9028,N_1204,N_4477);
nor U9029 (N_9029,N_4479,N_1841);
nand U9030 (N_9030,N_486,N_2637);
and U9031 (N_9031,N_1517,N_4762);
nor U9032 (N_9032,N_4362,N_4154);
xor U9033 (N_9033,N_3608,N_897);
xnor U9034 (N_9034,N_956,N_84);
nor U9035 (N_9035,N_4661,N_3412);
or U9036 (N_9036,N_4876,N_2310);
xnor U9037 (N_9037,N_4192,N_2977);
nand U9038 (N_9038,N_4246,N_2423);
nor U9039 (N_9039,N_2525,N_1688);
nand U9040 (N_9040,N_4923,N_1427);
xnor U9041 (N_9041,N_4194,N_4718);
or U9042 (N_9042,N_3115,N_529);
xor U9043 (N_9043,N_3777,N_3140);
nor U9044 (N_9044,N_3821,N_3583);
xnor U9045 (N_9045,N_474,N_4732);
nor U9046 (N_9046,N_186,N_808);
nand U9047 (N_9047,N_204,N_4165);
or U9048 (N_9048,N_3491,N_1361);
nor U9049 (N_9049,N_3122,N_1842);
or U9050 (N_9050,N_4610,N_535);
nand U9051 (N_9051,N_525,N_1569);
and U9052 (N_9052,N_4266,N_1058);
and U9053 (N_9053,N_3305,N_4232);
nand U9054 (N_9054,N_4400,N_2553);
and U9055 (N_9055,N_2697,N_1372);
xnor U9056 (N_9056,N_3965,N_3883);
xnor U9057 (N_9057,N_3969,N_2548);
nor U9058 (N_9058,N_820,N_1763);
xnor U9059 (N_9059,N_3384,N_4506);
nor U9060 (N_9060,N_25,N_2429);
nand U9061 (N_9061,N_4311,N_2756);
nor U9062 (N_9062,N_4141,N_1432);
nand U9063 (N_9063,N_3428,N_3649);
and U9064 (N_9064,N_4979,N_3287);
nor U9065 (N_9065,N_1015,N_395);
nand U9066 (N_9066,N_434,N_1068);
xnor U9067 (N_9067,N_3647,N_3238);
or U9068 (N_9068,N_310,N_4551);
nand U9069 (N_9069,N_4987,N_2661);
and U9070 (N_9070,N_4747,N_3685);
or U9071 (N_9071,N_3086,N_3412);
or U9072 (N_9072,N_4940,N_2994);
and U9073 (N_9073,N_1771,N_1850);
and U9074 (N_9074,N_660,N_1506);
and U9075 (N_9075,N_4819,N_3242);
nor U9076 (N_9076,N_2427,N_1683);
nor U9077 (N_9077,N_971,N_1410);
and U9078 (N_9078,N_4591,N_4538);
nand U9079 (N_9079,N_988,N_1052);
xnor U9080 (N_9080,N_4204,N_2850);
nand U9081 (N_9081,N_2731,N_2066);
nand U9082 (N_9082,N_1842,N_2563);
and U9083 (N_9083,N_255,N_2212);
nand U9084 (N_9084,N_4262,N_3522);
nor U9085 (N_9085,N_2982,N_2818);
or U9086 (N_9086,N_840,N_4160);
or U9087 (N_9087,N_169,N_1608);
nand U9088 (N_9088,N_2522,N_1311);
and U9089 (N_9089,N_3090,N_1001);
and U9090 (N_9090,N_1166,N_1390);
and U9091 (N_9091,N_4035,N_1575);
nor U9092 (N_9092,N_1820,N_364);
and U9093 (N_9093,N_4456,N_4962);
nor U9094 (N_9094,N_112,N_2219);
nand U9095 (N_9095,N_1284,N_3568);
nor U9096 (N_9096,N_2778,N_2477);
nor U9097 (N_9097,N_1196,N_4710);
xor U9098 (N_9098,N_2886,N_551);
or U9099 (N_9099,N_3304,N_4902);
nand U9100 (N_9100,N_1725,N_1056);
nand U9101 (N_9101,N_2338,N_3796);
nand U9102 (N_9102,N_2514,N_3385);
nor U9103 (N_9103,N_1227,N_3583);
nor U9104 (N_9104,N_3613,N_1986);
and U9105 (N_9105,N_2246,N_370);
or U9106 (N_9106,N_1044,N_1394);
or U9107 (N_9107,N_1333,N_374);
and U9108 (N_9108,N_3571,N_2073);
and U9109 (N_9109,N_1027,N_4078);
and U9110 (N_9110,N_4571,N_2228);
or U9111 (N_9111,N_2123,N_2519);
or U9112 (N_9112,N_4824,N_505);
nor U9113 (N_9113,N_1676,N_4462);
nand U9114 (N_9114,N_2538,N_615);
or U9115 (N_9115,N_3467,N_4019);
and U9116 (N_9116,N_1454,N_2591);
or U9117 (N_9117,N_881,N_1021);
nand U9118 (N_9118,N_881,N_3855);
and U9119 (N_9119,N_3297,N_3775);
nor U9120 (N_9120,N_4014,N_4389);
or U9121 (N_9121,N_4111,N_2075);
and U9122 (N_9122,N_2866,N_911);
nor U9123 (N_9123,N_2589,N_4839);
or U9124 (N_9124,N_3680,N_3040);
nor U9125 (N_9125,N_1927,N_3180);
nand U9126 (N_9126,N_4896,N_2082);
nand U9127 (N_9127,N_4137,N_1599);
nor U9128 (N_9128,N_2168,N_1086);
nand U9129 (N_9129,N_976,N_2586);
or U9130 (N_9130,N_764,N_1579);
and U9131 (N_9131,N_670,N_3403);
or U9132 (N_9132,N_1329,N_42);
and U9133 (N_9133,N_4297,N_482);
nand U9134 (N_9134,N_3133,N_1863);
nand U9135 (N_9135,N_1314,N_3724);
nor U9136 (N_9136,N_2789,N_157);
xnor U9137 (N_9137,N_2439,N_2229);
nand U9138 (N_9138,N_3470,N_2248);
nor U9139 (N_9139,N_533,N_1234);
and U9140 (N_9140,N_667,N_307);
nor U9141 (N_9141,N_3292,N_961);
nor U9142 (N_9142,N_1137,N_2663);
nand U9143 (N_9143,N_1420,N_3024);
xnor U9144 (N_9144,N_510,N_2279);
nor U9145 (N_9145,N_2174,N_1968);
or U9146 (N_9146,N_561,N_3600);
nor U9147 (N_9147,N_3305,N_3121);
nand U9148 (N_9148,N_2554,N_707);
nor U9149 (N_9149,N_1849,N_1373);
nor U9150 (N_9150,N_701,N_693);
nor U9151 (N_9151,N_1460,N_1094);
and U9152 (N_9152,N_2888,N_687);
nor U9153 (N_9153,N_783,N_4405);
nor U9154 (N_9154,N_4867,N_3780);
xor U9155 (N_9155,N_3968,N_1873);
or U9156 (N_9156,N_1927,N_3610);
and U9157 (N_9157,N_3729,N_4338);
xor U9158 (N_9158,N_4041,N_4949);
or U9159 (N_9159,N_610,N_4926);
or U9160 (N_9160,N_3502,N_2761);
nand U9161 (N_9161,N_1999,N_431);
and U9162 (N_9162,N_4033,N_2272);
nand U9163 (N_9163,N_2990,N_65);
nor U9164 (N_9164,N_2061,N_147);
xor U9165 (N_9165,N_1685,N_993);
nor U9166 (N_9166,N_409,N_4410);
and U9167 (N_9167,N_678,N_3934);
xnor U9168 (N_9168,N_756,N_3412);
or U9169 (N_9169,N_4788,N_2495);
or U9170 (N_9170,N_516,N_4425);
nor U9171 (N_9171,N_3795,N_3151);
nand U9172 (N_9172,N_816,N_3555);
nor U9173 (N_9173,N_3690,N_4791);
nor U9174 (N_9174,N_1733,N_2374);
nor U9175 (N_9175,N_574,N_2161);
nor U9176 (N_9176,N_1976,N_2365);
xnor U9177 (N_9177,N_1032,N_1847);
nand U9178 (N_9178,N_3003,N_3136);
or U9179 (N_9179,N_1811,N_1310);
xor U9180 (N_9180,N_1073,N_4053);
nand U9181 (N_9181,N_2194,N_146);
nand U9182 (N_9182,N_676,N_4545);
xnor U9183 (N_9183,N_1013,N_3352);
and U9184 (N_9184,N_846,N_841);
and U9185 (N_9185,N_3432,N_3604);
and U9186 (N_9186,N_214,N_1593);
nand U9187 (N_9187,N_3926,N_1446);
and U9188 (N_9188,N_1887,N_3548);
and U9189 (N_9189,N_1488,N_3271);
or U9190 (N_9190,N_425,N_4815);
xnor U9191 (N_9191,N_2912,N_2020);
xor U9192 (N_9192,N_1479,N_2522);
and U9193 (N_9193,N_4277,N_2839);
nor U9194 (N_9194,N_4243,N_292);
or U9195 (N_9195,N_3178,N_3001);
and U9196 (N_9196,N_3900,N_3046);
or U9197 (N_9197,N_3068,N_1904);
or U9198 (N_9198,N_216,N_2017);
and U9199 (N_9199,N_4040,N_4758);
nor U9200 (N_9200,N_3548,N_264);
nor U9201 (N_9201,N_3904,N_3319);
or U9202 (N_9202,N_2636,N_3797);
nor U9203 (N_9203,N_4929,N_4834);
nand U9204 (N_9204,N_3204,N_2368);
nor U9205 (N_9205,N_3409,N_3688);
nor U9206 (N_9206,N_1903,N_2970);
or U9207 (N_9207,N_1575,N_1095);
nand U9208 (N_9208,N_4853,N_3874);
and U9209 (N_9209,N_1592,N_3347);
nand U9210 (N_9210,N_797,N_2023);
or U9211 (N_9211,N_2814,N_1575);
nor U9212 (N_9212,N_2306,N_1344);
and U9213 (N_9213,N_1816,N_982);
and U9214 (N_9214,N_2681,N_4292);
or U9215 (N_9215,N_4614,N_3747);
and U9216 (N_9216,N_400,N_396);
and U9217 (N_9217,N_646,N_514);
or U9218 (N_9218,N_2085,N_1317);
xor U9219 (N_9219,N_4832,N_4935);
or U9220 (N_9220,N_3289,N_3001);
nand U9221 (N_9221,N_3142,N_1519);
nand U9222 (N_9222,N_375,N_2690);
nor U9223 (N_9223,N_1473,N_2865);
or U9224 (N_9224,N_4711,N_668);
or U9225 (N_9225,N_2378,N_3736);
xnor U9226 (N_9226,N_2693,N_1940);
or U9227 (N_9227,N_1024,N_3835);
nor U9228 (N_9228,N_3613,N_1164);
nand U9229 (N_9229,N_3829,N_4846);
or U9230 (N_9230,N_1733,N_3331);
nand U9231 (N_9231,N_163,N_3776);
and U9232 (N_9232,N_3076,N_2882);
and U9233 (N_9233,N_1164,N_3458);
nor U9234 (N_9234,N_2211,N_4509);
xnor U9235 (N_9235,N_4923,N_3307);
or U9236 (N_9236,N_4341,N_1853);
nand U9237 (N_9237,N_2704,N_1220);
nor U9238 (N_9238,N_96,N_2763);
or U9239 (N_9239,N_56,N_4068);
or U9240 (N_9240,N_1230,N_3630);
and U9241 (N_9241,N_3482,N_292);
nand U9242 (N_9242,N_2320,N_3172);
nor U9243 (N_9243,N_2706,N_3908);
and U9244 (N_9244,N_250,N_4704);
nor U9245 (N_9245,N_858,N_4218);
xnor U9246 (N_9246,N_1776,N_4549);
and U9247 (N_9247,N_42,N_650);
nand U9248 (N_9248,N_3635,N_2823);
and U9249 (N_9249,N_3842,N_982);
nand U9250 (N_9250,N_68,N_4291);
xnor U9251 (N_9251,N_984,N_2139);
xor U9252 (N_9252,N_997,N_3380);
xnor U9253 (N_9253,N_4389,N_2396);
xor U9254 (N_9254,N_3047,N_2917);
nand U9255 (N_9255,N_4135,N_895);
or U9256 (N_9256,N_2206,N_4324);
nand U9257 (N_9257,N_984,N_4313);
nand U9258 (N_9258,N_1222,N_2905);
nand U9259 (N_9259,N_2704,N_1677);
nor U9260 (N_9260,N_4894,N_1390);
nand U9261 (N_9261,N_2745,N_2142);
or U9262 (N_9262,N_2814,N_1187);
and U9263 (N_9263,N_783,N_2024);
xor U9264 (N_9264,N_2730,N_303);
nand U9265 (N_9265,N_2569,N_1015);
xnor U9266 (N_9266,N_2901,N_1574);
and U9267 (N_9267,N_706,N_2184);
nor U9268 (N_9268,N_4033,N_1311);
or U9269 (N_9269,N_666,N_1173);
xor U9270 (N_9270,N_4371,N_2782);
and U9271 (N_9271,N_1455,N_1417);
or U9272 (N_9272,N_2240,N_1271);
or U9273 (N_9273,N_3173,N_765);
nand U9274 (N_9274,N_3908,N_1154);
and U9275 (N_9275,N_2114,N_4252);
and U9276 (N_9276,N_3007,N_323);
nand U9277 (N_9277,N_1950,N_3507);
or U9278 (N_9278,N_4958,N_959);
xnor U9279 (N_9279,N_4980,N_3020);
and U9280 (N_9280,N_235,N_4880);
nand U9281 (N_9281,N_3605,N_4978);
nor U9282 (N_9282,N_2672,N_1500);
or U9283 (N_9283,N_3638,N_3463);
nor U9284 (N_9284,N_2761,N_297);
or U9285 (N_9285,N_1408,N_4877);
xnor U9286 (N_9286,N_3707,N_2401);
xor U9287 (N_9287,N_4423,N_2345);
or U9288 (N_9288,N_1987,N_1027);
xnor U9289 (N_9289,N_3865,N_967);
nor U9290 (N_9290,N_1507,N_4500);
or U9291 (N_9291,N_4931,N_1782);
xnor U9292 (N_9292,N_2054,N_498);
xor U9293 (N_9293,N_399,N_3896);
xor U9294 (N_9294,N_4934,N_3886);
and U9295 (N_9295,N_2782,N_4342);
and U9296 (N_9296,N_3078,N_922);
or U9297 (N_9297,N_2787,N_36);
nand U9298 (N_9298,N_2167,N_171);
nor U9299 (N_9299,N_1246,N_2997);
or U9300 (N_9300,N_555,N_234);
nand U9301 (N_9301,N_4257,N_4694);
nor U9302 (N_9302,N_329,N_2076);
xor U9303 (N_9303,N_4760,N_3192);
or U9304 (N_9304,N_4351,N_4808);
nand U9305 (N_9305,N_4272,N_1438);
or U9306 (N_9306,N_4394,N_2612);
nor U9307 (N_9307,N_2629,N_4516);
nand U9308 (N_9308,N_3807,N_502);
nor U9309 (N_9309,N_4286,N_2269);
nor U9310 (N_9310,N_3291,N_2743);
nor U9311 (N_9311,N_401,N_3740);
or U9312 (N_9312,N_3945,N_3711);
nor U9313 (N_9313,N_4385,N_2248);
nand U9314 (N_9314,N_4868,N_2280);
nor U9315 (N_9315,N_4527,N_4436);
nor U9316 (N_9316,N_3939,N_631);
or U9317 (N_9317,N_3831,N_1181);
nor U9318 (N_9318,N_4225,N_1973);
xnor U9319 (N_9319,N_4425,N_316);
nand U9320 (N_9320,N_3045,N_2801);
or U9321 (N_9321,N_1700,N_3911);
and U9322 (N_9322,N_296,N_716);
nand U9323 (N_9323,N_970,N_1620);
nor U9324 (N_9324,N_4695,N_548);
or U9325 (N_9325,N_3239,N_3678);
and U9326 (N_9326,N_2803,N_2034);
and U9327 (N_9327,N_722,N_1500);
xnor U9328 (N_9328,N_4240,N_687);
nand U9329 (N_9329,N_162,N_213);
and U9330 (N_9330,N_1447,N_3230);
and U9331 (N_9331,N_1138,N_3081);
nand U9332 (N_9332,N_710,N_559);
or U9333 (N_9333,N_3325,N_2000);
or U9334 (N_9334,N_4417,N_1101);
nor U9335 (N_9335,N_4345,N_2411);
nand U9336 (N_9336,N_1298,N_846);
or U9337 (N_9337,N_853,N_741);
xor U9338 (N_9338,N_364,N_1369);
xor U9339 (N_9339,N_3592,N_117);
nor U9340 (N_9340,N_4426,N_2583);
or U9341 (N_9341,N_463,N_3507);
xnor U9342 (N_9342,N_868,N_1603);
nand U9343 (N_9343,N_3717,N_4682);
nor U9344 (N_9344,N_445,N_4836);
and U9345 (N_9345,N_262,N_3654);
nor U9346 (N_9346,N_3446,N_2309);
and U9347 (N_9347,N_1247,N_3493);
xor U9348 (N_9348,N_4117,N_1561);
xor U9349 (N_9349,N_2229,N_334);
nand U9350 (N_9350,N_3641,N_4480);
nor U9351 (N_9351,N_1378,N_2684);
or U9352 (N_9352,N_4241,N_1052);
nor U9353 (N_9353,N_4717,N_974);
xor U9354 (N_9354,N_2842,N_3911);
nand U9355 (N_9355,N_4971,N_464);
nand U9356 (N_9356,N_3783,N_4734);
and U9357 (N_9357,N_973,N_2);
or U9358 (N_9358,N_3849,N_655);
and U9359 (N_9359,N_2301,N_2631);
xor U9360 (N_9360,N_3495,N_3595);
nor U9361 (N_9361,N_304,N_386);
and U9362 (N_9362,N_3027,N_906);
or U9363 (N_9363,N_3127,N_3474);
nand U9364 (N_9364,N_99,N_4307);
and U9365 (N_9365,N_1484,N_1660);
nor U9366 (N_9366,N_4370,N_3646);
nor U9367 (N_9367,N_3007,N_4501);
and U9368 (N_9368,N_418,N_3423);
xor U9369 (N_9369,N_3627,N_1982);
or U9370 (N_9370,N_3236,N_4992);
and U9371 (N_9371,N_2843,N_3801);
or U9372 (N_9372,N_2823,N_3346);
nor U9373 (N_9373,N_2394,N_3986);
nand U9374 (N_9374,N_2000,N_4979);
nand U9375 (N_9375,N_2283,N_4337);
xnor U9376 (N_9376,N_3869,N_1289);
nand U9377 (N_9377,N_3986,N_1573);
xnor U9378 (N_9378,N_730,N_4125);
nor U9379 (N_9379,N_4680,N_3380);
xnor U9380 (N_9380,N_1744,N_4668);
or U9381 (N_9381,N_1528,N_2420);
nor U9382 (N_9382,N_1961,N_3518);
or U9383 (N_9383,N_3352,N_664);
and U9384 (N_9384,N_4667,N_4853);
nor U9385 (N_9385,N_4355,N_4362);
nand U9386 (N_9386,N_4970,N_1032);
nor U9387 (N_9387,N_2165,N_1179);
nand U9388 (N_9388,N_3875,N_3443);
nor U9389 (N_9389,N_1954,N_2654);
nand U9390 (N_9390,N_1974,N_649);
xor U9391 (N_9391,N_3361,N_895);
nand U9392 (N_9392,N_4162,N_424);
nand U9393 (N_9393,N_2149,N_2429);
xor U9394 (N_9394,N_3645,N_1474);
and U9395 (N_9395,N_1808,N_3533);
xnor U9396 (N_9396,N_4771,N_634);
nand U9397 (N_9397,N_570,N_2726);
and U9398 (N_9398,N_495,N_2598);
or U9399 (N_9399,N_3460,N_3899);
nor U9400 (N_9400,N_4423,N_1839);
nor U9401 (N_9401,N_2368,N_1522);
and U9402 (N_9402,N_848,N_2571);
nand U9403 (N_9403,N_4855,N_3599);
or U9404 (N_9404,N_3070,N_3832);
or U9405 (N_9405,N_4482,N_546);
nand U9406 (N_9406,N_36,N_3631);
or U9407 (N_9407,N_845,N_2333);
or U9408 (N_9408,N_4341,N_3919);
nand U9409 (N_9409,N_3938,N_723);
and U9410 (N_9410,N_3560,N_3581);
and U9411 (N_9411,N_1859,N_4672);
nand U9412 (N_9412,N_1707,N_3763);
and U9413 (N_9413,N_1726,N_648);
xnor U9414 (N_9414,N_599,N_2236);
or U9415 (N_9415,N_2785,N_2791);
and U9416 (N_9416,N_2300,N_1277);
or U9417 (N_9417,N_1541,N_3570);
nand U9418 (N_9418,N_2533,N_4704);
nor U9419 (N_9419,N_3112,N_2112);
xor U9420 (N_9420,N_2523,N_1463);
nand U9421 (N_9421,N_4683,N_2487);
xnor U9422 (N_9422,N_2857,N_264);
nand U9423 (N_9423,N_1761,N_2627);
xnor U9424 (N_9424,N_3557,N_3321);
and U9425 (N_9425,N_3915,N_265);
xor U9426 (N_9426,N_4258,N_3158);
xor U9427 (N_9427,N_4585,N_3594);
or U9428 (N_9428,N_4109,N_2231);
or U9429 (N_9429,N_1978,N_2004);
xnor U9430 (N_9430,N_2776,N_1334);
or U9431 (N_9431,N_3781,N_4148);
xnor U9432 (N_9432,N_1159,N_3025);
and U9433 (N_9433,N_2348,N_2990);
xor U9434 (N_9434,N_4166,N_2878);
or U9435 (N_9435,N_3622,N_4885);
nand U9436 (N_9436,N_3547,N_3940);
nor U9437 (N_9437,N_467,N_4727);
and U9438 (N_9438,N_3617,N_1638);
or U9439 (N_9439,N_500,N_295);
and U9440 (N_9440,N_3494,N_4512);
and U9441 (N_9441,N_3649,N_4718);
nor U9442 (N_9442,N_4594,N_960);
nand U9443 (N_9443,N_4067,N_4084);
or U9444 (N_9444,N_708,N_1468);
nand U9445 (N_9445,N_1160,N_2841);
or U9446 (N_9446,N_4282,N_4946);
or U9447 (N_9447,N_473,N_3506);
and U9448 (N_9448,N_1537,N_3876);
xnor U9449 (N_9449,N_1578,N_9);
nor U9450 (N_9450,N_2464,N_2518);
or U9451 (N_9451,N_3860,N_3706);
nand U9452 (N_9452,N_2628,N_439);
and U9453 (N_9453,N_1398,N_3839);
and U9454 (N_9454,N_70,N_526);
nor U9455 (N_9455,N_2592,N_919);
or U9456 (N_9456,N_4084,N_3770);
and U9457 (N_9457,N_711,N_3620);
nand U9458 (N_9458,N_4057,N_2493);
xor U9459 (N_9459,N_2248,N_3933);
nor U9460 (N_9460,N_333,N_783);
or U9461 (N_9461,N_1704,N_1395);
nor U9462 (N_9462,N_4365,N_624);
and U9463 (N_9463,N_1917,N_4160);
and U9464 (N_9464,N_1698,N_3119);
nand U9465 (N_9465,N_3636,N_2834);
nor U9466 (N_9466,N_2482,N_3853);
nand U9467 (N_9467,N_1631,N_2503);
nand U9468 (N_9468,N_3424,N_3622);
nor U9469 (N_9469,N_1294,N_1140);
or U9470 (N_9470,N_1895,N_3199);
or U9471 (N_9471,N_31,N_2227);
or U9472 (N_9472,N_3715,N_4785);
and U9473 (N_9473,N_983,N_3568);
xnor U9474 (N_9474,N_862,N_2280);
nor U9475 (N_9475,N_2377,N_4214);
nor U9476 (N_9476,N_4925,N_938);
and U9477 (N_9477,N_2526,N_1711);
or U9478 (N_9478,N_715,N_2530);
xor U9479 (N_9479,N_4660,N_1826);
nand U9480 (N_9480,N_4332,N_1734);
nand U9481 (N_9481,N_2713,N_888);
xor U9482 (N_9482,N_2052,N_1259);
xor U9483 (N_9483,N_338,N_2541);
xnor U9484 (N_9484,N_3969,N_861);
nor U9485 (N_9485,N_1025,N_521);
nand U9486 (N_9486,N_2051,N_415);
xor U9487 (N_9487,N_4356,N_4193);
nand U9488 (N_9488,N_3544,N_2552);
or U9489 (N_9489,N_1069,N_1395);
and U9490 (N_9490,N_1010,N_1570);
nor U9491 (N_9491,N_2109,N_188);
xnor U9492 (N_9492,N_103,N_1117);
or U9493 (N_9493,N_3659,N_2433);
nor U9494 (N_9494,N_1065,N_3318);
nor U9495 (N_9495,N_4031,N_1968);
and U9496 (N_9496,N_2538,N_2591);
and U9497 (N_9497,N_1819,N_1260);
nand U9498 (N_9498,N_4231,N_3904);
xnor U9499 (N_9499,N_4005,N_1757);
or U9500 (N_9500,N_3839,N_4410);
or U9501 (N_9501,N_914,N_553);
or U9502 (N_9502,N_3095,N_3326);
nor U9503 (N_9503,N_1182,N_4655);
xnor U9504 (N_9504,N_2290,N_3949);
nor U9505 (N_9505,N_4151,N_3021);
and U9506 (N_9506,N_4745,N_3618);
and U9507 (N_9507,N_1329,N_4762);
nand U9508 (N_9508,N_3772,N_4325);
xor U9509 (N_9509,N_2868,N_504);
nor U9510 (N_9510,N_585,N_2647);
and U9511 (N_9511,N_3327,N_2364);
nand U9512 (N_9512,N_3680,N_2706);
nor U9513 (N_9513,N_673,N_2474);
nor U9514 (N_9514,N_3723,N_2657);
and U9515 (N_9515,N_3568,N_2500);
xnor U9516 (N_9516,N_336,N_1448);
nor U9517 (N_9517,N_3547,N_2448);
and U9518 (N_9518,N_1568,N_4971);
nor U9519 (N_9519,N_4670,N_3928);
nor U9520 (N_9520,N_1484,N_3396);
nand U9521 (N_9521,N_3717,N_4422);
and U9522 (N_9522,N_2864,N_3446);
nand U9523 (N_9523,N_3409,N_958);
nor U9524 (N_9524,N_4803,N_2777);
or U9525 (N_9525,N_4957,N_3094);
xor U9526 (N_9526,N_1891,N_3840);
or U9527 (N_9527,N_4382,N_1152);
and U9528 (N_9528,N_2202,N_3180);
nand U9529 (N_9529,N_2962,N_1019);
xor U9530 (N_9530,N_959,N_3267);
nor U9531 (N_9531,N_722,N_2854);
and U9532 (N_9532,N_4493,N_3065);
nand U9533 (N_9533,N_512,N_1911);
or U9534 (N_9534,N_2423,N_4270);
and U9535 (N_9535,N_4650,N_2854);
xnor U9536 (N_9536,N_4608,N_180);
and U9537 (N_9537,N_1999,N_2869);
or U9538 (N_9538,N_1091,N_1976);
nor U9539 (N_9539,N_2837,N_1666);
xor U9540 (N_9540,N_2553,N_3079);
or U9541 (N_9541,N_4051,N_3440);
and U9542 (N_9542,N_248,N_3694);
nor U9543 (N_9543,N_3442,N_2979);
or U9544 (N_9544,N_2099,N_780);
nor U9545 (N_9545,N_4859,N_1489);
and U9546 (N_9546,N_4739,N_4990);
nor U9547 (N_9547,N_768,N_4937);
nor U9548 (N_9548,N_175,N_2200);
or U9549 (N_9549,N_1096,N_2060);
nand U9550 (N_9550,N_87,N_1830);
nor U9551 (N_9551,N_4408,N_2025);
nand U9552 (N_9552,N_313,N_4041);
nor U9553 (N_9553,N_2423,N_230);
nor U9554 (N_9554,N_1831,N_1828);
xnor U9555 (N_9555,N_3974,N_1902);
or U9556 (N_9556,N_2444,N_1952);
xnor U9557 (N_9557,N_644,N_1515);
or U9558 (N_9558,N_4586,N_4868);
and U9559 (N_9559,N_2697,N_1867);
nor U9560 (N_9560,N_52,N_940);
nand U9561 (N_9561,N_4110,N_1068);
and U9562 (N_9562,N_2323,N_657);
xnor U9563 (N_9563,N_3549,N_2315);
nand U9564 (N_9564,N_4299,N_3514);
nor U9565 (N_9565,N_1325,N_1913);
nand U9566 (N_9566,N_1000,N_3866);
and U9567 (N_9567,N_4889,N_2366);
xnor U9568 (N_9568,N_2553,N_2448);
or U9569 (N_9569,N_761,N_3728);
nand U9570 (N_9570,N_2292,N_4907);
or U9571 (N_9571,N_2033,N_2059);
nand U9572 (N_9572,N_3566,N_4509);
or U9573 (N_9573,N_3329,N_530);
nand U9574 (N_9574,N_4484,N_348);
xnor U9575 (N_9575,N_2243,N_2010);
nor U9576 (N_9576,N_4882,N_1112);
xnor U9577 (N_9577,N_2882,N_3016);
xor U9578 (N_9578,N_2518,N_3836);
xnor U9579 (N_9579,N_1585,N_3137);
nor U9580 (N_9580,N_3486,N_3275);
or U9581 (N_9581,N_4044,N_4073);
and U9582 (N_9582,N_687,N_3424);
nor U9583 (N_9583,N_3633,N_4392);
xnor U9584 (N_9584,N_3507,N_1357);
and U9585 (N_9585,N_994,N_3736);
xnor U9586 (N_9586,N_1502,N_2329);
xor U9587 (N_9587,N_3442,N_4595);
and U9588 (N_9588,N_3148,N_643);
and U9589 (N_9589,N_3726,N_1904);
and U9590 (N_9590,N_3524,N_3817);
nor U9591 (N_9591,N_4732,N_3149);
or U9592 (N_9592,N_3707,N_489);
nand U9593 (N_9593,N_2994,N_3969);
nand U9594 (N_9594,N_3401,N_4091);
or U9595 (N_9595,N_4014,N_3592);
and U9596 (N_9596,N_1626,N_2821);
or U9597 (N_9597,N_3215,N_1109);
xnor U9598 (N_9598,N_573,N_3528);
nor U9599 (N_9599,N_1858,N_4371);
or U9600 (N_9600,N_3943,N_38);
nor U9601 (N_9601,N_1767,N_2810);
xor U9602 (N_9602,N_4848,N_3522);
or U9603 (N_9603,N_981,N_696);
nand U9604 (N_9604,N_302,N_550);
xor U9605 (N_9605,N_2526,N_1551);
nand U9606 (N_9606,N_2896,N_1565);
nor U9607 (N_9607,N_2556,N_2428);
nor U9608 (N_9608,N_2367,N_2710);
or U9609 (N_9609,N_2482,N_3648);
nor U9610 (N_9610,N_2697,N_3991);
and U9611 (N_9611,N_1673,N_2580);
or U9612 (N_9612,N_4378,N_2140);
nor U9613 (N_9613,N_1467,N_1838);
or U9614 (N_9614,N_142,N_2140);
xnor U9615 (N_9615,N_1964,N_3892);
nor U9616 (N_9616,N_325,N_2444);
xor U9617 (N_9617,N_1672,N_3042);
or U9618 (N_9618,N_3240,N_2614);
or U9619 (N_9619,N_1336,N_4970);
nand U9620 (N_9620,N_742,N_3057);
nor U9621 (N_9621,N_3345,N_782);
nor U9622 (N_9622,N_715,N_4650);
or U9623 (N_9623,N_1603,N_3957);
and U9624 (N_9624,N_3705,N_1272);
or U9625 (N_9625,N_4980,N_4476);
nor U9626 (N_9626,N_1998,N_3811);
and U9627 (N_9627,N_934,N_3423);
nor U9628 (N_9628,N_222,N_1581);
or U9629 (N_9629,N_1868,N_3473);
and U9630 (N_9630,N_1287,N_2505);
and U9631 (N_9631,N_426,N_3084);
and U9632 (N_9632,N_933,N_4905);
xnor U9633 (N_9633,N_340,N_70);
or U9634 (N_9634,N_3865,N_828);
or U9635 (N_9635,N_1575,N_1116);
xnor U9636 (N_9636,N_1356,N_3620);
nand U9637 (N_9637,N_107,N_956);
or U9638 (N_9638,N_4745,N_4645);
or U9639 (N_9639,N_1675,N_454);
nand U9640 (N_9640,N_2187,N_3704);
and U9641 (N_9641,N_2442,N_1229);
or U9642 (N_9642,N_4242,N_172);
nor U9643 (N_9643,N_2240,N_3736);
or U9644 (N_9644,N_630,N_1955);
and U9645 (N_9645,N_3047,N_3235);
xor U9646 (N_9646,N_2653,N_3658);
xor U9647 (N_9647,N_3351,N_1678);
xnor U9648 (N_9648,N_3176,N_3551);
nand U9649 (N_9649,N_2139,N_1990);
xor U9650 (N_9650,N_1114,N_4121);
nand U9651 (N_9651,N_2903,N_2739);
or U9652 (N_9652,N_4949,N_4204);
or U9653 (N_9653,N_864,N_862);
nor U9654 (N_9654,N_4804,N_2230);
nor U9655 (N_9655,N_2976,N_4778);
xor U9656 (N_9656,N_2329,N_1073);
or U9657 (N_9657,N_4545,N_1440);
nor U9658 (N_9658,N_3701,N_3521);
nor U9659 (N_9659,N_3460,N_3917);
or U9660 (N_9660,N_4309,N_880);
xor U9661 (N_9661,N_580,N_4637);
nor U9662 (N_9662,N_1758,N_4501);
and U9663 (N_9663,N_2773,N_1034);
and U9664 (N_9664,N_3859,N_4131);
nand U9665 (N_9665,N_2575,N_1792);
nor U9666 (N_9666,N_4881,N_3840);
nor U9667 (N_9667,N_433,N_1759);
or U9668 (N_9668,N_2136,N_4032);
and U9669 (N_9669,N_2413,N_3953);
nor U9670 (N_9670,N_3674,N_2626);
xnor U9671 (N_9671,N_2994,N_588);
and U9672 (N_9672,N_2345,N_1169);
nor U9673 (N_9673,N_1655,N_2063);
xor U9674 (N_9674,N_1248,N_1452);
xnor U9675 (N_9675,N_1325,N_303);
or U9676 (N_9676,N_905,N_2262);
nor U9677 (N_9677,N_800,N_3211);
nor U9678 (N_9678,N_1524,N_1040);
nor U9679 (N_9679,N_624,N_2902);
or U9680 (N_9680,N_2288,N_2165);
or U9681 (N_9681,N_929,N_3226);
nand U9682 (N_9682,N_2142,N_309);
or U9683 (N_9683,N_353,N_1802);
nand U9684 (N_9684,N_4532,N_1401);
or U9685 (N_9685,N_3167,N_647);
xor U9686 (N_9686,N_4023,N_1416);
or U9687 (N_9687,N_3906,N_3453);
or U9688 (N_9688,N_4725,N_3551);
and U9689 (N_9689,N_198,N_930);
or U9690 (N_9690,N_147,N_1187);
and U9691 (N_9691,N_3479,N_4798);
nand U9692 (N_9692,N_755,N_3976);
xor U9693 (N_9693,N_307,N_653);
and U9694 (N_9694,N_4990,N_2393);
and U9695 (N_9695,N_1155,N_4306);
nand U9696 (N_9696,N_3506,N_2794);
nor U9697 (N_9697,N_2265,N_3110);
and U9698 (N_9698,N_4801,N_3500);
and U9699 (N_9699,N_3716,N_4877);
or U9700 (N_9700,N_3596,N_2248);
xor U9701 (N_9701,N_1513,N_4032);
and U9702 (N_9702,N_2380,N_237);
xor U9703 (N_9703,N_4576,N_4202);
xor U9704 (N_9704,N_852,N_1933);
and U9705 (N_9705,N_3268,N_4037);
xor U9706 (N_9706,N_4767,N_4601);
nand U9707 (N_9707,N_2680,N_3660);
nor U9708 (N_9708,N_4155,N_3698);
or U9709 (N_9709,N_2160,N_3137);
nor U9710 (N_9710,N_3076,N_2649);
or U9711 (N_9711,N_4702,N_3443);
nor U9712 (N_9712,N_3865,N_1740);
and U9713 (N_9713,N_1448,N_2028);
nor U9714 (N_9714,N_2641,N_3238);
and U9715 (N_9715,N_1421,N_1486);
xnor U9716 (N_9716,N_1614,N_3061);
xor U9717 (N_9717,N_181,N_2268);
and U9718 (N_9718,N_3888,N_283);
and U9719 (N_9719,N_1970,N_4143);
xor U9720 (N_9720,N_4782,N_2754);
or U9721 (N_9721,N_2268,N_224);
and U9722 (N_9722,N_1608,N_1430);
nor U9723 (N_9723,N_2345,N_723);
or U9724 (N_9724,N_2700,N_1629);
nand U9725 (N_9725,N_2543,N_4743);
nand U9726 (N_9726,N_1855,N_2694);
or U9727 (N_9727,N_3930,N_4678);
and U9728 (N_9728,N_3745,N_585);
xor U9729 (N_9729,N_1551,N_3180);
nand U9730 (N_9730,N_1902,N_1956);
xor U9731 (N_9731,N_2121,N_3651);
or U9732 (N_9732,N_2619,N_804);
or U9733 (N_9733,N_795,N_4382);
xnor U9734 (N_9734,N_671,N_1155);
nor U9735 (N_9735,N_1249,N_1169);
nor U9736 (N_9736,N_4620,N_182);
and U9737 (N_9737,N_2659,N_983);
nand U9738 (N_9738,N_2677,N_1368);
and U9739 (N_9739,N_1528,N_4006);
xnor U9740 (N_9740,N_4433,N_2026);
xnor U9741 (N_9741,N_886,N_1548);
or U9742 (N_9742,N_3916,N_4094);
and U9743 (N_9743,N_3937,N_3315);
nand U9744 (N_9744,N_3453,N_935);
and U9745 (N_9745,N_4903,N_420);
nor U9746 (N_9746,N_368,N_353);
and U9747 (N_9747,N_2402,N_1960);
and U9748 (N_9748,N_3528,N_3276);
nor U9749 (N_9749,N_4985,N_1347);
nor U9750 (N_9750,N_4924,N_1537);
and U9751 (N_9751,N_530,N_3663);
nor U9752 (N_9752,N_3479,N_534);
and U9753 (N_9753,N_4668,N_606);
and U9754 (N_9754,N_1112,N_2753);
nand U9755 (N_9755,N_455,N_624);
nor U9756 (N_9756,N_2178,N_2815);
nand U9757 (N_9757,N_1930,N_3209);
xnor U9758 (N_9758,N_847,N_1268);
xnor U9759 (N_9759,N_1782,N_1469);
nand U9760 (N_9760,N_1869,N_3104);
and U9761 (N_9761,N_633,N_2831);
nand U9762 (N_9762,N_2519,N_1166);
nand U9763 (N_9763,N_3376,N_4431);
xor U9764 (N_9764,N_4495,N_2956);
nor U9765 (N_9765,N_3873,N_2747);
nand U9766 (N_9766,N_1495,N_1905);
xnor U9767 (N_9767,N_1986,N_347);
or U9768 (N_9768,N_2599,N_4069);
nor U9769 (N_9769,N_2055,N_2974);
nor U9770 (N_9770,N_3233,N_1077);
nor U9771 (N_9771,N_1366,N_1282);
and U9772 (N_9772,N_3605,N_2436);
or U9773 (N_9773,N_2927,N_2897);
nor U9774 (N_9774,N_2991,N_707);
and U9775 (N_9775,N_3289,N_2138);
nor U9776 (N_9776,N_4815,N_1212);
and U9777 (N_9777,N_4068,N_4172);
and U9778 (N_9778,N_4585,N_342);
nor U9779 (N_9779,N_2045,N_2671);
and U9780 (N_9780,N_1806,N_4371);
or U9781 (N_9781,N_1703,N_219);
or U9782 (N_9782,N_4704,N_2853);
nor U9783 (N_9783,N_2376,N_1871);
nor U9784 (N_9784,N_3208,N_2114);
or U9785 (N_9785,N_1931,N_4624);
xnor U9786 (N_9786,N_3463,N_4242);
and U9787 (N_9787,N_2579,N_1656);
or U9788 (N_9788,N_2950,N_4211);
nor U9789 (N_9789,N_4620,N_1561);
xor U9790 (N_9790,N_1926,N_4374);
xor U9791 (N_9791,N_2515,N_790);
or U9792 (N_9792,N_1125,N_405);
and U9793 (N_9793,N_2686,N_410);
or U9794 (N_9794,N_3924,N_1541);
nor U9795 (N_9795,N_126,N_1166);
and U9796 (N_9796,N_2609,N_3628);
nor U9797 (N_9797,N_684,N_3763);
or U9798 (N_9798,N_3125,N_3560);
and U9799 (N_9799,N_4670,N_4603);
nor U9800 (N_9800,N_583,N_1554);
and U9801 (N_9801,N_2999,N_3516);
or U9802 (N_9802,N_4314,N_3338);
nor U9803 (N_9803,N_298,N_1320);
nand U9804 (N_9804,N_4781,N_2303);
and U9805 (N_9805,N_484,N_4329);
and U9806 (N_9806,N_4436,N_1267);
and U9807 (N_9807,N_1099,N_4786);
nand U9808 (N_9808,N_2475,N_2255);
xnor U9809 (N_9809,N_3618,N_500);
nor U9810 (N_9810,N_1267,N_939);
and U9811 (N_9811,N_3035,N_2042);
nand U9812 (N_9812,N_4976,N_33);
nor U9813 (N_9813,N_239,N_3334);
xnor U9814 (N_9814,N_1180,N_77);
or U9815 (N_9815,N_130,N_4285);
and U9816 (N_9816,N_4521,N_1894);
and U9817 (N_9817,N_1782,N_4664);
or U9818 (N_9818,N_1642,N_2313);
and U9819 (N_9819,N_2104,N_4248);
xor U9820 (N_9820,N_2762,N_2205);
and U9821 (N_9821,N_2353,N_1509);
nand U9822 (N_9822,N_2046,N_3257);
nand U9823 (N_9823,N_672,N_3543);
xor U9824 (N_9824,N_847,N_3357);
nor U9825 (N_9825,N_4500,N_3062);
nand U9826 (N_9826,N_76,N_3623);
nor U9827 (N_9827,N_480,N_2941);
xnor U9828 (N_9828,N_2742,N_4410);
nand U9829 (N_9829,N_4820,N_4282);
xor U9830 (N_9830,N_3144,N_970);
xnor U9831 (N_9831,N_903,N_3247);
xnor U9832 (N_9832,N_1959,N_3358);
nor U9833 (N_9833,N_1101,N_842);
nand U9834 (N_9834,N_3494,N_3671);
nor U9835 (N_9835,N_4782,N_2271);
and U9836 (N_9836,N_2645,N_4728);
nor U9837 (N_9837,N_3811,N_1138);
xnor U9838 (N_9838,N_2897,N_3375);
nand U9839 (N_9839,N_2603,N_608);
or U9840 (N_9840,N_2000,N_2469);
and U9841 (N_9841,N_2619,N_4163);
nor U9842 (N_9842,N_4330,N_4528);
nand U9843 (N_9843,N_3854,N_290);
nand U9844 (N_9844,N_1962,N_2301);
nand U9845 (N_9845,N_1660,N_418);
nor U9846 (N_9846,N_2645,N_4482);
nand U9847 (N_9847,N_2072,N_2135);
nand U9848 (N_9848,N_3609,N_611);
nor U9849 (N_9849,N_1142,N_4945);
nand U9850 (N_9850,N_3205,N_3268);
or U9851 (N_9851,N_1346,N_3934);
or U9852 (N_9852,N_3496,N_690);
or U9853 (N_9853,N_1001,N_121);
and U9854 (N_9854,N_2803,N_4478);
or U9855 (N_9855,N_2721,N_4605);
or U9856 (N_9856,N_3990,N_4527);
xnor U9857 (N_9857,N_3228,N_989);
xor U9858 (N_9858,N_2954,N_2235);
xor U9859 (N_9859,N_3387,N_1773);
nand U9860 (N_9860,N_4032,N_4823);
or U9861 (N_9861,N_4441,N_4081);
or U9862 (N_9862,N_1383,N_3032);
or U9863 (N_9863,N_1112,N_4421);
and U9864 (N_9864,N_3425,N_4715);
nand U9865 (N_9865,N_3265,N_509);
or U9866 (N_9866,N_2143,N_1578);
nor U9867 (N_9867,N_930,N_3909);
or U9868 (N_9868,N_1251,N_3200);
or U9869 (N_9869,N_92,N_1254);
and U9870 (N_9870,N_1671,N_2114);
nor U9871 (N_9871,N_701,N_4210);
or U9872 (N_9872,N_4642,N_1227);
or U9873 (N_9873,N_4643,N_4443);
xor U9874 (N_9874,N_2817,N_412);
nand U9875 (N_9875,N_648,N_899);
nand U9876 (N_9876,N_2659,N_4549);
or U9877 (N_9877,N_797,N_3395);
nand U9878 (N_9878,N_2324,N_4223);
or U9879 (N_9879,N_18,N_3295);
or U9880 (N_9880,N_3271,N_3659);
nand U9881 (N_9881,N_2914,N_775);
nand U9882 (N_9882,N_1135,N_734);
xnor U9883 (N_9883,N_41,N_1538);
nor U9884 (N_9884,N_1816,N_2855);
nand U9885 (N_9885,N_642,N_4854);
xnor U9886 (N_9886,N_4543,N_3684);
nand U9887 (N_9887,N_3646,N_1368);
or U9888 (N_9888,N_2990,N_3585);
or U9889 (N_9889,N_978,N_3921);
nand U9890 (N_9890,N_3000,N_4448);
or U9891 (N_9891,N_4178,N_3846);
xnor U9892 (N_9892,N_3515,N_397);
xnor U9893 (N_9893,N_852,N_2931);
or U9894 (N_9894,N_2426,N_4786);
nor U9895 (N_9895,N_2523,N_4488);
nor U9896 (N_9896,N_733,N_4810);
nor U9897 (N_9897,N_3730,N_460);
nor U9898 (N_9898,N_230,N_1243);
nand U9899 (N_9899,N_1452,N_258);
xor U9900 (N_9900,N_1123,N_3986);
xor U9901 (N_9901,N_1760,N_4085);
nand U9902 (N_9902,N_553,N_2847);
nor U9903 (N_9903,N_4624,N_4438);
xor U9904 (N_9904,N_3959,N_2154);
or U9905 (N_9905,N_1287,N_2345);
xnor U9906 (N_9906,N_302,N_2429);
and U9907 (N_9907,N_903,N_3249);
xor U9908 (N_9908,N_3608,N_2986);
nand U9909 (N_9909,N_4004,N_743);
nor U9910 (N_9910,N_4061,N_4535);
or U9911 (N_9911,N_4794,N_1234);
and U9912 (N_9912,N_3410,N_1857);
and U9913 (N_9913,N_4995,N_917);
and U9914 (N_9914,N_1778,N_4691);
nor U9915 (N_9915,N_1481,N_1281);
and U9916 (N_9916,N_3708,N_4083);
or U9917 (N_9917,N_3158,N_3515);
or U9918 (N_9918,N_4102,N_4151);
or U9919 (N_9919,N_849,N_114);
or U9920 (N_9920,N_2592,N_1821);
xnor U9921 (N_9921,N_4592,N_4553);
or U9922 (N_9922,N_3101,N_1301);
xor U9923 (N_9923,N_3738,N_3440);
and U9924 (N_9924,N_4398,N_4840);
nor U9925 (N_9925,N_288,N_139);
and U9926 (N_9926,N_1019,N_3578);
and U9927 (N_9927,N_908,N_642);
nand U9928 (N_9928,N_3199,N_1881);
and U9929 (N_9929,N_4905,N_2344);
or U9930 (N_9930,N_3831,N_3833);
nor U9931 (N_9931,N_2301,N_2612);
and U9932 (N_9932,N_1151,N_1981);
xor U9933 (N_9933,N_1237,N_1727);
and U9934 (N_9934,N_897,N_3884);
or U9935 (N_9935,N_692,N_4950);
xnor U9936 (N_9936,N_1576,N_3582);
xnor U9937 (N_9937,N_4962,N_4332);
nor U9938 (N_9938,N_2033,N_4860);
nand U9939 (N_9939,N_3926,N_1728);
and U9940 (N_9940,N_4113,N_30);
xnor U9941 (N_9941,N_4715,N_3265);
xor U9942 (N_9942,N_1271,N_2486);
or U9943 (N_9943,N_2588,N_1946);
nor U9944 (N_9944,N_2439,N_2563);
or U9945 (N_9945,N_4927,N_2373);
xnor U9946 (N_9946,N_300,N_3222);
and U9947 (N_9947,N_2361,N_713);
nor U9948 (N_9948,N_2874,N_3166);
xnor U9949 (N_9949,N_3677,N_4278);
or U9950 (N_9950,N_3837,N_2257);
xor U9951 (N_9951,N_2602,N_1095);
or U9952 (N_9952,N_2909,N_202);
or U9953 (N_9953,N_2156,N_2007);
xor U9954 (N_9954,N_3403,N_3556);
xnor U9955 (N_9955,N_523,N_4407);
xnor U9956 (N_9956,N_1771,N_4401);
and U9957 (N_9957,N_2991,N_3715);
or U9958 (N_9958,N_2293,N_4115);
xor U9959 (N_9959,N_4894,N_2047);
and U9960 (N_9960,N_2613,N_140);
nor U9961 (N_9961,N_4327,N_1266);
or U9962 (N_9962,N_4632,N_2368);
and U9963 (N_9963,N_600,N_1581);
xor U9964 (N_9964,N_3957,N_2859);
nand U9965 (N_9965,N_1123,N_3319);
nor U9966 (N_9966,N_4333,N_1085);
nand U9967 (N_9967,N_1998,N_3700);
nor U9968 (N_9968,N_1052,N_2044);
nor U9969 (N_9969,N_527,N_4323);
nor U9970 (N_9970,N_1613,N_677);
nor U9971 (N_9971,N_4658,N_4692);
xor U9972 (N_9972,N_873,N_879);
nand U9973 (N_9973,N_2164,N_3600);
nor U9974 (N_9974,N_762,N_19);
xnor U9975 (N_9975,N_128,N_3948);
nand U9976 (N_9976,N_171,N_4400);
nand U9977 (N_9977,N_2922,N_1016);
nand U9978 (N_9978,N_3183,N_541);
and U9979 (N_9979,N_2539,N_2805);
and U9980 (N_9980,N_4969,N_1023);
and U9981 (N_9981,N_1502,N_593);
and U9982 (N_9982,N_2745,N_3252);
nor U9983 (N_9983,N_2428,N_374);
nor U9984 (N_9984,N_1781,N_3616);
nand U9985 (N_9985,N_2249,N_3351);
xnor U9986 (N_9986,N_1,N_2086);
nor U9987 (N_9987,N_3358,N_1844);
nand U9988 (N_9988,N_4278,N_1272);
and U9989 (N_9989,N_4841,N_2520);
and U9990 (N_9990,N_2540,N_2335);
xor U9991 (N_9991,N_375,N_2952);
and U9992 (N_9992,N_983,N_3241);
xor U9993 (N_9993,N_2561,N_3167);
and U9994 (N_9994,N_1217,N_3989);
nand U9995 (N_9995,N_184,N_129);
and U9996 (N_9996,N_1045,N_2954);
nor U9997 (N_9997,N_1002,N_4921);
or U9998 (N_9998,N_4627,N_1540);
or U9999 (N_9999,N_4067,N_3932);
nand U10000 (N_10000,N_6128,N_6111);
xnor U10001 (N_10001,N_8378,N_8860);
xor U10002 (N_10002,N_8356,N_8428);
nor U10003 (N_10003,N_5138,N_7520);
and U10004 (N_10004,N_8086,N_6260);
or U10005 (N_10005,N_9140,N_7007);
nand U10006 (N_10006,N_9153,N_7277);
xnor U10007 (N_10007,N_7889,N_8183);
nor U10008 (N_10008,N_6703,N_8655);
nand U10009 (N_10009,N_6993,N_5825);
xor U10010 (N_10010,N_8877,N_8986);
or U10011 (N_10011,N_7340,N_6289);
xor U10012 (N_10012,N_5802,N_6271);
and U10013 (N_10013,N_6667,N_6529);
or U10014 (N_10014,N_8452,N_8400);
nor U10015 (N_10015,N_9579,N_8711);
xor U10016 (N_10016,N_9951,N_6608);
nand U10017 (N_10017,N_7982,N_8505);
nand U10018 (N_10018,N_8257,N_8721);
or U10019 (N_10019,N_7505,N_9356);
xnor U10020 (N_10020,N_5700,N_8719);
nand U10021 (N_10021,N_6774,N_9978);
xnor U10022 (N_10022,N_5252,N_9134);
or U10023 (N_10023,N_9236,N_7790);
nor U10024 (N_10024,N_8493,N_8016);
xnor U10025 (N_10025,N_9173,N_6408);
nand U10026 (N_10026,N_8695,N_9872);
xnor U10027 (N_10027,N_6473,N_5328);
nand U10028 (N_10028,N_8218,N_8867);
xor U10029 (N_10029,N_5632,N_5892);
nor U10030 (N_10030,N_8529,N_8031);
xor U10031 (N_10031,N_7541,N_8756);
xor U10032 (N_10032,N_6579,N_9997);
and U10033 (N_10033,N_6445,N_9314);
xnor U10034 (N_10034,N_6093,N_8783);
nand U10035 (N_10035,N_9865,N_6297);
xor U10036 (N_10036,N_8386,N_5300);
xnor U10037 (N_10037,N_6736,N_8339);
nand U10038 (N_10038,N_7555,N_5239);
and U10039 (N_10039,N_7405,N_5666);
and U10040 (N_10040,N_7574,N_5908);
nand U10041 (N_10041,N_7977,N_6231);
and U10042 (N_10042,N_8114,N_6070);
and U10043 (N_10043,N_6734,N_6560);
nand U10044 (N_10044,N_6116,N_6317);
or U10045 (N_10045,N_5153,N_8311);
or U10046 (N_10046,N_5565,N_7699);
and U10047 (N_10047,N_7586,N_9499);
nand U10048 (N_10048,N_9386,N_8118);
nand U10049 (N_10049,N_5691,N_7479);
and U10050 (N_10050,N_5020,N_5453);
or U10051 (N_10051,N_5334,N_8952);
and U10052 (N_10052,N_9156,N_7421);
xnor U10053 (N_10053,N_6133,N_6810);
and U10054 (N_10054,N_7347,N_5600);
and U10055 (N_10055,N_7459,N_6363);
or U10056 (N_10056,N_8593,N_9383);
nand U10057 (N_10057,N_9910,N_8777);
nand U10058 (N_10058,N_5791,N_7095);
and U10059 (N_10059,N_8241,N_8602);
and U10060 (N_10060,N_8736,N_7538);
nor U10061 (N_10061,N_6991,N_6025);
and U10062 (N_10062,N_7083,N_7192);
or U10063 (N_10063,N_8545,N_9932);
or U10064 (N_10064,N_5952,N_5207);
nor U10065 (N_10065,N_6166,N_7697);
nor U10066 (N_10066,N_7758,N_9805);
nor U10067 (N_10067,N_5939,N_5276);
nand U10068 (N_10068,N_8355,N_9667);
xor U10069 (N_10069,N_8708,N_9034);
or U10070 (N_10070,N_7956,N_5529);
or U10071 (N_10071,N_6427,N_7952);
nor U10072 (N_10072,N_6031,N_9415);
or U10073 (N_10073,N_8781,N_8606);
nand U10074 (N_10074,N_9113,N_6321);
nand U10075 (N_10075,N_6891,N_8390);
nor U10076 (N_10076,N_7589,N_7104);
and U10077 (N_10077,N_9878,N_8525);
xnor U10078 (N_10078,N_9379,N_9715);
and U10079 (N_10079,N_8288,N_9995);
xor U10080 (N_10080,N_7341,N_7934);
nor U10081 (N_10081,N_8383,N_9248);
and U10082 (N_10082,N_5205,N_6165);
xnor U10083 (N_10083,N_9119,N_7848);
nor U10084 (N_10084,N_9183,N_9023);
nor U10085 (N_10085,N_8522,N_6203);
nand U10086 (N_10086,N_6252,N_5278);
nand U10087 (N_10087,N_5193,N_8481);
and U10088 (N_10088,N_7766,N_8673);
nor U10089 (N_10089,N_8296,N_5658);
or U10090 (N_10090,N_7513,N_5848);
and U10091 (N_10091,N_6670,N_5375);
xnor U10092 (N_10092,N_7649,N_8531);
nand U10093 (N_10093,N_7098,N_5832);
xnor U10094 (N_10094,N_5401,N_6362);
nor U10095 (N_10095,N_9365,N_9341);
nand U10096 (N_10096,N_8010,N_7799);
and U10097 (N_10097,N_6618,N_5521);
nand U10098 (N_10098,N_6054,N_8034);
and U10099 (N_10099,N_5436,N_5288);
and U10100 (N_10100,N_9010,N_5373);
nor U10101 (N_10101,N_7121,N_5245);
xor U10102 (N_10102,N_7248,N_9918);
nor U10103 (N_10103,N_6937,N_6151);
xnor U10104 (N_10104,N_6307,N_6443);
nor U10105 (N_10105,N_7967,N_7970);
nand U10106 (N_10106,N_7040,N_6860);
xnor U10107 (N_10107,N_7437,N_6533);
and U10108 (N_10108,N_5818,N_6622);
or U10109 (N_10109,N_7415,N_8855);
or U10110 (N_10110,N_9475,N_5940);
or U10111 (N_10111,N_8475,N_7033);
nor U10112 (N_10112,N_8432,N_6597);
or U10113 (N_10113,N_5315,N_5082);
nand U10114 (N_10114,N_6502,N_9988);
nor U10115 (N_10115,N_6370,N_5972);
nand U10116 (N_10116,N_5195,N_5306);
nand U10117 (N_10117,N_5819,N_9139);
and U10118 (N_10118,N_8157,N_7078);
nor U10119 (N_10119,N_5681,N_5651);
nor U10120 (N_10120,N_7351,N_7549);
xnor U10121 (N_10121,N_9403,N_9271);
nor U10122 (N_10122,N_8170,N_8261);
nand U10123 (N_10123,N_7572,N_6117);
or U10124 (N_10124,N_6309,N_9401);
and U10125 (N_10125,N_8312,N_8396);
or U10126 (N_10126,N_6832,N_9790);
xnor U10127 (N_10127,N_9275,N_7529);
nand U10128 (N_10128,N_7005,N_9874);
and U10129 (N_10129,N_7160,N_8836);
and U10130 (N_10130,N_5302,N_8388);
or U10131 (N_10131,N_6227,N_7317);
or U10132 (N_10132,N_7133,N_9381);
nand U10133 (N_10133,N_6061,N_8385);
nor U10134 (N_10134,N_9111,N_6994);
nand U10135 (N_10135,N_5022,N_8275);
xor U10136 (N_10136,N_9772,N_7516);
nand U10137 (N_10137,N_5606,N_6983);
or U10138 (N_10138,N_5714,N_9882);
xor U10139 (N_10139,N_5670,N_9570);
and U10140 (N_10140,N_6392,N_7680);
and U10141 (N_10141,N_8164,N_5978);
nor U10142 (N_10142,N_9098,N_7526);
nor U10143 (N_10143,N_5754,N_6696);
nor U10144 (N_10144,N_9443,N_5500);
or U10145 (N_10145,N_7226,N_5261);
nor U10146 (N_10146,N_8487,N_6848);
nor U10147 (N_10147,N_8319,N_6655);
and U10148 (N_10148,N_9900,N_8799);
nor U10149 (N_10149,N_9690,N_8773);
nor U10150 (N_10150,N_8917,N_8548);
or U10151 (N_10151,N_9618,N_7820);
and U10152 (N_10152,N_5965,N_8896);
or U10153 (N_10153,N_8080,N_7431);
nand U10154 (N_10154,N_6581,N_8091);
nand U10155 (N_10155,N_8539,N_9881);
nor U10156 (N_10156,N_5394,N_7748);
and U10157 (N_10157,N_6985,N_9843);
and U10158 (N_10158,N_7292,N_7857);
nor U10159 (N_10159,N_9869,N_5219);
nor U10160 (N_10160,N_5314,N_7044);
nor U10161 (N_10161,N_9873,N_8422);
or U10162 (N_10162,N_6114,N_8484);
and U10163 (N_10163,N_8746,N_6178);
xnor U10164 (N_10164,N_5976,N_7662);
and U10165 (N_10165,N_9174,N_5960);
or U10166 (N_10166,N_6112,N_8641);
nand U10167 (N_10167,N_5086,N_6910);
xnor U10168 (N_10168,N_7616,N_7822);
or U10169 (N_10169,N_5184,N_7197);
and U10170 (N_10170,N_9408,N_7238);
and U10171 (N_10171,N_5459,N_5602);
and U10172 (N_10172,N_5228,N_5788);
nand U10173 (N_10173,N_6426,N_9323);
xor U10174 (N_10174,N_9372,N_9244);
xnor U10175 (N_10175,N_5902,N_6024);
nor U10176 (N_10176,N_8216,N_9125);
xor U10177 (N_10177,N_8546,N_8612);
xnor U10178 (N_10178,N_9519,N_7612);
xor U10179 (N_10179,N_9016,N_8850);
xnor U10180 (N_10180,N_7972,N_8532);
xor U10181 (N_10181,N_8090,N_7788);
nor U10182 (N_10182,N_5857,N_6275);
xor U10183 (N_10183,N_9375,N_8151);
xor U10184 (N_10184,N_9544,N_6903);
xor U10185 (N_10185,N_9545,N_7890);
nor U10186 (N_10186,N_7548,N_7331);
or U10187 (N_10187,N_8067,N_5343);
nor U10188 (N_10188,N_5471,N_9378);
nor U10189 (N_10189,N_9482,N_6742);
nor U10190 (N_10190,N_8652,N_6123);
xor U10191 (N_10191,N_7774,N_5116);
nor U10192 (N_10192,N_9114,N_9661);
xor U10193 (N_10193,N_8175,N_7294);
and U10194 (N_10194,N_5094,N_6673);
or U10195 (N_10195,N_7569,N_8600);
and U10196 (N_10196,N_7462,N_8639);
xnor U10197 (N_10197,N_6242,N_9819);
and U10198 (N_10198,N_8139,N_9033);
xnor U10199 (N_10199,N_6998,N_8927);
nand U10200 (N_10200,N_9376,N_7079);
nand U10201 (N_10201,N_9404,N_6568);
and U10202 (N_10202,N_6838,N_7023);
nand U10203 (N_10203,N_9722,N_9250);
nor U10204 (N_10204,N_6907,N_9885);
xnor U10205 (N_10205,N_5784,N_5933);
nand U10206 (N_10206,N_9863,N_6319);
nor U10207 (N_10207,N_6603,N_7099);
or U10208 (N_10208,N_5554,N_5380);
nand U10209 (N_10209,N_6875,N_7198);
nor U10210 (N_10210,N_9556,N_6506);
xnor U10211 (N_10211,N_6060,N_9948);
xor U10212 (N_10212,N_7082,N_5849);
and U10213 (N_10213,N_9505,N_9812);
or U10214 (N_10214,N_7873,N_8054);
or U10215 (N_10215,N_8906,N_8370);
or U10216 (N_10216,N_8550,N_5174);
and U10217 (N_10217,N_8071,N_7831);
nor U10218 (N_10218,N_9669,N_5075);
nor U10219 (N_10219,N_5880,N_8498);
nand U10220 (N_10220,N_5937,N_7624);
or U10221 (N_10221,N_8298,N_6080);
or U10222 (N_10222,N_8039,N_7283);
or U10223 (N_10223,N_9480,N_5172);
or U10224 (N_10224,N_9421,N_5610);
nor U10225 (N_10225,N_5249,N_8795);
nand U10226 (N_10226,N_5585,N_7092);
nor U10227 (N_10227,N_8137,N_7655);
nor U10228 (N_10228,N_7853,N_6758);
or U10229 (N_10229,N_6806,N_8153);
nand U10230 (N_10230,N_8048,N_9827);
and U10231 (N_10231,N_8729,N_9781);
nand U10232 (N_10232,N_5864,N_9684);
and U10233 (N_10233,N_5445,N_7911);
nand U10234 (N_10234,N_5456,N_7753);
and U10235 (N_10235,N_5457,N_6627);
or U10236 (N_10236,N_5284,N_8231);
or U10237 (N_10237,N_8643,N_6600);
nor U10238 (N_10238,N_7707,N_5031);
or U10239 (N_10239,N_8625,N_7406);
xor U10240 (N_10240,N_7834,N_9464);
and U10241 (N_10241,N_6170,N_8975);
nand U10242 (N_10242,N_8154,N_9616);
nand U10243 (N_10243,N_7045,N_8905);
or U10244 (N_10244,N_6801,N_8021);
xnor U10245 (N_10245,N_5498,N_6259);
nand U10246 (N_10246,N_9693,N_6842);
and U10247 (N_10247,N_8540,N_7321);
nand U10248 (N_10248,N_8650,N_5046);
and U10249 (N_10249,N_9525,N_6872);
or U10250 (N_10250,N_7449,N_6167);
nand U10251 (N_10251,N_9506,N_7128);
xor U10252 (N_10252,N_7718,N_6660);
and U10253 (N_10253,N_8519,N_8660);
nor U10254 (N_10254,N_9591,N_8285);
nor U10255 (N_10255,N_6504,N_6045);
xnor U10256 (N_10256,N_9286,N_7690);
xor U10257 (N_10257,N_9603,N_9324);
xor U10258 (N_10258,N_9508,N_8250);
nand U10259 (N_10259,N_5487,N_7508);
xor U10260 (N_10260,N_9729,N_8063);
nor U10261 (N_10261,N_7393,N_8036);
nand U10262 (N_10262,N_8242,N_7071);
nor U10263 (N_10263,N_5566,N_6471);
or U10264 (N_10264,N_9867,N_7592);
nand U10265 (N_10265,N_9583,N_9766);
or U10266 (N_10266,N_5489,N_5021);
or U10267 (N_10267,N_8019,N_6247);
nor U10268 (N_10268,N_9122,N_8597);
nor U10269 (N_10269,N_5110,N_6966);
or U10270 (N_10270,N_6329,N_9943);
xnor U10271 (N_10271,N_5921,N_9337);
and U10272 (N_10272,N_6928,N_6953);
nand U10273 (N_10273,N_6301,N_7367);
or U10274 (N_10274,N_8784,N_9145);
nor U10275 (N_10275,N_8770,N_9413);
or U10276 (N_10276,N_6207,N_9334);
or U10277 (N_10277,N_9658,N_5834);
xor U10278 (N_10278,N_5597,N_7290);
nand U10279 (N_10279,N_9646,N_6556);
xnor U10280 (N_10280,N_7500,N_5291);
or U10281 (N_10281,N_9516,N_9014);
and U10282 (N_10282,N_7016,N_9130);
xor U10283 (N_10283,N_6629,N_7533);
or U10284 (N_10284,N_7635,N_5713);
xnor U10285 (N_10285,N_7135,N_9106);
or U10286 (N_10286,N_9309,N_8694);
or U10287 (N_10287,N_8566,N_8995);
or U10288 (N_10288,N_5214,N_5341);
xnor U10289 (N_10289,N_7936,N_8931);
nor U10290 (N_10290,N_6646,N_6083);
nand U10291 (N_10291,N_8480,N_7583);
nor U10292 (N_10292,N_6645,N_5366);
nor U10293 (N_10293,N_5782,N_7713);
nand U10294 (N_10294,N_9697,N_7828);
xor U10295 (N_10295,N_5707,N_5041);
or U10296 (N_10296,N_5320,N_5593);
xor U10297 (N_10297,N_8782,N_9594);
or U10298 (N_10298,N_7883,N_8789);
and U10299 (N_10299,N_9660,N_5582);
nor U10300 (N_10300,N_8834,N_6285);
nand U10301 (N_10301,N_6492,N_6740);
xor U10302 (N_10302,N_6725,N_6501);
or U10303 (N_10303,N_5798,N_9144);
nor U10304 (N_10304,N_7132,N_6187);
xor U10305 (N_10305,N_7755,N_5226);
nor U10306 (N_10306,N_7236,N_9118);
nand U10307 (N_10307,N_7839,N_6101);
nand U10308 (N_10308,N_6880,N_5614);
and U10309 (N_10309,N_9741,N_9186);
xor U10310 (N_10310,N_8172,N_8558);
nor U10311 (N_10311,N_9941,N_9531);
nor U10312 (N_10312,N_8828,N_8957);
or U10313 (N_10313,N_9619,N_5637);
or U10314 (N_10314,N_9171,N_6404);
or U10315 (N_10315,N_9216,N_6157);
and U10316 (N_10316,N_7084,N_6152);
nor U10317 (N_10317,N_5716,N_6480);
nor U10318 (N_10318,N_5257,N_5641);
or U10319 (N_10319,N_5406,N_8329);
xnor U10320 (N_10320,N_9026,N_7833);
nand U10321 (N_10321,N_5779,N_7225);
nand U10322 (N_10322,N_5999,N_9621);
or U10323 (N_10323,N_7352,N_8797);
xor U10324 (N_10324,N_7062,N_5166);
nor U10325 (N_10325,N_5522,N_6472);
xnor U10326 (N_10326,N_5390,N_7322);
xnor U10327 (N_10327,N_8538,N_8217);
nand U10328 (N_10328,N_9353,N_5561);
and U10329 (N_10329,N_7536,N_5063);
nand U10330 (N_10330,N_6510,N_5592);
nor U10331 (N_10331,N_7603,N_7478);
and U10332 (N_10332,N_7328,N_6639);
or U10333 (N_10333,N_9458,N_5411);
and U10334 (N_10334,N_8680,N_8992);
or U10335 (N_10335,N_8883,N_7058);
nand U10336 (N_10336,N_6677,N_9771);
nor U10337 (N_10337,N_6333,N_5118);
xnor U10338 (N_10338,N_5259,N_9461);
xnor U10339 (N_10339,N_6055,N_5034);
or U10340 (N_10340,N_5435,N_9636);
or U10341 (N_10341,N_9973,N_5845);
and U10342 (N_10342,N_7136,N_5956);
and U10343 (N_10343,N_9093,N_5155);
nor U10344 (N_10344,N_9340,N_5061);
and U10345 (N_10345,N_5254,N_8194);
nand U10346 (N_10346,N_6917,N_9154);
nor U10347 (N_10347,N_9031,N_5891);
nor U10348 (N_10348,N_9871,N_9756);
and U10349 (N_10349,N_6459,N_9041);
xnor U10350 (N_10350,N_7651,N_7167);
nand U10351 (N_10351,N_9860,N_7422);
nand U10352 (N_10352,N_8972,N_9816);
and U10353 (N_10353,N_8894,N_8690);
xor U10354 (N_10354,N_7195,N_8559);
and U10355 (N_10355,N_7960,N_7770);
xor U10356 (N_10356,N_9181,N_8577);
nor U10357 (N_10357,N_9813,N_7102);
xnor U10358 (N_10358,N_7971,N_9839);
nor U10359 (N_10359,N_7885,N_5270);
or U10360 (N_10360,N_6851,N_9203);
nor U10361 (N_10361,N_6914,N_8492);
nor U10362 (N_10362,N_5724,N_7836);
nor U10363 (N_10363,N_6893,N_8024);
or U10364 (N_10364,N_5769,N_9101);
and U10365 (N_10365,N_5431,N_8666);
nand U10366 (N_10366,N_7114,N_7560);
nand U10367 (N_10367,N_7912,N_7900);
nor U10368 (N_10368,N_9892,N_6511);
nor U10369 (N_10369,N_5867,N_8512);
nand U10370 (N_10370,N_5605,N_6044);
xnor U10371 (N_10371,N_9615,N_7204);
nor U10372 (N_10372,N_8045,N_7684);
and U10373 (N_10373,N_9933,N_6730);
nand U10374 (N_10374,N_9189,N_9653);
nand U10375 (N_10375,N_6652,N_7424);
xnor U10376 (N_10376,N_5630,N_7216);
nand U10377 (N_10377,N_9062,N_8207);
xnor U10378 (N_10378,N_6000,N_9185);
nor U10379 (N_10379,N_5621,N_8629);
nand U10380 (N_10380,N_5370,N_6718);
nand U10381 (N_10381,N_5383,N_5115);
or U10382 (N_10382,N_7097,N_5078);
or U10383 (N_10383,N_6246,N_6799);
nand U10384 (N_10384,N_7874,N_6513);
nand U10385 (N_10385,N_7053,N_8087);
and U10386 (N_10386,N_7762,N_9486);
nand U10387 (N_10387,N_9037,N_7069);
and U10388 (N_10388,N_9974,N_9430);
nor U10389 (N_10389,N_8989,N_7776);
nand U10390 (N_10390,N_9142,N_9553);
nor U10391 (N_10391,N_5145,N_7372);
nand U10392 (N_10392,N_6100,N_5823);
and U10393 (N_10393,N_6641,N_7947);
xor U10394 (N_10394,N_9074,N_7807);
or U10395 (N_10395,N_9412,N_8720);
nand U10396 (N_10396,N_8637,N_9162);
or U10397 (N_10397,N_6223,N_6784);
or U10398 (N_10398,N_8093,N_7801);
nand U10399 (N_10399,N_7208,N_5753);
nand U10400 (N_10400,N_8947,N_9352);
or U10401 (N_10401,N_8381,N_5255);
and U10402 (N_10402,N_5290,N_6591);
or U10403 (N_10403,N_5598,N_7050);
nand U10404 (N_10404,N_6381,N_8849);
and U10405 (N_10405,N_5203,N_6216);
nand U10406 (N_10406,N_6613,N_9363);
nor U10407 (N_10407,N_9972,N_6096);
nor U10408 (N_10408,N_5055,N_7810);
or U10409 (N_10409,N_6614,N_7716);
xnor U10410 (N_10410,N_5141,N_7983);
or U10411 (N_10411,N_8585,N_5603);
and U10412 (N_10412,N_7051,N_8671);
or U10413 (N_10413,N_5643,N_6302);
nor U10414 (N_10414,N_7476,N_7173);
nor U10415 (N_10415,N_9633,N_7995);
nand U10416 (N_10416,N_5745,N_7037);
or U10417 (N_10417,N_8700,N_5922);
nand U10418 (N_10418,N_7108,N_8333);
or U10419 (N_10419,N_5631,N_8057);
or U10420 (N_10420,N_7693,N_7920);
or U10421 (N_10421,N_9984,N_7361);
and U10422 (N_10422,N_9308,N_6382);
or U10423 (N_10423,N_9231,N_5690);
nor U10424 (N_10424,N_5757,N_7376);
nor U10425 (N_10425,N_7260,N_6457);
and U10426 (N_10426,N_8376,N_6509);
and U10427 (N_10427,N_7467,N_6724);
or U10428 (N_10428,N_6360,N_8739);
or U10429 (N_10429,N_7838,N_9893);
and U10430 (N_10430,N_6974,N_8027);
nor U10431 (N_10431,N_6159,N_6284);
nand U10432 (N_10432,N_8215,N_8657);
nor U10433 (N_10433,N_8392,N_9747);
and U10434 (N_10434,N_8664,N_7291);
and U10435 (N_10435,N_5865,N_7777);
xnor U10436 (N_10436,N_5579,N_9335);
xnor U10437 (N_10437,N_9573,N_5900);
nand U10438 (N_10438,N_6602,N_9280);
nor U10439 (N_10439,N_7217,N_8767);
xnor U10440 (N_10440,N_9422,N_7757);
xnor U10441 (N_10441,N_8703,N_6535);
nand U10442 (N_10442,N_9282,N_9802);
nand U10443 (N_10443,N_8845,N_9847);
and U10444 (N_10444,N_5243,N_9105);
xor U10445 (N_10445,N_8283,N_9907);
or U10446 (N_10446,N_8199,N_8049);
nand U10447 (N_10447,N_9205,N_7798);
nand U10448 (N_10448,N_8079,N_8617);
xnor U10449 (N_10449,N_8064,N_7360);
and U10450 (N_10450,N_8441,N_6103);
nor U10451 (N_10451,N_7987,N_7953);
nor U10452 (N_10452,N_8224,N_5201);
or U10453 (N_10453,N_5742,N_8421);
nor U10454 (N_10454,N_7120,N_9620);
or U10455 (N_10455,N_7751,N_7390);
xor U10456 (N_10456,N_6057,N_6200);
and U10457 (N_10457,N_6989,N_7116);
or U10458 (N_10458,N_6567,N_5295);
and U10459 (N_10459,N_9195,N_6834);
nand U10460 (N_10460,N_7886,N_9265);
xor U10461 (N_10461,N_9344,N_8884);
nand U10462 (N_10462,N_7392,N_9268);
nand U10463 (N_10463,N_8800,N_5797);
nand U10464 (N_10464,N_8366,N_7100);
xor U10465 (N_10465,N_9494,N_5995);
or U10466 (N_10466,N_9639,N_5869);
nor U10467 (N_10467,N_9698,N_7608);
nand U10468 (N_10468,N_7435,N_8791);
or U10469 (N_10469,N_9507,N_6499);
and U10470 (N_10470,N_6478,N_6446);
and U10471 (N_10471,N_8587,N_5329);
or U10472 (N_10472,N_7740,N_6279);
and U10473 (N_10473,N_7731,N_5191);
xnor U10474 (N_10474,N_5709,N_7319);
and U10475 (N_10475,N_5036,N_6750);
nor U10476 (N_10476,N_5267,N_5842);
xor U10477 (N_10477,N_5628,N_5164);
or U10478 (N_10478,N_9333,N_5948);
xor U10479 (N_10479,N_7324,N_9691);
nor U10480 (N_10480,N_6137,N_5331);
nor U10481 (N_10481,N_8935,N_5230);
nor U10482 (N_10482,N_7414,N_9002);
nor U10483 (N_10483,N_5599,N_9267);
and U10484 (N_10484,N_9318,N_9295);
and U10485 (N_10485,N_5755,N_6726);
and U10486 (N_10486,N_9021,N_9725);
or U10487 (N_10487,N_6265,N_9775);
nand U10488 (N_10488,N_7823,N_7932);
or U10489 (N_10489,N_8478,N_6868);
nand U10490 (N_10490,N_8802,N_7299);
nor U10491 (N_10491,N_9929,N_9252);
or U10492 (N_10492,N_8413,N_7105);
nand U10493 (N_10493,N_8469,N_8909);
nand U10494 (N_10494,N_5005,N_5781);
nor U10495 (N_10495,N_5987,N_7737);
nand U10496 (N_10496,N_6611,N_5231);
and U10497 (N_10497,N_9131,N_7539);
or U10498 (N_10498,N_7253,N_9825);
nor U10499 (N_10499,N_9814,N_5156);
and U10500 (N_10500,N_6245,N_9085);
or U10501 (N_10501,N_9659,N_6977);
xnor U10502 (N_10502,N_9928,N_7381);
xor U10503 (N_10503,N_6763,N_6512);
nand U10504 (N_10504,N_7072,N_8572);
nand U10505 (N_10505,N_8160,N_7382);
and U10506 (N_10506,N_6706,N_7937);
or U10507 (N_10507,N_8996,N_8042);
nand U10508 (N_10508,N_7587,N_5772);
nand U10509 (N_10509,N_9858,N_5543);
nor U10510 (N_10510,N_6470,N_5353);
xor U10511 (N_10511,N_9136,N_7993);
nor U10512 (N_10512,N_8462,N_6691);
or U10513 (N_10513,N_9470,N_6082);
xor U10514 (N_10514,N_9564,N_6104);
xor U10515 (N_10515,N_5897,N_5322);
or U10516 (N_10516,N_6308,N_9688);
and U10517 (N_10517,N_9696,N_6727);
and U10518 (N_10518,N_7418,N_7794);
xnor U10519 (N_10519,N_7343,N_7487);
nor U10520 (N_10520,N_5898,N_9924);
xnor U10521 (N_10521,N_8753,N_7146);
nor U10522 (N_10522,N_8483,N_5007);
nand U10523 (N_10523,N_8128,N_6355);
nand U10524 (N_10524,N_8106,N_7218);
and U10525 (N_10525,N_9079,N_5911);
nor U10526 (N_10526,N_7605,N_8276);
xor U10527 (N_10527,N_9733,N_6476);
nand U10528 (N_10528,N_9438,N_9567);
nor U10529 (N_10529,N_9107,N_7183);
nor U10530 (N_10530,N_9481,N_8638);
nand U10531 (N_10531,N_9483,N_6770);
and U10532 (N_10532,N_5106,N_7280);
or U10533 (N_10533,N_5378,N_6018);
and U10534 (N_10534,N_9009,N_7179);
nand U10535 (N_10535,N_5931,N_8623);
and U10536 (N_10536,N_7096,N_6160);
and U10537 (N_10537,N_6881,N_7949);
nor U10538 (N_10538,N_9479,N_9753);
and U10539 (N_10539,N_5072,N_5563);
or U10540 (N_10540,N_9543,N_6148);
xnor U10541 (N_10541,N_7139,N_5258);
and U10542 (N_10542,N_9495,N_9346);
and U10543 (N_10543,N_6757,N_5917);
nand U10544 (N_10544,N_9606,N_7611);
nor U10545 (N_10545,N_5833,N_7471);
and U10546 (N_10546,N_8969,N_9518);
nor U10547 (N_10547,N_5443,N_7318);
xnor U10548 (N_10548,N_8050,N_6354);
xor U10549 (N_10549,N_5250,N_5699);
xnor U10550 (N_10550,N_6658,N_5830);
nand U10551 (N_10551,N_8354,N_8131);
and U10552 (N_10552,N_8990,N_7270);
and U10553 (N_10553,N_8890,N_6515);
xnor U10554 (N_10554,N_6637,N_7711);
nor U10555 (N_10555,N_9754,N_9586);
and U10556 (N_10556,N_9498,N_5391);
or U10557 (N_10557,N_5475,N_8554);
nor U10558 (N_10558,N_8237,N_7312);
or U10559 (N_10559,N_7524,N_8830);
nand U10560 (N_10560,N_6030,N_6571);
and U10561 (N_10561,N_7369,N_6767);
xor U10562 (N_10562,N_8180,N_6978);
nand U10563 (N_10563,N_6743,N_8179);
and U10564 (N_10564,N_5696,N_5836);
and U10565 (N_10565,N_5402,N_8403);
xnor U10566 (N_10566,N_6379,N_7154);
nor U10567 (N_10567,N_6807,N_8052);
xor U10568 (N_10568,N_5119,N_7247);
nor U10569 (N_10569,N_6339,N_9896);
xnor U10570 (N_10570,N_9992,N_9230);
nor U10571 (N_10571,N_9032,N_7741);
or U10572 (N_10572,N_5015,N_8630);
and U10573 (N_10573,N_7905,N_8166);
nand U10574 (N_10574,N_7942,N_7903);
or U10575 (N_10575,N_9287,N_7618);
and U10576 (N_10576,N_9815,N_5604);
xor U10577 (N_10577,N_6206,N_8264);
xnor U10578 (N_10578,N_5170,N_8727);
and U10579 (N_10579,N_6999,N_5126);
xnor U10580 (N_10580,N_7599,N_8918);
nor U10581 (N_10581,N_9534,N_8107);
xnor U10582 (N_10582,N_8109,N_6884);
nor U10583 (N_10583,N_8099,N_9533);
or U10584 (N_10584,N_8426,N_5444);
and U10585 (N_10585,N_9926,N_9059);
and U10586 (N_10586,N_6984,N_7158);
or U10587 (N_10587,N_7149,N_6531);
nor U10588 (N_10588,N_5095,N_6589);
and U10589 (N_10589,N_9350,N_5074);
or U10590 (N_10590,N_6580,N_9785);
and U10591 (N_10591,N_9366,N_6433);
xor U10592 (N_10592,N_9898,N_5572);
or U10593 (N_10593,N_5958,N_6454);
and U10594 (N_10594,N_6812,N_8651);
and U10595 (N_10595,N_9414,N_6642);
or U10596 (N_10596,N_5874,N_5148);
nand U10597 (N_10597,N_8965,N_7815);
xnor U10598 (N_10598,N_5749,N_7131);
nand U10599 (N_10599,N_5312,N_9194);
xor U10600 (N_10600,N_7940,N_5455);
and U10601 (N_10601,N_8839,N_7320);
xor U10602 (N_10602,N_8959,N_6648);
nor U10603 (N_10603,N_5008,N_9990);
or U10604 (N_10604,N_8331,N_9406);
or U10605 (N_10605,N_9976,N_9739);
nand U10606 (N_10606,N_6697,N_7921);
nor U10607 (N_10607,N_7257,N_8675);
nor U10608 (N_10608,N_8258,N_6771);
nor U10609 (N_10609,N_6253,N_6712);
xnor U10610 (N_10610,N_6234,N_5440);
and U10611 (N_10611,N_6488,N_9612);
nor U10612 (N_10612,N_9610,N_6011);
nand U10613 (N_10613,N_6388,N_6650);
and U10614 (N_10614,N_5669,N_8167);
or U10615 (N_10615,N_5051,N_7152);
nor U10616 (N_10616,N_8389,N_9850);
nor U10617 (N_10617,N_8032,N_9724);
nand U10618 (N_10618,N_6605,N_7330);
nand U10619 (N_10619,N_6190,N_8330);
or U10620 (N_10620,N_8348,N_5645);
nand U10621 (N_10621,N_7075,N_7782);
or U10622 (N_10622,N_6038,N_9317);
nand U10623 (N_10623,N_6890,N_8809);
and U10624 (N_10624,N_6195,N_6986);
nand U10625 (N_10625,N_7189,N_9734);
xor U10626 (N_10626,N_9212,N_8584);
and U10627 (N_10627,N_9143,N_5197);
and U10628 (N_10628,N_5947,N_8780);
nand U10629 (N_10629,N_7284,N_7279);
or U10630 (N_10630,N_8912,N_7775);
and U10631 (N_10631,N_8749,N_8582);
or U10632 (N_10632,N_9744,N_9641);
xor U10633 (N_10633,N_7821,N_6340);
or U10634 (N_10634,N_8244,N_5426);
xor U10635 (N_10635,N_8399,N_9228);
and U10636 (N_10636,N_6258,N_8658);
nor U10637 (N_10637,N_7049,N_9991);
xor U10638 (N_10638,N_6003,N_7623);
or U10639 (N_10639,N_9735,N_7249);
nor U10640 (N_10640,N_5336,N_6437);
and U10641 (N_10641,N_8349,N_8859);
xnor U10642 (N_10642,N_8429,N_7955);
nand U10643 (N_10643,N_8916,N_6349);
xnor U10644 (N_10644,N_5540,N_9135);
nor U10645 (N_10645,N_5124,N_9737);
nor U10646 (N_10646,N_5915,N_6134);
and U10647 (N_10647,N_8615,N_9049);
nor U10648 (N_10648,N_8398,N_5052);
nor U10649 (N_10649,N_6653,N_9115);
nor U10650 (N_10650,N_7047,N_6813);
or U10651 (N_10651,N_9417,N_9213);
nand U10652 (N_10652,N_7577,N_6241);
xor U10653 (N_10653,N_5222,N_8431);
nand U10654 (N_10654,N_9150,N_8728);
or U10655 (N_10655,N_7534,N_9877);
nand U10656 (N_10656,N_9312,N_8454);
nand U10657 (N_10657,N_6251,N_8323);
nor U10658 (N_10658,N_9651,N_7984);
and U10659 (N_10659,N_7501,N_5535);
xor U10660 (N_10660,N_6274,N_7915);
xnor U10661 (N_10661,N_8380,N_6997);
nand U10662 (N_10662,N_7064,N_8000);
xnor U10663 (N_10663,N_5168,N_9076);
and U10664 (N_10664,N_9469,N_9713);
or U10665 (N_10665,N_8635,N_8033);
or U10666 (N_10666,N_5763,N_6145);
or U10667 (N_10667,N_9453,N_8281);
xnor U10668 (N_10668,N_5657,N_9915);
or U10669 (N_10669,N_8304,N_8243);
or U10670 (N_10670,N_8955,N_8162);
or U10671 (N_10671,N_7668,N_7032);
nand U10672 (N_10672,N_7304,N_8161);
xnor U10673 (N_10673,N_6584,N_9884);
nand U10674 (N_10674,N_8136,N_5728);
xor U10675 (N_10675,N_8299,N_8958);
xnor U10676 (N_10676,N_6343,N_8419);
nor U10677 (N_10677,N_5327,N_9081);
and U10678 (N_10678,N_5814,N_8901);
xor U10679 (N_10679,N_6982,N_5695);
or U10680 (N_10680,N_6563,N_6665);
or U10681 (N_10681,N_5629,N_7803);
nor U10682 (N_10682,N_6592,N_7281);
or U10683 (N_10683,N_6168,N_6293);
xnor U10684 (N_10684,N_9398,N_9001);
or U10685 (N_10685,N_6220,N_9833);
nand U10686 (N_10686,N_8534,N_7923);
and U10687 (N_10687,N_5293,N_7695);
nor U10688 (N_10688,N_6829,N_8458);
or U10689 (N_10689,N_8814,N_7460);
xor U10690 (N_10690,N_7151,N_6185);
and U10691 (N_10691,N_8778,N_8563);
xor U10692 (N_10692,N_7841,N_5286);
and U10693 (N_10693,N_8654,N_7582);
and U10694 (N_10694,N_9727,N_6463);
nand U10695 (N_10695,N_6410,N_5866);
nor U10696 (N_10696,N_5639,N_7200);
and U10697 (N_10697,N_9182,N_6164);
and U10698 (N_10698,N_8148,N_7009);
xor U10699 (N_10699,N_5003,N_9095);
xor U10700 (N_10700,N_9072,N_5189);
and U10701 (N_10701,N_5904,N_5640);
nor U10702 (N_10702,N_7250,N_6215);
and U10703 (N_10703,N_7496,N_8801);
nor U10704 (N_10704,N_8200,N_6546);
nand U10705 (N_10705,N_9804,N_8464);
or U10706 (N_10706,N_6788,N_8190);
or U10707 (N_10707,N_6485,N_9227);
nor U10708 (N_10708,N_9638,N_7687);
nor U10709 (N_10709,N_7242,N_6566);
and U10710 (N_10710,N_8122,N_6026);
nand U10711 (N_10711,N_7579,N_7667);
nor U10712 (N_10712,N_5861,N_5142);
nand U10713 (N_10713,N_6261,N_6442);
nor U10714 (N_10714,N_7945,N_7802);
nor U10715 (N_10715,N_9394,N_5547);
and U10716 (N_10716,N_9986,N_6106);
nand U10717 (N_10717,N_7025,N_6617);
and U10718 (N_10718,N_5549,N_9555);
xor U10719 (N_10719,N_7182,N_8440);
xor U10720 (N_10720,N_5750,N_7348);
nor U10721 (N_10721,N_5966,N_6412);
xor U10722 (N_10722,N_9502,N_5526);
nand U10723 (N_10723,N_9908,N_9758);
nand U10724 (N_10724,N_6228,N_7325);
nand U10725 (N_10725,N_8951,N_8196);
or U10726 (N_10726,N_6046,N_7630);
or U10727 (N_10727,N_6610,N_9166);
nor U10728 (N_10728,N_7441,N_9269);
xor U10729 (N_10729,N_6878,N_7337);
nand U10730 (N_10730,N_7617,N_7024);
xnor U10731 (N_10731,N_6599,N_9409);
xor U10732 (N_10732,N_5946,N_6222);
xnor U10733 (N_10733,N_5720,N_6077);
or U10734 (N_10734,N_7297,N_5042);
nand U10735 (N_10735,N_9906,N_8722);
xor U10736 (N_10736,N_9319,N_8324);
or U10737 (N_10737,N_6171,N_5981);
nand U10738 (N_10738,N_6720,N_5458);
or U10739 (N_10739,N_8993,N_6674);
or U10740 (N_10740,N_5425,N_6006);
xor U10741 (N_10741,N_9223,N_6544);
or U10742 (N_10742,N_8555,N_8576);
or U10743 (N_10743,N_7397,N_7004);
nor U10744 (N_10744,N_9266,N_6286);
xor U10745 (N_10745,N_6669,N_7170);
xnor U10746 (N_10746,N_7604,N_5613);
nand U10747 (N_10747,N_9224,N_8537);
nand U10748 (N_10748,N_5274,N_9400);
nor U10749 (N_10749,N_9054,N_5175);
nand U10750 (N_10750,N_9004,N_7504);
and U10751 (N_10751,N_9650,N_6897);
nand U10752 (N_10752,N_9522,N_9528);
and U10753 (N_10753,N_8111,N_6037);
nand U10754 (N_10754,N_6194,N_7580);
nor U10755 (N_10755,N_5377,N_7036);
or U10756 (N_10756,N_6398,N_7591);
xnor U10757 (N_10757,N_6021,N_6738);
nand U10758 (N_10758,N_8823,N_6102);
xor U10759 (N_10759,N_6453,N_8888);
and U10760 (N_10760,N_7825,N_8365);
nand U10761 (N_10761,N_7682,N_5906);
and U10762 (N_10762,N_5418,N_6428);
xnor U10763 (N_10763,N_5183,N_6126);
nand U10764 (N_10764,N_5485,N_7703);
nand U10765 (N_10765,N_5167,N_5423);
and U10766 (N_10766,N_8397,N_9473);
nor U10767 (N_10767,N_6127,N_7888);
nand U10768 (N_10768,N_7654,N_6889);
or U10769 (N_10769,N_8026,N_5693);
xor U10770 (N_10770,N_6539,N_5208);
and U10771 (N_10771,N_8206,N_5012);
nor U10772 (N_10772,N_9354,N_5516);
nor U10773 (N_10773,N_6305,N_9091);
nand U10774 (N_10774,N_8192,N_5744);
nor U10775 (N_10775,N_8163,N_6380);
xor U10776 (N_10776,N_5725,N_9146);
or U10777 (N_10777,N_7455,N_7285);
nand U10778 (N_10778,N_7726,N_6616);
and U10779 (N_10779,N_7796,N_5780);
and U10780 (N_10780,N_7867,N_7963);
or U10781 (N_10781,N_8803,N_8488);
nand U10782 (N_10782,N_6400,N_8640);
and U10783 (N_10783,N_8497,N_9757);
nor U10784 (N_10784,N_6951,N_9169);
and U10785 (N_10785,N_7566,N_5107);
nand U10786 (N_10786,N_6970,N_7458);
nand U10787 (N_10787,N_7689,N_6631);
or U10788 (N_10788,N_5963,N_9259);
xnor U10789 (N_10789,N_6162,N_6542);
nor U10790 (N_10790,N_5766,N_8202);
or U10791 (N_10791,N_8211,N_6013);
or U10792 (N_10792,N_8644,N_5574);
nand U10793 (N_10793,N_7275,N_6040);
nor U10794 (N_10794,N_7792,N_6793);
xor U10795 (N_10795,N_8669,N_5144);
nor U10796 (N_10796,N_6475,N_9315);
or U10797 (N_10797,N_7658,N_5176);
or U10798 (N_10798,N_7676,N_7223);
xor U10799 (N_10799,N_5710,N_9128);
or U10800 (N_10800,N_8309,N_7261);
xnor U10801 (N_10801,N_9431,N_9038);
or U10802 (N_10802,N_9770,N_8345);
nand U10803 (N_10803,N_9238,N_9155);
nor U10804 (N_10804,N_9748,N_9277);
and U10805 (N_10805,N_8415,N_9965);
and U10806 (N_10806,N_6822,N_6318);
and U10807 (N_10807,N_6828,N_7342);
or U10808 (N_10808,N_6198,N_8726);
or U10809 (N_10809,N_9761,N_6022);
nand U10810 (N_10810,N_8934,N_9046);
xor U10811 (N_10811,N_5680,N_5962);
nand U10812 (N_10812,N_9025,N_9336);
nand U10813 (N_10813,N_6762,N_9439);
nor U10814 (N_10814,N_5117,N_5277);
xnor U10815 (N_10815,N_7485,N_9226);
or U10816 (N_10816,N_9446,N_8482);
or U10817 (N_10817,N_8507,N_7003);
nor U10818 (N_10818,N_6933,N_8040);
xor U10819 (N_10819,N_6066,N_8910);
and U10820 (N_10820,N_5247,N_8844);
and U10821 (N_10821,N_9681,N_8515);
nor U10822 (N_10822,N_5178,N_8377);
nor U10823 (N_10823,N_8858,N_5149);
nand U10824 (N_10824,N_5828,N_9369);
nor U10825 (N_10825,N_9796,N_8123);
xnor U10826 (N_10826,N_9117,N_8158);
nand U10827 (N_10827,N_6780,N_8557);
xor U10828 (N_10828,N_6979,N_9755);
and U10829 (N_10829,N_5916,N_5337);
xnor U10830 (N_10830,N_7795,N_7314);
or U10831 (N_10831,N_8315,N_8564);
and U10832 (N_10832,N_5213,N_8065);
nor U10833 (N_10833,N_7329,N_7564);
nand U10834 (N_10834,N_9931,N_7975);
nand U10835 (N_10835,N_7518,N_9345);
or U10836 (N_10836,N_6396,N_7412);
and U10837 (N_10837,N_5491,N_7819);
nor U10838 (N_10838,N_7417,N_6193);
nand U10839 (N_10839,N_8527,N_9560);
nand U10840 (N_10840,N_5612,N_6825);
nor U10841 (N_10841,N_5241,N_6331);
xnor U10842 (N_10842,N_6948,N_8873);
and U10843 (N_10843,N_5979,N_6921);
xnor U10844 (N_10844,N_5556,N_8230);
xor U10845 (N_10845,N_9993,N_7484);
nand U10846 (N_10846,N_7207,N_9512);
and U10847 (N_10847,N_8936,N_5002);
and U10848 (N_10848,N_5820,N_7222);
and U10849 (N_10849,N_8372,N_7364);
xor U10850 (N_10850,N_6281,N_9731);
and U10851 (N_10851,N_5747,N_9665);
and U10852 (N_10852,N_7813,N_9405);
nand U10853 (N_10853,N_9311,N_7897);
nand U10854 (N_10854,N_7744,N_8226);
and U10855 (N_10855,N_5659,N_9500);
or U10856 (N_10856,N_5760,N_7391);
and U10857 (N_10857,N_9167,N_9856);
xnor U10858 (N_10858,N_9679,N_9423);
nand U10859 (N_10859,N_6522,N_8547);
xor U10860 (N_10860,N_7087,N_6047);
nand U10861 (N_10861,N_5502,N_7551);
or U10862 (N_10862,N_8500,N_9300);
xnor U10863 (N_10863,N_5688,N_6590);
nand U10864 (N_10864,N_9673,N_8596);
xor U10865 (N_10865,N_7293,N_7615);
and U10866 (N_10866,N_7276,N_6972);
nor U10867 (N_10867,N_5360,N_8165);
nor U10868 (N_10868,N_8130,N_6945);
or U10869 (N_10869,N_6325,N_6182);
nor U10870 (N_10870,N_7784,N_9395);
xnor U10871 (N_10871,N_5805,N_9656);
nor U10872 (N_10872,N_6892,N_9799);
or U10873 (N_10873,N_8827,N_5347);
nand U10874 (N_10874,N_9706,N_8286);
xnor U10875 (N_10875,N_7313,N_8266);
and U10876 (N_10876,N_8874,N_9728);
nand U10877 (N_10877,N_5729,N_6859);
nor U10878 (N_10878,N_7336,N_5488);
nand U10879 (N_10879,N_9313,N_6422);
nor U10880 (N_10880,N_6681,N_5804);
xor U10881 (N_10881,N_8930,N_7728);
and U10882 (N_10882,N_9187,N_9485);
or U10883 (N_10883,N_8956,N_7073);
xor U10884 (N_10884,N_8279,N_5844);
nor U10885 (N_10885,N_8846,N_7333);
nand U10886 (N_10886,N_6612,N_9511);
nand U10887 (N_10887,N_8028,N_8987);
or U10888 (N_10888,N_8634,N_7408);
xor U10889 (N_10889,N_9530,N_8822);
nand U10890 (N_10890,N_9424,N_8685);
or U10891 (N_10891,N_5244,N_9307);
xnor U10892 (N_10892,N_7598,N_5281);
and U10893 (N_10893,N_9890,N_5575);
nor U10894 (N_10894,N_5080,N_9640);
and U10895 (N_10895,N_9602,N_6448);
or U10896 (N_10896,N_5092,N_6615);
nor U10897 (N_10897,N_9963,N_5530);
xnor U10898 (N_10898,N_6455,N_8046);
nor U10899 (N_10899,N_9838,N_5079);
nor U10900 (N_10900,N_9407,N_8698);
or U10901 (N_10901,N_7315,N_5212);
xnor U10902 (N_10902,N_5664,N_8603);
nand U10903 (N_10903,N_6809,N_7423);
nor U10904 (N_10904,N_5047,N_5679);
or U10905 (N_10905,N_7057,N_6263);
nand U10906 (N_10906,N_9994,N_5321);
nor U10907 (N_10907,N_9912,N_8232);
nor U10908 (N_10908,N_7377,N_7878);
and U10909 (N_10909,N_8280,N_5103);
nand U10910 (N_10910,N_7679,N_9437);
xnor U10911 (N_10911,N_6888,N_9945);
nand U10912 (N_10912,N_5240,N_7155);
nor U10913 (N_10913,N_6395,N_7402);
and U10914 (N_10914,N_7166,N_8999);
and U10915 (N_10915,N_9909,N_8412);
and U10916 (N_10916,N_7661,N_5570);
xnor U10917 (N_10917,N_6585,N_8950);
nor U10918 (N_10918,N_7927,N_5953);
xor U10919 (N_10919,N_6855,N_5428);
nor U10920 (N_10920,N_5465,N_8908);
nor U10921 (N_10921,N_7483,N_6495);
and U10922 (N_10922,N_7127,N_5501);
and U10923 (N_10923,N_9861,N_9547);
or U10924 (N_10924,N_8631,N_8082);
nand U10925 (N_10925,N_7389,N_6419);
or U10926 (N_10926,N_8209,N_9459);
and U10927 (N_10927,N_8661,N_7126);
xnor U10928 (N_10928,N_8774,N_6464);
xnor U10929 (N_10929,N_9589,N_7666);
nand U10930 (N_10930,N_9901,N_9806);
nor U10931 (N_10931,N_7332,N_9961);
and U10932 (N_10932,N_5807,N_9028);
nor U10933 (N_10933,N_8621,N_7973);
nor U10934 (N_10934,N_6371,N_9100);
nand U10935 (N_10935,N_6795,N_7300);
nand U10936 (N_10936,N_6865,N_9410);
nor U10937 (N_10937,N_6779,N_7165);
and U10938 (N_10938,N_5060,N_9864);
xnor U10939 (N_10939,N_9875,N_8552);
or U10940 (N_10940,N_8648,N_8173);
xor U10941 (N_10941,N_8982,N_7962);
or U10942 (N_10942,N_7015,N_5793);
nand U10943 (N_10943,N_9559,N_5330);
nor U10944 (N_10944,N_5496,N_6802);
and U10945 (N_10945,N_8404,N_5179);
or U10946 (N_10946,N_6315,N_8178);
and U10947 (N_10947,N_6874,N_5450);
xnor U10948 (N_10948,N_9708,N_5069);
xnor U10949 (N_10949,N_6262,N_9053);
and U10950 (N_10950,N_8887,N_8994);
or U10951 (N_10951,N_5157,N_5775);
or U10952 (N_10952,N_7111,N_6877);
nand U10953 (N_10953,N_5035,N_6051);
and U10954 (N_10954,N_7442,N_6205);
and U10955 (N_10955,N_7672,N_8688);
or U10956 (N_10956,N_9642,N_5434);
and U10957 (N_10957,N_5140,N_7150);
or U10958 (N_10958,N_6411,N_6120);
xnor U10959 (N_10959,N_5594,N_7558);
or U10960 (N_10960,N_6377,N_8457);
or U10961 (N_10961,N_8465,N_9013);
nor U10962 (N_10962,N_6633,N_5469);
or U10963 (N_10963,N_6290,N_5359);
nor U10964 (N_10964,N_6484,N_8772);
nand U10965 (N_10965,N_8278,N_5158);
nand U10966 (N_10966,N_6657,N_6524);
or U10967 (N_10967,N_8368,N_7262);
xnor U10968 (N_10968,N_7013,N_9695);
and U10969 (N_10969,N_7639,N_9208);
and U10970 (N_10970,N_7241,N_8274);
nand U10971 (N_10971,N_8433,N_6925);
xnor U10972 (N_10972,N_7607,N_8265);
xnor U10973 (N_10973,N_7584,N_6424);
and U10974 (N_10974,N_5217,N_8081);
nand U10975 (N_10975,N_8308,N_9015);
nor U10976 (N_10976,N_7358,N_8251);
nor U10977 (N_10977,N_5362,N_7793);
nor U10978 (N_10978,N_8852,N_9540);
nor U10979 (N_10979,N_9720,N_8805);
nor U10980 (N_10980,N_5627,N_9977);
nand U10981 (N_10981,N_9765,N_8824);
or U10982 (N_10982,N_8588,N_6885);
nand U10983 (N_10983,N_5210,N_9355);
or U10984 (N_10984,N_9399,N_5925);
nand U10985 (N_10985,N_9957,N_7739);
and U10986 (N_10986,N_7110,N_7606);
nand U10987 (N_10987,N_8495,N_9159);
xor U10988 (N_10988,N_6596,N_5888);
nor U10989 (N_10989,N_9468,N_9920);
and U10990 (N_10990,N_9427,N_8303);
nor U10991 (N_10991,N_7089,N_5801);
xor U10992 (N_10992,N_8407,N_9832);
nand U10993 (N_10993,N_7884,N_8757);
or U10994 (N_10994,N_9463,N_7011);
nor U10995 (N_10995,N_6789,N_5907);
and U10996 (N_10996,N_8095,N_6393);
and U10997 (N_10997,N_8379,N_6447);
nor U10998 (N_10998,N_5357,N_7469);
nor U10999 (N_10999,N_6033,N_5211);
nor U11000 (N_11000,N_6300,N_8998);
xnor U11001 (N_11001,N_7627,N_7663);
nand U11002 (N_11002,N_5929,N_9291);
nor U11003 (N_11003,N_8926,N_7480);
and U11004 (N_11004,N_6635,N_6559);
xnor U11005 (N_11005,N_5057,N_5480);
and U11006 (N_11006,N_8518,N_7490);
and U11007 (N_11007,N_7338,N_9462);
or U11008 (N_11008,N_7239,N_6745);
and U11009 (N_11009,N_6935,N_8408);
nor U11010 (N_11010,N_6717,N_7048);
xnor U11011 (N_11011,N_8523,N_5136);
nor U11012 (N_11012,N_9449,N_7486);
nor U11013 (N_11013,N_7514,N_6403);
xor U11014 (N_11014,N_7206,N_8569);
nor U11015 (N_11015,N_7199,N_5448);
and U11016 (N_11016,N_8738,N_7156);
xor U11017 (N_11017,N_8056,N_5266);
nor U11018 (N_11018,N_7256,N_9384);
or U11019 (N_11019,N_6391,N_9493);
nand U11020 (N_11020,N_9163,N_7428);
nand U11021 (N_11021,N_9063,N_5694);
xnor U11022 (N_11022,N_7631,N_6224);
xnor U11023 (N_11023,N_7187,N_5251);
nor U11024 (N_11024,N_5589,N_5307);
and U11025 (N_11025,N_5371,N_7451);
or U11026 (N_11026,N_5309,N_7409);
nand U11027 (N_11027,N_7602,N_6140);
and U11028 (N_11028,N_8363,N_5216);
and U11029 (N_11029,N_9779,N_7252);
xnor U11030 (N_11030,N_8953,N_5088);
and U11031 (N_11031,N_6383,N_9980);
xor U11032 (N_11032,N_5412,N_5101);
or U11033 (N_11033,N_7379,N_5339);
nand U11034 (N_11034,N_7567,N_9718);
or U11035 (N_11035,N_7913,N_6034);
xor U11036 (N_11036,N_8439,N_8521);
xor U11037 (N_11037,N_6879,N_6735);
and U11038 (N_11038,N_5515,N_7553);
and U11039 (N_11039,N_8833,N_7387);
and U11040 (N_11040,N_9821,N_8245);
or U11041 (N_11041,N_8560,N_6746);
or U11042 (N_11042,N_7573,N_6507);
nand U11043 (N_11043,N_9807,N_8758);
nor U11044 (N_11044,N_6528,N_9738);
and U11045 (N_11045,N_6787,N_7398);
xor U11046 (N_11046,N_8420,N_6075);
nand U11047 (N_11047,N_9289,N_9253);
xnor U11048 (N_11048,N_8929,N_9061);
nand U11049 (N_11049,N_8068,N_7856);
or U11050 (N_11050,N_7621,N_5722);
nor U11051 (N_11051,N_9723,N_5954);
and U11052 (N_11052,N_8289,N_9342);
xor U11053 (N_11053,N_6537,N_5479);
nor U11054 (N_11054,N_6621,N_6693);
and U11055 (N_11055,N_9328,N_6064);
or U11056 (N_11056,N_6508,N_6957);
nand U11057 (N_11057,N_7706,N_5876);
xnor U11058 (N_11058,N_7145,N_5875);
nor U11059 (N_11059,N_9454,N_6558);
nand U11060 (N_11060,N_5555,N_9120);
nand U11061 (N_11061,N_8471,N_7530);
xnor U11062 (N_11062,N_9950,N_5253);
or U11063 (N_11063,N_6337,N_7395);
nor U11064 (N_11064,N_8751,N_6322);
nand U11065 (N_11065,N_9958,N_5048);
or U11066 (N_11066,N_5236,N_9699);
xnor U11067 (N_11067,N_7029,N_5517);
nor U11068 (N_11068,N_8072,N_8932);
xor U11069 (N_11069,N_5289,N_7374);
or U11070 (N_11070,N_9176,N_9585);
and U11071 (N_11071,N_7629,N_6638);
nor U11072 (N_11072,N_6817,N_8879);
or U11073 (N_11073,N_6773,N_9834);
nand U11074 (N_11074,N_5506,N_7473);
or U11075 (N_11075,N_9099,N_6132);
and U11076 (N_11076,N_5182,N_8463);
or U11077 (N_11077,N_9777,N_5340);
or U11078 (N_11078,N_7228,N_6541);
nor U11079 (N_11079,N_7106,N_8228);
and U11080 (N_11080,N_6486,N_8119);
nand U11081 (N_11081,N_8235,N_8541);
xnor U11082 (N_11082,N_9549,N_9952);
or U11083 (N_11083,N_6965,N_5634);
nand U11084 (N_11084,N_7020,N_5102);
nand U11085 (N_11085,N_9946,N_7378);
and U11086 (N_11086,N_7714,N_7026);
nor U11087 (N_11087,N_7211,N_7646);
or U11088 (N_11088,N_7055,N_5265);
and U11089 (N_11089,N_6169,N_5719);
nor U11090 (N_11090,N_9199,N_8171);
nor U11091 (N_11091,N_7419,N_9701);
or U11092 (N_11092,N_9824,N_9657);
nand U11093 (N_11093,N_8373,N_8434);
xor U11094 (N_11094,N_9168,N_9897);
nor U11095 (N_11095,N_7588,N_9769);
nor U11096 (N_11096,N_8813,N_5130);
nand U11097 (N_11097,N_5238,N_8717);
xnor U11098 (N_11098,N_7144,N_8945);
and U11099 (N_11099,N_9387,N_9178);
or U11100 (N_11100,N_6900,N_6532);
xnor U11101 (N_11101,N_8678,N_7452);
xor U11102 (N_11102,N_9382,N_6191);
xnor U11103 (N_11103,N_8646,N_8113);
xnor U11104 (N_11104,N_9184,N_6266);
nor U11105 (N_11105,N_9593,N_5246);
xor U11106 (N_11106,N_6444,N_6721);
and U11107 (N_11107,N_8583,N_8030);
and U11108 (N_11108,N_5885,N_9411);
nor U11109 (N_11109,N_7626,N_9562);
or U11110 (N_11110,N_9389,N_6926);
nor U11111 (N_11111,N_5829,N_5806);
nand U11112 (N_11112,N_7804,N_6909);
xor U11113 (N_11113,N_9127,N_6327);
and U11114 (N_11114,N_9234,N_7832);
nor U11115 (N_11115,N_8513,N_5190);
nor U11116 (N_11116,N_6493,N_7101);
xor U11117 (N_11117,N_6628,N_6676);
and U11118 (N_11118,N_6387,N_9109);
and U11119 (N_11119,N_6659,N_5560);
and U11120 (N_11120,N_9996,N_8271);
nand U11121 (N_11121,N_5025,N_8973);
and U11122 (N_11122,N_8938,N_6273);
nand U11123 (N_11123,N_6466,N_7596);
and U11124 (N_11124,N_7191,N_9241);
or U11125 (N_11125,N_9251,N_6341);
or U11126 (N_11126,N_8862,N_9301);
xnor U11127 (N_11127,N_7234,N_9445);
nor U11128 (N_11128,N_6708,N_8020);
or U11129 (N_11129,N_6326,N_8418);
or U11130 (N_11130,N_8831,N_7705);
nor U11131 (N_11131,N_8176,N_7609);
or U11132 (N_11132,N_6118,N_7696);
or U11133 (N_11133,N_8715,N_8302);
nand U11134 (N_11134,N_8707,N_6557);
and U11135 (N_11135,N_7070,N_7581);
or U11136 (N_11136,N_9206,N_9800);
xnor U11137 (N_11137,N_5682,N_6733);
nor U11138 (N_11138,N_7544,N_7998);
nor U11139 (N_11139,N_9829,N_8461);
nor U11140 (N_11140,N_6020,N_6764);
nand U11141 (N_11141,N_6039,N_8816);
nor U11142 (N_11142,N_8292,N_5053);
nand U11143 (N_11143,N_7468,N_8029);
and U11144 (N_11144,N_5218,N_6150);
nand U11145 (N_11145,N_8437,N_8628);
xor U11146 (N_11146,N_9239,N_5903);
xnor U11147 (N_11147,N_7829,N_9768);
or U11148 (N_11148,N_8282,N_7537);
nand U11149 (N_11149,N_8220,N_7830);
xor U11150 (N_11150,N_5044,N_5702);
and U11151 (N_11151,N_7858,N_6540);
nand U11152 (N_11152,N_6866,N_8198);
and U11153 (N_11153,N_8182,N_9605);
and U11154 (N_11154,N_5235,N_8035);
or U11155 (N_11155,N_6604,N_6483);
nand U11156 (N_11156,N_7493,N_5607);
or U11157 (N_11157,N_5557,N_7958);
and U11158 (N_11158,N_7525,N_7644);
nor U11159 (N_11159,N_9474,N_7877);
nand U11160 (N_11160,N_9192,N_8706);
and U11161 (N_11161,N_7445,N_6941);
or U11162 (N_11162,N_9007,N_5392);
xor U11163 (N_11163,N_8066,N_7103);
xor U11164 (N_11164,N_5056,N_5122);
or U11165 (N_11165,N_5173,N_5382);
nand U11166 (N_11166,N_8914,N_8893);
and U11167 (N_11167,N_5615,N_6517);
nand U11168 (N_11168,N_9164,N_7600);
or U11169 (N_11169,N_7557,N_9467);
nor U11170 (N_11170,N_8672,N_5712);
or U11171 (N_11171,N_7107,N_5134);
nor U11172 (N_11172,N_8915,N_9457);
nor U11173 (N_11173,N_8291,N_9784);
nand U11174 (N_11174,N_7746,N_9630);
nor U11175 (N_11175,N_9358,N_8486);
xor U11176 (N_11176,N_9604,N_8338);
nor U11177 (N_11177,N_9310,N_9456);
xor U11178 (N_11178,N_5815,N_6901);
xor U11179 (N_11179,N_9798,N_8542);
and U11180 (N_11180,N_6575,N_5860);
nor U11181 (N_11181,N_9548,N_5204);
or U11182 (N_11182,N_7808,N_5424);
nand U11183 (N_11183,N_6368,N_9635);
or U11184 (N_11184,N_9970,N_9132);
nand U11185 (N_11185,N_8451,N_7258);
nand U11186 (N_11186,N_8405,N_7980);
nor U11187 (N_11187,N_7303,N_9152);
and U11188 (N_11188,N_5983,N_7401);
nor U11189 (N_11189,N_8762,N_9674);
nand U11190 (N_11190,N_7691,N_5279);
nor U11191 (N_11191,N_5263,N_8116);
and U11192 (N_11192,N_7694,N_8943);
and U11193 (N_11193,N_5705,N_7659);
or U11194 (N_11194,N_9235,N_5332);
and U11195 (N_11195,N_5990,N_6282);
or U11196 (N_11196,N_7453,N_8832);
and U11197 (N_11197,N_8501,N_6179);
nand U11198 (N_11198,N_7440,N_9141);
or U11199 (N_11199,N_6854,N_8252);
nor U11200 (N_11200,N_7899,N_7169);
nor U11201 (N_11201,N_7664,N_5421);
nor U11202 (N_11202,N_8891,N_6154);
nand U11203 (N_11203,N_7432,N_6043);
and U11204 (N_11204,N_5272,N_9940);
xor U11205 (N_11205,N_8668,N_8713);
and U11206 (N_11206,N_7509,N_7729);
or U11207 (N_11207,N_7961,N_7908);
and U11208 (N_11208,N_7844,N_7891);
or U11209 (N_11209,N_8747,N_8960);
or U11210 (N_11210,N_7989,N_6731);
nor U11211 (N_11211,N_5388,N_7986);
xor U11212 (N_11212,N_5400,N_5084);
nand U11213 (N_11213,N_5275,N_5452);
nand U11214 (N_11214,N_8967,N_8336);
or U11215 (N_11215,N_7038,N_6183);
and U11216 (N_11216,N_6135,N_5449);
nand U11217 (N_11217,N_9260,N_5717);
and U11218 (N_11218,N_8589,N_5313);
nor U11219 (N_11219,N_7517,N_6534);
nand U11220 (N_11220,N_6625,N_5548);
nand U11221 (N_11221,N_7272,N_5533);
or U11222 (N_11222,N_5768,N_5111);
and U11223 (N_11223,N_5194,N_5206);
and U11224 (N_11224,N_8156,N_5562);
and U11225 (N_11225,N_6481,N_7041);
nor U11226 (N_11226,N_9568,N_7498);
or U11227 (N_11227,N_6161,N_7091);
and U11228 (N_11228,N_8195,N_7213);
nor U11229 (N_11229,N_5789,N_5813);
or U11230 (N_11230,N_9022,N_5595);
xor U11231 (N_11231,N_6685,N_7470);
nand U11232 (N_11232,N_5186,N_5029);
xnor U11233 (N_11233,N_7860,N_8256);
xor U11234 (N_11234,N_7778,N_7817);
nand U11235 (N_11235,N_6862,N_9752);
or U11236 (N_11236,N_8997,N_6798);
nand U11237 (N_11237,N_9710,N_9801);
and U11238 (N_11238,N_9221,N_9264);
xor U11239 (N_11239,N_9783,N_9842);
xnor U11240 (N_11240,N_6175,N_6141);
nand U11241 (N_11241,N_6858,N_9648);
xnor U11242 (N_11242,N_9172,N_9911);
or U11243 (N_11243,N_5131,N_9442);
and U11244 (N_11244,N_7130,N_7219);
nor U11245 (N_11245,N_8705,N_9561);
xnor U11246 (N_11246,N_9979,N_7511);
or U11247 (N_11247,N_6306,N_7138);
or U11248 (N_11248,N_5335,N_5809);
and U11249 (N_11249,N_7482,N_8150);
nand U11250 (N_11250,N_6549,N_5367);
xor U11251 (N_11251,N_5451,N_7488);
and U11252 (N_11252,N_6963,N_9904);
nand U11253 (N_11253,N_5667,N_8562);
xor U11254 (N_11254,N_5433,N_9574);
nor U11255 (N_11255,N_5523,N_5926);
nand U11256 (N_11256,N_8444,N_8337);
or U11257 (N_11257,N_8015,N_9200);
nand U11258 (N_11258,N_6450,N_9466);
and U11259 (N_11259,N_7356,N_6906);
nand U11260 (N_11260,N_5590,N_9782);
or U11261 (N_11261,N_7887,N_5350);
nor U11262 (N_11262,N_6482,N_6709);
nor U11263 (N_11263,N_8117,N_7643);
and U11264 (N_11264,N_6954,N_7907);
or U11265 (N_11265,N_6121,N_8724);
nor U11266 (N_11266,N_8120,N_6385);
and U11267 (N_11267,N_8949,N_6973);
and U11268 (N_11268,N_5233,N_8819);
xnor U11269 (N_11269,N_6846,N_7642);
xnor U11270 (N_11270,N_8159,N_9704);
or U11271 (N_11271,N_8320,N_8730);
or U11272 (N_11272,N_5395,N_6219);
or U11273 (N_11273,N_8733,N_6091);
nor U11274 (N_11274,N_7721,N_8249);
or U11275 (N_11275,N_8825,N_7781);
and U11276 (N_11276,N_7896,N_6845);
or U11277 (N_11277,N_9390,N_6777);
nand U11278 (N_11278,N_5863,N_9207);
xor U11279 (N_11279,N_7543,N_7443);
xor U11280 (N_11280,N_7571,N_6189);
nand U11281 (N_11281,N_9285,N_9542);
xnor U11282 (N_11282,N_6968,N_7610);
nand U11283 (N_11283,N_8684,N_7917);
xor U11284 (N_11284,N_9671,N_6561);
nor U11285 (N_11285,N_7704,N_7979);
and U11286 (N_11286,N_5967,N_8174);
xnor U11287 (N_11287,N_5553,N_6520);
nor U11288 (N_11288,N_6052,N_5199);
nand U11289 (N_11289,N_7590,N_7153);
or U11290 (N_11290,N_5912,N_8838);
nand U11291 (N_11291,N_5114,N_6074);
xor U11292 (N_11292,N_6911,N_6076);
nor U11293 (N_11293,N_8357,N_9578);
and U11294 (N_11294,N_6465,N_9703);
or U11295 (N_11295,N_5387,N_5854);
nor U11296 (N_11296,N_6230,N_8788);
xnor U11297 (N_11297,N_5941,N_7710);
or U11298 (N_11298,N_8435,N_5282);
nor U11299 (N_11299,N_7035,N_8221);
or U11300 (N_11300,N_7068,N_9571);
xor U11301 (N_11301,N_8047,N_7523);
or U11302 (N_11302,N_5853,N_8466);
or U11303 (N_11303,N_5992,N_8273);
and U11304 (N_11304,N_5345,N_9894);
xor U11305 (N_11305,N_9284,N_5311);
and U11306 (N_11306,N_5706,N_5649);
nand U11307 (N_11307,N_6138,N_6158);
or U11308 (N_11308,N_6671,N_8402);
nand U11309 (N_11309,N_9740,N_6505);
nand U11310 (N_11310,N_8806,N_5895);
nand U11311 (N_11311,N_6172,N_6969);
and U11312 (N_11312,N_9576,N_7345);
or U11313 (N_11313,N_8121,N_6458);
xnor U11314 (N_11314,N_7637,N_5856);
and U11315 (N_11315,N_8610,N_5242);
nand U11316 (N_11316,N_8911,N_5997);
or U11317 (N_11317,N_5123,N_9497);
and U11318 (N_11318,N_6238,N_9503);
or U11319 (N_11319,N_8649,N_7845);
nand U11320 (N_11320,N_9563,N_5146);
nand U11321 (N_11321,N_8477,N_5684);
and U11322 (N_11322,N_8616,N_9572);
nor U11323 (N_11323,N_5619,N_5073);
or U11324 (N_11324,N_5571,N_8919);
nand U11325 (N_11325,N_7355,N_9123);
or U11326 (N_11326,N_5352,N_5841);
nand U11327 (N_11327,N_6429,N_5503);
nor U11328 (N_11328,N_5871,N_6587);
and U11329 (N_11329,N_6330,N_7702);
or U11330 (N_11330,N_7386,N_5746);
and U11331 (N_11331,N_5369,N_6988);
xor U11332 (N_11332,N_8456,N_6781);
xnor U11333 (N_11333,N_9717,N_9712);
and U11334 (N_11334,N_9746,N_6594);
xnor U11335 (N_11335,N_8470,N_8143);
xnor U11336 (N_11336,N_7224,N_6582);
and U11337 (N_11337,N_6719,N_5927);
xnor U11338 (N_11338,N_9097,N_7472);
nor U11339 (N_11339,N_5135,N_9198);
nor U11340 (N_11340,N_6898,N_6196);
nor U11341 (N_11341,N_6578,N_7220);
xnor U11342 (N_11342,N_8535,N_7507);
nand U11343 (N_11343,N_9272,N_6023);
or U11344 (N_11344,N_5165,N_6536);
and U11345 (N_11345,N_7065,N_6288);
nand U11346 (N_11346,N_8359,N_7938);
xor U11347 (N_11347,N_7090,N_7786);
and U11348 (N_11348,N_9652,N_7870);
nand U11349 (N_11349,N_7859,N_8794);
xnor U11350 (N_11350,N_9565,N_5518);
or U11351 (N_11351,N_5476,N_6818);
nor U11352 (N_11352,N_5918,N_7939);
nand U11353 (N_11353,N_8321,N_6256);
nor U11354 (N_11354,N_5945,N_7894);
nor U11355 (N_11355,N_5655,N_7872);
nand U11356 (N_11356,N_5482,N_6407);
and U11357 (N_11357,N_5104,N_6678);
nand U11358 (N_11358,N_9557,N_6955);
and U11359 (N_11359,N_6915,N_5325);
nand U11360 (N_11360,N_6894,N_6139);
xnor U11361 (N_11361,N_5942,N_5346);
nand U11362 (N_11362,N_6960,N_8714);
or U11363 (N_11363,N_8089,N_7112);
nand U11364 (N_11364,N_5955,N_6538);
nor U11365 (N_11365,N_7570,N_5127);
xnor U11366 (N_11366,N_6792,N_7734);
xor U11367 (N_11367,N_5672,N_8417);
or U11368 (N_11368,N_9263,N_6521);
or U11369 (N_11369,N_6276,N_6012);
xor U11370 (N_11370,N_6359,N_9237);
and U11371 (N_11371,N_9989,N_9883);
xnor U11372 (N_11372,N_9071,N_7137);
or U11373 (N_11373,N_6311,N_9005);
xor U11374 (N_11374,N_8544,N_5028);
and U11375 (N_11375,N_7601,N_8290);
or U11376 (N_11376,N_5301,N_9887);
xnor U11377 (N_11377,N_6525,N_7444);
xnor U11378 (N_11378,N_6841,N_7168);
or U11379 (N_11379,N_8358,N_7640);
nor U11380 (N_11380,N_5638,N_9700);
nor U11381 (N_11381,N_8665,N_7180);
nand U11382 (N_11382,N_5878,N_5294);
nor U11383 (N_11383,N_8267,N_7634);
nor U11384 (N_11384,N_7388,N_7540);
xor U11385 (N_11385,N_5059,N_8092);
or U11386 (N_11386,N_6668,N_5090);
xnor U11387 (N_11387,N_5567,N_5777);
xor U11388 (N_11388,N_9110,N_5372);
nor U11389 (N_11389,N_9917,N_6716);
nor U11390 (N_11390,N_7365,N_9327);
nand U11391 (N_11391,N_8902,N_9218);
nand U11392 (N_11392,N_9998,N_7747);
nand U11393 (N_11393,N_5376,N_5920);
xnor U11394 (N_11394,N_7434,N_5318);
nor U11395 (N_11395,N_8619,N_8013);
nand U11396 (N_11396,N_8681,N_5580);
nor U11397 (N_11397,N_6710,N_7999);
or U11398 (N_11398,N_9614,N_5531);
xor U11399 (N_11399,N_9425,N_7411);
and U11400 (N_11400,N_7074,N_7499);
xnor U11401 (N_11401,N_8985,N_5062);
and U11402 (N_11402,N_7732,N_9096);
nand U11403 (N_11403,N_8350,N_6606);
or U11404 (N_11404,N_8101,N_7474);
and U11405 (N_11405,N_7948,N_5317);
nor U11406 (N_11406,N_8948,N_5887);
nor U11407 (N_11407,N_8841,N_8006);
xnor U11408 (N_11408,N_8044,N_6749);
nand U11409 (N_11409,N_6831,N_9320);
nand U11410 (N_11410,N_7944,N_9103);
or U11411 (N_11411,N_5735,N_6714);
nor U11412 (N_11412,N_6367,N_7190);
nand U11413 (N_11413,N_7030,N_9532);
xnor U11414 (N_11414,N_7812,N_5662);
xnor U11415 (N_11415,N_5356,N_9490);
nand U11416 (N_11416,N_9036,N_5232);
nor U11417 (N_11417,N_7791,N_9598);
or U11418 (N_11418,N_9513,N_6299);
or U11419 (N_11419,N_8313,N_5893);
xnor U11420 (N_11420,N_5616,N_5718);
or U11421 (N_11421,N_8689,N_6267);
nand U11422 (N_11422,N_7447,N_8472);
xnor U11423 (N_11423,N_6824,N_7628);
nor U11424 (N_11424,N_9416,N_6675);
nand U11425 (N_11425,N_8294,N_6050);
xor U11426 (N_11426,N_6294,N_7519);
or U11427 (N_11427,N_9960,N_5229);
xnor U11428 (N_11428,N_7316,N_7837);
nand U11429 (N_11429,N_8494,N_8246);
and U11430 (N_11430,N_6934,N_9647);
and U11431 (N_11431,N_6214,N_8155);
nand U11432 (N_11432,N_7783,N_5319);
or U11433 (N_11433,N_8300,N_7385);
nor U11434 (N_11434,N_5519,N_8096);
xnor U11435 (N_11435,N_7554,N_8899);
or U11436 (N_11436,N_8885,N_7761);
nand U11437 (N_11437,N_9489,N_6687);
nor U11438 (N_11438,N_9981,N_9451);
or U11439 (N_11439,N_6550,N_7502);
nor U11440 (N_11440,N_5470,N_6873);
nor U11441 (N_11441,N_7678,N_5432);
and U11442 (N_11442,N_5467,N_7282);
xnor U11443 (N_11443,N_7826,N_7843);
or U11444 (N_11444,N_6264,N_5674);
nor U11445 (N_11445,N_8693,N_6990);
nand U11446 (N_11446,N_5668,N_8318);
nand U11447 (N_11447,N_5379,N_9609);
or U11448 (N_11448,N_6839,N_5507);
xor U11449 (N_11449,N_8817,N_8132);
nand U11450 (N_11450,N_5273,N_9436);
or U11451 (N_11451,N_6369,N_6108);
xnor U11452 (N_11452,N_8353,N_9129);
nand U11453 (N_11453,N_8663,N_5936);
and U11454 (N_11454,N_7946,N_9558);
and U11455 (N_11455,N_8234,N_6389);
nand U11456 (N_11456,N_6816,N_5758);
nor U11457 (N_11457,N_7769,N_8342);
and U11458 (N_11458,N_7161,N_7448);
nand U11459 (N_11459,N_6649,N_8796);
xor U11460 (N_11460,N_8395,N_5049);
or U11461 (N_11461,N_9644,N_7871);
and U11462 (N_11462,N_6342,N_9429);
or U11463 (N_11463,N_5794,N_6073);
nand U11464 (N_11464,N_5264,N_9935);
or U11465 (N_11465,N_9491,N_8520);
xor U11466 (N_11466,N_6661,N_9000);
or U11467 (N_11467,N_8870,N_9905);
xnor U11468 (N_11468,N_7094,N_7066);
xor U11469 (N_11469,N_9848,N_8060);
or U11470 (N_11470,N_7717,N_8343);
or U11471 (N_11471,N_6826,N_5541);
xor U11472 (N_11472,N_9068,N_9347);
and U11473 (N_11473,N_9677,N_5070);
and U11474 (N_11474,N_9566,N_9551);
nand U11475 (N_11475,N_7088,N_7597);
and U11476 (N_11476,N_5268,N_9273);
nor U11477 (N_11477,N_9923,N_9692);
nand U11478 (N_11478,N_6063,N_6007);
nand U11479 (N_11479,N_6347,N_8255);
xnor U11480 (N_11480,N_8574,N_9759);
and U11481 (N_11481,N_6155,N_5838);
or U11482 (N_11482,N_5583,N_8732);
nand U11483 (N_11483,N_6243,N_5013);
nor U11484 (N_11484,N_7556,N_7384);
xnor U11485 (N_11485,N_6394,N_7785);
xor U11486 (N_11486,N_6778,N_7022);
or U11487 (N_11487,N_9541,N_8903);
or U11488 (N_11488,N_9514,N_5215);
or U11489 (N_11489,N_8430,N_8861);
xnor U11490 (N_11490,N_7056,N_5133);
nor U11491 (N_11491,N_7692,N_6350);
xor U11492 (N_11492,N_6086,N_8391);
nand U11493 (N_11493,N_8942,N_8146);
nor U11494 (N_11494,N_7866,N_5071);
nand U11495 (N_11495,N_8100,N_9662);
nand U11496 (N_11496,N_9326,N_7172);
nand U11497 (N_11497,N_8549,N_7565);
nor U11498 (N_11498,N_9089,N_7875);
nor U11499 (N_11499,N_9617,N_5625);
or U11500 (N_11500,N_6097,N_8889);
nor U11501 (N_11501,N_9537,N_6702);
or U11502 (N_11502,N_7542,N_8976);
and U11503 (N_11503,N_9956,N_9348);
nand U11504 (N_11504,N_6562,N_9121);
nand U11505 (N_11505,N_8575,N_9331);
nor U11506 (N_11506,N_8186,N_9133);
and U11507 (N_11507,N_5171,N_8284);
nor U11508 (N_11508,N_5305,N_7463);
and U11509 (N_11509,N_6113,N_7354);
nor U11510 (N_11510,N_8837,N_8627);
or U11511 (N_11511,N_8210,N_8270);
nor U11512 (N_11512,N_7660,N_5822);
xor U11513 (N_11513,N_7349,N_9209);
or U11514 (N_11514,N_6526,N_7806);
and U11515 (N_11515,N_6048,N_8423);
or U11516 (N_11516,N_5611,N_9939);
or U11517 (N_11517,N_5154,N_9338);
and U11518 (N_11518,N_8851,N_7712);
nand U11519 (N_11519,N_5024,N_6739);
nand U11520 (N_11520,N_8051,N_6715);
and U11521 (N_11521,N_5076,N_9581);
nor U11522 (N_11522,N_8406,N_5408);
nand U11523 (N_11523,N_6748,N_6240);
or U11524 (N_11524,N_7465,N_9370);
or U11525 (N_11525,N_5810,N_6397);
xnor U11526 (N_11526,N_9504,N_9786);
and U11527 (N_11527,N_5636,N_8253);
or U11528 (N_11528,N_5783,N_7966);
and U11529 (N_11529,N_5959,N_8966);
and U11530 (N_11530,N_5196,N_5894);
or U11531 (N_11531,N_6320,N_5739);
nand U11532 (N_11532,N_6269,N_5520);
nand U11533 (N_11533,N_5097,N_7593);
and U11534 (N_11534,N_5899,N_6869);
xnor U11535 (N_11535,N_7764,N_5398);
nand U11536 (N_11536,N_5151,N_7181);
and U11537 (N_11537,N_6479,N_5132);
xnor U11538 (N_11538,N_6852,N_6498);
nor U11539 (N_11539,N_9811,N_9774);
xor U11540 (N_11540,N_5943,N_6451);
xor U11541 (N_11541,N_5774,N_5977);
nand U11542 (N_11542,N_9204,N_7670);
nor U11543 (N_11543,N_8438,N_6068);
xnor U11544 (N_11544,N_7698,N_8490);
xnor U11545 (N_11545,N_5137,N_6940);
or U11546 (N_11546,N_8866,N_8954);
xnor U11547 (N_11547,N_7929,N_9450);
nor U11548 (N_11548,N_9964,N_6250);
and U11549 (N_11549,N_8197,N_6441);
xor U11550 (N_11550,N_8293,N_9006);
or U11551 (N_11551,N_9954,N_5650);
nor U11552 (N_11552,N_5740,N_7709);
nand U11553 (N_11553,N_9624,N_9817);
xnor U11554 (N_11554,N_5837,N_9870);
and U11555 (N_11555,N_8022,N_7656);
nand U11556 (N_11556,N_8448,N_9487);
xor U11557 (N_11557,N_9359,N_5839);
nor U11558 (N_11558,N_6815,N_8907);
and U11559 (N_11559,N_9148,N_5037);
and U11560 (N_11560,N_5108,N_5299);
xor U11561 (N_11561,N_8436,N_9078);
or U11562 (N_11562,N_6233,N_7772);
nand U11563 (N_11563,N_6729,N_9242);
xor U11564 (N_11564,N_9685,N_9051);
nand U11565 (N_11565,N_9018,N_8847);
xnor U11566 (N_11566,N_7429,N_5481);
nor U11567 (N_11567,N_8459,N_7148);
nand U11568 (N_11568,N_8335,N_8988);
nand U11569 (N_11569,N_8754,N_8449);
and U11570 (N_11570,N_6035,N_7308);
and U11571 (N_11571,N_9374,N_9886);
nand U11572 (N_11572,N_6722,N_7147);
nand U11573 (N_11573,N_6814,N_6679);
nor U11574 (N_11574,N_8360,N_5730);
nor U11575 (N_11575,N_7081,N_8394);
nand U11576 (N_11576,N_7491,N_7869);
xnor U11577 (N_11577,N_6129,N_8771);
and U11578 (N_11578,N_8219,N_8301);
nor U11579 (N_11579,N_5415,N_9930);
and U11580 (N_11580,N_5292,N_9803);
xnor U11581 (N_11581,N_9925,N_6105);
nor U11582 (N_11582,N_8510,N_8971);
nor U11583 (N_11583,N_7368,N_8375);
nand U11584 (N_11584,N_6500,N_6913);
nor U11585 (N_11585,N_9835,N_8189);
and U11586 (N_11586,N_6751,N_8453);
nand U11587 (N_11587,N_8147,N_7931);
or U11588 (N_11588,N_5656,N_5949);
xor U11589 (N_11589,N_8565,N_7648);
and U11590 (N_11590,N_6905,N_8592);
nand U11591 (N_11591,N_7561,N_9447);
nand U11592 (N_11592,N_7924,N_8037);
and U11593 (N_11593,N_6430,N_5683);
nor U11594 (N_11594,N_8516,N_9441);
nor U11595 (N_11595,N_8328,N_6056);
xnor U11596 (N_11596,N_5924,N_7140);
nor U11597 (N_11597,N_5399,N_8104);
nor U11598 (N_11598,N_7700,N_7157);
xor U11599 (N_11599,N_9944,N_8604);
nand U11600 (N_11600,N_5105,N_9243);
nand U11601 (N_11601,N_5647,N_5877);
nor U11602 (N_11602,N_9682,N_7773);
xnor U11603 (N_11603,N_7974,N_9043);
nor U11604 (N_11604,N_8622,N_9197);
nor U11605 (N_11605,N_9852,N_8263);
nor U11606 (N_11606,N_9188,N_5499);
xnor U11607 (N_11607,N_5493,N_8981);
nand U11608 (N_11608,N_7031,N_5030);
nand U11609 (N_11609,N_5410,N_5001);
or U11610 (N_11610,N_8384,N_8112);
xnor U11611 (N_11611,N_8636,N_7745);
and U11612 (N_11612,N_5180,N_5161);
nand U11613 (N_11613,N_6316,N_6004);
xnor U11614 (N_11614,N_5348,N_8863);
or U11615 (N_11615,N_6314,N_9851);
and U11616 (N_11616,N_9191,N_5004);
nor U11617 (N_11617,N_6908,N_8768);
nor U11618 (N_11618,N_6229,N_8509);
nor U11619 (N_11619,N_6518,N_5665);
or U11620 (N_11620,N_8578,N_8815);
and U11621 (N_11621,N_7842,N_9039);
xor U11622 (N_11622,N_5773,N_7657);
or U11623 (N_11623,N_9600,N_8667);
nand U11624 (N_11624,N_5660,N_8923);
nor U11625 (N_11625,N_9985,N_5139);
nand U11626 (N_11626,N_9232,N_8687);
xnor U11627 (N_11627,N_8970,N_8003);
or U11628 (N_11628,N_8526,N_6144);
and U11629 (N_11629,N_9967,N_5971);
nand U11630 (N_11630,N_5715,N_9791);
or U11631 (N_11631,N_6980,N_7008);
and U11632 (N_11632,N_5559,N_7674);
xnor U11633 (N_11633,N_7926,N_6570);
or U11634 (N_11634,N_9137,N_9045);
nand U11635 (N_11635,N_6225,N_9742);
or U11636 (N_11636,N_8499,N_9229);
nand U11637 (N_11637,N_9607,N_7688);
xnor U11638 (N_11638,N_7562,N_9857);
nor U11639 (N_11639,N_8605,N_9649);
and U11640 (N_11640,N_7210,N_8009);
or U11641 (N_11641,N_9255,N_5504);
xor U11642 (N_11642,N_5177,N_5081);
nand U11643 (N_11643,N_9057,N_6887);
or U11644 (N_11644,N_6049,N_6987);
nand U11645 (N_11645,N_7620,N_9380);
nor U11646 (N_11646,N_5221,N_7115);
or U11647 (N_11647,N_6805,N_5532);
xnor U11648 (N_11648,N_9288,N_6847);
nor U11649 (N_11649,N_5609,N_8305);
nand U11650 (N_11650,N_9902,N_6886);
xnor U11651 (N_11651,N_9396,N_8856);
nand U11652 (N_11652,N_5344,N_6460);
or U11653 (N_11653,N_6663,N_9736);
or U11654 (N_11654,N_8014,N_6836);
or U11655 (N_11655,N_9529,N_7497);
and U11656 (N_11656,N_8682,N_5998);
or U11657 (N_11657,N_7017,N_5422);
nand U11658 (N_11658,N_8807,N_6759);
or U11659 (N_11659,N_8247,N_8097);
and U11660 (N_11660,N_9371,N_5767);
or U11661 (N_11661,N_9011,N_6420);
nor U11662 (N_11662,N_7864,N_6844);
nand U11663 (N_11663,N_7295,N_7430);
and U11664 (N_11664,N_5970,N_5027);
or U11665 (N_11665,N_7214,N_5886);
nor U11666 (N_11666,N_5014,N_9060);
and U11667 (N_11667,N_7175,N_6956);
xor U11668 (N_11668,N_9283,N_8686);
xnor U11669 (N_11669,N_7178,N_5859);
xor U11670 (N_11670,N_9622,N_9180);
xor U11671 (N_11671,N_6876,N_8924);
nor U11672 (N_11672,N_5463,N_7492);
xnor U11673 (N_11673,N_6001,N_5050);
and U11674 (N_11674,N_7925,N_6569);
and U11675 (N_11675,N_8843,N_5298);
and U11676 (N_11676,N_8059,N_6672);
xor U11677 (N_11677,N_5727,N_5016);
and U11678 (N_11678,N_6833,N_7898);
nand U11679 (N_11679,N_7614,N_8571);
nand U11680 (N_11680,N_7876,N_7852);
nand U11681 (N_11681,N_5225,N_6975);
nand U11682 (N_11682,N_9959,N_5269);
or U11683 (N_11683,N_9517,N_7203);
xor U11684 (N_11684,N_6755,N_5323);
and U11685 (N_11685,N_6462,N_9362);
and U11686 (N_11686,N_9075,N_7042);
nor U11687 (N_11687,N_6768,N_6143);
nand U11688 (N_11688,N_9124,N_5536);
xor U11689 (N_11689,N_8755,N_6766);
and U11690 (N_11690,N_6634,N_6094);
nor U11691 (N_11691,N_5296,N_8314);
nor U11692 (N_11692,N_8001,N_7895);
and U11693 (N_11693,N_9837,N_9849);
nor U11694 (N_11694,N_6976,N_6015);
and U11695 (N_11695,N_6761,N_9019);
or U11696 (N_11696,N_6636,N_5438);
and U11697 (N_11697,N_6896,N_7334);
nand U11698 (N_11698,N_7001,N_5439);
nand U11699 (N_11699,N_5868,N_7943);
and U11700 (N_11700,N_8445,N_5944);
and U11701 (N_11701,N_9104,N_8083);
xnor U11702 (N_11702,N_7759,N_5338);
xnor U11703 (N_11703,N_7263,N_6861);
xor U11704 (N_11704,N_5011,N_9794);
or U11705 (N_11705,N_5466,N_8124);
and U11706 (N_11706,N_9613,N_6008);
xor U11707 (N_11707,N_9306,N_8725);
and U11708 (N_11708,N_5468,N_9418);
or U11709 (N_11709,N_7344,N_8991);
and U11710 (N_11710,N_5067,N_5778);
nor U11711 (N_11711,N_8473,N_7988);
nor U11712 (N_11712,N_7264,N_8875);
nor U11713 (N_11713,N_6079,N_7724);
xnor U11714 (N_11714,N_9008,N_7933);
nand U11715 (N_11715,N_5752,N_7880);
xnor U11716 (N_11716,N_5756,N_5351);
xor U11717 (N_11717,N_7550,N_9020);
xor U11718 (N_11718,N_9160,N_5840);
or U11719 (N_11719,N_6704,N_8041);
nand U11720 (N_11720,N_9854,N_7438);
nor U11721 (N_11721,N_5883,N_9210);
and U11722 (N_11722,N_8818,N_8573);
xnor U11723 (N_11723,N_5726,N_6689);
nor U11724 (N_11724,N_6752,N_8208);
or U11725 (N_11725,N_7235,N_6384);
nand U11726 (N_11726,N_7515,N_7535);
nor U11727 (N_11727,N_9056,N_5087);
or U11728 (N_11728,N_8152,N_7269);
nor U11729 (N_11729,N_6255,N_7779);
nand U11730 (N_11730,N_6728,N_7039);
and U11731 (N_11731,N_7805,N_8876);
or U11732 (N_11732,N_6942,N_6201);
xor U11733 (N_11733,N_6962,N_8077);
nor U11734 (N_11734,N_5698,N_8468);
nand U11735 (N_11735,N_5586,N_7085);
and U11736 (N_11736,N_9012,N_9705);
or U11737 (N_11737,N_6122,N_8737);
nand U11738 (N_11738,N_6236,N_6208);
or U11739 (N_11739,N_6364,N_8508);
nand U11740 (N_11740,N_9587,N_9880);
nor U11741 (N_11741,N_7494,N_8069);
nor U11742 (N_11742,N_8898,N_6930);
nor U11743 (N_11743,N_6199,N_6803);
nand U11744 (N_11744,N_7122,N_6085);
or U11745 (N_11745,N_8829,N_7638);
and U11746 (N_11746,N_9689,N_7231);
or U11747 (N_11747,N_8759,N_5831);
or U11748 (N_11748,N_6069,N_5913);
nand U11749 (N_11749,N_8787,N_8821);
and U11750 (N_11750,N_5648,N_6438);
nor U11751 (N_11751,N_9862,N_9763);
or U11752 (N_11752,N_6630,N_7715);
or U11753 (N_11753,N_8793,N_7043);
xnor U11754 (N_11754,N_9112,N_9214);
nand U11755 (N_11755,N_6576,N_7286);
nand U11756 (N_11756,N_8869,N_8670);
nand U11757 (N_11757,N_9428,N_9435);
nor U11758 (N_11758,N_9147,N_8233);
or U11759 (N_11759,N_6409,N_6467);
and U11760 (N_11760,N_6461,N_7059);
and U11761 (N_11761,N_5006,N_6664);
nand U11762 (N_11762,N_8591,N_8126);
and U11763 (N_11763,N_5152,N_6277);
and U11764 (N_11764,N_6335,N_9322);
and U11765 (N_11765,N_9879,N_8142);
or U11766 (N_11766,N_8474,N_8570);
nand U11767 (N_11767,N_7002,N_9597);
nor U11768 (N_11768,N_8601,N_9090);
and U11769 (N_11769,N_7797,N_8317);
xor U11770 (N_11770,N_5181,N_5862);
nor U11771 (N_11771,N_5909,N_9539);
or U11772 (N_11772,N_6695,N_6564);
and U11773 (N_11773,N_5704,N_7141);
xnor U11774 (N_11774,N_9299,N_5099);
xnor U11775 (N_11775,N_8222,N_8633);
xor U11776 (N_11776,N_9126,N_8683);
nor U11777 (N_11777,N_8533,N_5576);
and U11778 (N_11778,N_7288,N_5923);
and U11779 (N_11779,N_8062,N_6197);
nand U11780 (N_11780,N_5545,N_7240);
xor U11781 (N_11781,N_7922,N_7119);
nor U11782 (N_11782,N_5368,N_8865);
or U11783 (N_11783,N_8177,N_8240);
nand U11784 (N_11784,N_8326,N_5381);
nor U11785 (N_11785,N_8084,N_6019);
nand U11786 (N_11786,N_8790,N_9196);
nor U11787 (N_11787,N_5407,N_9170);
xor U11788 (N_11788,N_6142,N_8188);
or U11789 (N_11789,N_6916,N_6213);
and U11790 (N_11790,N_6099,N_6413);
nor U11791 (N_11791,N_7061,N_7400);
or U11792 (N_11792,N_6843,N_8702);
nor U11793 (N_11793,N_9247,N_7861);
and U11794 (N_11794,N_8414,N_6949);
and U11795 (N_11795,N_8760,N_9444);
or U11796 (N_11796,N_9158,N_5687);
nand U11797 (N_11797,N_8443,N_8798);
and U11798 (N_11798,N_7951,N_6268);
and U11799 (N_11799,N_6775,N_6084);
nor U11800 (N_11800,N_8144,N_5454);
nor U11801 (N_11801,N_6107,N_7046);
and U11802 (N_11802,N_8213,N_9675);
xnor U11803 (N_11803,N_5446,N_6468);
nor U11804 (N_11804,N_8503,N_5879);
nor U11805 (N_11805,N_5198,N_5528);
and U11806 (N_11806,N_8614,N_7346);
nor U11807 (N_11807,N_6680,N_7930);
xnor U11808 (N_11808,N_8595,N_8447);
or U11809 (N_11809,N_7855,N_5914);
or U11810 (N_11810,N_9903,N_9599);
xnor U11811 (N_11811,N_5618,N_5045);
or U11812 (N_11812,N_6146,N_5569);
xor U11813 (N_11813,N_9934,N_7990);
and U11814 (N_11814,N_6882,N_7708);
xor U11815 (N_11815,N_5733,N_9351);
and U11816 (N_11816,N_5100,N_5185);
xnor U11817 (N_11817,N_6062,N_9360);
xnor U11818 (N_11818,N_6323,N_6232);
nand U11819 (N_11819,N_9927,N_9222);
nand U11820 (N_11820,N_7811,N_5786);
nand U11821 (N_11821,N_8962,N_5285);
xnor U11822 (N_11822,N_5957,N_9789);
nor U11823 (N_11823,N_6405,N_6496);
nor U11824 (N_11824,N_5065,N_9330);
nand U11825 (N_11825,N_5743,N_6131);
nand U11826 (N_11826,N_5386,N_5961);
nor U11827 (N_11827,N_7359,N_6992);
xnor U11828 (N_11828,N_9391,N_7080);
xnor U11829 (N_11829,N_5993,N_6280);
and U11830 (N_11830,N_7653,N_5770);
and U11831 (N_11831,N_6626,N_5759);
xor U11832 (N_11832,N_9921,N_6783);
nor U11833 (N_11833,N_7162,N_5510);
and U11834 (N_11834,N_6772,N_6338);
nor U11835 (N_11835,N_7273,N_7006);
and U11836 (N_11836,N_7018,N_6931);
and U11837 (N_11837,N_5361,N_6088);
nand U11838 (N_11838,N_9293,N_6794);
or U11839 (N_11839,N_6163,N_7176);
and U11840 (N_11840,N_6548,N_9588);
or U11841 (N_11841,N_8442,N_9955);
and U11842 (N_11842,N_7918,N_7221);
or U11843 (N_11843,N_9820,N_8779);
nand U11844 (N_11844,N_6835,N_6922);
nor U11845 (N_11845,N_8743,N_5884);
xnor U11846 (N_11846,N_6820,N_8332);
nor U11847 (N_11847,N_6713,N_9719);
nand U11848 (N_11848,N_6378,N_6336);
nor U11849 (N_11849,N_6028,N_8699);
xnor U11850 (N_11850,N_5492,N_7311);
nand U11851 (N_11851,N_8236,N_5617);
nand U11852 (N_11852,N_9478,N_9249);
and U11853 (N_11853,N_8892,N_6551);
and U11854 (N_11854,N_9844,N_7720);
or U11855 (N_11855,N_5043,N_5721);
nor U11856 (N_11856,N_8946,N_9440);
xor U11857 (N_11857,N_5484,N_6386);
nor U11858 (N_11858,N_6959,N_9822);
nor U11859 (N_11859,N_5817,N_8567);
xnor U11860 (N_11860,N_8810,N_5461);
xnor U11861 (N_11861,N_6181,N_5163);
nor U11862 (N_11862,N_8744,N_9787);
or U11863 (N_11863,N_5623,N_7754);
nor U11864 (N_11864,N_8696,N_6358);
nor U11865 (N_11865,N_6701,N_6272);
or U11866 (N_11866,N_9397,N_6961);
nor U11867 (N_11867,N_8872,N_9003);
nand U11868 (N_11868,N_8105,N_9027);
nor U11869 (N_11869,N_5389,N_6032);
nor U11870 (N_11870,N_5129,N_7935);
xor U11871 (N_11871,N_5588,N_6421);
or U11872 (N_11872,N_7350,N_9711);
xnor U11873 (N_11873,N_7645,N_5112);
nor U11874 (N_11874,N_5220,N_6374);
nand U11875 (N_11875,N_6632,N_6699);
nor U11876 (N_11876,N_8011,N_9448);
xnor U11877 (N_11877,N_9055,N_5125);
nand U11878 (N_11878,N_5085,N_7142);
or U11879 (N_11879,N_7184,N_9116);
xnor U11880 (N_11880,N_6415,N_5527);
and U11881 (N_11881,N_8225,N_5564);
and U11882 (N_11882,N_8008,N_6583);
and U11883 (N_11883,N_9297,N_8327);
nand U11884 (N_11884,N_5827,N_7310);
xnor U11885 (N_11885,N_8055,N_8752);
nand U11886 (N_11886,N_7685,N_5525);
xor U11887 (N_11887,N_6497,N_8260);
and U11888 (N_11888,N_7850,N_9826);
nor U11889 (N_11889,N_6254,N_8214);
nor U11890 (N_11890,N_9393,N_7527);
or U11891 (N_11891,N_7650,N_6782);
or U11892 (N_11892,N_7233,N_7274);
nor U11893 (N_11893,N_8076,N_5901);
or U11894 (N_11894,N_9477,N_8607);
xnor U11895 (N_11895,N_9975,N_6372);
or U11896 (N_11896,N_6356,N_6683);
nand U11897 (N_11897,N_8496,N_8871);
or U11898 (N_11898,N_9596,N_7677);
nor U11899 (N_11899,N_8854,N_7765);
nor U11900 (N_11900,N_6545,N_7863);
nand U11901 (N_11901,N_6180,N_6662);
nor U11902 (N_11902,N_7559,N_5910);
and U11903 (N_11903,N_6110,N_6754);
xnor U11904 (N_11904,N_6296,N_9670);
and U11905 (N_11905,N_6821,N_8070);
xor U11906 (N_11906,N_7868,N_7410);
nand U11907 (N_11907,N_6173,N_8676);
and U11908 (N_11908,N_5723,N_9108);
and U11909 (N_11909,N_6996,N_8599);
nand U11910 (N_11910,N_7124,N_7034);
nor U11911 (N_11911,N_7809,N_9632);
xor U11912 (N_11912,N_9627,N_7464);
and U11913 (N_11913,N_5397,N_6577);
nand U11914 (N_11914,N_6598,N_8561);
nand U11915 (N_11915,N_6919,N_8551);
nor U11916 (N_11916,N_8979,N_8723);
and U11917 (N_11917,N_9501,N_6971);
nor U11918 (N_11918,N_6211,N_7404);
and U11919 (N_11919,N_6353,N_9764);
nor U11920 (N_11920,N_5928,N_7641);
or U11921 (N_11921,N_6741,N_8127);
or U11922 (N_11922,N_9262,N_6840);
nor U11923 (N_11923,N_9455,N_7904);
nor U11924 (N_11924,N_8361,N_6390);
nor U11925 (N_11925,N_6449,N_6078);
nand U11926 (N_11926,N_5546,N_7246);
and U11927 (N_11927,N_6530,N_8511);
nor U11928 (N_11928,N_8287,N_9982);
or U11929 (N_11929,N_8254,N_9349);
or U11930 (N_11930,N_8937,N_9217);
xnor U11931 (N_11931,N_6929,N_6348);
nand U11932 (N_11932,N_7323,N_5121);
and U11933 (N_11933,N_5881,N_6623);
nand U11934 (N_11934,N_5333,N_7370);
nor U11935 (N_11935,N_5761,N_7244);
xnor U11936 (N_11936,N_7636,N_5577);
nor U11937 (N_11937,N_8984,N_5738);
xnor U11938 (N_11938,N_8692,N_6932);
and U11939 (N_11939,N_9707,N_9179);
or U11940 (N_11940,N_9895,N_6837);
nor U11941 (N_11941,N_7163,N_8734);
and U11942 (N_11942,N_9702,N_8094);
and U11943 (N_11943,N_5919,N_9426);
and U11944 (N_11944,N_9432,N_5980);
nor U11945 (N_11945,N_5304,N_5009);
nor U11946 (N_11946,N_5550,N_8108);
nor U11947 (N_11947,N_7267,N_5975);
and U11948 (N_11948,N_7014,N_7416);
and U11949 (N_11949,N_9947,N_6328);
and U11950 (N_11950,N_7362,N_9058);
or U11951 (N_11951,N_8581,N_7433);
or U11952 (N_11952,N_6425,N_8786);
nor U11953 (N_11953,N_8502,N_7054);
and U11954 (N_11954,N_6210,N_7366);
and U11955 (N_11955,N_9067,N_9569);
and U11956 (N_11956,N_7595,N_5224);
xor U11957 (N_11957,N_5544,N_9550);
or U11958 (N_11958,N_6923,N_6324);
or U11959 (N_11959,N_5098,N_9048);
nand U11960 (N_11960,N_6188,N_5409);
and U11961 (N_11961,N_5324,N_6176);
nand U11962 (N_11962,N_8928,N_8347);
nor U11963 (N_11963,N_6756,N_6237);
nor U11964 (N_11964,N_6519,N_8735);
and U11965 (N_11965,N_5711,N_7622);
nand U11966 (N_11966,N_7647,N_7547);
and U11967 (N_11967,N_8811,N_6304);
xnor U11968 (N_11968,N_7457,N_7232);
xnor U11969 (N_11969,N_5663,N_9828);
nor U11970 (N_11970,N_6776,N_9233);
and U11971 (N_11971,N_9611,N_6686);
or U11972 (N_11972,N_9962,N_5447);
xnor U11973 (N_11973,N_9245,N_5635);
or U11974 (N_11974,N_6016,N_8506);
and U11975 (N_11975,N_5935,N_5018);
nand U11976 (N_11976,N_6283,N_9476);
or U11977 (N_11977,N_5771,N_5524);
and U11978 (N_11978,N_6554,N_8553);
nor U11979 (N_11979,N_8401,N_8134);
nand U11980 (N_11980,N_6723,N_5188);
xnor U11981 (N_11981,N_5785,N_6491);
or U11982 (N_11982,N_6147,N_8881);
and U11983 (N_11983,N_9044,N_6399);
nand U11984 (N_11984,N_8556,N_8460);
nand U11985 (N_11985,N_9634,N_9073);
nor U11986 (N_11986,N_8185,N_8489);
nor U11987 (N_11987,N_7675,N_9595);
nand U11988 (N_11988,N_5248,N_7851);
and U11989 (N_11989,N_5578,N_8141);
or U11990 (N_11990,N_6081,N_7396);
xor U11991 (N_11991,N_8073,N_5128);
or U11992 (N_11992,N_5620,N_9402);
nand U11993 (N_11993,N_7266,N_7522);
and U11994 (N_11994,N_8450,N_7265);
xnor U11995 (N_11995,N_5223,N_6029);
nand U11996 (N_11996,N_9240,N_5608);
nor U11997 (N_11997,N_8078,N_8963);
xor U11998 (N_11998,N_9788,N_5748);
nand U11999 (N_11999,N_6943,N_5835);
or U12000 (N_12000,N_7968,N_7339);
and U12001 (N_12001,N_5514,N_6313);
and U12002 (N_12002,N_8410,N_8642);
xor U12003 (N_12003,N_5405,N_5787);
or U12004 (N_12004,N_8115,N_7298);
and U12005 (N_12005,N_6310,N_9065);
and U12006 (N_12006,N_6895,N_8662);
nor U12007 (N_12007,N_6489,N_7086);
or U12008 (N_12008,N_8341,N_6431);
or U12009 (N_12009,N_9047,N_9969);
and U12010 (N_12010,N_9202,N_6964);
nand U12011 (N_12011,N_5581,N_5308);
xor U12012 (N_12012,N_6257,N_8882);
nor U12013 (N_12013,N_7077,N_8364);
xor U12014 (N_12014,N_6042,N_5414);
nand U12015 (N_12015,N_9749,N_7787);
or U12016 (N_12016,N_6747,N_8191);
and U12017 (N_12017,N_9211,N_8369);
nor U12018 (N_12018,N_7633,N_5765);
and U12019 (N_12019,N_8018,N_9797);
nand U12020 (N_12020,N_6947,N_5985);
or U12021 (N_12021,N_8921,N_5093);
nand U12022 (N_12022,N_7964,N_5384);
nand U12023 (N_12023,N_6688,N_9066);
nor U12024 (N_12024,N_6640,N_6366);
nand U12025 (N_12025,N_6593,N_9855);
or U12026 (N_12026,N_9357,N_6218);
nor U12027 (N_12027,N_7959,N_7928);
nor U12028 (N_12028,N_6226,N_5010);
xor U12029 (N_12029,N_9303,N_9582);
or U12030 (N_12030,N_6867,N_5342);
nor U12031 (N_12031,N_7254,N_7780);
and U12032 (N_12032,N_7827,N_6946);
and U12033 (N_12033,N_5764,N_7196);
nor U12034 (N_12034,N_8645,N_9830);
nand U12035 (N_12035,N_8005,N_5843);
xnor U12036 (N_12036,N_8900,N_5512);
nand U12037 (N_12037,N_5676,N_8620);
nor U12038 (N_12038,N_7965,N_9017);
and U12039 (N_12039,N_5762,N_8295);
nand U12040 (N_12040,N_8088,N_6027);
nor U12041 (N_12041,N_5808,N_9916);
or U12042 (N_12042,N_9030,N_9325);
nor U12043 (N_12043,N_7289,N_7730);
or U12044 (N_12044,N_5486,N_8920);
xor U12045 (N_12045,N_9818,N_5505);
xor U12046 (N_12046,N_9092,N_5162);
nor U12047 (N_12047,N_8653,N_7227);
or U12048 (N_12048,N_6682,N_8742);
xor U12049 (N_12049,N_9149,N_8374);
and U12050 (N_12050,N_6136,N_6503);
nand U12051 (N_12051,N_7301,N_8766);
xnor U12052 (N_12052,N_5462,N_5646);
and U12053 (N_12053,N_9292,N_7010);
and U12054 (N_12054,N_6278,N_7185);
and U12055 (N_12055,N_9523,N_8476);
nand U12056 (N_12056,N_7052,N_9845);
nor U12057 (N_12057,N_7427,N_9714);
xnor U12058 (N_12058,N_5542,N_8618);
and U12059 (N_12059,N_7202,N_7027);
nand U12060 (N_12060,N_8098,N_8925);
xor U12061 (N_12061,N_6212,N_8697);
or U12062 (N_12062,N_6573,N_8017);
nor U12063 (N_12063,N_7171,N_9278);
and U12064 (N_12064,N_6373,N_8004);
or U12065 (N_12065,N_7159,N_5234);
nor U12066 (N_12066,N_9538,N_5950);
xor U12067 (N_12067,N_9888,N_8334);
nor U12068 (N_12068,N_8586,N_8608);
nor U12069 (N_12069,N_9655,N_9795);
or U12070 (N_12070,N_6967,N_5227);
and U12071 (N_12071,N_7546,N_6270);
nor U12072 (N_12072,N_6435,N_9276);
and U12073 (N_12073,N_7425,N_7357);
nand U12074 (N_12074,N_7816,N_9836);
and U12075 (N_12075,N_7193,N_7575);
xor U12076 (N_12076,N_8933,N_5374);
xnor U12077 (N_12077,N_6036,N_7021);
xnor U12078 (N_12078,N_5591,N_7186);
nor U12079 (N_12079,N_6904,N_5568);
xnor U12080 (N_12080,N_6017,N_5497);
or U12081 (N_12081,N_6586,N_8895);
nand U12082 (N_12082,N_7818,N_5538);
nor U12083 (N_12083,N_7665,N_8340);
nor U12084 (N_12084,N_7296,N_6654);
or U12085 (N_12085,N_9329,N_7407);
nor U12086 (N_12086,N_6332,N_7882);
xor U12087 (N_12087,N_9953,N_8761);
nand U12088 (N_12088,N_5816,N_6827);
or U12089 (N_12089,N_8085,N_9750);
or U12090 (N_12090,N_8543,N_5905);
and U12091 (N_12091,N_7950,N_6494);
xnor U12092 (N_12092,N_8626,N_7910);
or U12093 (N_12093,N_8248,N_9290);
nand U12094 (N_12094,N_7997,N_9040);
nor U12095 (N_12095,N_6202,N_7652);
or U12096 (N_12096,N_5473,N_7906);
nor U12097 (N_12097,N_5058,N_8306);
and U12098 (N_12098,N_6217,N_9070);
xor U12099 (N_12099,N_7767,N_5256);
or U12100 (N_12100,N_7568,N_8961);
or U12101 (N_12101,N_6452,N_7914);
xnor U12102 (N_12102,N_8968,N_7531);
xnor U12103 (N_12103,N_7976,N_5889);
or U12104 (N_12104,N_8964,N_8594);
nand U12105 (N_12105,N_7506,N_9084);
and U12106 (N_12106,N_9726,N_7475);
or U12107 (N_12107,N_5932,N_7585);
nand U12108 (N_12108,N_9778,N_5737);
xor U12109 (N_12109,N_9157,N_7738);
nor U12110 (N_12110,N_6849,N_9215);
nand U12111 (N_12111,N_5209,N_7307);
nor U12112 (N_12112,N_8580,N_7686);
xor U12113 (N_12113,N_5882,N_9080);
xor U12114 (N_12114,N_6769,N_8731);
nor U12115 (N_12115,N_6753,N_8826);
nor U12116 (N_12116,N_9767,N_9257);
nor U12117 (N_12117,N_9368,N_9377);
or U12118 (N_12118,N_7978,N_9077);
and U12119 (N_12119,N_5303,N_7909);
and U12120 (N_12120,N_9509,N_7683);
xnor U12121 (N_12121,N_8193,N_9510);
nand U12122 (N_12122,N_9535,N_8168);
and U12123 (N_12123,N_9520,N_7671);
nand U12124 (N_12124,N_8129,N_9584);
nand U12125 (N_12125,N_6830,N_8239);
or U12126 (N_12126,N_8322,N_7113);
nor U12127 (N_12127,N_9546,N_9601);
or U12128 (N_12128,N_8886,N_8201);
nand U12129 (N_12129,N_6920,N_8074);
nand U12130 (N_12130,N_8691,N_9687);
and U12131 (N_12131,N_6357,N_6436);
or U12132 (N_12132,N_9913,N_5429);
or U12133 (N_12133,N_8922,N_8763);
and U12134 (N_12134,N_8446,N_5934);
nor U12135 (N_12135,N_6010,N_7594);
and U12136 (N_12136,N_9936,N_8135);
nand U12137 (N_12137,N_7619,N_6249);
xor U12138 (N_12138,N_5824,N_8277);
xor U12139 (N_12139,N_7456,N_9029);
or U12140 (N_12140,N_8344,N_9792);
xnor U12141 (N_12141,N_8259,N_7477);
xor U12142 (N_12142,N_6418,N_5989);
and U12143 (N_12143,N_7893,N_7719);
xnor U12144 (N_12144,N_5403,N_9840);
and U12145 (N_12145,N_8842,N_9452);
and U12146 (N_12146,N_8848,N_5792);
xnor U12147 (N_12147,N_5192,N_7251);
xnor U12148 (N_12148,N_5732,N_9258);
xnor U12149 (N_12149,N_6737,N_6711);
nor U12150 (N_12150,N_5038,N_6883);
nand U12151 (N_12151,N_8382,N_9219);
xor U12152 (N_12152,N_5951,N_7489);
nor U12153 (N_12153,N_5678,N_9088);
and U12154 (N_12154,N_6291,N_7268);
and U12155 (N_12155,N_9629,N_6130);
or U12156 (N_12156,N_7835,N_9086);
xor U12157 (N_12157,N_9745,N_5358);
xnor U12158 (N_12158,N_9971,N_8659);
nor U12159 (N_12159,N_8325,N_8205);
xor U12160 (N_12160,N_8792,N_6796);
nand U12161 (N_12161,N_5811,N_5430);
nand U12162 (N_12162,N_8820,N_8352);
xnor U12163 (N_12163,N_8624,N_8485);
and U12164 (N_12164,N_9694,N_8133);
nor U12165 (N_12165,N_9577,N_7824);
nor U12166 (N_12166,N_9716,N_8808);
and U12167 (N_12167,N_6115,N_5624);
nor U12168 (N_12168,N_9177,N_8748);
xor U12169 (N_12169,N_7177,N_5751);
nor U12170 (N_12170,N_7752,N_9680);
and U12171 (N_12171,N_8740,N_6981);
nand U12172 (N_12172,N_9793,N_5741);
and U12173 (N_12173,N_6924,N_5812);
and U12174 (N_12174,N_5736,N_5260);
nor U12175 (N_12175,N_7327,N_9676);
and U12176 (N_12176,N_8710,N_7019);
nor U12177 (N_12177,N_5364,N_5091);
xnor U12178 (N_12178,N_8590,N_5969);
or U12179 (N_12179,N_6192,N_7996);
xor U12180 (N_12180,N_8977,N_8367);
nor U12181 (N_12181,N_5472,N_9643);
nor U12182 (N_12182,N_8038,N_5677);
and U12183 (N_12183,N_6938,N_7768);
or U12184 (N_12184,N_8804,N_6184);
nor U12185 (N_12185,N_9064,N_9304);
or U12186 (N_12186,N_6487,N_8941);
nand U12187 (N_12187,N_9776,N_9846);
nor U12188 (N_12188,N_9721,N_6952);
nand U12189 (N_12189,N_8775,N_5416);
or U12190 (N_12190,N_7941,N_6899);
or U12191 (N_12191,N_6204,N_6439);
xnor U12192 (N_12192,N_6177,N_6871);
or U12193 (N_12193,N_9823,N_8125);
or U12194 (N_12194,N_9281,N_9524);
nand U12195 (N_12195,N_7512,N_5089);
nand U12196 (N_12196,N_8387,N_9859);
nor U12197 (N_12197,N_6823,N_7901);
and U12198 (N_12198,N_6927,N_7380);
nand U12199 (N_12199,N_7749,N_7403);
xnor U12200 (N_12200,N_8840,N_8940);
xor U12201 (N_12201,N_6918,N_8776);
nand U12202 (N_12202,N_9190,N_5159);
or U12203 (N_12203,N_5032,N_9279);
or U12204 (N_12204,N_8530,N_6555);
nor U12205 (N_12205,N_5150,N_5023);
and U12206 (N_12206,N_8656,N_8203);
and U12207 (N_12207,N_9949,N_9261);
nor U12208 (N_12208,N_5872,N_9666);
xor U12209 (N_12209,N_8409,N_6002);
or U12210 (N_12210,N_6644,N_8674);
nand U12211 (N_12211,N_6095,N_5326);
and U12212 (N_12212,N_6856,N_6490);
nor U12213 (N_12213,N_9914,N_6785);
nor U12214 (N_12214,N_7632,N_5513);
or U12215 (N_12215,N_9625,N_9332);
nor U12216 (N_12216,N_5964,N_7735);
xnor U12217 (N_12217,N_5661,N_9254);
nor U12218 (N_12218,N_5626,N_8007);
and U12219 (N_12219,N_5355,N_6572);
xor U12220 (N_12220,N_7212,N_5930);
nand U12221 (N_12221,N_8765,N_7725);
xor U12222 (N_12222,N_8424,N_6808);
and U12223 (N_12223,N_6552,N_6863);
nor U12224 (N_12224,N_6477,N_7373);
and U12225 (N_12225,N_7188,N_6797);
or U12226 (N_12226,N_5896,N_7902);
nor U12227 (N_12227,N_5644,N_8227);
xor U12228 (N_12228,N_8857,N_5622);
nor U12229 (N_12229,N_8110,N_7326);
xnor U12230 (N_12230,N_5873,N_7750);
or U12231 (N_12231,N_6149,N_7552);
nand U12232 (N_12232,N_7028,N_7760);
and U12233 (N_12233,N_5120,N_9841);
xor U12234 (N_12234,N_5287,N_5460);
nor U12235 (N_12235,N_5855,N_6819);
or U12236 (N_12236,N_5673,N_6375);
nor U12237 (N_12237,N_6647,N_7229);
or U12238 (N_12238,N_8716,N_6361);
xnor U12239 (N_12239,N_6705,N_9876);
nor U12240 (N_12240,N_5096,N_8075);
or U12241 (N_12241,N_7245,N_7237);
or U12242 (N_12242,N_8371,N_7881);
nand U12243 (N_12243,N_7394,N_9433);
or U12244 (N_12244,N_6239,N_6857);
and U12245 (N_12245,N_6936,N_9762);
or U12246 (N_12246,N_7969,N_6345);
nor U12247 (N_12247,N_7673,N_9628);
xnor U12248 (N_12248,N_5689,N_8145);
and U12249 (N_12249,N_7174,N_6700);
xnor U12250 (N_12250,N_8262,N_8769);
nor U12251 (N_12251,N_6574,N_8455);
nor U12252 (N_12252,N_7681,N_9919);
nand U12253 (N_12253,N_5363,N_5821);
nand U12254 (N_12254,N_5464,N_6067);
and U12255 (N_12255,N_8785,N_5846);
and U12256 (N_12256,N_9683,N_7012);
or U12257 (N_12257,N_5652,N_9554);
nand U12258 (N_12258,N_8712,N_5083);
nand U12259 (N_12259,N_9094,N_8268);
or U12260 (N_12260,N_6072,N_7309);
and U12261 (N_12261,N_9686,N_9521);
xor U12262 (N_12262,N_7143,N_7306);
or U12263 (N_12263,N_8297,N_5692);
and U12264 (N_12264,N_6041,N_7399);
or U12265 (N_12265,N_6344,N_6607);
nor U12266 (N_12266,N_8764,N_6553);
and U12267 (N_12267,N_7255,N_5202);
nor U12268 (N_12268,N_7383,N_8524);
xnor U12269 (N_12269,N_5283,N_5077);
and U12270 (N_12270,N_9536,N_6595);
nand U12271 (N_12271,N_5653,N_9138);
or U12272 (N_12272,N_9938,N_5169);
and U12273 (N_12273,N_7123,N_6474);
xnor U12274 (N_12274,N_9866,N_7991);
xnor U12275 (N_12275,N_8204,N_7259);
and U12276 (N_12276,N_6944,N_9419);
xnor U12277 (N_12277,N_9808,N_5776);
nor U12278 (N_12278,N_6853,N_5442);
xnor U12279 (N_12279,N_9942,N_6109);
or U12280 (N_12280,N_6588,N_7846);
xnor U12281 (N_12281,N_7436,N_9296);
xnor U12282 (N_12282,N_8138,N_8913);
or U12283 (N_12283,N_5847,N_6065);
and U12284 (N_12284,N_7563,N_7413);
xor U12285 (N_12285,N_8835,N_7454);
or U12286 (N_12286,N_8579,N_8187);
nand U12287 (N_12287,N_8504,N_7243);
and U12288 (N_12288,N_5982,N_5066);
nor U12289 (N_12289,N_8880,N_8853);
xor U12290 (N_12290,N_8467,N_8416);
nand U12291 (N_12291,N_5200,N_5483);
and U12292 (N_12292,N_8745,N_7521);
xnor U12293 (N_12293,N_7814,N_6009);
xnor U12294 (N_12294,N_6790,N_6912);
or U12295 (N_12295,N_7060,N_7763);
xnor U12296 (N_12296,N_9343,N_6406);
or U12297 (N_12297,N_6902,N_6124);
nand U12298 (N_12298,N_5551,N_8212);
and U12299 (N_12299,N_9678,N_6469);
nor U12300 (N_12300,N_6092,N_7278);
nor U12301 (N_12301,N_5413,N_5113);
xnor U12302 (N_12302,N_9937,N_8053);
or U12303 (N_12303,N_9672,N_5633);
xnor U12304 (N_12304,N_6119,N_7992);
or U12305 (N_12305,N_7129,N_9492);
nor U12306 (N_12306,N_6059,N_6014);
xnor U12307 (N_12307,N_7528,N_5994);
xnor U12308 (N_12308,N_7481,N_7503);
nand U12309 (N_12309,N_9024,N_6870);
or U12310 (N_12310,N_5596,N_6432);
xnor U12311 (N_12311,N_5991,N_9966);
nand U12312 (N_12312,N_8061,N_6619);
or U12313 (N_12313,N_9743,N_7625);
or U12314 (N_12314,N_8750,N_7862);
nand U12315 (N_12315,N_8002,N_8140);
or U12316 (N_12316,N_7957,N_5419);
xor U12317 (N_12317,N_8978,N_6850);
or U12318 (N_12318,N_9201,N_5996);
and U12319 (N_12319,N_6516,N_8427);
nor U12320 (N_12320,N_6456,N_6295);
and U12321 (N_12321,N_6744,N_8701);
nor U12322 (N_12322,N_7271,N_7847);
nand U12323 (N_12323,N_9575,N_5040);
nor U12324 (N_12324,N_6939,N_7576);
xor U12325 (N_12325,N_9069,N_7510);
xnor U12326 (N_12326,N_7076,N_7134);
nor U12327 (N_12327,N_9968,N_5671);
or U12328 (N_12328,N_7371,N_6864);
xor U12329 (N_12329,N_8149,N_8868);
nor U12330 (N_12330,N_5494,N_5349);
xor U12331 (N_12331,N_8184,N_7109);
nor U12332 (N_12332,N_9083,N_9460);
and U12333 (N_12333,N_7578,N_7733);
nor U12334 (N_12334,N_7736,N_5701);
nand U12335 (N_12335,N_9316,N_5968);
and U12336 (N_12336,N_6547,N_6666);
xor U12337 (N_12337,N_7230,N_9321);
nand U12338 (N_12338,N_9780,N_9102);
xor U12339 (N_12339,N_8223,N_5675);
xnor U12340 (N_12340,N_9623,N_5068);
or U12341 (N_12341,N_5297,N_8613);
and U12342 (N_12342,N_7743,N_5404);
xor U12343 (N_12343,N_7446,N_6656);
or U12344 (N_12344,N_8709,N_6527);
nand U12345 (N_12345,N_8169,N_5237);
nor U12346 (N_12346,N_8103,N_8598);
nor U12347 (N_12347,N_5858,N_6401);
xnor U12348 (N_12348,N_9496,N_9161);
xor U12349 (N_12349,N_9465,N_8272);
nand U12350 (N_12350,N_7164,N_6005);
nor U12351 (N_12351,N_6071,N_6209);
nand U12352 (N_12352,N_5365,N_7439);
nand U12353 (N_12353,N_8878,N_6811);
nor U12354 (N_12354,N_7892,N_7302);
xor U12355 (N_12355,N_5601,N_9225);
nand U12356 (N_12356,N_6732,N_7954);
nand U12357 (N_12357,N_9484,N_6292);
and U12358 (N_12358,N_6098,N_5890);
and U12359 (N_12359,N_8307,N_9165);
nor U12360 (N_12360,N_9637,N_6312);
nor U12361 (N_12361,N_6765,N_5054);
xnor U12362 (N_12362,N_9339,N_5573);
or U12363 (N_12363,N_8611,N_6346);
or U12364 (N_12364,N_9082,N_5417);
xor U12365 (N_12365,N_7545,N_5477);
nand U12366 (N_12366,N_9256,N_8346);
nor U12367 (N_12367,N_9654,N_5852);
nor U12368 (N_12368,N_6995,N_6684);
or U12369 (N_12369,N_8939,N_6543);
nor U12370 (N_12370,N_5803,N_6248);
nor U12371 (N_12371,N_6423,N_8568);
nand U12372 (N_12372,N_8491,N_9527);
nand U12373 (N_12373,N_6707,N_7865);
nand U12374 (N_12374,N_7985,N_6950);
or U12375 (N_12375,N_5685,N_8479);
or U12376 (N_12376,N_6609,N_5974);
nor U12377 (N_12377,N_8904,N_8647);
or U12378 (N_12378,N_5790,N_5017);
or U12379 (N_12379,N_8102,N_5160);
and U12380 (N_12380,N_5508,N_6786);
or U12381 (N_12381,N_8632,N_8536);
nor U12382 (N_12382,N_8517,N_7840);
xor U12383 (N_12383,N_9385,N_6692);
xnor U12384 (N_12384,N_5316,N_6804);
nor U12385 (N_12385,N_9608,N_8528);
nand U12386 (N_12386,N_9709,N_7117);
and U12387 (N_12387,N_9050,N_7532);
nor U12388 (N_12388,N_8023,N_9220);
nand U12389 (N_12389,N_6601,N_6089);
nor U12390 (N_12390,N_9270,N_9899);
xor U12391 (N_12391,N_6523,N_9302);
and U12392 (N_12392,N_7994,N_9922);
nor U12393 (N_12393,N_8310,N_9472);
xor U12394 (N_12394,N_5800,N_6303);
or U12395 (N_12395,N_7375,N_8677);
and U12396 (N_12396,N_5654,N_5731);
xor U12397 (N_12397,N_9831,N_7125);
xnor U12398 (N_12398,N_6694,N_5587);
xnor U12399 (N_12399,N_8351,N_9392);
nand U12400 (N_12400,N_5354,N_8043);
or U12401 (N_12401,N_9999,N_6643);
nand U12402 (N_12402,N_6153,N_7287);
and U12403 (N_12403,N_8609,N_7849);
or U12404 (N_12404,N_8944,N_6334);
nor U12405 (N_12405,N_5509,N_6235);
and U12406 (N_12406,N_9773,N_8058);
and U12407 (N_12407,N_8974,N_5796);
xnor U12408 (N_12408,N_5870,N_9388);
nor U12409 (N_12409,N_9052,N_7335);
nor U12410 (N_12410,N_6058,N_6760);
and U12411 (N_12411,N_5019,N_7879);
nor U12412 (N_12412,N_5310,N_8514);
xnor U12413 (N_12413,N_9035,N_5984);
and U12414 (N_12414,N_8269,N_8704);
and U12415 (N_12415,N_7669,N_5478);
and U12416 (N_12416,N_5795,N_5143);
and U12417 (N_12417,N_6651,N_7854);
xor U12418 (N_12418,N_6800,N_6376);
xnor U12419 (N_12419,N_5988,N_7067);
or U12420 (N_12420,N_6402,N_9373);
nor U12421 (N_12421,N_5064,N_9751);
xor U12422 (N_12422,N_9361,N_5703);
or U12423 (N_12423,N_7919,N_9809);
xor U12424 (N_12424,N_8238,N_5000);
or U12425 (N_12425,N_7194,N_6298);
or U12426 (N_12426,N_5420,N_6565);
nor U12427 (N_12427,N_5642,N_8897);
nand U12428 (N_12428,N_6620,N_5437);
nor U12429 (N_12429,N_5708,N_8316);
or U12430 (N_12430,N_7723,N_9526);
nand U12431 (N_12431,N_8679,N_6414);
nor U12432 (N_12432,N_9590,N_5534);
nor U12433 (N_12433,N_9631,N_5441);
nor U12434 (N_12434,N_7466,N_5427);
nand U12435 (N_12435,N_9305,N_5938);
xnor U12436 (N_12436,N_6053,N_9488);
xor U12437 (N_12437,N_5537,N_9367);
or U12438 (N_12438,N_8025,N_5271);
nor U12439 (N_12439,N_9515,N_7450);
and U12440 (N_12440,N_5385,N_6221);
nor U12441 (N_12441,N_8718,N_9274);
nor U12442 (N_12442,N_8181,N_5187);
and U12443 (N_12443,N_5147,N_5826);
or U12444 (N_12444,N_6417,N_9471);
xnor U12445 (N_12445,N_7215,N_5686);
nor U12446 (N_12446,N_5393,N_6365);
xnor U12447 (N_12447,N_6186,N_6690);
nor U12448 (N_12448,N_9298,N_6174);
or U12449 (N_12449,N_5552,N_7461);
or U12450 (N_12450,N_9434,N_9760);
nor U12451 (N_12451,N_7613,N_6624);
xnor U12452 (N_12452,N_7727,N_8980);
or U12453 (N_12453,N_7093,N_8229);
nand U12454 (N_12454,N_7000,N_6434);
nor U12455 (N_12455,N_7495,N_6514);
nor U12456 (N_12456,N_9151,N_5973);
or U12457 (N_12457,N_9294,N_9891);
or U12458 (N_12458,N_6791,N_9889);
or U12459 (N_12459,N_7981,N_8864);
xor U12460 (N_12460,N_9364,N_5280);
and U12461 (N_12461,N_9987,N_5396);
xnor U12462 (N_12462,N_7363,N_9868);
or U12463 (N_12463,N_6698,N_7800);
nor U12464 (N_12464,N_9810,N_5474);
and U12465 (N_12465,N_7201,N_6087);
xnor U12466 (N_12466,N_7771,N_9087);
and U12467 (N_12467,N_8411,N_5799);
nor U12468 (N_12468,N_5039,N_6352);
nand U12469 (N_12469,N_6287,N_8741);
or U12470 (N_12470,N_5851,N_7305);
nor U12471 (N_12471,N_9645,N_9175);
xor U12472 (N_12472,N_7722,N_8812);
nor U12473 (N_12473,N_9580,N_9853);
nor U12474 (N_12474,N_8393,N_5490);
nand U12475 (N_12475,N_6156,N_5033);
or U12476 (N_12476,N_9732,N_9246);
xor U12477 (N_12477,N_5558,N_7701);
or U12478 (N_12478,N_8983,N_5511);
and U12479 (N_12479,N_8362,N_9552);
xnor U12480 (N_12480,N_7118,N_9042);
or U12481 (N_12481,N_9592,N_5495);
xor U12482 (N_12482,N_9664,N_9983);
or U12483 (N_12483,N_5262,N_5734);
and U12484 (N_12484,N_6351,N_7353);
and U12485 (N_12485,N_9663,N_7742);
xor U12486 (N_12486,N_9420,N_7789);
xor U12487 (N_12487,N_9626,N_6416);
nor U12488 (N_12488,N_5539,N_5850);
or U12489 (N_12489,N_7205,N_5697);
and U12490 (N_12490,N_7756,N_7426);
nand U12491 (N_12491,N_8425,N_6958);
xor U12492 (N_12492,N_9730,N_7420);
nor U12493 (N_12493,N_7916,N_5986);
nor U12494 (N_12494,N_7063,N_5584);
xor U12495 (N_12495,N_8012,N_6125);
xnor U12496 (N_12496,N_5026,N_5109);
nor U12497 (N_12497,N_9193,N_6244);
and U12498 (N_12498,N_7209,N_9668);
xor U12499 (N_12499,N_6440,N_6090);
or U12500 (N_12500,N_9507,N_7937);
or U12501 (N_12501,N_7994,N_9955);
or U12502 (N_12502,N_5074,N_5678);
xnor U12503 (N_12503,N_9017,N_5969);
or U12504 (N_12504,N_6679,N_8629);
nor U12505 (N_12505,N_9382,N_8364);
or U12506 (N_12506,N_5867,N_5279);
and U12507 (N_12507,N_7138,N_5495);
or U12508 (N_12508,N_7327,N_9701);
nand U12509 (N_12509,N_5029,N_6664);
nand U12510 (N_12510,N_7007,N_9262);
xor U12511 (N_12511,N_6647,N_9667);
nand U12512 (N_12512,N_7452,N_6809);
nor U12513 (N_12513,N_5535,N_6945);
xnor U12514 (N_12514,N_8063,N_8026);
xor U12515 (N_12515,N_5685,N_8212);
xnor U12516 (N_12516,N_9735,N_8080);
xor U12517 (N_12517,N_9420,N_6527);
or U12518 (N_12518,N_8876,N_9618);
and U12519 (N_12519,N_5491,N_9892);
or U12520 (N_12520,N_9996,N_8242);
xor U12521 (N_12521,N_8408,N_7854);
nand U12522 (N_12522,N_7499,N_9238);
or U12523 (N_12523,N_8580,N_7137);
nor U12524 (N_12524,N_9494,N_5674);
xnor U12525 (N_12525,N_7820,N_7607);
or U12526 (N_12526,N_9947,N_5066);
and U12527 (N_12527,N_9302,N_7066);
xnor U12528 (N_12528,N_5702,N_8170);
or U12529 (N_12529,N_8542,N_6173);
and U12530 (N_12530,N_8189,N_6882);
or U12531 (N_12531,N_6955,N_6753);
and U12532 (N_12532,N_7306,N_9615);
nand U12533 (N_12533,N_9060,N_6437);
and U12534 (N_12534,N_5039,N_5268);
nor U12535 (N_12535,N_8505,N_9828);
and U12536 (N_12536,N_9609,N_8758);
nand U12537 (N_12537,N_8853,N_7586);
and U12538 (N_12538,N_7198,N_6155);
and U12539 (N_12539,N_5844,N_8944);
and U12540 (N_12540,N_9670,N_8412);
and U12541 (N_12541,N_5218,N_5240);
nor U12542 (N_12542,N_7746,N_5625);
xor U12543 (N_12543,N_8863,N_7547);
or U12544 (N_12544,N_8127,N_6064);
and U12545 (N_12545,N_8140,N_9386);
and U12546 (N_12546,N_8922,N_6557);
xor U12547 (N_12547,N_9237,N_8682);
nor U12548 (N_12548,N_6838,N_5968);
and U12549 (N_12549,N_9169,N_9355);
or U12550 (N_12550,N_8755,N_9345);
nand U12551 (N_12551,N_7939,N_7620);
nand U12552 (N_12552,N_5455,N_8427);
nand U12553 (N_12553,N_9204,N_7466);
xor U12554 (N_12554,N_9460,N_5543);
and U12555 (N_12555,N_7395,N_6085);
nand U12556 (N_12556,N_6358,N_8828);
nor U12557 (N_12557,N_9372,N_9083);
nand U12558 (N_12558,N_8913,N_9173);
or U12559 (N_12559,N_6704,N_9450);
nand U12560 (N_12560,N_7669,N_6415);
xor U12561 (N_12561,N_8308,N_6207);
xor U12562 (N_12562,N_7565,N_6435);
and U12563 (N_12563,N_7800,N_8224);
nand U12564 (N_12564,N_8686,N_6799);
and U12565 (N_12565,N_5335,N_5720);
xor U12566 (N_12566,N_9624,N_7447);
or U12567 (N_12567,N_5804,N_7116);
xnor U12568 (N_12568,N_7800,N_9576);
nand U12569 (N_12569,N_6400,N_9818);
or U12570 (N_12570,N_7586,N_6389);
and U12571 (N_12571,N_8403,N_7114);
nor U12572 (N_12572,N_5818,N_6057);
xor U12573 (N_12573,N_7813,N_5319);
nor U12574 (N_12574,N_5366,N_5986);
or U12575 (N_12575,N_5722,N_9430);
nand U12576 (N_12576,N_6216,N_9959);
and U12577 (N_12577,N_5120,N_9305);
and U12578 (N_12578,N_8555,N_8796);
nor U12579 (N_12579,N_9652,N_8721);
xor U12580 (N_12580,N_8419,N_7551);
xor U12581 (N_12581,N_5833,N_7668);
and U12582 (N_12582,N_8065,N_5782);
nor U12583 (N_12583,N_8029,N_9036);
nor U12584 (N_12584,N_7010,N_5964);
nand U12585 (N_12585,N_9016,N_5486);
xor U12586 (N_12586,N_6045,N_8282);
and U12587 (N_12587,N_8701,N_5812);
and U12588 (N_12588,N_6059,N_6834);
and U12589 (N_12589,N_8410,N_6952);
nor U12590 (N_12590,N_9436,N_7891);
nand U12591 (N_12591,N_7089,N_7544);
nand U12592 (N_12592,N_7935,N_9776);
or U12593 (N_12593,N_7197,N_9903);
or U12594 (N_12594,N_9883,N_7710);
xnor U12595 (N_12595,N_7292,N_6897);
and U12596 (N_12596,N_7100,N_7689);
nand U12597 (N_12597,N_9199,N_7921);
xnor U12598 (N_12598,N_5895,N_5496);
nand U12599 (N_12599,N_9196,N_5343);
nand U12600 (N_12600,N_5893,N_5810);
and U12601 (N_12601,N_8308,N_5568);
or U12602 (N_12602,N_5896,N_6069);
nand U12603 (N_12603,N_9074,N_6166);
xor U12604 (N_12604,N_6243,N_6647);
or U12605 (N_12605,N_7006,N_7621);
xnor U12606 (N_12606,N_7887,N_6902);
and U12607 (N_12607,N_6557,N_9371);
nor U12608 (N_12608,N_8609,N_6456);
nor U12609 (N_12609,N_7662,N_8678);
xnor U12610 (N_12610,N_9728,N_8463);
nand U12611 (N_12611,N_5551,N_9573);
xor U12612 (N_12612,N_6484,N_6763);
nor U12613 (N_12613,N_7683,N_9355);
or U12614 (N_12614,N_5467,N_8169);
nand U12615 (N_12615,N_8226,N_5174);
xnor U12616 (N_12616,N_5609,N_9742);
xnor U12617 (N_12617,N_5332,N_6826);
nand U12618 (N_12618,N_7331,N_8535);
nor U12619 (N_12619,N_5718,N_6911);
nand U12620 (N_12620,N_5495,N_6805);
xnor U12621 (N_12621,N_5746,N_5971);
or U12622 (N_12622,N_9446,N_9696);
and U12623 (N_12623,N_6337,N_9509);
nor U12624 (N_12624,N_5363,N_5101);
and U12625 (N_12625,N_9825,N_6041);
and U12626 (N_12626,N_8989,N_7170);
nor U12627 (N_12627,N_6362,N_7877);
or U12628 (N_12628,N_7529,N_7920);
nor U12629 (N_12629,N_5371,N_9178);
xnor U12630 (N_12630,N_5833,N_9307);
or U12631 (N_12631,N_5369,N_8953);
nor U12632 (N_12632,N_6741,N_7325);
xor U12633 (N_12633,N_5505,N_7419);
and U12634 (N_12634,N_5536,N_9423);
nor U12635 (N_12635,N_6433,N_7301);
or U12636 (N_12636,N_7487,N_6027);
nand U12637 (N_12637,N_7047,N_9200);
xor U12638 (N_12638,N_7423,N_5816);
nand U12639 (N_12639,N_8974,N_9656);
xnor U12640 (N_12640,N_6154,N_7397);
or U12641 (N_12641,N_5192,N_9274);
nor U12642 (N_12642,N_6624,N_9310);
or U12643 (N_12643,N_6338,N_7451);
and U12644 (N_12644,N_8117,N_6650);
and U12645 (N_12645,N_6893,N_7923);
and U12646 (N_12646,N_9699,N_9292);
nor U12647 (N_12647,N_8009,N_7135);
nor U12648 (N_12648,N_9622,N_9939);
or U12649 (N_12649,N_9737,N_8053);
nand U12650 (N_12650,N_8398,N_9032);
nand U12651 (N_12651,N_8920,N_9610);
nor U12652 (N_12652,N_6871,N_6132);
and U12653 (N_12653,N_5258,N_5507);
nand U12654 (N_12654,N_9903,N_8379);
xnor U12655 (N_12655,N_9387,N_8415);
xor U12656 (N_12656,N_5858,N_7960);
and U12657 (N_12657,N_6243,N_6223);
and U12658 (N_12658,N_5724,N_7770);
nand U12659 (N_12659,N_7428,N_7987);
nand U12660 (N_12660,N_9314,N_8668);
xor U12661 (N_12661,N_8795,N_9376);
or U12662 (N_12662,N_7650,N_6139);
and U12663 (N_12663,N_5677,N_7327);
or U12664 (N_12664,N_6781,N_8575);
or U12665 (N_12665,N_8939,N_5148);
or U12666 (N_12666,N_9456,N_9157);
xnor U12667 (N_12667,N_8878,N_9236);
or U12668 (N_12668,N_5221,N_6535);
or U12669 (N_12669,N_5980,N_8499);
and U12670 (N_12670,N_9232,N_5376);
nor U12671 (N_12671,N_9067,N_8836);
nand U12672 (N_12672,N_9727,N_9896);
xnor U12673 (N_12673,N_7946,N_7395);
nor U12674 (N_12674,N_7421,N_9121);
xor U12675 (N_12675,N_8772,N_5610);
nand U12676 (N_12676,N_9417,N_8535);
or U12677 (N_12677,N_8341,N_6949);
nand U12678 (N_12678,N_6309,N_5099);
nor U12679 (N_12679,N_9741,N_9046);
and U12680 (N_12680,N_7344,N_7093);
xnor U12681 (N_12681,N_9478,N_7950);
nor U12682 (N_12682,N_8045,N_7907);
xor U12683 (N_12683,N_5122,N_7506);
nand U12684 (N_12684,N_5372,N_9105);
xor U12685 (N_12685,N_5574,N_8028);
nand U12686 (N_12686,N_7948,N_9250);
nand U12687 (N_12687,N_5089,N_5452);
or U12688 (N_12688,N_6920,N_6820);
nand U12689 (N_12689,N_6400,N_9086);
and U12690 (N_12690,N_6358,N_6307);
or U12691 (N_12691,N_7040,N_9717);
or U12692 (N_12692,N_8967,N_9740);
or U12693 (N_12693,N_7574,N_9486);
and U12694 (N_12694,N_8964,N_7697);
or U12695 (N_12695,N_9226,N_7855);
or U12696 (N_12696,N_5330,N_5563);
and U12697 (N_12697,N_5052,N_6017);
nand U12698 (N_12698,N_8933,N_6900);
xor U12699 (N_12699,N_5025,N_8424);
and U12700 (N_12700,N_6281,N_8078);
nand U12701 (N_12701,N_5905,N_9662);
nand U12702 (N_12702,N_5399,N_8563);
xor U12703 (N_12703,N_5937,N_9034);
nor U12704 (N_12704,N_8045,N_7366);
or U12705 (N_12705,N_8826,N_7525);
and U12706 (N_12706,N_7824,N_7360);
or U12707 (N_12707,N_9397,N_5360);
and U12708 (N_12708,N_6263,N_7079);
xnor U12709 (N_12709,N_8969,N_9875);
nand U12710 (N_12710,N_9974,N_5214);
nand U12711 (N_12711,N_5692,N_8158);
or U12712 (N_12712,N_5748,N_8892);
nand U12713 (N_12713,N_6843,N_7921);
nor U12714 (N_12714,N_9383,N_5353);
xor U12715 (N_12715,N_6605,N_7787);
or U12716 (N_12716,N_5872,N_7473);
nand U12717 (N_12717,N_9697,N_5873);
xnor U12718 (N_12718,N_8943,N_8040);
and U12719 (N_12719,N_5567,N_7088);
xor U12720 (N_12720,N_7255,N_6524);
nor U12721 (N_12721,N_8724,N_7616);
nand U12722 (N_12722,N_5025,N_8760);
xor U12723 (N_12723,N_6877,N_8094);
and U12724 (N_12724,N_7057,N_9807);
nand U12725 (N_12725,N_6124,N_7377);
xnor U12726 (N_12726,N_7938,N_5582);
nand U12727 (N_12727,N_8504,N_8447);
and U12728 (N_12728,N_7023,N_8949);
nand U12729 (N_12729,N_6747,N_9127);
nor U12730 (N_12730,N_9452,N_9074);
and U12731 (N_12731,N_8733,N_8469);
nand U12732 (N_12732,N_8829,N_8554);
or U12733 (N_12733,N_8714,N_8934);
nand U12734 (N_12734,N_8624,N_7971);
or U12735 (N_12735,N_9460,N_9166);
or U12736 (N_12736,N_9080,N_5349);
xnor U12737 (N_12737,N_9840,N_9855);
xor U12738 (N_12738,N_5679,N_7391);
nand U12739 (N_12739,N_5086,N_5684);
nor U12740 (N_12740,N_9478,N_6346);
or U12741 (N_12741,N_7740,N_9660);
xor U12742 (N_12742,N_8586,N_5468);
or U12743 (N_12743,N_7133,N_8761);
nor U12744 (N_12744,N_9050,N_8751);
nand U12745 (N_12745,N_8220,N_9457);
or U12746 (N_12746,N_9930,N_7484);
and U12747 (N_12747,N_6200,N_8153);
xnor U12748 (N_12748,N_6139,N_7134);
nor U12749 (N_12749,N_9131,N_5386);
xnor U12750 (N_12750,N_9585,N_9125);
and U12751 (N_12751,N_9521,N_8581);
nand U12752 (N_12752,N_7867,N_8292);
nor U12753 (N_12753,N_7634,N_7129);
nor U12754 (N_12754,N_6229,N_6636);
xor U12755 (N_12755,N_9717,N_9247);
xnor U12756 (N_12756,N_5593,N_6931);
or U12757 (N_12757,N_9660,N_8481);
xnor U12758 (N_12758,N_9687,N_9254);
nand U12759 (N_12759,N_6751,N_5539);
nand U12760 (N_12760,N_9019,N_6025);
nand U12761 (N_12761,N_5945,N_5339);
nand U12762 (N_12762,N_9462,N_5730);
nand U12763 (N_12763,N_6338,N_6819);
nor U12764 (N_12764,N_5620,N_5340);
nand U12765 (N_12765,N_9368,N_5276);
nand U12766 (N_12766,N_6723,N_8303);
nand U12767 (N_12767,N_6557,N_5377);
xnor U12768 (N_12768,N_8054,N_7879);
and U12769 (N_12769,N_9536,N_8733);
nand U12770 (N_12770,N_8652,N_8034);
nand U12771 (N_12771,N_9451,N_7647);
nand U12772 (N_12772,N_8732,N_9720);
and U12773 (N_12773,N_5677,N_5131);
nand U12774 (N_12774,N_6428,N_5152);
or U12775 (N_12775,N_8264,N_6150);
or U12776 (N_12776,N_7789,N_5289);
or U12777 (N_12777,N_9102,N_6434);
xnor U12778 (N_12778,N_5830,N_6985);
and U12779 (N_12779,N_8831,N_7040);
nand U12780 (N_12780,N_6917,N_5500);
nand U12781 (N_12781,N_6311,N_7497);
nor U12782 (N_12782,N_5857,N_9160);
nand U12783 (N_12783,N_6086,N_5189);
or U12784 (N_12784,N_9464,N_7347);
or U12785 (N_12785,N_6444,N_5489);
nor U12786 (N_12786,N_5771,N_5170);
nand U12787 (N_12787,N_7787,N_6945);
nor U12788 (N_12788,N_8780,N_9282);
and U12789 (N_12789,N_5916,N_9486);
xor U12790 (N_12790,N_5906,N_7275);
and U12791 (N_12791,N_5037,N_5761);
nand U12792 (N_12792,N_7333,N_9156);
xnor U12793 (N_12793,N_9734,N_5829);
nor U12794 (N_12794,N_9511,N_7593);
or U12795 (N_12795,N_6188,N_8858);
nand U12796 (N_12796,N_5810,N_9493);
or U12797 (N_12797,N_7353,N_7128);
and U12798 (N_12798,N_7623,N_8068);
nand U12799 (N_12799,N_6810,N_5891);
and U12800 (N_12800,N_6839,N_6905);
and U12801 (N_12801,N_6331,N_5393);
nand U12802 (N_12802,N_8074,N_6914);
nor U12803 (N_12803,N_5220,N_7968);
or U12804 (N_12804,N_7323,N_8694);
nand U12805 (N_12805,N_6654,N_5613);
or U12806 (N_12806,N_7546,N_7673);
nand U12807 (N_12807,N_8214,N_5119);
nand U12808 (N_12808,N_6471,N_6257);
nor U12809 (N_12809,N_8237,N_5098);
or U12810 (N_12810,N_5150,N_8106);
xnor U12811 (N_12811,N_6349,N_6887);
and U12812 (N_12812,N_7733,N_9506);
and U12813 (N_12813,N_5820,N_9094);
xor U12814 (N_12814,N_5997,N_5470);
xnor U12815 (N_12815,N_5019,N_8771);
xor U12816 (N_12816,N_9598,N_9905);
nand U12817 (N_12817,N_5906,N_9086);
and U12818 (N_12818,N_5943,N_6339);
or U12819 (N_12819,N_6415,N_9160);
or U12820 (N_12820,N_9093,N_5769);
nand U12821 (N_12821,N_5281,N_7658);
and U12822 (N_12822,N_9991,N_9399);
and U12823 (N_12823,N_8499,N_7155);
nor U12824 (N_12824,N_5342,N_8288);
and U12825 (N_12825,N_7785,N_5411);
xnor U12826 (N_12826,N_7581,N_5178);
nand U12827 (N_12827,N_6874,N_5013);
nor U12828 (N_12828,N_6507,N_9980);
xor U12829 (N_12829,N_8863,N_9843);
and U12830 (N_12830,N_6193,N_9264);
xor U12831 (N_12831,N_7230,N_9601);
xor U12832 (N_12832,N_6058,N_8593);
and U12833 (N_12833,N_6364,N_8789);
nor U12834 (N_12834,N_5573,N_5596);
nand U12835 (N_12835,N_6953,N_9517);
and U12836 (N_12836,N_7698,N_6859);
xnor U12837 (N_12837,N_5925,N_6787);
nor U12838 (N_12838,N_7741,N_9286);
nor U12839 (N_12839,N_9221,N_9170);
and U12840 (N_12840,N_5359,N_8479);
xor U12841 (N_12841,N_7053,N_6854);
and U12842 (N_12842,N_6130,N_6063);
and U12843 (N_12843,N_7870,N_5302);
nand U12844 (N_12844,N_7022,N_5870);
nor U12845 (N_12845,N_7507,N_6865);
or U12846 (N_12846,N_9245,N_8812);
nor U12847 (N_12847,N_5763,N_5845);
and U12848 (N_12848,N_9652,N_7772);
xnor U12849 (N_12849,N_8879,N_8195);
and U12850 (N_12850,N_6105,N_5517);
xnor U12851 (N_12851,N_7571,N_6240);
nor U12852 (N_12852,N_8154,N_6525);
nand U12853 (N_12853,N_9657,N_9251);
and U12854 (N_12854,N_8129,N_9862);
and U12855 (N_12855,N_6629,N_5152);
or U12856 (N_12856,N_6997,N_5321);
xnor U12857 (N_12857,N_8496,N_5164);
xnor U12858 (N_12858,N_5869,N_8678);
or U12859 (N_12859,N_8853,N_5941);
or U12860 (N_12860,N_9471,N_9001);
xor U12861 (N_12861,N_8786,N_7428);
or U12862 (N_12862,N_5574,N_6818);
nand U12863 (N_12863,N_8052,N_6802);
or U12864 (N_12864,N_5625,N_5824);
nor U12865 (N_12865,N_9079,N_8580);
nand U12866 (N_12866,N_5115,N_7003);
nor U12867 (N_12867,N_7639,N_7257);
nor U12868 (N_12868,N_7165,N_6156);
nand U12869 (N_12869,N_6412,N_8795);
nand U12870 (N_12870,N_9472,N_6901);
nor U12871 (N_12871,N_9707,N_9819);
nand U12872 (N_12872,N_9013,N_5800);
or U12873 (N_12873,N_7095,N_8393);
xor U12874 (N_12874,N_8977,N_5568);
and U12875 (N_12875,N_6610,N_6236);
nor U12876 (N_12876,N_6609,N_9884);
or U12877 (N_12877,N_6796,N_8440);
and U12878 (N_12878,N_5287,N_9589);
nand U12879 (N_12879,N_7546,N_9447);
or U12880 (N_12880,N_9249,N_8755);
and U12881 (N_12881,N_9261,N_6490);
and U12882 (N_12882,N_5497,N_6833);
and U12883 (N_12883,N_7408,N_7286);
xnor U12884 (N_12884,N_8822,N_8264);
or U12885 (N_12885,N_7070,N_6446);
nor U12886 (N_12886,N_7665,N_8779);
or U12887 (N_12887,N_8438,N_5265);
or U12888 (N_12888,N_8481,N_7987);
and U12889 (N_12889,N_7646,N_6282);
and U12890 (N_12890,N_9979,N_6703);
nor U12891 (N_12891,N_8070,N_9702);
or U12892 (N_12892,N_7462,N_6108);
and U12893 (N_12893,N_9743,N_6505);
and U12894 (N_12894,N_7041,N_9545);
and U12895 (N_12895,N_6267,N_9485);
nor U12896 (N_12896,N_8608,N_6372);
nand U12897 (N_12897,N_9744,N_6425);
or U12898 (N_12898,N_7836,N_9796);
nand U12899 (N_12899,N_7129,N_7216);
and U12900 (N_12900,N_9989,N_7304);
nand U12901 (N_12901,N_7874,N_7195);
nor U12902 (N_12902,N_9541,N_8144);
and U12903 (N_12903,N_7870,N_5520);
nand U12904 (N_12904,N_5643,N_6758);
and U12905 (N_12905,N_9037,N_7824);
or U12906 (N_12906,N_8501,N_6116);
nand U12907 (N_12907,N_8960,N_7890);
xnor U12908 (N_12908,N_5240,N_8852);
nor U12909 (N_12909,N_6232,N_9607);
nand U12910 (N_12910,N_9057,N_8563);
or U12911 (N_12911,N_9189,N_9178);
xor U12912 (N_12912,N_7953,N_9118);
xor U12913 (N_12913,N_9856,N_7389);
xor U12914 (N_12914,N_6453,N_7067);
or U12915 (N_12915,N_6362,N_7212);
nand U12916 (N_12916,N_8976,N_7882);
nand U12917 (N_12917,N_6315,N_7993);
xor U12918 (N_12918,N_5272,N_9014);
and U12919 (N_12919,N_6693,N_6938);
or U12920 (N_12920,N_7665,N_7066);
or U12921 (N_12921,N_6732,N_6261);
or U12922 (N_12922,N_7870,N_8342);
or U12923 (N_12923,N_8473,N_8175);
or U12924 (N_12924,N_9132,N_8955);
xor U12925 (N_12925,N_6801,N_6255);
xor U12926 (N_12926,N_7239,N_6995);
nand U12927 (N_12927,N_5930,N_6125);
or U12928 (N_12928,N_6413,N_7025);
or U12929 (N_12929,N_7694,N_8679);
and U12930 (N_12930,N_6776,N_9750);
or U12931 (N_12931,N_6069,N_8868);
nor U12932 (N_12932,N_8059,N_8355);
nor U12933 (N_12933,N_8132,N_8135);
nor U12934 (N_12934,N_5577,N_8298);
or U12935 (N_12935,N_8138,N_7564);
xnor U12936 (N_12936,N_7746,N_8155);
and U12937 (N_12937,N_5501,N_7830);
or U12938 (N_12938,N_6175,N_9635);
and U12939 (N_12939,N_9477,N_6171);
and U12940 (N_12940,N_7667,N_5192);
nand U12941 (N_12941,N_9457,N_9448);
or U12942 (N_12942,N_6798,N_6146);
nor U12943 (N_12943,N_6068,N_9250);
and U12944 (N_12944,N_9885,N_7216);
nor U12945 (N_12945,N_6965,N_7686);
nand U12946 (N_12946,N_9035,N_9264);
or U12947 (N_12947,N_6218,N_8386);
nor U12948 (N_12948,N_8420,N_5946);
nand U12949 (N_12949,N_5958,N_6667);
nor U12950 (N_12950,N_9961,N_8704);
and U12951 (N_12951,N_5219,N_9129);
xor U12952 (N_12952,N_7090,N_7739);
nor U12953 (N_12953,N_9737,N_5253);
xor U12954 (N_12954,N_9121,N_5291);
xor U12955 (N_12955,N_9965,N_7955);
nand U12956 (N_12956,N_5162,N_8028);
nand U12957 (N_12957,N_9133,N_6302);
and U12958 (N_12958,N_7717,N_6726);
nand U12959 (N_12959,N_9030,N_8942);
nor U12960 (N_12960,N_6477,N_5330);
and U12961 (N_12961,N_6426,N_7242);
nor U12962 (N_12962,N_5127,N_9898);
and U12963 (N_12963,N_6202,N_7624);
or U12964 (N_12964,N_8146,N_6862);
or U12965 (N_12965,N_6188,N_7703);
and U12966 (N_12966,N_9956,N_9525);
or U12967 (N_12967,N_9571,N_8538);
xnor U12968 (N_12968,N_8474,N_6204);
xor U12969 (N_12969,N_7165,N_7272);
or U12970 (N_12970,N_5757,N_9627);
nand U12971 (N_12971,N_7449,N_9947);
xor U12972 (N_12972,N_8657,N_5649);
nor U12973 (N_12973,N_6268,N_5449);
or U12974 (N_12974,N_5197,N_5415);
nor U12975 (N_12975,N_5744,N_8907);
xnor U12976 (N_12976,N_7446,N_5848);
or U12977 (N_12977,N_6496,N_8044);
nor U12978 (N_12978,N_7064,N_6920);
nor U12979 (N_12979,N_9908,N_6513);
nand U12980 (N_12980,N_5840,N_7479);
xnor U12981 (N_12981,N_9640,N_6180);
or U12982 (N_12982,N_6888,N_9974);
or U12983 (N_12983,N_9801,N_5573);
and U12984 (N_12984,N_7689,N_8114);
or U12985 (N_12985,N_6807,N_8654);
nor U12986 (N_12986,N_7538,N_8543);
xor U12987 (N_12987,N_7878,N_6594);
nand U12988 (N_12988,N_7221,N_8347);
xnor U12989 (N_12989,N_7902,N_8033);
xor U12990 (N_12990,N_6265,N_6044);
xor U12991 (N_12991,N_6554,N_5330);
nor U12992 (N_12992,N_7611,N_5441);
xor U12993 (N_12993,N_8994,N_8448);
nor U12994 (N_12994,N_9734,N_8507);
nor U12995 (N_12995,N_7154,N_8908);
and U12996 (N_12996,N_5521,N_8326);
nor U12997 (N_12997,N_9514,N_7520);
nor U12998 (N_12998,N_5345,N_5567);
xor U12999 (N_12999,N_5437,N_9213);
or U13000 (N_13000,N_5635,N_6722);
nor U13001 (N_13001,N_8946,N_5481);
and U13002 (N_13002,N_6635,N_8807);
nor U13003 (N_13003,N_5503,N_9758);
nor U13004 (N_13004,N_6879,N_7475);
xor U13005 (N_13005,N_7732,N_7382);
xor U13006 (N_13006,N_6328,N_6570);
nor U13007 (N_13007,N_6980,N_6957);
nand U13008 (N_13008,N_7537,N_7069);
nor U13009 (N_13009,N_8246,N_9389);
nor U13010 (N_13010,N_7785,N_6321);
nor U13011 (N_13011,N_5181,N_8743);
nor U13012 (N_13012,N_5395,N_7241);
nand U13013 (N_13013,N_5715,N_6830);
nor U13014 (N_13014,N_8501,N_5446);
nor U13015 (N_13015,N_6413,N_5303);
and U13016 (N_13016,N_7727,N_5660);
or U13017 (N_13017,N_7044,N_7101);
and U13018 (N_13018,N_7188,N_9971);
or U13019 (N_13019,N_8692,N_6185);
xnor U13020 (N_13020,N_5192,N_8797);
or U13021 (N_13021,N_9101,N_9314);
xnor U13022 (N_13022,N_7996,N_9403);
or U13023 (N_13023,N_5619,N_6125);
xor U13024 (N_13024,N_5197,N_6277);
nor U13025 (N_13025,N_6660,N_6333);
nand U13026 (N_13026,N_9745,N_9726);
xnor U13027 (N_13027,N_8026,N_6566);
and U13028 (N_13028,N_7018,N_5015);
nor U13029 (N_13029,N_6703,N_7443);
nor U13030 (N_13030,N_5021,N_5589);
xor U13031 (N_13031,N_6665,N_9083);
nor U13032 (N_13032,N_6512,N_5457);
or U13033 (N_13033,N_7102,N_8425);
and U13034 (N_13034,N_6647,N_8734);
or U13035 (N_13035,N_6344,N_5383);
xnor U13036 (N_13036,N_6566,N_7184);
nand U13037 (N_13037,N_6926,N_9117);
xnor U13038 (N_13038,N_8488,N_7953);
xnor U13039 (N_13039,N_8485,N_9030);
xor U13040 (N_13040,N_9809,N_5586);
nand U13041 (N_13041,N_9157,N_5815);
or U13042 (N_13042,N_5582,N_6347);
xor U13043 (N_13043,N_6056,N_8329);
xnor U13044 (N_13044,N_6927,N_7376);
or U13045 (N_13045,N_7124,N_7629);
or U13046 (N_13046,N_6536,N_5361);
xnor U13047 (N_13047,N_5403,N_5810);
xor U13048 (N_13048,N_5550,N_7689);
and U13049 (N_13049,N_9910,N_7978);
nand U13050 (N_13050,N_9895,N_8226);
or U13051 (N_13051,N_6959,N_5646);
nand U13052 (N_13052,N_9426,N_7222);
xor U13053 (N_13053,N_9495,N_5841);
and U13054 (N_13054,N_5449,N_9815);
or U13055 (N_13055,N_8700,N_9746);
xnor U13056 (N_13056,N_8726,N_7799);
xor U13057 (N_13057,N_5299,N_9675);
nand U13058 (N_13058,N_7101,N_7386);
and U13059 (N_13059,N_7334,N_7976);
nor U13060 (N_13060,N_7254,N_8126);
xnor U13061 (N_13061,N_6751,N_8549);
xor U13062 (N_13062,N_9501,N_6074);
nor U13063 (N_13063,N_5555,N_5931);
or U13064 (N_13064,N_6939,N_7433);
or U13065 (N_13065,N_7353,N_6747);
xor U13066 (N_13066,N_9001,N_5252);
xor U13067 (N_13067,N_9077,N_7790);
nor U13068 (N_13068,N_6619,N_9061);
and U13069 (N_13069,N_7640,N_9637);
nor U13070 (N_13070,N_6657,N_9307);
xor U13071 (N_13071,N_5161,N_5980);
nor U13072 (N_13072,N_7937,N_7298);
or U13073 (N_13073,N_8786,N_8128);
or U13074 (N_13074,N_8743,N_8408);
and U13075 (N_13075,N_6879,N_5074);
nand U13076 (N_13076,N_5343,N_7469);
nor U13077 (N_13077,N_6531,N_7977);
nor U13078 (N_13078,N_8284,N_9003);
nor U13079 (N_13079,N_8730,N_6024);
nor U13080 (N_13080,N_6751,N_9832);
and U13081 (N_13081,N_6172,N_7939);
nand U13082 (N_13082,N_8224,N_5750);
nand U13083 (N_13083,N_5385,N_6235);
xor U13084 (N_13084,N_6595,N_5913);
nor U13085 (N_13085,N_7599,N_6276);
and U13086 (N_13086,N_6191,N_6513);
and U13087 (N_13087,N_9374,N_5784);
or U13088 (N_13088,N_8309,N_8413);
and U13089 (N_13089,N_6342,N_6965);
and U13090 (N_13090,N_7124,N_6213);
or U13091 (N_13091,N_7600,N_6043);
nor U13092 (N_13092,N_7090,N_8647);
nor U13093 (N_13093,N_9128,N_7423);
or U13094 (N_13094,N_5721,N_7397);
nor U13095 (N_13095,N_7668,N_8265);
nor U13096 (N_13096,N_8851,N_6005);
xor U13097 (N_13097,N_7292,N_9931);
or U13098 (N_13098,N_7647,N_8596);
xnor U13099 (N_13099,N_7629,N_5755);
nor U13100 (N_13100,N_7761,N_5098);
nor U13101 (N_13101,N_6557,N_9406);
and U13102 (N_13102,N_8532,N_5082);
or U13103 (N_13103,N_5128,N_7643);
xnor U13104 (N_13104,N_6852,N_7644);
nand U13105 (N_13105,N_9668,N_5645);
nor U13106 (N_13106,N_6452,N_7572);
xor U13107 (N_13107,N_8919,N_8903);
and U13108 (N_13108,N_9935,N_7254);
nor U13109 (N_13109,N_8044,N_7782);
xnor U13110 (N_13110,N_5789,N_8572);
or U13111 (N_13111,N_5776,N_9512);
nor U13112 (N_13112,N_9893,N_6089);
nand U13113 (N_13113,N_5481,N_6915);
nor U13114 (N_13114,N_6770,N_6049);
xor U13115 (N_13115,N_5012,N_9231);
nor U13116 (N_13116,N_8299,N_8402);
or U13117 (N_13117,N_9374,N_6401);
nor U13118 (N_13118,N_5836,N_6222);
nand U13119 (N_13119,N_7866,N_8616);
xor U13120 (N_13120,N_6283,N_7148);
or U13121 (N_13121,N_9826,N_5279);
nor U13122 (N_13122,N_9421,N_8716);
nor U13123 (N_13123,N_7076,N_6875);
nor U13124 (N_13124,N_6710,N_8248);
or U13125 (N_13125,N_9166,N_8998);
or U13126 (N_13126,N_9266,N_8673);
and U13127 (N_13127,N_6725,N_9944);
nor U13128 (N_13128,N_6749,N_8019);
xor U13129 (N_13129,N_9815,N_8719);
nor U13130 (N_13130,N_6508,N_6318);
xor U13131 (N_13131,N_8127,N_9266);
nand U13132 (N_13132,N_5482,N_9510);
nor U13133 (N_13133,N_5460,N_7127);
nand U13134 (N_13134,N_7504,N_8603);
nor U13135 (N_13135,N_5954,N_9795);
nand U13136 (N_13136,N_5616,N_5111);
or U13137 (N_13137,N_5616,N_6231);
nand U13138 (N_13138,N_5531,N_6106);
or U13139 (N_13139,N_6462,N_9569);
and U13140 (N_13140,N_8443,N_7399);
and U13141 (N_13141,N_7266,N_6589);
xor U13142 (N_13142,N_7933,N_8595);
xor U13143 (N_13143,N_6798,N_7055);
nor U13144 (N_13144,N_6613,N_5229);
or U13145 (N_13145,N_9480,N_7596);
nand U13146 (N_13146,N_6414,N_7996);
and U13147 (N_13147,N_5889,N_7398);
nand U13148 (N_13148,N_6714,N_8618);
and U13149 (N_13149,N_9030,N_9315);
nor U13150 (N_13150,N_5530,N_7559);
xnor U13151 (N_13151,N_6675,N_6237);
and U13152 (N_13152,N_9086,N_5758);
or U13153 (N_13153,N_9543,N_5901);
nor U13154 (N_13154,N_9352,N_6527);
xor U13155 (N_13155,N_6197,N_8692);
and U13156 (N_13156,N_5003,N_9523);
and U13157 (N_13157,N_9290,N_8727);
nand U13158 (N_13158,N_9009,N_9492);
nor U13159 (N_13159,N_7243,N_9039);
xnor U13160 (N_13160,N_9744,N_5389);
xnor U13161 (N_13161,N_6299,N_8520);
or U13162 (N_13162,N_9820,N_6953);
nand U13163 (N_13163,N_7003,N_5620);
or U13164 (N_13164,N_9907,N_5491);
xnor U13165 (N_13165,N_9421,N_7877);
nor U13166 (N_13166,N_6247,N_9541);
xnor U13167 (N_13167,N_9933,N_8773);
or U13168 (N_13168,N_5422,N_8941);
nand U13169 (N_13169,N_6947,N_6856);
nor U13170 (N_13170,N_9105,N_5596);
nand U13171 (N_13171,N_8531,N_8398);
and U13172 (N_13172,N_5747,N_6118);
xor U13173 (N_13173,N_9031,N_7693);
xnor U13174 (N_13174,N_5212,N_6580);
nor U13175 (N_13175,N_5608,N_5775);
xor U13176 (N_13176,N_5991,N_6452);
xnor U13177 (N_13177,N_9239,N_6267);
nand U13178 (N_13178,N_6460,N_5378);
and U13179 (N_13179,N_8993,N_8631);
or U13180 (N_13180,N_7654,N_6436);
nand U13181 (N_13181,N_5598,N_9971);
nor U13182 (N_13182,N_8239,N_8477);
xnor U13183 (N_13183,N_7916,N_6716);
and U13184 (N_13184,N_9426,N_9601);
or U13185 (N_13185,N_9257,N_6802);
xor U13186 (N_13186,N_5498,N_7138);
nand U13187 (N_13187,N_9260,N_9624);
xnor U13188 (N_13188,N_7168,N_6710);
nor U13189 (N_13189,N_6940,N_7454);
nand U13190 (N_13190,N_8476,N_8621);
nand U13191 (N_13191,N_7980,N_7635);
nand U13192 (N_13192,N_5276,N_9958);
nor U13193 (N_13193,N_6357,N_5919);
and U13194 (N_13194,N_8447,N_9110);
nor U13195 (N_13195,N_8641,N_9345);
or U13196 (N_13196,N_6908,N_5451);
and U13197 (N_13197,N_7327,N_7195);
and U13198 (N_13198,N_7513,N_6400);
or U13199 (N_13199,N_6266,N_8453);
nor U13200 (N_13200,N_7227,N_5111);
and U13201 (N_13201,N_9560,N_7953);
nor U13202 (N_13202,N_9573,N_9148);
nand U13203 (N_13203,N_6434,N_9554);
nand U13204 (N_13204,N_9956,N_5233);
nand U13205 (N_13205,N_6325,N_8901);
and U13206 (N_13206,N_5719,N_7312);
or U13207 (N_13207,N_7624,N_9668);
nor U13208 (N_13208,N_8810,N_8512);
xnor U13209 (N_13209,N_8349,N_7287);
or U13210 (N_13210,N_5920,N_7761);
or U13211 (N_13211,N_9620,N_9470);
nor U13212 (N_13212,N_7701,N_9042);
nor U13213 (N_13213,N_6140,N_8296);
and U13214 (N_13214,N_5073,N_9146);
xor U13215 (N_13215,N_6461,N_7269);
and U13216 (N_13216,N_5951,N_7202);
nand U13217 (N_13217,N_7133,N_6197);
nor U13218 (N_13218,N_5394,N_9098);
xor U13219 (N_13219,N_8530,N_6521);
and U13220 (N_13220,N_7188,N_6817);
or U13221 (N_13221,N_8322,N_6140);
and U13222 (N_13222,N_6437,N_9024);
and U13223 (N_13223,N_6655,N_7235);
nand U13224 (N_13224,N_5836,N_6415);
nor U13225 (N_13225,N_8366,N_5215);
nand U13226 (N_13226,N_5966,N_9152);
or U13227 (N_13227,N_5427,N_7213);
xnor U13228 (N_13228,N_7481,N_6213);
and U13229 (N_13229,N_6237,N_8460);
nor U13230 (N_13230,N_8519,N_8986);
nand U13231 (N_13231,N_5428,N_5952);
xnor U13232 (N_13232,N_7547,N_7057);
or U13233 (N_13233,N_9571,N_7217);
and U13234 (N_13234,N_9484,N_5273);
nor U13235 (N_13235,N_9937,N_9606);
and U13236 (N_13236,N_8893,N_7325);
and U13237 (N_13237,N_7722,N_6436);
xnor U13238 (N_13238,N_8192,N_7980);
xnor U13239 (N_13239,N_5223,N_5489);
xnor U13240 (N_13240,N_7833,N_8043);
xor U13241 (N_13241,N_8639,N_5807);
nor U13242 (N_13242,N_5590,N_8669);
and U13243 (N_13243,N_9003,N_6647);
nand U13244 (N_13244,N_5586,N_5800);
or U13245 (N_13245,N_6855,N_7308);
nand U13246 (N_13246,N_8081,N_8944);
nor U13247 (N_13247,N_5959,N_8288);
nor U13248 (N_13248,N_6508,N_7685);
and U13249 (N_13249,N_8259,N_7642);
and U13250 (N_13250,N_7605,N_7649);
and U13251 (N_13251,N_6609,N_8800);
xnor U13252 (N_13252,N_7809,N_9244);
xor U13253 (N_13253,N_8237,N_5438);
nor U13254 (N_13254,N_5439,N_5419);
nor U13255 (N_13255,N_8477,N_5165);
xor U13256 (N_13256,N_6055,N_5836);
and U13257 (N_13257,N_8412,N_6874);
nand U13258 (N_13258,N_9172,N_5157);
nand U13259 (N_13259,N_5073,N_8697);
or U13260 (N_13260,N_9284,N_7184);
or U13261 (N_13261,N_6981,N_5864);
nand U13262 (N_13262,N_8599,N_6646);
and U13263 (N_13263,N_7660,N_8801);
nand U13264 (N_13264,N_9551,N_5629);
xnor U13265 (N_13265,N_5329,N_5744);
nand U13266 (N_13266,N_9048,N_9891);
nor U13267 (N_13267,N_5217,N_5797);
nor U13268 (N_13268,N_5622,N_7476);
and U13269 (N_13269,N_8810,N_7104);
and U13270 (N_13270,N_7296,N_5281);
and U13271 (N_13271,N_9809,N_8885);
nand U13272 (N_13272,N_9651,N_8860);
nand U13273 (N_13273,N_7772,N_6831);
xnor U13274 (N_13274,N_9094,N_6748);
nand U13275 (N_13275,N_7513,N_8936);
nor U13276 (N_13276,N_9313,N_7714);
nor U13277 (N_13277,N_7115,N_7433);
nor U13278 (N_13278,N_9070,N_7732);
and U13279 (N_13279,N_5381,N_8711);
xnor U13280 (N_13280,N_9094,N_6906);
nor U13281 (N_13281,N_6864,N_6884);
or U13282 (N_13282,N_9232,N_9288);
and U13283 (N_13283,N_8676,N_8245);
nor U13284 (N_13284,N_7231,N_7133);
nor U13285 (N_13285,N_5887,N_6162);
xnor U13286 (N_13286,N_7998,N_7137);
xnor U13287 (N_13287,N_9121,N_5707);
nand U13288 (N_13288,N_6314,N_7144);
xor U13289 (N_13289,N_8552,N_8020);
or U13290 (N_13290,N_9454,N_6452);
xnor U13291 (N_13291,N_5794,N_9540);
nor U13292 (N_13292,N_9846,N_5939);
and U13293 (N_13293,N_6945,N_7373);
nor U13294 (N_13294,N_7485,N_5680);
nand U13295 (N_13295,N_6256,N_7410);
xnor U13296 (N_13296,N_5728,N_8138);
nand U13297 (N_13297,N_9128,N_5389);
or U13298 (N_13298,N_6820,N_5302);
or U13299 (N_13299,N_7730,N_6629);
or U13300 (N_13300,N_7564,N_5174);
nor U13301 (N_13301,N_6706,N_8793);
or U13302 (N_13302,N_6268,N_8376);
or U13303 (N_13303,N_5719,N_6274);
and U13304 (N_13304,N_5967,N_6836);
nor U13305 (N_13305,N_6931,N_6697);
nand U13306 (N_13306,N_9651,N_7799);
and U13307 (N_13307,N_7431,N_5212);
and U13308 (N_13308,N_9416,N_6025);
or U13309 (N_13309,N_8134,N_7655);
nor U13310 (N_13310,N_9829,N_7136);
or U13311 (N_13311,N_6786,N_5559);
nor U13312 (N_13312,N_6736,N_9735);
or U13313 (N_13313,N_8734,N_9643);
or U13314 (N_13314,N_5352,N_5769);
nand U13315 (N_13315,N_5160,N_7681);
or U13316 (N_13316,N_9457,N_7872);
or U13317 (N_13317,N_8389,N_7084);
and U13318 (N_13318,N_7347,N_5960);
nand U13319 (N_13319,N_7084,N_7932);
xor U13320 (N_13320,N_8827,N_5700);
xor U13321 (N_13321,N_6915,N_5222);
nand U13322 (N_13322,N_7895,N_9509);
or U13323 (N_13323,N_9187,N_5301);
nor U13324 (N_13324,N_5121,N_9060);
nand U13325 (N_13325,N_6645,N_9892);
nand U13326 (N_13326,N_8535,N_6571);
or U13327 (N_13327,N_7770,N_8536);
nor U13328 (N_13328,N_8471,N_8016);
nor U13329 (N_13329,N_5115,N_7425);
nor U13330 (N_13330,N_5794,N_7188);
or U13331 (N_13331,N_8656,N_8021);
xor U13332 (N_13332,N_8187,N_9359);
and U13333 (N_13333,N_6577,N_7455);
xor U13334 (N_13334,N_7654,N_6587);
and U13335 (N_13335,N_5576,N_9170);
nand U13336 (N_13336,N_8811,N_8618);
nor U13337 (N_13337,N_5945,N_9844);
xnor U13338 (N_13338,N_8846,N_6380);
or U13339 (N_13339,N_5780,N_9036);
nor U13340 (N_13340,N_5597,N_8863);
nor U13341 (N_13341,N_6831,N_8512);
nand U13342 (N_13342,N_9559,N_5239);
and U13343 (N_13343,N_6978,N_9134);
nand U13344 (N_13344,N_8537,N_5063);
and U13345 (N_13345,N_7351,N_7502);
and U13346 (N_13346,N_8430,N_9345);
and U13347 (N_13347,N_6689,N_5691);
nor U13348 (N_13348,N_8447,N_9783);
nor U13349 (N_13349,N_6299,N_6132);
nand U13350 (N_13350,N_6953,N_8892);
nand U13351 (N_13351,N_6149,N_5355);
nor U13352 (N_13352,N_7431,N_6679);
and U13353 (N_13353,N_5728,N_7092);
nand U13354 (N_13354,N_9566,N_6957);
or U13355 (N_13355,N_7565,N_8197);
nor U13356 (N_13356,N_9060,N_8758);
nor U13357 (N_13357,N_6305,N_6878);
nand U13358 (N_13358,N_7696,N_6793);
and U13359 (N_13359,N_5184,N_5917);
and U13360 (N_13360,N_6313,N_7509);
xnor U13361 (N_13361,N_5773,N_5310);
nand U13362 (N_13362,N_5172,N_8274);
or U13363 (N_13363,N_7801,N_7944);
nand U13364 (N_13364,N_6132,N_9853);
nor U13365 (N_13365,N_9609,N_5999);
xor U13366 (N_13366,N_5549,N_5454);
nand U13367 (N_13367,N_7084,N_9892);
and U13368 (N_13368,N_7992,N_5495);
nand U13369 (N_13369,N_5784,N_7405);
or U13370 (N_13370,N_6612,N_5483);
or U13371 (N_13371,N_7669,N_8555);
nor U13372 (N_13372,N_5953,N_7900);
or U13373 (N_13373,N_7509,N_9275);
and U13374 (N_13374,N_8419,N_8461);
nand U13375 (N_13375,N_9306,N_5941);
xnor U13376 (N_13376,N_7848,N_8688);
or U13377 (N_13377,N_5975,N_5803);
nor U13378 (N_13378,N_8470,N_9980);
xnor U13379 (N_13379,N_5635,N_9311);
and U13380 (N_13380,N_9853,N_7299);
or U13381 (N_13381,N_9567,N_9492);
nand U13382 (N_13382,N_6948,N_7122);
xor U13383 (N_13383,N_6541,N_6273);
nor U13384 (N_13384,N_5428,N_9854);
and U13385 (N_13385,N_7217,N_5231);
xor U13386 (N_13386,N_8908,N_8672);
or U13387 (N_13387,N_9643,N_8274);
nor U13388 (N_13388,N_5886,N_7859);
xnor U13389 (N_13389,N_8990,N_6846);
and U13390 (N_13390,N_5155,N_6281);
xor U13391 (N_13391,N_7358,N_7528);
or U13392 (N_13392,N_6682,N_8746);
nor U13393 (N_13393,N_8349,N_7956);
nor U13394 (N_13394,N_5548,N_7682);
nand U13395 (N_13395,N_6294,N_5415);
nor U13396 (N_13396,N_5012,N_9606);
or U13397 (N_13397,N_7415,N_7194);
nor U13398 (N_13398,N_8128,N_6385);
or U13399 (N_13399,N_8240,N_9536);
xor U13400 (N_13400,N_8444,N_9604);
or U13401 (N_13401,N_9264,N_8491);
nand U13402 (N_13402,N_9290,N_8762);
nor U13403 (N_13403,N_6350,N_9167);
nor U13404 (N_13404,N_7685,N_8331);
xor U13405 (N_13405,N_6455,N_5801);
and U13406 (N_13406,N_8691,N_7127);
nor U13407 (N_13407,N_7431,N_5742);
nor U13408 (N_13408,N_9451,N_6143);
and U13409 (N_13409,N_8737,N_9737);
or U13410 (N_13410,N_6966,N_5613);
xor U13411 (N_13411,N_7910,N_6675);
or U13412 (N_13412,N_8166,N_6862);
xor U13413 (N_13413,N_6323,N_7610);
xnor U13414 (N_13414,N_5435,N_9517);
nor U13415 (N_13415,N_8587,N_7092);
nand U13416 (N_13416,N_9076,N_6643);
or U13417 (N_13417,N_7058,N_9537);
or U13418 (N_13418,N_9110,N_9940);
nor U13419 (N_13419,N_6559,N_5470);
xnor U13420 (N_13420,N_6753,N_6700);
xnor U13421 (N_13421,N_6106,N_8899);
xnor U13422 (N_13422,N_9024,N_5712);
or U13423 (N_13423,N_5113,N_8873);
nand U13424 (N_13424,N_9426,N_6880);
nor U13425 (N_13425,N_5858,N_7136);
and U13426 (N_13426,N_6466,N_6670);
nand U13427 (N_13427,N_5293,N_5762);
xor U13428 (N_13428,N_8313,N_8695);
nor U13429 (N_13429,N_8827,N_6679);
xor U13430 (N_13430,N_7889,N_9571);
nand U13431 (N_13431,N_9924,N_7552);
nand U13432 (N_13432,N_8626,N_7834);
nand U13433 (N_13433,N_8403,N_5578);
or U13434 (N_13434,N_5495,N_5572);
xnor U13435 (N_13435,N_5790,N_6501);
nor U13436 (N_13436,N_9122,N_5635);
nor U13437 (N_13437,N_7281,N_5040);
xor U13438 (N_13438,N_8528,N_9332);
xnor U13439 (N_13439,N_8105,N_9092);
xor U13440 (N_13440,N_8338,N_6450);
nand U13441 (N_13441,N_7660,N_6974);
nor U13442 (N_13442,N_9715,N_7043);
nor U13443 (N_13443,N_5495,N_5397);
nand U13444 (N_13444,N_8458,N_8269);
nand U13445 (N_13445,N_6753,N_8861);
xnor U13446 (N_13446,N_6872,N_7146);
xnor U13447 (N_13447,N_5926,N_9760);
xnor U13448 (N_13448,N_9394,N_6853);
nor U13449 (N_13449,N_7215,N_6885);
and U13450 (N_13450,N_7494,N_6009);
nor U13451 (N_13451,N_6556,N_7641);
nand U13452 (N_13452,N_7323,N_5652);
and U13453 (N_13453,N_6090,N_6092);
nor U13454 (N_13454,N_5082,N_5129);
xor U13455 (N_13455,N_6127,N_5796);
nand U13456 (N_13456,N_6375,N_5601);
xnor U13457 (N_13457,N_9982,N_6007);
or U13458 (N_13458,N_7618,N_8036);
xnor U13459 (N_13459,N_8357,N_6453);
and U13460 (N_13460,N_8827,N_8725);
and U13461 (N_13461,N_6468,N_8414);
or U13462 (N_13462,N_7739,N_6837);
xor U13463 (N_13463,N_5242,N_6437);
or U13464 (N_13464,N_7690,N_6770);
nor U13465 (N_13465,N_6621,N_9386);
nand U13466 (N_13466,N_6290,N_8766);
or U13467 (N_13467,N_8993,N_7592);
nand U13468 (N_13468,N_8298,N_7885);
and U13469 (N_13469,N_6544,N_5302);
nand U13470 (N_13470,N_6938,N_8012);
and U13471 (N_13471,N_5585,N_9148);
nor U13472 (N_13472,N_9471,N_6411);
nand U13473 (N_13473,N_5762,N_8379);
xor U13474 (N_13474,N_5689,N_9315);
nand U13475 (N_13475,N_9365,N_5537);
nand U13476 (N_13476,N_7009,N_7777);
xor U13477 (N_13477,N_7221,N_8077);
and U13478 (N_13478,N_9193,N_6627);
nor U13479 (N_13479,N_9536,N_8473);
nand U13480 (N_13480,N_5885,N_9125);
xor U13481 (N_13481,N_5010,N_7118);
and U13482 (N_13482,N_5332,N_5125);
nand U13483 (N_13483,N_8075,N_8253);
xnor U13484 (N_13484,N_9212,N_7289);
nor U13485 (N_13485,N_8979,N_7772);
nor U13486 (N_13486,N_5607,N_9449);
and U13487 (N_13487,N_9067,N_9436);
nand U13488 (N_13488,N_8722,N_7429);
and U13489 (N_13489,N_8101,N_8530);
xor U13490 (N_13490,N_9085,N_7718);
and U13491 (N_13491,N_6641,N_5231);
or U13492 (N_13492,N_6314,N_6572);
nor U13493 (N_13493,N_7452,N_5287);
xnor U13494 (N_13494,N_5592,N_6257);
nand U13495 (N_13495,N_9382,N_8468);
or U13496 (N_13496,N_8235,N_7973);
xnor U13497 (N_13497,N_7685,N_6559);
nand U13498 (N_13498,N_7409,N_8744);
and U13499 (N_13499,N_9699,N_6160);
and U13500 (N_13500,N_5300,N_9605);
or U13501 (N_13501,N_6816,N_9276);
and U13502 (N_13502,N_8050,N_7931);
xor U13503 (N_13503,N_9654,N_6247);
nand U13504 (N_13504,N_8877,N_7646);
nor U13505 (N_13505,N_6488,N_6417);
nor U13506 (N_13506,N_7720,N_8148);
nand U13507 (N_13507,N_7467,N_6468);
nor U13508 (N_13508,N_8486,N_6789);
and U13509 (N_13509,N_5242,N_6730);
nor U13510 (N_13510,N_8116,N_5247);
and U13511 (N_13511,N_7610,N_9490);
or U13512 (N_13512,N_5857,N_7050);
or U13513 (N_13513,N_9563,N_7571);
nand U13514 (N_13514,N_5532,N_5625);
nor U13515 (N_13515,N_8604,N_6772);
or U13516 (N_13516,N_8444,N_6483);
xor U13517 (N_13517,N_5139,N_5713);
or U13518 (N_13518,N_7119,N_6230);
and U13519 (N_13519,N_9657,N_5878);
nand U13520 (N_13520,N_8695,N_8209);
xor U13521 (N_13521,N_9319,N_5731);
xor U13522 (N_13522,N_5818,N_6273);
xor U13523 (N_13523,N_6466,N_8222);
xor U13524 (N_13524,N_8172,N_7900);
nor U13525 (N_13525,N_9837,N_7600);
nor U13526 (N_13526,N_8187,N_8682);
xor U13527 (N_13527,N_6373,N_7606);
or U13528 (N_13528,N_8849,N_9465);
nand U13529 (N_13529,N_5964,N_8864);
xor U13530 (N_13530,N_7949,N_5160);
nand U13531 (N_13531,N_8530,N_9570);
xnor U13532 (N_13532,N_7667,N_7725);
nand U13533 (N_13533,N_8386,N_7359);
xor U13534 (N_13534,N_6254,N_8588);
xor U13535 (N_13535,N_9864,N_9458);
and U13536 (N_13536,N_7357,N_7383);
nand U13537 (N_13537,N_6812,N_7966);
nand U13538 (N_13538,N_5248,N_9070);
and U13539 (N_13539,N_7588,N_9108);
nand U13540 (N_13540,N_5212,N_8206);
nand U13541 (N_13541,N_7072,N_7763);
nand U13542 (N_13542,N_9147,N_9644);
nor U13543 (N_13543,N_5881,N_8795);
xor U13544 (N_13544,N_6326,N_6166);
or U13545 (N_13545,N_8499,N_9857);
nor U13546 (N_13546,N_8320,N_5436);
nor U13547 (N_13547,N_6193,N_8119);
xnor U13548 (N_13548,N_7378,N_9904);
nand U13549 (N_13549,N_6552,N_6691);
and U13550 (N_13550,N_8492,N_6994);
nand U13551 (N_13551,N_6283,N_5390);
or U13552 (N_13552,N_6837,N_9427);
nor U13553 (N_13553,N_8723,N_5636);
xnor U13554 (N_13554,N_6879,N_6919);
nand U13555 (N_13555,N_7348,N_9017);
nor U13556 (N_13556,N_5619,N_9903);
nor U13557 (N_13557,N_7679,N_5739);
nand U13558 (N_13558,N_6963,N_9707);
nand U13559 (N_13559,N_6766,N_5050);
nand U13560 (N_13560,N_6341,N_9012);
nor U13561 (N_13561,N_6968,N_6052);
nand U13562 (N_13562,N_6229,N_8001);
or U13563 (N_13563,N_5875,N_5228);
xnor U13564 (N_13564,N_9586,N_9378);
and U13565 (N_13565,N_6868,N_9915);
and U13566 (N_13566,N_9965,N_8617);
nand U13567 (N_13567,N_9702,N_6929);
nand U13568 (N_13568,N_9950,N_6216);
or U13569 (N_13569,N_6046,N_6989);
nand U13570 (N_13570,N_5503,N_7881);
nand U13571 (N_13571,N_5945,N_7718);
and U13572 (N_13572,N_6098,N_7070);
or U13573 (N_13573,N_9484,N_7069);
nor U13574 (N_13574,N_5778,N_5976);
nor U13575 (N_13575,N_7561,N_7250);
and U13576 (N_13576,N_8781,N_6154);
nand U13577 (N_13577,N_7596,N_9221);
nor U13578 (N_13578,N_6442,N_8152);
nand U13579 (N_13579,N_6336,N_8275);
xor U13580 (N_13580,N_8171,N_9227);
nor U13581 (N_13581,N_5285,N_8473);
and U13582 (N_13582,N_7061,N_9481);
and U13583 (N_13583,N_7921,N_9753);
and U13584 (N_13584,N_6645,N_9544);
nand U13585 (N_13585,N_7780,N_8192);
and U13586 (N_13586,N_9927,N_5663);
or U13587 (N_13587,N_8475,N_8767);
nor U13588 (N_13588,N_7652,N_9879);
nor U13589 (N_13589,N_5151,N_8282);
xnor U13590 (N_13590,N_9847,N_9003);
and U13591 (N_13591,N_6862,N_9882);
xnor U13592 (N_13592,N_6665,N_9918);
xor U13593 (N_13593,N_7106,N_5703);
xnor U13594 (N_13594,N_8802,N_7700);
and U13595 (N_13595,N_8016,N_9826);
xnor U13596 (N_13596,N_5476,N_6754);
nor U13597 (N_13597,N_9509,N_5878);
and U13598 (N_13598,N_9522,N_8309);
nor U13599 (N_13599,N_6608,N_7972);
or U13600 (N_13600,N_8647,N_9811);
nand U13601 (N_13601,N_7881,N_7904);
nand U13602 (N_13602,N_9195,N_7885);
and U13603 (N_13603,N_8036,N_8398);
nand U13604 (N_13604,N_7712,N_7822);
or U13605 (N_13605,N_8662,N_6584);
xor U13606 (N_13606,N_7740,N_9817);
xor U13607 (N_13607,N_9391,N_9814);
nor U13608 (N_13608,N_9547,N_7162);
nor U13609 (N_13609,N_5610,N_5833);
or U13610 (N_13610,N_5190,N_8916);
and U13611 (N_13611,N_5354,N_6520);
nor U13612 (N_13612,N_7672,N_5881);
and U13613 (N_13613,N_6950,N_7501);
xnor U13614 (N_13614,N_9034,N_5406);
xnor U13615 (N_13615,N_8524,N_6749);
and U13616 (N_13616,N_8834,N_8186);
xnor U13617 (N_13617,N_9772,N_8315);
xor U13618 (N_13618,N_5658,N_7912);
or U13619 (N_13619,N_6950,N_8656);
xor U13620 (N_13620,N_7276,N_8891);
xnor U13621 (N_13621,N_7796,N_6271);
xor U13622 (N_13622,N_8610,N_9386);
nand U13623 (N_13623,N_9959,N_8346);
and U13624 (N_13624,N_8882,N_9255);
and U13625 (N_13625,N_7834,N_8441);
and U13626 (N_13626,N_8752,N_6575);
nand U13627 (N_13627,N_5812,N_9431);
xnor U13628 (N_13628,N_7632,N_5929);
nand U13629 (N_13629,N_5266,N_9921);
nor U13630 (N_13630,N_9789,N_5587);
or U13631 (N_13631,N_6582,N_5903);
and U13632 (N_13632,N_6938,N_7548);
or U13633 (N_13633,N_9102,N_9264);
or U13634 (N_13634,N_7675,N_9996);
nand U13635 (N_13635,N_8911,N_5920);
nor U13636 (N_13636,N_7422,N_6096);
nand U13637 (N_13637,N_7180,N_8728);
nand U13638 (N_13638,N_9876,N_8817);
or U13639 (N_13639,N_8233,N_7212);
nand U13640 (N_13640,N_9090,N_8030);
nor U13641 (N_13641,N_6251,N_7544);
nor U13642 (N_13642,N_9600,N_5134);
xor U13643 (N_13643,N_7855,N_7067);
xnor U13644 (N_13644,N_5204,N_7768);
or U13645 (N_13645,N_7550,N_7602);
nor U13646 (N_13646,N_6915,N_9544);
nand U13647 (N_13647,N_9189,N_5988);
or U13648 (N_13648,N_6356,N_8514);
nand U13649 (N_13649,N_5159,N_6659);
xor U13650 (N_13650,N_9322,N_6589);
nor U13651 (N_13651,N_5711,N_9652);
and U13652 (N_13652,N_8099,N_6874);
nand U13653 (N_13653,N_5100,N_7851);
or U13654 (N_13654,N_6769,N_6256);
nand U13655 (N_13655,N_6912,N_8000);
or U13656 (N_13656,N_9993,N_8920);
nor U13657 (N_13657,N_9891,N_5969);
xor U13658 (N_13658,N_9996,N_9601);
or U13659 (N_13659,N_7066,N_9163);
and U13660 (N_13660,N_7821,N_6439);
and U13661 (N_13661,N_6879,N_8102);
nor U13662 (N_13662,N_5516,N_7058);
and U13663 (N_13663,N_9170,N_7797);
or U13664 (N_13664,N_8709,N_8652);
xnor U13665 (N_13665,N_9949,N_8990);
and U13666 (N_13666,N_8935,N_8200);
nand U13667 (N_13667,N_7716,N_5562);
nand U13668 (N_13668,N_9977,N_8822);
and U13669 (N_13669,N_9610,N_5312);
nor U13670 (N_13670,N_7962,N_5777);
or U13671 (N_13671,N_5678,N_6030);
nor U13672 (N_13672,N_7032,N_6068);
or U13673 (N_13673,N_9825,N_6403);
nand U13674 (N_13674,N_5178,N_9938);
nand U13675 (N_13675,N_7132,N_6333);
or U13676 (N_13676,N_8892,N_7036);
nand U13677 (N_13677,N_7810,N_6353);
and U13678 (N_13678,N_8847,N_9432);
nor U13679 (N_13679,N_9204,N_6413);
nor U13680 (N_13680,N_7010,N_7957);
xnor U13681 (N_13681,N_9539,N_6205);
xor U13682 (N_13682,N_9218,N_6216);
xor U13683 (N_13683,N_7494,N_7844);
nand U13684 (N_13684,N_5864,N_8922);
nor U13685 (N_13685,N_9721,N_6470);
nor U13686 (N_13686,N_8040,N_5955);
nand U13687 (N_13687,N_9740,N_7481);
nand U13688 (N_13688,N_9002,N_8638);
xnor U13689 (N_13689,N_5656,N_9126);
or U13690 (N_13690,N_6864,N_6096);
nor U13691 (N_13691,N_5269,N_5397);
or U13692 (N_13692,N_5910,N_5810);
nor U13693 (N_13693,N_8803,N_6891);
nand U13694 (N_13694,N_9266,N_7411);
and U13695 (N_13695,N_7301,N_5104);
nor U13696 (N_13696,N_5325,N_9271);
or U13697 (N_13697,N_6629,N_7733);
nand U13698 (N_13698,N_6360,N_6184);
nand U13699 (N_13699,N_8869,N_8319);
xor U13700 (N_13700,N_5063,N_6736);
and U13701 (N_13701,N_8448,N_5056);
or U13702 (N_13702,N_7724,N_5094);
and U13703 (N_13703,N_5403,N_7307);
or U13704 (N_13704,N_9458,N_5875);
or U13705 (N_13705,N_5057,N_8414);
nand U13706 (N_13706,N_8348,N_8853);
and U13707 (N_13707,N_9725,N_9627);
or U13708 (N_13708,N_8106,N_9758);
or U13709 (N_13709,N_9744,N_9143);
nand U13710 (N_13710,N_5062,N_5201);
nor U13711 (N_13711,N_7555,N_8975);
nor U13712 (N_13712,N_9058,N_6867);
and U13713 (N_13713,N_5382,N_5582);
nand U13714 (N_13714,N_9735,N_7714);
or U13715 (N_13715,N_9498,N_5298);
and U13716 (N_13716,N_9182,N_7780);
nor U13717 (N_13717,N_8504,N_5164);
or U13718 (N_13718,N_7205,N_6408);
nor U13719 (N_13719,N_7852,N_9337);
nor U13720 (N_13720,N_9779,N_8223);
nor U13721 (N_13721,N_5733,N_8186);
nor U13722 (N_13722,N_7689,N_5328);
nand U13723 (N_13723,N_9446,N_7372);
or U13724 (N_13724,N_8950,N_6645);
xnor U13725 (N_13725,N_8654,N_5683);
xor U13726 (N_13726,N_9402,N_7079);
nand U13727 (N_13727,N_7145,N_9305);
and U13728 (N_13728,N_9982,N_8716);
nor U13729 (N_13729,N_6943,N_9570);
or U13730 (N_13730,N_6596,N_9643);
nor U13731 (N_13731,N_9903,N_9074);
and U13732 (N_13732,N_5242,N_9697);
xnor U13733 (N_13733,N_7433,N_6694);
or U13734 (N_13734,N_6234,N_5197);
or U13735 (N_13735,N_7097,N_6480);
and U13736 (N_13736,N_8656,N_8100);
and U13737 (N_13737,N_7591,N_9222);
and U13738 (N_13738,N_8367,N_5775);
xnor U13739 (N_13739,N_5802,N_9548);
nand U13740 (N_13740,N_8271,N_9364);
xnor U13741 (N_13741,N_8902,N_5320);
nor U13742 (N_13742,N_7151,N_8719);
xor U13743 (N_13743,N_5270,N_8014);
and U13744 (N_13744,N_7969,N_9147);
and U13745 (N_13745,N_7240,N_7753);
or U13746 (N_13746,N_7447,N_9235);
xnor U13747 (N_13747,N_8850,N_6561);
and U13748 (N_13748,N_5139,N_7891);
or U13749 (N_13749,N_8012,N_6070);
nand U13750 (N_13750,N_8300,N_6015);
nand U13751 (N_13751,N_5061,N_6953);
xor U13752 (N_13752,N_6022,N_7568);
xnor U13753 (N_13753,N_9699,N_6358);
nand U13754 (N_13754,N_7259,N_5962);
or U13755 (N_13755,N_5582,N_8262);
or U13756 (N_13756,N_5742,N_9750);
nor U13757 (N_13757,N_9887,N_5817);
or U13758 (N_13758,N_6912,N_9997);
and U13759 (N_13759,N_7781,N_6850);
nor U13760 (N_13760,N_9927,N_7935);
nand U13761 (N_13761,N_6496,N_8362);
nor U13762 (N_13762,N_7688,N_9732);
xor U13763 (N_13763,N_8042,N_6067);
nand U13764 (N_13764,N_6036,N_6953);
nand U13765 (N_13765,N_6248,N_9727);
nor U13766 (N_13766,N_7463,N_5760);
or U13767 (N_13767,N_7230,N_9362);
nand U13768 (N_13768,N_7081,N_6172);
xnor U13769 (N_13769,N_9281,N_9779);
nand U13770 (N_13770,N_9868,N_9572);
xor U13771 (N_13771,N_9051,N_8967);
and U13772 (N_13772,N_7465,N_8027);
or U13773 (N_13773,N_6834,N_9001);
and U13774 (N_13774,N_5532,N_7769);
or U13775 (N_13775,N_9461,N_7859);
or U13776 (N_13776,N_9191,N_7579);
or U13777 (N_13777,N_9406,N_8955);
and U13778 (N_13778,N_8095,N_5328);
xor U13779 (N_13779,N_9494,N_8315);
nand U13780 (N_13780,N_8625,N_5362);
xor U13781 (N_13781,N_7877,N_6746);
and U13782 (N_13782,N_7176,N_5390);
or U13783 (N_13783,N_5017,N_7541);
and U13784 (N_13784,N_6880,N_9344);
nand U13785 (N_13785,N_9731,N_8034);
nor U13786 (N_13786,N_8896,N_6637);
or U13787 (N_13787,N_9401,N_7157);
or U13788 (N_13788,N_8322,N_6340);
and U13789 (N_13789,N_7559,N_5563);
xor U13790 (N_13790,N_9466,N_6365);
and U13791 (N_13791,N_5845,N_5492);
nand U13792 (N_13792,N_6531,N_8626);
or U13793 (N_13793,N_5091,N_7639);
or U13794 (N_13794,N_6701,N_7696);
xnor U13795 (N_13795,N_5271,N_8435);
nand U13796 (N_13796,N_5449,N_9660);
nand U13797 (N_13797,N_7470,N_7627);
nor U13798 (N_13798,N_6891,N_6258);
xnor U13799 (N_13799,N_6649,N_7832);
xor U13800 (N_13800,N_5863,N_7297);
and U13801 (N_13801,N_8909,N_9261);
or U13802 (N_13802,N_5900,N_9537);
or U13803 (N_13803,N_7256,N_8343);
and U13804 (N_13804,N_7649,N_8823);
or U13805 (N_13805,N_5728,N_6932);
nor U13806 (N_13806,N_6872,N_6464);
nor U13807 (N_13807,N_6089,N_7532);
and U13808 (N_13808,N_9138,N_6240);
and U13809 (N_13809,N_7412,N_5576);
and U13810 (N_13810,N_7166,N_6637);
xnor U13811 (N_13811,N_7907,N_6897);
nand U13812 (N_13812,N_8454,N_8664);
xor U13813 (N_13813,N_6778,N_5618);
or U13814 (N_13814,N_5607,N_5663);
nand U13815 (N_13815,N_5040,N_9544);
nor U13816 (N_13816,N_9168,N_5735);
xnor U13817 (N_13817,N_9953,N_9168);
nor U13818 (N_13818,N_6804,N_9424);
or U13819 (N_13819,N_6203,N_5098);
or U13820 (N_13820,N_5100,N_7431);
xnor U13821 (N_13821,N_8209,N_5594);
and U13822 (N_13822,N_8831,N_8484);
nor U13823 (N_13823,N_8362,N_7052);
or U13824 (N_13824,N_9975,N_5492);
nor U13825 (N_13825,N_9525,N_8846);
nor U13826 (N_13826,N_7603,N_7489);
or U13827 (N_13827,N_6392,N_8331);
and U13828 (N_13828,N_9492,N_6718);
nor U13829 (N_13829,N_7142,N_6809);
nor U13830 (N_13830,N_9754,N_7722);
xnor U13831 (N_13831,N_8771,N_6411);
or U13832 (N_13832,N_6295,N_5199);
xnor U13833 (N_13833,N_6138,N_6249);
nand U13834 (N_13834,N_8537,N_8389);
and U13835 (N_13835,N_7171,N_5685);
xnor U13836 (N_13836,N_6170,N_5370);
or U13837 (N_13837,N_8376,N_8211);
and U13838 (N_13838,N_8212,N_6675);
xor U13839 (N_13839,N_5087,N_6390);
or U13840 (N_13840,N_8189,N_8305);
or U13841 (N_13841,N_7087,N_5362);
or U13842 (N_13842,N_9856,N_5725);
xnor U13843 (N_13843,N_7334,N_6026);
xor U13844 (N_13844,N_9605,N_9691);
nor U13845 (N_13845,N_9393,N_8398);
or U13846 (N_13846,N_8288,N_6002);
xnor U13847 (N_13847,N_5694,N_9728);
or U13848 (N_13848,N_8763,N_7625);
nand U13849 (N_13849,N_7867,N_8377);
nor U13850 (N_13850,N_6269,N_9356);
nor U13851 (N_13851,N_7898,N_6271);
nand U13852 (N_13852,N_7649,N_8687);
or U13853 (N_13853,N_7092,N_7906);
nor U13854 (N_13854,N_8052,N_6266);
nand U13855 (N_13855,N_7217,N_5578);
nand U13856 (N_13856,N_8625,N_9607);
and U13857 (N_13857,N_9680,N_9863);
and U13858 (N_13858,N_9542,N_5831);
xor U13859 (N_13859,N_7314,N_6052);
and U13860 (N_13860,N_8983,N_7895);
nand U13861 (N_13861,N_9793,N_6516);
nor U13862 (N_13862,N_7180,N_6816);
and U13863 (N_13863,N_5139,N_9002);
xnor U13864 (N_13864,N_9589,N_6927);
or U13865 (N_13865,N_9447,N_6333);
and U13866 (N_13866,N_9118,N_6023);
nand U13867 (N_13867,N_7220,N_9337);
nor U13868 (N_13868,N_5341,N_8816);
nor U13869 (N_13869,N_8805,N_6452);
nand U13870 (N_13870,N_9407,N_8893);
or U13871 (N_13871,N_6066,N_5799);
nor U13872 (N_13872,N_7393,N_9356);
and U13873 (N_13873,N_5163,N_5769);
nor U13874 (N_13874,N_5965,N_8492);
xor U13875 (N_13875,N_9228,N_8973);
or U13876 (N_13876,N_7126,N_7272);
nor U13877 (N_13877,N_6654,N_9715);
xor U13878 (N_13878,N_7006,N_9712);
or U13879 (N_13879,N_6630,N_8573);
xnor U13880 (N_13880,N_6646,N_9325);
or U13881 (N_13881,N_6143,N_7538);
nand U13882 (N_13882,N_9767,N_9149);
nor U13883 (N_13883,N_6416,N_7181);
nor U13884 (N_13884,N_9305,N_7799);
and U13885 (N_13885,N_7939,N_5679);
nand U13886 (N_13886,N_8762,N_8938);
nand U13887 (N_13887,N_7245,N_7662);
or U13888 (N_13888,N_9255,N_9601);
and U13889 (N_13889,N_6335,N_5906);
and U13890 (N_13890,N_7368,N_7807);
or U13891 (N_13891,N_9402,N_8029);
nand U13892 (N_13892,N_7609,N_8992);
or U13893 (N_13893,N_7884,N_9519);
nand U13894 (N_13894,N_8911,N_6781);
nand U13895 (N_13895,N_5824,N_9772);
nand U13896 (N_13896,N_7230,N_5160);
nand U13897 (N_13897,N_5540,N_5028);
xnor U13898 (N_13898,N_5843,N_5427);
nor U13899 (N_13899,N_6110,N_8308);
xnor U13900 (N_13900,N_7042,N_6567);
and U13901 (N_13901,N_7526,N_6748);
xor U13902 (N_13902,N_5995,N_6677);
or U13903 (N_13903,N_6462,N_5038);
xnor U13904 (N_13904,N_6571,N_7033);
nand U13905 (N_13905,N_8243,N_5546);
nor U13906 (N_13906,N_9662,N_9381);
xnor U13907 (N_13907,N_5683,N_7313);
xor U13908 (N_13908,N_9248,N_6263);
nand U13909 (N_13909,N_6517,N_6082);
or U13910 (N_13910,N_8583,N_7627);
nand U13911 (N_13911,N_9737,N_9904);
nor U13912 (N_13912,N_5979,N_9787);
or U13913 (N_13913,N_8899,N_6156);
xor U13914 (N_13914,N_8406,N_8779);
xnor U13915 (N_13915,N_7515,N_8288);
nor U13916 (N_13916,N_5347,N_6276);
or U13917 (N_13917,N_7994,N_7416);
and U13918 (N_13918,N_6600,N_8494);
and U13919 (N_13919,N_7903,N_8839);
xor U13920 (N_13920,N_9586,N_9165);
or U13921 (N_13921,N_7781,N_9397);
xor U13922 (N_13922,N_8185,N_5145);
xor U13923 (N_13923,N_5109,N_8977);
nand U13924 (N_13924,N_9477,N_5622);
or U13925 (N_13925,N_5693,N_9620);
and U13926 (N_13926,N_9155,N_5874);
or U13927 (N_13927,N_5573,N_5256);
or U13928 (N_13928,N_8932,N_9569);
nand U13929 (N_13929,N_5554,N_8203);
or U13930 (N_13930,N_6464,N_8064);
nand U13931 (N_13931,N_7332,N_7878);
nor U13932 (N_13932,N_8230,N_7421);
or U13933 (N_13933,N_6054,N_7536);
or U13934 (N_13934,N_7021,N_9610);
xor U13935 (N_13935,N_9682,N_6579);
or U13936 (N_13936,N_9054,N_9013);
or U13937 (N_13937,N_6654,N_8976);
nor U13938 (N_13938,N_9184,N_7617);
nand U13939 (N_13939,N_9209,N_9291);
nor U13940 (N_13940,N_7516,N_8182);
or U13941 (N_13941,N_5884,N_8512);
xor U13942 (N_13942,N_5360,N_6469);
and U13943 (N_13943,N_9042,N_5745);
xnor U13944 (N_13944,N_7547,N_6571);
and U13945 (N_13945,N_9833,N_9459);
or U13946 (N_13946,N_8255,N_7784);
or U13947 (N_13947,N_5818,N_6041);
or U13948 (N_13948,N_9120,N_5829);
and U13949 (N_13949,N_6392,N_5902);
xnor U13950 (N_13950,N_8399,N_7822);
and U13951 (N_13951,N_6170,N_9961);
and U13952 (N_13952,N_9635,N_7898);
nor U13953 (N_13953,N_9352,N_8264);
xor U13954 (N_13954,N_7572,N_6432);
nor U13955 (N_13955,N_9287,N_7535);
xor U13956 (N_13956,N_5765,N_9419);
and U13957 (N_13957,N_8635,N_6965);
or U13958 (N_13958,N_8199,N_7416);
nor U13959 (N_13959,N_6260,N_9409);
nand U13960 (N_13960,N_9223,N_7973);
and U13961 (N_13961,N_8411,N_5705);
nand U13962 (N_13962,N_9450,N_8427);
nand U13963 (N_13963,N_7126,N_7427);
and U13964 (N_13964,N_8583,N_7472);
xnor U13965 (N_13965,N_5382,N_7554);
nand U13966 (N_13966,N_9866,N_9487);
xnor U13967 (N_13967,N_5642,N_9729);
xor U13968 (N_13968,N_8481,N_6295);
and U13969 (N_13969,N_7962,N_7005);
xnor U13970 (N_13970,N_9327,N_5020);
and U13971 (N_13971,N_8445,N_5171);
or U13972 (N_13972,N_7375,N_9555);
or U13973 (N_13973,N_9791,N_6638);
xor U13974 (N_13974,N_7715,N_7610);
and U13975 (N_13975,N_7203,N_5487);
xnor U13976 (N_13976,N_7940,N_9713);
nand U13977 (N_13977,N_6842,N_8565);
or U13978 (N_13978,N_6244,N_6855);
or U13979 (N_13979,N_7552,N_7149);
or U13980 (N_13980,N_6973,N_9284);
nor U13981 (N_13981,N_6798,N_8694);
nor U13982 (N_13982,N_7452,N_7662);
nor U13983 (N_13983,N_9517,N_5133);
xor U13984 (N_13984,N_5788,N_7464);
xor U13985 (N_13985,N_8328,N_7404);
xnor U13986 (N_13986,N_5203,N_6319);
nor U13987 (N_13987,N_9475,N_9206);
nor U13988 (N_13988,N_7670,N_6628);
nand U13989 (N_13989,N_5522,N_7418);
nor U13990 (N_13990,N_7989,N_9873);
nor U13991 (N_13991,N_9090,N_7858);
nor U13992 (N_13992,N_7975,N_7827);
or U13993 (N_13993,N_9387,N_7989);
nor U13994 (N_13994,N_8278,N_9957);
and U13995 (N_13995,N_5768,N_6407);
nand U13996 (N_13996,N_8296,N_5566);
xnor U13997 (N_13997,N_8074,N_8615);
nand U13998 (N_13998,N_6495,N_9885);
and U13999 (N_13999,N_5650,N_6557);
nand U14000 (N_14000,N_5595,N_7607);
and U14001 (N_14001,N_9550,N_8678);
and U14002 (N_14002,N_6487,N_6158);
xnor U14003 (N_14003,N_7851,N_8700);
and U14004 (N_14004,N_6406,N_6139);
xnor U14005 (N_14005,N_8569,N_6685);
nor U14006 (N_14006,N_7138,N_5683);
nor U14007 (N_14007,N_7214,N_6325);
or U14008 (N_14008,N_9710,N_5270);
nand U14009 (N_14009,N_7410,N_6244);
or U14010 (N_14010,N_6893,N_5920);
nor U14011 (N_14011,N_5553,N_9355);
nor U14012 (N_14012,N_7379,N_6183);
nor U14013 (N_14013,N_8182,N_6018);
nor U14014 (N_14014,N_9549,N_7299);
xnor U14015 (N_14015,N_5452,N_5012);
or U14016 (N_14016,N_6891,N_5646);
nor U14017 (N_14017,N_8587,N_6868);
and U14018 (N_14018,N_8381,N_8605);
xor U14019 (N_14019,N_7912,N_6422);
xor U14020 (N_14020,N_8892,N_9865);
nor U14021 (N_14021,N_5057,N_8633);
and U14022 (N_14022,N_9325,N_7962);
nor U14023 (N_14023,N_6836,N_6782);
and U14024 (N_14024,N_7519,N_6005);
or U14025 (N_14025,N_7770,N_6661);
or U14026 (N_14026,N_5372,N_7484);
nor U14027 (N_14027,N_9284,N_7031);
nand U14028 (N_14028,N_8945,N_5263);
nor U14029 (N_14029,N_9311,N_6408);
xor U14030 (N_14030,N_5743,N_8486);
and U14031 (N_14031,N_6864,N_9318);
xor U14032 (N_14032,N_9362,N_5518);
and U14033 (N_14033,N_8276,N_9672);
xor U14034 (N_14034,N_8715,N_7642);
and U14035 (N_14035,N_9093,N_5055);
or U14036 (N_14036,N_8657,N_5275);
nor U14037 (N_14037,N_6347,N_9548);
nor U14038 (N_14038,N_8883,N_9528);
nand U14039 (N_14039,N_7472,N_5300);
or U14040 (N_14040,N_9667,N_9267);
nand U14041 (N_14041,N_9317,N_5294);
nand U14042 (N_14042,N_7463,N_8942);
xnor U14043 (N_14043,N_6198,N_6975);
xor U14044 (N_14044,N_5097,N_5047);
nor U14045 (N_14045,N_7733,N_5495);
nor U14046 (N_14046,N_6304,N_6590);
xor U14047 (N_14047,N_7934,N_9027);
nor U14048 (N_14048,N_9433,N_9823);
nor U14049 (N_14049,N_9686,N_7521);
or U14050 (N_14050,N_5464,N_6214);
or U14051 (N_14051,N_9331,N_6739);
or U14052 (N_14052,N_7239,N_9451);
or U14053 (N_14053,N_8621,N_6767);
nand U14054 (N_14054,N_5200,N_9708);
nand U14055 (N_14055,N_5765,N_9103);
xnor U14056 (N_14056,N_8319,N_8880);
and U14057 (N_14057,N_9574,N_6489);
xnor U14058 (N_14058,N_5935,N_6957);
and U14059 (N_14059,N_5269,N_5424);
xnor U14060 (N_14060,N_6518,N_6583);
nor U14061 (N_14061,N_8833,N_5234);
nor U14062 (N_14062,N_9188,N_6747);
nand U14063 (N_14063,N_6937,N_5783);
or U14064 (N_14064,N_6911,N_5776);
xor U14065 (N_14065,N_9041,N_9781);
nor U14066 (N_14066,N_7323,N_9378);
nand U14067 (N_14067,N_5791,N_6975);
or U14068 (N_14068,N_5082,N_5433);
and U14069 (N_14069,N_8984,N_6974);
nor U14070 (N_14070,N_9050,N_9577);
nor U14071 (N_14071,N_6638,N_8787);
or U14072 (N_14072,N_9837,N_6210);
and U14073 (N_14073,N_6042,N_5827);
or U14074 (N_14074,N_8908,N_5411);
xor U14075 (N_14075,N_5328,N_6527);
nand U14076 (N_14076,N_6988,N_8993);
and U14077 (N_14077,N_8972,N_9796);
xnor U14078 (N_14078,N_7631,N_6630);
xnor U14079 (N_14079,N_9045,N_5485);
nor U14080 (N_14080,N_6984,N_6864);
nand U14081 (N_14081,N_9871,N_7290);
nor U14082 (N_14082,N_5509,N_6505);
xor U14083 (N_14083,N_6242,N_5234);
nand U14084 (N_14084,N_5689,N_5516);
nor U14085 (N_14085,N_6087,N_6759);
and U14086 (N_14086,N_9055,N_5552);
nand U14087 (N_14087,N_5174,N_9215);
and U14088 (N_14088,N_5910,N_8501);
nand U14089 (N_14089,N_7832,N_7222);
and U14090 (N_14090,N_8098,N_8965);
nand U14091 (N_14091,N_6397,N_8879);
xor U14092 (N_14092,N_6177,N_6702);
nand U14093 (N_14093,N_7468,N_8451);
xor U14094 (N_14094,N_5762,N_9365);
and U14095 (N_14095,N_9093,N_9813);
xnor U14096 (N_14096,N_6432,N_8483);
nand U14097 (N_14097,N_8493,N_6924);
xor U14098 (N_14098,N_6588,N_6308);
nor U14099 (N_14099,N_6676,N_6643);
nand U14100 (N_14100,N_8673,N_9185);
xnor U14101 (N_14101,N_7193,N_6761);
and U14102 (N_14102,N_8008,N_6436);
nor U14103 (N_14103,N_8589,N_6680);
nor U14104 (N_14104,N_8361,N_5563);
xnor U14105 (N_14105,N_7512,N_9994);
or U14106 (N_14106,N_6018,N_8440);
nor U14107 (N_14107,N_8885,N_7446);
xnor U14108 (N_14108,N_6596,N_9466);
nand U14109 (N_14109,N_7387,N_6418);
xnor U14110 (N_14110,N_8639,N_7641);
nand U14111 (N_14111,N_6666,N_7748);
and U14112 (N_14112,N_8743,N_9309);
xor U14113 (N_14113,N_9771,N_9018);
and U14114 (N_14114,N_5141,N_7797);
nor U14115 (N_14115,N_7983,N_6081);
and U14116 (N_14116,N_8872,N_8466);
and U14117 (N_14117,N_5573,N_8866);
nand U14118 (N_14118,N_8742,N_7471);
xor U14119 (N_14119,N_5126,N_5262);
xor U14120 (N_14120,N_7078,N_7662);
nor U14121 (N_14121,N_9534,N_5958);
and U14122 (N_14122,N_5929,N_7245);
nor U14123 (N_14123,N_6727,N_6755);
nor U14124 (N_14124,N_9602,N_8235);
xor U14125 (N_14125,N_8036,N_9793);
or U14126 (N_14126,N_5948,N_5786);
nand U14127 (N_14127,N_5503,N_8522);
or U14128 (N_14128,N_6430,N_6891);
or U14129 (N_14129,N_9497,N_9595);
and U14130 (N_14130,N_8201,N_6728);
or U14131 (N_14131,N_7219,N_7975);
and U14132 (N_14132,N_6073,N_6053);
nor U14133 (N_14133,N_5565,N_6290);
nor U14134 (N_14134,N_5421,N_6926);
nor U14135 (N_14135,N_9077,N_7652);
or U14136 (N_14136,N_5428,N_7372);
nand U14137 (N_14137,N_7311,N_6730);
nor U14138 (N_14138,N_9675,N_8872);
or U14139 (N_14139,N_6722,N_5085);
or U14140 (N_14140,N_6507,N_6745);
xor U14141 (N_14141,N_8308,N_9656);
nand U14142 (N_14142,N_6339,N_9081);
nand U14143 (N_14143,N_8000,N_6322);
xnor U14144 (N_14144,N_9768,N_6652);
xor U14145 (N_14145,N_6686,N_8267);
and U14146 (N_14146,N_5827,N_9803);
xnor U14147 (N_14147,N_6349,N_8231);
nand U14148 (N_14148,N_9183,N_5420);
or U14149 (N_14149,N_6563,N_7040);
or U14150 (N_14150,N_5477,N_5737);
nand U14151 (N_14151,N_5672,N_6980);
nor U14152 (N_14152,N_6801,N_9755);
nand U14153 (N_14153,N_7865,N_9904);
nor U14154 (N_14154,N_9796,N_6131);
or U14155 (N_14155,N_7867,N_8557);
xnor U14156 (N_14156,N_7402,N_6858);
and U14157 (N_14157,N_6484,N_9844);
nand U14158 (N_14158,N_7439,N_6327);
nand U14159 (N_14159,N_7952,N_6980);
or U14160 (N_14160,N_8250,N_6295);
nand U14161 (N_14161,N_7853,N_5214);
and U14162 (N_14162,N_5990,N_7675);
and U14163 (N_14163,N_8143,N_6852);
or U14164 (N_14164,N_6167,N_5742);
xor U14165 (N_14165,N_9257,N_6645);
nand U14166 (N_14166,N_6663,N_8593);
nand U14167 (N_14167,N_6183,N_5459);
nor U14168 (N_14168,N_8661,N_7962);
or U14169 (N_14169,N_8873,N_8126);
nand U14170 (N_14170,N_6483,N_6053);
nand U14171 (N_14171,N_5746,N_7250);
nor U14172 (N_14172,N_9251,N_7055);
nor U14173 (N_14173,N_7574,N_9785);
or U14174 (N_14174,N_7526,N_9488);
and U14175 (N_14175,N_8887,N_7239);
nand U14176 (N_14176,N_8137,N_9392);
xor U14177 (N_14177,N_9100,N_7001);
nor U14178 (N_14178,N_6441,N_5015);
and U14179 (N_14179,N_9737,N_7222);
xnor U14180 (N_14180,N_6895,N_8343);
xnor U14181 (N_14181,N_8332,N_7148);
and U14182 (N_14182,N_7242,N_5422);
xnor U14183 (N_14183,N_8176,N_7169);
nand U14184 (N_14184,N_6533,N_9046);
nor U14185 (N_14185,N_8924,N_5755);
or U14186 (N_14186,N_8251,N_8111);
nand U14187 (N_14187,N_9247,N_8929);
and U14188 (N_14188,N_7830,N_8326);
nor U14189 (N_14189,N_7148,N_8181);
or U14190 (N_14190,N_6320,N_6287);
nand U14191 (N_14191,N_9912,N_7031);
and U14192 (N_14192,N_6225,N_7265);
or U14193 (N_14193,N_6874,N_8221);
or U14194 (N_14194,N_6422,N_9029);
xor U14195 (N_14195,N_9413,N_7760);
or U14196 (N_14196,N_9647,N_7743);
xor U14197 (N_14197,N_6573,N_7316);
nor U14198 (N_14198,N_8627,N_7642);
and U14199 (N_14199,N_7743,N_7789);
and U14200 (N_14200,N_5417,N_7847);
and U14201 (N_14201,N_8166,N_9481);
and U14202 (N_14202,N_6808,N_6715);
nand U14203 (N_14203,N_9511,N_7720);
xor U14204 (N_14204,N_7986,N_9382);
nand U14205 (N_14205,N_8688,N_7614);
or U14206 (N_14206,N_7423,N_5435);
nor U14207 (N_14207,N_8612,N_9477);
or U14208 (N_14208,N_5942,N_5608);
or U14209 (N_14209,N_8017,N_6426);
and U14210 (N_14210,N_8073,N_5115);
or U14211 (N_14211,N_8805,N_6859);
or U14212 (N_14212,N_5263,N_6811);
xor U14213 (N_14213,N_5753,N_6701);
nand U14214 (N_14214,N_7003,N_7615);
xor U14215 (N_14215,N_9548,N_9590);
xor U14216 (N_14216,N_5167,N_5760);
nand U14217 (N_14217,N_7551,N_5973);
or U14218 (N_14218,N_7625,N_8266);
xor U14219 (N_14219,N_9088,N_7283);
xor U14220 (N_14220,N_7070,N_6896);
nor U14221 (N_14221,N_6582,N_7190);
and U14222 (N_14222,N_5588,N_6039);
nor U14223 (N_14223,N_8430,N_5640);
nor U14224 (N_14224,N_8917,N_6913);
or U14225 (N_14225,N_5058,N_9436);
nand U14226 (N_14226,N_5075,N_9367);
nand U14227 (N_14227,N_9207,N_9316);
nor U14228 (N_14228,N_7256,N_6915);
nand U14229 (N_14229,N_8532,N_7162);
and U14230 (N_14230,N_8160,N_8015);
or U14231 (N_14231,N_7805,N_8458);
xnor U14232 (N_14232,N_9689,N_6738);
nand U14233 (N_14233,N_9871,N_5117);
or U14234 (N_14234,N_5743,N_6618);
nand U14235 (N_14235,N_9735,N_5092);
nor U14236 (N_14236,N_9811,N_6476);
nor U14237 (N_14237,N_8909,N_5755);
nand U14238 (N_14238,N_8835,N_6679);
or U14239 (N_14239,N_6599,N_8670);
xor U14240 (N_14240,N_7994,N_5935);
and U14241 (N_14241,N_6699,N_9613);
xor U14242 (N_14242,N_9445,N_8708);
and U14243 (N_14243,N_9856,N_9747);
nand U14244 (N_14244,N_9545,N_6962);
and U14245 (N_14245,N_8715,N_7661);
and U14246 (N_14246,N_9100,N_6870);
xor U14247 (N_14247,N_7634,N_8866);
nor U14248 (N_14248,N_5263,N_9535);
xnor U14249 (N_14249,N_9494,N_7251);
xor U14250 (N_14250,N_8075,N_9929);
and U14251 (N_14251,N_9749,N_7343);
or U14252 (N_14252,N_6264,N_7747);
or U14253 (N_14253,N_8578,N_9592);
nor U14254 (N_14254,N_6440,N_5705);
nand U14255 (N_14255,N_8809,N_8667);
nand U14256 (N_14256,N_6167,N_6004);
nor U14257 (N_14257,N_8698,N_7297);
nand U14258 (N_14258,N_9064,N_5541);
xnor U14259 (N_14259,N_6669,N_9542);
or U14260 (N_14260,N_9493,N_6748);
or U14261 (N_14261,N_9325,N_5006);
nand U14262 (N_14262,N_6072,N_9420);
xor U14263 (N_14263,N_6414,N_8438);
xor U14264 (N_14264,N_9633,N_6935);
nor U14265 (N_14265,N_7097,N_8567);
xor U14266 (N_14266,N_6470,N_9966);
nor U14267 (N_14267,N_8495,N_9133);
nand U14268 (N_14268,N_5920,N_9497);
nor U14269 (N_14269,N_9997,N_9290);
nor U14270 (N_14270,N_7612,N_7501);
xnor U14271 (N_14271,N_7708,N_7774);
and U14272 (N_14272,N_7769,N_6465);
xnor U14273 (N_14273,N_5651,N_5442);
and U14274 (N_14274,N_6331,N_7325);
nor U14275 (N_14275,N_8444,N_9763);
xor U14276 (N_14276,N_6296,N_7013);
nand U14277 (N_14277,N_7014,N_5968);
or U14278 (N_14278,N_5596,N_9592);
nor U14279 (N_14279,N_8008,N_6519);
nand U14280 (N_14280,N_7578,N_7601);
or U14281 (N_14281,N_9156,N_5381);
xor U14282 (N_14282,N_9206,N_8596);
or U14283 (N_14283,N_6607,N_8788);
nand U14284 (N_14284,N_7765,N_6631);
or U14285 (N_14285,N_6420,N_6128);
and U14286 (N_14286,N_9744,N_7873);
xnor U14287 (N_14287,N_9357,N_6411);
nand U14288 (N_14288,N_7491,N_7211);
or U14289 (N_14289,N_8606,N_9584);
nand U14290 (N_14290,N_7601,N_5456);
nand U14291 (N_14291,N_5599,N_5785);
nand U14292 (N_14292,N_9994,N_8212);
nor U14293 (N_14293,N_6854,N_6915);
xor U14294 (N_14294,N_7124,N_9782);
nand U14295 (N_14295,N_8620,N_6225);
nor U14296 (N_14296,N_7783,N_9961);
and U14297 (N_14297,N_9113,N_6340);
xnor U14298 (N_14298,N_9273,N_7836);
or U14299 (N_14299,N_5018,N_5697);
and U14300 (N_14300,N_5826,N_9695);
and U14301 (N_14301,N_6323,N_9982);
nand U14302 (N_14302,N_6139,N_9287);
or U14303 (N_14303,N_7551,N_5998);
and U14304 (N_14304,N_7762,N_9326);
or U14305 (N_14305,N_9343,N_8244);
nor U14306 (N_14306,N_9676,N_9998);
nor U14307 (N_14307,N_9133,N_8957);
and U14308 (N_14308,N_7196,N_9877);
nor U14309 (N_14309,N_7313,N_6927);
and U14310 (N_14310,N_8256,N_8192);
nand U14311 (N_14311,N_8644,N_8722);
nand U14312 (N_14312,N_6329,N_5479);
nand U14313 (N_14313,N_5078,N_9613);
or U14314 (N_14314,N_5845,N_9405);
xnor U14315 (N_14315,N_5412,N_5492);
or U14316 (N_14316,N_9692,N_6344);
nor U14317 (N_14317,N_7038,N_7317);
xor U14318 (N_14318,N_9104,N_9353);
xor U14319 (N_14319,N_5050,N_6819);
xor U14320 (N_14320,N_6550,N_8845);
or U14321 (N_14321,N_6941,N_7034);
nand U14322 (N_14322,N_7822,N_5127);
xnor U14323 (N_14323,N_8280,N_6229);
nand U14324 (N_14324,N_9931,N_6035);
and U14325 (N_14325,N_6608,N_7914);
and U14326 (N_14326,N_6704,N_7241);
or U14327 (N_14327,N_9510,N_9465);
xnor U14328 (N_14328,N_9741,N_5676);
and U14329 (N_14329,N_8207,N_7989);
nand U14330 (N_14330,N_5588,N_6635);
or U14331 (N_14331,N_8180,N_8350);
nand U14332 (N_14332,N_9239,N_6252);
xnor U14333 (N_14333,N_5788,N_9023);
or U14334 (N_14334,N_8379,N_6219);
xnor U14335 (N_14335,N_6783,N_7060);
xor U14336 (N_14336,N_7741,N_5831);
and U14337 (N_14337,N_9370,N_6280);
xor U14338 (N_14338,N_5454,N_8500);
nand U14339 (N_14339,N_5932,N_7483);
nand U14340 (N_14340,N_8186,N_5693);
xnor U14341 (N_14341,N_9617,N_8997);
and U14342 (N_14342,N_5267,N_5664);
nand U14343 (N_14343,N_7414,N_9361);
or U14344 (N_14344,N_7343,N_6764);
and U14345 (N_14345,N_9175,N_5041);
xnor U14346 (N_14346,N_5596,N_9248);
and U14347 (N_14347,N_9095,N_9387);
nand U14348 (N_14348,N_9650,N_5343);
nand U14349 (N_14349,N_6976,N_8798);
nand U14350 (N_14350,N_9462,N_5785);
xnor U14351 (N_14351,N_9990,N_9727);
and U14352 (N_14352,N_7547,N_8618);
xor U14353 (N_14353,N_5673,N_6938);
nor U14354 (N_14354,N_5440,N_9961);
nand U14355 (N_14355,N_9213,N_6201);
nand U14356 (N_14356,N_6046,N_5823);
nor U14357 (N_14357,N_5164,N_5427);
or U14358 (N_14358,N_6052,N_6652);
and U14359 (N_14359,N_6808,N_9715);
nor U14360 (N_14360,N_8431,N_9990);
or U14361 (N_14361,N_6795,N_8548);
or U14362 (N_14362,N_7538,N_7720);
and U14363 (N_14363,N_8603,N_6630);
or U14364 (N_14364,N_8959,N_9954);
xor U14365 (N_14365,N_8766,N_8982);
and U14366 (N_14366,N_8084,N_5841);
or U14367 (N_14367,N_6836,N_7566);
nor U14368 (N_14368,N_9789,N_6775);
and U14369 (N_14369,N_9730,N_5676);
and U14370 (N_14370,N_9091,N_7696);
nor U14371 (N_14371,N_9833,N_5375);
and U14372 (N_14372,N_5327,N_8185);
nor U14373 (N_14373,N_7522,N_8967);
nand U14374 (N_14374,N_8248,N_8924);
nand U14375 (N_14375,N_8795,N_8638);
nor U14376 (N_14376,N_5273,N_9698);
and U14377 (N_14377,N_9005,N_6749);
and U14378 (N_14378,N_7682,N_5081);
or U14379 (N_14379,N_6248,N_6713);
or U14380 (N_14380,N_9338,N_6807);
or U14381 (N_14381,N_5272,N_7288);
and U14382 (N_14382,N_9233,N_7550);
nand U14383 (N_14383,N_5776,N_8268);
xor U14384 (N_14384,N_5900,N_7204);
nor U14385 (N_14385,N_7687,N_6058);
xor U14386 (N_14386,N_7134,N_8590);
nor U14387 (N_14387,N_8203,N_6816);
xnor U14388 (N_14388,N_5614,N_8896);
or U14389 (N_14389,N_8575,N_7068);
and U14390 (N_14390,N_7619,N_9616);
xor U14391 (N_14391,N_8790,N_7665);
or U14392 (N_14392,N_8676,N_7962);
and U14393 (N_14393,N_5151,N_8197);
and U14394 (N_14394,N_8882,N_9550);
nand U14395 (N_14395,N_9720,N_9973);
or U14396 (N_14396,N_8189,N_5130);
or U14397 (N_14397,N_8234,N_6486);
or U14398 (N_14398,N_8348,N_7407);
or U14399 (N_14399,N_5427,N_8535);
xor U14400 (N_14400,N_9033,N_5599);
or U14401 (N_14401,N_6749,N_9319);
nor U14402 (N_14402,N_9915,N_5200);
or U14403 (N_14403,N_6202,N_6678);
nand U14404 (N_14404,N_8904,N_9853);
nor U14405 (N_14405,N_8161,N_7695);
nor U14406 (N_14406,N_6526,N_8482);
nor U14407 (N_14407,N_9684,N_8052);
nand U14408 (N_14408,N_6727,N_9733);
nor U14409 (N_14409,N_7258,N_6382);
xor U14410 (N_14410,N_6743,N_5402);
nand U14411 (N_14411,N_5724,N_7053);
and U14412 (N_14412,N_6570,N_5442);
nand U14413 (N_14413,N_6489,N_9471);
xor U14414 (N_14414,N_6227,N_6187);
nand U14415 (N_14415,N_9298,N_9777);
nand U14416 (N_14416,N_7488,N_8806);
nor U14417 (N_14417,N_9664,N_9565);
nand U14418 (N_14418,N_8707,N_7890);
nand U14419 (N_14419,N_5947,N_9916);
and U14420 (N_14420,N_5772,N_6780);
or U14421 (N_14421,N_7694,N_5849);
xor U14422 (N_14422,N_5193,N_6612);
or U14423 (N_14423,N_8990,N_5309);
or U14424 (N_14424,N_7490,N_7565);
nor U14425 (N_14425,N_5519,N_7965);
and U14426 (N_14426,N_6636,N_6973);
nand U14427 (N_14427,N_6601,N_6335);
nor U14428 (N_14428,N_5980,N_5841);
nor U14429 (N_14429,N_7246,N_7950);
nand U14430 (N_14430,N_6917,N_5915);
xnor U14431 (N_14431,N_7143,N_5704);
or U14432 (N_14432,N_6603,N_6026);
nand U14433 (N_14433,N_6995,N_5258);
or U14434 (N_14434,N_8724,N_8875);
or U14435 (N_14435,N_9486,N_8105);
and U14436 (N_14436,N_9691,N_5641);
and U14437 (N_14437,N_5030,N_8968);
or U14438 (N_14438,N_7594,N_7236);
or U14439 (N_14439,N_5553,N_9175);
nor U14440 (N_14440,N_9411,N_9362);
nor U14441 (N_14441,N_6326,N_5526);
or U14442 (N_14442,N_6262,N_8946);
nor U14443 (N_14443,N_8628,N_8344);
or U14444 (N_14444,N_6826,N_7882);
xnor U14445 (N_14445,N_8439,N_9114);
xor U14446 (N_14446,N_8584,N_6291);
xnor U14447 (N_14447,N_7534,N_8606);
nor U14448 (N_14448,N_8893,N_7306);
xnor U14449 (N_14449,N_7895,N_8788);
nor U14450 (N_14450,N_6310,N_6169);
nand U14451 (N_14451,N_8696,N_7411);
and U14452 (N_14452,N_8689,N_9003);
xor U14453 (N_14453,N_5582,N_6018);
or U14454 (N_14454,N_7278,N_8476);
and U14455 (N_14455,N_8905,N_8352);
or U14456 (N_14456,N_7305,N_9677);
xor U14457 (N_14457,N_5144,N_6387);
xnor U14458 (N_14458,N_6959,N_9628);
nand U14459 (N_14459,N_6153,N_7643);
nor U14460 (N_14460,N_5423,N_8360);
and U14461 (N_14461,N_5925,N_9612);
nor U14462 (N_14462,N_9323,N_5587);
and U14463 (N_14463,N_7205,N_9708);
xor U14464 (N_14464,N_8229,N_6529);
nor U14465 (N_14465,N_6748,N_7299);
or U14466 (N_14466,N_7744,N_6043);
nand U14467 (N_14467,N_8595,N_5831);
nor U14468 (N_14468,N_8310,N_8498);
nand U14469 (N_14469,N_8653,N_6289);
xor U14470 (N_14470,N_5550,N_7488);
nor U14471 (N_14471,N_8791,N_6157);
nand U14472 (N_14472,N_7045,N_8476);
nor U14473 (N_14473,N_7932,N_5577);
nand U14474 (N_14474,N_6911,N_8976);
and U14475 (N_14475,N_8496,N_5666);
nand U14476 (N_14476,N_8957,N_8159);
nand U14477 (N_14477,N_7800,N_6369);
nor U14478 (N_14478,N_9637,N_8659);
and U14479 (N_14479,N_5776,N_8733);
or U14480 (N_14480,N_9189,N_7717);
nand U14481 (N_14481,N_6734,N_6337);
and U14482 (N_14482,N_6971,N_9869);
nor U14483 (N_14483,N_5941,N_7173);
nor U14484 (N_14484,N_6741,N_8977);
nand U14485 (N_14485,N_8170,N_8837);
nor U14486 (N_14486,N_5340,N_9659);
nand U14487 (N_14487,N_9084,N_5827);
nand U14488 (N_14488,N_5015,N_7184);
and U14489 (N_14489,N_5098,N_9328);
and U14490 (N_14490,N_6101,N_8195);
and U14491 (N_14491,N_9075,N_8402);
nor U14492 (N_14492,N_6758,N_6076);
xnor U14493 (N_14493,N_9192,N_8019);
nand U14494 (N_14494,N_8997,N_5629);
nand U14495 (N_14495,N_9102,N_8323);
nor U14496 (N_14496,N_6093,N_9979);
xnor U14497 (N_14497,N_5357,N_9331);
nor U14498 (N_14498,N_9637,N_6852);
xnor U14499 (N_14499,N_9149,N_5545);
and U14500 (N_14500,N_5356,N_7262);
xnor U14501 (N_14501,N_9707,N_5957);
xnor U14502 (N_14502,N_5345,N_6558);
nand U14503 (N_14503,N_5880,N_6823);
nor U14504 (N_14504,N_7402,N_7842);
and U14505 (N_14505,N_5547,N_7467);
and U14506 (N_14506,N_9819,N_9314);
or U14507 (N_14507,N_9084,N_7148);
nand U14508 (N_14508,N_7390,N_6572);
and U14509 (N_14509,N_7959,N_8732);
or U14510 (N_14510,N_7061,N_8283);
and U14511 (N_14511,N_9815,N_6107);
nor U14512 (N_14512,N_5995,N_8068);
or U14513 (N_14513,N_9461,N_8055);
or U14514 (N_14514,N_6638,N_5441);
or U14515 (N_14515,N_5772,N_6750);
or U14516 (N_14516,N_5445,N_5098);
xor U14517 (N_14517,N_8774,N_6184);
or U14518 (N_14518,N_6731,N_8115);
and U14519 (N_14519,N_8617,N_6818);
or U14520 (N_14520,N_8073,N_8946);
and U14521 (N_14521,N_6528,N_8038);
nor U14522 (N_14522,N_7474,N_9458);
nor U14523 (N_14523,N_5645,N_7146);
xor U14524 (N_14524,N_6113,N_8624);
or U14525 (N_14525,N_7759,N_8827);
or U14526 (N_14526,N_9558,N_7127);
xor U14527 (N_14527,N_7807,N_7825);
nand U14528 (N_14528,N_7040,N_8581);
nand U14529 (N_14529,N_6810,N_6681);
xnor U14530 (N_14530,N_8091,N_9697);
and U14531 (N_14531,N_7619,N_6062);
xnor U14532 (N_14532,N_5383,N_7646);
or U14533 (N_14533,N_6418,N_7794);
nand U14534 (N_14534,N_5541,N_5703);
or U14535 (N_14535,N_7652,N_8967);
and U14536 (N_14536,N_9488,N_9022);
nor U14537 (N_14537,N_8382,N_6548);
and U14538 (N_14538,N_7506,N_7329);
and U14539 (N_14539,N_6820,N_5149);
nand U14540 (N_14540,N_8376,N_8922);
or U14541 (N_14541,N_5219,N_9453);
or U14542 (N_14542,N_9785,N_7237);
nand U14543 (N_14543,N_6570,N_5474);
xnor U14544 (N_14544,N_6620,N_7161);
nor U14545 (N_14545,N_8403,N_6621);
or U14546 (N_14546,N_7896,N_5409);
xnor U14547 (N_14547,N_9842,N_5816);
nand U14548 (N_14548,N_8963,N_6223);
nand U14549 (N_14549,N_7259,N_9431);
nor U14550 (N_14550,N_9076,N_5013);
or U14551 (N_14551,N_8928,N_6598);
or U14552 (N_14552,N_5919,N_8739);
nand U14553 (N_14553,N_8190,N_5541);
nor U14554 (N_14554,N_9452,N_6413);
xor U14555 (N_14555,N_8673,N_6261);
xnor U14556 (N_14556,N_8897,N_7159);
or U14557 (N_14557,N_7210,N_5087);
and U14558 (N_14558,N_9627,N_6930);
nor U14559 (N_14559,N_8100,N_6151);
xnor U14560 (N_14560,N_9960,N_5013);
or U14561 (N_14561,N_5005,N_9368);
xnor U14562 (N_14562,N_5456,N_5906);
nand U14563 (N_14563,N_8430,N_8711);
nor U14564 (N_14564,N_7420,N_9412);
and U14565 (N_14565,N_7335,N_5916);
or U14566 (N_14566,N_6743,N_8070);
nand U14567 (N_14567,N_6706,N_5513);
nor U14568 (N_14568,N_9990,N_6716);
nor U14569 (N_14569,N_9628,N_5256);
xor U14570 (N_14570,N_8162,N_8209);
and U14571 (N_14571,N_6049,N_9308);
nor U14572 (N_14572,N_5623,N_8287);
and U14573 (N_14573,N_8522,N_9364);
nand U14574 (N_14574,N_6715,N_9831);
nor U14575 (N_14575,N_5247,N_5876);
nor U14576 (N_14576,N_8388,N_6223);
or U14577 (N_14577,N_6518,N_8476);
nor U14578 (N_14578,N_8595,N_5100);
xnor U14579 (N_14579,N_8185,N_6006);
or U14580 (N_14580,N_9313,N_8149);
nor U14581 (N_14581,N_9499,N_7422);
or U14582 (N_14582,N_9425,N_8102);
xor U14583 (N_14583,N_5819,N_7018);
xor U14584 (N_14584,N_7914,N_8399);
xnor U14585 (N_14585,N_8204,N_9567);
xnor U14586 (N_14586,N_6463,N_6175);
nor U14587 (N_14587,N_7215,N_8112);
nand U14588 (N_14588,N_8141,N_9215);
nand U14589 (N_14589,N_7185,N_7143);
nand U14590 (N_14590,N_7126,N_6462);
nor U14591 (N_14591,N_5299,N_5272);
nand U14592 (N_14592,N_6112,N_7090);
xor U14593 (N_14593,N_6436,N_8300);
nor U14594 (N_14594,N_7465,N_7253);
nor U14595 (N_14595,N_9142,N_8322);
nor U14596 (N_14596,N_7790,N_6736);
or U14597 (N_14597,N_8009,N_9867);
nand U14598 (N_14598,N_9528,N_9252);
nor U14599 (N_14599,N_5804,N_6123);
nand U14600 (N_14600,N_7624,N_8069);
xor U14601 (N_14601,N_8135,N_8004);
or U14602 (N_14602,N_7059,N_7546);
xor U14603 (N_14603,N_6450,N_5056);
and U14604 (N_14604,N_5025,N_8312);
or U14605 (N_14605,N_9945,N_6048);
nand U14606 (N_14606,N_8333,N_9088);
nand U14607 (N_14607,N_5753,N_9941);
and U14608 (N_14608,N_9956,N_6259);
or U14609 (N_14609,N_6096,N_7127);
or U14610 (N_14610,N_7397,N_9269);
or U14611 (N_14611,N_7982,N_6968);
nand U14612 (N_14612,N_7071,N_9740);
or U14613 (N_14613,N_6198,N_8701);
nand U14614 (N_14614,N_9908,N_8619);
or U14615 (N_14615,N_9246,N_7483);
nor U14616 (N_14616,N_9552,N_5192);
and U14617 (N_14617,N_5031,N_5762);
or U14618 (N_14618,N_6655,N_8831);
and U14619 (N_14619,N_8668,N_6248);
xnor U14620 (N_14620,N_9664,N_6476);
xnor U14621 (N_14621,N_8479,N_6386);
or U14622 (N_14622,N_9639,N_5014);
xor U14623 (N_14623,N_9998,N_6884);
nand U14624 (N_14624,N_5588,N_6852);
nand U14625 (N_14625,N_6839,N_7125);
nand U14626 (N_14626,N_6406,N_8417);
or U14627 (N_14627,N_6708,N_8059);
or U14628 (N_14628,N_9236,N_6016);
and U14629 (N_14629,N_7700,N_6852);
nor U14630 (N_14630,N_7608,N_5025);
nor U14631 (N_14631,N_9995,N_5429);
and U14632 (N_14632,N_5002,N_7034);
nor U14633 (N_14633,N_9789,N_9529);
and U14634 (N_14634,N_9707,N_8993);
nor U14635 (N_14635,N_9790,N_7972);
xnor U14636 (N_14636,N_5047,N_6430);
nand U14637 (N_14637,N_6846,N_7582);
and U14638 (N_14638,N_5830,N_8479);
xor U14639 (N_14639,N_5454,N_6603);
nor U14640 (N_14640,N_8813,N_6258);
xor U14641 (N_14641,N_7039,N_8528);
xor U14642 (N_14642,N_8730,N_8931);
xor U14643 (N_14643,N_5291,N_6807);
or U14644 (N_14644,N_8932,N_6005);
and U14645 (N_14645,N_6623,N_5328);
xor U14646 (N_14646,N_8212,N_5045);
or U14647 (N_14647,N_8296,N_6003);
nand U14648 (N_14648,N_9118,N_8384);
or U14649 (N_14649,N_9134,N_5374);
nand U14650 (N_14650,N_8719,N_5047);
or U14651 (N_14651,N_6955,N_9662);
nand U14652 (N_14652,N_7235,N_5372);
or U14653 (N_14653,N_5611,N_5598);
xor U14654 (N_14654,N_8929,N_7277);
nor U14655 (N_14655,N_9731,N_7823);
xor U14656 (N_14656,N_5878,N_7103);
and U14657 (N_14657,N_5975,N_8655);
nor U14658 (N_14658,N_7181,N_7085);
or U14659 (N_14659,N_8335,N_6646);
nor U14660 (N_14660,N_8541,N_7017);
nand U14661 (N_14661,N_7781,N_5336);
and U14662 (N_14662,N_8802,N_6989);
xnor U14663 (N_14663,N_5645,N_5855);
nor U14664 (N_14664,N_9543,N_5194);
and U14665 (N_14665,N_7957,N_9984);
nor U14666 (N_14666,N_5247,N_8224);
and U14667 (N_14667,N_6327,N_8589);
or U14668 (N_14668,N_8443,N_8575);
xor U14669 (N_14669,N_6423,N_7832);
xnor U14670 (N_14670,N_9707,N_9198);
nand U14671 (N_14671,N_6702,N_9461);
xnor U14672 (N_14672,N_9145,N_9013);
xor U14673 (N_14673,N_7895,N_9239);
xor U14674 (N_14674,N_6790,N_9256);
or U14675 (N_14675,N_6401,N_7147);
and U14676 (N_14676,N_7258,N_5831);
and U14677 (N_14677,N_7330,N_9821);
nor U14678 (N_14678,N_9815,N_6443);
xor U14679 (N_14679,N_9631,N_7123);
and U14680 (N_14680,N_9926,N_8525);
and U14681 (N_14681,N_7972,N_7642);
nor U14682 (N_14682,N_7687,N_6254);
or U14683 (N_14683,N_5866,N_9552);
or U14684 (N_14684,N_8681,N_8253);
or U14685 (N_14685,N_9981,N_7439);
nand U14686 (N_14686,N_5435,N_5722);
nand U14687 (N_14687,N_9706,N_6932);
nor U14688 (N_14688,N_5112,N_9817);
or U14689 (N_14689,N_8759,N_8455);
xnor U14690 (N_14690,N_9137,N_6113);
or U14691 (N_14691,N_9256,N_6628);
xnor U14692 (N_14692,N_6764,N_9501);
xnor U14693 (N_14693,N_7724,N_8829);
nor U14694 (N_14694,N_6421,N_5266);
nor U14695 (N_14695,N_7804,N_6747);
nor U14696 (N_14696,N_8797,N_5829);
nor U14697 (N_14697,N_9588,N_7723);
xor U14698 (N_14698,N_5355,N_7464);
nand U14699 (N_14699,N_7905,N_7436);
nand U14700 (N_14700,N_7348,N_7272);
nor U14701 (N_14701,N_5779,N_7986);
nor U14702 (N_14702,N_8526,N_5894);
nand U14703 (N_14703,N_5177,N_7429);
nor U14704 (N_14704,N_9391,N_5034);
or U14705 (N_14705,N_5070,N_5770);
xnor U14706 (N_14706,N_6404,N_6926);
nand U14707 (N_14707,N_9610,N_7453);
nand U14708 (N_14708,N_7373,N_8523);
or U14709 (N_14709,N_7765,N_9309);
nand U14710 (N_14710,N_8602,N_5450);
nand U14711 (N_14711,N_9103,N_6096);
nor U14712 (N_14712,N_9506,N_7111);
xnor U14713 (N_14713,N_9231,N_6927);
nand U14714 (N_14714,N_8106,N_8471);
xor U14715 (N_14715,N_9787,N_8117);
nand U14716 (N_14716,N_9946,N_7980);
or U14717 (N_14717,N_7278,N_9722);
and U14718 (N_14718,N_8037,N_6388);
or U14719 (N_14719,N_5177,N_8163);
nor U14720 (N_14720,N_5142,N_7113);
nor U14721 (N_14721,N_7688,N_7486);
xor U14722 (N_14722,N_5606,N_6365);
nor U14723 (N_14723,N_8493,N_9018);
or U14724 (N_14724,N_6757,N_8075);
nor U14725 (N_14725,N_7897,N_9138);
nand U14726 (N_14726,N_5611,N_9615);
xnor U14727 (N_14727,N_8579,N_7398);
nand U14728 (N_14728,N_9443,N_7413);
xnor U14729 (N_14729,N_7685,N_8601);
nand U14730 (N_14730,N_6161,N_8187);
nor U14731 (N_14731,N_7325,N_7549);
or U14732 (N_14732,N_9280,N_9834);
nor U14733 (N_14733,N_6791,N_9635);
nand U14734 (N_14734,N_9918,N_5158);
or U14735 (N_14735,N_7808,N_6973);
nand U14736 (N_14736,N_5852,N_7594);
and U14737 (N_14737,N_5516,N_9142);
xnor U14738 (N_14738,N_7639,N_8987);
or U14739 (N_14739,N_8274,N_9308);
and U14740 (N_14740,N_6196,N_8419);
and U14741 (N_14741,N_7858,N_9913);
and U14742 (N_14742,N_8597,N_9475);
or U14743 (N_14743,N_9322,N_6383);
nand U14744 (N_14744,N_5064,N_8702);
or U14745 (N_14745,N_5467,N_9296);
and U14746 (N_14746,N_9527,N_7295);
xor U14747 (N_14747,N_7797,N_5229);
xnor U14748 (N_14748,N_9782,N_7671);
or U14749 (N_14749,N_6939,N_8835);
nand U14750 (N_14750,N_8815,N_5140);
nand U14751 (N_14751,N_9651,N_8548);
or U14752 (N_14752,N_9643,N_7837);
or U14753 (N_14753,N_8291,N_6069);
nor U14754 (N_14754,N_5881,N_5648);
nor U14755 (N_14755,N_5988,N_8963);
nand U14756 (N_14756,N_6440,N_5171);
and U14757 (N_14757,N_5913,N_8634);
or U14758 (N_14758,N_7762,N_8343);
nor U14759 (N_14759,N_7554,N_9467);
and U14760 (N_14760,N_8654,N_9693);
nand U14761 (N_14761,N_6742,N_8606);
nand U14762 (N_14762,N_5423,N_5836);
xnor U14763 (N_14763,N_8318,N_5945);
or U14764 (N_14764,N_7155,N_8958);
and U14765 (N_14765,N_7674,N_8870);
xnor U14766 (N_14766,N_5320,N_5110);
or U14767 (N_14767,N_8651,N_6097);
or U14768 (N_14768,N_9929,N_7714);
and U14769 (N_14769,N_7109,N_6676);
xor U14770 (N_14770,N_6322,N_9795);
nor U14771 (N_14771,N_5295,N_9300);
nor U14772 (N_14772,N_8516,N_7482);
or U14773 (N_14773,N_5115,N_9736);
xor U14774 (N_14774,N_8288,N_7458);
xor U14775 (N_14775,N_8075,N_7277);
xnor U14776 (N_14776,N_9486,N_7675);
nand U14777 (N_14777,N_6132,N_7738);
or U14778 (N_14778,N_8492,N_6566);
nand U14779 (N_14779,N_6933,N_9731);
nand U14780 (N_14780,N_9620,N_7103);
nor U14781 (N_14781,N_7559,N_9999);
nand U14782 (N_14782,N_6181,N_8568);
xnor U14783 (N_14783,N_5463,N_8049);
xor U14784 (N_14784,N_7915,N_8993);
or U14785 (N_14785,N_7309,N_6426);
nor U14786 (N_14786,N_6379,N_5892);
nand U14787 (N_14787,N_6383,N_7269);
xnor U14788 (N_14788,N_6668,N_7414);
nor U14789 (N_14789,N_5952,N_6726);
xnor U14790 (N_14790,N_5704,N_7348);
or U14791 (N_14791,N_5674,N_8617);
and U14792 (N_14792,N_9589,N_9837);
nand U14793 (N_14793,N_5152,N_7958);
nor U14794 (N_14794,N_7974,N_7718);
or U14795 (N_14795,N_8318,N_6314);
nor U14796 (N_14796,N_9287,N_5717);
nand U14797 (N_14797,N_8417,N_5488);
and U14798 (N_14798,N_6057,N_8776);
xnor U14799 (N_14799,N_6580,N_8965);
xor U14800 (N_14800,N_6105,N_6337);
and U14801 (N_14801,N_8359,N_7272);
and U14802 (N_14802,N_8992,N_8662);
and U14803 (N_14803,N_5709,N_6863);
xor U14804 (N_14804,N_7780,N_8919);
xnor U14805 (N_14805,N_9918,N_5790);
nor U14806 (N_14806,N_6439,N_5915);
nor U14807 (N_14807,N_6386,N_9743);
and U14808 (N_14808,N_5405,N_8196);
or U14809 (N_14809,N_7581,N_6562);
or U14810 (N_14810,N_6641,N_6557);
or U14811 (N_14811,N_9725,N_6044);
nand U14812 (N_14812,N_6877,N_7458);
xor U14813 (N_14813,N_9338,N_8126);
and U14814 (N_14814,N_7061,N_9191);
nand U14815 (N_14815,N_9239,N_7468);
nand U14816 (N_14816,N_5941,N_6677);
nor U14817 (N_14817,N_5161,N_6032);
nor U14818 (N_14818,N_7601,N_8069);
nand U14819 (N_14819,N_9542,N_8313);
and U14820 (N_14820,N_7634,N_5489);
nor U14821 (N_14821,N_9313,N_6129);
or U14822 (N_14822,N_9021,N_8185);
nor U14823 (N_14823,N_8774,N_9611);
or U14824 (N_14824,N_7215,N_9863);
nand U14825 (N_14825,N_9851,N_7421);
and U14826 (N_14826,N_7147,N_6700);
xor U14827 (N_14827,N_7583,N_9811);
or U14828 (N_14828,N_9126,N_8491);
and U14829 (N_14829,N_8076,N_8783);
or U14830 (N_14830,N_8913,N_5306);
or U14831 (N_14831,N_6948,N_6957);
and U14832 (N_14832,N_5461,N_6837);
nor U14833 (N_14833,N_8693,N_6853);
nor U14834 (N_14834,N_7027,N_7600);
nor U14835 (N_14835,N_8343,N_8308);
nor U14836 (N_14836,N_6401,N_7562);
or U14837 (N_14837,N_5809,N_9890);
xnor U14838 (N_14838,N_9990,N_8725);
nor U14839 (N_14839,N_8688,N_5990);
xor U14840 (N_14840,N_8325,N_7207);
or U14841 (N_14841,N_7396,N_9228);
or U14842 (N_14842,N_5077,N_6262);
and U14843 (N_14843,N_8908,N_6803);
xnor U14844 (N_14844,N_7526,N_9844);
and U14845 (N_14845,N_8095,N_9646);
nor U14846 (N_14846,N_9224,N_7581);
xnor U14847 (N_14847,N_9572,N_7880);
nand U14848 (N_14848,N_7193,N_8975);
nand U14849 (N_14849,N_6306,N_7957);
nor U14850 (N_14850,N_5429,N_7534);
and U14851 (N_14851,N_5707,N_8465);
nor U14852 (N_14852,N_7420,N_6190);
xor U14853 (N_14853,N_5781,N_5335);
xor U14854 (N_14854,N_8537,N_7611);
nand U14855 (N_14855,N_6946,N_7424);
xnor U14856 (N_14856,N_6849,N_7047);
nand U14857 (N_14857,N_6690,N_9045);
nand U14858 (N_14858,N_9901,N_9797);
nor U14859 (N_14859,N_7898,N_9588);
nor U14860 (N_14860,N_5852,N_8936);
or U14861 (N_14861,N_8566,N_9309);
or U14862 (N_14862,N_6332,N_8132);
xnor U14863 (N_14863,N_5014,N_6741);
or U14864 (N_14864,N_5405,N_6255);
and U14865 (N_14865,N_9857,N_9294);
nor U14866 (N_14866,N_6922,N_9697);
or U14867 (N_14867,N_6755,N_9605);
xor U14868 (N_14868,N_9852,N_9982);
and U14869 (N_14869,N_8002,N_9906);
nor U14870 (N_14870,N_5258,N_5754);
nor U14871 (N_14871,N_7661,N_8617);
xnor U14872 (N_14872,N_6082,N_9608);
nand U14873 (N_14873,N_7119,N_7927);
nor U14874 (N_14874,N_8763,N_5365);
or U14875 (N_14875,N_8624,N_9267);
and U14876 (N_14876,N_5588,N_7419);
nand U14877 (N_14877,N_7258,N_5660);
or U14878 (N_14878,N_9520,N_6655);
or U14879 (N_14879,N_7889,N_5256);
xor U14880 (N_14880,N_8652,N_5611);
and U14881 (N_14881,N_6503,N_7053);
and U14882 (N_14882,N_7023,N_9449);
and U14883 (N_14883,N_9861,N_8754);
nand U14884 (N_14884,N_7461,N_7989);
xor U14885 (N_14885,N_9701,N_6151);
nand U14886 (N_14886,N_8243,N_6779);
nor U14887 (N_14887,N_5475,N_8544);
nor U14888 (N_14888,N_6886,N_8237);
nand U14889 (N_14889,N_5943,N_6616);
nand U14890 (N_14890,N_5621,N_8062);
xnor U14891 (N_14891,N_6826,N_5079);
and U14892 (N_14892,N_9357,N_7642);
nor U14893 (N_14893,N_8166,N_8498);
xnor U14894 (N_14894,N_9679,N_7650);
xnor U14895 (N_14895,N_5515,N_9417);
nor U14896 (N_14896,N_6683,N_8137);
xnor U14897 (N_14897,N_9146,N_7482);
nand U14898 (N_14898,N_9767,N_9469);
or U14899 (N_14899,N_8079,N_9726);
or U14900 (N_14900,N_7067,N_8252);
xor U14901 (N_14901,N_7615,N_5191);
or U14902 (N_14902,N_9267,N_9478);
xor U14903 (N_14903,N_8207,N_8506);
and U14904 (N_14904,N_5716,N_6082);
nor U14905 (N_14905,N_9377,N_6656);
nor U14906 (N_14906,N_6798,N_8780);
xor U14907 (N_14907,N_8472,N_9041);
nor U14908 (N_14908,N_5911,N_8696);
and U14909 (N_14909,N_6533,N_9794);
xor U14910 (N_14910,N_8733,N_5417);
or U14911 (N_14911,N_7244,N_9151);
nand U14912 (N_14912,N_5509,N_6979);
nand U14913 (N_14913,N_8685,N_6269);
or U14914 (N_14914,N_7099,N_7313);
and U14915 (N_14915,N_9053,N_5913);
or U14916 (N_14916,N_7992,N_8337);
nand U14917 (N_14917,N_7641,N_5516);
nand U14918 (N_14918,N_6991,N_5985);
and U14919 (N_14919,N_7666,N_5001);
or U14920 (N_14920,N_5964,N_5501);
nand U14921 (N_14921,N_5801,N_7691);
xnor U14922 (N_14922,N_9473,N_5059);
or U14923 (N_14923,N_8832,N_9482);
and U14924 (N_14924,N_8914,N_6580);
or U14925 (N_14925,N_8201,N_7363);
nor U14926 (N_14926,N_8498,N_6068);
nor U14927 (N_14927,N_5096,N_8920);
or U14928 (N_14928,N_5485,N_9713);
xnor U14929 (N_14929,N_7188,N_8156);
and U14930 (N_14930,N_6549,N_7978);
nand U14931 (N_14931,N_5672,N_6280);
or U14932 (N_14932,N_5741,N_5783);
and U14933 (N_14933,N_9493,N_8025);
nand U14934 (N_14934,N_9370,N_6502);
or U14935 (N_14935,N_7001,N_7297);
and U14936 (N_14936,N_5345,N_7992);
xor U14937 (N_14937,N_8853,N_7292);
and U14938 (N_14938,N_8256,N_8839);
and U14939 (N_14939,N_6212,N_7372);
or U14940 (N_14940,N_7390,N_6380);
or U14941 (N_14941,N_6823,N_5683);
xor U14942 (N_14942,N_6291,N_9754);
and U14943 (N_14943,N_7796,N_5691);
or U14944 (N_14944,N_9647,N_7631);
or U14945 (N_14945,N_9224,N_8216);
or U14946 (N_14946,N_8708,N_8683);
nand U14947 (N_14947,N_6957,N_6075);
xor U14948 (N_14948,N_9010,N_7377);
xnor U14949 (N_14949,N_7244,N_8144);
and U14950 (N_14950,N_6606,N_8503);
and U14951 (N_14951,N_9341,N_5813);
or U14952 (N_14952,N_5763,N_5433);
xor U14953 (N_14953,N_7411,N_6572);
xor U14954 (N_14954,N_5858,N_9655);
nor U14955 (N_14955,N_5705,N_8761);
xnor U14956 (N_14956,N_9651,N_7462);
nand U14957 (N_14957,N_9781,N_6528);
or U14958 (N_14958,N_8901,N_8187);
xnor U14959 (N_14959,N_7881,N_7972);
or U14960 (N_14960,N_7198,N_7264);
or U14961 (N_14961,N_6041,N_6938);
and U14962 (N_14962,N_9138,N_8994);
nor U14963 (N_14963,N_5861,N_7817);
nand U14964 (N_14964,N_7952,N_9071);
or U14965 (N_14965,N_6963,N_5126);
and U14966 (N_14966,N_6163,N_9567);
nand U14967 (N_14967,N_9324,N_8479);
and U14968 (N_14968,N_7729,N_5351);
xnor U14969 (N_14969,N_7950,N_7205);
and U14970 (N_14970,N_8423,N_7687);
nand U14971 (N_14971,N_9799,N_6689);
and U14972 (N_14972,N_7766,N_6985);
and U14973 (N_14973,N_7552,N_7347);
or U14974 (N_14974,N_8841,N_9864);
nor U14975 (N_14975,N_6445,N_9889);
nor U14976 (N_14976,N_9596,N_6812);
nor U14977 (N_14977,N_9915,N_7566);
nand U14978 (N_14978,N_9670,N_7106);
nand U14979 (N_14979,N_7348,N_6824);
or U14980 (N_14980,N_9915,N_9634);
nand U14981 (N_14981,N_9491,N_8662);
or U14982 (N_14982,N_9177,N_5715);
nand U14983 (N_14983,N_9534,N_5842);
and U14984 (N_14984,N_9693,N_8399);
nor U14985 (N_14985,N_8365,N_7339);
or U14986 (N_14986,N_6734,N_9399);
or U14987 (N_14987,N_6206,N_9866);
and U14988 (N_14988,N_7822,N_5409);
xnor U14989 (N_14989,N_6136,N_6227);
nor U14990 (N_14990,N_8991,N_7509);
or U14991 (N_14991,N_7075,N_5468);
nor U14992 (N_14992,N_6985,N_7854);
nor U14993 (N_14993,N_9866,N_8624);
nor U14994 (N_14994,N_7485,N_7531);
nand U14995 (N_14995,N_8436,N_5516);
nor U14996 (N_14996,N_8081,N_5302);
and U14997 (N_14997,N_9847,N_5646);
or U14998 (N_14998,N_6937,N_7266);
xor U14999 (N_14999,N_8435,N_6008);
xnor U15000 (N_15000,N_12788,N_14150);
nor U15001 (N_15001,N_10069,N_13372);
nand U15002 (N_15002,N_10033,N_13830);
nand U15003 (N_15003,N_12896,N_10180);
nand U15004 (N_15004,N_13245,N_11525);
or U15005 (N_15005,N_11251,N_10052);
xor U15006 (N_15006,N_11383,N_12488);
and U15007 (N_15007,N_10325,N_12376);
and U15008 (N_15008,N_14996,N_12502);
nand U15009 (N_15009,N_13144,N_13772);
nor U15010 (N_15010,N_13623,N_11536);
and U15011 (N_15011,N_13053,N_12406);
nor U15012 (N_15012,N_13803,N_14367);
xnor U15013 (N_15013,N_14222,N_12057);
or U15014 (N_15014,N_12589,N_11656);
or U15015 (N_15015,N_10875,N_14346);
or U15016 (N_15016,N_10584,N_13018);
nand U15017 (N_15017,N_11569,N_14784);
nand U15018 (N_15018,N_12869,N_14662);
nor U15019 (N_15019,N_12775,N_13233);
and U15020 (N_15020,N_12021,N_14431);
nand U15021 (N_15021,N_13371,N_12316);
and U15022 (N_15022,N_10400,N_10267);
nor U15023 (N_15023,N_13346,N_12417);
xor U15024 (N_15024,N_12452,N_14679);
or U15025 (N_15025,N_11979,N_13883);
nor U15026 (N_15026,N_11909,N_10038);
nand U15027 (N_15027,N_14539,N_13219);
and U15028 (N_15028,N_11688,N_14142);
xnor U15029 (N_15029,N_10906,N_10174);
nor U15030 (N_15030,N_10064,N_14554);
or U15031 (N_15031,N_14318,N_12912);
nor U15032 (N_15032,N_12301,N_11555);
nor U15033 (N_15033,N_11967,N_14430);
or U15034 (N_15034,N_12424,N_11067);
xnor U15035 (N_15035,N_13939,N_12458);
nand U15036 (N_15036,N_11476,N_11778);
nand U15037 (N_15037,N_14719,N_12296);
or U15038 (N_15038,N_13596,N_11657);
xor U15039 (N_15039,N_12430,N_12249);
or U15040 (N_15040,N_14130,N_14504);
nor U15041 (N_15041,N_10465,N_10931);
nor U15042 (N_15042,N_11617,N_12046);
or U15043 (N_15043,N_13204,N_14588);
nor U15044 (N_15044,N_10153,N_14332);
or U15045 (N_15045,N_13866,N_14102);
and U15046 (N_15046,N_14824,N_11256);
xnor U15047 (N_15047,N_11660,N_14201);
xor U15048 (N_15048,N_12169,N_11087);
xor U15049 (N_15049,N_10573,N_10547);
or U15050 (N_15050,N_14811,N_14803);
nor U15051 (N_15051,N_11043,N_11771);
nand U15052 (N_15052,N_11182,N_10973);
or U15053 (N_15053,N_13446,N_12489);
nor U15054 (N_15054,N_14747,N_12996);
and U15055 (N_15055,N_12661,N_10299);
and U15056 (N_15056,N_14184,N_12528);
nand U15057 (N_15057,N_14756,N_13416);
nand U15058 (N_15058,N_12813,N_11744);
and U15059 (N_15059,N_10082,N_12780);
and U15060 (N_15060,N_13466,N_10874);
nor U15061 (N_15061,N_13438,N_12393);
or U15062 (N_15062,N_11009,N_13203);
or U15063 (N_15063,N_13636,N_13960);
nand U15064 (N_15064,N_10125,N_10716);
nor U15065 (N_15065,N_14211,N_10763);
or U15066 (N_15066,N_12960,N_13294);
xor U15067 (N_15067,N_10133,N_10755);
xor U15068 (N_15068,N_13914,N_13609);
xor U15069 (N_15069,N_14113,N_14037);
nand U15070 (N_15070,N_14826,N_12673);
and U15071 (N_15071,N_11540,N_12124);
or U15072 (N_15072,N_13603,N_14191);
nand U15073 (N_15073,N_14185,N_12276);
and U15074 (N_15074,N_11075,N_12320);
nor U15075 (N_15075,N_10712,N_11102);
xor U15076 (N_15076,N_11783,N_11456);
and U15077 (N_15077,N_14638,N_11554);
nor U15078 (N_15078,N_14182,N_10621);
xnor U15079 (N_15079,N_13793,N_13486);
xor U15080 (N_15080,N_11761,N_12705);
nor U15081 (N_15081,N_13526,N_14505);
or U15082 (N_15082,N_14010,N_14770);
and U15083 (N_15083,N_11840,N_14343);
and U15084 (N_15084,N_13520,N_13248);
xnor U15085 (N_15085,N_14393,N_12179);
or U15086 (N_15086,N_10076,N_12829);
nor U15087 (N_15087,N_13759,N_10784);
or U15088 (N_15088,N_13176,N_13473);
nand U15089 (N_15089,N_11079,N_14816);
nand U15090 (N_15090,N_12596,N_11244);
nand U15091 (N_15091,N_12364,N_14727);
and U15092 (N_15092,N_13207,N_13511);
nor U15093 (N_15093,N_11213,N_13317);
or U15094 (N_15094,N_10120,N_12041);
xnor U15095 (N_15095,N_10667,N_11833);
nand U15096 (N_15096,N_14058,N_11805);
nand U15097 (N_15097,N_14020,N_11943);
xor U15098 (N_15098,N_13396,N_13357);
and U15099 (N_15099,N_12107,N_13071);
and U15100 (N_15100,N_10121,N_13592);
nor U15101 (N_15101,N_14138,N_14992);
nand U15102 (N_15102,N_10756,N_11799);
xor U15103 (N_15103,N_14087,N_13938);
xnor U15104 (N_15104,N_13318,N_12837);
xnor U15105 (N_15105,N_13354,N_14589);
nand U15106 (N_15106,N_10708,N_10697);
nand U15107 (N_15107,N_12740,N_13987);
xor U15108 (N_15108,N_13404,N_11626);
and U15109 (N_15109,N_10955,N_11165);
or U15110 (N_15110,N_10163,N_13135);
and U15111 (N_15111,N_10845,N_11685);
nand U15112 (N_15112,N_12300,N_10889);
and U15113 (N_15113,N_10105,N_13947);
xor U15114 (N_15114,N_11049,N_12663);
xnor U15115 (N_15115,N_11792,N_11291);
or U15116 (N_15116,N_12384,N_10006);
xnor U15117 (N_15117,N_13693,N_14698);
xor U15118 (N_15118,N_11320,N_12302);
and U15119 (N_15119,N_12470,N_13213);
nor U15120 (N_15120,N_10903,N_10855);
nand U15121 (N_15121,N_10783,N_12591);
nor U15122 (N_15122,N_12793,N_13591);
nor U15123 (N_15123,N_14750,N_11773);
xor U15124 (N_15124,N_12381,N_11463);
and U15125 (N_15125,N_14487,N_11366);
or U15126 (N_15126,N_11263,N_13068);
and U15127 (N_15127,N_12728,N_10202);
xnor U15128 (N_15128,N_14533,N_12219);
nand U15129 (N_15129,N_12997,N_13870);
or U15130 (N_15130,N_12892,N_10691);
or U15131 (N_15131,N_13661,N_14524);
nand U15132 (N_15132,N_11679,N_11516);
and U15133 (N_15133,N_13033,N_11851);
nor U15134 (N_15134,N_10479,N_11574);
nand U15135 (N_15135,N_11264,N_14891);
or U15136 (N_15136,N_14534,N_14099);
xnor U15137 (N_15137,N_10405,N_10637);
or U15138 (N_15138,N_12361,N_13170);
nor U15139 (N_15139,N_12394,N_11502);
or U15140 (N_15140,N_12861,N_14796);
or U15141 (N_15141,N_10692,N_13902);
nor U15142 (N_15142,N_11892,N_14492);
or U15143 (N_15143,N_10509,N_10902);
nor U15144 (N_15144,N_10936,N_13680);
and U15145 (N_15145,N_11363,N_10251);
nand U15146 (N_15146,N_12943,N_14563);
nor U15147 (N_15147,N_13600,N_14093);
nor U15148 (N_15148,N_13659,N_10575);
nor U15149 (N_15149,N_10438,N_13403);
xor U15150 (N_15150,N_11396,N_13199);
nor U15151 (N_15151,N_12322,N_13295);
nand U15152 (N_15152,N_13079,N_10217);
and U15153 (N_15153,N_10188,N_12333);
nor U15154 (N_15154,N_10235,N_10680);
xnor U15155 (N_15155,N_14388,N_13013);
nand U15156 (N_15156,N_11083,N_12423);
nor U15157 (N_15157,N_10071,N_13517);
nor U15158 (N_15158,N_13804,N_10036);
nor U15159 (N_15159,N_13181,N_11785);
and U15160 (N_15160,N_11157,N_14830);
nor U15161 (N_15161,N_11905,N_14241);
nand U15162 (N_15162,N_13730,N_12863);
nor U15163 (N_15163,N_12592,N_10950);
or U15164 (N_15164,N_13221,N_12771);
and U15165 (N_15165,N_14836,N_14468);
nor U15166 (N_15166,N_12583,N_12483);
nand U15167 (N_15167,N_13386,N_14415);
or U15168 (N_15168,N_10834,N_10679);
xnor U15169 (N_15169,N_11277,N_10425);
nand U15170 (N_15170,N_10754,N_14014);
and U15171 (N_15171,N_12557,N_10363);
and U15172 (N_15172,N_10720,N_10238);
or U15173 (N_15173,N_12641,N_12081);
xnor U15174 (N_15174,N_10780,N_13877);
and U15175 (N_15175,N_11381,N_12188);
nor U15176 (N_15176,N_14118,N_10682);
or U15177 (N_15177,N_14190,N_12246);
and U15178 (N_15178,N_13224,N_12182);
nor U15179 (N_15179,N_11346,N_13822);
nand U15180 (N_15180,N_12429,N_10740);
nand U15181 (N_15181,N_11241,N_11404);
and U15182 (N_15182,N_11261,N_14527);
nand U15183 (N_15183,N_11423,N_11269);
nor U15184 (N_15184,N_10256,N_10811);
and U15185 (N_15185,N_10896,N_12737);
and U15186 (N_15186,N_10976,N_14954);
and U15187 (N_15187,N_10778,N_12602);
nor U15188 (N_15188,N_10618,N_10767);
nand U15189 (N_15189,N_11254,N_12253);
nand U15190 (N_15190,N_11776,N_13900);
xnor U15191 (N_15191,N_12251,N_12939);
and U15192 (N_15192,N_10693,N_11658);
or U15193 (N_15193,N_12030,N_11941);
or U15194 (N_15194,N_10303,N_11844);
xor U15195 (N_15195,N_13749,N_10961);
and U15196 (N_15196,N_10476,N_12946);
or U15197 (N_15197,N_10883,N_14316);
nand U15198 (N_15198,N_14667,N_10964);
and U15199 (N_15199,N_12297,N_11561);
xor U15200 (N_15200,N_10246,N_13310);
or U15201 (N_15201,N_13143,N_10499);
xor U15202 (N_15202,N_10869,N_14874);
xor U15203 (N_15203,N_10321,N_11141);
nor U15204 (N_15204,N_11565,N_12797);
xnor U15205 (N_15205,N_12212,N_14204);
xnor U15206 (N_15206,N_13745,N_11861);
or U15207 (N_15207,N_13364,N_11206);
xor U15208 (N_15208,N_14506,N_13392);
or U15209 (N_15209,N_13918,N_14322);
nand U15210 (N_15210,N_10164,N_14351);
nand U15211 (N_15211,N_14977,N_13202);
or U15212 (N_15212,N_10422,N_10047);
nor U15213 (N_15213,N_10137,N_13530);
nand U15214 (N_15214,N_14270,N_11188);
and U15215 (N_15215,N_13714,N_11236);
xor U15216 (N_15216,N_13559,N_11559);
and U15217 (N_15217,N_10797,N_13996);
nand U15218 (N_15218,N_12126,N_11202);
nand U15219 (N_15219,N_13655,N_12926);
or U15220 (N_15220,N_12461,N_13195);
and U15221 (N_15221,N_13454,N_10265);
xor U15222 (N_15222,N_14911,N_14976);
nand U15223 (N_15223,N_11237,N_10209);
xor U15224 (N_15224,N_11191,N_12530);
nand U15225 (N_15225,N_12236,N_10021);
nor U15226 (N_15226,N_11537,N_10404);
nor U15227 (N_15227,N_13741,N_13103);
nand U15228 (N_15228,N_12418,N_11640);
nor U15229 (N_15229,N_10612,N_10140);
xnor U15230 (N_15230,N_12239,N_10090);
nand U15231 (N_15231,N_11281,N_13919);
and U15232 (N_15232,N_13982,N_11039);
nand U15233 (N_15233,N_13828,N_10398);
nand U15234 (N_15234,N_10409,N_12113);
and U15235 (N_15235,N_13905,N_14942);
and U15236 (N_15236,N_14602,N_13481);
xnor U15237 (N_15237,N_10428,N_10451);
or U15238 (N_15238,N_14434,N_11276);
and U15239 (N_15239,N_10578,N_13235);
xnor U15240 (N_15240,N_14147,N_12642);
or U15241 (N_15241,N_11508,N_14407);
or U15242 (N_15242,N_13840,N_12637);
nor U15243 (N_15243,N_14512,N_10887);
xor U15244 (N_15244,N_11158,N_11221);
and U15245 (N_15245,N_14908,N_11216);
nor U15246 (N_15246,N_13732,N_10450);
nand U15247 (N_15247,N_13425,N_14511);
nand U15248 (N_15248,N_12687,N_12761);
xnor U15249 (N_15249,N_11295,N_11161);
nor U15250 (N_15250,N_11430,N_13039);
xnor U15251 (N_15251,N_12688,N_14286);
or U15252 (N_15252,N_14383,N_14484);
and U15253 (N_15253,N_12338,N_12866);
or U15254 (N_15254,N_14497,N_10282);
or U15255 (N_15255,N_12501,N_13588);
nand U15256 (N_15256,N_14298,N_11332);
xnor U15257 (N_15257,N_13196,N_13338);
nor U15258 (N_15258,N_13073,N_12975);
or U15259 (N_15259,N_12092,N_12180);
or U15260 (N_15260,N_13509,N_14002);
or U15261 (N_15261,N_14692,N_12938);
nor U15262 (N_15262,N_12103,N_11451);
nor U15263 (N_15263,N_14793,N_14724);
or U15264 (N_15264,N_13391,N_10255);
or U15265 (N_15265,N_12617,N_13412);
nand U15266 (N_15266,N_10714,N_12587);
nor U15267 (N_15267,N_12466,N_12879);
or U15268 (N_15268,N_13956,N_13989);
nand U15269 (N_15269,N_14556,N_12324);
and U15270 (N_15270,N_12094,N_10628);
nand U15271 (N_15271,N_12250,N_12507);
or U15272 (N_15272,N_14257,N_13689);
and U15273 (N_15273,N_13555,N_14689);
or U15274 (N_15274,N_14305,N_11808);
nand U15275 (N_15275,N_11105,N_11866);
and U15276 (N_15276,N_10656,N_13529);
and U15277 (N_15277,N_14810,N_14635);
and U15278 (N_15278,N_12010,N_13988);
nor U15279 (N_15279,N_11974,N_12901);
and U15280 (N_15280,N_10603,N_11839);
nor U15281 (N_15281,N_14210,N_11318);
xor U15282 (N_15282,N_11448,N_14799);
nand U15283 (N_15283,N_10305,N_12726);
or U15284 (N_15284,N_11961,N_13893);
xnor U15285 (N_15285,N_10349,N_11192);
nand U15286 (N_15286,N_13834,N_13615);
nor U15287 (N_15287,N_14256,N_13972);
and U15288 (N_15288,N_10135,N_12791);
nor U15289 (N_15289,N_13777,N_13970);
xor U15290 (N_15290,N_13270,N_10934);
xnor U15291 (N_15291,N_10542,N_13604);
and U15292 (N_15292,N_10226,N_13858);
xor U15293 (N_15293,N_12841,N_14986);
or U15294 (N_15294,N_12991,N_10608);
nor U15295 (N_15295,N_12291,N_14938);
xor U15296 (N_15296,N_12881,N_11872);
xor U15297 (N_15297,N_11946,N_12431);
xnor U15298 (N_15298,N_10704,N_13131);
xor U15299 (N_15299,N_14955,N_14880);
xnor U15300 (N_15300,N_11735,N_14139);
nor U15301 (N_15301,N_11817,N_10207);
nand U15302 (N_15302,N_10622,N_14043);
xor U15303 (N_15303,N_11501,N_10475);
nand U15304 (N_15304,N_10978,N_13393);
or U15305 (N_15305,N_12303,N_12905);
nor U15306 (N_15306,N_10841,N_12538);
nand U15307 (N_15307,N_13080,N_10706);
and U15308 (N_15308,N_13798,N_12803);
and U15309 (N_15309,N_12290,N_12950);
nor U15310 (N_15310,N_13581,N_14086);
or U15311 (N_15311,N_11696,N_12197);
nand U15312 (N_15312,N_13617,N_12590);
xnor U15313 (N_15313,N_11958,N_11870);
nor U15314 (N_15314,N_12897,N_12511);
and U15315 (N_15315,N_11292,N_10387);
xnor U15316 (N_15316,N_10910,N_10825);
xor U15317 (N_15317,N_11354,N_10997);
nand U15318 (N_15318,N_14744,N_12422);
or U15319 (N_15319,N_10962,N_11010);
and U15320 (N_15320,N_12478,N_14514);
and U15321 (N_15321,N_12559,N_10766);
or U15322 (N_15322,N_10624,N_12217);
nor U15323 (N_15323,N_14605,N_11891);
and U15324 (N_15324,N_11217,N_11889);
or U15325 (N_15325,N_12809,N_11527);
or U15326 (N_15326,N_14075,N_12156);
xor U15327 (N_15327,N_13247,N_12555);
and U15328 (N_15328,N_12521,N_14910);
nand U15329 (N_15329,N_13713,N_13369);
nand U15330 (N_15330,N_10132,N_11123);
or U15331 (N_15331,N_14861,N_12252);
xnor U15332 (N_15332,N_10331,N_13983);
nor U15333 (N_15333,N_11235,N_14819);
or U15334 (N_15334,N_14453,N_13380);
and U15335 (N_15335,N_11890,N_11164);
and U15336 (N_15336,N_13193,N_11519);
or U15337 (N_15337,N_10686,N_13326);
and U15338 (N_15338,N_10635,N_14443);
or U15339 (N_15339,N_12416,N_10231);
or U15340 (N_15340,N_13375,N_14537);
or U15341 (N_15341,N_12595,N_13276);
nand U15342 (N_15342,N_12556,N_11386);
nand U15343 (N_15343,N_11481,N_11014);
nand U15344 (N_15344,N_10354,N_14179);
and U15345 (N_15345,N_13150,N_12289);
xnor U15346 (N_15346,N_10956,N_12875);
nor U15347 (N_15347,N_14577,N_12213);
or U15348 (N_15348,N_11026,N_14798);
nand U15349 (N_15349,N_10676,N_14215);
nor U15350 (N_15350,N_12762,N_13546);
or U15351 (N_15351,N_14091,N_12585);
nor U15352 (N_15352,N_13721,N_14934);
and U15353 (N_15353,N_12676,N_14162);
and U15354 (N_15354,N_13493,N_14859);
nand U15355 (N_15355,N_14302,N_10980);
or U15356 (N_15356,N_14140,N_13389);
nor U15357 (N_15357,N_10419,N_10543);
and U15358 (N_15358,N_11822,N_14032);
nand U15359 (N_15359,N_14876,N_14599);
or U15360 (N_15360,N_12083,N_11841);
nand U15361 (N_15361,N_13427,N_13360);
nand U15362 (N_15362,N_10045,N_12553);
nor U15363 (N_15363,N_11506,N_10343);
and U15364 (N_15364,N_10641,N_13497);
or U15365 (N_15365,N_10292,N_11030);
nor U15366 (N_15366,N_12307,N_10681);
nand U15367 (N_15367,N_14732,N_14248);
nor U15368 (N_15368,N_10017,N_12751);
nor U15369 (N_15369,N_11942,N_12698);
nor U15370 (N_15370,N_13077,N_11945);
nor U15371 (N_15371,N_12039,N_10489);
or U15372 (N_15372,N_10487,N_13498);
xnor U15373 (N_15373,N_10690,N_14483);
nor U15374 (N_15374,N_13643,N_11917);
or U15375 (N_15375,N_11862,N_12961);
or U15376 (N_15376,N_14787,N_10553);
nor U15377 (N_15377,N_13334,N_10083);
or U15378 (N_15378,N_12765,N_11743);
nor U15379 (N_15379,N_13808,N_12980);
nand U15380 (N_15380,N_13776,N_12815);
nand U15381 (N_15381,N_10525,N_12703);
xor U15382 (N_15382,N_10652,N_13907);
xnor U15383 (N_15383,N_11755,N_10629);
nand U15384 (N_15384,N_11690,N_14011);
and U15385 (N_15385,N_13917,N_12082);
and U15386 (N_15386,N_11677,N_12562);
nor U15387 (N_15387,N_10408,N_13835);
or U15388 (N_15388,N_13107,N_12646);
nand U15389 (N_15389,N_10861,N_13031);
and U15390 (N_15390,N_12216,N_10673);
and U15391 (N_15391,N_14209,N_12163);
or U15392 (N_15392,N_10898,N_10600);
nand U15393 (N_15393,N_14656,N_11697);
nand U15394 (N_15394,N_10663,N_11166);
nor U15395 (N_15395,N_14720,N_12386);
and U15396 (N_15396,N_14661,N_12155);
nor U15397 (N_15397,N_13631,N_14167);
nor U15398 (N_15398,N_13946,N_11932);
and U15399 (N_15399,N_14441,N_13344);
and U15400 (N_15400,N_10148,N_12790);
nor U15401 (N_15401,N_12228,N_10427);
xnor U15402 (N_15402,N_14133,N_12999);
and U15403 (N_15403,N_14247,N_10779);
nand U15404 (N_15404,N_11603,N_11751);
and U15405 (N_15405,N_12257,N_12379);
nor U15406 (N_15406,N_12223,N_14989);
or U15407 (N_15407,N_12924,N_14212);
xor U15408 (N_15408,N_14766,N_14643);
xnor U15409 (N_15409,N_13618,N_14923);
or U15410 (N_15410,N_11107,N_10154);
nand U15411 (N_15411,N_12639,N_10182);
nor U15412 (N_15412,N_14684,N_13865);
xor U15413 (N_15413,N_14096,N_10417);
nand U15414 (N_15414,N_10725,N_12810);
nand U15415 (N_15415,N_12165,N_14403);
and U15416 (N_15416,N_14186,N_12904);
nor U15417 (N_15417,N_13041,N_13428);
nor U15418 (N_15418,N_14314,N_11093);
nand U15419 (N_15419,N_14366,N_12884);
or U15420 (N_15420,N_14956,N_10243);
nor U15421 (N_15421,N_12594,N_14603);
and U15422 (N_15422,N_12078,N_10620);
nand U15423 (N_15423,N_10420,N_13190);
nor U15424 (N_15424,N_13851,N_12352);
and U15425 (N_15425,N_11865,N_14786);
or U15426 (N_15426,N_12874,N_13370);
nand U15427 (N_15427,N_13432,N_12178);
or U15428 (N_15428,N_13521,N_11002);
xnor U15429 (N_15429,N_10377,N_13172);
nand U15430 (N_15430,N_14872,N_14894);
and U15431 (N_15431,N_12481,N_11408);
xor U15432 (N_15432,N_14097,N_11678);
and U15433 (N_15433,N_14871,N_10440);
nand U15434 (N_15434,N_10880,N_11976);
or U15435 (N_15435,N_11368,N_12467);
and U15436 (N_15436,N_11667,N_11117);
xor U15437 (N_15437,N_13482,N_14848);
nand U15438 (N_15438,N_13695,N_10029);
nor U15439 (N_15439,N_12260,N_13343);
nor U15440 (N_15440,N_12789,N_13515);
or U15441 (N_15441,N_13846,N_14561);
nand U15442 (N_15442,N_11411,N_12578);
nor U15443 (N_15443,N_12334,N_11307);
and U15444 (N_15444,N_13538,N_11172);
nor U15445 (N_15445,N_10241,N_12383);
nand U15446 (N_15446,N_13789,N_13161);
nor U15447 (N_15447,N_14838,N_14448);
or U15448 (N_15448,N_13435,N_10967);
and U15449 (N_15449,N_10602,N_11643);
nand U15450 (N_15450,N_13129,N_14862);
nand U15451 (N_15451,N_13264,N_10555);
xor U15452 (N_15452,N_11471,N_12060);
and U15453 (N_15453,N_14926,N_14957);
nor U15454 (N_15454,N_12568,N_10213);
or U15455 (N_15455,N_14410,N_12505);
and U15456 (N_15456,N_12032,N_10518);
or U15457 (N_15457,N_14583,N_12317);
or U15458 (N_15458,N_11431,N_14893);
and U15459 (N_15459,N_14852,N_13166);
nor U15460 (N_15460,N_11018,N_12330);
and U15461 (N_15461,N_12206,N_14892);
xor U15462 (N_15462,N_12957,N_10070);
nor U15463 (N_15463,N_11683,N_12143);
xnor U15464 (N_15464,N_11350,N_12597);
and U15465 (N_15465,N_14356,N_10131);
nor U15466 (N_15466,N_13899,N_14450);
nand U15467 (N_15467,N_12826,N_10591);
nand U15468 (N_15468,N_11072,N_10722);
nand U15469 (N_15469,N_11314,N_10101);
or U15470 (N_15470,N_14154,N_12369);
nand U15471 (N_15471,N_13095,N_14801);
nor U15472 (N_15472,N_13927,N_13374);
and U15473 (N_15473,N_13975,N_14660);
nor U15474 (N_15474,N_11092,N_12994);
or U15475 (N_15475,N_14921,N_13358);
or U15476 (N_15476,N_11689,N_13234);
nor U15477 (N_15477,N_12284,N_11127);
nand U15478 (N_15478,N_10796,N_11855);
nor U15479 (N_15479,N_13925,N_14885);
xnor U15480 (N_15480,N_11077,N_12106);
or U15481 (N_15481,N_12857,N_10276);
nor U15482 (N_15482,N_14835,N_12350);
nor U15483 (N_15483,N_11806,N_11106);
or U15484 (N_15484,N_13205,N_10007);
nor U15485 (N_15485,N_11982,N_12552);
xor U15486 (N_15486,N_11168,N_12550);
nor U15487 (N_15487,N_11813,N_10711);
or U15488 (N_15488,N_12231,N_11154);
xnor U15489 (N_15489,N_10183,N_11146);
xor U15490 (N_15490,N_14279,N_14128);
xnor U15491 (N_15491,N_14604,N_10842);
and U15492 (N_15492,N_12007,N_13398);
nand U15493 (N_15493,N_12139,N_14884);
nor U15494 (N_15494,N_13026,N_13385);
nand U15495 (N_15495,N_14110,N_12400);
xnor U15496 (N_15496,N_14777,N_12579);
nor U15497 (N_15497,N_12209,N_13342);
xnor U15498 (N_15498,N_14646,N_13121);
nand U15499 (N_15499,N_14163,N_14092);
xnor U15500 (N_15500,N_13171,N_13449);
nor U15501 (N_15501,N_12234,N_14708);
nand U15502 (N_15502,N_14621,N_14311);
or U15503 (N_15503,N_12640,N_13941);
nand U15504 (N_15504,N_10758,N_13256);
or U15505 (N_15505,N_11091,N_10388);
nor U15506 (N_15506,N_10802,N_10933);
nor U15507 (N_15507,N_11334,N_12779);
and U15508 (N_15508,N_11910,N_10286);
or U15509 (N_15509,N_13770,N_14300);
and U15510 (N_15510,N_10564,N_13118);
or U15511 (N_15511,N_11712,N_12069);
nand U15512 (N_15512,N_12541,N_11991);
nand U15513 (N_15513,N_10483,N_11372);
nor U15514 (N_15514,N_14570,N_10165);
nor U15515 (N_15515,N_11081,N_10645);
xnor U15516 (N_15516,N_12491,N_10151);
and U15517 (N_15517,N_13839,N_11258);
xnor U15518 (N_15518,N_13341,N_13191);
or U15519 (N_15519,N_14760,N_10866);
nand U15520 (N_15520,N_11472,N_11283);
and U15521 (N_15521,N_14691,N_14584);
and U15522 (N_15522,N_13045,N_12248);
nand U15523 (N_15523,N_12110,N_11209);
nor U15524 (N_15524,N_11315,N_10049);
or U15525 (N_15525,N_13903,N_12095);
or U15526 (N_15526,N_13101,N_13353);
xnor U15527 (N_15527,N_14931,N_10998);
and U15528 (N_15528,N_14077,N_11969);
nor U15529 (N_15529,N_12715,N_14674);
and U15530 (N_15530,N_12045,N_12099);
or U15531 (N_15531,N_12434,N_10689);
or U15532 (N_15532,N_14595,N_12337);
nand U15533 (N_15533,N_14263,N_11710);
xor U15534 (N_15534,N_14797,N_14508);
nand U15535 (N_15535,N_13720,N_14575);
xnor U15536 (N_15536,N_12985,N_12159);
or U15537 (N_15537,N_11611,N_11450);
and U15538 (N_15538,N_11324,N_13864);
or U15539 (N_15539,N_11487,N_10585);
xor U15540 (N_15540,N_12079,N_11968);
or U15541 (N_15541,N_11308,N_12494);
xor U15542 (N_15542,N_13309,N_12536);
xor U15543 (N_15543,N_11867,N_11940);
nor U15544 (N_15544,N_11538,N_12878);
and U15545 (N_15545,N_13536,N_10149);
or U15546 (N_15546,N_10252,N_12354);
nor U15547 (N_15547,N_10275,N_11800);
and U15548 (N_15548,N_12098,N_14175);
nand U15549 (N_15549,N_12199,N_12956);
nor U15550 (N_15550,N_11918,N_13630);
and U15551 (N_15551,N_14739,N_13758);
nor U15552 (N_15552,N_13016,N_12405);
xnor U15553 (N_15553,N_11378,N_13258);
nand U15554 (N_15554,N_12653,N_10434);
nor U15555 (N_15555,N_14420,N_12665);
nand U15556 (N_15556,N_10872,N_12627);
xnor U15557 (N_15557,N_10738,N_11464);
xor U15558 (N_15558,N_13136,N_12480);
xor U15559 (N_15559,N_14073,N_14569);
nor U15560 (N_15560,N_13554,N_11842);
xnor U15561 (N_15561,N_13155,N_14672);
nand U15562 (N_15562,N_10744,N_14008);
and U15563 (N_15563,N_10567,N_14006);
or U15564 (N_15564,N_10819,N_10609);
nand U15565 (N_15565,N_12210,N_12743);
nand U15566 (N_15566,N_11486,N_10785);
and U15567 (N_15567,N_11210,N_13599);
or U15568 (N_15568,N_12498,N_11271);
nand U15569 (N_15569,N_13913,N_12971);
xnor U15570 (N_15570,N_12911,N_14552);
or U15571 (N_15571,N_10185,N_12170);
and U15572 (N_15572,N_14728,N_14353);
and U15573 (N_15573,N_11859,N_10671);
nand U15574 (N_15574,N_12226,N_12667);
xnor U15575 (N_15575,N_11041,N_10088);
and U15576 (N_15576,N_11605,N_10858);
and U15577 (N_15577,N_10820,N_10195);
and U15578 (N_15578,N_14670,N_14009);
xnor U15579 (N_15579,N_13868,N_13186);
nand U15580 (N_15580,N_10118,N_13842);
or U15581 (N_15581,N_10930,N_12012);
nor U15582 (N_15582,N_12456,N_10373);
and U15583 (N_15583,N_11478,N_12222);
nand U15584 (N_15584,N_10821,N_13873);
xor U15585 (N_15585,N_14232,N_11375);
or U15586 (N_15586,N_13333,N_13518);
nor U15587 (N_15587,N_12712,N_11775);
and U15588 (N_15588,N_14357,N_11507);
and U15589 (N_15589,N_10953,N_13516);
nor U15590 (N_15590,N_14540,N_13701);
and U15591 (N_15591,N_14049,N_12133);
and U15592 (N_15592,N_14948,N_11061);
xnor U15593 (N_15593,N_13650,N_11809);
and U15594 (N_15594,N_11440,N_10472);
nand U15595 (N_15595,N_10885,N_10982);
nand U15596 (N_15596,N_12802,N_10074);
nand U15597 (N_15597,N_11068,N_13010);
and U15598 (N_15598,N_12732,N_10386);
nand U15599 (N_15599,N_14509,N_12745);
nand U15600 (N_15600,N_12218,N_14249);
and U15601 (N_15601,N_14461,N_11391);
or U15602 (N_15602,N_13106,N_11766);
or U15603 (N_15603,N_13262,N_12177);
xnor U15604 (N_15604,N_12907,N_11461);
nor U15605 (N_15605,N_10636,N_11734);
nor U15606 (N_15606,N_14711,N_12273);
and U15607 (N_15607,N_10648,N_10644);
or U15608 (N_15608,N_13577,N_14890);
and U15609 (N_15609,N_13117,N_10436);
and U15610 (N_15610,N_11429,N_12607);
nor U15611 (N_15611,N_11058,N_10848);
nand U15612 (N_15612,N_10201,N_10749);
nand U15613 (N_15613,N_10664,N_11233);
nor U15614 (N_15614,N_10190,N_10989);
or U15615 (N_15615,N_13763,N_11143);
nor U15616 (N_15616,N_12845,N_14642);
or U15617 (N_15617,N_11384,N_10053);
and U15618 (N_15618,N_10186,N_13263);
nand U15619 (N_15619,N_13743,N_12824);
xnor U15620 (N_15620,N_12649,N_14294);
xnor U15621 (N_15621,N_13500,N_10776);
xor U15622 (N_15622,N_11073,N_14391);
xnor U15623 (N_15623,N_10854,N_10304);
or U15624 (N_15624,N_10338,N_13257);
nor U15625 (N_15625,N_10775,N_11063);
nor U15626 (N_15626,N_14390,N_11133);
and U15627 (N_15627,N_13861,N_10557);
xor U15628 (N_15628,N_10882,N_13109);
or U15629 (N_15629,N_13854,N_12168);
and U15630 (N_15630,N_13894,N_13197);
nand U15631 (N_15631,N_10089,N_12784);
or U15632 (N_15632,N_11995,N_14429);
nor U15633 (N_15633,N_13816,N_13102);
and U15634 (N_15634,N_14896,N_13069);
or U15635 (N_15635,N_10329,N_13908);
nor U15636 (N_15636,N_12657,N_12516);
or U15637 (N_15637,N_11704,N_11497);
or U15638 (N_15638,N_10081,N_14280);
or U15639 (N_15639,N_13088,N_10345);
nand U15640 (N_15640,N_11654,N_12402);
or U15641 (N_15641,N_12056,N_10562);
xnor U15642 (N_15642,N_12409,N_11369);
or U15643 (N_15643,N_14292,N_10916);
nand U15644 (N_15644,N_14015,N_13407);
nor U15645 (N_15645,N_14800,N_11948);
and U15646 (N_15646,N_14445,N_11419);
and U15647 (N_15647,N_13635,N_13047);
or U15648 (N_15648,N_14206,N_12914);
xor U15649 (N_15649,N_13212,N_11257);
or U15650 (N_15650,N_13692,N_12117);
nor U15651 (N_15651,N_11124,N_10340);
xnor U15652 (N_15652,N_13504,N_10546);
nand U15653 (N_15653,N_13980,N_14053);
and U15654 (N_15654,N_13653,N_14628);
nand U15655 (N_15655,N_13209,N_14433);
nand U15656 (N_15656,N_14914,N_12894);
and U15657 (N_15657,N_14993,N_11584);
and U15658 (N_15658,N_11847,N_13638);
or U15659 (N_15659,N_10096,N_14273);
and U15660 (N_15660,N_13046,N_12127);
xor U15661 (N_15661,N_13718,N_13268);
or U15662 (N_15662,N_11186,N_14377);
or U15663 (N_15663,N_13531,N_13133);
nand U15664 (N_15664,N_14571,N_11820);
nor U15665 (N_15665,N_10347,N_13002);
nand U15666 (N_15666,N_14276,N_13152);
xor U15667 (N_15667,N_14253,N_10958);
and U15668 (N_15668,N_11682,N_13594);
and U15669 (N_15669,N_11035,N_13814);
nand U15670 (N_15670,N_14134,N_13290);
or U15671 (N_15671,N_13569,N_12723);
nor U15672 (N_15672,N_11627,N_13489);
nand U15673 (N_15673,N_12741,N_12269);
xor U15674 (N_15674,N_10192,N_12717);
xor U15675 (N_15675,N_13885,N_12807);
and U15676 (N_15676,N_10670,N_11115);
or U15677 (N_15677,N_11551,N_10742);
xnor U15678 (N_15678,N_11632,N_12343);
and U15679 (N_15679,N_11051,N_10710);
nand U15680 (N_15680,N_13510,N_10856);
or U15681 (N_15681,N_10490,N_10996);
and U15682 (N_15682,N_12420,N_11728);
nor U15683 (N_15683,N_10753,N_13361);
and U15684 (N_15684,N_12920,N_10468);
xnor U15685 (N_15685,N_11298,N_13440);
xor U15686 (N_15686,N_12535,N_13462);
and U15687 (N_15687,N_12638,N_13859);
or U15688 (N_15688,N_10103,N_13791);
xor U15689 (N_15689,N_11056,N_14342);
nand U15690 (N_15690,N_11279,N_10326);
or U15691 (N_15691,N_13784,N_11764);
xnor U15692 (N_15692,N_12834,N_10056);
and U15693 (N_15693,N_10457,N_12811);
xnor U15694 (N_15694,N_13750,N_12382);
or U15695 (N_15695,N_12136,N_14974);
xor U15696 (N_15696,N_11090,N_12839);
and U15697 (N_15697,N_11479,N_10402);
nand U15698 (N_15698,N_14693,N_13847);
and U15699 (N_15699,N_10293,N_10253);
xor U15700 (N_15700,N_14736,N_12708);
nand U15701 (N_15701,N_13349,N_12711);
nor U15702 (N_15702,N_13725,N_10556);
and U15703 (N_15703,N_14454,N_11175);
xor U15704 (N_15704,N_12392,N_11513);
nor U15705 (N_15705,N_10215,N_10804);
or U15706 (N_15706,N_12782,N_13111);
and U15707 (N_15707,N_14669,N_12859);
or U15708 (N_15708,N_14768,N_12927);
nor U15709 (N_15709,N_11700,N_11114);
or U15710 (N_15710,N_14194,N_10311);
xor U15711 (N_15711,N_10113,N_10289);
xnor U15712 (N_15712,N_10581,N_11219);
nand U15713 (N_15713,N_14917,N_11021);
nor U15714 (N_15714,N_11729,N_14502);
nand U15715 (N_15715,N_14496,N_14141);
nand U15716 (N_15716,N_12929,N_12942);
nand U15717 (N_15717,N_14233,N_14068);
or U15718 (N_15718,N_13716,N_11373);
nand U15719 (N_15719,N_11745,N_12995);
nor U15720 (N_15720,N_13229,N_11121);
nand U15721 (N_15721,N_13583,N_12518);
nor U15722 (N_15722,N_13739,N_13356);
nand U15723 (N_15723,N_11784,N_13831);
xor U15724 (N_15724,N_10550,N_10884);
xnor U15725 (N_15725,N_14109,N_13395);
or U15726 (N_15726,N_11005,N_10571);
and U15727 (N_15727,N_12174,N_13242);
nand U15728 (N_15728,N_14423,N_11923);
nand U15729 (N_15729,N_10244,N_11407);
nor U15730 (N_15730,N_11814,N_14617);
or U15731 (N_15731,N_14939,N_14452);
and U15732 (N_15732,N_12508,N_13036);
xnor U15733 (N_15733,N_10097,N_11663);
or U15734 (N_15734,N_11400,N_12035);
nand U15735 (N_15735,N_14323,N_14650);
nor U15736 (N_15736,N_10206,N_11054);
nor U15737 (N_15737,N_14022,N_14869);
nand U15738 (N_15738,N_10528,N_12247);
nor U15739 (N_15739,N_10694,N_11297);
xnor U15740 (N_15740,N_10294,N_14773);
or U15741 (N_15741,N_12261,N_14550);
or U15742 (N_15742,N_13066,N_10886);
and U15743 (N_15743,N_10010,N_14112);
nand U15744 (N_15744,N_11260,N_12970);
nor U15745 (N_15745,N_13104,N_13433);
nand U15746 (N_15746,N_14426,N_13645);
nor U15747 (N_15747,N_14153,N_10979);
nand U15748 (N_15748,N_13676,N_11211);
nor U15749 (N_15749,N_14358,N_13123);
or U15750 (N_15750,N_10020,N_12224);
xnor U15751 (N_15751,N_12264,N_14372);
nand U15752 (N_15752,N_13681,N_13062);
nand U15753 (N_15753,N_13723,N_14718);
nor U15754 (N_15754,N_12062,N_13843);
xnor U15755 (N_15755,N_14776,N_11869);
and U15756 (N_15756,N_12982,N_11126);
or U15757 (N_15757,N_11171,N_14516);
xnor U15758 (N_15758,N_14199,N_11934);
nor U15759 (N_15759,N_13619,N_14677);
and U15760 (N_15760,N_12972,N_14350);
nor U15761 (N_15761,N_10551,N_14227);
and U15762 (N_15762,N_10561,N_12085);
nand U15763 (N_15763,N_12860,N_11252);
nand U15764 (N_15764,N_14295,N_13587);
nand U15765 (N_15765,N_10392,N_10833);
nand U15766 (N_15766,N_14903,N_13365);
nor U15767 (N_15767,N_14854,N_10590);
nand U15768 (N_15768,N_11578,N_12476);
xnor U15769 (N_15769,N_11649,N_14207);
or U15770 (N_15770,N_14401,N_11698);
nor U15771 (N_15771,N_11136,N_13932);
nor U15772 (N_15772,N_12820,N_11435);
nor U15773 (N_15773,N_10757,N_10344);
and U15774 (N_15774,N_13421,N_10279);
xor U15775 (N_15775,N_11212,N_10939);
nand U15776 (N_15776,N_13447,N_11492);
and U15777 (N_15777,N_14521,N_13898);
nor U15778 (N_15778,N_14034,N_14513);
xor U15779 (N_15779,N_11893,N_13651);
or U15780 (N_15780,N_12080,N_11128);
nand U15781 (N_15781,N_10999,N_12315);
or U15782 (N_15782,N_12065,N_13476);
or U15783 (N_15783,N_11548,N_11490);
and U15784 (N_15784,N_11336,N_13128);
nor U15785 (N_15785,N_11240,N_13802);
xor U15786 (N_15786,N_10895,N_10891);
and U15787 (N_15787,N_11912,N_14875);
nand U15788 (N_15788,N_13699,N_11480);
xor U15789 (N_15789,N_10351,N_10396);
nand U15790 (N_15790,N_10342,N_10516);
xor U15791 (N_15791,N_10972,N_11392);
xor U15792 (N_15792,N_14613,N_10589);
xnor U15793 (N_15793,N_10161,N_12933);
xnor U15794 (N_15794,N_10091,N_10018);
or U15795 (N_15795,N_14655,N_10280);
xnor U15796 (N_15796,N_10868,N_14769);
and U15797 (N_15797,N_11185,N_12767);
nand U15798 (N_15798,N_12577,N_11006);
nand U15799 (N_15799,N_12191,N_10565);
xnor U15800 (N_15800,N_11130,N_10307);
and U15801 (N_15801,N_11402,N_13513);
nand U15802 (N_15802,N_13967,N_12504);
and U15803 (N_15803,N_11085,N_12532);
nand U15804 (N_15804,N_14526,N_14726);
nand U15805 (N_15805,N_14754,N_14159);
nand U15806 (N_15806,N_11097,N_10899);
and U15807 (N_15807,N_10965,N_10734);
or U15808 (N_15808,N_11355,N_10110);
and U15809 (N_15809,N_10583,N_10537);
nor U15810 (N_15810,N_13682,N_11846);
and U15811 (N_15811,N_13426,N_11984);
and U15812 (N_15812,N_11265,N_11770);
or U15813 (N_15813,N_11349,N_14335);
and U15814 (N_15814,N_11184,N_13070);
or U15815 (N_15815,N_14239,N_11330);
nand U15816 (N_15816,N_11142,N_14145);
nor U15817 (N_15817,N_10860,N_13690);
and U15818 (N_15818,N_14764,N_14594);
or U15819 (N_15819,N_11250,N_13231);
or U15820 (N_15820,N_12678,N_11189);
and U15821 (N_15821,N_12034,N_11939);
or U15822 (N_15822,N_12949,N_12852);
xnor U15823 (N_15823,N_14161,N_12812);
and U15824 (N_15824,N_12948,N_14297);
and U15825 (N_15825,N_13024,N_10701);
xnor U15826 (N_15826,N_12629,N_13078);
nor U15827 (N_15827,N_13757,N_11112);
xnor U15828 (N_15828,N_10055,N_13265);
or U15829 (N_15829,N_13534,N_13085);
xnor U15830 (N_15830,N_12636,N_13911);
xnor U15831 (N_15831,N_10699,N_12913);
nand U15832 (N_15832,N_12674,N_13003);
xor U15833 (N_15833,N_12087,N_12195);
and U15834 (N_15834,N_10510,N_13336);
and U15835 (N_15835,N_10432,N_12605);
and U15836 (N_15836,N_13998,N_11489);
nor U15837 (N_15837,N_10981,N_13005);
and U15838 (N_15838,N_13856,N_14856);
nor U15839 (N_15839,N_14841,N_11438);
nand U15840 (N_15840,N_11303,N_10482);
nor U15841 (N_15841,N_14244,N_12644);
xnor U15842 (N_15842,N_14775,N_10807);
and U15843 (N_15843,N_11340,N_11759);
nor U15844 (N_15844,N_14345,N_13138);
nand U15845 (N_15845,N_11541,N_10484);
and U15846 (N_15846,N_11230,N_12372);
nand U15847 (N_15847,N_14782,N_12974);
or U15848 (N_15848,N_12214,N_13384);
xor U15849 (N_15849,N_10065,N_14396);
nor U15850 (N_15850,N_10803,N_11824);
nand U15851 (N_15851,N_12005,N_10502);
and U15852 (N_15852,N_14688,N_12356);
xor U15853 (N_15853,N_11229,N_11526);
nand U15854 (N_15854,N_10677,N_10829);
nor U15855 (N_15855,N_11153,N_12515);
or U15856 (N_15856,N_10200,N_12808);
nor U15857 (N_15857,N_13054,N_14122);
nand U15858 (N_15858,N_13823,N_11978);
and U15859 (N_15859,N_11076,N_14664);
nand U15860 (N_15860,N_14173,N_14733);
nor U15861 (N_15861,N_10669,N_12371);
and U15862 (N_15862,N_10414,N_13875);
nor U15863 (N_15863,N_12531,N_13141);
nand U15864 (N_15864,N_14127,N_14172);
nand U15865 (N_15865,N_10793,N_13411);
and U15866 (N_15866,N_13735,N_14045);
nor U15867 (N_15867,N_13278,N_12003);
nor U15868 (N_15868,N_10897,N_11223);
nand U15869 (N_15869,N_13206,N_11239);
nand U15870 (N_15870,N_10831,N_14258);
or U15871 (N_15871,N_10260,N_11563);
nor U15872 (N_15872,N_10724,N_10384);
nand U15873 (N_15873,N_10631,N_13548);
nand U15874 (N_15874,N_10129,N_14831);
xnor U15875 (N_15875,N_14899,N_10034);
nand U15876 (N_15876,N_11017,N_13857);
and U15877 (N_15877,N_13185,N_13580);
xnor U15878 (N_15878,N_13475,N_11278);
and U15879 (N_15879,N_10274,N_14517);
or U15880 (N_15880,N_14399,N_13335);
nor U15881 (N_15881,N_12363,N_11529);
or U15882 (N_15882,N_11666,N_13633);
xor U15883 (N_15883,N_10665,N_12061);
or U15884 (N_15884,N_11452,N_11518);
xor U15885 (N_15885,N_12527,N_13551);
nor U15886 (N_15886,N_10799,N_10594);
or U15887 (N_15887,N_12699,N_11718);
xnor U15888 (N_15888,N_12204,N_10403);
nand U15889 (N_15889,N_11804,N_14932);
xor U15890 (N_15890,N_10816,N_12414);
nand U15891 (N_15891,N_11034,N_12537);
nor U15892 (N_15892,N_13487,N_10728);
nor U15893 (N_15893,N_10177,N_10878);
or U15894 (N_15894,N_13805,N_14070);
nand U15895 (N_15895,N_14230,N_11737);
nor U15896 (N_15896,N_10517,N_12001);
xnor U15897 (N_15897,N_14648,N_11533);
and U15898 (N_15898,N_10471,N_12814);
nand U15899 (N_15899,N_12736,N_10375);
nand U15900 (N_15900,N_10078,N_13429);
and U15901 (N_15901,N_13821,N_12669);
nor U15902 (N_15902,N_13292,N_14181);
nand U15903 (N_15903,N_12058,N_13139);
or U15904 (N_15904,N_10957,N_13480);
or U15905 (N_15905,N_13576,N_14649);
and U15906 (N_15906,N_12026,N_11875);
xor U15907 (N_15907,N_14228,N_12015);
nand U15908 (N_15908,N_14808,N_10367);
xor U15909 (N_15909,N_12819,N_10615);
xor U15910 (N_15910,N_13921,N_10040);
nor U15911 (N_15911,N_13922,N_13874);
nand U15912 (N_15912,N_11220,N_13094);
nand U15913 (N_15913,N_10291,N_10838);
nand U15914 (N_15914,N_13465,N_10577);
xnor U15915 (N_15915,N_13841,N_14013);
nor U15916 (N_15916,N_13367,N_12362);
nor U15917 (N_15917,N_11854,N_11467);
or U15918 (N_15918,N_14746,N_11858);
nand U15919 (N_15919,N_13059,N_11987);
nand U15920 (N_15920,N_14544,N_12725);
or U15921 (N_15921,N_13568,N_12471);
nor U15922 (N_15922,N_10224,N_13355);
or U15923 (N_15923,N_12840,N_13082);
and U15924 (N_15924,N_13064,N_10114);
nand U15925 (N_15925,N_11359,N_14143);
nor U15926 (N_15926,N_14216,N_10315);
and U15927 (N_15927,N_12668,N_11730);
xor U15928 (N_15928,N_12131,N_12166);
or U15929 (N_15929,N_13153,N_11294);
and U15930 (N_15930,N_12108,N_13657);
and U15931 (N_15931,N_11389,N_13646);
nand U15932 (N_15932,N_12014,N_13964);
and U15933 (N_15933,N_13648,N_14486);
nand U15934 (N_15934,N_13639,N_14380);
nor U15935 (N_15935,N_11610,N_14193);
and U15936 (N_15936,N_10314,N_11790);
nand U15937 (N_15937,N_14115,N_11545);
nand U15938 (N_15938,N_11195,N_13994);
nor U15939 (N_15939,N_14472,N_14229);
and U15940 (N_15940,N_14160,N_11746);
xor U15941 (N_15941,N_14290,N_10355);
nor U15942 (N_15942,N_13833,N_11607);
xor U15943 (N_15943,N_13072,N_12490);
and U15944 (N_15944,N_11662,N_10374);
and U15945 (N_15945,N_12691,N_11342);
nand U15946 (N_15946,N_12831,N_10625);
and U15947 (N_15947,N_10474,N_14721);
or U15948 (N_15948,N_13673,N_11963);
and U15949 (N_15949,N_11491,N_13008);
and U15950 (N_15950,N_12380,N_13297);
xor U15951 (N_15951,N_10568,N_14999);
and U15952 (N_15952,N_11780,N_13519);
and U15953 (N_15953,N_12692,N_10205);
or U15954 (N_15954,N_11664,N_14967);
nor U15955 (N_15955,N_11769,N_10041);
nor U15956 (N_15956,N_12773,N_12374);
and U15957 (N_15957,N_11422,N_13752);
and U15958 (N_15958,N_11426,N_13968);
nand U15959 (N_15959,N_10228,N_11364);
xnor U15960 (N_15960,N_12953,N_12318);
or U15961 (N_15961,N_13175,N_11403);
nand U15962 (N_15962,N_14416,N_13165);
xor U15963 (N_15963,N_10444,N_12277);
xor U15964 (N_15964,N_10046,N_10923);
and U15965 (N_15965,N_11980,N_10806);
xor U15966 (N_15966,N_12237,N_14278);
and U15967 (N_15967,N_10991,N_14622);
xnor U15968 (N_15968,N_13656,N_10063);
or U15969 (N_15969,N_12121,N_14137);
xor U15970 (N_15970,N_14881,N_14218);
nand U15971 (N_15971,N_12298,N_11811);
xor U15972 (N_15972,N_13252,N_13601);
and U15973 (N_15973,N_10545,N_10169);
nor U15974 (N_15974,N_10951,N_13658);
nand U15975 (N_15975,N_14155,N_11835);
nor U15976 (N_15976,N_11639,N_13316);
nor U15977 (N_15977,N_10385,N_10705);
or U15978 (N_15978,N_13606,N_13729);
or U15979 (N_15979,N_14818,N_14059);
nor U15980 (N_15980,N_11510,N_14639);
nand U15981 (N_15981,N_13413,N_11238);
or U15982 (N_15982,N_11572,N_10623);
nor U15983 (N_15983,N_12347,N_12522);
and U15984 (N_15984,N_10339,N_11398);
or U15985 (N_15985,N_12485,N_14125);
nand U15986 (N_15986,N_10143,N_13140);
xor U15987 (N_15987,N_13460,N_10515);
or U15988 (N_15988,N_14889,N_13424);
or U15989 (N_15989,N_13216,N_11059);
xor U15990 (N_15990,N_11874,N_13312);
xnor U15991 (N_15991,N_14041,N_14421);
and U15992 (N_15992,N_10859,N_14730);
nand U15993 (N_15993,N_14406,N_14455);
nand U15994 (N_15994,N_12479,N_13456);
nor U15995 (N_15995,N_12570,N_14477);
and U15996 (N_15996,N_10873,N_10617);
or U15997 (N_15997,N_10707,N_11177);
and U15998 (N_15998,N_13419,N_13366);
and U15999 (N_15999,N_13775,N_13289);
xor U16000 (N_16000,N_10334,N_11843);
nor U16001 (N_16001,N_13350,N_13997);
nor U16002 (N_16002,N_14902,N_11152);
nor U16003 (N_16003,N_10781,N_13853);
or U16004 (N_16004,N_11782,N_11145);
xor U16005 (N_16005,N_14565,N_11618);
or U16006 (N_16006,N_12947,N_12462);
nand U16007 (N_16007,N_13373,N_13293);
nand U16008 (N_16008,N_11834,N_11753);
xor U16009 (N_16009,N_12656,N_10601);
and U16010 (N_16010,N_14418,N_14714);
nand U16011 (N_16011,N_10287,N_12190);
or U16012 (N_16012,N_10000,N_14909);
nand U16013 (N_16013,N_13314,N_13151);
nor U16014 (N_16014,N_13649,N_11993);
or U16015 (N_16015,N_11871,N_14729);
or U16016 (N_16016,N_14240,N_13662);
nand U16017 (N_16017,N_11485,N_10817);
nand U16018 (N_16018,N_11007,N_13124);
nand U16019 (N_16019,N_11337,N_10147);
or U16020 (N_16020,N_11960,N_10795);
and U16021 (N_16021,N_10333,N_13957);
nor U16022 (N_16022,N_13837,N_12387);
nor U16023 (N_16023,N_13990,N_11567);
nand U16024 (N_16024,N_14467,N_14555);
and U16025 (N_16025,N_10748,N_10513);
or U16026 (N_16026,N_10219,N_13812);
nand U16027 (N_16027,N_11815,N_13572);
or U16028 (N_16028,N_13299,N_13915);
and U16029 (N_16029,N_13844,N_11935);
and U16030 (N_16030,N_13086,N_10520);
xnor U16031 (N_16031,N_14855,N_13445);
nor U16032 (N_16032,N_12144,N_13158);
nor U16033 (N_16033,N_11985,N_12599);
nor U16034 (N_16034,N_11591,N_10921);
and U16035 (N_16035,N_13090,N_13704);
nor U16036 (N_16036,N_10269,N_14333);
nand U16037 (N_16037,N_13738,N_10002);
nor U16038 (N_16038,N_14202,N_14238);
nor U16039 (N_16039,N_12399,N_12730);
xnor U16040 (N_16040,N_12707,N_10187);
xor U16041 (N_16041,N_10809,N_11406);
xor U16042 (N_16042,N_10013,N_13755);
nor U16043 (N_16043,N_11242,N_13891);
xnor U16044 (N_16044,N_10801,N_13953);
and U16045 (N_16045,N_14148,N_10592);
or U16046 (N_16046,N_14562,N_13920);
xnor U16047 (N_16047,N_11031,N_13969);
or U16048 (N_16048,N_13838,N_13458);
and U16049 (N_16049,N_13637,N_10117);
and U16050 (N_16050,N_11267,N_13300);
xnor U16051 (N_16051,N_10918,N_11331);
or U16052 (N_16052,N_14742,N_10443);
nand U16053 (N_16053,N_12664,N_14791);
xor U16054 (N_16054,N_14470,N_14374);
or U16055 (N_16055,N_14007,N_11290);
and U16056 (N_16056,N_14817,N_13545);
xor U16057 (N_16057,N_14676,N_10077);
or U16058 (N_16058,N_13785,N_11319);
or U16059 (N_16059,N_12827,N_13553);
xor U16060 (N_16060,N_14339,N_10660);
nand U16061 (N_16061,N_12067,N_14289);
or U16062 (N_16062,N_14381,N_12724);
xnor U16063 (N_16063,N_10092,N_12036);
or U16064 (N_16064,N_14471,N_10654);
or U16065 (N_16065,N_10765,N_13959);
and U16066 (N_16066,N_12053,N_12357);
or U16067 (N_16067,N_12321,N_14860);
or U16068 (N_16068,N_12871,N_10762);
nor U16069 (N_16069,N_14900,N_14094);
or U16070 (N_16070,N_10718,N_10166);
nor U16071 (N_16071,N_10350,N_10062);
xnor U16072 (N_16072,N_10948,N_14260);
nor U16073 (N_16073,N_13719,N_13654);
nand U16074 (N_16074,N_13543,N_12754);
xor U16075 (N_16075,N_10433,N_12828);
or U16076 (N_16076,N_12503,N_12930);
nand U16077 (N_16077,N_12763,N_14462);
nand U16078 (N_16078,N_12800,N_11405);
xor U16079 (N_16079,N_14063,N_14359);
nand U16080 (N_16080,N_14904,N_14990);
xnor U16081 (N_16081,N_14336,N_13985);
and U16082 (N_16082,N_12854,N_12279);
xnor U16083 (N_16083,N_10808,N_12395);
xnor U16084 (N_16084,N_12013,N_11262);
nor U16085 (N_16085,N_12146,N_14633);
and U16086 (N_16086,N_10535,N_13715);
nand U16087 (N_16087,N_14054,N_12928);
and U16088 (N_16088,N_12652,N_10379);
or U16089 (N_16089,N_11050,N_11036);
or U16090 (N_16090,N_13501,N_14363);
or U16091 (N_16091,N_11708,N_14442);
xnor U16092 (N_16092,N_10301,N_11088);
or U16093 (N_16093,N_12282,N_10005);
and U16094 (N_16094,N_10769,N_10890);
nand U16095 (N_16095,N_13677,N_12189);
and U16096 (N_16096,N_12348,N_12129);
nand U16097 (N_16097,N_13782,N_11199);
and U16098 (N_16098,N_12310,N_14944);
and U16099 (N_16099,N_14641,N_12184);
nand U16100 (N_16100,N_14828,N_12685);
or U16101 (N_16101,N_10030,N_14370);
nor U16102 (N_16102,N_12153,N_11488);
xor U16103 (N_16103,N_12281,N_10947);
nand U16104 (N_16104,N_10211,N_10352);
nand U16105 (N_16105,N_11901,N_13028);
nor U16106 (N_16106,N_14040,N_12908);
xnor U16107 (N_16107,N_14036,N_14004);
xnor U16108 (N_16108,N_12308,N_13686);
nand U16109 (N_16109,N_13034,N_10262);
nand U16110 (N_16110,N_11915,N_12447);
xnor U16111 (N_16111,N_11289,N_11460);
and U16112 (N_16112,N_12128,N_10595);
nor U16113 (N_16113,N_13328,N_12569);
nor U16114 (N_16114,N_10574,N_12979);
nand U16115 (N_16115,N_10668,N_12066);
or U16116 (N_16116,N_14593,N_11621);
and U16117 (N_16117,N_14779,N_13605);
and U16118 (N_16118,N_11316,N_12891);
nor U16119 (N_16119,N_14717,N_11971);
nor U16120 (N_16120,N_14789,N_11613);
nand U16121 (N_16121,N_11911,N_14197);
and U16122 (N_16122,N_13533,N_12981);
and U16123 (N_16123,N_13277,N_14183);
nor U16124 (N_16124,N_14103,N_11925);
nor U16125 (N_16125,N_12358,N_11011);
or U16126 (N_16126,N_11779,N_10942);
nand U16127 (N_16127,N_13348,N_13267);
xnor U16128 (N_16128,N_14581,N_10907);
and U16129 (N_16129,N_13463,N_11335);
or U16130 (N_16130,N_11374,N_12091);
nor U16131 (N_16131,N_13795,N_11637);
or U16132 (N_16132,N_11266,N_14304);
and U16133 (N_16133,N_10531,N_14833);
nand U16134 (N_16134,N_10746,N_12415);
and U16135 (N_16135,N_13944,N_10786);
or U16136 (N_16136,N_14494,N_11619);
or U16137 (N_16137,N_10473,N_13415);
and U16138 (N_16138,N_10607,N_14574);
xor U16139 (N_16139,N_11920,N_11620);
nor U16140 (N_16140,N_12868,N_14972);
nor U16141 (N_16141,N_13130,N_10798);
nor U16142 (N_16142,N_12786,N_11740);
nand U16143 (N_16143,N_10446,N_12647);
or U16144 (N_16144,N_13556,N_12690);
nor U16145 (N_16145,N_11789,N_10470);
nor U16146 (N_16146,N_13558,N_11762);
or U16147 (N_16147,N_11837,N_10521);
or U16148 (N_16148,N_11310,N_11864);
or U16149 (N_16149,N_10098,N_10563);
nand U16150 (N_16150,N_10102,N_12683);
and U16151 (N_16151,N_12130,N_13174);
and U16152 (N_16152,N_10455,N_12547);
nor U16153 (N_16153,N_13388,N_14048);
xnor U16154 (N_16154,N_10042,N_10879);
nand U16155 (N_16155,N_13164,N_14878);
and U16156 (N_16156,N_12862,N_12689);
and U16157 (N_16157,N_12631,N_14205);
nand U16158 (N_16158,N_14072,N_12571);
nor U16159 (N_16159,N_10439,N_11338);
xor U16160 (N_16160,N_10627,N_14277);
nor U16161 (N_16161,N_14330,N_11752);
or U16162 (N_16162,N_14226,N_13006);
nor U16163 (N_16163,N_11444,N_14331);
or U16164 (N_16164,N_13178,N_13627);
xnor U16165 (N_16165,N_12662,N_14251);
xor U16166 (N_16166,N_13075,N_10463);
and U16167 (N_16167,N_10827,N_10826);
nor U16168 (N_16168,N_12509,N_13571);
nor U16169 (N_16169,N_10008,N_14344);
or U16170 (N_16170,N_11902,N_10932);
nor U16171 (N_16171,N_10271,N_14469);
or U16172 (N_16172,N_13522,N_13376);
and U16173 (N_16173,N_13746,N_11116);
nand U16174 (N_16174,N_13801,N_10684);
and U16175 (N_16175,N_14888,N_12835);
nand U16176 (N_16176,N_10968,N_11101);
and U16177 (N_16177,N_14365,N_11553);
or U16178 (N_16178,N_10911,N_10643);
nor U16179 (N_16179,N_13792,N_13971);
and U16180 (N_16180,N_14432,N_14269);
nand U16181 (N_16181,N_10168,N_10155);
nand U16182 (N_16182,N_11104,N_11544);
nor U16183 (N_16183,N_11274,N_12704);
and U16184 (N_16184,N_10505,N_12389);
nand U16185 (N_16185,N_13942,N_14507);
xor U16186 (N_16186,N_10975,N_12314);
nor U16187 (N_16187,N_13931,N_14963);
nor U16188 (N_16188,N_11309,N_13514);
or U16189 (N_16189,N_14090,N_10395);
xnor U16190 (N_16190,N_13912,N_10383);
and U16191 (N_16191,N_14897,N_14857);
xnor U16192 (N_16192,N_11147,N_12235);
nor U16193 (N_16193,N_10399,N_14601);
nand U16194 (N_16194,N_12339,N_10969);
and U16195 (N_16195,N_11818,N_14121);
nor U16196 (N_16196,N_11996,N_11760);
or U16197 (N_16197,N_12781,N_11181);
and U16198 (N_16198,N_10862,N_13220);
nor U16199 (N_16199,N_14474,N_14644);
nand U16200 (N_16200,N_11125,N_12630);
or U16201 (N_16201,N_10970,N_12513);
and U16202 (N_16202,N_11564,N_11707);
xnor U16203 (N_16203,N_14375,N_13986);
or U16204 (N_16204,N_11880,N_11601);
and U16205 (N_16205,N_13552,N_11135);
nand U16206 (N_16206,N_14411,N_11898);
or U16207 (N_16207,N_14039,N_14067);
nor U16208 (N_16208,N_12993,N_14785);
xnor U16209 (N_16209,N_13055,N_13105);
or U16210 (N_16210,N_11661,N_13464);
or U16211 (N_16211,N_11715,N_14958);
nand U16212 (N_16212,N_10582,N_13226);
xor U16213 (N_16213,N_14531,N_14632);
nor U16214 (N_16214,N_12906,N_14157);
or U16215 (N_16215,N_11756,N_14023);
and U16216 (N_16216,N_12370,N_14827);
nor U16217 (N_16217,N_13826,N_13115);
xor U16218 (N_16218,N_11395,N_12450);
nor U16219 (N_16219,N_13401,N_12727);
xor U16220 (N_16220,N_14424,N_12670);
and U16221 (N_16221,N_13022,N_10016);
xor U16222 (N_16222,N_14498,N_12658);
xnor U16223 (N_16223,N_12492,N_14376);
nand U16224 (N_16224,N_11176,N_12794);
and U16225 (N_16225,N_12325,N_11748);
and U16226 (N_16226,N_10361,N_11592);
nor U16227 (N_16227,N_10111,N_12373);
and U16228 (N_16228,N_14362,N_10814);
and U16229 (N_16229,N_11950,N_12601);
nand U16230 (N_16230,N_14379,N_11615);
or U16231 (N_16231,N_11692,N_13076);
nand U16232 (N_16232,N_11962,N_14865);
or U16233 (N_16233,N_13232,N_12412);
nand U16234 (N_16234,N_12955,N_10310);
nor U16235 (N_16235,N_14916,N_13182);
and U16236 (N_16236,N_13783,N_10486);
nor U16237 (N_16237,N_14493,N_10922);
and U16238 (N_16238,N_12969,N_11924);
and U16239 (N_16239,N_13132,N_13223);
nor U16240 (N_16240,N_11957,N_13722);
nor U16241 (N_16241,N_10032,N_14338);
and U16242 (N_16242,N_10130,N_11831);
xnor U16243 (N_16243,N_12900,N_11470);
nor U16244 (N_16244,N_13589,N_12198);
nand U16245 (N_16245,N_11606,N_14499);
xor U16246 (N_16246,N_10549,N_12421);
xnor U16247 (N_16247,N_11414,N_10322);
or U16248 (N_16248,N_12331,N_11904);
xor U16249 (N_16249,N_13706,N_10596);
nor U16250 (N_16250,N_11863,N_11027);
nor U16251 (N_16251,N_13339,N_10302);
and U16252 (N_16252,N_12801,N_14645);
nor U16253 (N_16253,N_11717,N_14518);
and U16254 (N_16254,N_10678,N_14591);
nand U16255 (N_16255,N_14312,N_13806);
or U16256 (N_16256,N_12183,N_14960);
or U16257 (N_16257,N_14082,N_13282);
or U16258 (N_16258,N_13255,N_10061);
nand U16259 (N_16259,N_13431,N_13324);
nor U16260 (N_16260,N_10336,N_14030);
nor U16261 (N_16261,N_14707,N_12047);
xor U16262 (N_16262,N_10093,N_13450);
or U16263 (N_16263,N_14610,N_14299);
and U16264 (N_16264,N_14844,N_13329);
and U16265 (N_16265,N_10966,N_12759);
xor U16266 (N_16266,N_14913,N_13924);
nor U16267 (N_16267,N_12326,N_11883);
xor U16268 (N_16268,N_13087,N_13269);
nor U16269 (N_16269,N_14459,N_14659);
nor U16270 (N_16270,N_14480,N_11713);
nor U16271 (N_16271,N_13001,N_12432);
nand U16272 (N_16272,N_12564,N_13067);
xor U16273 (N_16273,N_12221,N_10559);
or U16274 (N_16274,N_11499,N_13628);
nand U16275 (N_16275,N_14168,N_10466);
nor U16276 (N_16276,N_10493,N_10421);
and U16277 (N_16277,N_11025,N_12072);
and U16278 (N_16278,N_11530,N_14373);
or U16279 (N_16279,N_12768,N_14282);
nor U16280 (N_16280,N_10054,N_11037);
xnor U16281 (N_16281,N_11964,N_10501);
or U16282 (N_16282,N_12517,N_11816);
xnor U16283 (N_16283,N_12286,N_14285);
or U16284 (N_16284,N_14626,N_12580);
nand U16285 (N_16285,N_12378,N_14126);
or U16286 (N_16286,N_11503,N_12112);
and U16287 (N_16287,N_14815,N_11356);
xnor U16288 (N_16288,N_13208,N_12561);
nand U16289 (N_16289,N_13525,N_13110);
and U16290 (N_16290,N_10368,N_12147);
nor U16291 (N_16291,N_10530,N_13950);
nor U16292 (N_16292,N_10372,N_13670);
xor U16293 (N_16293,N_14704,N_10067);
and U16294 (N_16294,N_11647,N_12208);
nor U16295 (N_16295,N_14598,N_10713);
nor U16296 (N_16296,N_13405,N_14284);
xor U16297 (N_16297,N_12267,N_13965);
and U16298 (N_16298,N_14743,N_14624);
and U16299 (N_16299,N_10364,N_11113);
nand U16300 (N_16300,N_12157,N_14984);
nor U16301 (N_16301,N_11604,N_14940);
xnor U16302 (N_16302,N_13162,N_12551);
and U16303 (N_16303,N_14371,N_12375);
nand U16304 (N_16304,N_10481,N_12731);
xnor U16305 (N_16305,N_10971,N_13570);
nor U16306 (N_16306,N_12574,N_13575);
or U16307 (N_16307,N_13740,N_10813);
or U16308 (N_16308,N_14446,N_13845);
nand U16309 (N_16309,N_12719,N_14196);
xor U16310 (N_16310,N_12917,N_12453);
and U16311 (N_16311,N_10218,N_13993);
and U16312 (N_16312,N_11703,N_14501);
xnor U16313 (N_16313,N_14823,N_14104);
nor U16314 (N_16314,N_11282,N_11137);
and U16315 (N_16315,N_13037,N_13218);
xor U16316 (N_16316,N_10685,N_10416);
and U16317 (N_16317,N_10938,N_11259);
and U16318 (N_16318,N_10295,N_13897);
nand U16319 (N_16319,N_10024,N_11227);
or U16320 (N_16320,N_10974,N_13301);
nand U16321 (N_16321,N_13966,N_13327);
nor U16322 (N_16322,N_11232,N_12870);
and U16323 (N_16323,N_10141,N_12686);
and U16324 (N_16324,N_11305,N_12806);
nand U16325 (N_16325,N_11173,N_13566);
xor U16326 (N_16326,N_10323,N_12563);
and U16327 (N_16327,N_14549,N_10044);
nand U16328 (N_16328,N_12027,N_14763);
or U16329 (N_16329,N_13756,N_11907);
nor U16330 (N_16330,N_11614,N_13582);
nor U16331 (N_16331,N_12336,N_14473);
nor U16332 (N_16332,N_13451,N_12753);
and U16333 (N_16333,N_13112,N_13958);
nand U16334 (N_16334,N_12359,N_10839);
xor U16335 (N_16335,N_14255,N_14303);
xnor U16336 (N_16336,N_10184,N_14627);
or U16337 (N_16337,N_13436,N_11345);
or U16338 (N_16338,N_13098,N_11646);
nor U16339 (N_16339,N_11878,N_11906);
and U16340 (N_16340,N_11549,N_13287);
nand U16341 (N_16341,N_13286,N_10249);
nand U16342 (N_16342,N_13114,N_12992);
nand U16343 (N_16343,N_10214,N_14695);
and U16344 (N_16344,N_13527,N_11956);
and U16345 (N_16345,N_10532,N_12161);
nand U16346 (N_16346,N_11099,N_11162);
or U16347 (N_16347,N_12200,N_13173);
nor U16348 (N_16348,N_11071,N_13325);
or U16349 (N_16349,N_14106,N_12164);
or U16350 (N_16350,N_12017,N_13940);
nand U16351 (N_16351,N_13272,N_10524);
nor U16352 (N_16352,N_14879,N_11156);
or U16353 (N_16353,N_11208,N_14320);
xnor U16354 (N_16354,N_11272,N_12546);
xor U16355 (N_16355,N_11015,N_13625);
or U16356 (N_16356,N_10197,N_13285);
and U16357 (N_16357,N_10630,N_13038);
and U16358 (N_16358,N_10480,N_11379);
or U16359 (N_16359,N_13660,N_11899);
or U16360 (N_16360,N_12196,N_11339);
or U16361 (N_16361,N_12624,N_11494);
nor U16362 (N_16362,N_10732,N_10534);
nand U16363 (N_16363,N_12694,N_11498);
nand U16364 (N_16364,N_12990,N_10284);
and U16365 (N_16365,N_14873,N_12778);
or U16366 (N_16366,N_14943,N_14447);
nand U16367 (N_16367,N_11194,N_10019);
or U16368 (N_16368,N_12512,N_14665);
xor U16369 (N_16369,N_14725,N_13879);
nor U16370 (N_16370,N_12346,N_10993);
or U16371 (N_16371,N_13528,N_11684);
and U16372 (N_16372,N_12202,N_14028);
nand U16373 (N_16373,N_11455,N_14745);
and U16374 (N_16374,N_13945,N_12028);
nand U16375 (N_16375,N_10158,N_14165);
and U16376 (N_16376,N_11810,N_10167);
or U16377 (N_16377,N_13189,N_11377);
nand U16378 (N_16378,N_13383,N_10944);
and U16379 (N_16379,N_10415,N_13236);
nand U16380 (N_16380,N_12455,N_13305);
xnor U16381 (N_16381,N_13788,N_14840);
xor U16382 (N_16382,N_10031,N_12446);
nor U16383 (N_16383,N_12162,N_13093);
xnor U16384 (N_16384,N_14952,N_10401);
xor U16385 (N_16385,N_13616,N_14340);
and U16386 (N_16386,N_13836,N_12962);
nor U16387 (N_16387,N_10514,N_11575);
xnor U16388 (N_16388,N_13726,N_12987);
and U16389 (N_16389,N_14623,N_14024);
nor U16390 (N_16390,N_12573,N_12777);
nand U16391 (N_16391,N_14837,N_13244);
nand U16392 (N_16392,N_14795,N_12849);
xnor U16393 (N_16393,N_14055,N_13177);
nand U16394 (N_16394,N_11560,N_11468);
xor U16395 (N_16395,N_14741,N_12111);
nor U16396 (N_16396,N_10945,N_11774);
nor U16397 (N_16397,N_10634,N_12064);
nor U16398 (N_16398,N_11231,N_11791);
nand U16399 (N_16399,N_12006,N_13779);
nand U16400 (N_16400,N_10043,N_11542);
nor U16401 (N_16401,N_10050,N_13963);
or U16402 (N_16402,N_11983,N_10012);
xor U16403 (N_16403,N_11955,N_14449);
nor U16404 (N_16404,N_14224,N_11807);
nor U16405 (N_16405,N_14176,N_10393);
and U16406 (N_16406,N_11534,N_10523);
and U16407 (N_16407,N_10306,N_14400);
and U16408 (N_16408,N_12816,N_10646);
and U16409 (N_16409,N_14080,N_13377);
xor U16410 (N_16410,N_14296,N_14044);
xnor U16411 (N_16411,N_10469,N_12533);
nor U16412 (N_16412,N_12804,N_11635);
and U16413 (N_16413,N_11325,N_14166);
nor U16414 (N_16414,N_14337,N_13443);
and U16415 (N_16415,N_11048,N_12693);
or U16416 (N_16416,N_10181,N_11686);
xor U16417 (N_16417,N_12396,N_12899);
or U16418 (N_16418,N_14254,N_10657);
and U16419 (N_16419,N_13127,N_10139);
or U16420 (N_16420,N_11311,N_10022);
nor U16421 (N_16421,N_10319,N_12931);
xnor U16422 (N_16422,N_12548,N_12102);
or U16423 (N_16423,N_11204,N_13937);
and U16424 (N_16424,N_11409,N_13188);
nand U16425 (N_16425,N_10027,N_13544);
and U16426 (N_16426,N_10369,N_11749);
nor U16427 (N_16427,N_11951,N_14219);
or U16428 (N_16428,N_12436,N_10828);
and U16429 (N_16429,N_14061,N_13797);
nand U16430 (N_16430,N_11623,N_14412);
nand U16431 (N_16431,N_12390,N_14500);
and U16432 (N_16432,N_12019,N_13179);
xnor U16433 (N_16433,N_14425,N_12940);
and U16434 (N_16434,N_12774,N_11676);
xnor U16435 (N_16435,N_14710,N_12910);
or U16436 (N_16436,N_14834,N_10281);
xnor U16437 (N_16437,N_13766,N_14066);
and U16438 (N_16438,N_13564,N_13467);
or U16439 (N_16439,N_13017,N_11856);
or U16440 (N_16440,N_13832,N_11023);
or U16441 (N_16441,N_12893,N_14038);
and U16442 (N_16442,N_10462,N_13948);
nor U16443 (N_16443,N_13992,N_14117);
nand U16444 (N_16444,N_12922,N_10170);
or U16445 (N_16445,N_12073,N_12437);
nand U16446 (N_16446,N_13535,N_14767);
nand U16447 (N_16447,N_14920,N_13708);
xnor U16448 (N_16448,N_14307,N_12150);
or U16449 (N_16449,N_13753,N_14616);
and U16450 (N_16450,N_11343,N_14845);
xnor U16451 (N_16451,N_10576,N_14129);
or U16452 (N_16452,N_13979,N_11702);
xor U16453 (N_16453,N_12048,N_14436);
nand U16454 (N_16454,N_11312,N_10844);
and U16455 (N_16455,N_10675,N_13291);
xnor U16456 (N_16456,N_11462,N_13379);
and U16457 (N_16457,N_14680,N_12675);
xor U16458 (N_16458,N_11823,N_12090);
xor U16459 (N_16459,N_14525,N_10109);
nor U16460 (N_16460,N_13890,N_12850);
nand U16461 (N_16461,N_10494,N_12484);
or U16462 (N_16462,N_12964,N_13813);
nand U16463 (N_16463,N_12576,N_14225);
and U16464 (N_16464,N_11437,N_13815);
xnor U16465 (N_16465,N_13977,N_10662);
nor U16466 (N_16466,N_14755,N_13142);
nor U16467 (N_16467,N_11469,N_14709);
nand U16468 (N_16468,N_11317,N_10060);
xnor U16469 (N_16469,N_10850,N_12706);
nor U16470 (N_16470,N_14169,N_11293);
nor U16471 (N_16471,N_12137,N_14481);
xnor U16472 (N_16472,N_11709,N_10760);
nand U16473 (N_16473,N_11509,N_12848);
nor U16474 (N_16474,N_12718,N_14378);
or U16475 (N_16475,N_10366,N_14982);
xor U16476 (N_16476,N_14759,N_12193);
nand U16477 (N_16477,N_11358,N_12951);
nand U16478 (N_16478,N_13194,N_12620);
or U16479 (N_16479,N_13991,N_13728);
or U16480 (N_16480,N_10745,N_11118);
and U16481 (N_16481,N_13590,N_10619);
and U16482 (N_16482,N_12444,N_13871);
and U16483 (N_16483,N_13886,N_12989);
nand U16484 (N_16484,N_13829,N_14849);
and U16485 (N_16485,N_14100,N_12846);
nand U16486 (N_16486,N_11714,N_12983);
xor U16487 (N_16487,N_11552,N_13027);
or U16488 (N_16488,N_11246,N_14820);
xor U16489 (N_16489,N_10498,N_14262);
nor U16490 (N_16490,N_11586,N_13241);
nor U16491 (N_16491,N_12886,N_12477);
nor U16492 (N_16492,N_14457,N_10178);
and U16493 (N_16493,N_10313,N_14398);
or U16494 (N_16494,N_11765,N_11300);
xor U16495 (N_16495,N_14988,N_12076);
nor U16496 (N_16496,N_14637,N_14653);
or U16497 (N_16497,N_14124,N_12398);
or U16498 (N_16498,N_13896,N_13483);
xor U16499 (N_16499,N_10413,N_12016);
nor U16500 (N_16500,N_10099,N_14485);
and U16501 (N_16501,N_14465,N_14832);
xnor U16502 (N_16502,N_10009,N_10341);
xnor U16503 (N_16503,N_11196,N_12040);
or U16504 (N_16504,N_11515,N_11042);
nand U16505 (N_16505,N_12283,N_11981);
nor U16506 (N_16506,N_14579,N_11938);
and U16507 (N_16507,N_14866,N_11053);
xor U16508 (N_16508,N_13748,N_14352);
or U16509 (N_16509,N_12739,N_10452);
and U16510 (N_16510,N_12973,N_10437);
xor U16511 (N_16511,N_12474,N_13512);
nor U16512 (N_16512,N_11631,N_13626);
and U16513 (N_16513,N_12120,N_14324);
nor U16514 (N_16514,N_11095,N_11802);
xor U16515 (N_16515,N_12294,N_12454);
and U16516 (N_16516,N_14019,N_11868);
or U16517 (N_16517,N_12254,N_10512);
or U16518 (N_16518,N_12856,N_14566);
and U16519 (N_16519,N_13298,N_12089);
xnor U16520 (N_16520,N_11884,N_14387);
and U16521 (N_16521,N_12457,N_13820);
or U16522 (N_16522,N_14069,N_13768);
nor U16523 (N_16523,N_14428,N_11845);
nor U16524 (N_16524,N_14609,N_14699);
nand U16525 (N_16525,N_12211,N_13227);
or U16526 (N_16526,N_14164,N_11415);
nor U16527 (N_16527,N_10915,N_10810);
nor U16528 (N_16528,N_12329,N_12873);
or U16529 (N_16529,N_10836,N_10086);
nand U16530 (N_16530,N_12545,N_14267);
and U16531 (N_16531,N_10912,N_10824);
or U16532 (N_16532,N_10330,N_14135);
nand U16533 (N_16533,N_13306,N_11992);
and U16534 (N_16534,N_11449,N_13323);
or U16535 (N_16535,N_14519,N_10359);
and U16536 (N_16536,N_13254,N_10867);
or U16537 (N_16537,N_10717,N_12976);
xnor U16538 (N_16538,N_10126,N_12883);
or U16539 (N_16539,N_14000,N_10233);
nand U16540 (N_16540,N_14272,N_14870);
xor U16541 (N_16541,N_14863,N_13827);
nor U16542 (N_16542,N_14084,N_12051);
xor U16543 (N_16543,N_11119,N_12403);
nor U16544 (N_16544,N_10529,N_11013);
and U16545 (N_16545,N_12292,N_13168);
and U16546 (N_16546,N_14293,N_14288);
nor U16547 (N_16547,N_14309,N_10658);
xnor U16548 (N_16548,N_10460,N_11388);
nand U16549 (N_16549,N_12681,N_13097);
nand U16550 (N_16550,N_12116,N_10316);
nand U16551 (N_16551,N_11695,N_11655);
nand U16552 (N_16552,N_14682,N_14631);
nor U16553 (N_16553,N_12275,N_13058);
xnor U16554 (N_16554,N_10703,N_11570);
or U16555 (N_16555,N_13083,N_14151);
or U16556 (N_16556,N_14203,N_12176);
or U16557 (N_16557,N_14221,N_12622);
or U16558 (N_16558,N_10371,N_12695);
or U16559 (N_16559,N_13790,N_14573);
and U16560 (N_16560,N_11908,N_11587);
nand U16561 (N_16561,N_14696,N_14576);
and U16562 (N_16562,N_11794,N_11131);
or U16563 (N_16563,N_10004,N_10247);
and U16564 (N_16564,N_12243,N_13122);
xnor U16565 (N_16565,N_14758,N_13200);
and U16566 (N_16566,N_10242,N_14615);
xor U16567 (N_16567,N_12151,N_14545);
and U16568 (N_16568,N_10426,N_12407);
nor U16569 (N_16569,N_14076,N_14405);
xnor U16570 (N_16570,N_12109,N_14047);
and U16571 (N_16571,N_10122,N_12497);
nand U16572 (N_16572,N_14364,N_14287);
and U16573 (N_16573,N_13381,N_10229);
nand U16574 (N_16574,N_11671,N_10380);
nor U16575 (N_16575,N_13052,N_11046);
nor U16576 (N_16576,N_11417,N_10028);
nor U16577 (N_16577,N_10835,N_11225);
xnor U16578 (N_16578,N_11433,N_14451);
xnor U16579 (N_16579,N_13134,N_11496);
or U16580 (N_16580,N_10566,N_14636);
or U16581 (N_16581,N_13283,N_10633);
nand U16582 (N_16582,N_11110,N_10283);
xor U16583 (N_16583,N_10123,N_11517);
and U16584 (N_16584,N_13995,N_11057);
xor U16585 (N_16585,N_14572,N_14611);
nor U16586 (N_16586,N_11144,N_14056);
xor U16587 (N_16587,N_12451,N_11022);
nand U16588 (N_16588,N_13850,N_12766);
nand U16589 (N_16589,N_13532,N_14548);
nand U16590 (N_16590,N_13961,N_11597);
nor U16591 (N_16591,N_10865,N_13537);
nand U16592 (N_16592,N_11341,N_14095);
and U16593 (N_16593,N_13417,N_13624);
and U16594 (N_16594,N_11653,N_13869);
xor U16595 (N_16595,N_13817,N_10586);
nor U16596 (N_16596,N_10736,N_13573);
nand U16597 (N_16597,N_14887,N_14814);
and U16598 (N_16598,N_14029,N_11594);
or U16599 (N_16599,N_13198,N_14114);
xnor U16600 (N_16600,N_11247,N_14980);
nor U16601 (N_16601,N_11795,N_11876);
and U16602 (N_16602,N_12499,N_11581);
nor U16603 (N_16603,N_11812,N_13461);
and U16604 (N_16604,N_13279,N_12293);
nand U16605 (N_16605,N_12581,N_13249);
and U16606 (N_16606,N_14180,N_10558);
nor U16607 (N_16607,N_11970,N_13707);
nor U16608 (N_16608,N_14657,N_11585);
and U16609 (N_16609,N_12520,N_14600);
nor U16610 (N_16610,N_14458,N_11576);
xnor U16611 (N_16611,N_10985,N_11763);
xnor U16612 (N_16612,N_11504,N_13754);
xor U16613 (N_16613,N_13824,N_10661);
or U16614 (N_16614,N_10389,N_12101);
and U16615 (N_16615,N_13387,N_11937);
nand U16616 (N_16616,N_14690,N_12610);
and U16617 (N_16617,N_14543,N_11483);
or U16618 (N_16618,N_10454,N_11328);
nand U16619 (N_16619,N_11167,N_12233);
and U16620 (N_16620,N_13674,N_13420);
nor U16621 (N_16621,N_12984,N_12105);
nor U16622 (N_16622,N_13760,N_11326);
and U16623 (N_16623,N_14607,N_12651);
nand U16624 (N_16624,N_12052,N_12071);
nor U16625 (N_16625,N_12411,N_12783);
nor U16626 (N_16626,N_11882,N_10519);
nor U16627 (N_16627,N_14946,N_14107);
and U16628 (N_16628,N_11457,N_10495);
nand U16629 (N_16629,N_10015,N_12805);
nor U16630 (N_16630,N_13712,N_12472);
xor U16631 (N_16631,N_14538,N_11353);
nand U16632 (N_16632,N_12635,N_14535);
nand U16633 (N_16633,N_13929,N_11207);
and U16634 (N_16634,N_11888,N_12148);
nand U16635 (N_16635,N_13084,N_10411);
and U16636 (N_16636,N_10764,N_13215);
nand U16637 (N_16637,N_14116,N_13684);
and U16638 (N_16638,N_14111,N_13884);
xor U16639 (N_16639,N_12889,N_11838);
nor U16640 (N_16640,N_12401,N_14523);
or U16641 (N_16641,N_11566,N_12934);
or U16642 (N_16642,N_12353,N_14783);
nor U16643 (N_16643,N_14463,N_11634);
and U16644 (N_16644,N_12288,N_12459);
nor U16645 (N_16645,N_11205,N_13678);
and U16646 (N_16646,N_14867,N_13154);
nor U16647 (N_16647,N_10073,N_12795);
nand U16648 (N_16648,N_13021,N_11694);
xor U16649 (N_16649,N_10277,N_12123);
xnor U16650 (N_16650,N_11367,N_10952);
and U16651 (N_16651,N_14553,N_13470);
nand U16652 (N_16652,N_10216,N_13237);
and U16653 (N_16653,N_12278,N_11301);
nor U16654 (N_16654,N_13771,N_12709);
nor U16655 (N_16655,N_13382,N_10852);
xor U16656 (N_16656,N_11629,N_14083);
or U16657 (N_16657,N_10358,N_11754);
nor U16658 (N_16658,N_13547,N_12648);
or U16659 (N_16659,N_14847,N_12328);
xnor U16660 (N_16660,N_13000,N_14805);
nand U16661 (N_16661,N_12677,N_10461);
nand U16662 (N_16662,N_14970,N_11885);
nor U16663 (N_16663,N_11060,N_13394);
xor U16664 (N_16664,N_12566,N_13540);
xor U16665 (N_16665,N_12268,N_10579);
and U16666 (N_16666,N_10288,N_12843);
nand U16667 (N_16667,N_10124,N_12671);
nand U16668 (N_16668,N_13724,N_13146);
xor U16669 (N_16669,N_12238,N_13505);
xor U16670 (N_16670,N_12659,N_11693);
or U16671 (N_16671,N_11781,N_12628);
nor U16672 (N_16672,N_13457,N_14557);
or U16673 (N_16673,N_12588,N_13685);
nand U16674 (N_16674,N_14074,N_11648);
or U16675 (N_16675,N_11273,N_13762);
xor U16676 (N_16676,N_12921,N_13145);
xor U16677 (N_16677,N_10239,N_11084);
and U16678 (N_16678,N_12460,N_11952);
nor U16679 (N_16679,N_11599,N_14317);
nand U16680 (N_16680,N_12049,N_12830);
and U16681 (N_16681,N_14559,N_10394);
nor U16682 (N_16682,N_12902,N_12755);
nand U16683 (N_16683,N_14440,N_13120);
nor U16684 (N_16684,N_14774,N_11390);
and U16685 (N_16685,N_12367,N_13474);
xor U16686 (N_16686,N_10203,N_11410);
xor U16687 (N_16687,N_14918,N_13238);
nor U16688 (N_16688,N_13711,N_13455);
or U16689 (N_16689,N_14315,N_13452);
xor U16690 (N_16690,N_12744,N_11416);
and U16691 (N_16691,N_14018,N_11159);
nand U16692 (N_16692,N_11524,N_10988);
and U16693 (N_16693,N_13644,N_11286);
nand U16694 (N_16694,N_13508,N_10626);
nor U16695 (N_16695,N_11609,N_14264);
and U16696 (N_16696,N_11636,N_10504);
xor U16697 (N_16697,N_14788,N_11742);
or U16698 (N_16698,N_10449,N_13882);
xnor U16699 (N_16699,N_14460,N_10992);
xor U16700 (N_16700,N_13495,N_10442);
nand U16701 (N_16701,N_12853,N_11922);
nor U16702 (N_16702,N_13032,N_14329);
and U16703 (N_16703,N_11849,N_14630);
nand U16704 (N_16704,N_10913,N_12798);
and U16705 (N_16705,N_10904,N_13878);
nand U16706 (N_16706,N_11826,N_12441);
xnor U16707 (N_16707,N_14901,N_10290);
or U16708 (N_16708,N_10812,N_12280);
and U16709 (N_16709,N_11681,N_13368);
or U16710 (N_16710,N_11020,N_13881);
or U16711 (N_16711,N_11454,N_13108);
xnor U16712 (N_16712,N_10266,N_14567);
xor U16713 (N_16713,N_12944,N_13488);
nand U16714 (N_16714,N_10107,N_14722);
nor U16715 (N_16715,N_10227,N_14762);
nor U16716 (N_16716,N_11180,N_10095);
and U16717 (N_16717,N_10733,N_13251);
xor U16718 (N_16718,N_12611,N_14629);
or U16719 (N_16719,N_13116,N_12823);
nand U16720 (N_16720,N_10327,N_14187);
xor U16721 (N_16721,N_12232,N_11788);
or U16722 (N_16722,N_12757,N_10709);
and U16723 (N_16723,N_14192,N_10001);
nor U16724 (N_16724,N_10240,N_13747);
nand U16725 (N_16725,N_12613,N_12368);
nor U16726 (N_16726,N_10638,N_11900);
nor U16727 (N_16727,N_13978,N_14716);
nor U16728 (N_16728,N_14283,N_13437);
and U16729 (N_16729,N_12449,N_13705);
and U16730 (N_16730,N_13999,N_10741);
nand U16731 (N_16731,N_10554,N_11512);
nor U16732 (N_16732,N_11418,N_12720);
or U16733 (N_16733,N_10759,N_14275);
and U16734 (N_16734,N_13702,N_13453);
or U16735 (N_16735,N_12408,N_10357);
or U16736 (N_16736,N_14479,N_11065);
or U16737 (N_16737,N_12075,N_14156);
nand U16738 (N_16738,N_12923,N_10152);
nand U16739 (N_16739,N_11711,N_12287);
or U16740 (N_16740,N_14590,N_13148);
xor U16741 (N_16741,N_13974,N_13092);
xnor U16742 (N_16742,N_12054,N_11532);
and U16743 (N_16743,N_10407,N_14582);
or U16744 (N_16744,N_11659,N_11903);
and U16745 (N_16745,N_11879,N_14208);
nand U16746 (N_16746,N_12227,N_11004);
or U16747 (N_16747,N_11224,N_13230);
nand U16748 (N_16748,N_13872,N_11916);
xnor U16749 (N_16749,N_11024,N_11348);
xor U16750 (N_16750,N_14027,N_11111);
xor U16751 (N_16751,N_11473,N_12936);
or U16752 (N_16752,N_11616,N_12608);
nor U16753 (N_16753,N_11475,N_14587);
nand U16754 (N_16754,N_11387,N_11786);
nand U16755 (N_16755,N_11493,N_12776);
and U16756 (N_16756,N_12002,N_14422);
nor U16757 (N_16757,N_10309,N_13271);
nor U16758 (N_16758,N_12440,N_13892);
xnor U16759 (N_16759,N_11644,N_14751);
and U16760 (N_16760,N_10672,N_12033);
and U16761 (N_16761,N_12388,N_14541);
or U16762 (N_16762,N_12140,N_12799);
xnor U16763 (N_16763,N_10598,N_13736);
or U16764 (N_16764,N_11673,N_10894);
or U16765 (N_16765,N_14547,N_14936);
nor U16766 (N_16766,N_13020,N_14994);
and U16767 (N_16767,N_13319,N_12241);
or U16768 (N_16768,N_13442,N_12100);
xnor U16769 (N_16769,N_11096,N_14953);
nand U16770 (N_16770,N_11160,N_10221);
xnor U16771 (N_16771,N_12696,N_13260);
or U16772 (N_16772,N_10853,N_14195);
xnor U16773 (N_16773,N_14546,N_14252);
xnor U16774 (N_16774,N_10397,N_11327);
nor U16775 (N_16775,N_11047,N_13916);
nand U16776 (N_16776,N_10026,N_11000);
and U16777 (N_16777,N_14057,N_12025);
nor U16778 (N_16778,N_10544,N_14925);
and U16779 (N_16779,N_11351,N_10935);
and U16780 (N_16780,N_14912,N_13930);
xor U16781 (N_16781,N_11801,N_13737);
nor U16782 (N_16782,N_11850,N_14495);
and U16783 (N_16783,N_12890,N_11723);
xor U16784 (N_16784,N_13477,N_14051);
nor U16785 (N_16785,N_12225,N_11044);
and U16786 (N_16786,N_12145,N_13423);
nand U16787 (N_16787,N_12341,N_10145);
or U16788 (N_16788,N_12009,N_13019);
xnor U16789 (N_16789,N_10003,N_10146);
nor U16790 (N_16790,N_14951,N_12487);
xnor U16791 (N_16791,N_13668,N_10871);
nor U16792 (N_16792,N_14654,N_13786);
and U16793 (N_16793,N_11886,N_14625);
xor U16794 (N_16794,N_14308,N_12274);
nand U16795 (N_16795,N_10023,N_13672);
nor U16796 (N_16796,N_11148,N_14735);
nor U16797 (N_16797,N_14895,N_13764);
and U16798 (N_16798,N_10726,N_13557);
or U16799 (N_16799,N_14435,N_14088);
nor U16800 (N_16800,N_13778,N_14596);
nor U16801 (N_16801,N_11360,N_11986);
or U16802 (N_16802,N_12442,N_11589);
and U16803 (N_16803,N_10424,N_12898);
and U16804 (N_16804,N_12514,N_11990);
nor U16805 (N_16805,N_10731,N_14757);
nand U16806 (N_16806,N_13691,N_12270);
xnor U16807 (N_16807,N_12916,N_13683);
nor U16808 (N_16808,N_10647,N_11642);
or U16809 (N_16809,N_12919,N_12832);
and U16810 (N_16810,N_13562,N_12542);
or U16811 (N_16811,N_10917,N_12365);
xor U16812 (N_16812,N_12134,N_13579);
and U16813 (N_16813,N_11138,N_14385);
and U16814 (N_16814,N_10485,N_13409);
nand U16815 (N_16815,N_14131,N_10503);
and U16816 (N_16816,N_11949,N_14319);
nand U16817 (N_16817,N_11687,N_12713);
nand U16818 (N_16818,N_14780,N_11089);
xor U16819 (N_16819,N_10459,N_14243);
nor U16820 (N_16820,N_12865,N_10453);
nand U16821 (N_16821,N_12619,N_12063);
nor U16822 (N_16822,N_12822,N_13347);
xor U16823 (N_16823,N_10116,N_14864);
xnor U16824 (N_16824,N_13563,N_13439);
nor U16825 (N_16825,N_14964,N_10650);
nor U16826 (N_16826,N_11556,N_12271);
nand U16827 (N_16827,N_14806,N_14017);
nand U16828 (N_16828,N_10572,N_10604);
nand U16829 (N_16829,N_14327,N_13613);
or U16830 (N_16830,N_10430,N_14937);
nand U16831 (N_16831,N_14713,N_10640);
or U16832 (N_16832,N_12175,N_11966);
nand U16833 (N_16833,N_14369,N_10927);
or U16834 (N_16834,N_11832,N_11972);
and U16835 (N_16835,N_12645,N_10080);
and U16836 (N_16836,N_13049,N_14685);
and U16837 (N_16837,N_14392,N_10541);
or U16838 (N_16838,N_14419,N_14060);
nor U16839 (N_16839,N_14001,N_10317);
nand U16840 (N_16840,N_14409,N_13490);
and U16841 (N_16841,N_10881,N_12425);
and U16842 (N_16842,N_11203,N_10193);
xnor U16843 (N_16843,N_13734,N_14647);
nor U16844 (N_16844,N_11394,N_12963);
nand U16845 (N_16845,N_12756,N_13359);
or U16846 (N_16846,N_11821,N_13586);
xor U16847 (N_16847,N_10406,N_10508);
or U16848 (N_16848,N_14738,N_10223);
or U16849 (N_16849,N_12486,N_12716);
or U16850 (N_16850,N_12575,N_11691);
and U16851 (N_16851,N_13611,N_12510);
and U16852 (N_16852,N_14408,N_12952);
xnor U16853 (N_16853,N_11361,N_12769);
xor U16854 (N_16854,N_10774,N_14050);
xor U16855 (N_16855,N_10893,N_14108);
and U16856 (N_16856,N_13523,N_14382);
or U16857 (N_16857,N_12586,N_14214);
xor U16858 (N_16858,N_13160,N_13250);
xor U16859 (N_16859,N_11200,N_10616);
and U16860 (N_16860,N_12876,N_14510);
nor U16861 (N_16861,N_11255,N_10467);
xor U16862 (N_16862,N_12285,N_14851);
nor U16863 (N_16863,N_13315,N_14402);
xnor U16864 (N_16864,N_12171,N_10084);
xnor U16865 (N_16865,N_12742,N_13042);
and U16866 (N_16866,N_13597,N_14306);
nand U16867 (N_16867,N_13642,N_11881);
nor U16868 (N_16868,N_10066,N_10659);
or U16869 (N_16869,N_10057,N_10456);
nand U16870 (N_16870,N_13060,N_11427);
or U16871 (N_16871,N_10418,N_13184);
nand U16872 (N_16872,N_11215,N_11573);
nor U16873 (N_16873,N_14052,N_10750);
and U16874 (N_16874,N_13799,N_13228);
xor U16875 (N_16875,N_12941,N_10925);
or U16876 (N_16876,N_12614,N_10588);
xor U16877 (N_16877,N_11120,N_14979);
and U16878 (N_16878,N_14737,N_11638);
xnor U16879 (N_16879,N_12351,N_12473);
xor U16880 (N_16880,N_11736,N_14702);
xor U16881 (N_16881,N_10196,N_11557);
nand U16882 (N_16882,N_14634,N_12008);
and U16883 (N_16883,N_12847,N_10772);
and U16884 (N_16884,N_12965,N_13700);
and U16885 (N_16885,N_14949,N_14749);
nor U16886 (N_16886,N_13284,N_10928);
xnor U16887 (N_16887,N_10264,N_14941);
xor U16888 (N_16888,N_14404,N_12660);
nand U16889 (N_16889,N_10210,N_13261);
and U16890 (N_16890,N_12448,N_11796);
nor U16891 (N_16891,N_14064,N_11919);
and U16892 (N_16892,N_11382,N_12385);
nand U16893 (N_16893,N_12142,N_13029);
or U16894 (N_16894,N_14983,N_11362);
xor U16895 (N_16895,N_14551,N_12524);
xnor U16896 (N_16896,N_13503,N_13909);
nor U16897 (N_16897,N_13962,N_11197);
nor U16898 (N_16898,N_12821,N_10360);
nor U16899 (N_16899,N_10014,N_11583);
nand U16900 (N_16900,N_11514,N_12495);
nand U16901 (N_16901,N_10378,N_13524);
nor U16902 (N_16902,N_11965,N_14438);
nor U16903 (N_16903,N_13641,N_12029);
nand U16904 (N_16904,N_10157,N_13345);
xor U16905 (N_16905,N_10870,N_11371);
or U16906 (N_16906,N_13542,N_14437);
and U16907 (N_16907,N_10237,N_14105);
nand U16908 (N_16908,N_13099,N_10431);
nand U16909 (N_16909,N_13313,N_10068);
and U16910 (N_16910,N_11988,N_11927);
nand U16911 (N_16911,N_10674,N_13499);
xnor U16912 (N_16912,N_14734,N_10273);
nor U16913 (N_16913,N_11719,N_11214);
nor U16914 (N_16914,N_11929,N_14842);
nand U16915 (N_16915,N_10025,N_11571);
xnor U16916 (N_16916,N_11151,N_10179);
and U16917 (N_16917,N_10995,N_12312);
nand U16918 (N_16918,N_11716,N_10771);
and U16919 (N_16919,N_10448,N_13378);
xor U16920 (N_16920,N_11750,N_11064);
or U16921 (N_16921,N_12958,N_10199);
nand U16922 (N_16922,N_14807,N_11595);
nor U16923 (N_16923,N_13984,N_11645);
xnor U16924 (N_16924,N_14189,N_13274);
and U16925 (N_16925,N_10391,N_10892);
xor U16926 (N_16926,N_14261,N_11287);
nand U16927 (N_16927,N_11446,N_10075);
nand U16928 (N_16928,N_11055,N_14731);
nand U16929 (N_16929,N_10642,N_10653);
xnor U16930 (N_16930,N_13043,N_10613);
or U16931 (N_16931,N_10300,N_13901);
or U16932 (N_16932,N_12355,N_13469);
nand U16933 (N_16933,N_11672,N_14929);
nor U16934 (N_16934,N_12633,N_14250);
nand U16935 (N_16935,N_10011,N_12729);
nand U16936 (N_16936,N_14906,N_10818);
nand U16937 (N_16937,N_14868,N_12672);
nand U16938 (N_16938,N_10789,N_11412);
nand U16939 (N_16939,N_11149,N_10320);
nand U16940 (N_16940,N_13091,N_12413);
nor U16941 (N_16941,N_12734,N_12903);
or U16942 (N_16942,N_11528,N_12496);
or U16943 (N_16943,N_13448,N_13943);
nand U16944 (N_16944,N_11322,N_12702);
or U16945 (N_16945,N_13201,N_13794);
or U16946 (N_16946,N_13011,N_10250);
or U16947 (N_16947,N_13561,N_12463);
and U16948 (N_16948,N_13113,N_10507);
nand U16949 (N_16949,N_12149,N_12097);
xor U16950 (N_16950,N_13050,N_10729);
or U16951 (N_16951,N_13266,N_12867);
xor U16952 (N_16952,N_13614,N_14821);
and U16953 (N_16953,N_14620,N_14663);
nand U16954 (N_16954,N_11590,N_10940);
xor U16955 (N_16955,N_11376,N_11701);
and U16956 (N_16956,N_11074,N_10312);
nor U16957 (N_16957,N_10719,N_10846);
nor U16958 (N_16958,N_11819,N_13981);
nand U16959 (N_16959,N_11588,N_10739);
nand U16960 (N_16960,N_10429,N_13934);
nor U16961 (N_16961,N_10136,N_14476);
and U16962 (N_16962,N_12410,N_10059);
nand U16963 (N_16963,N_10639,N_12093);
or U16964 (N_16964,N_14933,N_10723);
nor U16965 (N_16965,N_14978,N_14170);
or U16966 (N_16966,N_11877,N_14678);
and U16967 (N_16967,N_14341,N_13506);
nor U16968 (N_16968,N_13926,N_11947);
or U16969 (N_16969,N_14995,N_10830);
and U16970 (N_16970,N_13679,N_12523);
nand U16971 (N_16971,N_12697,N_12044);
nand U16972 (N_16972,N_11086,N_13273);
nor U16973 (N_16973,N_11190,N_13163);
nand U16974 (N_16974,N_10610,N_14491);
xor U16975 (N_16975,N_12625,N_11857);
and U16976 (N_16976,N_13192,N_11129);
or U16977 (N_16977,N_12086,N_13225);
and U16978 (N_16978,N_11333,N_11443);
nor U16979 (N_16979,N_12070,N_10112);
xor U16980 (N_16980,N_11887,N_10072);
and U16981 (N_16981,N_14177,N_14761);
nor U16982 (N_16982,N_10651,N_12023);
nor U16983 (N_16983,N_10815,N_10730);
xor U16984 (N_16984,N_13578,N_11370);
or U16985 (N_16985,N_11665,N_14813);
nor U16986 (N_16986,N_10943,N_11562);
nor U16987 (N_16987,N_14368,N_11705);
xor U16988 (N_16988,N_14771,N_12042);
nand U16989 (N_16989,N_11651,N_13340);
xnor U16990 (N_16990,N_13620,N_12554);
nor U16991 (N_16991,N_12792,N_11747);
nand U16992 (N_16992,N_14697,N_11624);
nor U16993 (N_16993,N_14886,N_11848);
and U16994 (N_16994,N_12377,N_14395);
nor U16995 (N_16995,N_13157,N_12266);
nor U16996 (N_16996,N_12332,N_10926);
xor U16997 (N_16997,N_12038,N_14360);
xor U16998 (N_16998,N_11600,N_14928);
xnor U16999 (N_16999,N_12187,N_12519);
xor U17000 (N_17000,N_12543,N_13663);
and U17001 (N_17001,N_12132,N_14924);
xnor U17002 (N_17002,N_12772,N_11482);
or U17003 (N_17003,N_10987,N_13671);
nor U17004 (N_17004,N_12895,N_11029);
and U17005 (N_17005,N_12616,N_10790);
nand U17006 (N_17006,N_11453,N_10506);
or U17007 (N_17007,N_10773,N_10536);
and U17008 (N_17008,N_12750,N_11772);
nor U17009 (N_17009,N_11323,N_11675);
and U17010 (N_17010,N_12785,N_13061);
and U17011 (N_17011,N_13056,N_10248);
nand U17012 (N_17012,N_12141,N_11432);
and U17013 (N_17013,N_13243,N_10259);
xor U17014 (N_17014,N_12154,N_14301);
nand U17015 (N_17015,N_11428,N_12345);
or U17016 (N_17016,N_11445,N_11511);
xnor U17017 (N_17017,N_11830,N_13478);
xnor U17018 (N_17018,N_12909,N_13222);
nand U17019 (N_17019,N_11028,N_13397);
nand U17020 (N_17020,N_10847,N_14586);
and U17021 (N_17021,N_10937,N_13973);
nand U17022 (N_17022,N_14687,N_13025);
nand U17023 (N_17023,N_12967,N_10127);
nor U17024 (N_17024,N_12059,N_12135);
and U17025 (N_17025,N_10905,N_12468);
nor U17026 (N_17026,N_14065,N_10548);
or U17027 (N_17027,N_12998,N_14686);
nor U17028 (N_17028,N_11393,N_11926);
or U17029 (N_17029,N_10959,N_13302);
nand U17030 (N_17030,N_13239,N_12593);
nand U17031 (N_17031,N_12349,N_13288);
or U17032 (N_17032,N_11930,N_11914);
or U17033 (N_17033,N_13731,N_10751);
nor U17034 (N_17034,N_13852,N_13167);
nor U17035 (N_17035,N_13051,N_12634);
and U17036 (N_17036,N_10611,N_12710);
and U17037 (N_17037,N_11270,N_12796);
and U17038 (N_17038,N_14384,N_12618);
xnor U17039 (N_17039,N_10929,N_12031);
nor U17040 (N_17040,N_13337,N_12037);
xnor U17041 (N_17041,N_12327,N_12700);
or U17042 (N_17042,N_12230,N_12323);
nand U17043 (N_17043,N_10715,N_10296);
nand U17044 (N_17044,N_14564,N_12084);
xnor U17045 (N_17045,N_12115,N_13399);
and U17046 (N_17046,N_11625,N_13696);
nor U17047 (N_17047,N_11380,N_13585);
nand U17048 (N_17048,N_14046,N_11546);
and U17049 (N_17049,N_12262,N_13634);
or U17050 (N_17050,N_13159,N_10580);
or U17051 (N_17051,N_12265,N_11226);
nand U17052 (N_17052,N_12205,N_10727);
nor U17053 (N_17053,N_12885,N_14772);
and U17054 (N_17054,N_10849,N_11352);
nand U17055 (N_17055,N_10225,N_12968);
nand U17056 (N_17056,N_10285,N_12194);
xnor U17057 (N_17057,N_12011,N_12650);
and U17058 (N_17058,N_10526,N_10100);
and U17059 (N_17059,N_13665,N_14397);
nor U17060 (N_17060,N_14618,N_10362);
xnor U17061 (N_17061,N_12340,N_13259);
or U17062 (N_17062,N_13612,N_10960);
xnor U17063 (N_17063,N_10605,N_13608);
and U17064 (N_17064,N_10522,N_12397);
nand U17065 (N_17065,N_11668,N_11313);
or U17066 (N_17066,N_10191,N_12245);
or U17067 (N_17067,N_11477,N_10791);
and U17068 (N_17068,N_12978,N_14265);
nor U17069 (N_17069,N_11413,N_12701);
and U17070 (N_17070,N_13040,N_11268);
nand U17071 (N_17071,N_12229,N_12604);
or U17072 (N_17072,N_11997,N_12582);
and U17073 (N_17073,N_14850,N_11082);
and U17074 (N_17074,N_10777,N_10688);
nor U17075 (N_17075,N_11630,N_13434);
and U17076 (N_17076,N_10805,N_14675);
or U17077 (N_17077,N_10144,N_10156);
and U17078 (N_17078,N_12203,N_14417);
or U17079 (N_17079,N_12074,N_11183);
and U17080 (N_17080,N_14119,N_11860);
nand U17081 (N_17081,N_11458,N_11078);
nand U17082 (N_17082,N_10308,N_12242);
nand U17083 (N_17083,N_13895,N_14965);
xnor U17084 (N_17084,N_11577,N_13550);
nor U17085 (N_17085,N_10410,N_13936);
and U17086 (N_17086,N_13687,N_14703);
xor U17087 (N_17087,N_13214,N_12864);
or U17088 (N_17088,N_11484,N_14348);
xnor U17089 (N_17089,N_10843,N_13800);
and U17090 (N_17090,N_14877,N_11222);
xnor U17091 (N_17091,N_14313,N_13009);
nor U17092 (N_17092,N_14464,N_14858);
nand U17093 (N_17093,N_11669,N_11733);
nor U17094 (N_17094,N_13602,N_11344);
nor U17095 (N_17095,N_11465,N_12746);
xor U17096 (N_17096,N_11201,N_14608);
nand U17097 (N_17097,N_10994,N_14560);
xor U17098 (N_17098,N_13281,N_11522);
xnor U17099 (N_17099,N_14245,N_12004);
or U17100 (N_17100,N_13418,N_12256);
and U17101 (N_17101,N_12842,N_13330);
xnor U17102 (N_17102,N_14475,N_10552);
and U17103 (N_17103,N_10497,N_12626);
and U17104 (N_17104,N_12918,N_14098);
xor U17105 (N_17105,N_11302,N_12954);
nor U17106 (N_17106,N_13819,N_10941);
nand U17107 (N_17107,N_11758,N_10743);
or U17108 (N_17108,N_11652,N_14003);
xor U17109 (N_17109,N_13210,N_13906);
or U17110 (N_17110,N_11732,N_12825);
or U17111 (N_17111,N_11187,N_13363);
xnor U17112 (N_17112,N_11720,N_12258);
nor U17113 (N_17113,N_10445,N_10104);
nand U17114 (N_17114,N_10488,N_10698);
xnor U17115 (N_17115,N_10119,N_12207);
nand U17116 (N_17116,N_13811,N_13767);
and U17117 (N_17117,N_11954,N_14580);
xor U17118 (N_17118,N_14792,N_11134);
nand U17119 (N_17119,N_10198,N_11280);
xnor U17120 (N_17120,N_13607,N_13667);
nor U17121 (N_17121,N_14804,N_11150);
or U17122 (N_17122,N_11520,N_11304);
and U17123 (N_17123,N_10051,N_14991);
xor U17124 (N_17124,N_13352,N_10356);
nor U17125 (N_17125,N_13675,N_10990);
xnor U17126 (N_17126,N_10094,N_14016);
nor U17127 (N_17127,N_11424,N_14198);
nand U17128 (N_17128,N_11040,N_10752);
xor U17129 (N_17129,N_10832,N_11003);
nor U17130 (N_17130,N_13444,N_14089);
or U17131 (N_17131,N_11523,N_14152);
xor U17132 (N_17132,N_10696,N_12465);
xnor U17133 (N_17133,N_13744,N_12311);
nor U17134 (N_17134,N_11108,N_12844);
nor U17135 (N_17135,N_11193,N_14413);
nor U17136 (N_17136,N_12525,N_12068);
nor U17137 (N_17137,N_14898,N_11122);
nor U17138 (N_17138,N_14532,N_14915);
nand U17139 (N_17139,N_11568,N_14536);
nand U17140 (N_17140,N_14606,N_11032);
or U17141 (N_17141,N_10138,N_11170);
or U17142 (N_17142,N_12539,N_13491);
nor U17143 (N_17143,N_10423,N_14922);
or U17144 (N_17144,N_11803,N_12122);
or U17145 (N_17145,N_11895,N_12240);
nor U17146 (N_17146,N_11953,N_10702);
nor U17147 (N_17147,N_11650,N_10222);
and U17148 (N_17148,N_14666,N_11425);
nand U17149 (N_17149,N_11439,N_10851);
nor U17150 (N_17150,N_14158,N_13015);
xnor U17151 (N_17151,N_10173,N_13502);
nor U17152 (N_17152,N_12735,N_10533);
xor U17153 (N_17153,N_11275,N_10597);
nand U17154 (N_17154,N_13598,N_12426);
nor U17155 (N_17155,N_11069,N_14520);
xnor U17156 (N_17156,N_13935,N_13773);
xor U17157 (N_17157,N_12464,N_12603);
and U17158 (N_17158,N_12077,N_10261);
or U17159 (N_17159,N_14740,N_10160);
and U17160 (N_17160,N_11767,N_12770);
or U17161 (N_17161,N_10254,N_11401);
nor U17162 (N_17162,N_13560,N_14414);
nor U17163 (N_17163,N_11680,N_12167);
and U17164 (N_17164,N_14822,N_14444);
nand U17165 (N_17165,N_12977,N_13818);
nor U17166 (N_17166,N_14489,N_14515);
or U17167 (N_17167,N_11329,N_10963);
nand U17168 (N_17168,N_14223,N_13949);
or U17169 (N_17169,N_11296,N_11944);
xor U17170 (N_17170,N_13459,N_12438);
and U17171 (N_17171,N_14268,N_11998);
or U17172 (N_17172,N_10381,N_12682);
and U17173 (N_17173,N_13622,N_12114);
nand U17174 (N_17174,N_13253,N_12152);
xor U17175 (N_17175,N_11500,N_13479);
and U17176 (N_17176,N_11062,N_11829);
or U17177 (N_17177,N_13860,N_12606);
nor U17178 (N_17178,N_14274,N_13584);
nor U17179 (N_17179,N_10492,N_13035);
or U17180 (N_17180,N_10212,N_14062);
or U17181 (N_17181,N_14658,N_14542);
nand U17182 (N_17182,N_14809,N_12565);
xor U17183 (N_17183,N_12684,N_12925);
nand U17184 (N_17184,N_11768,N_10822);
and U17185 (N_17185,N_10496,N_11385);
and U17186 (N_17186,N_13402,N_14640);
or U17187 (N_17187,N_11070,N_13089);
nor U17188 (N_17188,N_12945,N_11521);
or U17189 (N_17189,N_13275,N_12096);
nand U17190 (N_17190,N_14271,N_12600);
nor U17191 (N_17191,N_10230,N_11738);
nor U17192 (N_17192,N_14217,N_10954);
xnor U17193 (N_17193,N_11793,N_12872);
nor U17194 (N_17194,N_12439,N_11633);
nand U17195 (N_17195,N_12787,N_11731);
nand U17196 (N_17196,N_10412,N_14558);
nor U17197 (N_17197,N_11397,N_13848);
nor U17198 (N_17198,N_13951,N_14612);
or U17199 (N_17199,N_14619,N_12855);
and U17200 (N_17200,N_11284,N_14694);
or U17201 (N_17201,N_10176,N_10920);
or U17202 (N_17202,N_14673,N_13063);
xor U17203 (N_17203,N_10792,N_12419);
xor U17204 (N_17204,N_14585,N_12752);
and U17205 (N_17205,N_11420,N_14237);
xnor U17206 (N_17206,N_10478,N_13574);
nor U17207 (N_17207,N_13065,N_11248);
or U17208 (N_17208,N_13709,N_13471);
xnor U17209 (N_17209,N_14079,N_13496);
xnor U17210 (N_17210,N_13595,N_12138);
nand U17211 (N_17211,N_12428,N_11787);
nand U17212 (N_17212,N_10079,N_12482);
or U17213 (N_17213,N_14752,N_13217);
nor U17214 (N_17214,N_11012,N_10695);
or U17215 (N_17215,N_12932,N_10761);
or U17216 (N_17216,N_14242,N_14325);
and U17217 (N_17217,N_12255,N_13125);
nor U17218 (N_17218,N_12748,N_14012);
xor U17219 (N_17219,N_14651,N_10172);
and U17220 (N_17220,N_14829,N_14310);
and U17221 (N_17221,N_13933,N_13862);
xor U17222 (N_17222,N_11598,N_14482);
and U17223 (N_17223,N_13867,N_10035);
or U17224 (N_17224,N_12158,N_10587);
nand U17225 (N_17225,N_10500,N_11896);
and U17226 (N_17226,N_13694,N_11928);
or U17227 (N_17227,N_11100,N_10171);
or U17228 (N_17228,N_12986,N_10085);
and U17229 (N_17229,N_10924,N_12309);
nor U17230 (N_17230,N_14171,N_12733);
and U17231 (N_17231,N_13652,N_12877);
nand U17232 (N_17232,N_13180,N_10983);
nand U17233 (N_17233,N_10747,N_10593);
and U17234 (N_17234,N_12598,N_12722);
and U17235 (N_17235,N_13849,N_14578);
nor U17236 (N_17236,N_13796,N_14781);
nor U17237 (N_17237,N_13710,N_12469);
xor U17238 (N_17238,N_14349,N_11612);
and U17239 (N_17239,N_10234,N_12220);
and U17240 (N_17240,N_12567,N_10128);
and U17241 (N_17241,N_14753,N_12344);
xnor U17242 (N_17242,N_10236,N_13321);
nand U17243 (N_17243,N_10700,N_11913);
xor U17244 (N_17244,N_12215,N_14178);
nand U17245 (N_17245,N_12534,N_10606);
nand U17246 (N_17246,N_14025,N_14971);
and U17247 (N_17247,N_10348,N_12506);
and U17248 (N_17248,N_13717,N_14812);
nor U17249 (N_17249,N_13410,N_13697);
xnor U17250 (N_17250,N_14748,N_12935);
or U17251 (N_17251,N_11436,N_14882);
nand U17252 (N_17252,N_13549,N_11228);
and U17253 (N_17253,N_10048,N_12887);
nand U17254 (N_17254,N_14101,N_13593);
and U17255 (N_17255,N_10263,N_12572);
nor U17256 (N_17256,N_10087,N_10946);
and U17257 (N_17257,N_10540,N_11140);
nor U17258 (N_17258,N_12181,N_13765);
nor U17259 (N_17259,N_14174,N_13322);
xnor U17260 (N_17260,N_10823,N_12020);
and U17261 (N_17261,N_11038,N_10370);
nand U17262 (N_17262,N_14326,N_14790);
nor U17263 (N_17263,N_11174,N_12201);
or U17264 (N_17264,N_14522,N_11179);
or U17265 (N_17265,N_14355,N_11539);
nor U17266 (N_17266,N_13351,N_10857);
xor U17267 (N_17267,N_10977,N_14478);
nor U17268 (N_17268,N_11825,N_13855);
and U17269 (N_17269,N_11066,N_14236);
xor U17270 (N_17270,N_14259,N_10208);
and U17271 (N_17271,N_12000,N_12119);
or U17272 (N_17272,N_11797,N_13632);
nor U17273 (N_17273,N_14132,N_14794);
xor U17274 (N_17274,N_12623,N_11365);
and U17275 (N_17275,N_11550,N_11243);
nor U17276 (N_17276,N_10175,N_11827);
nor U17277 (N_17277,N_14973,N_11016);
nor U17278 (N_17278,N_14071,N_13012);
or U17279 (N_17279,N_11558,N_10232);
xnor U17280 (N_17280,N_14712,N_13889);
xnor U17281 (N_17281,N_11602,N_13825);
nor U17282 (N_17282,N_10863,N_11045);
and U17283 (N_17283,N_13468,N_10721);
nor U17284 (N_17284,N_13807,N_14078);
nand U17285 (N_17285,N_10569,N_14706);
xnor U17286 (N_17286,N_11357,N_12263);
nor U17287 (N_17287,N_11999,N_11777);
or U17288 (N_17288,N_13928,N_14778);
and U17289 (N_17289,N_13809,N_12526);
or U17290 (N_17290,N_10382,N_14220);
xor U17291 (N_17291,N_13246,N_11741);
nor U17292 (N_17292,N_12427,N_14361);
xnor U17293 (N_17293,N_13954,N_13774);
or U17294 (N_17294,N_14683,N_14846);
or U17295 (N_17295,N_11447,N_14136);
and U17296 (N_17296,N_11080,N_12558);
or U17297 (N_17297,N_11994,N_11739);
or U17298 (N_17298,N_13280,N_13910);
nand U17299 (N_17299,N_11727,N_14386);
or U17300 (N_17300,N_11628,N_12615);
nor U17301 (N_17301,N_13390,N_11674);
nor U17302 (N_17302,N_10840,N_13311);
nor U17303 (N_17303,N_12433,N_14723);
nor U17304 (N_17304,N_10511,N_14614);
or U17305 (N_17305,N_11288,N_13810);
xor U17306 (N_17306,N_12529,N_10337);
nand U17307 (N_17307,N_14715,N_14883);
xnor U17308 (N_17308,N_11535,N_13004);
and U17309 (N_17309,N_14701,N_12621);
and U17310 (N_17310,N_14930,N_12714);
and U17311 (N_17311,N_10538,N_12747);
and U17312 (N_17312,N_14839,N_13742);
nor U17313 (N_17313,N_11399,N_14328);
nand U17314 (N_17314,N_11582,N_13888);
nor U17315 (N_17315,N_11977,N_14389);
nand U17316 (N_17316,N_12018,N_11109);
xor U17317 (N_17317,N_13472,N_12540);
xor U17318 (N_17318,N_10297,N_12335);
or U17319 (N_17319,N_11757,N_12342);
or U17320 (N_17320,N_13876,N_10435);
or U17321 (N_17321,N_11641,N_11434);
xnor U17322 (N_17322,N_11959,N_11596);
or U17323 (N_17323,N_11531,N_14700);
and U17324 (N_17324,N_10737,N_12966);
xor U17325 (N_17325,N_10318,N_14213);
xor U17326 (N_17326,N_10919,N_12937);
and U17327 (N_17327,N_11579,N_11019);
nand U17328 (N_17328,N_14439,N_12360);
xnor U17329 (N_17329,N_14334,N_13952);
or U17330 (N_17330,N_13621,N_12838);
and U17331 (N_17331,N_12679,N_11852);
and U17332 (N_17332,N_14081,N_13539);
nand U17333 (N_17333,N_10477,N_13308);
nand U17334 (N_17334,N_10376,N_12758);
xnor U17335 (N_17335,N_11706,N_11008);
xnor U17336 (N_17336,N_13629,N_10162);
nand U17337 (N_17337,N_11442,N_14231);
and U17338 (N_17338,N_12549,N_11001);
and U17339 (N_17339,N_11725,N_10900);
nand U17340 (N_17340,N_10888,N_13484);
or U17341 (N_17341,N_13769,N_12500);
nand U17342 (N_17342,N_13669,N_14969);
xor U17343 (N_17343,N_11033,N_10332);
xor U17344 (N_17344,N_12654,N_11163);
nand U17345 (N_17345,N_12404,N_14950);
nor U17346 (N_17346,N_12306,N_10570);
nor U17347 (N_17347,N_14802,N_13664);
nor U17348 (N_17348,N_11853,N_13647);
nand U17349 (N_17349,N_11441,N_13149);
nand U17350 (N_17350,N_12443,N_13307);
nand U17351 (N_17351,N_11505,N_11306);
xor U17352 (N_17352,N_10464,N_11139);
nand U17353 (N_17353,N_12836,N_14466);
xor U17354 (N_17354,N_14597,N_13100);
xnor U17355 (N_17355,N_14394,N_11098);
nand U17356 (N_17356,N_10328,N_10194);
nand U17357 (N_17357,N_13863,N_14853);
nor U17358 (N_17358,N_14321,N_13414);
and U17359 (N_17359,N_12088,N_12680);
nor U17360 (N_17360,N_10655,N_12721);
nor U17361 (N_17361,N_13688,N_10189);
nor U17362 (N_17362,N_13565,N_12666);
and U17363 (N_17363,N_13781,N_10683);
and U17364 (N_17364,N_12888,N_13147);
nand U17365 (N_17365,N_13923,N_14530);
nor U17366 (N_17366,N_12173,N_11973);
nor U17367 (N_17367,N_12186,N_13057);
nor U17368 (N_17368,N_14681,N_14354);
nor U17369 (N_17369,N_10353,N_10666);
xor U17370 (N_17370,N_14919,N_11547);
nand U17371 (N_17371,N_14035,N_10949);
or U17372 (N_17372,N_10800,N_13096);
nand U17373 (N_17373,N_12544,N_10447);
nor U17374 (N_17374,N_13610,N_12988);
or U17375 (N_17375,N_14975,N_10134);
and U17376 (N_17376,N_11931,N_13240);
xor U17377 (N_17377,N_11421,N_13169);
xnor U17378 (N_17378,N_13187,N_14529);
nand U17379 (N_17379,N_13074,N_13492);
nand U17380 (N_17380,N_13507,N_13494);
xnor U17381 (N_17381,N_13007,N_13044);
nand U17382 (N_17382,N_11155,N_13955);
nor U17383 (N_17383,N_12022,N_13400);
xor U17384 (N_17384,N_13640,N_14981);
xnor U17385 (N_17385,N_14568,N_13698);
nand U17386 (N_17386,N_14347,N_13119);
and U17387 (N_17387,N_13787,N_10270);
nor U17388 (N_17388,N_11894,N_12259);
nor U17389 (N_17389,N_13320,N_10876);
or U17390 (N_17390,N_11989,N_10258);
and U17391 (N_17391,N_11245,N_12612);
and U17392 (N_17392,N_10864,N_14825);
and U17393 (N_17393,N_14959,N_12445);
and U17394 (N_17394,N_13081,N_13422);
and U17395 (N_17395,N_12833,N_10560);
or U17396 (N_17396,N_10150,N_12915);
nor U17397 (N_17397,N_11622,N_14144);
nand U17398 (N_17398,N_10527,N_12738);
and U17399 (N_17399,N_11873,N_12304);
and U17400 (N_17400,N_10986,N_12609);
or U17401 (N_17401,N_11593,N_13048);
xor U17402 (N_17402,N_14503,N_14671);
or U17403 (N_17403,N_10441,N_13126);
nor U17404 (N_17404,N_13211,N_13137);
or U17405 (N_17405,N_11198,N_12749);
and U17406 (N_17406,N_10324,N_10787);
xor U17407 (N_17407,N_10782,N_10768);
xnor U17408 (N_17408,N_11721,N_14592);
or U17409 (N_17409,N_12366,N_14200);
and U17410 (N_17410,N_12818,N_10491);
or U17411 (N_17411,N_13303,N_13156);
xor U17412 (N_17412,N_13183,N_13408);
and U17413 (N_17413,N_11103,N_11178);
nor U17414 (N_17414,N_11132,N_14456);
xnor U17415 (N_17415,N_12959,N_13030);
nor U17416 (N_17416,N_11828,N_14927);
xor U17417 (N_17417,N_14085,N_10837);
nor U17418 (N_17418,N_12244,N_14998);
nand U17419 (N_17419,N_14987,N_13727);
nor U17420 (N_17420,N_10108,N_11975);
nor U17421 (N_17421,N_11321,N_12295);
and U17422 (N_17422,N_14962,N_10614);
xnor U17423 (N_17423,N_14246,N_14005);
nand U17424 (N_17424,N_14120,N_11724);
or U17425 (N_17425,N_13880,N_12185);
nand U17426 (N_17426,N_10220,N_11699);
or U17427 (N_17427,N_10037,N_14427);
nor U17428 (N_17428,N_10539,N_14668);
and U17429 (N_17429,N_10204,N_11936);
or U17430 (N_17430,N_11798,N_11253);
or U17431 (N_17431,N_14907,N_12817);
and U17432 (N_17432,N_14188,N_14997);
and U17433 (N_17433,N_13567,N_14935);
nor U17434 (N_17434,N_14985,N_11169);
nand U17435 (N_17435,N_13362,N_13541);
xor U17436 (N_17436,N_11474,N_10914);
or U17437 (N_17437,N_13023,N_13751);
nor U17438 (N_17438,N_10735,N_14281);
xor U17439 (N_17439,N_10272,N_10159);
or U17440 (N_17440,N_11459,N_11285);
and U17441 (N_17441,N_13904,N_10687);
nand U17442 (N_17442,N_10245,N_10106);
and U17443 (N_17443,N_12055,N_11921);
nor U17444 (N_17444,N_14235,N_10278);
xnor U17445 (N_17445,N_10335,N_11299);
nand U17446 (N_17446,N_13485,N_12313);
or U17447 (N_17447,N_10142,N_14765);
nand U17448 (N_17448,N_13666,N_10909);
xor U17449 (N_17449,N_12391,N_10599);
and U17450 (N_17450,N_14905,N_12435);
xnor U17451 (N_17451,N_12851,N_12024);
nor U17452 (N_17452,N_13304,N_11052);
and U17453 (N_17453,N_11543,N_13331);
nand U17454 (N_17454,N_11722,N_13703);
or U17455 (N_17455,N_14488,N_12160);
xor U17456 (N_17456,N_11249,N_12319);
or U17457 (N_17457,N_14945,N_12192);
xor U17458 (N_17458,N_13976,N_11094);
or U17459 (N_17459,N_12858,N_14042);
nor U17460 (N_17460,N_14528,N_12760);
and U17461 (N_17461,N_13296,N_14149);
nand U17462 (N_17462,N_12655,N_12299);
nor U17463 (N_17463,N_14291,N_10365);
or U17464 (N_17464,N_14966,N_12632);
nor U17465 (N_17465,N_13430,N_12118);
nor U17466 (N_17466,N_13406,N_12305);
xnor U17467 (N_17467,N_10058,N_13761);
xor U17468 (N_17468,N_14266,N_10268);
and U17469 (N_17469,N_14961,N_10632);
or U17470 (N_17470,N_14026,N_14021);
or U17471 (N_17471,N_11933,N_13014);
or U17472 (N_17472,N_13887,N_14968);
or U17473 (N_17473,N_14843,N_14490);
nor U17474 (N_17474,N_12584,N_11608);
xor U17475 (N_17475,N_10346,N_13441);
xnor U17476 (N_17476,N_14033,N_12104);
nor U17477 (N_17477,N_10039,N_14234);
and U17478 (N_17478,N_11580,N_14947);
xnor U17479 (N_17479,N_10770,N_14146);
nand U17480 (N_17480,N_11726,N_12493);
and U17481 (N_17481,N_14031,N_10901);
or U17482 (N_17482,N_10458,N_12172);
or U17483 (N_17483,N_10877,N_10984);
and U17484 (N_17484,N_14705,N_12882);
nand U17485 (N_17485,N_13733,N_14123);
xnor U17486 (N_17486,N_14652,N_11347);
and U17487 (N_17487,N_12272,N_11495);
nand U17488 (N_17488,N_11466,N_12880);
or U17489 (N_17489,N_11234,N_12125);
nor U17490 (N_17490,N_11670,N_10115);
and U17491 (N_17491,N_12475,N_10257);
and U17492 (N_17492,N_11897,N_11836);
and U17493 (N_17493,N_11218,N_10649);
xnor U17494 (N_17494,N_10788,N_12643);
nand U17495 (N_17495,N_12043,N_12560);
nor U17496 (N_17496,N_12050,N_10298);
xnor U17497 (N_17497,N_10390,N_13332);
or U17498 (N_17498,N_10908,N_13780);
and U17499 (N_17499,N_10794,N_12764);
nor U17500 (N_17500,N_10507,N_12284);
and U17501 (N_17501,N_10334,N_14133);
xor U17502 (N_17502,N_12260,N_12695);
nor U17503 (N_17503,N_14447,N_12009);
xor U17504 (N_17504,N_14520,N_14757);
or U17505 (N_17505,N_10106,N_11271);
and U17506 (N_17506,N_11612,N_13848);
nor U17507 (N_17507,N_14886,N_14011);
nor U17508 (N_17508,N_11699,N_11706);
or U17509 (N_17509,N_10706,N_11613);
nand U17510 (N_17510,N_10241,N_13782);
nor U17511 (N_17511,N_14756,N_11323);
xor U17512 (N_17512,N_11676,N_12532);
and U17513 (N_17513,N_14630,N_11519);
nand U17514 (N_17514,N_14853,N_12455);
xor U17515 (N_17515,N_12417,N_14567);
or U17516 (N_17516,N_11966,N_11726);
and U17517 (N_17517,N_10218,N_13683);
xnor U17518 (N_17518,N_11933,N_10879);
nand U17519 (N_17519,N_14168,N_12825);
nand U17520 (N_17520,N_10439,N_11273);
nor U17521 (N_17521,N_10285,N_14725);
or U17522 (N_17522,N_10751,N_11419);
xor U17523 (N_17523,N_12136,N_14481);
and U17524 (N_17524,N_14313,N_10937);
nor U17525 (N_17525,N_14220,N_12565);
xnor U17526 (N_17526,N_14773,N_10740);
nor U17527 (N_17527,N_12667,N_12001);
or U17528 (N_17528,N_12117,N_10526);
nor U17529 (N_17529,N_11928,N_12820);
or U17530 (N_17530,N_12863,N_13211);
or U17531 (N_17531,N_14137,N_12968);
nand U17532 (N_17532,N_10577,N_10104);
and U17533 (N_17533,N_12381,N_11380);
nor U17534 (N_17534,N_13232,N_10784);
nand U17535 (N_17535,N_12869,N_13118);
and U17536 (N_17536,N_11673,N_10855);
nand U17537 (N_17537,N_14838,N_12889);
nand U17538 (N_17538,N_12637,N_14480);
xnor U17539 (N_17539,N_14059,N_11858);
and U17540 (N_17540,N_12315,N_10950);
or U17541 (N_17541,N_13273,N_12708);
and U17542 (N_17542,N_10280,N_10115);
nand U17543 (N_17543,N_14646,N_13241);
nor U17544 (N_17544,N_12514,N_14401);
nor U17545 (N_17545,N_12601,N_13255);
or U17546 (N_17546,N_12365,N_13865);
and U17547 (N_17547,N_11127,N_14022);
or U17548 (N_17548,N_14982,N_14973);
xnor U17549 (N_17549,N_14309,N_14446);
and U17550 (N_17550,N_13723,N_14582);
nor U17551 (N_17551,N_11320,N_13957);
or U17552 (N_17552,N_11846,N_10443);
or U17553 (N_17553,N_14634,N_12352);
and U17554 (N_17554,N_13338,N_13057);
and U17555 (N_17555,N_13029,N_12354);
and U17556 (N_17556,N_13143,N_10320);
or U17557 (N_17557,N_11381,N_13026);
xnor U17558 (N_17558,N_13775,N_13996);
and U17559 (N_17559,N_14379,N_10364);
nand U17560 (N_17560,N_12707,N_10183);
and U17561 (N_17561,N_12310,N_10403);
xnor U17562 (N_17562,N_13531,N_12461);
and U17563 (N_17563,N_11527,N_13026);
xnor U17564 (N_17564,N_14604,N_11473);
or U17565 (N_17565,N_14225,N_14368);
or U17566 (N_17566,N_10783,N_14928);
nor U17567 (N_17567,N_11336,N_14819);
and U17568 (N_17568,N_10055,N_12946);
and U17569 (N_17569,N_11972,N_14665);
xnor U17570 (N_17570,N_13368,N_12877);
nand U17571 (N_17571,N_11054,N_12107);
xnor U17572 (N_17572,N_10218,N_12174);
or U17573 (N_17573,N_11935,N_10984);
nand U17574 (N_17574,N_14436,N_13115);
or U17575 (N_17575,N_12411,N_12950);
nand U17576 (N_17576,N_14290,N_10489);
nand U17577 (N_17577,N_12005,N_12546);
nor U17578 (N_17578,N_11524,N_10330);
nand U17579 (N_17579,N_12751,N_11415);
and U17580 (N_17580,N_11538,N_10781);
nand U17581 (N_17581,N_12992,N_14874);
nor U17582 (N_17582,N_12133,N_14475);
or U17583 (N_17583,N_14819,N_12492);
nand U17584 (N_17584,N_14375,N_13507);
xor U17585 (N_17585,N_11235,N_11231);
nand U17586 (N_17586,N_14605,N_11805);
nor U17587 (N_17587,N_13335,N_11290);
xor U17588 (N_17588,N_12619,N_13255);
and U17589 (N_17589,N_12584,N_12305);
and U17590 (N_17590,N_10339,N_10089);
and U17591 (N_17591,N_10808,N_11826);
or U17592 (N_17592,N_14878,N_10538);
and U17593 (N_17593,N_12335,N_12395);
and U17594 (N_17594,N_14126,N_12497);
and U17595 (N_17595,N_13579,N_12715);
and U17596 (N_17596,N_10431,N_12856);
nand U17597 (N_17597,N_14578,N_12508);
and U17598 (N_17598,N_11955,N_11303);
nand U17599 (N_17599,N_14755,N_11707);
and U17600 (N_17600,N_13504,N_10602);
or U17601 (N_17601,N_12640,N_10997);
or U17602 (N_17602,N_12104,N_13312);
nor U17603 (N_17603,N_13759,N_14022);
xnor U17604 (N_17604,N_12910,N_10975);
nand U17605 (N_17605,N_13350,N_14850);
nor U17606 (N_17606,N_14733,N_11092);
or U17607 (N_17607,N_14950,N_11037);
or U17608 (N_17608,N_14089,N_13483);
nor U17609 (N_17609,N_11986,N_13679);
or U17610 (N_17610,N_10098,N_13639);
and U17611 (N_17611,N_14432,N_13561);
nand U17612 (N_17612,N_11663,N_10370);
and U17613 (N_17613,N_13808,N_11017);
nand U17614 (N_17614,N_13814,N_11031);
nand U17615 (N_17615,N_11539,N_12427);
or U17616 (N_17616,N_14763,N_14175);
nor U17617 (N_17617,N_10494,N_12352);
and U17618 (N_17618,N_13344,N_10526);
nor U17619 (N_17619,N_10718,N_14680);
nor U17620 (N_17620,N_11747,N_13720);
or U17621 (N_17621,N_11912,N_14051);
nor U17622 (N_17622,N_13143,N_11043);
and U17623 (N_17623,N_10655,N_10441);
and U17624 (N_17624,N_14602,N_13033);
and U17625 (N_17625,N_14810,N_13435);
nor U17626 (N_17626,N_10820,N_12734);
xnor U17627 (N_17627,N_11313,N_14983);
and U17628 (N_17628,N_10185,N_13998);
nand U17629 (N_17629,N_12371,N_14632);
or U17630 (N_17630,N_11194,N_14253);
xnor U17631 (N_17631,N_12225,N_12390);
xnor U17632 (N_17632,N_14134,N_10507);
nor U17633 (N_17633,N_10979,N_10716);
nor U17634 (N_17634,N_14203,N_13484);
xnor U17635 (N_17635,N_12903,N_11071);
and U17636 (N_17636,N_13849,N_12645);
nand U17637 (N_17637,N_11006,N_11081);
nand U17638 (N_17638,N_14559,N_10656);
xnor U17639 (N_17639,N_13352,N_12784);
nor U17640 (N_17640,N_13530,N_11969);
xor U17641 (N_17641,N_14695,N_14213);
xor U17642 (N_17642,N_10030,N_14049);
nand U17643 (N_17643,N_14225,N_13436);
nand U17644 (N_17644,N_12576,N_11350);
nor U17645 (N_17645,N_13927,N_11989);
and U17646 (N_17646,N_10216,N_13621);
nor U17647 (N_17647,N_11424,N_12299);
or U17648 (N_17648,N_11634,N_13363);
and U17649 (N_17649,N_10030,N_10372);
xor U17650 (N_17650,N_14711,N_13600);
xor U17651 (N_17651,N_13649,N_13777);
nor U17652 (N_17652,N_11445,N_14718);
nand U17653 (N_17653,N_13318,N_14480);
and U17654 (N_17654,N_12288,N_12380);
or U17655 (N_17655,N_13576,N_12791);
nand U17656 (N_17656,N_14268,N_12405);
nor U17657 (N_17657,N_14900,N_13297);
or U17658 (N_17658,N_10767,N_10293);
nor U17659 (N_17659,N_11449,N_13897);
xor U17660 (N_17660,N_12446,N_14827);
nand U17661 (N_17661,N_14467,N_13435);
or U17662 (N_17662,N_13587,N_12191);
xnor U17663 (N_17663,N_14174,N_12415);
or U17664 (N_17664,N_14365,N_11188);
nand U17665 (N_17665,N_12417,N_13751);
or U17666 (N_17666,N_10361,N_13019);
xnor U17667 (N_17667,N_12349,N_11631);
or U17668 (N_17668,N_13565,N_14418);
nor U17669 (N_17669,N_11785,N_14482);
and U17670 (N_17670,N_13195,N_12613);
nor U17671 (N_17671,N_13262,N_12190);
xor U17672 (N_17672,N_10850,N_11117);
and U17673 (N_17673,N_12783,N_10618);
nand U17674 (N_17674,N_10165,N_13146);
nor U17675 (N_17675,N_11365,N_10499);
xnor U17676 (N_17676,N_11962,N_13858);
nand U17677 (N_17677,N_13032,N_10365);
nand U17678 (N_17678,N_14152,N_11070);
nand U17679 (N_17679,N_12766,N_14594);
xnor U17680 (N_17680,N_14829,N_14601);
nand U17681 (N_17681,N_11398,N_14442);
xnor U17682 (N_17682,N_13894,N_10574);
xor U17683 (N_17683,N_13738,N_14198);
nand U17684 (N_17684,N_13725,N_10856);
xor U17685 (N_17685,N_12701,N_14257);
xor U17686 (N_17686,N_10908,N_10916);
nor U17687 (N_17687,N_10777,N_12733);
xnor U17688 (N_17688,N_13906,N_10592);
or U17689 (N_17689,N_14358,N_13542);
and U17690 (N_17690,N_12570,N_14488);
nand U17691 (N_17691,N_10325,N_14239);
nor U17692 (N_17692,N_10225,N_14571);
or U17693 (N_17693,N_14119,N_13259);
nor U17694 (N_17694,N_11697,N_10146);
or U17695 (N_17695,N_13665,N_14675);
xor U17696 (N_17696,N_14437,N_14363);
nor U17697 (N_17697,N_12306,N_10665);
nor U17698 (N_17698,N_14733,N_13456);
or U17699 (N_17699,N_10585,N_10067);
nand U17700 (N_17700,N_11472,N_13124);
xnor U17701 (N_17701,N_13870,N_14722);
nor U17702 (N_17702,N_10753,N_12610);
nand U17703 (N_17703,N_11194,N_10852);
xnor U17704 (N_17704,N_10133,N_10582);
nor U17705 (N_17705,N_12737,N_11277);
xnor U17706 (N_17706,N_11420,N_11812);
nor U17707 (N_17707,N_14316,N_11078);
nor U17708 (N_17708,N_10869,N_14476);
xnor U17709 (N_17709,N_13225,N_13822);
and U17710 (N_17710,N_11088,N_14692);
nand U17711 (N_17711,N_10978,N_14863);
nor U17712 (N_17712,N_11589,N_14917);
and U17713 (N_17713,N_10617,N_12986);
xor U17714 (N_17714,N_12345,N_10457);
nand U17715 (N_17715,N_14006,N_10525);
nor U17716 (N_17716,N_13621,N_13229);
and U17717 (N_17717,N_13971,N_14676);
nor U17718 (N_17718,N_11237,N_10840);
xor U17719 (N_17719,N_10548,N_14486);
xnor U17720 (N_17720,N_13775,N_11177);
or U17721 (N_17721,N_12173,N_10056);
nand U17722 (N_17722,N_13020,N_12004);
nor U17723 (N_17723,N_12401,N_12540);
xnor U17724 (N_17724,N_11360,N_11696);
or U17725 (N_17725,N_12590,N_13258);
xor U17726 (N_17726,N_11113,N_12475);
xnor U17727 (N_17727,N_13984,N_13348);
and U17728 (N_17728,N_14114,N_14603);
nor U17729 (N_17729,N_14873,N_12187);
nor U17730 (N_17730,N_14689,N_13112);
xor U17731 (N_17731,N_13333,N_10317);
xor U17732 (N_17732,N_14585,N_12550);
nand U17733 (N_17733,N_10326,N_13966);
or U17734 (N_17734,N_14089,N_10898);
nor U17735 (N_17735,N_12764,N_11188);
nand U17736 (N_17736,N_13234,N_11602);
nor U17737 (N_17737,N_14862,N_12208);
xor U17738 (N_17738,N_12038,N_10664);
or U17739 (N_17739,N_11694,N_11912);
xor U17740 (N_17740,N_11911,N_13036);
or U17741 (N_17741,N_12452,N_14604);
xnor U17742 (N_17742,N_10844,N_13106);
nor U17743 (N_17743,N_14652,N_13299);
xnor U17744 (N_17744,N_14002,N_11448);
nand U17745 (N_17745,N_13051,N_11730);
xnor U17746 (N_17746,N_10536,N_10736);
nor U17747 (N_17747,N_14603,N_12546);
nand U17748 (N_17748,N_12467,N_13934);
nor U17749 (N_17749,N_10761,N_12384);
xnor U17750 (N_17750,N_10939,N_11539);
or U17751 (N_17751,N_11993,N_10648);
nand U17752 (N_17752,N_13922,N_13829);
nor U17753 (N_17753,N_14900,N_13546);
and U17754 (N_17754,N_14888,N_14663);
or U17755 (N_17755,N_13526,N_11472);
and U17756 (N_17756,N_10727,N_11695);
nor U17757 (N_17757,N_13658,N_12297);
xnor U17758 (N_17758,N_12061,N_13395);
or U17759 (N_17759,N_11629,N_12538);
nand U17760 (N_17760,N_13160,N_14560);
or U17761 (N_17761,N_11923,N_12639);
nand U17762 (N_17762,N_13972,N_12240);
nand U17763 (N_17763,N_13379,N_11860);
nand U17764 (N_17764,N_12014,N_12702);
or U17765 (N_17765,N_10182,N_13151);
and U17766 (N_17766,N_10504,N_12268);
xor U17767 (N_17767,N_14954,N_12913);
nand U17768 (N_17768,N_13082,N_14163);
nor U17769 (N_17769,N_14939,N_13842);
xor U17770 (N_17770,N_13014,N_14718);
nor U17771 (N_17771,N_10198,N_11562);
or U17772 (N_17772,N_10040,N_14464);
and U17773 (N_17773,N_11972,N_11462);
or U17774 (N_17774,N_14234,N_11312);
xor U17775 (N_17775,N_14601,N_11399);
nand U17776 (N_17776,N_12432,N_11601);
nand U17777 (N_17777,N_12618,N_11465);
or U17778 (N_17778,N_12748,N_11369);
xnor U17779 (N_17779,N_11504,N_12450);
and U17780 (N_17780,N_10303,N_14982);
and U17781 (N_17781,N_12574,N_10457);
xnor U17782 (N_17782,N_14249,N_13533);
xnor U17783 (N_17783,N_14755,N_12941);
or U17784 (N_17784,N_12483,N_13762);
nor U17785 (N_17785,N_12943,N_14540);
nand U17786 (N_17786,N_12885,N_13864);
xor U17787 (N_17787,N_12840,N_14793);
or U17788 (N_17788,N_10436,N_11680);
nand U17789 (N_17789,N_14837,N_12105);
nor U17790 (N_17790,N_13124,N_14793);
or U17791 (N_17791,N_11962,N_14366);
and U17792 (N_17792,N_13938,N_14110);
or U17793 (N_17793,N_12887,N_14041);
and U17794 (N_17794,N_11960,N_12758);
xor U17795 (N_17795,N_12157,N_12782);
nor U17796 (N_17796,N_10262,N_12012);
nor U17797 (N_17797,N_13144,N_11769);
and U17798 (N_17798,N_13602,N_10085);
and U17799 (N_17799,N_11075,N_14728);
nand U17800 (N_17800,N_11671,N_13345);
xor U17801 (N_17801,N_10989,N_10647);
xnor U17802 (N_17802,N_10171,N_13456);
nor U17803 (N_17803,N_12584,N_11528);
nor U17804 (N_17804,N_13213,N_14843);
and U17805 (N_17805,N_11884,N_12315);
or U17806 (N_17806,N_13569,N_10294);
nor U17807 (N_17807,N_11297,N_13610);
or U17808 (N_17808,N_13491,N_10259);
and U17809 (N_17809,N_11990,N_10704);
xor U17810 (N_17810,N_13149,N_13568);
xnor U17811 (N_17811,N_10764,N_10471);
or U17812 (N_17812,N_10397,N_14050);
xor U17813 (N_17813,N_13502,N_12487);
or U17814 (N_17814,N_13313,N_13613);
and U17815 (N_17815,N_10971,N_13674);
or U17816 (N_17816,N_14252,N_13168);
and U17817 (N_17817,N_12938,N_10743);
or U17818 (N_17818,N_12544,N_10853);
nand U17819 (N_17819,N_11400,N_14884);
and U17820 (N_17820,N_12797,N_13521);
nand U17821 (N_17821,N_10680,N_13162);
xor U17822 (N_17822,N_13578,N_13047);
and U17823 (N_17823,N_14682,N_10894);
and U17824 (N_17824,N_11201,N_11870);
or U17825 (N_17825,N_10512,N_12895);
nand U17826 (N_17826,N_12384,N_12814);
xnor U17827 (N_17827,N_12040,N_10033);
and U17828 (N_17828,N_12627,N_12236);
xor U17829 (N_17829,N_13845,N_14788);
nand U17830 (N_17830,N_12389,N_12268);
and U17831 (N_17831,N_13329,N_13862);
or U17832 (N_17832,N_12742,N_14079);
xor U17833 (N_17833,N_13245,N_14832);
xnor U17834 (N_17834,N_12690,N_11992);
xnor U17835 (N_17835,N_13193,N_10220);
and U17836 (N_17836,N_13412,N_11164);
and U17837 (N_17837,N_10048,N_11758);
xor U17838 (N_17838,N_11408,N_13159);
nand U17839 (N_17839,N_11152,N_13063);
or U17840 (N_17840,N_14158,N_11028);
nand U17841 (N_17841,N_11582,N_11515);
or U17842 (N_17842,N_13149,N_14863);
or U17843 (N_17843,N_10677,N_13245);
or U17844 (N_17844,N_13932,N_11168);
and U17845 (N_17845,N_12254,N_12644);
nor U17846 (N_17846,N_13646,N_11611);
nor U17847 (N_17847,N_10964,N_12828);
nor U17848 (N_17848,N_12678,N_12047);
or U17849 (N_17849,N_11692,N_14509);
nor U17850 (N_17850,N_12457,N_10905);
or U17851 (N_17851,N_14932,N_14648);
nand U17852 (N_17852,N_14338,N_12657);
nor U17853 (N_17853,N_12438,N_12208);
or U17854 (N_17854,N_14099,N_13564);
or U17855 (N_17855,N_14167,N_13614);
nor U17856 (N_17856,N_13975,N_14579);
nand U17857 (N_17857,N_14740,N_14790);
nor U17858 (N_17858,N_10634,N_13686);
nor U17859 (N_17859,N_13816,N_10153);
xnor U17860 (N_17860,N_13758,N_12586);
or U17861 (N_17861,N_12098,N_10677);
nand U17862 (N_17862,N_11640,N_14428);
and U17863 (N_17863,N_14613,N_13435);
nor U17864 (N_17864,N_10023,N_13755);
nand U17865 (N_17865,N_12494,N_13301);
and U17866 (N_17866,N_12901,N_14681);
or U17867 (N_17867,N_14391,N_11897);
nand U17868 (N_17868,N_10716,N_10246);
and U17869 (N_17869,N_11082,N_10378);
nand U17870 (N_17870,N_10903,N_13939);
and U17871 (N_17871,N_13345,N_13507);
and U17872 (N_17872,N_12404,N_10169);
and U17873 (N_17873,N_12933,N_10740);
xor U17874 (N_17874,N_14018,N_14665);
nor U17875 (N_17875,N_14987,N_12990);
or U17876 (N_17876,N_12191,N_10171);
and U17877 (N_17877,N_10541,N_13672);
or U17878 (N_17878,N_12437,N_13868);
nor U17879 (N_17879,N_11282,N_10541);
nor U17880 (N_17880,N_11578,N_10785);
nor U17881 (N_17881,N_14830,N_14760);
and U17882 (N_17882,N_10391,N_13867);
and U17883 (N_17883,N_13086,N_13316);
nor U17884 (N_17884,N_11060,N_13097);
nor U17885 (N_17885,N_12281,N_13216);
or U17886 (N_17886,N_11371,N_12784);
or U17887 (N_17887,N_14528,N_12376);
xor U17888 (N_17888,N_10109,N_10865);
and U17889 (N_17889,N_10262,N_12285);
nand U17890 (N_17890,N_12374,N_11779);
and U17891 (N_17891,N_12759,N_10767);
or U17892 (N_17892,N_10414,N_14469);
nor U17893 (N_17893,N_13261,N_12886);
nor U17894 (N_17894,N_13650,N_14094);
nand U17895 (N_17895,N_12416,N_10273);
or U17896 (N_17896,N_10801,N_10459);
xor U17897 (N_17897,N_10278,N_11244);
xor U17898 (N_17898,N_14913,N_14269);
or U17899 (N_17899,N_13518,N_14688);
and U17900 (N_17900,N_12346,N_13601);
and U17901 (N_17901,N_13463,N_11828);
nor U17902 (N_17902,N_11018,N_12699);
and U17903 (N_17903,N_12285,N_10596);
and U17904 (N_17904,N_13187,N_14707);
xor U17905 (N_17905,N_12366,N_14341);
and U17906 (N_17906,N_10804,N_12554);
nand U17907 (N_17907,N_11958,N_12782);
nand U17908 (N_17908,N_14904,N_14927);
or U17909 (N_17909,N_13649,N_12526);
xnor U17910 (N_17910,N_10742,N_14082);
nand U17911 (N_17911,N_12477,N_11009);
nor U17912 (N_17912,N_10126,N_13071);
nand U17913 (N_17913,N_12573,N_10696);
nand U17914 (N_17914,N_10666,N_12510);
or U17915 (N_17915,N_10962,N_10040);
nand U17916 (N_17916,N_14812,N_14082);
nand U17917 (N_17917,N_11565,N_10791);
nand U17918 (N_17918,N_14829,N_12915);
or U17919 (N_17919,N_10326,N_14115);
or U17920 (N_17920,N_11625,N_13275);
nor U17921 (N_17921,N_11007,N_14242);
or U17922 (N_17922,N_11319,N_10395);
or U17923 (N_17923,N_14873,N_12924);
and U17924 (N_17924,N_11519,N_11582);
xnor U17925 (N_17925,N_11100,N_10212);
xnor U17926 (N_17926,N_10982,N_13611);
nand U17927 (N_17927,N_13338,N_13170);
and U17928 (N_17928,N_14072,N_10663);
xor U17929 (N_17929,N_11453,N_10911);
xor U17930 (N_17930,N_13841,N_10824);
and U17931 (N_17931,N_10639,N_14982);
nand U17932 (N_17932,N_12259,N_14111);
nand U17933 (N_17933,N_11552,N_10494);
and U17934 (N_17934,N_10029,N_13043);
nand U17935 (N_17935,N_13749,N_13130);
nand U17936 (N_17936,N_13288,N_12324);
nand U17937 (N_17937,N_13437,N_12556);
nand U17938 (N_17938,N_14509,N_11562);
or U17939 (N_17939,N_11905,N_14690);
and U17940 (N_17940,N_11790,N_11593);
xor U17941 (N_17941,N_12508,N_13731);
or U17942 (N_17942,N_12834,N_12004);
or U17943 (N_17943,N_14238,N_11894);
nor U17944 (N_17944,N_12370,N_11118);
and U17945 (N_17945,N_10944,N_14376);
nand U17946 (N_17946,N_14531,N_13321);
nand U17947 (N_17947,N_13156,N_11625);
nor U17948 (N_17948,N_14278,N_13531);
nand U17949 (N_17949,N_11517,N_11322);
xor U17950 (N_17950,N_14400,N_14804);
and U17951 (N_17951,N_14900,N_12581);
nand U17952 (N_17952,N_11261,N_11908);
nor U17953 (N_17953,N_14471,N_14209);
nor U17954 (N_17954,N_13262,N_10304);
or U17955 (N_17955,N_13786,N_13689);
nor U17956 (N_17956,N_12371,N_12777);
nand U17957 (N_17957,N_13031,N_13959);
xnor U17958 (N_17958,N_10641,N_10531);
xor U17959 (N_17959,N_10275,N_14102);
and U17960 (N_17960,N_10887,N_11856);
and U17961 (N_17961,N_10448,N_11840);
and U17962 (N_17962,N_13018,N_11523);
xor U17963 (N_17963,N_10744,N_10396);
nor U17964 (N_17964,N_10237,N_11227);
nor U17965 (N_17965,N_11365,N_14138);
and U17966 (N_17966,N_12770,N_13438);
xor U17967 (N_17967,N_13878,N_12758);
nor U17968 (N_17968,N_12597,N_10506);
xor U17969 (N_17969,N_11851,N_13012);
and U17970 (N_17970,N_14556,N_13524);
xnor U17971 (N_17971,N_10195,N_12546);
nor U17972 (N_17972,N_10379,N_12865);
nor U17973 (N_17973,N_10560,N_13532);
nand U17974 (N_17974,N_13268,N_11284);
xor U17975 (N_17975,N_12159,N_12816);
nor U17976 (N_17976,N_13813,N_13925);
and U17977 (N_17977,N_13857,N_13762);
nor U17978 (N_17978,N_13732,N_10623);
nand U17979 (N_17979,N_12086,N_11419);
xnor U17980 (N_17980,N_11258,N_13362);
xor U17981 (N_17981,N_13052,N_10434);
nor U17982 (N_17982,N_13939,N_10325);
nand U17983 (N_17983,N_14609,N_12990);
or U17984 (N_17984,N_11459,N_12158);
nor U17985 (N_17985,N_11740,N_13858);
and U17986 (N_17986,N_13237,N_12390);
and U17987 (N_17987,N_13577,N_10035);
nand U17988 (N_17988,N_11494,N_12569);
nand U17989 (N_17989,N_11973,N_11681);
or U17990 (N_17990,N_12079,N_12992);
and U17991 (N_17991,N_10792,N_13720);
nand U17992 (N_17992,N_13548,N_10002);
or U17993 (N_17993,N_11514,N_14724);
xor U17994 (N_17994,N_12520,N_12464);
nand U17995 (N_17995,N_12767,N_13563);
nand U17996 (N_17996,N_10075,N_12281);
xor U17997 (N_17997,N_11389,N_12550);
nand U17998 (N_17998,N_11199,N_10233);
or U17999 (N_17999,N_14824,N_13894);
nor U18000 (N_18000,N_14928,N_10489);
or U18001 (N_18001,N_14305,N_12387);
xnor U18002 (N_18002,N_11070,N_12709);
xnor U18003 (N_18003,N_13514,N_12549);
xnor U18004 (N_18004,N_10608,N_10468);
xnor U18005 (N_18005,N_11049,N_13034);
nor U18006 (N_18006,N_14430,N_10642);
nor U18007 (N_18007,N_10678,N_11801);
or U18008 (N_18008,N_10827,N_13209);
and U18009 (N_18009,N_13869,N_13887);
or U18010 (N_18010,N_13328,N_10005);
or U18011 (N_18011,N_12207,N_13344);
nor U18012 (N_18012,N_11343,N_11714);
nor U18013 (N_18013,N_14909,N_11390);
nor U18014 (N_18014,N_12653,N_11924);
nor U18015 (N_18015,N_13780,N_13676);
and U18016 (N_18016,N_11761,N_12777);
nand U18017 (N_18017,N_10707,N_11588);
and U18018 (N_18018,N_11377,N_13248);
and U18019 (N_18019,N_12370,N_13151);
and U18020 (N_18020,N_11541,N_13813);
and U18021 (N_18021,N_14050,N_12863);
and U18022 (N_18022,N_12612,N_10661);
or U18023 (N_18023,N_11143,N_11726);
and U18024 (N_18024,N_10886,N_12137);
nor U18025 (N_18025,N_13272,N_14694);
nor U18026 (N_18026,N_12526,N_14180);
nor U18027 (N_18027,N_12339,N_14273);
or U18028 (N_18028,N_13355,N_10167);
or U18029 (N_18029,N_13707,N_14166);
nor U18030 (N_18030,N_10845,N_14554);
nand U18031 (N_18031,N_10335,N_14172);
nand U18032 (N_18032,N_14055,N_11417);
xnor U18033 (N_18033,N_12390,N_13343);
or U18034 (N_18034,N_12214,N_13070);
nand U18035 (N_18035,N_14436,N_13397);
xnor U18036 (N_18036,N_13752,N_10444);
nor U18037 (N_18037,N_11943,N_12104);
nor U18038 (N_18038,N_10096,N_14921);
nand U18039 (N_18039,N_13816,N_11208);
xor U18040 (N_18040,N_14273,N_14216);
nand U18041 (N_18041,N_14816,N_13424);
or U18042 (N_18042,N_13824,N_14267);
or U18043 (N_18043,N_10495,N_10350);
nand U18044 (N_18044,N_14327,N_14649);
xor U18045 (N_18045,N_11454,N_12684);
or U18046 (N_18046,N_14050,N_11215);
nand U18047 (N_18047,N_14736,N_13447);
and U18048 (N_18048,N_13238,N_11698);
or U18049 (N_18049,N_11871,N_12768);
and U18050 (N_18050,N_10613,N_14007);
or U18051 (N_18051,N_10308,N_13997);
xnor U18052 (N_18052,N_12569,N_13134);
nand U18053 (N_18053,N_12989,N_10172);
and U18054 (N_18054,N_13924,N_10283);
or U18055 (N_18055,N_11244,N_12285);
nand U18056 (N_18056,N_11298,N_14796);
xor U18057 (N_18057,N_11461,N_10030);
nor U18058 (N_18058,N_10073,N_12227);
nor U18059 (N_18059,N_12778,N_10337);
xor U18060 (N_18060,N_13520,N_10897);
nor U18061 (N_18061,N_11232,N_11669);
xnor U18062 (N_18062,N_12450,N_12616);
and U18063 (N_18063,N_11026,N_14654);
nor U18064 (N_18064,N_10802,N_12195);
nor U18065 (N_18065,N_14905,N_12167);
and U18066 (N_18066,N_12706,N_13131);
or U18067 (N_18067,N_11739,N_11557);
nor U18068 (N_18068,N_14522,N_10234);
or U18069 (N_18069,N_10640,N_10968);
xor U18070 (N_18070,N_13078,N_10740);
nand U18071 (N_18071,N_12673,N_14383);
nor U18072 (N_18072,N_11496,N_11343);
nor U18073 (N_18073,N_12322,N_12765);
and U18074 (N_18074,N_13381,N_13254);
xor U18075 (N_18075,N_12635,N_14798);
and U18076 (N_18076,N_13945,N_10501);
nand U18077 (N_18077,N_14731,N_10048);
xor U18078 (N_18078,N_13711,N_10466);
xor U18079 (N_18079,N_12469,N_13272);
and U18080 (N_18080,N_14833,N_12815);
or U18081 (N_18081,N_12617,N_11068);
xnor U18082 (N_18082,N_10334,N_13303);
and U18083 (N_18083,N_10577,N_12243);
nor U18084 (N_18084,N_14397,N_10869);
xnor U18085 (N_18085,N_13862,N_14992);
xor U18086 (N_18086,N_11108,N_14228);
and U18087 (N_18087,N_12611,N_11281);
nand U18088 (N_18088,N_14655,N_13208);
or U18089 (N_18089,N_14973,N_11422);
or U18090 (N_18090,N_13146,N_11541);
xor U18091 (N_18091,N_12535,N_12879);
nor U18092 (N_18092,N_12910,N_12917);
nor U18093 (N_18093,N_11522,N_13037);
nand U18094 (N_18094,N_10093,N_10425);
and U18095 (N_18095,N_12772,N_12357);
nor U18096 (N_18096,N_10185,N_14374);
nor U18097 (N_18097,N_11549,N_14932);
nor U18098 (N_18098,N_10491,N_11159);
or U18099 (N_18099,N_10026,N_11437);
and U18100 (N_18100,N_10251,N_10588);
and U18101 (N_18101,N_13708,N_10746);
xnor U18102 (N_18102,N_14120,N_12700);
xnor U18103 (N_18103,N_10775,N_11830);
and U18104 (N_18104,N_13511,N_13558);
xnor U18105 (N_18105,N_14727,N_14010);
nor U18106 (N_18106,N_11067,N_11919);
nand U18107 (N_18107,N_10245,N_13061);
nor U18108 (N_18108,N_11330,N_11044);
xor U18109 (N_18109,N_12996,N_11607);
nor U18110 (N_18110,N_14585,N_14614);
nand U18111 (N_18111,N_10142,N_12241);
or U18112 (N_18112,N_12929,N_13449);
xnor U18113 (N_18113,N_14751,N_13329);
xor U18114 (N_18114,N_14562,N_12863);
nand U18115 (N_18115,N_10254,N_12233);
and U18116 (N_18116,N_10426,N_14615);
xnor U18117 (N_18117,N_14243,N_11905);
nand U18118 (N_18118,N_11733,N_12395);
and U18119 (N_18119,N_11244,N_10034);
nor U18120 (N_18120,N_11459,N_10122);
nand U18121 (N_18121,N_12241,N_10606);
or U18122 (N_18122,N_13479,N_11990);
and U18123 (N_18123,N_13106,N_12228);
or U18124 (N_18124,N_14184,N_12816);
or U18125 (N_18125,N_10016,N_12276);
and U18126 (N_18126,N_14796,N_14386);
and U18127 (N_18127,N_11213,N_11440);
nand U18128 (N_18128,N_10134,N_13558);
and U18129 (N_18129,N_12973,N_10677);
and U18130 (N_18130,N_11490,N_10419);
and U18131 (N_18131,N_13023,N_14975);
nor U18132 (N_18132,N_12569,N_13071);
or U18133 (N_18133,N_14805,N_11721);
xor U18134 (N_18134,N_10089,N_11831);
nand U18135 (N_18135,N_10120,N_13150);
nand U18136 (N_18136,N_11296,N_12067);
and U18137 (N_18137,N_10125,N_13737);
and U18138 (N_18138,N_10774,N_10056);
or U18139 (N_18139,N_14039,N_13685);
or U18140 (N_18140,N_13807,N_13465);
or U18141 (N_18141,N_11148,N_12414);
xnor U18142 (N_18142,N_13616,N_14383);
and U18143 (N_18143,N_10029,N_13956);
and U18144 (N_18144,N_14133,N_13425);
xor U18145 (N_18145,N_10515,N_12023);
xor U18146 (N_18146,N_13938,N_10374);
and U18147 (N_18147,N_13323,N_11848);
or U18148 (N_18148,N_10465,N_12973);
and U18149 (N_18149,N_11314,N_11223);
or U18150 (N_18150,N_11881,N_11116);
and U18151 (N_18151,N_11864,N_12953);
nand U18152 (N_18152,N_14720,N_13112);
xor U18153 (N_18153,N_14143,N_12112);
nor U18154 (N_18154,N_10355,N_13070);
xnor U18155 (N_18155,N_14513,N_12623);
and U18156 (N_18156,N_13941,N_13656);
nand U18157 (N_18157,N_10235,N_11502);
nor U18158 (N_18158,N_10586,N_14208);
or U18159 (N_18159,N_11126,N_11756);
nor U18160 (N_18160,N_14443,N_10129);
and U18161 (N_18161,N_12562,N_13308);
and U18162 (N_18162,N_12285,N_11417);
nor U18163 (N_18163,N_11184,N_10693);
or U18164 (N_18164,N_10997,N_10931);
or U18165 (N_18165,N_10439,N_11989);
xnor U18166 (N_18166,N_10876,N_12958);
nor U18167 (N_18167,N_14176,N_12245);
or U18168 (N_18168,N_13110,N_11339);
or U18169 (N_18169,N_12771,N_10861);
and U18170 (N_18170,N_11740,N_10737);
nand U18171 (N_18171,N_10256,N_14106);
nand U18172 (N_18172,N_10964,N_12342);
nand U18173 (N_18173,N_14573,N_13757);
nor U18174 (N_18174,N_10913,N_14166);
or U18175 (N_18175,N_14583,N_11960);
or U18176 (N_18176,N_14238,N_11088);
nand U18177 (N_18177,N_12559,N_14527);
or U18178 (N_18178,N_12591,N_11321);
or U18179 (N_18179,N_10329,N_13891);
and U18180 (N_18180,N_10429,N_12361);
nor U18181 (N_18181,N_11266,N_12246);
nand U18182 (N_18182,N_11498,N_12939);
and U18183 (N_18183,N_12100,N_14986);
xnor U18184 (N_18184,N_10827,N_12143);
xor U18185 (N_18185,N_10560,N_14991);
or U18186 (N_18186,N_10663,N_14528);
nand U18187 (N_18187,N_14325,N_12332);
xor U18188 (N_18188,N_10617,N_13705);
nand U18189 (N_18189,N_14270,N_13602);
and U18190 (N_18190,N_11894,N_11038);
and U18191 (N_18191,N_10775,N_13682);
nand U18192 (N_18192,N_10627,N_13539);
nor U18193 (N_18193,N_11707,N_13743);
and U18194 (N_18194,N_11639,N_13434);
nand U18195 (N_18195,N_10632,N_13973);
and U18196 (N_18196,N_14966,N_11385);
and U18197 (N_18197,N_10692,N_10604);
xnor U18198 (N_18198,N_13219,N_11137);
xor U18199 (N_18199,N_13071,N_10276);
xor U18200 (N_18200,N_13858,N_12835);
or U18201 (N_18201,N_10906,N_13813);
or U18202 (N_18202,N_12721,N_13000);
or U18203 (N_18203,N_11536,N_12262);
and U18204 (N_18204,N_13641,N_12835);
nand U18205 (N_18205,N_11362,N_11283);
nor U18206 (N_18206,N_14052,N_11638);
or U18207 (N_18207,N_10490,N_13365);
or U18208 (N_18208,N_12769,N_10828);
nor U18209 (N_18209,N_13648,N_11743);
or U18210 (N_18210,N_11985,N_12990);
and U18211 (N_18211,N_14003,N_12202);
xor U18212 (N_18212,N_12979,N_10779);
or U18213 (N_18213,N_11346,N_11449);
and U18214 (N_18214,N_14484,N_13264);
and U18215 (N_18215,N_11708,N_14657);
and U18216 (N_18216,N_12563,N_11333);
nand U18217 (N_18217,N_12363,N_14820);
and U18218 (N_18218,N_13094,N_13655);
nor U18219 (N_18219,N_10510,N_14820);
nor U18220 (N_18220,N_14792,N_12492);
or U18221 (N_18221,N_14266,N_14289);
or U18222 (N_18222,N_12170,N_13094);
xor U18223 (N_18223,N_12073,N_12989);
or U18224 (N_18224,N_12083,N_11704);
or U18225 (N_18225,N_10454,N_14361);
and U18226 (N_18226,N_12919,N_11617);
nand U18227 (N_18227,N_14510,N_10682);
or U18228 (N_18228,N_11857,N_13682);
or U18229 (N_18229,N_11343,N_13351);
and U18230 (N_18230,N_11752,N_13310);
and U18231 (N_18231,N_14261,N_12031);
nor U18232 (N_18232,N_11050,N_11955);
nand U18233 (N_18233,N_14005,N_13378);
nand U18234 (N_18234,N_12065,N_14611);
nor U18235 (N_18235,N_12247,N_11756);
and U18236 (N_18236,N_14616,N_10983);
nor U18237 (N_18237,N_10564,N_13077);
and U18238 (N_18238,N_13161,N_14747);
xnor U18239 (N_18239,N_10616,N_10283);
xnor U18240 (N_18240,N_14291,N_14364);
nor U18241 (N_18241,N_11602,N_11860);
nor U18242 (N_18242,N_13111,N_14952);
xnor U18243 (N_18243,N_10673,N_11444);
and U18244 (N_18244,N_12633,N_10876);
nand U18245 (N_18245,N_14552,N_14562);
xor U18246 (N_18246,N_13891,N_10637);
xor U18247 (N_18247,N_14355,N_11985);
nand U18248 (N_18248,N_11732,N_10697);
xnor U18249 (N_18249,N_13266,N_14375);
xnor U18250 (N_18250,N_13036,N_10136);
or U18251 (N_18251,N_13321,N_11778);
xnor U18252 (N_18252,N_13774,N_12811);
nor U18253 (N_18253,N_13208,N_11150);
or U18254 (N_18254,N_11679,N_14286);
nor U18255 (N_18255,N_10463,N_10179);
nor U18256 (N_18256,N_12686,N_13927);
or U18257 (N_18257,N_13322,N_12060);
or U18258 (N_18258,N_10969,N_11040);
nor U18259 (N_18259,N_11409,N_14789);
nor U18260 (N_18260,N_12873,N_10756);
nor U18261 (N_18261,N_14783,N_10002);
or U18262 (N_18262,N_10441,N_12180);
nand U18263 (N_18263,N_11962,N_10913);
nand U18264 (N_18264,N_11653,N_11128);
or U18265 (N_18265,N_12798,N_14385);
xor U18266 (N_18266,N_10406,N_10561);
nor U18267 (N_18267,N_14977,N_10304);
xnor U18268 (N_18268,N_13334,N_10903);
nor U18269 (N_18269,N_14290,N_13211);
nor U18270 (N_18270,N_13644,N_11837);
xnor U18271 (N_18271,N_13084,N_13991);
or U18272 (N_18272,N_10744,N_13231);
nand U18273 (N_18273,N_14954,N_12882);
nor U18274 (N_18274,N_12940,N_14416);
and U18275 (N_18275,N_11465,N_14209);
and U18276 (N_18276,N_14806,N_10833);
xor U18277 (N_18277,N_12013,N_11020);
xnor U18278 (N_18278,N_14210,N_12290);
nand U18279 (N_18279,N_11607,N_11888);
and U18280 (N_18280,N_10651,N_13146);
or U18281 (N_18281,N_13602,N_12648);
nor U18282 (N_18282,N_14719,N_13906);
and U18283 (N_18283,N_11943,N_10151);
and U18284 (N_18284,N_14303,N_14136);
and U18285 (N_18285,N_13578,N_13234);
or U18286 (N_18286,N_11973,N_13159);
nand U18287 (N_18287,N_11350,N_11659);
nand U18288 (N_18288,N_14922,N_12644);
nor U18289 (N_18289,N_14606,N_10900);
nand U18290 (N_18290,N_12442,N_12194);
nor U18291 (N_18291,N_13550,N_10328);
nor U18292 (N_18292,N_13672,N_11502);
xnor U18293 (N_18293,N_12173,N_13694);
and U18294 (N_18294,N_12117,N_13822);
and U18295 (N_18295,N_11199,N_12775);
xnor U18296 (N_18296,N_13174,N_10599);
or U18297 (N_18297,N_13565,N_13435);
nand U18298 (N_18298,N_11718,N_10132);
nand U18299 (N_18299,N_10019,N_12545);
xor U18300 (N_18300,N_14883,N_12001);
and U18301 (N_18301,N_13440,N_10094);
nand U18302 (N_18302,N_11646,N_10735);
nor U18303 (N_18303,N_13350,N_13144);
or U18304 (N_18304,N_13348,N_11334);
and U18305 (N_18305,N_12348,N_10659);
and U18306 (N_18306,N_12997,N_10918);
nand U18307 (N_18307,N_13610,N_13506);
xor U18308 (N_18308,N_14514,N_13501);
nand U18309 (N_18309,N_11049,N_11614);
or U18310 (N_18310,N_14147,N_13759);
nand U18311 (N_18311,N_12507,N_12487);
or U18312 (N_18312,N_11349,N_14004);
or U18313 (N_18313,N_11415,N_14713);
and U18314 (N_18314,N_10406,N_12330);
xnor U18315 (N_18315,N_11405,N_13131);
or U18316 (N_18316,N_12369,N_10686);
nand U18317 (N_18317,N_10210,N_12983);
nand U18318 (N_18318,N_11708,N_14844);
and U18319 (N_18319,N_14484,N_13426);
and U18320 (N_18320,N_12729,N_11665);
nor U18321 (N_18321,N_11206,N_12690);
xor U18322 (N_18322,N_11707,N_11788);
nand U18323 (N_18323,N_14291,N_10876);
or U18324 (N_18324,N_13355,N_11666);
nor U18325 (N_18325,N_11958,N_14382);
or U18326 (N_18326,N_10028,N_14345);
and U18327 (N_18327,N_13408,N_12785);
nor U18328 (N_18328,N_14390,N_13191);
nor U18329 (N_18329,N_11241,N_13137);
nand U18330 (N_18330,N_10375,N_10951);
or U18331 (N_18331,N_12215,N_14380);
xnor U18332 (N_18332,N_12466,N_13085);
xnor U18333 (N_18333,N_14238,N_14565);
or U18334 (N_18334,N_10920,N_14024);
nor U18335 (N_18335,N_14636,N_11710);
or U18336 (N_18336,N_13963,N_11616);
nor U18337 (N_18337,N_14964,N_11054);
and U18338 (N_18338,N_10422,N_10436);
and U18339 (N_18339,N_14199,N_13486);
and U18340 (N_18340,N_12328,N_12875);
nand U18341 (N_18341,N_12005,N_12495);
and U18342 (N_18342,N_11272,N_13533);
nand U18343 (N_18343,N_12261,N_13885);
nor U18344 (N_18344,N_14546,N_12961);
or U18345 (N_18345,N_14659,N_11120);
or U18346 (N_18346,N_10246,N_13613);
xnor U18347 (N_18347,N_13920,N_10221);
nand U18348 (N_18348,N_11429,N_11244);
nor U18349 (N_18349,N_13556,N_14681);
or U18350 (N_18350,N_12075,N_12999);
xnor U18351 (N_18351,N_14328,N_13461);
xnor U18352 (N_18352,N_14364,N_11218);
xnor U18353 (N_18353,N_13449,N_10194);
nor U18354 (N_18354,N_14249,N_11759);
nand U18355 (N_18355,N_13585,N_11645);
or U18356 (N_18356,N_12924,N_12703);
nor U18357 (N_18357,N_13511,N_11684);
nand U18358 (N_18358,N_10650,N_12013);
nand U18359 (N_18359,N_10273,N_12634);
xnor U18360 (N_18360,N_11770,N_10651);
or U18361 (N_18361,N_12188,N_11994);
and U18362 (N_18362,N_12402,N_12061);
and U18363 (N_18363,N_10806,N_11144);
nand U18364 (N_18364,N_10440,N_13201);
nor U18365 (N_18365,N_12600,N_14429);
nand U18366 (N_18366,N_10292,N_13345);
or U18367 (N_18367,N_12273,N_12194);
nor U18368 (N_18368,N_10818,N_13172);
nand U18369 (N_18369,N_12802,N_12923);
xor U18370 (N_18370,N_11938,N_12443);
nand U18371 (N_18371,N_12392,N_10185);
or U18372 (N_18372,N_10018,N_14972);
xnor U18373 (N_18373,N_11253,N_11375);
nor U18374 (N_18374,N_12778,N_14848);
nor U18375 (N_18375,N_13839,N_12758);
or U18376 (N_18376,N_14264,N_14294);
or U18377 (N_18377,N_14606,N_13562);
xnor U18378 (N_18378,N_11210,N_13735);
and U18379 (N_18379,N_14652,N_10227);
xnor U18380 (N_18380,N_12873,N_14481);
nand U18381 (N_18381,N_10092,N_13571);
nor U18382 (N_18382,N_12847,N_14744);
nor U18383 (N_18383,N_11317,N_14323);
or U18384 (N_18384,N_14148,N_11590);
or U18385 (N_18385,N_13019,N_10659);
xnor U18386 (N_18386,N_14443,N_10501);
nor U18387 (N_18387,N_14124,N_12496);
nand U18388 (N_18388,N_11336,N_13135);
or U18389 (N_18389,N_12830,N_11272);
xor U18390 (N_18390,N_14692,N_11534);
xor U18391 (N_18391,N_14833,N_13218);
xnor U18392 (N_18392,N_12987,N_11653);
or U18393 (N_18393,N_10367,N_10045);
and U18394 (N_18394,N_13420,N_13713);
xor U18395 (N_18395,N_13416,N_10120);
xnor U18396 (N_18396,N_13276,N_11514);
nand U18397 (N_18397,N_11970,N_12967);
nor U18398 (N_18398,N_11060,N_13630);
xor U18399 (N_18399,N_12686,N_13037);
xnor U18400 (N_18400,N_13743,N_12796);
xnor U18401 (N_18401,N_14683,N_12010);
nand U18402 (N_18402,N_10064,N_14992);
and U18403 (N_18403,N_10063,N_14789);
nand U18404 (N_18404,N_10147,N_10282);
nor U18405 (N_18405,N_11667,N_10836);
or U18406 (N_18406,N_11991,N_11401);
nor U18407 (N_18407,N_10073,N_13197);
and U18408 (N_18408,N_11619,N_11483);
or U18409 (N_18409,N_14316,N_11904);
xnor U18410 (N_18410,N_11038,N_12847);
nand U18411 (N_18411,N_14299,N_14162);
nand U18412 (N_18412,N_10931,N_14090);
or U18413 (N_18413,N_12565,N_10613);
nand U18414 (N_18414,N_10217,N_11596);
xnor U18415 (N_18415,N_11450,N_13046);
or U18416 (N_18416,N_14885,N_13964);
nand U18417 (N_18417,N_12557,N_10966);
nand U18418 (N_18418,N_13525,N_13302);
xor U18419 (N_18419,N_12113,N_11860);
nand U18420 (N_18420,N_13355,N_14950);
xor U18421 (N_18421,N_14734,N_11895);
xor U18422 (N_18422,N_12321,N_13726);
and U18423 (N_18423,N_11020,N_14614);
nand U18424 (N_18424,N_11588,N_10613);
or U18425 (N_18425,N_13374,N_13809);
or U18426 (N_18426,N_12226,N_13432);
or U18427 (N_18427,N_11877,N_10968);
xor U18428 (N_18428,N_11111,N_12989);
nor U18429 (N_18429,N_12242,N_11615);
nand U18430 (N_18430,N_13953,N_13739);
nand U18431 (N_18431,N_13883,N_13658);
xor U18432 (N_18432,N_11512,N_13072);
xnor U18433 (N_18433,N_11685,N_10604);
or U18434 (N_18434,N_12240,N_11700);
and U18435 (N_18435,N_14536,N_13559);
nor U18436 (N_18436,N_10546,N_11069);
nor U18437 (N_18437,N_11916,N_11900);
nand U18438 (N_18438,N_11092,N_12550);
nand U18439 (N_18439,N_13515,N_14634);
xor U18440 (N_18440,N_14919,N_11508);
nand U18441 (N_18441,N_14436,N_10749);
nor U18442 (N_18442,N_14642,N_14380);
nand U18443 (N_18443,N_10966,N_10978);
nand U18444 (N_18444,N_10644,N_13943);
xor U18445 (N_18445,N_13858,N_13608);
or U18446 (N_18446,N_11791,N_10237);
nor U18447 (N_18447,N_13550,N_12202);
or U18448 (N_18448,N_12258,N_10444);
or U18449 (N_18449,N_11187,N_14089);
and U18450 (N_18450,N_10814,N_13920);
nand U18451 (N_18451,N_13443,N_10267);
or U18452 (N_18452,N_10550,N_13148);
nor U18453 (N_18453,N_11934,N_10100);
xnor U18454 (N_18454,N_13157,N_14962);
nor U18455 (N_18455,N_14167,N_12103);
and U18456 (N_18456,N_11313,N_13130);
or U18457 (N_18457,N_10441,N_10109);
nand U18458 (N_18458,N_13522,N_14910);
or U18459 (N_18459,N_10845,N_14673);
xnor U18460 (N_18460,N_12330,N_10374);
or U18461 (N_18461,N_10496,N_10909);
or U18462 (N_18462,N_14420,N_12823);
xnor U18463 (N_18463,N_10240,N_13820);
and U18464 (N_18464,N_12794,N_11008);
xor U18465 (N_18465,N_14120,N_10467);
nand U18466 (N_18466,N_14525,N_14233);
and U18467 (N_18467,N_11299,N_12307);
or U18468 (N_18468,N_12680,N_12188);
nand U18469 (N_18469,N_14128,N_10138);
nor U18470 (N_18470,N_14452,N_13044);
nand U18471 (N_18471,N_12470,N_12914);
nor U18472 (N_18472,N_11988,N_14321);
or U18473 (N_18473,N_12667,N_13412);
nor U18474 (N_18474,N_14877,N_10097);
xor U18475 (N_18475,N_11005,N_10839);
or U18476 (N_18476,N_13658,N_10367);
and U18477 (N_18477,N_14615,N_10160);
or U18478 (N_18478,N_11878,N_14846);
and U18479 (N_18479,N_10668,N_14325);
and U18480 (N_18480,N_13396,N_11306);
nand U18481 (N_18481,N_11262,N_10460);
xor U18482 (N_18482,N_10805,N_12424);
xnor U18483 (N_18483,N_14945,N_13610);
and U18484 (N_18484,N_11654,N_14249);
or U18485 (N_18485,N_10990,N_12568);
or U18486 (N_18486,N_14515,N_14022);
and U18487 (N_18487,N_11005,N_14735);
and U18488 (N_18488,N_11438,N_12961);
or U18489 (N_18489,N_12720,N_14315);
nand U18490 (N_18490,N_14343,N_11431);
nor U18491 (N_18491,N_11830,N_12497);
nand U18492 (N_18492,N_11869,N_10014);
or U18493 (N_18493,N_13429,N_13300);
nor U18494 (N_18494,N_13878,N_13676);
nand U18495 (N_18495,N_13193,N_14477);
nand U18496 (N_18496,N_14080,N_13357);
xor U18497 (N_18497,N_12882,N_13217);
and U18498 (N_18498,N_14745,N_10637);
and U18499 (N_18499,N_12129,N_10630);
nand U18500 (N_18500,N_14877,N_10843);
xor U18501 (N_18501,N_10256,N_12701);
xnor U18502 (N_18502,N_11305,N_10378);
or U18503 (N_18503,N_14859,N_11948);
or U18504 (N_18504,N_12355,N_11945);
xnor U18505 (N_18505,N_12048,N_14800);
nand U18506 (N_18506,N_10075,N_10135);
xor U18507 (N_18507,N_14164,N_13994);
or U18508 (N_18508,N_14981,N_13778);
nand U18509 (N_18509,N_13003,N_12208);
nand U18510 (N_18510,N_13735,N_11593);
and U18511 (N_18511,N_11256,N_13867);
nor U18512 (N_18512,N_13082,N_10723);
nand U18513 (N_18513,N_14381,N_12092);
nand U18514 (N_18514,N_13982,N_13222);
xor U18515 (N_18515,N_14765,N_14155);
nor U18516 (N_18516,N_12064,N_12305);
xnor U18517 (N_18517,N_10830,N_12474);
nor U18518 (N_18518,N_12959,N_11868);
and U18519 (N_18519,N_11396,N_14284);
xnor U18520 (N_18520,N_14611,N_12659);
nor U18521 (N_18521,N_12739,N_11482);
nand U18522 (N_18522,N_13965,N_14868);
or U18523 (N_18523,N_13564,N_12007);
or U18524 (N_18524,N_11662,N_12265);
and U18525 (N_18525,N_12424,N_12356);
nand U18526 (N_18526,N_13667,N_14070);
nor U18527 (N_18527,N_13791,N_11593);
and U18528 (N_18528,N_10786,N_11565);
xor U18529 (N_18529,N_14010,N_14019);
nor U18530 (N_18530,N_12102,N_13351);
nor U18531 (N_18531,N_10851,N_11443);
nor U18532 (N_18532,N_10213,N_10252);
nand U18533 (N_18533,N_14312,N_14849);
and U18534 (N_18534,N_12043,N_10310);
xor U18535 (N_18535,N_13465,N_13966);
nor U18536 (N_18536,N_10140,N_13275);
nor U18537 (N_18537,N_13689,N_14309);
nor U18538 (N_18538,N_13099,N_11250);
and U18539 (N_18539,N_10102,N_14452);
and U18540 (N_18540,N_11246,N_11510);
and U18541 (N_18541,N_13873,N_11991);
xor U18542 (N_18542,N_11389,N_12225);
nor U18543 (N_18543,N_14087,N_12257);
and U18544 (N_18544,N_13146,N_13618);
xnor U18545 (N_18545,N_14299,N_11608);
and U18546 (N_18546,N_11496,N_11628);
or U18547 (N_18547,N_11820,N_11198);
nand U18548 (N_18548,N_11910,N_14111);
xor U18549 (N_18549,N_13518,N_12148);
nand U18550 (N_18550,N_10596,N_11159);
nand U18551 (N_18551,N_13491,N_14462);
nor U18552 (N_18552,N_12286,N_14323);
xnor U18553 (N_18553,N_13608,N_10001);
or U18554 (N_18554,N_10057,N_13893);
xnor U18555 (N_18555,N_11164,N_13143);
nand U18556 (N_18556,N_13943,N_12761);
xnor U18557 (N_18557,N_11862,N_12134);
nor U18558 (N_18558,N_10160,N_13176);
or U18559 (N_18559,N_10994,N_14431);
nor U18560 (N_18560,N_10664,N_14056);
nor U18561 (N_18561,N_14514,N_12650);
or U18562 (N_18562,N_12509,N_11774);
and U18563 (N_18563,N_12762,N_14484);
nand U18564 (N_18564,N_10731,N_11779);
nand U18565 (N_18565,N_13432,N_14544);
xnor U18566 (N_18566,N_12732,N_13408);
xor U18567 (N_18567,N_11379,N_11500);
and U18568 (N_18568,N_11622,N_13823);
or U18569 (N_18569,N_11462,N_14576);
nor U18570 (N_18570,N_10048,N_13900);
and U18571 (N_18571,N_13369,N_14794);
nand U18572 (N_18572,N_14879,N_12893);
and U18573 (N_18573,N_10230,N_11125);
xnor U18574 (N_18574,N_12190,N_10931);
or U18575 (N_18575,N_13297,N_13008);
xnor U18576 (N_18576,N_12123,N_14448);
xor U18577 (N_18577,N_14059,N_11276);
nand U18578 (N_18578,N_13501,N_12015);
or U18579 (N_18579,N_14033,N_13619);
nand U18580 (N_18580,N_10619,N_14527);
nor U18581 (N_18581,N_14338,N_10764);
nor U18582 (N_18582,N_10360,N_12661);
nand U18583 (N_18583,N_11160,N_10350);
nor U18584 (N_18584,N_12837,N_13189);
or U18585 (N_18585,N_12156,N_11637);
and U18586 (N_18586,N_12360,N_11770);
nand U18587 (N_18587,N_12784,N_12642);
nand U18588 (N_18588,N_10295,N_13554);
xnor U18589 (N_18589,N_12862,N_13698);
nand U18590 (N_18590,N_10537,N_14853);
nand U18591 (N_18591,N_13333,N_11488);
and U18592 (N_18592,N_13018,N_12359);
nand U18593 (N_18593,N_10268,N_10798);
or U18594 (N_18594,N_10841,N_11729);
nor U18595 (N_18595,N_10806,N_12486);
xor U18596 (N_18596,N_14529,N_10116);
xnor U18597 (N_18597,N_14937,N_12278);
and U18598 (N_18598,N_12678,N_13982);
and U18599 (N_18599,N_13941,N_11180);
nor U18600 (N_18600,N_11175,N_13600);
or U18601 (N_18601,N_13415,N_10168);
nor U18602 (N_18602,N_13516,N_12043);
xnor U18603 (N_18603,N_14077,N_14391);
nand U18604 (N_18604,N_13862,N_10347);
nand U18605 (N_18605,N_13604,N_10089);
xnor U18606 (N_18606,N_12658,N_13667);
nand U18607 (N_18607,N_10997,N_14785);
nor U18608 (N_18608,N_10184,N_14729);
or U18609 (N_18609,N_10562,N_14839);
and U18610 (N_18610,N_11155,N_13564);
nor U18611 (N_18611,N_12132,N_12987);
or U18612 (N_18612,N_11999,N_11021);
nor U18613 (N_18613,N_14623,N_13327);
nor U18614 (N_18614,N_12757,N_10914);
nor U18615 (N_18615,N_13312,N_14896);
or U18616 (N_18616,N_12702,N_14504);
or U18617 (N_18617,N_10874,N_13965);
or U18618 (N_18618,N_13254,N_12713);
and U18619 (N_18619,N_11545,N_11363);
nand U18620 (N_18620,N_11920,N_13354);
xor U18621 (N_18621,N_13561,N_14733);
nor U18622 (N_18622,N_12508,N_13885);
or U18623 (N_18623,N_14657,N_14757);
nor U18624 (N_18624,N_12805,N_13597);
and U18625 (N_18625,N_10596,N_14536);
nor U18626 (N_18626,N_10515,N_11576);
nand U18627 (N_18627,N_13320,N_11436);
or U18628 (N_18628,N_10630,N_14944);
nand U18629 (N_18629,N_10242,N_14587);
nand U18630 (N_18630,N_13970,N_13288);
nor U18631 (N_18631,N_14879,N_14512);
and U18632 (N_18632,N_10090,N_10783);
xor U18633 (N_18633,N_12427,N_14111);
nor U18634 (N_18634,N_14525,N_11553);
and U18635 (N_18635,N_14070,N_11161);
nor U18636 (N_18636,N_11201,N_13000);
nand U18637 (N_18637,N_11448,N_10951);
nand U18638 (N_18638,N_13167,N_11399);
and U18639 (N_18639,N_12613,N_11095);
nor U18640 (N_18640,N_12185,N_11886);
nor U18641 (N_18641,N_10599,N_12582);
xor U18642 (N_18642,N_10549,N_14464);
or U18643 (N_18643,N_10083,N_13221);
and U18644 (N_18644,N_12992,N_13380);
xor U18645 (N_18645,N_11932,N_11141);
xnor U18646 (N_18646,N_12419,N_13330);
or U18647 (N_18647,N_10164,N_10705);
nor U18648 (N_18648,N_14747,N_13805);
and U18649 (N_18649,N_12326,N_11075);
and U18650 (N_18650,N_13446,N_13989);
and U18651 (N_18651,N_14216,N_12503);
or U18652 (N_18652,N_10548,N_13564);
or U18653 (N_18653,N_11212,N_13398);
and U18654 (N_18654,N_11640,N_14531);
nor U18655 (N_18655,N_11816,N_11576);
nor U18656 (N_18656,N_13154,N_11715);
and U18657 (N_18657,N_13682,N_10623);
and U18658 (N_18658,N_13467,N_10212);
and U18659 (N_18659,N_10620,N_10557);
nand U18660 (N_18660,N_10774,N_13512);
xor U18661 (N_18661,N_10431,N_14210);
or U18662 (N_18662,N_12220,N_14660);
or U18663 (N_18663,N_12138,N_10573);
or U18664 (N_18664,N_11102,N_13630);
xor U18665 (N_18665,N_14630,N_11039);
nor U18666 (N_18666,N_11370,N_13856);
and U18667 (N_18667,N_14196,N_13955);
and U18668 (N_18668,N_12638,N_10623);
and U18669 (N_18669,N_13535,N_13838);
xor U18670 (N_18670,N_11789,N_10402);
nand U18671 (N_18671,N_11366,N_14077);
nor U18672 (N_18672,N_14048,N_11812);
nor U18673 (N_18673,N_12461,N_11133);
and U18674 (N_18674,N_14259,N_10812);
and U18675 (N_18675,N_13699,N_14257);
nand U18676 (N_18676,N_11886,N_14385);
or U18677 (N_18677,N_13607,N_14746);
xor U18678 (N_18678,N_11808,N_14611);
and U18679 (N_18679,N_13752,N_12441);
or U18680 (N_18680,N_13506,N_14611);
nor U18681 (N_18681,N_11599,N_12334);
nor U18682 (N_18682,N_11300,N_14274);
or U18683 (N_18683,N_14153,N_10798);
nand U18684 (N_18684,N_11424,N_12840);
and U18685 (N_18685,N_11431,N_14955);
nand U18686 (N_18686,N_13726,N_12246);
nor U18687 (N_18687,N_13168,N_11602);
nor U18688 (N_18688,N_14379,N_12629);
nor U18689 (N_18689,N_13890,N_14464);
and U18690 (N_18690,N_14853,N_14365);
nor U18691 (N_18691,N_13396,N_14535);
nand U18692 (N_18692,N_13963,N_11570);
nand U18693 (N_18693,N_10185,N_11410);
nand U18694 (N_18694,N_10648,N_10901);
nor U18695 (N_18695,N_10477,N_11731);
or U18696 (N_18696,N_14332,N_11116);
or U18697 (N_18697,N_12250,N_12841);
or U18698 (N_18698,N_10963,N_11238);
and U18699 (N_18699,N_13959,N_14720);
or U18700 (N_18700,N_12387,N_14645);
nor U18701 (N_18701,N_12997,N_12538);
nor U18702 (N_18702,N_11529,N_12096);
nor U18703 (N_18703,N_13963,N_14818);
or U18704 (N_18704,N_10586,N_12454);
xnor U18705 (N_18705,N_14875,N_10593);
nand U18706 (N_18706,N_11376,N_11155);
xnor U18707 (N_18707,N_13407,N_12703);
nor U18708 (N_18708,N_12304,N_12138);
xnor U18709 (N_18709,N_13620,N_11379);
xor U18710 (N_18710,N_13093,N_10392);
xor U18711 (N_18711,N_11585,N_10324);
xor U18712 (N_18712,N_10011,N_12324);
nand U18713 (N_18713,N_14965,N_10902);
xnor U18714 (N_18714,N_12175,N_12324);
nor U18715 (N_18715,N_12841,N_12496);
xnor U18716 (N_18716,N_13731,N_12159);
nand U18717 (N_18717,N_10922,N_12146);
or U18718 (N_18718,N_14590,N_12253);
or U18719 (N_18719,N_14942,N_13169);
nand U18720 (N_18720,N_14716,N_12019);
or U18721 (N_18721,N_14203,N_14694);
or U18722 (N_18722,N_10084,N_12123);
and U18723 (N_18723,N_10536,N_10691);
nor U18724 (N_18724,N_10241,N_11505);
nor U18725 (N_18725,N_12172,N_13133);
nor U18726 (N_18726,N_11463,N_10538);
xnor U18727 (N_18727,N_12934,N_14845);
xor U18728 (N_18728,N_11547,N_11112);
or U18729 (N_18729,N_14198,N_12932);
nand U18730 (N_18730,N_11727,N_14522);
nor U18731 (N_18731,N_14167,N_11713);
or U18732 (N_18732,N_13333,N_11823);
nand U18733 (N_18733,N_12358,N_11178);
nor U18734 (N_18734,N_11151,N_11084);
nand U18735 (N_18735,N_10105,N_11622);
nor U18736 (N_18736,N_14998,N_14496);
nor U18737 (N_18737,N_11637,N_11208);
and U18738 (N_18738,N_13283,N_12842);
and U18739 (N_18739,N_12312,N_13016);
or U18740 (N_18740,N_10498,N_10220);
nand U18741 (N_18741,N_14487,N_11408);
or U18742 (N_18742,N_13128,N_13190);
nor U18743 (N_18743,N_13254,N_11889);
nor U18744 (N_18744,N_12513,N_13283);
nand U18745 (N_18745,N_10378,N_11340);
nand U18746 (N_18746,N_12543,N_13902);
and U18747 (N_18747,N_11729,N_10688);
xnor U18748 (N_18748,N_12654,N_11024);
xnor U18749 (N_18749,N_14396,N_12437);
and U18750 (N_18750,N_14366,N_10526);
xor U18751 (N_18751,N_14517,N_11444);
xnor U18752 (N_18752,N_11966,N_12772);
nor U18753 (N_18753,N_13428,N_11683);
or U18754 (N_18754,N_12629,N_12668);
nand U18755 (N_18755,N_11575,N_14139);
and U18756 (N_18756,N_12114,N_12667);
or U18757 (N_18757,N_11295,N_14564);
xnor U18758 (N_18758,N_13751,N_11012);
nand U18759 (N_18759,N_11181,N_12851);
and U18760 (N_18760,N_10042,N_14003);
nor U18761 (N_18761,N_14637,N_10669);
or U18762 (N_18762,N_12090,N_12275);
and U18763 (N_18763,N_13156,N_13309);
and U18764 (N_18764,N_10638,N_12100);
xor U18765 (N_18765,N_14252,N_11595);
nor U18766 (N_18766,N_12376,N_14688);
nand U18767 (N_18767,N_11026,N_10633);
and U18768 (N_18768,N_14153,N_10486);
and U18769 (N_18769,N_13226,N_14465);
nand U18770 (N_18770,N_14439,N_13272);
nand U18771 (N_18771,N_14741,N_11303);
nor U18772 (N_18772,N_12426,N_14354);
nor U18773 (N_18773,N_12200,N_10443);
xnor U18774 (N_18774,N_11696,N_11032);
and U18775 (N_18775,N_10508,N_14621);
xor U18776 (N_18776,N_10825,N_12096);
or U18777 (N_18777,N_12068,N_14491);
xnor U18778 (N_18778,N_10569,N_11365);
nand U18779 (N_18779,N_13634,N_13630);
nand U18780 (N_18780,N_13573,N_12178);
nand U18781 (N_18781,N_10957,N_14654);
and U18782 (N_18782,N_10150,N_11569);
or U18783 (N_18783,N_12459,N_10437);
nand U18784 (N_18784,N_14010,N_10864);
nand U18785 (N_18785,N_11701,N_11481);
nor U18786 (N_18786,N_13599,N_10900);
or U18787 (N_18787,N_13145,N_13013);
xor U18788 (N_18788,N_14766,N_10715);
or U18789 (N_18789,N_12751,N_13249);
nor U18790 (N_18790,N_11120,N_14935);
xor U18791 (N_18791,N_14676,N_11688);
xnor U18792 (N_18792,N_10251,N_10518);
and U18793 (N_18793,N_14831,N_11928);
or U18794 (N_18794,N_13611,N_14970);
nor U18795 (N_18795,N_11393,N_13425);
and U18796 (N_18796,N_10487,N_13449);
xor U18797 (N_18797,N_12098,N_14838);
or U18798 (N_18798,N_12065,N_14212);
or U18799 (N_18799,N_14079,N_12298);
xor U18800 (N_18800,N_12766,N_13691);
nand U18801 (N_18801,N_10202,N_14994);
nor U18802 (N_18802,N_12676,N_14815);
xor U18803 (N_18803,N_10504,N_10818);
nor U18804 (N_18804,N_12153,N_14201);
nor U18805 (N_18805,N_12326,N_11307);
nor U18806 (N_18806,N_10685,N_13119);
xnor U18807 (N_18807,N_14058,N_12282);
and U18808 (N_18808,N_11040,N_12468);
nand U18809 (N_18809,N_13937,N_11042);
and U18810 (N_18810,N_11126,N_12612);
and U18811 (N_18811,N_11845,N_10423);
and U18812 (N_18812,N_12891,N_11309);
or U18813 (N_18813,N_11457,N_11297);
and U18814 (N_18814,N_11781,N_10741);
nor U18815 (N_18815,N_12489,N_10527);
xor U18816 (N_18816,N_13266,N_13085);
and U18817 (N_18817,N_11446,N_13793);
xnor U18818 (N_18818,N_12034,N_14676);
nor U18819 (N_18819,N_14879,N_11161);
and U18820 (N_18820,N_11298,N_12593);
nor U18821 (N_18821,N_11847,N_14561);
and U18822 (N_18822,N_12133,N_13993);
and U18823 (N_18823,N_10396,N_13504);
xor U18824 (N_18824,N_13137,N_11994);
nor U18825 (N_18825,N_11403,N_14794);
nor U18826 (N_18826,N_11530,N_14966);
nor U18827 (N_18827,N_12823,N_13732);
nor U18828 (N_18828,N_12565,N_13078);
xor U18829 (N_18829,N_12453,N_14252);
and U18830 (N_18830,N_11854,N_13072);
or U18831 (N_18831,N_12404,N_10103);
nor U18832 (N_18832,N_13687,N_12956);
or U18833 (N_18833,N_11902,N_11738);
nand U18834 (N_18834,N_11691,N_14090);
nand U18835 (N_18835,N_12426,N_11227);
or U18836 (N_18836,N_10116,N_12313);
nor U18837 (N_18837,N_14838,N_13526);
or U18838 (N_18838,N_14556,N_10772);
nor U18839 (N_18839,N_11502,N_14447);
nor U18840 (N_18840,N_10132,N_14306);
nor U18841 (N_18841,N_12646,N_14979);
nand U18842 (N_18842,N_12936,N_13570);
xnor U18843 (N_18843,N_10684,N_11472);
or U18844 (N_18844,N_12300,N_10295);
xnor U18845 (N_18845,N_13833,N_10880);
nand U18846 (N_18846,N_11518,N_14265);
xor U18847 (N_18847,N_10558,N_13034);
xnor U18848 (N_18848,N_13115,N_10065);
nand U18849 (N_18849,N_12318,N_14976);
nor U18850 (N_18850,N_14551,N_10700);
xnor U18851 (N_18851,N_11550,N_14272);
or U18852 (N_18852,N_13739,N_10248);
and U18853 (N_18853,N_10749,N_11962);
xnor U18854 (N_18854,N_11132,N_10633);
nand U18855 (N_18855,N_12776,N_11189);
and U18856 (N_18856,N_11069,N_11298);
nor U18857 (N_18857,N_10001,N_14169);
nor U18858 (N_18858,N_14773,N_11895);
xor U18859 (N_18859,N_10314,N_13174);
xor U18860 (N_18860,N_10327,N_10642);
xnor U18861 (N_18861,N_10833,N_12336);
nor U18862 (N_18862,N_12157,N_12137);
xor U18863 (N_18863,N_12631,N_14200);
xnor U18864 (N_18864,N_14945,N_13122);
or U18865 (N_18865,N_10218,N_13915);
and U18866 (N_18866,N_12861,N_14808);
nand U18867 (N_18867,N_13466,N_12263);
and U18868 (N_18868,N_10959,N_11628);
nand U18869 (N_18869,N_11802,N_12286);
and U18870 (N_18870,N_13662,N_13954);
nor U18871 (N_18871,N_13059,N_14719);
or U18872 (N_18872,N_11167,N_12489);
and U18873 (N_18873,N_14868,N_12768);
and U18874 (N_18874,N_13122,N_14556);
xnor U18875 (N_18875,N_11128,N_12205);
xnor U18876 (N_18876,N_11994,N_14274);
nor U18877 (N_18877,N_12893,N_14301);
or U18878 (N_18878,N_12481,N_12733);
nor U18879 (N_18879,N_11496,N_13967);
or U18880 (N_18880,N_10769,N_12019);
xor U18881 (N_18881,N_14194,N_11917);
nor U18882 (N_18882,N_13278,N_13519);
nor U18883 (N_18883,N_10888,N_11601);
nor U18884 (N_18884,N_10824,N_13004);
nor U18885 (N_18885,N_11905,N_14432);
nor U18886 (N_18886,N_13113,N_11477);
and U18887 (N_18887,N_10707,N_12947);
nand U18888 (N_18888,N_13957,N_12204);
and U18889 (N_18889,N_13494,N_11764);
and U18890 (N_18890,N_14280,N_11174);
or U18891 (N_18891,N_12723,N_10314);
nand U18892 (N_18892,N_11103,N_11221);
nand U18893 (N_18893,N_12249,N_11529);
and U18894 (N_18894,N_13849,N_10326);
or U18895 (N_18895,N_10642,N_12878);
xnor U18896 (N_18896,N_14822,N_11180);
nor U18897 (N_18897,N_14746,N_12700);
or U18898 (N_18898,N_13952,N_13215);
nand U18899 (N_18899,N_14293,N_14794);
and U18900 (N_18900,N_11325,N_14732);
or U18901 (N_18901,N_11850,N_11188);
nor U18902 (N_18902,N_12335,N_11193);
nand U18903 (N_18903,N_14061,N_10314);
nand U18904 (N_18904,N_14299,N_11545);
xor U18905 (N_18905,N_10622,N_10314);
or U18906 (N_18906,N_11519,N_12727);
and U18907 (N_18907,N_11047,N_14517);
nand U18908 (N_18908,N_10096,N_12292);
nand U18909 (N_18909,N_12536,N_12663);
xnor U18910 (N_18910,N_13461,N_14718);
xnor U18911 (N_18911,N_13558,N_13459);
xor U18912 (N_18912,N_11722,N_13981);
nor U18913 (N_18913,N_14903,N_12989);
xnor U18914 (N_18914,N_12641,N_13889);
nor U18915 (N_18915,N_13256,N_11111);
or U18916 (N_18916,N_13365,N_10349);
xor U18917 (N_18917,N_11799,N_12495);
and U18918 (N_18918,N_11543,N_14721);
and U18919 (N_18919,N_10671,N_13175);
nor U18920 (N_18920,N_11662,N_11688);
nand U18921 (N_18921,N_14859,N_13751);
nor U18922 (N_18922,N_12631,N_11625);
and U18923 (N_18923,N_10185,N_10527);
nand U18924 (N_18924,N_10872,N_11431);
xnor U18925 (N_18925,N_10037,N_14089);
or U18926 (N_18926,N_13940,N_13768);
nand U18927 (N_18927,N_14179,N_13688);
nand U18928 (N_18928,N_13640,N_11930);
and U18929 (N_18929,N_10223,N_14812);
and U18930 (N_18930,N_10561,N_14276);
nand U18931 (N_18931,N_11172,N_10209);
and U18932 (N_18932,N_10314,N_11402);
nor U18933 (N_18933,N_14826,N_10687);
nor U18934 (N_18934,N_12261,N_10305);
and U18935 (N_18935,N_12724,N_14160);
xnor U18936 (N_18936,N_14617,N_14515);
and U18937 (N_18937,N_11287,N_10936);
nand U18938 (N_18938,N_11098,N_10064);
xor U18939 (N_18939,N_13900,N_10985);
nand U18940 (N_18940,N_14259,N_12649);
nor U18941 (N_18941,N_10930,N_14444);
and U18942 (N_18942,N_11546,N_12040);
and U18943 (N_18943,N_13992,N_13491);
xor U18944 (N_18944,N_14173,N_11200);
and U18945 (N_18945,N_12559,N_10405);
and U18946 (N_18946,N_11951,N_10207);
xnor U18947 (N_18947,N_13678,N_12212);
nor U18948 (N_18948,N_12358,N_10521);
or U18949 (N_18949,N_11928,N_13319);
or U18950 (N_18950,N_13665,N_13633);
nor U18951 (N_18951,N_14714,N_12962);
nand U18952 (N_18952,N_14246,N_14363);
or U18953 (N_18953,N_13842,N_14467);
nor U18954 (N_18954,N_12122,N_12658);
and U18955 (N_18955,N_12150,N_11278);
nand U18956 (N_18956,N_14233,N_14713);
nor U18957 (N_18957,N_13932,N_10685);
and U18958 (N_18958,N_12077,N_14480);
xor U18959 (N_18959,N_11283,N_14064);
or U18960 (N_18960,N_14499,N_11370);
or U18961 (N_18961,N_10043,N_14326);
or U18962 (N_18962,N_14590,N_11617);
xnor U18963 (N_18963,N_11009,N_10927);
or U18964 (N_18964,N_14698,N_11425);
and U18965 (N_18965,N_11579,N_10405);
xnor U18966 (N_18966,N_10758,N_12620);
xnor U18967 (N_18967,N_13597,N_11966);
nor U18968 (N_18968,N_11845,N_14433);
nand U18969 (N_18969,N_14166,N_10573);
nor U18970 (N_18970,N_14620,N_11290);
nor U18971 (N_18971,N_10122,N_11727);
and U18972 (N_18972,N_10043,N_11932);
or U18973 (N_18973,N_12750,N_14626);
nand U18974 (N_18974,N_13694,N_10476);
xnor U18975 (N_18975,N_14989,N_10429);
and U18976 (N_18976,N_13583,N_10960);
or U18977 (N_18977,N_12048,N_14950);
or U18978 (N_18978,N_12575,N_13562);
or U18979 (N_18979,N_12660,N_11249);
and U18980 (N_18980,N_14035,N_12162);
xnor U18981 (N_18981,N_13971,N_14203);
nor U18982 (N_18982,N_10650,N_10755);
or U18983 (N_18983,N_12995,N_13008);
xor U18984 (N_18984,N_10921,N_12654);
nor U18985 (N_18985,N_11321,N_11662);
xor U18986 (N_18986,N_11395,N_14291);
or U18987 (N_18987,N_13076,N_10676);
nand U18988 (N_18988,N_10338,N_10913);
nand U18989 (N_18989,N_10446,N_10696);
nand U18990 (N_18990,N_10481,N_11604);
nand U18991 (N_18991,N_14356,N_14213);
xnor U18992 (N_18992,N_10913,N_13091);
xnor U18993 (N_18993,N_10484,N_10718);
nor U18994 (N_18994,N_11563,N_12559);
xnor U18995 (N_18995,N_14324,N_13195);
nand U18996 (N_18996,N_12740,N_14546);
xor U18997 (N_18997,N_12583,N_10692);
xor U18998 (N_18998,N_11629,N_13613);
or U18999 (N_18999,N_14048,N_10275);
and U19000 (N_19000,N_14757,N_11553);
xnor U19001 (N_19001,N_11703,N_10104);
or U19002 (N_19002,N_14849,N_10765);
and U19003 (N_19003,N_11768,N_13497);
and U19004 (N_19004,N_12982,N_14972);
and U19005 (N_19005,N_14332,N_12019);
or U19006 (N_19006,N_14486,N_12060);
nor U19007 (N_19007,N_14715,N_13454);
xor U19008 (N_19008,N_10876,N_13195);
nand U19009 (N_19009,N_10419,N_11657);
xor U19010 (N_19010,N_13718,N_10214);
xor U19011 (N_19011,N_10698,N_13705);
xor U19012 (N_19012,N_10798,N_11523);
xnor U19013 (N_19013,N_14600,N_10606);
and U19014 (N_19014,N_13117,N_13868);
nor U19015 (N_19015,N_10316,N_13374);
and U19016 (N_19016,N_12806,N_13037);
nor U19017 (N_19017,N_11770,N_11698);
and U19018 (N_19018,N_10641,N_11022);
nand U19019 (N_19019,N_10569,N_11432);
and U19020 (N_19020,N_14269,N_14258);
or U19021 (N_19021,N_14266,N_12735);
nor U19022 (N_19022,N_13528,N_11692);
xor U19023 (N_19023,N_10991,N_12403);
nor U19024 (N_19024,N_13393,N_13079);
and U19025 (N_19025,N_12896,N_10442);
or U19026 (N_19026,N_10879,N_11184);
and U19027 (N_19027,N_11718,N_13401);
or U19028 (N_19028,N_12056,N_10514);
or U19029 (N_19029,N_13140,N_14095);
or U19030 (N_19030,N_10573,N_14783);
xor U19031 (N_19031,N_13656,N_11450);
nor U19032 (N_19032,N_10840,N_11483);
nor U19033 (N_19033,N_11035,N_11096);
nor U19034 (N_19034,N_13443,N_11835);
or U19035 (N_19035,N_12325,N_13446);
xnor U19036 (N_19036,N_13246,N_11525);
nand U19037 (N_19037,N_13377,N_12221);
xnor U19038 (N_19038,N_13778,N_14034);
or U19039 (N_19039,N_14733,N_11252);
nand U19040 (N_19040,N_13520,N_10324);
and U19041 (N_19041,N_12096,N_12163);
nand U19042 (N_19042,N_14635,N_13585);
and U19043 (N_19043,N_11284,N_14741);
nor U19044 (N_19044,N_14173,N_14957);
nand U19045 (N_19045,N_12943,N_11052);
and U19046 (N_19046,N_11522,N_13540);
nand U19047 (N_19047,N_11120,N_12242);
xor U19048 (N_19048,N_12505,N_11904);
nand U19049 (N_19049,N_12214,N_14854);
nand U19050 (N_19050,N_14154,N_10337);
nand U19051 (N_19051,N_12954,N_14742);
xor U19052 (N_19052,N_14473,N_11040);
xor U19053 (N_19053,N_12414,N_10474);
nand U19054 (N_19054,N_11942,N_13196);
nand U19055 (N_19055,N_14070,N_10114);
or U19056 (N_19056,N_13943,N_13781);
nor U19057 (N_19057,N_13908,N_10956);
nor U19058 (N_19058,N_12300,N_13897);
nor U19059 (N_19059,N_11194,N_13110);
nor U19060 (N_19060,N_12038,N_11034);
nand U19061 (N_19061,N_13921,N_10541);
or U19062 (N_19062,N_12179,N_13504);
or U19063 (N_19063,N_12212,N_13092);
or U19064 (N_19064,N_13410,N_10455);
nand U19065 (N_19065,N_13109,N_13439);
or U19066 (N_19066,N_11187,N_11947);
xnor U19067 (N_19067,N_11926,N_11277);
nand U19068 (N_19068,N_11817,N_11009);
nand U19069 (N_19069,N_11362,N_10298);
nand U19070 (N_19070,N_10914,N_12882);
or U19071 (N_19071,N_11517,N_11079);
xor U19072 (N_19072,N_14119,N_10184);
and U19073 (N_19073,N_12554,N_10857);
and U19074 (N_19074,N_13137,N_11710);
nor U19075 (N_19075,N_11359,N_13441);
nand U19076 (N_19076,N_13796,N_12075);
nand U19077 (N_19077,N_14920,N_10109);
nand U19078 (N_19078,N_13763,N_12227);
nor U19079 (N_19079,N_11138,N_14217);
xnor U19080 (N_19080,N_10547,N_13794);
xor U19081 (N_19081,N_14220,N_11579);
or U19082 (N_19082,N_12872,N_12084);
nand U19083 (N_19083,N_11935,N_11444);
or U19084 (N_19084,N_11536,N_14278);
and U19085 (N_19085,N_11099,N_11728);
nand U19086 (N_19086,N_10800,N_12001);
or U19087 (N_19087,N_14246,N_13658);
or U19088 (N_19088,N_13257,N_10205);
nor U19089 (N_19089,N_10824,N_14536);
and U19090 (N_19090,N_11052,N_12036);
nand U19091 (N_19091,N_12663,N_11084);
xnor U19092 (N_19092,N_10227,N_14282);
xor U19093 (N_19093,N_11850,N_11984);
nor U19094 (N_19094,N_14192,N_13790);
nor U19095 (N_19095,N_14284,N_12489);
and U19096 (N_19096,N_10097,N_10404);
or U19097 (N_19097,N_14239,N_10162);
nand U19098 (N_19098,N_13032,N_10308);
nand U19099 (N_19099,N_12568,N_12205);
or U19100 (N_19100,N_12178,N_13488);
or U19101 (N_19101,N_12150,N_13162);
xor U19102 (N_19102,N_13328,N_13132);
xor U19103 (N_19103,N_10359,N_13982);
xor U19104 (N_19104,N_11074,N_12520);
and U19105 (N_19105,N_14724,N_10769);
nor U19106 (N_19106,N_13749,N_11159);
or U19107 (N_19107,N_10770,N_11248);
nand U19108 (N_19108,N_14236,N_12925);
and U19109 (N_19109,N_11347,N_14732);
or U19110 (N_19110,N_14709,N_12942);
xor U19111 (N_19111,N_11789,N_12347);
or U19112 (N_19112,N_13547,N_13888);
and U19113 (N_19113,N_12264,N_11703);
nand U19114 (N_19114,N_10757,N_10023);
nor U19115 (N_19115,N_13706,N_12336);
or U19116 (N_19116,N_11589,N_14410);
nor U19117 (N_19117,N_12437,N_11008);
nor U19118 (N_19118,N_12675,N_13769);
nand U19119 (N_19119,N_10655,N_10735);
or U19120 (N_19120,N_13855,N_12659);
and U19121 (N_19121,N_13971,N_11621);
xnor U19122 (N_19122,N_14372,N_10839);
xor U19123 (N_19123,N_13985,N_14131);
xor U19124 (N_19124,N_12847,N_10878);
and U19125 (N_19125,N_13548,N_10705);
and U19126 (N_19126,N_13657,N_11209);
xor U19127 (N_19127,N_12434,N_10291);
xnor U19128 (N_19128,N_11713,N_14361);
xnor U19129 (N_19129,N_14949,N_14267);
xnor U19130 (N_19130,N_11338,N_12147);
or U19131 (N_19131,N_10451,N_14908);
nor U19132 (N_19132,N_10663,N_10436);
and U19133 (N_19133,N_10622,N_13529);
xor U19134 (N_19134,N_14728,N_11444);
and U19135 (N_19135,N_11435,N_13408);
and U19136 (N_19136,N_10538,N_11793);
xnor U19137 (N_19137,N_10705,N_13993);
or U19138 (N_19138,N_14027,N_11575);
or U19139 (N_19139,N_12849,N_11533);
nand U19140 (N_19140,N_13692,N_13940);
nor U19141 (N_19141,N_13291,N_13277);
nor U19142 (N_19142,N_10888,N_11026);
nor U19143 (N_19143,N_11293,N_14590);
xor U19144 (N_19144,N_10383,N_10372);
nand U19145 (N_19145,N_14596,N_12540);
or U19146 (N_19146,N_11394,N_10845);
xnor U19147 (N_19147,N_10452,N_12082);
xor U19148 (N_19148,N_13711,N_13251);
nor U19149 (N_19149,N_12074,N_11217);
nand U19150 (N_19150,N_11850,N_10000);
xnor U19151 (N_19151,N_14757,N_12230);
and U19152 (N_19152,N_13536,N_14270);
xnor U19153 (N_19153,N_14704,N_10583);
nor U19154 (N_19154,N_11127,N_14277);
or U19155 (N_19155,N_12928,N_11086);
xor U19156 (N_19156,N_14154,N_10819);
nor U19157 (N_19157,N_13405,N_12896);
and U19158 (N_19158,N_10344,N_12413);
or U19159 (N_19159,N_11331,N_13937);
or U19160 (N_19160,N_13328,N_13545);
or U19161 (N_19161,N_14884,N_12025);
and U19162 (N_19162,N_13450,N_11308);
nor U19163 (N_19163,N_14947,N_12362);
nor U19164 (N_19164,N_10870,N_14703);
and U19165 (N_19165,N_13734,N_12504);
xor U19166 (N_19166,N_11698,N_14617);
nor U19167 (N_19167,N_10233,N_14522);
nand U19168 (N_19168,N_10463,N_13319);
xor U19169 (N_19169,N_14806,N_14447);
or U19170 (N_19170,N_11727,N_14331);
nor U19171 (N_19171,N_13615,N_13238);
and U19172 (N_19172,N_11184,N_14276);
or U19173 (N_19173,N_10685,N_14424);
and U19174 (N_19174,N_13644,N_14379);
and U19175 (N_19175,N_13336,N_13752);
or U19176 (N_19176,N_11825,N_11976);
nand U19177 (N_19177,N_14079,N_10118);
or U19178 (N_19178,N_11254,N_12941);
xor U19179 (N_19179,N_14521,N_13085);
and U19180 (N_19180,N_13982,N_10584);
nor U19181 (N_19181,N_10318,N_12336);
nand U19182 (N_19182,N_13309,N_11876);
xor U19183 (N_19183,N_10125,N_12988);
xor U19184 (N_19184,N_10108,N_14652);
nand U19185 (N_19185,N_10230,N_10747);
nand U19186 (N_19186,N_11102,N_13180);
and U19187 (N_19187,N_12210,N_14583);
or U19188 (N_19188,N_14525,N_10014);
or U19189 (N_19189,N_13807,N_13148);
nand U19190 (N_19190,N_14724,N_13214);
nor U19191 (N_19191,N_12003,N_10393);
or U19192 (N_19192,N_14884,N_11381);
nand U19193 (N_19193,N_11869,N_13351);
xor U19194 (N_19194,N_14566,N_13849);
xnor U19195 (N_19195,N_10419,N_14652);
or U19196 (N_19196,N_10105,N_10320);
xor U19197 (N_19197,N_13800,N_12265);
nor U19198 (N_19198,N_11752,N_11830);
nor U19199 (N_19199,N_12426,N_14195);
or U19200 (N_19200,N_13241,N_12767);
nand U19201 (N_19201,N_14315,N_12394);
nor U19202 (N_19202,N_10350,N_12589);
xnor U19203 (N_19203,N_11127,N_10013);
nor U19204 (N_19204,N_11045,N_12314);
or U19205 (N_19205,N_12600,N_10862);
nor U19206 (N_19206,N_14432,N_13302);
nand U19207 (N_19207,N_12429,N_11172);
nand U19208 (N_19208,N_14034,N_12208);
and U19209 (N_19209,N_14065,N_13215);
or U19210 (N_19210,N_12024,N_14745);
nand U19211 (N_19211,N_13397,N_10338);
xnor U19212 (N_19212,N_14313,N_14425);
or U19213 (N_19213,N_12882,N_11484);
or U19214 (N_19214,N_12054,N_13214);
xnor U19215 (N_19215,N_11941,N_10384);
and U19216 (N_19216,N_10873,N_14249);
or U19217 (N_19217,N_14021,N_13770);
xnor U19218 (N_19218,N_10975,N_12604);
xor U19219 (N_19219,N_11392,N_11175);
or U19220 (N_19220,N_11408,N_12814);
or U19221 (N_19221,N_13635,N_12169);
and U19222 (N_19222,N_11300,N_13840);
nor U19223 (N_19223,N_10762,N_12318);
or U19224 (N_19224,N_11483,N_10046);
nand U19225 (N_19225,N_13032,N_11867);
nand U19226 (N_19226,N_10106,N_13080);
nand U19227 (N_19227,N_10521,N_13704);
xnor U19228 (N_19228,N_14612,N_12825);
and U19229 (N_19229,N_12255,N_11573);
and U19230 (N_19230,N_11428,N_14030);
xnor U19231 (N_19231,N_11007,N_12106);
and U19232 (N_19232,N_12757,N_13889);
nand U19233 (N_19233,N_14178,N_11910);
xnor U19234 (N_19234,N_13132,N_10825);
and U19235 (N_19235,N_12496,N_13252);
and U19236 (N_19236,N_10520,N_14823);
nor U19237 (N_19237,N_14717,N_12067);
or U19238 (N_19238,N_13023,N_10808);
and U19239 (N_19239,N_13301,N_11769);
xnor U19240 (N_19240,N_11138,N_12971);
nor U19241 (N_19241,N_11446,N_12210);
or U19242 (N_19242,N_14964,N_10069);
nand U19243 (N_19243,N_11665,N_10706);
or U19244 (N_19244,N_12105,N_11371);
or U19245 (N_19245,N_11008,N_10490);
and U19246 (N_19246,N_11416,N_11223);
or U19247 (N_19247,N_14767,N_11951);
nand U19248 (N_19248,N_10924,N_11072);
or U19249 (N_19249,N_14054,N_13629);
xor U19250 (N_19250,N_14456,N_10829);
and U19251 (N_19251,N_11462,N_13328);
nand U19252 (N_19252,N_10814,N_10496);
nor U19253 (N_19253,N_10308,N_14110);
xor U19254 (N_19254,N_10092,N_11101);
nand U19255 (N_19255,N_14424,N_14817);
nand U19256 (N_19256,N_13782,N_14556);
xor U19257 (N_19257,N_11623,N_10633);
or U19258 (N_19258,N_12223,N_14448);
xnor U19259 (N_19259,N_11307,N_10503);
or U19260 (N_19260,N_13917,N_12156);
or U19261 (N_19261,N_12528,N_12337);
and U19262 (N_19262,N_11677,N_12829);
and U19263 (N_19263,N_12984,N_12037);
or U19264 (N_19264,N_10075,N_11287);
xnor U19265 (N_19265,N_10315,N_14445);
and U19266 (N_19266,N_10677,N_10837);
nand U19267 (N_19267,N_11006,N_12254);
nand U19268 (N_19268,N_12828,N_10260);
nor U19269 (N_19269,N_14485,N_11839);
xnor U19270 (N_19270,N_11146,N_11766);
nor U19271 (N_19271,N_10457,N_10124);
nor U19272 (N_19272,N_14937,N_11060);
and U19273 (N_19273,N_10010,N_13297);
and U19274 (N_19274,N_11003,N_11932);
nand U19275 (N_19275,N_13927,N_14435);
or U19276 (N_19276,N_11058,N_12895);
nand U19277 (N_19277,N_10490,N_13497);
or U19278 (N_19278,N_10070,N_14682);
or U19279 (N_19279,N_13240,N_14486);
xnor U19280 (N_19280,N_10649,N_10794);
nor U19281 (N_19281,N_12620,N_10399);
or U19282 (N_19282,N_14524,N_10392);
xnor U19283 (N_19283,N_14679,N_12238);
xnor U19284 (N_19284,N_12984,N_13649);
nand U19285 (N_19285,N_12923,N_14891);
or U19286 (N_19286,N_14367,N_11025);
xnor U19287 (N_19287,N_13332,N_12279);
or U19288 (N_19288,N_12922,N_14360);
or U19289 (N_19289,N_11515,N_10619);
or U19290 (N_19290,N_13394,N_12992);
xnor U19291 (N_19291,N_14216,N_13038);
nor U19292 (N_19292,N_14330,N_12364);
nor U19293 (N_19293,N_11365,N_11124);
xnor U19294 (N_19294,N_14006,N_14843);
xnor U19295 (N_19295,N_14536,N_10147);
or U19296 (N_19296,N_10610,N_14075);
and U19297 (N_19297,N_11390,N_12191);
nor U19298 (N_19298,N_12937,N_14153);
xnor U19299 (N_19299,N_13876,N_12360);
or U19300 (N_19300,N_13199,N_13526);
or U19301 (N_19301,N_10010,N_13660);
and U19302 (N_19302,N_14145,N_12809);
and U19303 (N_19303,N_11807,N_11939);
xnor U19304 (N_19304,N_12289,N_12366);
nor U19305 (N_19305,N_14019,N_11926);
or U19306 (N_19306,N_12461,N_10628);
nor U19307 (N_19307,N_14910,N_11208);
xor U19308 (N_19308,N_10921,N_11955);
or U19309 (N_19309,N_12437,N_14795);
or U19310 (N_19310,N_14285,N_14127);
xnor U19311 (N_19311,N_14844,N_11122);
nand U19312 (N_19312,N_10204,N_11579);
nand U19313 (N_19313,N_14349,N_13612);
or U19314 (N_19314,N_10607,N_12547);
or U19315 (N_19315,N_14193,N_10989);
and U19316 (N_19316,N_10508,N_13360);
and U19317 (N_19317,N_10882,N_14447);
xnor U19318 (N_19318,N_13635,N_12816);
nand U19319 (N_19319,N_14080,N_14450);
nor U19320 (N_19320,N_11241,N_12978);
xnor U19321 (N_19321,N_10072,N_13929);
and U19322 (N_19322,N_10521,N_11196);
or U19323 (N_19323,N_10229,N_11390);
nor U19324 (N_19324,N_10633,N_14135);
nand U19325 (N_19325,N_10092,N_13954);
nor U19326 (N_19326,N_11153,N_12877);
nor U19327 (N_19327,N_13921,N_12777);
and U19328 (N_19328,N_10216,N_11946);
xnor U19329 (N_19329,N_12004,N_11266);
nor U19330 (N_19330,N_11797,N_13345);
nor U19331 (N_19331,N_14977,N_11874);
xor U19332 (N_19332,N_11041,N_12875);
nor U19333 (N_19333,N_11875,N_14109);
nor U19334 (N_19334,N_12955,N_13819);
xnor U19335 (N_19335,N_12323,N_11301);
nor U19336 (N_19336,N_13931,N_13819);
and U19337 (N_19337,N_12419,N_10692);
nor U19338 (N_19338,N_10137,N_11440);
and U19339 (N_19339,N_11986,N_10112);
nor U19340 (N_19340,N_10917,N_14964);
and U19341 (N_19341,N_12751,N_13227);
and U19342 (N_19342,N_13810,N_11062);
nor U19343 (N_19343,N_14241,N_14117);
nor U19344 (N_19344,N_10238,N_10914);
and U19345 (N_19345,N_11409,N_11545);
xor U19346 (N_19346,N_14742,N_13278);
nor U19347 (N_19347,N_10697,N_11311);
and U19348 (N_19348,N_13702,N_10674);
nand U19349 (N_19349,N_13438,N_13737);
or U19350 (N_19350,N_11841,N_14866);
xnor U19351 (N_19351,N_12268,N_14078);
or U19352 (N_19352,N_10394,N_12790);
xor U19353 (N_19353,N_11770,N_10524);
nor U19354 (N_19354,N_11820,N_12914);
nand U19355 (N_19355,N_14582,N_14150);
and U19356 (N_19356,N_14587,N_12396);
nand U19357 (N_19357,N_10488,N_11292);
nor U19358 (N_19358,N_13075,N_14564);
and U19359 (N_19359,N_10538,N_14683);
or U19360 (N_19360,N_14645,N_12748);
and U19361 (N_19361,N_13756,N_10090);
nor U19362 (N_19362,N_10083,N_12414);
nand U19363 (N_19363,N_14642,N_10717);
nor U19364 (N_19364,N_10057,N_12108);
or U19365 (N_19365,N_10034,N_14673);
or U19366 (N_19366,N_10798,N_14023);
nor U19367 (N_19367,N_10651,N_11121);
and U19368 (N_19368,N_11994,N_11825);
and U19369 (N_19369,N_13325,N_13071);
xnor U19370 (N_19370,N_13035,N_13496);
xor U19371 (N_19371,N_13751,N_12680);
and U19372 (N_19372,N_14680,N_14306);
nand U19373 (N_19373,N_11487,N_11377);
nor U19374 (N_19374,N_11173,N_13814);
xnor U19375 (N_19375,N_10964,N_14917);
or U19376 (N_19376,N_12136,N_14262);
nand U19377 (N_19377,N_11547,N_11962);
xor U19378 (N_19378,N_12199,N_13185);
nor U19379 (N_19379,N_14238,N_13422);
and U19380 (N_19380,N_13865,N_12175);
and U19381 (N_19381,N_11202,N_10948);
and U19382 (N_19382,N_14717,N_13855);
nor U19383 (N_19383,N_12437,N_14518);
nor U19384 (N_19384,N_11343,N_12901);
or U19385 (N_19385,N_10177,N_12807);
or U19386 (N_19386,N_11808,N_14003);
or U19387 (N_19387,N_12216,N_11311);
nand U19388 (N_19388,N_10185,N_10336);
and U19389 (N_19389,N_10920,N_14350);
xnor U19390 (N_19390,N_10471,N_14538);
nor U19391 (N_19391,N_12463,N_13909);
nand U19392 (N_19392,N_12586,N_11612);
nor U19393 (N_19393,N_11735,N_13128);
or U19394 (N_19394,N_14106,N_11618);
or U19395 (N_19395,N_10892,N_13351);
nor U19396 (N_19396,N_13626,N_11368);
nand U19397 (N_19397,N_13346,N_10369);
and U19398 (N_19398,N_13121,N_14218);
xnor U19399 (N_19399,N_10402,N_12868);
nor U19400 (N_19400,N_10651,N_14324);
nor U19401 (N_19401,N_13760,N_11403);
nand U19402 (N_19402,N_12573,N_14050);
or U19403 (N_19403,N_11583,N_14361);
nor U19404 (N_19404,N_11165,N_14852);
or U19405 (N_19405,N_10987,N_11914);
or U19406 (N_19406,N_12593,N_13952);
xnor U19407 (N_19407,N_12909,N_12005);
nor U19408 (N_19408,N_13929,N_12454);
nand U19409 (N_19409,N_11634,N_14902);
and U19410 (N_19410,N_13142,N_11585);
and U19411 (N_19411,N_12053,N_10319);
nor U19412 (N_19412,N_10745,N_11599);
nand U19413 (N_19413,N_10932,N_12481);
and U19414 (N_19414,N_11710,N_11341);
nor U19415 (N_19415,N_14486,N_13592);
nor U19416 (N_19416,N_13920,N_14979);
or U19417 (N_19417,N_11283,N_11156);
nand U19418 (N_19418,N_11735,N_14424);
nor U19419 (N_19419,N_11542,N_12252);
or U19420 (N_19420,N_11565,N_11507);
or U19421 (N_19421,N_11284,N_14804);
xnor U19422 (N_19422,N_10293,N_12953);
or U19423 (N_19423,N_10813,N_12622);
and U19424 (N_19424,N_14315,N_14262);
and U19425 (N_19425,N_12639,N_14794);
nor U19426 (N_19426,N_12551,N_10366);
nor U19427 (N_19427,N_10476,N_12808);
xor U19428 (N_19428,N_11106,N_11697);
nor U19429 (N_19429,N_11177,N_10808);
or U19430 (N_19430,N_10892,N_14338);
or U19431 (N_19431,N_12719,N_11491);
nor U19432 (N_19432,N_11594,N_10531);
xnor U19433 (N_19433,N_12224,N_14423);
xor U19434 (N_19434,N_13603,N_14769);
xor U19435 (N_19435,N_14316,N_11803);
or U19436 (N_19436,N_14752,N_14233);
xor U19437 (N_19437,N_13501,N_14289);
and U19438 (N_19438,N_13267,N_11648);
nand U19439 (N_19439,N_13600,N_12282);
or U19440 (N_19440,N_11657,N_13964);
or U19441 (N_19441,N_11183,N_13155);
nand U19442 (N_19442,N_13353,N_12759);
or U19443 (N_19443,N_14264,N_14682);
nand U19444 (N_19444,N_13846,N_13782);
and U19445 (N_19445,N_12674,N_11931);
or U19446 (N_19446,N_11873,N_10174);
xor U19447 (N_19447,N_11039,N_10506);
nand U19448 (N_19448,N_14966,N_10683);
xnor U19449 (N_19449,N_11232,N_12306);
xnor U19450 (N_19450,N_11502,N_10709);
xnor U19451 (N_19451,N_12335,N_10112);
and U19452 (N_19452,N_14878,N_12307);
xnor U19453 (N_19453,N_12766,N_12555);
and U19454 (N_19454,N_11124,N_11635);
or U19455 (N_19455,N_14045,N_11800);
xnor U19456 (N_19456,N_11491,N_13843);
and U19457 (N_19457,N_13582,N_13527);
nand U19458 (N_19458,N_12226,N_11969);
xor U19459 (N_19459,N_11790,N_14205);
nor U19460 (N_19460,N_10489,N_12946);
nor U19461 (N_19461,N_14642,N_11666);
xnor U19462 (N_19462,N_14507,N_13072);
or U19463 (N_19463,N_12878,N_13061);
and U19464 (N_19464,N_13586,N_11984);
xor U19465 (N_19465,N_13948,N_12705);
and U19466 (N_19466,N_10979,N_11569);
and U19467 (N_19467,N_13352,N_10538);
nand U19468 (N_19468,N_10420,N_12600);
xor U19469 (N_19469,N_14258,N_12855);
or U19470 (N_19470,N_11031,N_11826);
nand U19471 (N_19471,N_14411,N_10451);
xnor U19472 (N_19472,N_10992,N_10368);
and U19473 (N_19473,N_13290,N_11552);
nand U19474 (N_19474,N_11552,N_13821);
xnor U19475 (N_19475,N_11577,N_13483);
or U19476 (N_19476,N_14223,N_10996);
or U19477 (N_19477,N_12403,N_13084);
xnor U19478 (N_19478,N_14307,N_13172);
and U19479 (N_19479,N_13688,N_13345);
and U19480 (N_19480,N_14571,N_13142);
xor U19481 (N_19481,N_12467,N_14521);
xnor U19482 (N_19482,N_11107,N_10042);
nor U19483 (N_19483,N_11009,N_10410);
xor U19484 (N_19484,N_14385,N_10664);
nor U19485 (N_19485,N_14248,N_12159);
or U19486 (N_19486,N_11528,N_10597);
nand U19487 (N_19487,N_14356,N_13925);
nor U19488 (N_19488,N_10673,N_11107);
xnor U19489 (N_19489,N_10623,N_11331);
nand U19490 (N_19490,N_14012,N_14416);
xnor U19491 (N_19491,N_14895,N_14869);
nand U19492 (N_19492,N_13788,N_11566);
nor U19493 (N_19493,N_13378,N_11191);
nand U19494 (N_19494,N_12816,N_11808);
nand U19495 (N_19495,N_10886,N_13632);
and U19496 (N_19496,N_10574,N_12496);
or U19497 (N_19497,N_14493,N_11942);
and U19498 (N_19498,N_10240,N_10818);
nand U19499 (N_19499,N_11390,N_11717);
or U19500 (N_19500,N_14667,N_13611);
xor U19501 (N_19501,N_11325,N_12315);
nor U19502 (N_19502,N_14682,N_12529);
and U19503 (N_19503,N_12265,N_11616);
nand U19504 (N_19504,N_12814,N_10559);
and U19505 (N_19505,N_12745,N_12873);
nor U19506 (N_19506,N_12079,N_14013);
nand U19507 (N_19507,N_12650,N_12245);
xor U19508 (N_19508,N_10860,N_14979);
nand U19509 (N_19509,N_11553,N_11994);
nor U19510 (N_19510,N_13931,N_11457);
and U19511 (N_19511,N_12585,N_12103);
xnor U19512 (N_19512,N_10450,N_12095);
xor U19513 (N_19513,N_10806,N_12601);
nand U19514 (N_19514,N_12129,N_13376);
or U19515 (N_19515,N_12904,N_13532);
xnor U19516 (N_19516,N_13468,N_14861);
nor U19517 (N_19517,N_11786,N_12039);
or U19518 (N_19518,N_14395,N_13687);
and U19519 (N_19519,N_13286,N_14477);
xor U19520 (N_19520,N_13901,N_13108);
nor U19521 (N_19521,N_14805,N_14637);
nor U19522 (N_19522,N_10863,N_11071);
and U19523 (N_19523,N_12069,N_12406);
or U19524 (N_19524,N_11695,N_13160);
xnor U19525 (N_19525,N_10731,N_11782);
nor U19526 (N_19526,N_12176,N_14801);
nand U19527 (N_19527,N_14835,N_12128);
and U19528 (N_19528,N_14558,N_10589);
or U19529 (N_19529,N_14477,N_14796);
nor U19530 (N_19530,N_12740,N_14513);
or U19531 (N_19531,N_12051,N_12382);
nor U19532 (N_19532,N_11934,N_12484);
or U19533 (N_19533,N_10865,N_11023);
and U19534 (N_19534,N_12863,N_12354);
xor U19535 (N_19535,N_12809,N_11679);
nor U19536 (N_19536,N_12853,N_13129);
xor U19537 (N_19537,N_12062,N_12867);
nor U19538 (N_19538,N_12691,N_13760);
and U19539 (N_19539,N_10073,N_10311);
xnor U19540 (N_19540,N_13801,N_11675);
and U19541 (N_19541,N_10502,N_10547);
xor U19542 (N_19542,N_10267,N_13978);
nand U19543 (N_19543,N_12061,N_12965);
and U19544 (N_19544,N_14307,N_11859);
nor U19545 (N_19545,N_11252,N_14051);
or U19546 (N_19546,N_14091,N_13027);
or U19547 (N_19547,N_13574,N_11470);
or U19548 (N_19548,N_10844,N_14355);
xnor U19549 (N_19549,N_10956,N_11441);
nand U19550 (N_19550,N_10560,N_13549);
xnor U19551 (N_19551,N_14739,N_14275);
and U19552 (N_19552,N_13696,N_13204);
and U19553 (N_19553,N_10284,N_12429);
nor U19554 (N_19554,N_11336,N_13177);
or U19555 (N_19555,N_10259,N_13049);
or U19556 (N_19556,N_10693,N_13529);
xor U19557 (N_19557,N_10151,N_11428);
xor U19558 (N_19558,N_14735,N_11981);
or U19559 (N_19559,N_10065,N_12903);
or U19560 (N_19560,N_14935,N_13015);
nand U19561 (N_19561,N_11946,N_12179);
and U19562 (N_19562,N_11913,N_14357);
nor U19563 (N_19563,N_12460,N_12186);
or U19564 (N_19564,N_11175,N_10156);
and U19565 (N_19565,N_13982,N_14835);
nand U19566 (N_19566,N_13287,N_10411);
xnor U19567 (N_19567,N_10947,N_14834);
or U19568 (N_19568,N_10411,N_10514);
nor U19569 (N_19569,N_11661,N_12849);
xor U19570 (N_19570,N_12167,N_10554);
nand U19571 (N_19571,N_14587,N_14970);
and U19572 (N_19572,N_10734,N_14895);
xor U19573 (N_19573,N_12627,N_10027);
or U19574 (N_19574,N_10057,N_13189);
nand U19575 (N_19575,N_12321,N_10105);
nor U19576 (N_19576,N_12652,N_11019);
nand U19577 (N_19577,N_10143,N_10182);
and U19578 (N_19578,N_14635,N_14584);
and U19579 (N_19579,N_12537,N_13710);
and U19580 (N_19580,N_12233,N_14657);
nand U19581 (N_19581,N_12019,N_13084);
nor U19582 (N_19582,N_10047,N_12504);
or U19583 (N_19583,N_10055,N_10545);
nor U19584 (N_19584,N_13934,N_13735);
and U19585 (N_19585,N_11845,N_10603);
nor U19586 (N_19586,N_10377,N_11384);
nand U19587 (N_19587,N_13388,N_13525);
nor U19588 (N_19588,N_13363,N_14976);
and U19589 (N_19589,N_13838,N_10303);
nand U19590 (N_19590,N_11908,N_11631);
xor U19591 (N_19591,N_13988,N_14283);
or U19592 (N_19592,N_13126,N_13840);
or U19593 (N_19593,N_10724,N_11415);
or U19594 (N_19594,N_14533,N_12771);
xor U19595 (N_19595,N_12103,N_13644);
nor U19596 (N_19596,N_14445,N_12195);
xor U19597 (N_19597,N_12475,N_12499);
or U19598 (N_19598,N_11315,N_10676);
nor U19599 (N_19599,N_14642,N_11400);
xor U19600 (N_19600,N_14429,N_13135);
nand U19601 (N_19601,N_11834,N_14894);
nand U19602 (N_19602,N_11513,N_11553);
nor U19603 (N_19603,N_13249,N_11973);
nor U19604 (N_19604,N_14250,N_12811);
and U19605 (N_19605,N_10910,N_14048);
nor U19606 (N_19606,N_11927,N_14818);
nor U19607 (N_19607,N_12205,N_12793);
xnor U19608 (N_19608,N_11512,N_12214);
nor U19609 (N_19609,N_13912,N_13173);
nand U19610 (N_19610,N_11049,N_13350);
xor U19611 (N_19611,N_12889,N_14841);
nor U19612 (N_19612,N_10046,N_10925);
xnor U19613 (N_19613,N_10413,N_11901);
and U19614 (N_19614,N_14946,N_10739);
nand U19615 (N_19615,N_11692,N_13748);
nand U19616 (N_19616,N_14127,N_13371);
xor U19617 (N_19617,N_11461,N_13396);
or U19618 (N_19618,N_13502,N_10904);
xnor U19619 (N_19619,N_10084,N_14020);
nand U19620 (N_19620,N_14230,N_10469);
nor U19621 (N_19621,N_13822,N_13238);
xor U19622 (N_19622,N_14317,N_13820);
nand U19623 (N_19623,N_10993,N_10344);
nor U19624 (N_19624,N_12764,N_12315);
or U19625 (N_19625,N_14410,N_10970);
and U19626 (N_19626,N_10823,N_11005);
or U19627 (N_19627,N_14788,N_11799);
nand U19628 (N_19628,N_13392,N_11740);
nand U19629 (N_19629,N_12275,N_11680);
xor U19630 (N_19630,N_14453,N_10630);
and U19631 (N_19631,N_11402,N_13825);
or U19632 (N_19632,N_12541,N_11558);
nand U19633 (N_19633,N_14338,N_11415);
nand U19634 (N_19634,N_11532,N_12894);
nand U19635 (N_19635,N_14994,N_10914);
nor U19636 (N_19636,N_13387,N_12594);
xnor U19637 (N_19637,N_12242,N_14228);
xnor U19638 (N_19638,N_11777,N_13288);
nand U19639 (N_19639,N_12692,N_14192);
nand U19640 (N_19640,N_13029,N_13670);
nand U19641 (N_19641,N_13043,N_13197);
xor U19642 (N_19642,N_14997,N_13835);
and U19643 (N_19643,N_11108,N_13784);
and U19644 (N_19644,N_13757,N_14928);
or U19645 (N_19645,N_12273,N_11949);
and U19646 (N_19646,N_11219,N_12887);
or U19647 (N_19647,N_12225,N_14602);
xor U19648 (N_19648,N_11582,N_12233);
and U19649 (N_19649,N_11768,N_13018);
or U19650 (N_19650,N_13314,N_12577);
nand U19651 (N_19651,N_10155,N_11264);
nor U19652 (N_19652,N_12686,N_12178);
nor U19653 (N_19653,N_11666,N_11943);
nor U19654 (N_19654,N_13108,N_11946);
xnor U19655 (N_19655,N_12166,N_11795);
nand U19656 (N_19656,N_11114,N_12509);
nor U19657 (N_19657,N_14344,N_10641);
nand U19658 (N_19658,N_11884,N_10263);
or U19659 (N_19659,N_11963,N_12257);
nor U19660 (N_19660,N_13969,N_13668);
and U19661 (N_19661,N_14782,N_10459);
xor U19662 (N_19662,N_14857,N_13212);
nand U19663 (N_19663,N_11223,N_12539);
nand U19664 (N_19664,N_10781,N_13044);
nand U19665 (N_19665,N_13702,N_13979);
or U19666 (N_19666,N_13189,N_11280);
nor U19667 (N_19667,N_13352,N_10215);
or U19668 (N_19668,N_13673,N_11688);
nor U19669 (N_19669,N_10747,N_14101);
xnor U19670 (N_19670,N_10085,N_11872);
xnor U19671 (N_19671,N_11236,N_12691);
nor U19672 (N_19672,N_12952,N_10928);
xor U19673 (N_19673,N_14126,N_14860);
nor U19674 (N_19674,N_13387,N_12122);
and U19675 (N_19675,N_13136,N_11830);
nand U19676 (N_19676,N_14724,N_10467);
or U19677 (N_19677,N_11446,N_11215);
and U19678 (N_19678,N_13516,N_10978);
and U19679 (N_19679,N_14494,N_13132);
nand U19680 (N_19680,N_11783,N_10339);
nand U19681 (N_19681,N_11123,N_13315);
xnor U19682 (N_19682,N_10024,N_12084);
nand U19683 (N_19683,N_14344,N_14006);
nor U19684 (N_19684,N_14234,N_14024);
or U19685 (N_19685,N_12338,N_11686);
nor U19686 (N_19686,N_13950,N_10436);
nor U19687 (N_19687,N_11558,N_12098);
xor U19688 (N_19688,N_13670,N_14819);
nor U19689 (N_19689,N_10992,N_12559);
xor U19690 (N_19690,N_13228,N_11586);
or U19691 (N_19691,N_14796,N_12973);
nor U19692 (N_19692,N_11454,N_11734);
xnor U19693 (N_19693,N_13213,N_11716);
nor U19694 (N_19694,N_10594,N_10024);
nand U19695 (N_19695,N_14056,N_13708);
nor U19696 (N_19696,N_10989,N_10006);
nand U19697 (N_19697,N_10870,N_10665);
xor U19698 (N_19698,N_14507,N_10615);
or U19699 (N_19699,N_10949,N_10487);
and U19700 (N_19700,N_13651,N_13111);
nand U19701 (N_19701,N_14168,N_10931);
nor U19702 (N_19702,N_11197,N_10632);
nand U19703 (N_19703,N_11739,N_13973);
nand U19704 (N_19704,N_10134,N_14434);
and U19705 (N_19705,N_13435,N_10545);
nand U19706 (N_19706,N_10488,N_12742);
nand U19707 (N_19707,N_12121,N_10744);
or U19708 (N_19708,N_12767,N_12991);
or U19709 (N_19709,N_12726,N_13343);
or U19710 (N_19710,N_13060,N_12203);
and U19711 (N_19711,N_12509,N_12728);
nor U19712 (N_19712,N_14163,N_14247);
and U19713 (N_19713,N_11115,N_14493);
nand U19714 (N_19714,N_13882,N_11914);
xor U19715 (N_19715,N_13643,N_13953);
nor U19716 (N_19716,N_13566,N_10647);
and U19717 (N_19717,N_14848,N_13457);
nor U19718 (N_19718,N_10844,N_11269);
and U19719 (N_19719,N_10931,N_13574);
nor U19720 (N_19720,N_13023,N_13298);
or U19721 (N_19721,N_10724,N_12973);
xnor U19722 (N_19722,N_11612,N_11154);
xor U19723 (N_19723,N_10798,N_13710);
and U19724 (N_19724,N_14447,N_12387);
or U19725 (N_19725,N_10360,N_12636);
and U19726 (N_19726,N_11537,N_11510);
xor U19727 (N_19727,N_12505,N_14462);
or U19728 (N_19728,N_13848,N_10618);
nor U19729 (N_19729,N_10326,N_13887);
xor U19730 (N_19730,N_13774,N_13754);
nand U19731 (N_19731,N_10309,N_13156);
or U19732 (N_19732,N_14042,N_13788);
and U19733 (N_19733,N_13229,N_13672);
xnor U19734 (N_19734,N_12994,N_13536);
or U19735 (N_19735,N_12121,N_11485);
nor U19736 (N_19736,N_10396,N_13771);
nor U19737 (N_19737,N_11632,N_14065);
nor U19738 (N_19738,N_13692,N_11461);
nor U19739 (N_19739,N_12108,N_11974);
and U19740 (N_19740,N_14027,N_11892);
nor U19741 (N_19741,N_12934,N_14288);
nand U19742 (N_19742,N_10659,N_11051);
or U19743 (N_19743,N_11182,N_14894);
or U19744 (N_19744,N_13320,N_10737);
nand U19745 (N_19745,N_13775,N_12469);
nand U19746 (N_19746,N_14980,N_11578);
nand U19747 (N_19747,N_10317,N_13323);
xnor U19748 (N_19748,N_10739,N_11802);
and U19749 (N_19749,N_13149,N_12638);
nor U19750 (N_19750,N_12688,N_12180);
or U19751 (N_19751,N_13744,N_11681);
nor U19752 (N_19752,N_12467,N_11147);
xnor U19753 (N_19753,N_11955,N_13474);
and U19754 (N_19754,N_11576,N_13238);
and U19755 (N_19755,N_10295,N_14427);
xnor U19756 (N_19756,N_10635,N_11688);
nor U19757 (N_19757,N_14948,N_14231);
and U19758 (N_19758,N_13412,N_12269);
or U19759 (N_19759,N_12631,N_12356);
or U19760 (N_19760,N_11535,N_14844);
xnor U19761 (N_19761,N_12713,N_14813);
and U19762 (N_19762,N_12658,N_11290);
or U19763 (N_19763,N_13837,N_10083);
or U19764 (N_19764,N_13860,N_14266);
and U19765 (N_19765,N_14622,N_12452);
or U19766 (N_19766,N_10475,N_12532);
xnor U19767 (N_19767,N_13099,N_13813);
nor U19768 (N_19768,N_11664,N_12177);
nand U19769 (N_19769,N_14143,N_11610);
and U19770 (N_19770,N_10535,N_13401);
xor U19771 (N_19771,N_12610,N_14964);
nand U19772 (N_19772,N_11659,N_10039);
or U19773 (N_19773,N_10041,N_10979);
nor U19774 (N_19774,N_11058,N_11309);
xor U19775 (N_19775,N_12960,N_12157);
or U19776 (N_19776,N_12789,N_10659);
xnor U19777 (N_19777,N_10063,N_10549);
and U19778 (N_19778,N_11824,N_14822);
nand U19779 (N_19779,N_11130,N_14899);
and U19780 (N_19780,N_11576,N_14624);
or U19781 (N_19781,N_11772,N_14200);
nand U19782 (N_19782,N_13860,N_13020);
or U19783 (N_19783,N_14553,N_13142);
and U19784 (N_19784,N_10600,N_11594);
or U19785 (N_19785,N_11789,N_14514);
or U19786 (N_19786,N_11030,N_11689);
nor U19787 (N_19787,N_11477,N_12722);
or U19788 (N_19788,N_12528,N_10680);
nor U19789 (N_19789,N_10382,N_11695);
xor U19790 (N_19790,N_11681,N_10540);
nand U19791 (N_19791,N_13451,N_14363);
nor U19792 (N_19792,N_10434,N_14926);
nand U19793 (N_19793,N_11666,N_12556);
and U19794 (N_19794,N_12309,N_12909);
nor U19795 (N_19795,N_11201,N_14345);
and U19796 (N_19796,N_11880,N_12555);
nor U19797 (N_19797,N_13958,N_13792);
nand U19798 (N_19798,N_11554,N_12638);
nor U19799 (N_19799,N_11551,N_13610);
nand U19800 (N_19800,N_10096,N_14567);
or U19801 (N_19801,N_14517,N_11090);
nor U19802 (N_19802,N_11283,N_13157);
xor U19803 (N_19803,N_10992,N_13098);
and U19804 (N_19804,N_10680,N_12503);
xnor U19805 (N_19805,N_14685,N_12556);
xnor U19806 (N_19806,N_10167,N_13387);
or U19807 (N_19807,N_14152,N_11605);
or U19808 (N_19808,N_11424,N_14992);
nand U19809 (N_19809,N_13130,N_13977);
nor U19810 (N_19810,N_14712,N_13148);
and U19811 (N_19811,N_10964,N_10205);
nand U19812 (N_19812,N_13129,N_12556);
nor U19813 (N_19813,N_12783,N_10467);
nor U19814 (N_19814,N_12773,N_13384);
nor U19815 (N_19815,N_14383,N_10286);
and U19816 (N_19816,N_11594,N_13638);
and U19817 (N_19817,N_13215,N_11635);
and U19818 (N_19818,N_12419,N_10218);
nand U19819 (N_19819,N_10738,N_11243);
or U19820 (N_19820,N_12203,N_12012);
or U19821 (N_19821,N_11752,N_10936);
nor U19822 (N_19822,N_13243,N_10562);
nand U19823 (N_19823,N_12227,N_11233);
nor U19824 (N_19824,N_10636,N_14863);
and U19825 (N_19825,N_14998,N_13909);
or U19826 (N_19826,N_10648,N_10071);
nand U19827 (N_19827,N_13039,N_11486);
and U19828 (N_19828,N_13659,N_14662);
and U19829 (N_19829,N_12937,N_12412);
xnor U19830 (N_19830,N_14183,N_12293);
and U19831 (N_19831,N_12977,N_13611);
nor U19832 (N_19832,N_13610,N_14641);
nand U19833 (N_19833,N_13872,N_11845);
nand U19834 (N_19834,N_11957,N_14156);
nor U19835 (N_19835,N_12154,N_12105);
and U19836 (N_19836,N_13890,N_13026);
and U19837 (N_19837,N_14398,N_13632);
or U19838 (N_19838,N_11945,N_12479);
nand U19839 (N_19839,N_14310,N_14814);
or U19840 (N_19840,N_12780,N_14646);
nand U19841 (N_19841,N_13438,N_11031);
and U19842 (N_19842,N_10672,N_11399);
and U19843 (N_19843,N_14779,N_13906);
or U19844 (N_19844,N_10853,N_11338);
and U19845 (N_19845,N_12873,N_10777);
nor U19846 (N_19846,N_13850,N_10595);
and U19847 (N_19847,N_14886,N_13944);
or U19848 (N_19848,N_14502,N_11399);
nand U19849 (N_19849,N_10574,N_11350);
or U19850 (N_19850,N_10303,N_13335);
and U19851 (N_19851,N_12762,N_13722);
nor U19852 (N_19852,N_10934,N_10123);
nand U19853 (N_19853,N_13487,N_13923);
xor U19854 (N_19854,N_12792,N_12128);
nor U19855 (N_19855,N_11991,N_12789);
xor U19856 (N_19856,N_13446,N_10476);
nand U19857 (N_19857,N_13322,N_12579);
nor U19858 (N_19858,N_14790,N_11035);
and U19859 (N_19859,N_11509,N_12379);
xnor U19860 (N_19860,N_10962,N_11134);
or U19861 (N_19861,N_10532,N_11932);
and U19862 (N_19862,N_12438,N_12907);
and U19863 (N_19863,N_10832,N_11765);
nor U19864 (N_19864,N_12690,N_11178);
nand U19865 (N_19865,N_10138,N_12614);
xor U19866 (N_19866,N_12102,N_10328);
nor U19867 (N_19867,N_10420,N_11225);
nor U19868 (N_19868,N_13875,N_10147);
or U19869 (N_19869,N_12958,N_10016);
nor U19870 (N_19870,N_10178,N_12383);
or U19871 (N_19871,N_10452,N_12555);
and U19872 (N_19872,N_13451,N_10413);
nor U19873 (N_19873,N_12310,N_14309);
and U19874 (N_19874,N_14752,N_11898);
nand U19875 (N_19875,N_10434,N_13535);
or U19876 (N_19876,N_13591,N_13634);
or U19877 (N_19877,N_12536,N_13824);
nor U19878 (N_19878,N_14545,N_14159);
and U19879 (N_19879,N_14360,N_12990);
and U19880 (N_19880,N_12421,N_13065);
or U19881 (N_19881,N_14459,N_13414);
and U19882 (N_19882,N_12940,N_12460);
nor U19883 (N_19883,N_11170,N_12253);
or U19884 (N_19884,N_10265,N_10159);
nor U19885 (N_19885,N_12764,N_11278);
or U19886 (N_19886,N_11243,N_11791);
and U19887 (N_19887,N_12198,N_11919);
and U19888 (N_19888,N_10963,N_13968);
nor U19889 (N_19889,N_11918,N_11051);
and U19890 (N_19890,N_11821,N_11678);
or U19891 (N_19891,N_14921,N_10326);
or U19892 (N_19892,N_12709,N_14946);
and U19893 (N_19893,N_10361,N_13301);
and U19894 (N_19894,N_10594,N_10206);
nand U19895 (N_19895,N_13788,N_10824);
or U19896 (N_19896,N_11935,N_14689);
xor U19897 (N_19897,N_11390,N_13405);
nand U19898 (N_19898,N_12960,N_11600);
xnor U19899 (N_19899,N_12164,N_13042);
xor U19900 (N_19900,N_13394,N_12311);
or U19901 (N_19901,N_12912,N_12563);
nor U19902 (N_19902,N_11657,N_11255);
nand U19903 (N_19903,N_10834,N_14970);
xnor U19904 (N_19904,N_13947,N_14766);
nand U19905 (N_19905,N_14211,N_14537);
nor U19906 (N_19906,N_12898,N_12473);
xor U19907 (N_19907,N_10833,N_10977);
and U19908 (N_19908,N_12150,N_13477);
nor U19909 (N_19909,N_10873,N_12712);
and U19910 (N_19910,N_12574,N_10898);
or U19911 (N_19911,N_10264,N_13445);
or U19912 (N_19912,N_12793,N_11823);
nand U19913 (N_19913,N_12893,N_12585);
or U19914 (N_19914,N_12586,N_13335);
and U19915 (N_19915,N_12698,N_11691);
nor U19916 (N_19916,N_12599,N_14726);
nor U19917 (N_19917,N_13340,N_11833);
and U19918 (N_19918,N_13934,N_13793);
nand U19919 (N_19919,N_13967,N_12158);
xnor U19920 (N_19920,N_13186,N_12988);
nor U19921 (N_19921,N_10406,N_10442);
and U19922 (N_19922,N_14001,N_10512);
xnor U19923 (N_19923,N_10743,N_13861);
nor U19924 (N_19924,N_12774,N_10585);
xnor U19925 (N_19925,N_13265,N_10532);
nor U19926 (N_19926,N_11300,N_10463);
nor U19927 (N_19927,N_12532,N_14370);
nor U19928 (N_19928,N_10531,N_13562);
nand U19929 (N_19929,N_13564,N_10030);
nand U19930 (N_19930,N_14995,N_14138);
and U19931 (N_19931,N_10518,N_14249);
and U19932 (N_19932,N_14605,N_13019);
nor U19933 (N_19933,N_14068,N_11944);
nand U19934 (N_19934,N_13646,N_10213);
xnor U19935 (N_19935,N_10080,N_12180);
nand U19936 (N_19936,N_10563,N_12081);
nand U19937 (N_19937,N_10127,N_14812);
nand U19938 (N_19938,N_10283,N_12462);
nand U19939 (N_19939,N_10997,N_10187);
xor U19940 (N_19940,N_10718,N_12366);
or U19941 (N_19941,N_10181,N_10094);
nor U19942 (N_19942,N_10496,N_10093);
nand U19943 (N_19943,N_11352,N_12736);
and U19944 (N_19944,N_12390,N_13224);
or U19945 (N_19945,N_13219,N_14132);
or U19946 (N_19946,N_14853,N_13814);
nor U19947 (N_19947,N_13253,N_14354);
and U19948 (N_19948,N_14101,N_13127);
nor U19949 (N_19949,N_10512,N_11253);
and U19950 (N_19950,N_12795,N_11713);
and U19951 (N_19951,N_12700,N_10978);
nand U19952 (N_19952,N_12550,N_10603);
and U19953 (N_19953,N_13128,N_14975);
xor U19954 (N_19954,N_14223,N_12606);
xor U19955 (N_19955,N_12980,N_13431);
or U19956 (N_19956,N_14675,N_14517);
or U19957 (N_19957,N_13393,N_11935);
nor U19958 (N_19958,N_11083,N_13203);
or U19959 (N_19959,N_13254,N_12675);
and U19960 (N_19960,N_10459,N_12888);
xor U19961 (N_19961,N_14335,N_14167);
nand U19962 (N_19962,N_13739,N_14488);
nand U19963 (N_19963,N_12582,N_12183);
nor U19964 (N_19964,N_11673,N_13869);
nor U19965 (N_19965,N_13684,N_13483);
and U19966 (N_19966,N_12291,N_14448);
nand U19967 (N_19967,N_14592,N_13432);
or U19968 (N_19968,N_10091,N_14620);
or U19969 (N_19969,N_11556,N_13467);
nand U19970 (N_19970,N_10520,N_11559);
xor U19971 (N_19971,N_11372,N_11204);
xor U19972 (N_19972,N_13676,N_12791);
nand U19973 (N_19973,N_12351,N_14764);
nand U19974 (N_19974,N_11697,N_12239);
or U19975 (N_19975,N_13106,N_11109);
nor U19976 (N_19976,N_14084,N_14154);
or U19977 (N_19977,N_11994,N_10506);
nand U19978 (N_19978,N_14407,N_11304);
xnor U19979 (N_19979,N_13309,N_10577);
xnor U19980 (N_19980,N_11911,N_14460);
nor U19981 (N_19981,N_14950,N_14981);
or U19982 (N_19982,N_13632,N_11969);
and U19983 (N_19983,N_10260,N_12297);
nand U19984 (N_19984,N_11929,N_11114);
and U19985 (N_19985,N_10905,N_11793);
nand U19986 (N_19986,N_11405,N_12771);
or U19987 (N_19987,N_14326,N_10766);
nand U19988 (N_19988,N_11771,N_14956);
or U19989 (N_19989,N_12855,N_12074);
nor U19990 (N_19990,N_13948,N_14635);
xnor U19991 (N_19991,N_13573,N_14361);
xnor U19992 (N_19992,N_14620,N_12409);
xnor U19993 (N_19993,N_12925,N_10832);
and U19994 (N_19994,N_11928,N_10747);
nor U19995 (N_19995,N_14632,N_11869);
xnor U19996 (N_19996,N_14437,N_13729);
or U19997 (N_19997,N_12415,N_12608);
or U19998 (N_19998,N_12667,N_14762);
nand U19999 (N_19999,N_13157,N_14387);
xnor U20000 (N_20000,N_16822,N_15190);
nand U20001 (N_20001,N_19272,N_15887);
nor U20002 (N_20002,N_15373,N_16746);
or U20003 (N_20003,N_17399,N_19777);
nand U20004 (N_20004,N_19736,N_17319);
nor U20005 (N_20005,N_15990,N_18759);
and U20006 (N_20006,N_19717,N_17520);
nand U20007 (N_20007,N_19543,N_15950);
nand U20008 (N_20008,N_19087,N_15678);
and U20009 (N_20009,N_15390,N_17643);
xor U20010 (N_20010,N_16071,N_16692);
or U20011 (N_20011,N_19515,N_15502);
or U20012 (N_20012,N_19806,N_18347);
and U20013 (N_20013,N_18994,N_19747);
nand U20014 (N_20014,N_19999,N_19456);
xor U20015 (N_20015,N_18081,N_17408);
xor U20016 (N_20016,N_17404,N_18802);
nor U20017 (N_20017,N_15668,N_17533);
nand U20018 (N_20018,N_17452,N_15590);
or U20019 (N_20019,N_19270,N_15568);
nor U20020 (N_20020,N_15429,N_17709);
xor U20021 (N_20021,N_19205,N_17612);
xnor U20022 (N_20022,N_17460,N_18602);
or U20023 (N_20023,N_19018,N_15387);
or U20024 (N_20024,N_18865,N_16848);
nand U20025 (N_20025,N_15236,N_17896);
nor U20026 (N_20026,N_15501,N_18575);
and U20027 (N_20027,N_18888,N_18911);
or U20028 (N_20028,N_16913,N_17106);
or U20029 (N_20029,N_18177,N_16806);
or U20030 (N_20030,N_16695,N_18954);
nand U20031 (N_20031,N_19923,N_16081);
and U20032 (N_20032,N_18705,N_17316);
or U20033 (N_20033,N_18357,N_17848);
or U20034 (N_20034,N_16982,N_19036);
nor U20035 (N_20035,N_17818,N_17051);
and U20036 (N_20036,N_15873,N_17807);
or U20037 (N_20037,N_17658,N_16386);
nor U20038 (N_20038,N_18023,N_18734);
xnor U20039 (N_20039,N_15483,N_15603);
or U20040 (N_20040,N_16669,N_19006);
nor U20041 (N_20041,N_17145,N_17207);
nand U20042 (N_20042,N_18387,N_19871);
nor U20043 (N_20043,N_18735,N_15948);
and U20044 (N_20044,N_18298,N_17115);
or U20045 (N_20045,N_17457,N_16618);
or U20046 (N_20046,N_15230,N_19130);
xor U20047 (N_20047,N_15855,N_16204);
and U20048 (N_20048,N_17366,N_17999);
nand U20049 (N_20049,N_18946,N_19697);
nor U20050 (N_20050,N_18979,N_19255);
xor U20051 (N_20051,N_15033,N_19132);
or U20052 (N_20052,N_17560,N_18579);
or U20053 (N_20053,N_19307,N_17799);
and U20054 (N_20054,N_15181,N_16581);
nand U20055 (N_20055,N_19296,N_15465);
nand U20056 (N_20056,N_18282,N_19724);
or U20057 (N_20057,N_15388,N_19888);
or U20058 (N_20058,N_18074,N_18538);
or U20059 (N_20059,N_17356,N_18601);
and U20060 (N_20060,N_16169,N_17912);
and U20061 (N_20061,N_19640,N_17859);
nor U20062 (N_20062,N_19176,N_17708);
and U20063 (N_20063,N_19941,N_15958);
and U20064 (N_20064,N_16475,N_17814);
xnor U20065 (N_20065,N_18267,N_16999);
or U20066 (N_20066,N_17063,N_16390);
and U20067 (N_20067,N_17285,N_15244);
and U20068 (N_20068,N_15679,N_16510);
nor U20069 (N_20069,N_19774,N_17043);
nand U20070 (N_20070,N_15667,N_18928);
and U20071 (N_20071,N_19044,N_17338);
and U20072 (N_20072,N_17586,N_18892);
nand U20073 (N_20073,N_18346,N_18804);
xnor U20074 (N_20074,N_19797,N_18006);
nand U20075 (N_20075,N_15787,N_19787);
or U20076 (N_20076,N_19580,N_15112);
nand U20077 (N_20077,N_16102,N_15402);
or U20078 (N_20078,N_16128,N_17378);
xnor U20079 (N_20079,N_16380,N_18855);
and U20080 (N_20080,N_16662,N_16236);
xnor U20081 (N_20081,N_17751,N_18783);
nor U20082 (N_20082,N_15509,N_18243);
and U20083 (N_20083,N_16644,N_18902);
xor U20084 (N_20084,N_17244,N_19361);
or U20085 (N_20085,N_15774,N_18240);
nand U20086 (N_20086,N_18525,N_18196);
or U20087 (N_20087,N_18609,N_16768);
nand U20088 (N_20088,N_19303,N_17716);
nor U20089 (N_20089,N_16868,N_17987);
or U20090 (N_20090,N_19162,N_16246);
xnor U20091 (N_20091,N_19293,N_16221);
xnor U20092 (N_20092,N_17868,N_18161);
and U20093 (N_20093,N_17477,N_17744);
and U20094 (N_20094,N_15286,N_19064);
xnor U20095 (N_20095,N_18148,N_19744);
nor U20096 (N_20096,N_18051,N_17531);
nand U20097 (N_20097,N_17522,N_18955);
nand U20098 (N_20098,N_16203,N_15857);
xnor U20099 (N_20099,N_15179,N_19665);
nor U20100 (N_20100,N_18683,N_19514);
nor U20101 (N_20101,N_17937,N_16804);
nand U20102 (N_20102,N_19156,N_18369);
nand U20103 (N_20103,N_15938,N_16328);
and U20104 (N_20104,N_16192,N_16084);
nor U20105 (N_20105,N_19037,N_17895);
nor U20106 (N_20106,N_18645,N_19125);
xor U20107 (N_20107,N_16834,N_15091);
xnor U20108 (N_20108,N_15757,N_19577);
nand U20109 (N_20109,N_16055,N_17939);
nand U20110 (N_20110,N_16991,N_18682);
nand U20111 (N_20111,N_15370,N_15520);
and U20112 (N_20112,N_15722,N_17314);
nor U20113 (N_20113,N_17032,N_15783);
or U20114 (N_20114,N_17927,N_17405);
or U20115 (N_20115,N_15718,N_15413);
nand U20116 (N_20116,N_16816,N_15002);
or U20117 (N_20117,N_17669,N_15551);
nor U20118 (N_20118,N_15635,N_15926);
or U20119 (N_20119,N_15115,N_17216);
nand U20120 (N_20120,N_15310,N_19373);
nand U20121 (N_20121,N_16395,N_16326);
nor U20122 (N_20122,N_18944,N_17031);
nand U20123 (N_20123,N_18329,N_15619);
nand U20124 (N_20124,N_16653,N_18750);
and U20125 (N_20125,N_18001,N_18215);
or U20126 (N_20126,N_19557,N_19025);
or U20127 (N_20127,N_16279,N_19939);
xor U20128 (N_20128,N_15694,N_18030);
nand U20129 (N_20129,N_19406,N_15817);
nor U20130 (N_20130,N_15297,N_18303);
xnor U20131 (N_20131,N_19096,N_17144);
nand U20132 (N_20132,N_18122,N_16638);
nand U20133 (N_20133,N_15562,N_15629);
xnor U20134 (N_20134,N_17002,N_17220);
and U20135 (N_20135,N_16770,N_15442);
nand U20136 (N_20136,N_19019,N_16785);
or U20137 (N_20137,N_18751,N_17424);
or U20138 (N_20138,N_16428,N_15738);
xor U20139 (N_20139,N_16803,N_19108);
or U20140 (N_20140,N_19190,N_17458);
xnor U20141 (N_20141,N_17943,N_18638);
nor U20142 (N_20142,N_18146,N_17132);
xnor U20143 (N_20143,N_17577,N_18862);
nand U20144 (N_20144,N_17579,N_18179);
nand U20145 (N_20145,N_18908,N_15263);
xor U20146 (N_20146,N_19181,N_19880);
nor U20147 (N_20147,N_17642,N_16301);
and U20148 (N_20148,N_16443,N_15627);
xor U20149 (N_20149,N_17961,N_19741);
xnor U20150 (N_20150,N_17160,N_18969);
nand U20151 (N_20151,N_17760,N_19524);
or U20152 (N_20152,N_19139,N_16099);
nand U20153 (N_20153,N_15784,N_17802);
and U20154 (N_20154,N_15352,N_16844);
nor U20155 (N_20155,N_19035,N_19384);
nor U20156 (N_20156,N_18721,N_19615);
or U20157 (N_20157,N_15209,N_18269);
or U20158 (N_20158,N_18772,N_15847);
nand U20159 (N_20159,N_16241,N_19437);
nand U20160 (N_20160,N_15126,N_18322);
and U20161 (N_20161,N_17867,N_16562);
and U20162 (N_20162,N_18571,N_19206);
xnor U20163 (N_20163,N_18847,N_18117);
and U20164 (N_20164,N_19761,N_15906);
xor U20165 (N_20165,N_15257,N_18684);
and U20166 (N_20166,N_18868,N_15985);
or U20167 (N_20167,N_19111,N_19386);
nand U20168 (N_20168,N_15377,N_16008);
and U20169 (N_20169,N_15290,N_17982);
nor U20170 (N_20170,N_17434,N_15059);
or U20171 (N_20171,N_17364,N_18510);
nor U20172 (N_20172,N_18389,N_17650);
nand U20173 (N_20173,N_19983,N_18664);
or U20174 (N_20174,N_18031,N_18596);
or U20175 (N_20175,N_15835,N_18691);
nor U20176 (N_20176,N_15626,N_15131);
xnor U20177 (N_20177,N_16597,N_15177);
xor U20178 (N_20178,N_17855,N_16742);
xor U20179 (N_20179,N_17615,N_16795);
nand U20180 (N_20180,N_17093,N_16687);
and U20181 (N_20181,N_18677,N_18229);
xnor U20182 (N_20182,N_18416,N_15136);
and U20183 (N_20183,N_19267,N_15127);
and U20184 (N_20184,N_18015,N_17371);
xnor U20185 (N_20185,N_19829,N_18268);
and U20186 (N_20186,N_18660,N_19369);
nand U20187 (N_20187,N_18084,N_15902);
or U20188 (N_20188,N_18489,N_15300);
nand U20189 (N_20189,N_16971,N_19565);
nand U20190 (N_20190,N_18864,N_18569);
or U20191 (N_20191,N_19608,N_16318);
xor U20192 (N_20192,N_18440,N_19695);
and U20193 (N_20193,N_18290,N_15765);
nor U20194 (N_20194,N_15803,N_18710);
and U20195 (N_20195,N_16787,N_16234);
and U20196 (N_20196,N_18737,N_16256);
nor U20197 (N_20197,N_16727,N_18766);
and U20198 (N_20198,N_19357,N_17813);
nand U20199 (N_20199,N_19663,N_18483);
nand U20200 (N_20200,N_18174,N_18408);
or U20201 (N_20201,N_17360,N_18560);
nand U20202 (N_20202,N_16181,N_17571);
xnor U20203 (N_20203,N_16867,N_15448);
or U20204 (N_20204,N_15322,N_19789);
xor U20205 (N_20205,N_17887,N_17077);
nand U20206 (N_20206,N_16996,N_18678);
or U20207 (N_20207,N_18997,N_18021);
nand U20208 (N_20208,N_16048,N_18400);
or U20209 (N_20209,N_16492,N_19593);
and U20210 (N_20210,N_19144,N_17480);
xnor U20211 (N_20211,N_15278,N_17521);
xor U20212 (N_20212,N_15797,N_18296);
or U20213 (N_20213,N_19168,N_16201);
or U20214 (N_20214,N_18851,N_18548);
xor U20215 (N_20215,N_18674,N_17990);
nand U20216 (N_20216,N_16665,N_18258);
nor U20217 (N_20217,N_15695,N_19988);
nor U20218 (N_20218,N_15224,N_15576);
nand U20219 (N_20219,N_19844,N_19688);
or U20220 (N_20220,N_17346,N_15953);
nand U20221 (N_20221,N_17465,N_17635);
or U20222 (N_20222,N_15168,N_17556);
xnor U20223 (N_20223,N_18890,N_16752);
or U20224 (N_20224,N_17253,N_19031);
nand U20225 (N_20225,N_19862,N_15995);
nor U20226 (N_20226,N_19196,N_16704);
nor U20227 (N_20227,N_16956,N_19447);
or U20228 (N_20228,N_16864,N_17245);
xor U20229 (N_20229,N_18506,N_17047);
xnor U20230 (N_20230,N_15885,N_15480);
xnor U20231 (N_20231,N_17840,N_16045);
nor U20232 (N_20232,N_18756,N_15640);
nand U20233 (N_20233,N_16725,N_18663);
nor U20234 (N_20234,N_18564,N_18849);
nand U20235 (N_20235,N_17841,N_17241);
or U20236 (N_20236,N_15537,N_15994);
nand U20237 (N_20237,N_15727,N_16713);
xnor U20238 (N_20238,N_18667,N_17210);
nand U20239 (N_20239,N_19734,N_18948);
or U20240 (N_20240,N_18673,N_15092);
nand U20241 (N_20241,N_17454,N_19269);
or U20242 (N_20242,N_19332,N_19194);
or U20243 (N_20243,N_15226,N_18566);
or U20244 (N_20244,N_15759,N_15383);
nor U20245 (N_20245,N_15820,N_17232);
nand U20246 (N_20246,N_19364,N_15407);
xor U20247 (N_20247,N_18463,N_17380);
xnor U20248 (N_20248,N_17731,N_16321);
nor U20249 (N_20249,N_18671,N_18532);
nor U20250 (N_20250,N_15398,N_19216);
xor U20251 (N_20251,N_15612,N_15066);
nand U20252 (N_20252,N_16347,N_17200);
and U20253 (N_20253,N_19881,N_18881);
and U20254 (N_20254,N_16745,N_17379);
xnor U20255 (N_20255,N_16862,N_16780);
and U20256 (N_20256,N_16556,N_16657);
xor U20257 (N_20257,N_16635,N_18017);
or U20258 (N_20258,N_17069,N_18989);
and U20259 (N_20259,N_19564,N_17934);
nand U20260 (N_20260,N_19897,N_17971);
or U20261 (N_20261,N_18546,N_19199);
nor U20262 (N_20262,N_17595,N_17020);
xor U20263 (N_20263,N_15529,N_19596);
and U20264 (N_20264,N_15072,N_19843);
nand U20265 (N_20265,N_19195,N_16130);
xor U20266 (N_20266,N_18061,N_19276);
nand U20267 (N_20267,N_15745,N_18261);
xor U20268 (N_20268,N_17886,N_15645);
and U20269 (N_20269,N_16271,N_17869);
nand U20270 (N_20270,N_15366,N_18741);
or U20271 (N_20271,N_15221,N_16056);
nand U20272 (N_20272,N_18966,N_15621);
and U20273 (N_20273,N_15458,N_17564);
nand U20274 (N_20274,N_19799,N_15690);
and U20275 (N_20275,N_19165,N_15818);
and U20276 (N_20276,N_19291,N_16266);
or U20277 (N_20277,N_15686,N_16616);
nor U20278 (N_20278,N_15683,N_18696);
nor U20279 (N_20279,N_19992,N_16085);
nand U20280 (N_20280,N_18689,N_19151);
or U20281 (N_20281,N_19951,N_19649);
nor U20282 (N_20282,N_19424,N_18505);
and U20283 (N_20283,N_18839,N_15862);
or U20284 (N_20284,N_17900,N_17935);
or U20285 (N_20285,N_16031,N_17365);
or U20286 (N_20286,N_19468,N_15085);
and U20287 (N_20287,N_19956,N_16276);
nand U20288 (N_20288,N_17459,N_19572);
nor U20289 (N_20289,N_15550,N_15897);
nor U20290 (N_20290,N_15564,N_16132);
nand U20291 (N_20291,N_15010,N_19810);
or U20292 (N_20292,N_18438,N_17570);
nor U20293 (N_20293,N_16212,N_17491);
and U20294 (N_20294,N_18809,N_19922);
and U20295 (N_20295,N_18411,N_17254);
nor U20296 (N_20296,N_18402,N_17870);
or U20297 (N_20297,N_19484,N_17598);
xnor U20298 (N_20298,N_16512,N_15761);
xor U20299 (N_20299,N_15535,N_16574);
nor U20300 (N_20300,N_17389,N_17786);
or U20301 (N_20301,N_18796,N_18617);
xor U20302 (N_20302,N_17332,N_16587);
xnor U20303 (N_20303,N_16916,N_15907);
nor U20304 (N_20304,N_15239,N_15280);
xor U20305 (N_20305,N_19657,N_18018);
nor U20306 (N_20306,N_16182,N_17211);
nand U20307 (N_20307,N_16066,N_19105);
and U20308 (N_20308,N_18845,N_15277);
nand U20309 (N_20309,N_19017,N_16352);
nand U20310 (N_20310,N_16503,N_16603);
or U20311 (N_20311,N_17262,N_17784);
nand U20312 (N_20312,N_19847,N_15998);
nor U20313 (N_20313,N_17624,N_19141);
xor U20314 (N_20314,N_16940,N_15531);
nor U20315 (N_20315,N_17357,N_17794);
or U20316 (N_20316,N_16546,N_17916);
xnor U20317 (N_20317,N_17849,N_15736);
or U20318 (N_20318,N_18711,N_17269);
xor U20319 (N_20319,N_15315,N_18434);
nand U20320 (N_20320,N_19807,N_17268);
xnor U20321 (N_20321,N_17967,N_15254);
xor U20322 (N_20322,N_17436,N_19508);
nand U20323 (N_20323,N_16720,N_18764);
and U20324 (N_20324,N_19429,N_15067);
or U20325 (N_20325,N_18150,N_18668);
nand U20326 (N_20326,N_19979,N_16756);
or U20327 (N_20327,N_16280,N_18284);
or U20328 (N_20328,N_19065,N_16420);
or U20329 (N_20329,N_18273,N_15628);
and U20330 (N_20330,N_17300,N_19840);
nor U20331 (N_20331,N_16566,N_15997);
nand U20332 (N_20332,N_17532,N_15336);
nand U20333 (N_20333,N_15712,N_15427);
and U20334 (N_20334,N_19242,N_16604);
xor U20335 (N_20335,N_16539,N_15342);
or U20336 (N_20336,N_16708,N_18950);
nand U20337 (N_20337,N_15034,N_19319);
or U20338 (N_20338,N_15511,N_17625);
xor U20339 (N_20339,N_19791,N_19057);
and U20340 (N_20340,N_17054,N_17774);
and U20341 (N_20341,N_16507,N_18022);
and U20342 (N_20342,N_16789,N_17178);
nor U20343 (N_20343,N_18155,N_16039);
and U20344 (N_20344,N_18878,N_16230);
nor U20345 (N_20345,N_16423,N_17746);
nand U20346 (N_20346,N_19491,N_19232);
nand U20347 (N_20347,N_16870,N_18531);
nand U20348 (N_20348,N_15436,N_16038);
or U20349 (N_20349,N_19820,N_18493);
and U20350 (N_20350,N_15378,N_18289);
and U20351 (N_20351,N_18610,N_18144);
nand U20352 (N_20352,N_16035,N_16490);
nand U20353 (N_20353,N_15586,N_18028);
xnor U20354 (N_20354,N_17899,N_18497);
nand U20355 (N_20355,N_19738,N_19315);
or U20356 (N_20356,N_18317,N_17315);
or U20357 (N_20357,N_15552,N_18653);
nand U20358 (N_20358,N_19839,N_16437);
and U20359 (N_20359,N_17536,N_15494);
nor U20360 (N_20360,N_15606,N_19574);
xnor U20361 (N_20361,N_17552,N_15984);
nand U20362 (N_20362,N_16627,N_16027);
or U20363 (N_20363,N_15065,N_15934);
and U20364 (N_20364,N_15397,N_19215);
and U20365 (N_20365,N_19909,N_19609);
xor U20366 (N_20366,N_15415,N_16124);
nand U20367 (N_20367,N_15982,N_15993);
xor U20368 (N_20368,N_15949,N_15574);
xnor U20369 (N_20369,N_18520,N_19028);
nand U20370 (N_20370,N_16922,N_19834);
nand U20371 (N_20371,N_18744,N_17363);
and U20372 (N_20372,N_18372,N_18473);
nor U20373 (N_20373,N_15350,N_18134);
xnor U20374 (N_20374,N_19085,N_18648);
and U20375 (N_20375,N_16023,N_15148);
xnor U20376 (N_20376,N_16337,N_18374);
xnor U20377 (N_20377,N_16491,N_15634);
and U20378 (N_20378,N_15571,N_17293);
nor U20379 (N_20379,N_15567,N_15910);
nor U20380 (N_20380,N_19803,N_18462);
nand U20381 (N_20381,N_19549,N_17837);
nor U20382 (N_20382,N_19214,N_18293);
nand U20383 (N_20383,N_16223,N_15861);
nor U20384 (N_20384,N_19800,N_16598);
xnor U20385 (N_20385,N_16125,N_18488);
nand U20386 (N_20386,N_15393,N_17894);
nor U20387 (N_20387,N_15255,N_19821);
nor U20388 (N_20388,N_16480,N_16849);
xor U20389 (N_20389,N_18657,N_15332);
or U20390 (N_20390,N_17715,N_18821);
or U20391 (N_20391,N_18315,N_18328);
or U20392 (N_20392,N_16393,N_19547);
nand U20393 (N_20393,N_15304,N_17329);
xor U20394 (N_20394,N_19305,N_16655);
nor U20395 (N_20395,N_19174,N_18020);
and U20396 (N_20396,N_15104,N_16133);
nand U20397 (N_20397,N_19090,N_19230);
and U20398 (N_20398,N_18382,N_17500);
xor U20399 (N_20399,N_17511,N_17645);
xor U20400 (N_20400,N_19262,N_16036);
nor U20401 (N_20401,N_19379,N_17791);
and U20402 (N_20402,N_16483,N_15705);
xor U20403 (N_20403,N_16680,N_19505);
and U20404 (N_20404,N_17089,N_19611);
or U20405 (N_20405,N_19323,N_15565);
nand U20406 (N_20406,N_19772,N_18194);
or U20407 (N_20407,N_16178,N_19107);
and U20408 (N_20408,N_15295,N_16406);
nor U20409 (N_20409,N_17242,N_15778);
nand U20410 (N_20410,N_19353,N_19630);
nand U20411 (N_20411,N_17473,N_16494);
or U20412 (N_20412,N_19180,N_18234);
nand U20413 (N_20413,N_15828,N_17071);
or U20414 (N_20414,N_19118,N_17629);
nor U20415 (N_20415,N_17128,N_19752);
xor U20416 (N_20416,N_18728,N_16544);
or U20417 (N_20417,N_15368,N_16506);
xor U20418 (N_20418,N_19240,N_15120);
nor U20419 (N_20419,N_19189,N_15713);
or U20420 (N_20420,N_16533,N_16398);
nand U20421 (N_20421,N_18025,N_18976);
nor U20422 (N_20422,N_15076,N_17163);
or U20423 (N_20423,N_18854,N_15566);
nor U20424 (N_20424,N_17888,N_18454);
xnor U20425 (N_20425,N_19336,N_19627);
or U20426 (N_20426,N_18938,N_18339);
nand U20427 (N_20427,N_16359,N_17718);
or U20428 (N_20428,N_16896,N_17429);
nor U20429 (N_20429,N_19004,N_18056);
nor U20430 (N_20430,N_18259,N_18407);
nor U20431 (N_20431,N_15622,N_18565);
or U20432 (N_20432,N_18904,N_17024);
nor U20433 (N_20433,N_16830,N_19275);
nor U20434 (N_20434,N_16317,N_17117);
nor U20435 (N_20435,N_19792,N_16555);
nor U20436 (N_20436,N_17636,N_19977);
and U20437 (N_20437,N_15401,N_15681);
nor U20438 (N_20438,N_18567,N_18661);
xor U20439 (N_20439,N_18385,N_16654);
nor U20440 (N_20440,N_15486,N_17602);
and U20441 (N_20441,N_18633,N_17798);
or U20442 (N_20442,N_18104,N_15262);
nand U20443 (N_20443,N_15070,N_16154);
and U20444 (N_20444,N_16067,N_15959);
xor U20445 (N_20445,N_15197,N_18067);
and U20446 (N_20446,N_19867,N_18043);
nor U20447 (N_20447,N_15754,N_16243);
xor U20448 (N_20448,N_15886,N_16100);
or U20449 (N_20449,N_15813,N_17442);
xnor U20450 (N_20450,N_16632,N_16877);
or U20451 (N_20451,N_16002,N_19200);
xor U20452 (N_20452,N_19119,N_17305);
xor U20453 (N_20453,N_15175,N_15455);
nand U20454 (N_20454,N_16387,N_15514);
or U20455 (N_20455,N_17957,N_16573);
and U20456 (N_20456,N_17509,N_15101);
or U20457 (N_20457,N_15268,N_17167);
nor U20458 (N_20458,N_15250,N_19971);
and U20459 (N_20459,N_15203,N_19614);
nand U20460 (N_20460,N_16794,N_19521);
or U20461 (N_20461,N_17843,N_16377);
nand U20462 (N_20462,N_15253,N_17359);
nor U20463 (N_20463,N_15100,N_16348);
and U20464 (N_20464,N_16880,N_16466);
nand U20465 (N_20465,N_16268,N_17409);
or U20466 (N_20466,N_19338,N_17638);
xor U20467 (N_20467,N_15408,N_17376);
or U20468 (N_20468,N_19591,N_19055);
nor U20469 (N_20469,N_19928,N_18354);
xor U20470 (N_20470,N_16073,N_19525);
xnor U20471 (N_20471,N_15411,N_17324);
nand U20472 (N_20472,N_17411,N_17391);
nor U20473 (N_20473,N_16362,N_17893);
nand U20474 (N_20474,N_18699,N_16621);
xnor U20475 (N_20475,N_16783,N_17616);
xor U20476 (N_20476,N_19446,N_19914);
xor U20477 (N_20477,N_16227,N_18130);
nor U20478 (N_20478,N_18464,N_17809);
or U20479 (N_20479,N_18848,N_16438);
nor U20480 (N_20480,N_17001,N_18870);
nand U20481 (N_20481,N_19570,N_16840);
xnor U20482 (N_20482,N_17204,N_18096);
nand U20483 (N_20483,N_17852,N_18882);
xnor U20484 (N_20484,N_16802,N_19069);
nor U20485 (N_20485,N_19355,N_15663);
or U20486 (N_20486,N_19405,N_19399);
or U20487 (N_20487,N_17604,N_18014);
nor U20488 (N_20488,N_16297,N_19628);
or U20489 (N_20489,N_18647,N_15184);
nor U20490 (N_20490,N_17238,N_16949);
or U20491 (N_20491,N_15275,N_15962);
nand U20492 (N_20492,N_15559,N_15737);
and U20493 (N_20493,N_18223,N_18693);
nor U20494 (N_20494,N_19801,N_19394);
nor U20495 (N_20495,N_17696,N_16292);
nor U20496 (N_20496,N_16965,N_17052);
nand U20497 (N_20497,N_18311,N_16174);
and U20498 (N_20498,N_15578,N_17277);
xor U20499 (N_20499,N_18987,N_19532);
and U20500 (N_20500,N_19646,N_15488);
nand U20501 (N_20501,N_19449,N_17671);
xor U20502 (N_20502,N_15602,N_15016);
xnor U20503 (N_20503,N_17589,N_19997);
and U20504 (N_20504,N_15008,N_15173);
and U20505 (N_20505,N_18256,N_16514);
and U20506 (N_20506,N_18630,N_19845);
or U20507 (N_20507,N_18947,N_16208);
or U20508 (N_20508,N_16467,N_17419);
and U20509 (N_20509,N_17712,N_17014);
or U20510 (N_20510,N_19982,N_16945);
xor U20511 (N_20511,N_19599,N_18283);
and U20512 (N_20512,N_18698,N_15056);
xnor U20513 (N_20513,N_15762,N_15425);
xnor U20514 (N_20514,N_19773,N_17037);
nor U20515 (N_20515,N_16298,N_18222);
nor U20516 (N_20516,N_19371,N_19516);
or U20517 (N_20517,N_17392,N_19546);
nor U20518 (N_20518,N_19755,N_15721);
and U20519 (N_20519,N_16837,N_17435);
or U20520 (N_20520,N_15354,N_18088);
nor U20521 (N_20521,N_15426,N_18388);
xor U20522 (N_20522,N_18823,N_18091);
nand U20523 (N_20523,N_19340,N_15047);
and U20524 (N_20524,N_15804,N_17481);
or U20525 (N_20525,N_19664,N_16640);
and U20526 (N_20526,N_16656,N_16329);
nor U20527 (N_20527,N_15191,N_15517);
nand U20528 (N_20528,N_15205,N_16005);
xor U20529 (N_20529,N_16367,N_19605);
and U20530 (N_20530,N_17279,N_18112);
and U20531 (N_20531,N_15633,N_15889);
xor U20532 (N_20532,N_18594,N_18059);
and U20533 (N_20533,N_16237,N_17367);
nor U20534 (N_20534,N_17149,N_16898);
xnor U20535 (N_20535,N_17622,N_17381);
or U20536 (N_20536,N_15491,N_17667);
and U20537 (N_20537,N_18192,N_19226);
or U20538 (N_20538,N_17447,N_16260);
or U20539 (N_20539,N_16902,N_17013);
xnor U20540 (N_20540,N_16150,N_19387);
nand U20541 (N_20541,N_17239,N_18512);
and U20542 (N_20542,N_15605,N_18461);
nor U20543 (N_20543,N_18866,N_19227);
nor U20544 (N_20544,N_15081,N_17621);
and U20545 (N_20545,N_17078,N_19354);
or U20546 (N_20546,N_15850,N_15308);
nand U20547 (N_20547,N_17915,N_15728);
or U20548 (N_20548,N_17516,N_19783);
and U20549 (N_20549,N_16046,N_15655);
xor U20550 (N_20550,N_18108,N_16123);
nor U20551 (N_20551,N_15689,N_17066);
xor U20552 (N_20552,N_19294,N_18906);
xor U20553 (N_20553,N_18396,N_15826);
and U20554 (N_20554,N_18863,N_19957);
nor U20555 (N_20555,N_19131,N_16033);
nand U20556 (N_20556,N_15903,N_18611);
and U20557 (N_20557,N_17095,N_18384);
and U20558 (N_20558,N_19251,N_18316);
nor U20559 (N_20559,N_15319,N_17573);
or U20560 (N_20560,N_18869,N_16617);
or U20561 (N_20561,N_15298,N_17593);
nand U20562 (N_20562,N_18037,N_17444);
and U20563 (N_20563,N_18123,N_18419);
xnor U20564 (N_20564,N_17467,N_19968);
xnor U20565 (N_20565,N_16262,N_16757);
nand U20566 (N_20566,N_16968,N_16460);
nand U20567 (N_20567,N_16979,N_15068);
nor U20568 (N_20568,N_15942,N_16434);
xnor U20569 (N_20569,N_18800,N_15752);
nor U20570 (N_20570,N_17180,N_17572);
nand U20571 (N_20571,N_17755,N_17012);
nor U20572 (N_20572,N_15036,N_16863);
nor U20573 (N_20573,N_18719,N_17942);
or U20574 (N_20574,N_16436,N_16927);
and U20575 (N_20575,N_16924,N_15199);
nand U20576 (N_20576,N_18195,N_17865);
nor U20577 (N_20577,N_17428,N_16088);
xor U20578 (N_20578,N_19687,N_18920);
or U20579 (N_20579,N_16011,N_19212);
nand U20580 (N_20580,N_15140,N_16548);
nor U20581 (N_20581,N_15808,N_18871);
nor U20582 (N_20582,N_15302,N_19128);
nor U20583 (N_20583,N_15549,N_18079);
and U20584 (N_20584,N_17781,N_18136);
nor U20585 (N_20585,N_17331,N_16610);
and U20586 (N_20586,N_18139,N_17683);
nor U20587 (N_20587,N_17307,N_15475);
nor U20588 (N_20588,N_18115,N_15641);
nand U20589 (N_20589,N_17926,N_16733);
nor U20590 (N_20590,N_16338,N_17133);
nand U20591 (N_20591,N_18746,N_19879);
or U20592 (N_20592,N_15305,N_19071);
xnor U20593 (N_20593,N_15492,N_16184);
nor U20594 (N_20594,N_15595,N_15581);
or U20595 (N_20595,N_19470,N_18141);
or U20596 (N_20596,N_15933,N_19900);
xor U20597 (N_20597,N_15323,N_15132);
xor U20598 (N_20598,N_19893,N_17989);
xnor U20599 (N_20599,N_15150,N_16515);
and U20600 (N_20600,N_15137,N_19188);
nor U20601 (N_20601,N_19952,N_19855);
or U20602 (N_20602,N_17681,N_16057);
nand U20603 (N_20603,N_16198,N_18518);
nand U20604 (N_20604,N_18185,N_16247);
or U20605 (N_20605,N_18919,N_18356);
and U20606 (N_20606,N_17361,N_16500);
xnor U20607 (N_20607,N_16274,N_19647);
nor U20608 (N_20608,N_16136,N_19802);
nor U20609 (N_20609,N_16288,N_17995);
nand U20610 (N_20610,N_16092,N_16137);
or U20611 (N_20611,N_15296,N_18618);
xnor U20612 (N_20612,N_19086,N_16739);
xnor U20613 (N_20613,N_18032,N_18996);
nor U20614 (N_20614,N_15548,N_15742);
or U20615 (N_20615,N_19947,N_16164);
or U20616 (N_20616,N_16818,N_16007);
or U20617 (N_20617,N_15815,N_17606);
nand U20618 (N_20618,N_15283,N_18978);
xnor U20619 (N_20619,N_15212,N_17779);
nand U20620 (N_20620,N_17192,N_18053);
or U20621 (N_20621,N_19966,N_17910);
and U20622 (N_20622,N_18367,N_18982);
nand U20623 (N_20623,N_19503,N_18080);
nor U20624 (N_20624,N_15452,N_17000);
or U20625 (N_20625,N_17079,N_16791);
xnor U20626 (N_20626,N_19253,N_16098);
and U20627 (N_20627,N_17825,N_18713);
xor U20628 (N_20628,N_18580,N_18365);
and U20629 (N_20629,N_15698,N_19089);
xor U20630 (N_20630,N_17256,N_16645);
and U20631 (N_20631,N_19460,N_16391);
nand U20632 (N_20632,N_18544,N_19094);
or U20633 (N_20633,N_15834,N_15023);
and U20634 (N_20634,N_15631,N_19158);
or U20635 (N_20635,N_17727,N_18167);
nor U20636 (N_20636,N_17785,N_16072);
nor U20637 (N_20637,N_19281,N_15810);
xnor U20638 (N_20638,N_17864,N_15404);
xnor U20639 (N_20639,N_19644,N_16026);
nor U20640 (N_20640,N_18650,N_15071);
xnor U20641 (N_20641,N_17130,N_18055);
and U20642 (N_20642,N_17390,N_19967);
or U20643 (N_20643,N_15259,N_16439);
or U20644 (N_20644,N_19260,N_19382);
and U20645 (N_20645,N_16053,N_15499);
xor U20646 (N_20646,N_19776,N_19049);
or U20647 (N_20647,N_17749,N_15992);
or U20648 (N_20648,N_18655,N_17383);
nor U20649 (N_20649,N_17567,N_16074);
nand U20650 (N_20650,N_16418,N_16340);
xor U20651 (N_20651,N_15487,N_19906);
xnor U20652 (N_20652,N_16248,N_18239);
or U20653 (N_20653,N_16217,N_17131);
nor U20654 (N_20654,N_16962,N_18040);
xnor U20655 (N_20655,N_15607,N_17815);
and U20656 (N_20656,N_19770,N_19523);
nor U20657 (N_20657,N_15052,N_17113);
and U20658 (N_20658,N_16077,N_18118);
or U20659 (N_20659,N_15747,N_19699);
or U20660 (N_20660,N_18490,N_19040);
nor U20661 (N_20661,N_19632,N_17684);
nand U20662 (N_20662,N_17605,N_17124);
and U20663 (N_20663,N_17766,N_15766);
nand U20664 (N_20664,N_16134,N_17523);
nor U20665 (N_20665,N_17998,N_18252);
or U20666 (N_20666,N_16762,N_17545);
nand U20667 (N_20667,N_16817,N_15417);
xor U20668 (N_20668,N_18861,N_18593);
or U20669 (N_20669,N_19217,N_15208);
xor U20670 (N_20670,N_19436,N_16309);
or U20671 (N_20671,N_19273,N_15749);
xor U20672 (N_20672,N_18158,N_18867);
and U20673 (N_20673,N_19155,N_16674);
nor U20674 (N_20674,N_18441,N_19707);
nand U20675 (N_20675,N_17395,N_18401);
nor U20676 (N_20676,N_19563,N_18831);
xnor U20677 (N_20677,N_18156,N_19346);
xor U20678 (N_20678,N_15348,N_15543);
or U20679 (N_20679,N_18833,N_18499);
nor U20680 (N_20680,N_19625,N_18875);
nand U20681 (N_20681,N_15146,N_15812);
and U20682 (N_20682,N_19754,N_15963);
nand U20683 (N_20683,N_19877,N_16828);
and U20684 (N_20684,N_18859,N_17590);
nand U20685 (N_20685,N_19713,N_16214);
and U20686 (N_20686,N_18126,N_19700);
xnor U20687 (N_20687,N_15077,N_15405);
xnor U20688 (N_20688,N_15706,N_18585);
nor U20689 (N_20689,N_16866,N_15796);
nor U20690 (N_20690,N_18324,N_15453);
or U20691 (N_20691,N_16517,N_16455);
nor U20692 (N_20692,N_18077,N_19742);
nand U20693 (N_20693,N_19530,N_18926);
nand U20694 (N_20694,N_16559,N_16911);
and U20695 (N_20695,N_18923,N_15665);
nand U20696 (N_20696,N_17485,N_17275);
or U20697 (N_20697,N_16485,N_17343);
xnor U20698 (N_20698,N_17495,N_16853);
xnor U20699 (N_20699,N_18551,N_16951);
nor U20700 (N_20700,N_19626,N_19674);
nand U20701 (N_20701,N_16964,N_19835);
nand U20702 (N_20702,N_18333,N_15000);
xnor U20703 (N_20703,N_18535,N_18165);
nand U20704 (N_20704,N_19106,N_18318);
nor U20705 (N_20705,N_17951,N_18487);
nand U20706 (N_20706,N_17246,N_16932);
nor U20707 (N_20707,N_16758,N_15096);
or U20708 (N_20708,N_17721,N_15868);
or U20709 (N_20709,N_17187,N_18299);
xor U20710 (N_20710,N_19555,N_19014);
nand U20711 (N_20711,N_18477,N_18708);
and U20712 (N_20712,N_18453,N_16353);
xor U20713 (N_20713,N_18206,N_16948);
and U20714 (N_20714,N_17845,N_17041);
nor U20715 (N_20715,N_15159,N_15584);
nand U20716 (N_20716,N_15374,N_18265);
nor U20717 (N_20717,N_19012,N_18176);
nand U20718 (N_20718,N_19471,N_16478);
or U20719 (N_20719,N_16146,N_17639);
nand U20720 (N_20720,N_16385,N_19415);
and U20721 (N_20721,N_15616,N_15943);
and U20722 (N_20722,N_16706,N_18092);
nor U20723 (N_20723,N_18332,N_16993);
or U20724 (N_20724,N_18577,N_15055);
nand U20725 (N_20725,N_16567,N_16369);
xnor U20726 (N_20726,N_18730,N_15053);
nor U20727 (N_20727,N_18236,N_16101);
nand U20728 (N_20728,N_19606,N_18909);
xnor U20729 (N_20729,N_15838,N_15913);
xor U20730 (N_20730,N_16589,N_15260);
and U20731 (N_20731,N_15504,N_18643);
nor U20732 (N_20732,N_18457,N_15185);
nand U20733 (N_20733,N_15961,N_16021);
and U20734 (N_20734,N_16113,N_15320);
nor U20735 (N_20735,N_17762,N_15554);
or U20736 (N_20736,N_16354,N_16740);
nand U20737 (N_20737,N_19345,N_18805);
or U20738 (N_20738,N_16550,N_16376);
or U20739 (N_20739,N_18992,N_15845);
nand U20740 (N_20740,N_16814,N_16462);
nor U20741 (N_20741,N_15284,N_16222);
nand U20742 (N_20742,N_17203,N_19074);
and U20743 (N_20743,N_18286,N_18065);
nor U20744 (N_20744,N_19875,N_19712);
and U20745 (N_20745,N_15666,N_18319);
nand U20746 (N_20746,N_16670,N_15134);
and U20747 (N_20747,N_16554,N_16717);
nor U20748 (N_20748,N_15716,N_18550);
and U20749 (N_20749,N_15447,N_17687);
xnor U20750 (N_20750,N_15693,N_17296);
or U20751 (N_20751,N_17640,N_16142);
or U20752 (N_20752,N_17737,N_18274);
nand U20753 (N_20753,N_15243,N_16601);
and U20754 (N_20754,N_18707,N_19766);
or U20755 (N_20755,N_15888,N_17061);
and U20756 (N_20756,N_15597,N_15133);
nand U20757 (N_20757,N_16175,N_16191);
and U20758 (N_20758,N_15895,N_18012);
xnor U20759 (N_20759,N_16479,N_16839);
xnor U20760 (N_20760,N_15505,N_17931);
xor U20761 (N_20761,N_19254,N_15877);
nor U20762 (N_20762,N_19274,N_17873);
xor U20763 (N_20763,N_18767,N_16831);
xnor U20764 (N_20764,N_15764,N_16832);
nand U20765 (N_20765,N_16957,N_16935);
and U20766 (N_20766,N_19073,N_18748);
or U20767 (N_20767,N_19009,N_15746);
nand U20768 (N_20768,N_19537,N_18540);
and U20769 (N_20769,N_19883,N_18069);
and U20770 (N_20770,N_17952,N_17723);
nor U20771 (N_20771,N_15900,N_15031);
nor U20772 (N_20772,N_16499,N_19899);
and U20773 (N_20773,N_17219,N_19866);
or U20774 (N_20774,N_18302,N_17905);
and U20775 (N_20775,N_16187,N_18945);
xnor U20776 (N_20776,N_18242,N_18491);
xor U20777 (N_20777,N_19327,N_19497);
or U20778 (N_20778,N_15182,N_15708);
nor U20779 (N_20779,N_18999,N_17947);
nand U20780 (N_20780,N_19691,N_17081);
nor U20781 (N_20781,N_19701,N_19109);
or U20782 (N_20782,N_18977,N_17354);
nand U20783 (N_20783,N_18429,N_18478);
or U20784 (N_20784,N_16064,N_15688);
or U20785 (N_20785,N_17596,N_17212);
nor U20786 (N_20786,N_17055,N_18597);
nor U20787 (N_20787,N_17286,N_19476);
and U20788 (N_20788,N_16051,N_16792);
nand U20789 (N_20789,N_18883,N_15015);
nor U20790 (N_20790,N_15572,N_19329);
or U20791 (N_20791,N_15012,N_17568);
or U20792 (N_20792,N_15901,N_16985);
and U20793 (N_20793,N_16270,N_16570);
and U20794 (N_20794,N_18216,N_16311);
and U20795 (N_20795,N_18113,N_18701);
or U20796 (N_20796,N_17691,N_18717);
nor U20797 (N_20797,N_19585,N_17188);
xnor U20798 (N_20798,N_17171,N_16213);
nand U20799 (N_20799,N_18980,N_18094);
nor U20800 (N_20800,N_15247,N_19653);
nand U20801 (N_20801,N_17208,N_15266);
or U20802 (N_20802,N_15856,N_19192);
nand U20803 (N_20803,N_17034,N_15496);
or U20804 (N_20804,N_18940,N_18033);
and U20805 (N_20805,N_19452,N_17221);
and U20806 (N_20806,N_19680,N_16812);
nand U20807 (N_20807,N_19590,N_18616);
xnor U20808 (N_20808,N_18917,N_19495);
nor U20809 (N_20809,N_19417,N_16703);
or U20810 (N_20810,N_19159,N_17729);
xnor U20811 (N_20811,N_16983,N_15235);
nand U20812 (N_20812,N_17312,N_19804);
nor U20813 (N_20813,N_19735,N_16875);
nand U20814 (N_20814,N_17311,N_19072);
nand U20815 (N_20815,N_18576,N_17919);
xnor U20816 (N_20816,N_19654,N_19024);
nand U20817 (N_20817,N_17652,N_16219);
nand U20818 (N_20818,N_18771,N_19290);
and U20819 (N_20819,N_17892,N_18095);
nand U20820 (N_20820,N_16349,N_18172);
or U20821 (N_20821,N_17377,N_19473);
nand U20822 (N_20822,N_17747,N_16796);
or U20823 (N_20823,N_17617,N_17806);
xnor U20824 (N_20824,N_19358,N_17340);
nor U20825 (N_20825,N_17375,N_19235);
nor U20826 (N_20826,N_15211,N_19220);
and U20827 (N_20827,N_18439,N_18459);
and U20828 (N_20828,N_18656,N_16889);
and U20829 (N_20829,N_17613,N_15980);
nor U20830 (N_20830,N_15451,N_18011);
xor U20831 (N_20831,N_15316,N_19612);
xnor U20832 (N_20832,N_17678,N_18960);
xnor U20833 (N_20833,N_18383,N_17660);
xor U20834 (N_20834,N_16660,N_18853);
xor U20835 (N_20835,N_15966,N_19034);
and U20836 (N_20836,N_19138,N_17028);
nand U20837 (N_20837,N_15345,N_15083);
nor U20838 (N_20838,N_15054,N_18466);
nand U20839 (N_20839,N_19601,N_16760);
or U20840 (N_20840,N_18723,N_16044);
or U20841 (N_20841,N_18391,N_18305);
nor U20842 (N_20842,N_16180,N_18019);
nor U20843 (N_20843,N_15359,N_18386);
nor U20844 (N_20844,N_19607,N_15261);
and U20845 (N_20845,N_16509,N_16915);
xor U20846 (N_20846,N_16905,N_19425);
xnor U20847 (N_20847,N_18729,N_15702);
nor U20848 (N_20848,N_17288,N_18287);
and U20849 (N_20849,N_16663,N_19575);
xor U20850 (N_20850,N_16879,N_17417);
and U20851 (N_20851,N_16341,N_19292);
nand U20852 (N_20852,N_19366,N_18198);
xor U20853 (N_20853,N_19864,N_17833);
nand U20854 (N_20854,N_19683,N_15521);
nand U20855 (N_20855,N_18642,N_19257);
and U20856 (N_20856,N_15414,N_19309);
or U20857 (N_20857,N_18230,N_16861);
nor U20858 (N_20858,N_17431,N_18712);
xor U20859 (N_20859,N_17795,N_16228);
nor U20860 (N_20860,N_16189,N_18076);
xor U20861 (N_20861,N_16790,N_19308);
and U20862 (N_20862,N_17432,N_19624);
nand U20863 (N_20863,N_15293,N_19280);
nor U20864 (N_20864,N_19868,N_19825);
xor U20865 (N_20865,N_17783,N_15573);
or U20866 (N_20866,N_17217,N_18193);
and U20867 (N_20867,N_15986,N_18101);
nor U20868 (N_20868,N_15360,N_18704);
xnor U20869 (N_20869,N_15242,N_19767);
or U20870 (N_20870,N_19258,N_18237);
and U20871 (N_20871,N_19295,N_16296);
or U20872 (N_20872,N_19328,N_15317);
xnor U20873 (N_20873,N_15279,N_15237);
nor U20874 (N_20874,N_18715,N_18481);
and U20875 (N_20875,N_19414,N_18157);
nor U20876 (N_20876,N_15227,N_16264);
and U20877 (N_20877,N_15213,N_15842);
nor U20878 (N_20878,N_16457,N_19413);
nor U20879 (N_20879,N_17974,N_19703);
nor U20880 (N_20880,N_17854,N_16363);
or U20881 (N_20881,N_18679,N_18785);
nand U20882 (N_20882,N_15928,N_16343);
xor U20883 (N_20883,N_17597,N_19187);
or U20884 (N_20884,N_19428,N_15540);
xor U20885 (N_20885,N_15863,N_17958);
and U20886 (N_20886,N_18545,N_18353);
nand U20887 (N_20887,N_19769,N_18739);
xor U20888 (N_20888,N_19650,N_19686);
or U20889 (N_20889,N_17198,N_17317);
xor U20890 (N_20890,N_16310,N_16159);
nand U20891 (N_20891,N_17110,N_15512);
and U20892 (N_20892,N_18732,N_16624);
nand U20893 (N_20893,N_17105,N_18942);
nor U20894 (N_20894,N_15837,N_15624);
or U20895 (N_20895,N_19554,N_19439);
or U20896 (N_20896,N_19553,N_19518);
and U20897 (N_20897,N_17804,N_17539);
nor U20898 (N_20898,N_17932,N_15144);
and U20899 (N_20899,N_19682,N_15271);
xnor U20900 (N_20900,N_17118,N_15977);
nor U20901 (N_20901,N_15630,N_19403);
xor U20902 (N_20902,N_16661,N_15207);
nand U20903 (N_20903,N_15734,N_15195);
or U20904 (N_20904,N_16028,N_18670);
nor U20905 (N_20905,N_17879,N_15334);
xor U20906 (N_20906,N_18818,N_19147);
or U20907 (N_20907,N_17748,N_18747);
and U20908 (N_20908,N_18631,N_19768);
or U20909 (N_20909,N_18627,N_16767);
nor U20910 (N_20910,N_18188,N_19318);
nor U20911 (N_20911,N_15814,N_19985);
or U20912 (N_20912,N_16699,N_15830);
xor U20913 (N_20913,N_16676,N_19812);
xor U20914 (N_20914,N_17342,N_17918);
and U20915 (N_20915,N_17954,N_16784);
nor U20916 (N_20916,N_18826,N_16405);
and U20917 (N_20917,N_18087,N_17243);
nor U20918 (N_20918,N_15158,N_17714);
nand U20919 (N_20919,N_15241,N_19221);
nand U20920 (N_20920,N_19779,N_17778);
nand U20921 (N_20921,N_18676,N_19136);
and U20922 (N_20922,N_19182,N_17827);
and U20923 (N_20923,N_19137,N_17828);
and U20924 (N_20924,N_17226,N_15924);
nand U20925 (N_20925,N_19143,N_18846);
and U20926 (N_20926,N_17165,N_19958);
or U20927 (N_20927,N_19479,N_19715);
or U20928 (N_20928,N_16580,N_18320);
or U20929 (N_20929,N_17583,N_15500);
or U20930 (N_20930,N_19860,N_17120);
nor U20931 (N_20931,N_18583,N_19116);
nor U20932 (N_20932,N_17580,N_17964);
xor U20933 (N_20933,N_16854,N_15793);
xor U20934 (N_20934,N_15970,N_15858);
nor U20935 (N_20935,N_19842,N_19716);
xnor U20936 (N_20936,N_19283,N_18685);
nand U20937 (N_20937,N_17557,N_15026);
xnor U20938 (N_20938,N_16320,N_18953);
nand U20939 (N_20939,N_18390,N_16892);
xor U20940 (N_20940,N_17701,N_18241);
nor U20941 (N_20941,N_18447,N_18331);
and U20942 (N_20942,N_15623,N_16719);
and U20943 (N_20943,N_18620,N_15028);
nor U20944 (N_20944,N_15439,N_16083);
nor U20945 (N_20945,N_17656,N_16931);
xor U20946 (N_20946,N_15719,N_16006);
nor U20947 (N_20947,N_16540,N_15341);
and U20948 (N_20948,N_17373,N_17768);
xor U20949 (N_20949,N_19120,N_17690);
and U20950 (N_20950,N_18581,N_19539);
or U20951 (N_20951,N_15064,N_18394);
nor U20952 (N_20952,N_16112,N_15152);
or U20953 (N_20953,N_16402,N_19892);
or U20954 (N_20954,N_16231,N_18366);
xnor U20955 (N_20955,N_18437,N_19512);
nand U20956 (N_20956,N_18731,N_19763);
xnor U20957 (N_20957,N_17249,N_18034);
and U20958 (N_20958,N_17453,N_16392);
or U20959 (N_20959,N_19613,N_16613);
nand U20960 (N_20960,N_16003,N_16049);
nand U20961 (N_20961,N_19854,N_16012);
or U20962 (N_20962,N_18433,N_18397);
nand U20963 (N_20963,N_16557,N_15128);
xnor U20964 (N_20964,N_18456,N_18467);
nand U20965 (N_20965,N_18836,N_17139);
xor U20966 (N_20966,N_16923,N_18937);
or U20967 (N_20967,N_16970,N_19561);
or U20968 (N_20968,N_15106,N_16308);
and U20969 (N_20969,N_18991,N_16325);
xnor U20970 (N_20970,N_18417,N_19377);
or U20971 (N_20971,N_18873,N_15240);
and U20972 (N_20972,N_15468,N_17327);
nand U20973 (N_20973,N_17808,N_17740);
and U20974 (N_20974,N_18039,N_15684);
nand U20975 (N_20975,N_15632,N_16568);
nand U20976 (N_20976,N_15078,N_17476);
nand U20977 (N_20977,N_15432,N_19638);
and U20978 (N_20978,N_19434,N_18743);
or U20979 (N_20979,N_17680,N_18513);
xor U20980 (N_20980,N_18686,N_19396);
nor U20981 (N_20981,N_15831,N_15991);
nor U20982 (N_20982,N_19337,N_18436);
and U20983 (N_20983,N_15874,N_15391);
nor U20984 (N_20984,N_17148,N_19984);
and U20985 (N_20985,N_19083,N_16921);
or U20986 (N_20986,N_17674,N_16293);
and U20987 (N_20987,N_16743,N_18956);
nor U20988 (N_20988,N_19059,N_17722);
nand U20989 (N_20989,N_16939,N_16998);
xor U20990 (N_20990,N_16122,N_16771);
and U20991 (N_20991,N_19482,N_19265);
nor U20992 (N_20992,N_18857,N_18608);
nand U20993 (N_20993,N_17776,N_17282);
or U20994 (N_20994,N_17403,N_18445);
nand U20995 (N_20995,N_18561,N_17488);
nand U20996 (N_20996,N_16721,N_19015);
xnor U20997 (N_20997,N_17274,N_16177);
or U20998 (N_20998,N_19725,N_17554);
and U20999 (N_20999,N_17152,N_15865);
or U21000 (N_21000,N_15040,N_15711);
nand U21001 (N_21001,N_18168,N_18929);
nor U21002 (N_21002,N_17183,N_17803);
nand U21003 (N_21003,N_17309,N_18103);
and U21004 (N_21004,N_16282,N_18662);
nor U21005 (N_21005,N_15020,N_17292);
xor U21006 (N_21006,N_18724,N_19581);
or U21007 (N_21007,N_18381,N_16170);
and U21008 (N_21008,N_19896,N_18002);
nand U21009 (N_21009,N_17810,N_19448);
and U21010 (N_21010,N_18524,N_18993);
xor U21011 (N_21011,N_18523,N_19823);
nor U21012 (N_21012,N_17787,N_19148);
nand U21013 (N_21013,N_15692,N_19419);
xnor U21014 (N_21014,N_17487,N_15021);
nor U21015 (N_21015,N_16104,N_18279);
nor U21016 (N_21016,N_18024,N_16679);
xnor U21017 (N_21017,N_18102,N_15878);
nand U21018 (N_21018,N_16145,N_17026);
and U21019 (N_21019,N_18337,N_17575);
xnor U21020 (N_21020,N_19041,N_17472);
nor U21021 (N_21021,N_18709,N_19693);
xnor U21022 (N_21022,N_16205,N_15046);
and U21023 (N_21023,N_18280,N_16442);
xnor U21024 (N_21024,N_16156,N_18952);
nand U21025 (N_21025,N_16211,N_17662);
xnor U21026 (N_21026,N_18700,N_15324);
xnor U21027 (N_21027,N_17626,N_18178);
nand U21028 (N_21028,N_15433,N_17503);
nor U21029 (N_21029,N_17273,N_18646);
xnor U21030 (N_21030,N_16050,N_19186);
nand U21031 (N_21031,N_19088,N_18635);
and U21032 (N_21032,N_17334,N_16876);
nor U21033 (N_21033,N_15095,N_17587);
nor U21034 (N_21034,N_18838,N_18220);
xnor U21035 (N_21035,N_18166,N_18856);
nor U21036 (N_21036,N_19841,N_19302);
xor U21037 (N_21037,N_16799,N_19099);
and U21038 (N_21038,N_18841,N_16765);
xor U21039 (N_21039,N_17551,N_15779);
or U21040 (N_21040,N_18465,N_18541);
nor U21041 (N_21041,N_18309,N_18782);
nor U21042 (N_21042,N_19264,N_15600);
or U21043 (N_21043,N_17394,N_18184);
nor U21044 (N_21044,N_15099,N_16781);
or U21045 (N_21045,N_19786,N_15615);
nor U21046 (N_21046,N_16882,N_19021);
and U21047 (N_21047,N_16360,N_17763);
xnor U21048 (N_21048,N_16766,N_18812);
nor U21049 (N_21049,N_17099,N_19400);
nor U21050 (N_21050,N_15589,N_15037);
xnor U21051 (N_21051,N_18967,N_18129);
nand U21052 (N_21052,N_16037,N_17489);
or U21053 (N_21053,N_19135,N_15073);
nor U21054 (N_21054,N_16389,N_18874);
or U21055 (N_21055,N_19622,N_19542);
xor U21056 (N_21056,N_15604,N_15273);
and U21057 (N_21057,N_16681,N_17461);
nand U21058 (N_21058,N_16775,N_16906);
nor U21059 (N_21059,N_18288,N_16926);
nor U21060 (N_21060,N_15658,N_15139);
xor U21061 (N_21061,N_18272,N_16305);
or U21062 (N_21062,N_19832,N_17227);
nand U21063 (N_21063,N_19757,N_18170);
nand U21064 (N_21064,N_17930,N_19426);
or U21065 (N_21065,N_18927,N_17251);
or U21066 (N_21066,N_18553,N_15267);
xor U21067 (N_21067,N_17664,N_19042);
nand U21068 (N_21068,N_19097,N_16671);
nand U21069 (N_21069,N_17534,N_15880);
nor U21070 (N_21070,N_19365,N_19994);
xor U21071 (N_21071,N_16833,N_15035);
and U21072 (N_21072,N_15503,N_16415);
nand U21073 (N_21073,N_15795,N_18227);
nand U21074 (N_21074,N_18558,N_19410);
or U21075 (N_21075,N_16797,N_18837);
or U21076 (N_21076,N_19764,N_19727);
and U21077 (N_21077,N_17992,N_19149);
nor U21078 (N_21078,N_19324,N_15032);
or U21079 (N_21079,N_15335,N_15912);
or U21080 (N_21080,N_19905,N_18985);
nand U21081 (N_21081,N_15186,N_16024);
and U21082 (N_21082,N_16350,N_18089);
or U21083 (N_21083,N_19183,N_16368);
or U21084 (N_21084,N_15672,N_16773);
nand U21085 (N_21085,N_15063,N_18572);
nand U21086 (N_21086,N_17159,N_18082);
xnor U21087 (N_21087,N_17953,N_17558);
nand U21088 (N_21088,N_17663,N_16251);
nand U21089 (N_21089,N_15084,N_15449);
and U21090 (N_21090,N_16530,N_19288);
nand U21091 (N_21091,N_17563,N_17527);
or U21092 (N_21092,N_17440,N_17441);
nand U21093 (N_21093,N_19166,N_17724);
or U21094 (N_21094,N_17726,N_18790);
and U21095 (N_21095,N_15108,N_19457);
nand U21096 (N_21096,N_15344,N_17641);
xor U21097 (N_21097,N_16257,N_18301);
xor U21098 (N_21098,N_16522,N_16078);
and U21099 (N_21099,N_17839,N_16399);
nand U21100 (N_21100,N_15775,N_19668);
and U21101 (N_21101,N_19350,N_19671);
xor U21102 (N_21102,N_15833,N_15467);
or U21103 (N_21103,N_19891,N_17039);
and U21104 (N_21104,N_16643,N_16652);
xnor U21105 (N_21105,N_16978,N_19243);
nand U21106 (N_21106,N_18214,N_16397);
nor U21107 (N_21107,N_19389,N_17035);
or U21108 (N_21108,N_15309,N_17559);
xor U21109 (N_21109,N_17614,N_19910);
nor U21110 (N_21110,N_19256,N_19836);
nand U21111 (N_21111,N_18380,N_16825);
xor U21112 (N_21112,N_15339,N_15697);
nand U21113 (N_21113,N_19782,N_17817);
or U21114 (N_21114,N_18338,N_18905);
xor U21115 (N_21115,N_17834,N_16878);
and U21116 (N_21116,N_15041,N_15786);
xnor U21117 (N_21117,N_17074,N_16728);
or U21118 (N_21118,N_15931,N_18832);
and U21119 (N_21119,N_16689,N_15098);
and U21120 (N_21120,N_16620,N_17466);
xor U21121 (N_21121,N_18435,N_19916);
nand U21122 (N_21122,N_19204,N_18263);
xnor U21123 (N_21123,N_17108,N_19157);
nor U21124 (N_21124,N_15039,N_17252);
and U21125 (N_21125,N_17299,N_15019);
and U21126 (N_21126,N_19571,N_19201);
and U21127 (N_21127,N_17250,N_19661);
xnor U21128 (N_21128,N_16119,N_17860);
and U21129 (N_21129,N_15088,N_19209);
and U21130 (N_21130,N_16333,N_17796);
or U21131 (N_21131,N_16736,N_15009);
nand U21132 (N_21132,N_18200,N_18547);
or U21133 (N_21133,N_19213,N_16453);
or U21134 (N_21134,N_15124,N_18218);
xor U21135 (N_21135,N_18171,N_17842);
or U21136 (N_21136,N_17965,N_18639);
or U21137 (N_21137,N_15915,N_18903);
xor U21138 (N_21138,N_16989,N_18536);
xnor U21139 (N_21139,N_16786,N_18669);
xor U21140 (N_21140,N_18508,N_16440);
nor U21141 (N_21141,N_16565,N_16030);
nand U21142 (N_21142,N_18132,N_16459);
nand U21143 (N_21143,N_17443,N_18934);
xnor U21144 (N_21144,N_16412,N_18654);
or U21145 (N_21145,N_18000,N_15939);
nand U21146 (N_21146,N_17199,N_15380);
nor U21147 (N_21147,N_16541,N_16209);
nor U21148 (N_21148,N_19830,N_15153);
or U21149 (N_21149,N_19178,N_16850);
and U21150 (N_21150,N_17906,N_16197);
nor U21151 (N_21151,N_15891,N_15643);
nand U21152 (N_21152,N_18341,N_17182);
nand U21153 (N_21153,N_16218,N_18765);
or U21154 (N_21154,N_16090,N_17386);
or U21155 (N_21155,N_15969,N_16995);
nand U21156 (N_21156,N_17326,N_19467);
nand U21157 (N_21157,N_15904,N_18990);
or U21158 (N_21158,N_18658,N_17156);
xnor U21159 (N_21159,N_16937,N_19237);
and U21160 (N_21160,N_19517,N_19022);
and U21161 (N_21161,N_17505,N_15406);
and U21162 (N_21162,N_15164,N_19124);
and U21163 (N_21163,N_18474,N_17350);
nor U21164 (N_21164,N_19719,N_15246);
and U21165 (N_21165,N_16592,N_18364);
or U21166 (N_21166,N_19368,N_19937);
and U21167 (N_21167,N_19478,N_16059);
nor U21168 (N_21168,N_17176,N_18312);
and U21169 (N_21169,N_17109,N_19878);
nand U21170 (N_21170,N_19146,N_18404);
nor U21171 (N_21171,N_17141,N_19326);
or U21172 (N_21172,N_16447,N_19310);
and U21173 (N_21173,N_19339,N_16718);
nand U21174 (N_21174,N_19170,N_18557);
nand U21175 (N_21175,N_15717,N_16267);
or U21176 (N_21176,N_15556,N_17512);
or U21177 (N_21177,N_15882,N_18925);
nand U21178 (N_21178,N_19526,N_18326);
or U21179 (N_21179,N_16058,N_17866);
or U21180 (N_21180,N_18421,N_17448);
nand U21181 (N_21181,N_18680,N_15617);
nand U21182 (N_21182,N_16446,N_15591);
nand U21183 (N_21183,N_18154,N_15172);
or U21184 (N_21184,N_18797,N_16572);
nand U21185 (N_21185,N_15109,N_17742);
and U21186 (N_21186,N_19536,N_18690);
and U21187 (N_21187,N_15976,N_16682);
nand U21188 (N_21188,N_17097,N_17540);
nand U21189 (N_21189,N_18514,N_15206);
xnor U21190 (N_21190,N_17091,N_17272);
and U21191 (N_21191,N_16897,N_18109);
nand U21192 (N_21192,N_16966,N_18451);
nand U21193 (N_21193,N_19039,N_16872);
or U21194 (N_21194,N_15647,N_17884);
nand U21195 (N_21195,N_16162,N_19316);
nand U21196 (N_21196,N_19805,N_15791);
and U21197 (N_21197,N_15141,N_15785);
nand U21198 (N_21198,N_18774,N_16498);
nand U21199 (N_21199,N_15733,N_18554);
or U21200 (N_21200,N_16043,N_15288);
xor U21201 (N_21201,N_17064,N_15157);
nor U21202 (N_21202,N_19743,N_16800);
or U21203 (N_21203,N_19092,N_19920);
nor U21204 (N_21204,N_16821,N_17861);
or U21205 (N_21205,N_19603,N_19395);
nor U21206 (N_21206,N_16856,N_17853);
or U21207 (N_21207,N_17553,N_19986);
nand U21208 (N_21208,N_15014,N_18897);
or U21209 (N_21209,N_19076,N_16735);
nor U21210 (N_21210,N_16087,N_17847);
or U21211 (N_21211,N_19912,N_15829);
nor U21212 (N_21212,N_17138,N_19930);
nand U21213 (N_21213,N_16358,N_15062);
nor U21214 (N_21214,N_16824,N_18834);
nor U21215 (N_21215,N_19964,N_17574);
nor U21216 (N_21216,N_15637,N_17765);
xor U21217 (N_21217,N_18933,N_15735);
and U21218 (N_21218,N_19160,N_19499);
nor U21219 (N_21219,N_17928,N_15905);
xnor U21220 (N_21220,N_19819,N_17260);
nand U21221 (N_21221,N_16845,N_18238);
nor U21222 (N_21222,N_16158,N_18556);
nor U21223 (N_21223,N_16615,N_18736);
or U21224 (N_21224,N_19435,N_16675);
xor U21225 (N_21225,N_16342,N_16990);
and U21226 (N_21226,N_18480,N_17276);
nand U21227 (N_21227,N_16612,N_19048);
nor U21228 (N_21228,N_16593,N_18876);
and U21229 (N_21229,N_18613,N_19304);
nand U21230 (N_21230,N_19583,N_15176);
or U21231 (N_21231,N_18057,N_16934);
or U21232 (N_21232,N_15802,N_17295);
xor U21233 (N_21233,N_19067,N_16452);
xor U21234 (N_21234,N_17682,N_17628);
nand U21235 (N_21235,N_19973,N_17423);
xor U21236 (N_21236,N_16336,N_16852);
and U21237 (N_21237,N_18877,N_18752);
and U21238 (N_21238,N_16678,N_18294);
or U21239 (N_21239,N_16994,N_17733);
nand U21240 (N_21240,N_16461,N_16131);
or U21241 (N_21241,N_19248,N_16300);
nor U21242 (N_21242,N_16901,N_18244);
or U21243 (N_21243,N_17770,N_15516);
xnor U21244 (N_21244,N_19714,N_18007);
and U21245 (N_21245,N_15598,N_15057);
xnor U21246 (N_21246,N_15358,N_15007);
and U21247 (N_21247,N_17541,N_16366);
or U21248 (N_21248,N_18921,N_15852);
or U21249 (N_21249,N_15642,N_18586);
or U21250 (N_21250,N_19374,N_17608);
nor U21251 (N_21251,N_15848,N_19352);
xnor U21252 (N_21252,N_17526,N_18896);
nor U21253 (N_21253,N_19995,N_15780);
xnor U21254 (N_21254,N_17154,N_16772);
and U21255 (N_21255,N_17398,N_19211);
nand U21256 (N_21256,N_16685,N_19925);
xnor U21257 (N_21257,N_19538,N_19442);
nor U21258 (N_21258,N_16183,N_18511);
and U21259 (N_21259,N_17835,N_17388);
or U21260 (N_21260,N_19987,N_19894);
and U21261 (N_21261,N_15445,N_18449);
or U21262 (N_21262,N_17033,N_17175);
nor U21263 (N_21263,N_16696,N_16532);
and U21264 (N_21264,N_16495,N_17463);
and U21265 (N_21265,N_19778,N_18359);
nor U21266 (N_21266,N_16986,N_15303);
and U21267 (N_21267,N_17944,N_18412);
xnor U21268 (N_21268,N_15282,N_17223);
or U21269 (N_21269,N_15893,N_16955);
or U21270 (N_21270,N_15553,N_17076);
nand U21271 (N_21271,N_17056,N_15497);
and U21272 (N_21272,N_17822,N_19642);
xor U21273 (N_21273,N_17831,N_18169);
and U21274 (N_21274,N_17418,N_16534);
and U21275 (N_21275,N_18183,N_19756);
or U21276 (N_21276,N_16749,N_16942);
xor U21277 (N_21277,N_16488,N_15620);
or U21278 (N_21278,N_15093,N_19579);
or U21279 (N_21279,N_17792,N_17228);
and U21280 (N_21280,N_17499,N_16885);
or U21281 (N_21281,N_19670,N_18010);
nor U21282 (N_21282,N_15362,N_19874);
and U21283 (N_21283,N_16793,N_16666);
nor U21284 (N_21284,N_16472,N_18591);
nor U21285 (N_21285,N_18245,N_19588);
nand U21286 (N_21286,N_19513,N_15601);
nand U21287 (N_21287,N_16095,N_15743);
nand U21288 (N_21288,N_17882,N_18515);
or U21289 (N_21289,N_17507,N_19498);
and U21290 (N_21290,N_19722,N_15669);
or U21291 (N_21291,N_18468,N_18075);
xnor U21292 (N_21292,N_19474,N_16684);
nand U21293 (N_21293,N_18064,N_16118);
and U21294 (N_21294,N_17661,N_15776);
nor U21295 (N_21295,N_19718,N_16672);
xnor U21296 (N_21296,N_18135,N_17938);
nand U21297 (N_21297,N_15533,N_16477);
and U21298 (N_21298,N_19210,N_15704);
xnor U21299 (N_21299,N_18850,N_17665);
and U21300 (N_21300,N_17719,N_16413);
nor U21301 (N_21301,N_18355,N_17325);
or U21302 (N_21302,N_19463,N_15768);
nand U21303 (N_21303,N_19882,N_19876);
nor U21304 (N_21304,N_15384,N_18811);
nand U21305 (N_21305,N_15005,N_17101);
nand U21306 (N_21306,N_16060,N_15222);
xor U21307 (N_21307,N_17772,N_17562);
and U21308 (N_21308,N_19917,N_16070);
xor U21309 (N_21309,N_18555,N_17857);
xor U21310 (N_21310,N_18574,N_15143);
or U21311 (N_21311,N_16900,N_17349);
xnor U21312 (N_21312,N_16105,N_18111);
and U21313 (N_21313,N_15507,N_15696);
xor U21314 (N_21314,N_19461,N_16153);
xor U21315 (N_21315,N_19793,N_17224);
nor U21316 (N_21316,N_18235,N_16294);
or U21317 (N_21317,N_19225,N_16421);
nor U21318 (N_21318,N_15196,N_19333);
nand U21319 (N_21319,N_19852,N_16152);
nor U21320 (N_21320,N_17451,N_17289);
and U21321 (N_21321,N_17264,N_15954);
nand U21322 (N_21322,N_19548,N_19431);
and U21323 (N_21323,N_15723,N_19050);
nand U21324 (N_21324,N_18180,N_16891);
xor U21325 (N_21325,N_15238,N_15051);
xor U21326 (N_21326,N_15022,N_15180);
and U21327 (N_21327,N_16958,N_19278);
or U21328 (N_21328,N_17529,N_15430);
xnor U21329 (N_21329,N_16988,N_17686);
nand U21330 (N_21330,N_17700,N_16917);
xor U21331 (N_21331,N_19032,N_15466);
nor U21332 (N_21332,N_16759,N_19975);
xnor U21333 (N_21333,N_16414,N_16019);
xor U21334 (N_21334,N_18330,N_17053);
and U21335 (N_21335,N_16371,N_15524);
nand U21336 (N_21336,N_16303,N_18226);
or U21337 (N_21337,N_18842,N_17581);
and U21338 (N_21338,N_16578,N_18773);
nor U21339 (N_21339,N_15670,N_18519);
xor U21340 (N_21340,N_18005,N_16193);
nand U21341 (N_21341,N_15561,N_19858);
nor U21342 (N_21342,N_17090,N_18716);
nor U21343 (N_21343,N_16561,N_16138);
nand U21344 (N_21344,N_18062,N_19963);
and U21345 (N_21345,N_16427,N_19271);
xor U21346 (N_21346,N_15703,N_17677);
or U21347 (N_21347,N_15975,N_16583);
nand U21348 (N_21348,N_18446,N_18219);
or U21349 (N_21349,N_18504,N_16609);
or U21350 (N_21350,N_17736,N_17535);
and U21351 (N_21351,N_16904,N_18965);
xor U21352 (N_21352,N_19167,N_15750);
xor U21353 (N_21353,N_16858,N_16284);
and U21354 (N_21354,N_18190,N_17036);
and U21355 (N_21355,N_16899,N_18795);
or U21356 (N_21356,N_18313,N_19198);
xor U21357 (N_21357,N_19811,N_18281);
xnor U21358 (N_21358,N_17236,N_19857);
nand U21359 (N_21359,N_15103,N_19759);
nand U21360 (N_21360,N_16167,N_19047);
and U21361 (N_21361,N_19164,N_17445);
and U21362 (N_21362,N_16147,N_19082);
xor U21363 (N_21363,N_17302,N_16173);
and U21364 (N_21364,N_19692,N_17694);
and U21365 (N_21365,N_15327,N_16518);
or U21366 (N_21366,N_19104,N_17741);
nor U21367 (N_21367,N_19207,N_17029);
and U21368 (N_21368,N_17267,N_16912);
and U21369 (N_21369,N_17100,N_15232);
xnor U21370 (N_21370,N_17632,N_16185);
nand U21371 (N_21371,N_17758,N_15219);
or U21372 (N_21372,N_17561,N_17846);
and U21373 (N_21373,N_15788,N_19066);
nor U21374 (N_21374,N_18221,N_19990);
nand U21375 (N_21375,N_15165,N_19228);
and U21376 (N_21376,N_17655,N_16869);
nor U21377 (N_21377,N_15145,N_18377);
or U21378 (N_21378,N_17140,N_18127);
and U21379 (N_21379,N_17490,N_17610);
xnor U21380 (N_21380,N_17607,N_15972);
xor U21381 (N_21381,N_16594,N_18050);
nor U21382 (N_21382,N_16202,N_17107);
and U21383 (N_21383,N_19095,N_19259);
or U21384 (N_21384,N_19266,N_18595);
nand U21385 (N_21385,N_15385,N_17693);
nor U21386 (N_21386,N_19586,N_15519);
or U21387 (N_21387,N_17284,N_17936);
or U21388 (N_21388,N_16549,N_15849);
and U21389 (N_21389,N_15476,N_18291);
and U21390 (N_21390,N_15231,N_18503);
nand U21391 (N_21391,N_17475,N_16449);
and U21392 (N_21392,N_19965,N_17406);
nand U21393 (N_21393,N_15372,N_19356);
and U21394 (N_21394,N_16525,N_15707);
or U21395 (N_21395,N_16482,N_16552);
and U21396 (N_21396,N_19475,N_19038);
and U21397 (N_21397,N_15114,N_15122);
nor U21398 (N_21398,N_16315,N_19690);
nand U21399 (N_21399,N_16020,N_15193);
or U21400 (N_21400,N_19306,N_15527);
or U21401 (N_21401,N_19507,N_15822);
and U21402 (N_21402,N_16836,N_19816);
or U21403 (N_21403,N_18681,N_19931);
and U21404 (N_21404,N_18573,N_17017);
and U21405 (N_21405,N_15951,N_17382);
xnor U21406 (N_21406,N_17283,N_17819);
nor U21407 (N_21407,N_18745,N_19127);
and U21408 (N_21408,N_18784,N_16404);
nor U21409 (N_21409,N_16429,N_17710);
nor U21410 (N_21410,N_19886,N_17384);
nor U21411 (N_21411,N_15161,N_18899);
xor U21412 (N_21412,N_15909,N_18563);
xor U21413 (N_21413,N_15102,N_17676);
xor U21414 (N_21414,N_15960,N_17266);
nor U21415 (N_21415,N_16529,N_19114);
and U21416 (N_21416,N_16963,N_19416);
and U21417 (N_21417,N_19224,N_19943);
nand U21418 (N_21418,N_15456,N_19651);
or U21419 (N_21419,N_15459,N_19331);
nor U21420 (N_21420,N_15069,N_16881);
or U21421 (N_21421,N_19568,N_18974);
or U21422 (N_21422,N_17970,N_16015);
xor U21423 (N_21423,N_17112,N_18786);
nor U21424 (N_21424,N_18375,N_19558);
or U21425 (N_21425,N_16259,N_19317);
nor U21426 (N_21426,N_16061,N_18114);
nor U21427 (N_21427,N_16388,N_18498);
xnor U21428 (N_21428,N_16639,N_18957);
xnor U21429 (N_21429,N_17975,N_18791);
nand U21430 (N_21430,N_17303,N_19016);
nand U21431 (N_21431,N_19241,N_15592);
or U21432 (N_21432,N_18886,N_16992);
and U21433 (N_21433,N_16871,N_17328);
and U21434 (N_21434,N_15753,N_15382);
or U21435 (N_21435,N_18727,N_19794);
and U21436 (N_21436,N_16941,N_17501);
or U21437 (N_21437,N_16079,N_19208);
xor U21438 (N_21438,N_15935,N_19751);
xnor U21439 (N_21439,N_18549,N_17225);
and U21440 (N_21440,N_19974,N_18810);
xnor U21441 (N_21441,N_19527,N_19172);
or U21442 (N_21442,N_18623,N_17695);
xnor U21443 (N_21443,N_19134,N_16226);
or U21444 (N_21444,N_17871,N_15045);
or U21445 (N_21445,N_18587,N_16032);
nand U21446 (N_21446,N_16809,N_17474);
xor U21447 (N_21447,N_15528,N_15547);
or U21448 (N_21448,N_18121,N_19753);
nand U21449 (N_21449,N_19710,N_18559);
nor U21450 (N_21450,N_19962,N_18798);
or U21451 (N_21451,N_15911,N_19817);
and U21452 (N_21452,N_19506,N_17764);
xor U21453 (N_21453,N_19454,N_18277);
nor U21454 (N_21454,N_16859,N_19745);
or U21455 (N_21455,N_15326,N_18598);
nor U21456 (N_21456,N_15599,N_17197);
and U21457 (N_21457,N_17976,N_17902);
nor U21458 (N_21458,N_15170,N_16960);
xor U21459 (N_21459,N_16815,N_16748);
or U21460 (N_21460,N_19197,N_17004);
or U21461 (N_21461,N_18476,N_16409);
and U21462 (N_21462,N_19179,N_18255);
xnor U21463 (N_21463,N_18726,N_15805);
xnor U21464 (N_21464,N_15422,N_17119);
xnor U21465 (N_21465,N_17903,N_16287);
or U21466 (N_21466,N_19388,N_18247);
and U21467 (N_21467,N_17215,N_16528);
nor U21468 (N_21468,N_18624,N_15252);
nor U21469 (N_21469,N_15755,N_16722);
nand U21470 (N_21470,N_16712,N_17121);
and U21471 (N_21471,N_18807,N_17161);
and U21472 (N_21472,N_18251,N_16106);
and U21473 (N_21473,N_19370,N_18578);
and U21474 (N_21474,N_15361,N_16820);
nand U21475 (N_21475,N_15147,N_19093);
xor U21476 (N_21476,N_17933,N_19940);
nor U21477 (N_21477,N_17956,N_16445);
nand U21478 (N_21478,N_19696,N_19885);
xnor U21479 (N_21479,N_16502,N_18399);
or U21480 (N_21480,N_19020,N_15654);
and U21481 (N_21481,N_15318,N_15557);
or U21482 (N_21482,N_19932,N_19398);
and U21483 (N_21483,N_18528,N_17027);
nand U21484 (N_21484,N_19330,N_19154);
and U21485 (N_21485,N_16332,N_15988);
xnor U21486 (N_21486,N_16465,N_15811);
nor U21487 (N_21487,N_15720,N_17449);
or U21488 (N_21488,N_15472,N_18187);
xnor U21489 (N_21489,N_19597,N_19784);
or U21490 (N_21490,N_16382,N_17761);
nand U21491 (N_21491,N_16065,N_19444);
and U21492 (N_21492,N_15463,N_15353);
nand U21493 (N_21493,N_18840,N_15932);
or U21494 (N_21494,N_19079,N_19030);
nor U21495 (N_21495,N_15094,N_16602);
and U21496 (N_21496,N_18151,N_15836);
or U21497 (N_21497,N_18395,N_15685);
nor U21498 (N_21498,N_16093,N_17576);
xnor U21499 (N_21499,N_19169,N_16903);
xnor U21500 (N_21500,N_17308,N_16560);
and U21501 (N_21501,N_18590,N_18334);
nor U21502 (N_21502,N_19602,N_18981);
xor U21503 (N_21503,N_19091,N_17883);
xnor U21504 (N_21504,N_18414,N_19815);
xnor U21505 (N_21505,N_16693,N_17137);
and U21506 (N_21506,N_16141,N_16394);
nor U21507 (N_21507,N_15570,N_15223);
or U21508 (N_21508,N_17732,N_19702);
xnor U21509 (N_21509,N_19101,N_18442);
xor U21510 (N_21510,N_17544,N_16289);
nand U21511 (N_21511,N_16416,N_17072);
nand U21512 (N_21512,N_18808,N_15169);
or U21513 (N_21513,N_18495,N_18325);
or U21514 (N_21514,N_19948,N_16474);
or U21515 (N_21515,N_17067,N_16034);
or U21516 (N_21516,N_17672,N_15003);
nand U21517 (N_21517,N_17400,N_16435);
and U21518 (N_21518,N_18516,N_18482);
or U21519 (N_21519,N_18884,N_16384);
and U21520 (N_21520,N_16179,N_15450);
or U21521 (N_21521,N_16513,N_17821);
or U21522 (N_21522,N_15462,N_19550);
nand U21523 (N_21523,N_15798,N_18983);
and U21524 (N_21524,N_18829,N_15922);
and U21525 (N_21525,N_16313,N_17789);
and U21526 (N_21526,N_15652,N_18054);
nor U21527 (N_21527,N_19629,N_16254);
xnor U21528 (N_21528,N_17170,N_16944);
nor U21529 (N_21529,N_17771,N_17688);
xor U21530 (N_21530,N_16144,N_17569);
nor U21531 (N_21531,N_19998,N_17528);
or U21532 (N_21532,N_19945,N_19496);
or U21533 (N_21533,N_18621,N_16444);
or U21534 (N_21534,N_16631,N_16890);
xnor U21535 (N_21535,N_19748,N_18703);
xor U21536 (N_21536,N_19459,N_17856);
and U21537 (N_21537,N_18951,N_15930);
nand U21538 (N_21538,N_18393,N_15356);
and U21539 (N_21539,N_18292,N_15265);
xor U21540 (N_21540,N_17185,N_17248);
xor U21541 (N_21541,N_19145,N_17752);
nor U21542 (N_21542,N_18542,N_17983);
or U21543 (N_21543,N_18431,N_18432);
nand U21544 (N_21544,N_18455,N_15650);
xor U21545 (N_21545,N_17548,N_17707);
nand U21546 (N_21546,N_15090,N_15614);
xnor U21547 (N_21547,N_15080,N_18149);
nand U21548 (N_21548,N_18152,N_19407);
xor U21549 (N_21549,N_17980,N_15424);
or U21550 (N_21550,N_18964,N_15824);
xnor U21551 (N_21551,N_16959,N_15651);
xnor U21552 (N_21552,N_19185,N_18425);
xor U21553 (N_21553,N_17318,N_15917);
or U21554 (N_21554,N_17484,N_19102);
or U21555 (N_21555,N_19218,N_15588);
xnor U21556 (N_21556,N_17142,N_16981);
xnor U21557 (N_21557,N_15201,N_16143);
xnor U21558 (N_21558,N_19007,N_15839);
and U21559 (N_21559,N_19433,N_18885);
or U21560 (N_21560,N_15135,N_19223);
nand U21561 (N_21561,N_18343,N_16383);
nand U21562 (N_21562,N_19284,N_16441);
nand U21563 (N_21563,N_19060,N_17753);
or U21564 (N_21564,N_16827,N_17773);
and U21565 (N_21565,N_18534,N_15832);
nand U21566 (N_21566,N_15234,N_17816);
and U21567 (N_21567,N_16764,N_18777);
nor U21568 (N_21568,N_16946,N_17462);
and U21569 (N_21569,N_17966,N_16925);
xnor U21570 (N_21570,N_16751,N_19935);
xor U21571 (N_21571,N_15853,N_19904);
or U21572 (N_21572,N_19440,N_16025);
nor U21573 (N_21573,N_19519,N_19383);
nand U21574 (N_21574,N_16984,N_18936);
and U21575 (N_21575,N_19865,N_17482);
nor U21576 (N_21576,N_17297,N_18131);
nor U21577 (N_21577,N_15163,N_17044);
or U21578 (N_21578,N_17492,N_16476);
nor U21579 (N_21579,N_15899,N_18475);
nand U21580 (N_21580,N_16625,N_19500);
xor U21581 (N_21581,N_16887,N_15892);
nor U21582 (N_21582,N_16972,N_16199);
and U21583 (N_21583,N_18004,N_19859);
or U21584 (N_21584,N_19153,N_17517);
xor U21585 (N_21585,N_16710,N_19535);
nor U21586 (N_21586,N_16486,N_16686);
nand U21587 (N_21587,N_18824,N_19391);
nand U21588 (N_21588,N_17735,N_17008);
nor U21589 (N_21589,N_16165,N_19013);
and U21590 (N_21590,N_18844,N_16484);
xor U21591 (N_21591,N_15801,N_16281);
or U21592 (N_21592,N_15659,N_15585);
nand U21593 (N_21593,N_16052,N_19645);
and U21594 (N_21594,N_18970,N_17634);
nand U21595 (N_21595,N_16563,N_15739);
xnor U21596 (N_21596,N_16697,N_16373);
nor U21597 (N_21597,N_16929,N_18097);
or U21598 (N_21598,N_17908,N_18860);
xnor U21599 (N_21599,N_16086,N_17525);
xor U21600 (N_21600,N_16551,N_15125);
and U21601 (N_21601,N_19861,N_15200);
xnor U21602 (N_21602,N_16424,N_16683);
xnor U21603 (N_21603,N_17355,N_15575);
or U21604 (N_21604,N_15495,N_17337);
or U21605 (N_21605,N_16364,N_16531);
xnor U21606 (N_21606,N_18086,N_18806);
xor U21607 (N_21607,N_18110,N_15154);
or U21608 (N_21608,N_17191,N_19869);
xor U21609 (N_21609,N_18047,N_18537);
nand U21610 (N_21610,N_16216,N_17889);
nand U21611 (N_21611,N_19246,N_19780);
or U21612 (N_21612,N_17603,N_19863);
nor U21613 (N_21613,N_17401,N_18182);
xor U21614 (N_21614,N_17301,N_18894);
nand U21615 (N_21615,N_19432,N_16691);
xor U21616 (N_21616,N_15680,N_17909);
xor U21617 (N_21617,N_18307,N_15936);
nor U21618 (N_21618,N_18327,N_18036);
and U21619 (N_21619,N_19704,N_15981);
and U21620 (N_21620,N_15777,N_16464);
xor U21621 (N_21621,N_18368,N_17913);
or U21622 (N_21622,N_18958,N_16062);
and U21623 (N_21623,N_18879,N_17087);
xor U21624 (N_21624,N_18543,N_16774);
nand U21625 (N_21625,N_19980,N_17891);
nor U21626 (N_21626,N_15312,N_15846);
or U21627 (N_21627,N_16595,N_19619);
nand U21628 (N_21628,N_17126,N_19676);
nor U21629 (N_21629,N_16732,N_15649);
xor U21630 (N_21630,N_16954,N_16741);
nand U21631 (N_21631,N_18738,N_17397);
and U21632 (N_21632,N_19924,N_16433);
and U21633 (N_21633,N_17666,N_17166);
xor U21634 (N_21634,N_16641,N_17757);
xnor U21635 (N_21635,N_17294,N_16451);
nor U21636 (N_21636,N_15896,N_18348);
nand U21637 (N_21637,N_19944,N_15940);
nor U21638 (N_21638,N_16114,N_19976);
and U21639 (N_21639,N_16857,N_19989);
nor U21640 (N_21640,N_17673,N_19397);
nor U21641 (N_21641,N_16245,N_19926);
or U21642 (N_21642,N_15225,N_17885);
and U21643 (N_21643,N_17049,N_17439);
or U21644 (N_21644,N_19598,N_18507);
nand U21645 (N_21645,N_16626,N_18742);
and U21646 (N_21646,N_15409,N_15074);
xor U21647 (N_21647,N_15744,N_17685);
nor U21648 (N_21648,N_15412,N_18702);
or U21649 (N_21649,N_16648,N_17257);
nand U21650 (N_21650,N_17769,N_17728);
nor U21651 (N_21651,N_16127,N_16973);
nor U21652 (N_21652,N_19490,N_18038);
nand U21653 (N_21653,N_16107,N_19582);
or U21654 (N_21654,N_16374,N_19730);
or U21655 (N_21655,N_17730,N_16980);
xor U21656 (N_21656,N_18285,N_17830);
and U21657 (N_21657,N_15434,N_17205);
or U21658 (N_21658,N_19658,N_15389);
and U21659 (N_21659,N_18207,N_19140);
nand U21660 (N_21660,N_19412,N_16194);
xor U21661 (N_21661,N_15473,N_16450);
and U21662 (N_21662,N_17019,N_17057);
xnor U21663 (N_21663,N_18614,N_19486);
nand U21664 (N_21664,N_16724,N_15687);
or U21665 (N_21665,N_19075,N_17179);
nor U21666 (N_21666,N_19152,N_17155);
or U21667 (N_21667,N_19808,N_17255);
or U21668 (N_21668,N_15919,N_16082);
xnor U21669 (N_21669,N_19453,N_19635);
or U21670 (N_21670,N_16016,N_19184);
xnor U21671 (N_21671,N_15188,N_18972);
nand U21672 (N_21672,N_18212,N_15821);
nor U21673 (N_21673,N_17456,N_16080);
or U21674 (N_21674,N_17310,N_18048);
nor U21675 (N_21675,N_16788,N_16089);
xnor U21676 (N_21676,N_16355,N_18778);
and U21677 (N_21677,N_16263,N_19051);
nor U21678 (N_21678,N_15532,N_16419);
and U21679 (N_21679,N_19913,N_17920);
xnor U21680 (N_21680,N_18138,N_19681);
or U21681 (N_21681,N_16250,N_19023);
and U21682 (N_21682,N_19029,N_18058);
or U21683 (N_21683,N_16591,N_17921);
and U21684 (N_21684,N_16582,N_18939);
and U21685 (N_21685,N_18350,N_18962);
nand U21686 (N_21686,N_17675,N_16747);
nand U21687 (N_21687,N_19950,N_17697);
and U21688 (N_21688,N_17464,N_16454);
xor U21689 (N_21689,N_19837,N_19685);
nand U21690 (N_21690,N_17358,N_16239);
nand U21691 (N_21691,N_15149,N_17196);
xor U21692 (N_21692,N_17437,N_17599);
xor U21693 (N_21693,N_16599,N_19677);
and U21694 (N_21694,N_15258,N_15217);
nand U21695 (N_21695,N_15113,N_18085);
or U21696 (N_21696,N_18373,N_17271);
nand U21697 (N_21697,N_15515,N_18073);
nor U21698 (N_21698,N_18426,N_19477);
xor U21699 (N_21699,N_16677,N_16275);
and U21700 (N_21700,N_18907,N_15044);
and U21701 (N_21701,N_15167,N_17788);
xor U21702 (N_21702,N_19408,N_16969);
nand U21703 (N_21703,N_16976,N_18415);
nor U21704 (N_21704,N_18458,N_15331);
xnor U21705 (N_21705,N_16651,N_19509);
nand U21706 (N_21706,N_18789,N_18336);
xor U21707 (N_21707,N_17979,N_18349);
nand U21708 (N_21708,N_18201,N_16731);
and U21709 (N_21709,N_19520,N_16157);
nor U21710 (N_21710,N_16040,N_18232);
nor U21711 (N_21711,N_18046,N_19641);
or U21712 (N_21712,N_17351,N_15555);
and U21713 (N_21713,N_16527,N_16407);
and U21714 (N_21714,N_18706,N_17015);
xor U21715 (N_21715,N_15989,N_18898);
nor U21716 (N_21716,N_15416,N_17007);
xor U21717 (N_21717,N_17945,N_17955);
or U21718 (N_21718,N_15441,N_18344);
xor U21719 (N_21719,N_15097,N_15435);
and U21720 (N_21720,N_18589,N_19576);
nor U21721 (N_21721,N_15215,N_17993);
or U21722 (N_21722,N_18164,N_16705);
and U21723 (N_21723,N_16063,N_16709);
xor U21724 (N_21724,N_16894,N_17195);
nand U21725 (N_21725,N_19360,N_15656);
and U21726 (N_21726,N_17940,N_17162);
or U21727 (N_21727,N_18208,N_16823);
nor U21728 (N_21728,N_19061,N_16715);
and U21729 (N_21729,N_18027,N_18760);
or U21730 (N_21730,N_15769,N_19287);
or U21731 (N_21731,N_17972,N_18816);
nor U21732 (N_21732,N_18424,N_17048);
or U21733 (N_21733,N_16961,N_19359);
nand U21734 (N_21734,N_18984,N_17059);
or U21735 (N_21735,N_19485,N_19848);
and U21736 (N_21736,N_18517,N_18801);
nand U21737 (N_21737,N_16847,N_19652);
and U21738 (N_21738,N_15773,N_19234);
and U21739 (N_21739,N_16010,N_18820);
and U21740 (N_21740,N_15513,N_16473);
nor U21741 (N_21741,N_19249,N_16166);
xor U21742 (N_21742,N_19098,N_17922);
or U21743 (N_21743,N_15927,N_19788);
nand U21744 (N_21744,N_17206,N_17782);
or U21745 (N_21745,N_15946,N_17174);
nor U21746 (N_21746,N_16777,N_19907);
nor U21747 (N_21747,N_15461,N_17258);
or U21748 (N_21748,N_19393,N_15767);
nor U21749 (N_21749,N_18189,N_16314);
nor U21750 (N_21750,N_16410,N_15691);
nand U21751 (N_21751,N_16425,N_15337);
or U21752 (N_21752,N_15610,N_19451);
xnor U21753 (N_21753,N_18733,N_18160);
and U21754 (N_21754,N_18787,N_16628);
nor U21755 (N_21755,N_18262,N_15740);
or U21756 (N_21756,N_19362,N_19510);
and U21757 (N_21757,N_17186,N_17407);
nor U21758 (N_21758,N_17767,N_18248);
and U21759 (N_21759,N_16430,N_15060);
and U21760 (N_21760,N_19872,N_16225);
or U21761 (N_21761,N_17986,N_19219);
nor U21762 (N_21762,N_15364,N_17734);
xor U21763 (N_21763,N_17169,N_15204);
and U21764 (N_21764,N_16543,N_19458);
nand U21765 (N_21765,N_19720,N_15194);
and U21766 (N_21766,N_18403,N_15929);
xnor U21767 (N_21767,N_16761,N_18278);
nand U21768 (N_21768,N_16571,N_16750);
xor U21769 (N_21769,N_18321,N_15871);
nor U21770 (N_21770,N_19487,N_15042);
nor U21771 (N_21771,N_18562,N_18211);
nand U21772 (N_21772,N_17633,N_18612);
xnor U21773 (N_21773,N_18210,N_18749);
xnor U21774 (N_21774,N_17425,N_19846);
and U21775 (N_21775,N_18757,N_16579);
nor U21776 (N_21776,N_15048,N_16711);
nand U21777 (N_21777,N_17890,N_17725);
and U21778 (N_21778,N_15792,N_17478);
and U21779 (N_21779,N_19643,N_19261);
xor U21780 (N_21780,N_18770,N_17959);
and U21781 (N_21781,N_18191,N_18422);
nor U21782 (N_21782,N_16195,N_15151);
xnor U21783 (N_21783,N_19052,N_18484);
and U21784 (N_21784,N_18605,N_18071);
nor U21785 (N_21785,N_15890,N_17065);
or U21786 (N_21786,N_19282,N_19559);
and U21787 (N_21787,N_17422,N_17618);
nor U21788 (N_21788,N_18687,N_16826);
xnor U21789 (N_21789,N_15957,N_17336);
xnor U21790 (N_21790,N_16252,N_19729);
or U21791 (N_21791,N_18052,N_16664);
nand U21792 (N_21792,N_19567,N_15117);
and U21793 (N_21793,N_15228,N_16047);
or U21794 (N_21794,N_18029,N_19955);
and U21795 (N_21795,N_17016,N_19732);
or U21796 (N_21796,N_18762,N_15974);
xnor U21797 (N_21797,N_17335,N_16754);
or U21798 (N_21798,N_18799,N_17647);
nor U21799 (N_21799,N_18652,N_17348);
nor U21800 (N_21800,N_19161,N_17209);
and U21801 (N_21801,N_16883,N_16379);
and U21802 (N_21802,N_15440,N_17184);
and U21803 (N_21803,N_17780,N_17450);
nor U21804 (N_21804,N_15860,N_16622);
and U21805 (N_21805,N_16378,N_18788);
or U21806 (N_21806,N_18345,N_15198);
xnor U21807 (N_21807,N_18140,N_16375);
nand U21808 (N_21808,N_15202,N_16206);
or U21809 (N_21809,N_15854,N_16838);
and U21810 (N_21810,N_15454,N_15371);
xnor U21811 (N_21811,N_18755,N_16649);
nor U21812 (N_21812,N_19689,N_18827);
xnor U21813 (N_21813,N_16938,N_17591);
nor U21814 (N_21814,N_19760,N_19466);
and U21815 (N_21815,N_15269,N_16108);
nand U21816 (N_21816,N_16607,N_18405);
xnor U21817 (N_21817,N_19818,N_16295);
and U21818 (N_21818,N_16967,N_19279);
xnor U21819 (N_21819,N_18615,N_18592);
or U21820 (N_21820,N_19100,N_19103);
nand U21821 (N_21821,N_19010,N_19334);
nand U21822 (N_21822,N_15968,N_15174);
nor U21823 (N_21823,N_17969,N_15130);
nand U21824 (N_21824,N_19202,N_17611);
nor U21825 (N_21825,N_17498,N_17651);
or U21826 (N_21826,N_19533,N_19781);
xor U21827 (N_21827,N_15428,N_15321);
and U21828 (N_21828,N_16707,N_19390);
and U21829 (N_21829,N_16737,N_19363);
and U21830 (N_21830,N_16690,N_19684);
xor U21831 (N_21831,N_16129,N_17438);
nand U21832 (N_21832,N_15178,N_15027);
nand U21833 (N_21833,N_16307,N_15971);
or U21834 (N_21834,N_19600,N_15675);
nor U21835 (N_21835,N_17201,N_15367);
nor U21836 (N_21836,N_15270,N_19890);
or U21837 (N_21837,N_15724,N_18420);
and U21838 (N_21838,N_16215,N_15823);
nor U21839 (N_21839,N_18665,N_15479);
nand U21840 (N_21840,N_15192,N_18035);
xor U21841 (N_21841,N_16345,N_16489);
xor U21842 (N_21842,N_19728,N_18628);
nor U21843 (N_21843,N_15800,N_15872);
or U21844 (N_21844,N_16168,N_16843);
and U21845 (N_21845,N_17929,N_16523);
and U21846 (N_21846,N_19277,N_15715);
or U21847 (N_21847,N_19229,N_18697);
nand U21848 (N_21848,N_19566,N_19541);
xnor U21849 (N_21849,N_16501,N_16068);
nor U21850 (N_21850,N_17793,N_17005);
nor U21851 (N_21851,N_19001,N_19325);
nor U21852 (N_21852,N_19347,N_16726);
xor U21853 (N_21853,N_17050,N_15251);
or U21854 (N_21854,N_19322,N_18363);
or U21855 (N_21855,N_19385,N_17281);
and U21856 (N_21856,N_15123,N_15816);
and U21857 (N_21857,N_19443,N_18641);
nor U21858 (N_21858,N_16537,N_18159);
and U21859 (N_21859,N_18093,N_15116);
nor U21860 (N_21860,N_18173,N_17917);
nand U21861 (N_21861,N_15908,N_16526);
nor U21862 (N_21862,N_16469,N_18398);
and U21863 (N_21863,N_15593,N_16186);
nor U21864 (N_21864,N_19502,N_16121);
nand U21865 (N_21865,N_15210,N_17322);
or U21866 (N_21866,N_19343,N_16249);
and U21867 (N_21867,N_19056,N_18637);
and U21868 (N_21868,N_15596,N_16801);
or U21869 (N_21869,N_19633,N_18068);
nor U21870 (N_21870,N_19263,N_17518);
and U21871 (N_21871,N_18217,N_15018);
nand U21872 (N_21872,N_19960,N_15376);
xnor U21873 (N_21873,N_19961,N_16753);
nand U21874 (N_21874,N_18197,N_16542);
xnor U21875 (N_21875,N_19631,N_15827);
xnor U21876 (N_21876,N_17668,N_19430);
or U21877 (N_21877,N_17082,N_15731);
and U21878 (N_21878,N_18500,N_16240);
or U21879 (N_21879,N_15050,N_17387);
and U21880 (N_21880,N_17030,N_19545);
or U21881 (N_21881,N_15075,N_16908);
and U21882 (N_21882,N_19244,N_18225);
nor U21883 (N_21883,N_16493,N_19991);
nand U21884 (N_21884,N_17230,N_19175);
or U21885 (N_21885,N_18427,N_19312);
or U21886 (N_21886,N_15058,N_16716);
nor U21887 (N_21887,N_16403,N_18688);
and U21888 (N_21888,N_18666,N_17164);
nand U21889 (N_21889,N_18203,N_17543);
nor U21890 (N_21890,N_18042,N_17530);
nand U21891 (N_21891,N_16564,N_19464);
or U21892 (N_21892,N_18918,N_15851);
and U21893 (N_21893,N_16524,N_17754);
nor U21894 (N_21894,N_17104,N_19648);
nand U21895 (N_21895,N_17981,N_18584);
nand U21896 (N_21896,N_19483,N_19402);
nand U21897 (N_21897,N_17231,N_19421);
xnor U21898 (N_21898,N_18430,N_17948);
nand U21899 (N_21899,N_16895,N_19110);
xor U21900 (N_21900,N_19409,N_17739);
xnor U21901 (N_21901,N_16608,N_17588);
or U21902 (N_21902,N_17508,N_19870);
nor U21903 (N_21903,N_16611,N_15682);
nor U21904 (N_21904,N_15291,N_15526);
nor U21905 (N_21905,N_15256,N_16694);
nor U21906 (N_21906,N_18260,N_17654);
or U21907 (N_21907,N_18257,N_19711);
or U21908 (N_21908,N_19659,N_15187);
nand U21909 (N_21909,N_17497,N_19084);
and U21910 (N_21910,N_16636,N_19173);
and U21911 (N_21911,N_18915,N_15183);
or U21912 (N_21912,N_16109,N_19534);
nor U21913 (N_21913,N_16323,N_17698);
nor U21914 (N_21914,N_19824,N_17988);
nor U21915 (N_21915,N_18013,N_19054);
nand U21916 (N_21916,N_15807,N_19427);
and U21917 (N_21917,N_16538,N_15648);
nor U21918 (N_21918,N_15464,N_17812);
and U21919 (N_21919,N_15965,N_18582);
and U21920 (N_21920,N_15403,N_19798);
nand U21921 (N_21921,N_15446,N_19068);
and U21922 (N_21922,N_16851,N_19765);
nand U21923 (N_21923,N_18310,N_19610);
or U21924 (N_21924,N_19231,N_17923);
nor U21925 (N_21925,N_19771,N_17018);
and U21926 (N_21926,N_19445,N_18448);
xor U21927 (N_21927,N_19833,N_19469);
nor U21928 (N_21928,N_17080,N_15841);
and U21929 (N_21929,N_17515,N_15474);
and U21930 (N_21930,N_17352,N_16351);
nand U21931 (N_21931,N_17538,N_15920);
nor U21932 (N_21932,N_19367,N_17136);
nor U21933 (N_21933,N_19081,N_15333);
and U21934 (N_21934,N_16734,N_15489);
and U21935 (N_21935,N_16481,N_18835);
and U21936 (N_21936,N_17997,N_17345);
nand U21937 (N_21937,N_16238,N_17046);
nor U21938 (N_21938,N_16907,N_17116);
nand U21939 (N_21939,N_16778,N_16269);
nor U21940 (N_21940,N_15937,N_16361);
xnor U21941 (N_21941,N_18124,N_15840);
nor U21942 (N_21942,N_17237,N_17321);
xnor U21943 (N_21943,N_16041,N_19901);
and U21944 (N_21944,N_15522,N_18142);
nor U21945 (N_21945,N_17190,N_16096);
and U21946 (N_21946,N_18814,N_18887);
nor U21947 (N_21947,N_16519,N_19540);
or U21948 (N_21948,N_16110,N_17832);
and U21949 (N_21949,N_16782,N_15314);
nor U21950 (N_21950,N_16520,N_17333);
nor U21951 (N_21951,N_19342,N_18963);
xnor U21952 (N_21952,N_15477,N_18675);
nor U21953 (N_21953,N_15082,N_17863);
xor U21954 (N_21954,N_19005,N_19737);
and U21955 (N_21955,N_15460,N_16235);
or U21956 (N_21956,N_19749,N_18472);
nor U21957 (N_21957,N_16431,N_16000);
nor U21958 (N_21958,N_18246,N_18792);
or U21959 (N_21959,N_17330,N_19236);
or U21960 (N_21960,N_18758,N_18228);
nand U21961 (N_21961,N_15883,N_16738);
nand U21962 (N_21962,N_19245,N_19584);
and U21963 (N_21963,N_18889,N_18063);
nand U21964 (N_21964,N_17127,N_19942);
or U21965 (N_21965,N_19511,N_19587);
and U21966 (N_21966,N_17287,N_19133);
nand U21967 (N_21967,N_16330,N_18125);
nand U21968 (N_21968,N_18045,N_16600);
xnor U21969 (N_21969,N_19344,N_19239);
and U21970 (N_21970,N_16920,N_18186);
and U21971 (N_21971,N_19666,N_15534);
and U21972 (N_21972,N_15898,N_17911);
xor U21973 (N_21973,N_16258,N_17876);
xor U21974 (N_21974,N_16558,N_16140);
nand U21975 (N_21975,N_15983,N_18910);
nand U21976 (N_21976,N_18202,N_17811);
xor U21977 (N_21977,N_19981,N_19078);
nand U21978 (N_21978,N_16013,N_17978);
and U21979 (N_21979,N_19902,N_17925);
and U21980 (N_21980,N_15653,N_19569);
xnor U21981 (N_21981,N_16810,N_16575);
xor U21982 (N_21982,N_15539,N_18070);
nand U21983 (N_21983,N_16755,N_18622);
nor U21984 (N_21984,N_16261,N_16210);
or U21985 (N_21985,N_17872,N_16148);
nor U21986 (N_21986,N_18406,N_18626);
and U21987 (N_21987,N_19247,N_18452);
nor U21988 (N_21988,N_15484,N_16798);
nor U21989 (N_21989,N_19851,N_16135);
and U21990 (N_21990,N_17151,N_19401);
nor U21991 (N_21991,N_17085,N_16614);
xnor U21992 (N_21992,N_15119,N_19268);
nor U21993 (N_21993,N_18308,N_17114);
or U21994 (N_21994,N_18026,N_19544);
xnor U21995 (N_21995,N_17609,N_18779);
nand U21996 (N_21996,N_18209,N_19062);
or U21997 (N_21997,N_17430,N_19822);
and U21998 (N_21998,N_16933,N_15870);
nand U21999 (N_21999,N_17009,N_17172);
xnor U22000 (N_22000,N_15644,N_16188);
xnor U22001 (N_22001,N_16029,N_19775);
and U22002 (N_22002,N_15249,N_17627);
xor U22003 (N_22003,N_18264,N_15229);
nand U22004 (N_22004,N_16470,N_18413);
nand U22005 (N_22005,N_15613,N_16835);
xor U22006 (N_22006,N_15536,N_18253);
or U22007 (N_22007,N_19126,N_17555);
or U22008 (N_22008,N_15274,N_19655);
or U22009 (N_22009,N_19494,N_16521);
and U22010 (N_22010,N_16411,N_19492);
xnor U22011 (N_22011,N_17229,N_16974);
and U22012 (N_22012,N_17703,N_17646);
xor U22013 (N_22013,N_17949,N_15493);
and U22014 (N_22014,N_15558,N_17858);
or U22015 (N_22015,N_17657,N_18213);
xnor U22016 (N_22016,N_18986,N_19392);
nor U22017 (N_22017,N_17125,N_19341);
xnor U22018 (N_22018,N_16813,N_17743);
or U22019 (N_22019,N_18009,N_17353);
xor U22020 (N_22020,N_18276,N_16255);
and U22021 (N_22021,N_15790,N_19335);
or U22022 (N_22022,N_17720,N_18794);
nand U22023 (N_22023,N_19562,N_16365);
and U22024 (N_22024,N_17468,N_19286);
nor U22025 (N_22025,N_17038,N_15287);
or U22026 (N_22026,N_15276,N_18852);
or U22027 (N_22027,N_15329,N_19884);
xnor U22028 (N_22028,N_15338,N_19070);
xnor U22029 (N_22029,N_15921,N_16763);
or U22030 (N_22030,N_18199,N_19993);
xor U22031 (N_22031,N_17592,N_17075);
and U22032 (N_22032,N_15843,N_15806);
and U22033 (N_22033,N_15325,N_17222);
xor U22034 (N_22034,N_18530,N_15330);
or U22035 (N_22035,N_16947,N_16272);
nor U22036 (N_22036,N_15510,N_16606);
nand U22037 (N_22037,N_16417,N_15281);
and U22038 (N_22038,N_19938,N_17094);
xnor U22039 (N_22039,N_18423,N_17025);
nor U22040 (N_22040,N_17021,N_15138);
nand U22041 (N_22041,N_15725,N_19996);
xor U22042 (N_22042,N_19828,N_18314);
nor U22043 (N_22043,N_15714,N_16091);
nor U22044 (N_22044,N_16596,N_18205);
nor U22045 (N_22045,N_19008,N_15038);
xor U22046 (N_22046,N_19501,N_16171);
xnor U22047 (N_22047,N_17446,N_16623);
xnor U22048 (N_22048,N_16344,N_18378);
and U22049 (N_22049,N_16339,N_19634);
xnor U22050 (N_22050,N_16987,N_18175);
or U22051 (N_22051,N_16536,N_18342);
xnor U22052 (N_22052,N_17259,N_15967);
and U22053 (N_22053,N_19252,N_19573);
or U22054 (N_22054,N_18360,N_19972);
nand U22055 (N_22055,N_19637,N_15061);
xnor U22056 (N_22056,N_17306,N_17504);
or U22057 (N_22057,N_16200,N_17421);
and U22058 (N_22058,N_16730,N_16285);
nand U22059 (N_22059,N_19027,N_16422);
nand U22060 (N_22060,N_18941,N_19933);
or U22061 (N_22061,N_17566,N_17537);
and U22062 (N_22062,N_18931,N_16111);
nand U22063 (N_22063,N_18479,N_19739);
nor U22064 (N_22064,N_18644,N_18410);
nor U22065 (N_22065,N_17088,N_15379);
xnor U22066 (N_22066,N_15638,N_15608);
and U22067 (N_22067,N_16290,N_18659);
or U22068 (N_22068,N_17011,N_15583);
and U22069 (N_22069,N_18444,N_18973);
nor U22070 (N_22070,N_18636,N_19705);
xnor U22071 (N_22071,N_18570,N_18943);
or U22072 (N_22072,N_17550,N_15947);
or U22073 (N_22073,N_15952,N_19679);
nor U22074 (N_22074,N_19080,N_16356);
and U22075 (N_22075,N_15421,N_17800);
nor U22076 (N_22076,N_19620,N_17756);
nand U22077 (N_22077,N_17844,N_15110);
or U22078 (N_22078,N_16928,N_16888);
nor U22079 (N_22079,N_16505,N_16463);
xor U22080 (N_22080,N_18753,N_15925);
or U22081 (N_22081,N_17070,N_19375);
xor U22082 (N_22082,N_15478,N_17578);
and U22083 (N_22083,N_19970,N_15662);
or U22084 (N_22084,N_15923,N_15730);
or U22085 (N_22085,N_19918,N_16322);
nor U22086 (N_22086,N_15011,N_17304);
nor U22087 (N_22087,N_15916,N_17826);
and U22088 (N_22088,N_16229,N_15973);
nor U22089 (N_22089,N_15508,N_15544);
xnor U22090 (N_22090,N_19669,N_15782);
nand U22091 (N_22091,N_15313,N_19297);
nand U22092 (N_22092,N_16667,N_15875);
nand U22093 (N_22093,N_18998,N_19675);
or U22094 (N_22094,N_17820,N_16283);
or U22095 (N_22095,N_15700,N_16841);
xor U22096 (N_22096,N_19723,N_15881);
and U22097 (N_22097,N_15869,N_16605);
xor U22098 (N_22098,N_16634,N_15365);
or U22099 (N_22099,N_18893,N_15311);
nand U22100 (N_22100,N_17585,N_18409);
nor U22101 (N_22101,N_19522,N_17414);
xor U22102 (N_22102,N_17143,N_19831);
and U22103 (N_22103,N_16508,N_15357);
nand U22104 (N_22104,N_15636,N_18603);
nor U22105 (N_22105,N_19418,N_19969);
nor U22106 (N_22106,N_19616,N_17111);
or U22107 (N_22107,N_16004,N_17402);
nand U22108 (N_22108,N_18916,N_15245);
or U22109 (N_22109,N_16372,N_16151);
xor U22110 (N_22110,N_16846,N_15506);
and U22111 (N_22111,N_19298,N_18775);
nor U22112 (N_22112,N_19908,N_18119);
or U22113 (N_22113,N_15594,N_19321);
nand U22114 (N_22114,N_17877,N_19746);
xor U22115 (N_22115,N_15024,N_19504);
nand U22116 (N_22116,N_16458,N_17261);
nand U22117 (N_22117,N_19740,N_16155);
nor U22118 (N_22118,N_19694,N_16253);
and U22119 (N_22119,N_16163,N_17129);
or U22120 (N_22120,N_17150,N_16207);
and U22121 (N_22121,N_15546,N_19556);
and U22122 (N_22122,N_18362,N_17235);
xor U22123 (N_22123,N_17594,N_17946);
or U22124 (N_22124,N_17278,N_15340);
and U22125 (N_22125,N_16629,N_15674);
nor U22126 (N_22126,N_17510,N_15609);
and U22127 (N_22127,N_19678,N_15709);
nor U22128 (N_22128,N_18496,N_19887);
xnor U22129 (N_22129,N_19191,N_16291);
nand U22130 (N_22130,N_16698,N_16302);
nor U22131 (N_22131,N_19488,N_16588);
or U22132 (N_22132,N_19058,N_17897);
nor U22133 (N_22133,N_19708,N_18692);
or U22134 (N_22134,N_15660,N_17630);
or U22135 (N_22135,N_18822,N_19043);
xor U22136 (N_22136,N_15978,N_15579);
or U22137 (N_22137,N_15671,N_15086);
nor U22138 (N_22138,N_18304,N_17985);
xor U22139 (N_22139,N_19796,N_18720);
xor U22140 (N_22140,N_15918,N_17829);
nand U22141 (N_22141,N_19129,N_18825);
xnor U22142 (N_22142,N_19381,N_17623);
xnor U22143 (N_22143,N_16535,N_16273);
xor U22144 (N_22144,N_17823,N_16094);
xnor U22145 (N_22145,N_17963,N_15485);
and U22146 (N_22146,N_18722,N_16673);
xor U22147 (N_22147,N_18776,N_15079);
xnor U22148 (N_22148,N_17801,N_15563);
and U22149 (N_22149,N_15518,N_17189);
nand U22150 (N_22150,N_16312,N_19113);
xor U22151 (N_22151,N_17941,N_15560);
nand U22152 (N_22152,N_17631,N_16914);
nor U22153 (N_22153,N_17416,N_19662);
nor U22154 (N_22154,N_18358,N_17455);
or U22155 (N_22155,N_17705,N_16776);
nand U22156 (N_22156,N_17370,N_15029);
or U22157 (N_22157,N_17805,N_15864);
or U22158 (N_22158,N_17874,N_17717);
or U22159 (N_22159,N_16569,N_15289);
and U22160 (N_22160,N_18815,N_17040);
nor U22161 (N_22161,N_18858,N_17973);
and U22162 (N_22162,N_19853,N_18975);
xnor U22163 (N_22163,N_18588,N_17193);
or U22164 (N_22164,N_16014,N_15729);
nand U22165 (N_22165,N_17924,N_19709);
nand U22166 (N_22166,N_16496,N_15530);
nor U22167 (N_22167,N_18204,N_16511);
xor U22168 (N_22168,N_19480,N_17659);
xor U22169 (N_22169,N_17135,N_18924);
or U22170 (N_22170,N_18995,N_17410);
nor U22171 (N_22171,N_16769,N_19621);
nand U22172 (N_22172,N_17649,N_15819);
or U22173 (N_22173,N_18935,N_19706);
or U22174 (N_22174,N_19077,N_15156);
and U22175 (N_22175,N_16647,N_15996);
and U22176 (N_22176,N_15582,N_18959);
and U22177 (N_22177,N_19813,N_19450);
and U22178 (N_22178,N_16471,N_18370);
xnor U22179 (N_22179,N_17514,N_15400);
nor U22180 (N_22180,N_17042,N_19455);
nand U22181 (N_22181,N_16456,N_15541);
and U22182 (N_22182,N_19529,N_15004);
or U22183 (N_22183,N_16723,N_17240);
nand U22184 (N_22184,N_16701,N_18501);
nor U22185 (N_22185,N_16811,N_17496);
nand U22186 (N_22186,N_18016,N_18769);
nor U22187 (N_22187,N_19978,N_17234);
xnor U22188 (N_22188,N_15306,N_17968);
xor U22189 (N_22189,N_17102,N_18083);
xor U22190 (N_22190,N_15770,N_19311);
and U22191 (N_22191,N_16001,N_19809);
and U22192 (N_22192,N_16400,N_16873);
nor U22193 (N_22193,N_18640,N_16952);
xor U22194 (N_22194,N_18817,N_19376);
nand U22195 (N_22195,N_15748,N_19726);
and U22196 (N_22196,N_19404,N_18502);
nand U22197 (N_22197,N_18469,N_16286);
nand U22198 (N_22198,N_18568,N_15343);
or U22199 (N_22199,N_19856,N_18714);
xnor U22200 (N_22200,N_18351,N_15756);
xor U22201 (N_22201,N_15171,N_16172);
nor U22202 (N_22202,N_15160,N_19758);
xor U22203 (N_22203,N_18725,N_18625);
nand U22204 (N_22204,N_15347,N_19423);
or U22205 (N_22205,N_16149,N_18137);
or U22206 (N_22206,N_16909,N_16584);
and U22207 (N_22207,N_16658,N_17265);
or U22208 (N_22208,N_18044,N_17010);
nand U22209 (N_22209,N_17704,N_16097);
or U22210 (N_22210,N_18099,N_18371);
xnor U22211 (N_22211,N_18107,N_18522);
nor U22212 (N_22212,N_19493,N_17542);
and U22213 (N_22213,N_17073,N_15538);
or U22214 (N_22214,N_17280,N_19911);
and U22215 (N_22215,N_17369,N_19000);
xor U22216 (N_22216,N_15884,N_15677);
xnor U22217 (N_22217,N_19462,N_15945);
nand U22218 (N_22218,N_16975,N_16808);
and U22219 (N_22219,N_17086,N_15914);
and U22220 (N_22220,N_17513,N_15490);
xor U22221 (N_22221,N_17263,N_17565);
nand U22222 (N_22222,N_16117,N_19250);
or U22223 (N_22223,N_19122,N_17851);
xor U22224 (N_22224,N_19233,N_17233);
nor U22225 (N_22225,N_17368,N_18619);
nand U22226 (N_22226,N_16346,N_17341);
xor U22227 (N_22227,N_19919,N_18900);
or U22228 (N_22228,N_15726,N_18932);
or U22229 (N_22229,N_15469,N_16120);
and U22230 (N_22230,N_16324,N_18922);
nand U22231 (N_22231,N_15618,N_19320);
nand U22232 (N_22232,N_17084,N_15789);
or U22233 (N_22233,N_18604,N_18971);
or U22234 (N_22234,N_18392,N_19946);
or U22235 (N_22235,N_18803,N_15142);
or U22236 (N_22236,N_16116,N_17323);
nand U22237 (N_22237,N_18335,N_17824);
nor U22238 (N_22238,N_18694,N_19889);
nor U22239 (N_22239,N_15941,N_15580);
or U22240 (N_22240,N_18485,N_17471);
xnor U22241 (N_22241,N_15569,N_17134);
and U22242 (N_22242,N_15844,N_15420);
xor U22243 (N_22243,N_15523,N_18297);
nand U22244 (N_22244,N_18509,N_15438);
nand U22245 (N_22245,N_18930,N_16401);
and U22246 (N_22246,N_18098,N_17122);
nand U22247 (N_22247,N_17313,N_16017);
and U22248 (N_22248,N_17600,N_18649);
or U22249 (N_22249,N_17092,N_16357);
and U22250 (N_22250,N_18133,N_19481);
nor U22251 (N_22251,N_16516,N_19150);
and U22252 (N_22252,N_19639,N_16316);
and U22253 (N_22253,N_19721,N_15944);
and U22254 (N_22254,N_18049,N_15292);
or U22255 (N_22255,N_15043,N_15363);
nand U22256 (N_22256,N_18128,N_18003);
xnor U22257 (N_22257,N_17881,N_15049);
or U22258 (N_22258,N_16918,N_19838);
or U22259 (N_22259,N_17904,N_16306);
nand U22260 (N_22260,N_19795,N_17797);
nand U22261 (N_22261,N_17344,N_15162);
or U22262 (N_22262,N_15328,N_19551);
nor U22263 (N_22263,N_15437,N_17880);
nor U22264 (N_22264,N_15166,N_17045);
or U22265 (N_22265,N_19898,N_19115);
nor U22266 (N_22266,N_16232,N_18632);
or U22267 (N_22267,N_16953,N_19903);
or U22268 (N_22268,N_17991,N_17706);
or U22269 (N_22269,N_18443,N_15399);
xor U22270 (N_22270,N_19953,N_15825);
nand U22271 (N_22271,N_15664,N_18306);
xor U22272 (N_22272,N_18895,N_18901);
and U22273 (N_22273,N_15299,N_16855);
or U22274 (N_22274,N_15760,N_19915);
nor U22275 (N_22275,N_19673,N_17962);
nor U22276 (N_22276,N_18891,N_16729);
nand U22277 (N_22277,N_19849,N_19289);
xnor U22278 (N_22278,N_17374,N_16432);
or U22279 (N_22279,N_19349,N_18486);
and U22280 (N_22280,N_18629,N_17173);
or U22281 (N_22281,N_16176,N_18780);
or U22282 (N_22282,N_18106,N_18275);
nand U22283 (N_22283,N_17214,N_17546);
nor U22284 (N_22284,N_15867,N_18361);
or U22285 (N_22285,N_18607,N_19959);
xor U22286 (N_22286,N_19441,N_15625);
and U22287 (N_22287,N_19380,N_15866);
nand U22288 (N_22288,N_17218,N_17298);
nand U22289 (N_22289,N_19163,N_19026);
nor U22290 (N_22290,N_17096,N_15395);
or U22291 (N_22291,N_15233,N_18526);
xnor U22292 (N_22292,N_15657,N_19827);
or U22293 (N_22293,N_17702,N_17413);
or U22294 (N_22294,N_15525,N_15307);
nor U22295 (N_22295,N_15220,N_15423);
or U22296 (N_22296,N_18529,N_17584);
xor U22297 (N_22297,N_15089,N_18988);
nor U22298 (N_22298,N_15482,N_16160);
xnor U22299 (N_22299,N_17168,N_19411);
nor U22300 (N_22300,N_16997,N_16426);
and U22301 (N_22301,N_18880,N_19667);
or U22302 (N_22302,N_19045,N_16042);
nand U22303 (N_22303,N_16977,N_15741);
nand U22304 (N_22304,N_19123,N_17547);
and U22305 (N_22305,N_19378,N_17153);
nor U22306 (N_22306,N_18066,N_15396);
and U22307 (N_22307,N_16860,N_16190);
and U22308 (N_22308,N_17347,N_17759);
xnor U22309 (N_22309,N_15294,N_17058);
or U22310 (N_22310,N_17738,N_17385);
xor U22311 (N_22311,N_16408,N_15457);
xor U22312 (N_22312,N_19142,N_19301);
and U22313 (N_22313,N_19750,N_18606);
nand U22314 (N_22314,N_17838,N_16319);
nor U22315 (N_22315,N_16126,N_15129);
xor U22316 (N_22316,N_17060,N_18740);
and U22317 (N_22317,N_15673,N_15214);
or U22318 (N_22318,N_18379,N_16224);
nor U22319 (N_22319,N_18781,N_19785);
and U22320 (N_22320,N_17862,N_16265);
nand U22321 (N_22321,N_17486,N_19002);
or U22322 (N_22322,N_18695,N_16304);
nor U22323 (N_22323,N_15758,N_16139);
and U22324 (N_22324,N_16779,N_18949);
and U22325 (N_22325,N_19314,N_19053);
or U22326 (N_22326,N_16381,N_18533);
nand U22327 (N_22327,N_16865,N_19604);
and U22328 (N_22328,N_16590,N_15661);
or U22329 (N_22329,N_19033,N_19873);
xnor U22330 (N_22330,N_16075,N_19528);
nor U22331 (N_22331,N_15013,N_19472);
nor U22332 (N_22332,N_16585,N_15118);
nor U22333 (N_22333,N_19299,N_17068);
or U22334 (N_22334,N_15876,N_19121);
and U22335 (N_22335,N_19063,N_18552);
and U22336 (N_22336,N_18224,N_16448);
xnor U22337 (N_22337,N_18162,N_15431);
and U22338 (N_22338,N_17098,N_18153);
and U22339 (N_22339,N_16805,N_18145);
or U22340 (N_22340,N_19617,N_18231);
nor U22341 (N_22341,N_19422,N_15030);
nor U22342 (N_22342,N_19171,N_16331);
and U22343 (N_22343,N_17679,N_18599);
xor U22344 (N_22344,N_18521,N_19552);
or U22345 (N_22345,N_19112,N_16744);
nand U22346 (N_22346,N_17213,N_17637);
and U22347 (N_22347,N_19300,N_17470);
xnor U22348 (N_22348,N_17670,N_15772);
nor U22349 (N_22349,N_15155,N_15763);
nor U22350 (N_22350,N_15587,N_16242);
and U22351 (N_22351,N_18961,N_15121);
nor U22352 (N_22352,N_18340,N_17415);
nor U22353 (N_22353,N_15394,N_18843);
xnor U22354 (N_22354,N_19790,N_17396);
nand U22355 (N_22355,N_18271,N_16076);
or U22356 (N_22356,N_18718,N_17247);
or U22357 (N_22357,N_18471,N_17750);
xor U22358 (N_22358,N_18143,N_15386);
xnor U22359 (N_22359,N_18181,N_19595);
and U22360 (N_22360,N_19193,N_18376);
xor U22361 (N_22361,N_16196,N_17977);
and U22362 (N_22362,N_16018,N_15676);
nand U22363 (N_22363,N_16161,N_15443);
or U22364 (N_22364,N_15105,N_16874);
xnor U22365 (N_22365,N_16220,N_15732);
and U22366 (N_22366,N_19656,N_18527);
and U22367 (N_22367,N_15956,N_18163);
nand U22368 (N_22368,N_16370,N_15639);
or U22369 (N_22369,N_15611,N_16714);
xnor U22370 (N_22370,N_18060,N_19733);
and U22371 (N_22371,N_17123,N_16702);
or U22372 (N_22372,N_19814,N_18754);
and U22373 (N_22373,N_18100,N_18828);
xor U22374 (N_22374,N_17290,N_18300);
nand U22375 (N_22375,N_17878,N_16327);
or U22376 (N_22376,N_17996,N_15001);
xnor U22377 (N_22377,N_17901,N_15381);
nand U22378 (N_22378,N_15248,N_15781);
or U22379 (N_22379,N_17850,N_18090);
nor U22380 (N_22380,N_19927,N_16619);
and U22381 (N_22381,N_17023,N_19177);
and U22382 (N_22382,N_18105,N_15545);
and U22383 (N_22383,N_19285,N_18147);
nand U22384 (N_22384,N_17960,N_15351);
nand U22385 (N_22385,N_19826,N_19594);
and U22386 (N_22386,N_17103,N_15799);
xor U22387 (N_22387,N_17519,N_18295);
xnor U22388 (N_22388,N_17157,N_18249);
nand U22389 (N_22389,N_18914,N_17713);
nand U22390 (N_22390,N_15879,N_16642);
and U22391 (N_22391,N_18968,N_18470);
or U22392 (N_22392,N_18672,N_15025);
nor U22393 (N_22393,N_18830,N_15859);
or U22394 (N_22394,N_19623,N_19351);
and U22395 (N_22395,N_18634,N_15471);
or U22396 (N_22396,N_15577,N_19578);
nor U22397 (N_22397,N_18494,N_17483);
xnor U22398 (N_22398,N_16943,N_16884);
and U22399 (N_22399,N_17146,N_15987);
nor U22400 (N_22400,N_18120,N_19731);
nand U22401 (N_22401,N_15964,N_17711);
xnor U22402 (N_22402,N_16646,N_18233);
xor U22403 (N_22403,N_17003,N_19921);
nor U22404 (N_22404,N_17619,N_15794);
nand U22405 (N_22405,N_15355,N_16886);
and U22406 (N_22406,N_18072,N_18450);
or U22407 (N_22407,N_15189,N_17648);
and U22408 (N_22408,N_16334,N_17270);
nand U22409 (N_22409,N_15955,N_15410);
or U22410 (N_22410,N_18352,N_19560);
nand U22411 (N_22411,N_16842,N_16545);
or U22412 (N_22412,N_15369,N_18460);
or U22413 (N_22413,N_18813,N_16277);
xor U22414 (N_22414,N_19531,N_15418);
and U22415 (N_22415,N_17582,N_18270);
or U22416 (N_22416,N_17006,N_19660);
nor U22417 (N_22417,N_15809,N_16910);
xor U22418 (N_22418,N_17984,N_16807);
nand U22419 (N_22419,N_16547,N_15710);
and U22420 (N_22420,N_16650,N_17898);
and U22421 (N_22421,N_16504,N_19372);
nand U22422 (N_22422,N_17147,N_16278);
or U22423 (N_22423,N_15979,N_15419);
nor U22424 (N_22424,N_15481,N_18913);
nor U22425 (N_22425,N_17177,N_18872);
xnor U22426 (N_22426,N_17502,N_16919);
nor U22427 (N_22427,N_19489,N_17549);
nor U22428 (N_22428,N_19698,N_15107);
and U22429 (N_22429,N_15771,N_15006);
xnor U22430 (N_22430,N_16233,N_19936);
nand U22431 (N_22431,N_18254,N_18078);
nand U22432 (N_22432,N_19313,N_18600);
and U22433 (N_22433,N_16468,N_18250);
nand U22434 (N_22434,N_17914,N_19003);
or U22435 (N_22435,N_18041,N_16659);
xor U22436 (N_22436,N_17083,N_17158);
and U22437 (N_22437,N_17062,N_17493);
and U22438 (N_22438,N_19895,N_15542);
nor U22439 (N_22439,N_17181,N_19850);
nand U22440 (N_22440,N_17469,N_19011);
and U22441 (N_22441,N_19465,N_18651);
and U22442 (N_22442,N_16936,N_19117);
and U22443 (N_22443,N_17950,N_15751);
nand U22444 (N_22444,N_15218,N_16819);
or U22445 (N_22445,N_17339,N_18912);
xor U22446 (N_22446,N_15216,N_18323);
nor U22447 (N_22447,N_16115,N_17427);
or U22448 (N_22448,N_17689,N_16700);
nand U22449 (N_22449,N_16009,N_15444);
or U22450 (N_22450,N_17420,N_19203);
or U22451 (N_22451,N_18418,N_15470);
nor U22452 (N_22452,N_17907,N_16299);
nor U22453 (N_22453,N_19589,N_19238);
and U22454 (N_22454,N_15498,N_15285);
nor U22455 (N_22455,N_19636,N_15346);
or U22456 (N_22456,N_16688,N_17506);
xnor U22457 (N_22457,N_16054,N_15999);
xor U22458 (N_22458,N_17790,N_18768);
or U22459 (N_22459,N_17775,N_15017);
xor U22460 (N_22460,N_16930,N_16069);
nor U22461 (N_22461,N_17022,N_17393);
nor U22462 (N_22462,N_17777,N_17836);
nand U22463 (N_22463,N_19592,N_15111);
nor U22464 (N_22464,N_15894,N_16497);
and U22465 (N_22465,N_16244,N_19672);
or U22466 (N_22466,N_17202,N_15392);
or U22467 (N_22467,N_19348,N_17433);
or U22468 (N_22468,N_16577,N_19420);
and U22469 (N_22469,N_16633,N_17745);
nand U22470 (N_22470,N_17479,N_17875);
nand U22471 (N_22471,N_18428,N_16893);
or U22472 (N_22472,N_15375,N_19222);
and U22473 (N_22473,N_16487,N_15349);
and U22474 (N_22474,N_18763,N_17601);
xnor U22475 (N_22475,N_19046,N_18492);
nand U22476 (N_22476,N_16396,N_17494);
nand U22477 (N_22477,N_17692,N_19438);
and U22478 (N_22478,N_16103,N_19762);
xor U22479 (N_22479,N_17653,N_18761);
and U22480 (N_22480,N_17194,N_15301);
nor U22481 (N_22481,N_19949,N_15646);
and U22482 (N_22482,N_16950,N_16630);
or U22483 (N_22483,N_17644,N_15701);
nand U22484 (N_22484,N_15272,N_15699);
or U22485 (N_22485,N_15087,N_18819);
nand U22486 (N_22486,N_18008,N_16335);
or U22487 (N_22487,N_19954,N_17291);
or U22488 (N_22488,N_16586,N_18266);
nand U22489 (N_22489,N_19618,N_18793);
nand U22490 (N_22490,N_17412,N_18539);
nand U22491 (N_22491,N_16553,N_17994);
or U22492 (N_22492,N_17620,N_17699);
nand U22493 (N_22493,N_16022,N_16668);
xnor U22494 (N_22494,N_19929,N_17426);
and U22495 (N_22495,N_15264,N_19934);
xor U22496 (N_22496,N_17362,N_17524);
or U22497 (N_22497,N_16829,N_17372);
and U22498 (N_22498,N_18116,N_16576);
xor U22499 (N_22499,N_16637,N_17320);
xor U22500 (N_22500,N_16801,N_19535);
nand U22501 (N_22501,N_19471,N_15145);
or U22502 (N_22502,N_15941,N_16275);
nor U22503 (N_22503,N_17469,N_16426);
and U22504 (N_22504,N_15182,N_18167);
nand U22505 (N_22505,N_16894,N_19371);
nor U22506 (N_22506,N_15193,N_16171);
xnor U22507 (N_22507,N_19703,N_19629);
nand U22508 (N_22508,N_17073,N_15822);
or U22509 (N_22509,N_15358,N_18308);
nor U22510 (N_22510,N_17772,N_18756);
nor U22511 (N_22511,N_17982,N_18306);
and U22512 (N_22512,N_15557,N_18761);
xnor U22513 (N_22513,N_19662,N_19863);
nand U22514 (N_22514,N_15091,N_17745);
xnor U22515 (N_22515,N_17246,N_18991);
nand U22516 (N_22516,N_18789,N_16894);
and U22517 (N_22517,N_18581,N_15524);
nor U22518 (N_22518,N_16930,N_17974);
nand U22519 (N_22519,N_15431,N_15944);
or U22520 (N_22520,N_17293,N_15324);
xor U22521 (N_22521,N_17121,N_19736);
xor U22522 (N_22522,N_19706,N_19484);
or U22523 (N_22523,N_15495,N_15282);
or U22524 (N_22524,N_16554,N_15146);
nor U22525 (N_22525,N_15417,N_15100);
nor U22526 (N_22526,N_16982,N_17702);
nand U22527 (N_22527,N_17846,N_18475);
nor U22528 (N_22528,N_15237,N_16368);
or U22529 (N_22529,N_19311,N_18835);
xnor U22530 (N_22530,N_15160,N_15736);
and U22531 (N_22531,N_15270,N_16466);
nand U22532 (N_22532,N_18159,N_15670);
nand U22533 (N_22533,N_15734,N_18434);
nor U22534 (N_22534,N_19181,N_16465);
nand U22535 (N_22535,N_18637,N_15366);
and U22536 (N_22536,N_15897,N_17804);
and U22537 (N_22537,N_15534,N_18883);
and U22538 (N_22538,N_17773,N_17613);
or U22539 (N_22539,N_15253,N_17825);
nor U22540 (N_22540,N_15441,N_19289);
xnor U22541 (N_22541,N_18966,N_18845);
xnor U22542 (N_22542,N_17519,N_19137);
nor U22543 (N_22543,N_18196,N_17244);
or U22544 (N_22544,N_17717,N_17365);
nand U22545 (N_22545,N_18711,N_19901);
and U22546 (N_22546,N_17897,N_17289);
and U22547 (N_22547,N_18874,N_17620);
or U22548 (N_22548,N_17612,N_19581);
xor U22549 (N_22549,N_15570,N_17752);
nand U22550 (N_22550,N_15877,N_16326);
nand U22551 (N_22551,N_17445,N_19766);
xnor U22552 (N_22552,N_18523,N_15466);
and U22553 (N_22553,N_19250,N_16667);
nor U22554 (N_22554,N_18329,N_19867);
nor U22555 (N_22555,N_19752,N_18478);
nor U22556 (N_22556,N_15938,N_15015);
nand U22557 (N_22557,N_17087,N_19034);
and U22558 (N_22558,N_15482,N_17476);
xor U22559 (N_22559,N_17207,N_18301);
xnor U22560 (N_22560,N_18739,N_16208);
or U22561 (N_22561,N_15355,N_16917);
or U22562 (N_22562,N_16254,N_15637);
nand U22563 (N_22563,N_15853,N_19211);
xnor U22564 (N_22564,N_15236,N_17185);
or U22565 (N_22565,N_18758,N_19636);
and U22566 (N_22566,N_16881,N_19270);
nand U22567 (N_22567,N_18198,N_16954);
nand U22568 (N_22568,N_16467,N_18391);
and U22569 (N_22569,N_15148,N_17649);
nor U22570 (N_22570,N_18436,N_17645);
and U22571 (N_22571,N_18799,N_19360);
nand U22572 (N_22572,N_17341,N_16751);
or U22573 (N_22573,N_17752,N_19719);
xor U22574 (N_22574,N_15530,N_16138);
nor U22575 (N_22575,N_18148,N_15929);
nand U22576 (N_22576,N_18881,N_15852);
or U22577 (N_22577,N_18090,N_15429);
nor U22578 (N_22578,N_19616,N_15857);
or U22579 (N_22579,N_16269,N_17947);
and U22580 (N_22580,N_15325,N_18607);
and U22581 (N_22581,N_15924,N_18218);
nor U22582 (N_22582,N_15636,N_16018);
xnor U22583 (N_22583,N_17800,N_18112);
nand U22584 (N_22584,N_19547,N_17141);
or U22585 (N_22585,N_16813,N_18626);
or U22586 (N_22586,N_19963,N_15295);
xnor U22587 (N_22587,N_15123,N_18144);
xor U22588 (N_22588,N_19878,N_19096);
and U22589 (N_22589,N_16703,N_15230);
and U22590 (N_22590,N_17810,N_18424);
or U22591 (N_22591,N_18260,N_19194);
or U22592 (N_22592,N_16038,N_16854);
or U22593 (N_22593,N_18611,N_15885);
xnor U22594 (N_22594,N_18768,N_15749);
nor U22595 (N_22595,N_15287,N_15315);
nor U22596 (N_22596,N_15528,N_15982);
or U22597 (N_22597,N_16257,N_18312);
or U22598 (N_22598,N_16249,N_19080);
and U22599 (N_22599,N_15124,N_16374);
nor U22600 (N_22600,N_18232,N_17454);
and U22601 (N_22601,N_18073,N_19910);
or U22602 (N_22602,N_19218,N_17504);
nand U22603 (N_22603,N_18077,N_15803);
nand U22604 (N_22604,N_18701,N_18917);
or U22605 (N_22605,N_18927,N_18162);
nor U22606 (N_22606,N_17592,N_17299);
nor U22607 (N_22607,N_16012,N_18617);
nand U22608 (N_22608,N_17456,N_15177);
xor U22609 (N_22609,N_19078,N_19487);
xor U22610 (N_22610,N_17253,N_19475);
nor U22611 (N_22611,N_17789,N_17276);
xnor U22612 (N_22612,N_15647,N_15726);
nor U22613 (N_22613,N_19746,N_15653);
or U22614 (N_22614,N_15290,N_19991);
and U22615 (N_22615,N_19940,N_16573);
and U22616 (N_22616,N_15987,N_15383);
and U22617 (N_22617,N_18753,N_19556);
and U22618 (N_22618,N_16087,N_19379);
nor U22619 (N_22619,N_16793,N_15106);
or U22620 (N_22620,N_19019,N_17217);
xor U22621 (N_22621,N_18479,N_18250);
nor U22622 (N_22622,N_19113,N_16982);
xor U22623 (N_22623,N_17008,N_19344);
xnor U22624 (N_22624,N_16340,N_15989);
nand U22625 (N_22625,N_19526,N_16037);
nor U22626 (N_22626,N_15896,N_18606);
nor U22627 (N_22627,N_18542,N_16791);
nor U22628 (N_22628,N_15272,N_16794);
nand U22629 (N_22629,N_18812,N_16732);
xor U22630 (N_22630,N_15231,N_16521);
nand U22631 (N_22631,N_18451,N_15574);
nor U22632 (N_22632,N_17150,N_19563);
and U22633 (N_22633,N_18593,N_16598);
nand U22634 (N_22634,N_15885,N_19636);
nand U22635 (N_22635,N_15295,N_19767);
xnor U22636 (N_22636,N_18117,N_18786);
and U22637 (N_22637,N_19118,N_16221);
and U22638 (N_22638,N_16169,N_17532);
nand U22639 (N_22639,N_16040,N_19809);
nor U22640 (N_22640,N_17522,N_17292);
and U22641 (N_22641,N_18239,N_17722);
nand U22642 (N_22642,N_16828,N_18841);
xor U22643 (N_22643,N_18622,N_17718);
nand U22644 (N_22644,N_15489,N_16390);
and U22645 (N_22645,N_16769,N_16320);
and U22646 (N_22646,N_15085,N_16667);
or U22647 (N_22647,N_16583,N_15727);
nand U22648 (N_22648,N_18091,N_16693);
and U22649 (N_22649,N_16253,N_18550);
and U22650 (N_22650,N_15815,N_16708);
nor U22651 (N_22651,N_16501,N_18260);
nand U22652 (N_22652,N_18513,N_16703);
or U22653 (N_22653,N_17038,N_18600);
and U22654 (N_22654,N_19689,N_17056);
nor U22655 (N_22655,N_19309,N_17878);
xor U22656 (N_22656,N_15434,N_19680);
xor U22657 (N_22657,N_18152,N_19655);
nor U22658 (N_22658,N_17977,N_19463);
nand U22659 (N_22659,N_15324,N_18713);
xor U22660 (N_22660,N_15661,N_15242);
and U22661 (N_22661,N_18455,N_18942);
nand U22662 (N_22662,N_19424,N_19867);
nor U22663 (N_22663,N_15252,N_16343);
nor U22664 (N_22664,N_16714,N_15495);
nor U22665 (N_22665,N_17362,N_16396);
nor U22666 (N_22666,N_16620,N_18267);
nor U22667 (N_22667,N_18630,N_18253);
nor U22668 (N_22668,N_19521,N_15982);
nor U22669 (N_22669,N_17950,N_16143);
nor U22670 (N_22670,N_17795,N_18189);
nor U22671 (N_22671,N_16218,N_17109);
or U22672 (N_22672,N_19976,N_16965);
nand U22673 (N_22673,N_19402,N_18151);
nand U22674 (N_22674,N_18356,N_18558);
or U22675 (N_22675,N_15267,N_17637);
xnor U22676 (N_22676,N_16115,N_19761);
nand U22677 (N_22677,N_18698,N_16737);
xor U22678 (N_22678,N_18611,N_19424);
xor U22679 (N_22679,N_16709,N_16609);
or U22680 (N_22680,N_19633,N_16991);
xnor U22681 (N_22681,N_19453,N_19988);
nand U22682 (N_22682,N_19388,N_15857);
nand U22683 (N_22683,N_17089,N_18028);
and U22684 (N_22684,N_15631,N_18171);
or U22685 (N_22685,N_17027,N_15364);
xnor U22686 (N_22686,N_15314,N_16866);
and U22687 (N_22687,N_17342,N_16034);
and U22688 (N_22688,N_16217,N_17805);
xnor U22689 (N_22689,N_19922,N_18328);
xor U22690 (N_22690,N_19865,N_18347);
xor U22691 (N_22691,N_18314,N_16697);
or U22692 (N_22692,N_18649,N_17212);
xnor U22693 (N_22693,N_19003,N_18200);
xnor U22694 (N_22694,N_17050,N_16729);
nor U22695 (N_22695,N_15371,N_15877);
nor U22696 (N_22696,N_16544,N_15284);
xnor U22697 (N_22697,N_15898,N_19483);
nor U22698 (N_22698,N_18813,N_15428);
nor U22699 (N_22699,N_19872,N_18752);
nor U22700 (N_22700,N_15604,N_15299);
or U22701 (N_22701,N_16879,N_17190);
or U22702 (N_22702,N_15932,N_19626);
nand U22703 (N_22703,N_18739,N_16527);
nor U22704 (N_22704,N_16375,N_19701);
or U22705 (N_22705,N_18566,N_18913);
or U22706 (N_22706,N_17060,N_19046);
xor U22707 (N_22707,N_19895,N_18667);
nand U22708 (N_22708,N_17771,N_17097);
nor U22709 (N_22709,N_19092,N_15828);
nand U22710 (N_22710,N_18215,N_17916);
xnor U22711 (N_22711,N_15028,N_18222);
xnor U22712 (N_22712,N_18120,N_19807);
and U22713 (N_22713,N_16312,N_17079);
or U22714 (N_22714,N_18058,N_16586);
and U22715 (N_22715,N_15459,N_19443);
or U22716 (N_22716,N_18246,N_16879);
and U22717 (N_22717,N_19565,N_19006);
nand U22718 (N_22718,N_15042,N_16521);
or U22719 (N_22719,N_16939,N_17251);
or U22720 (N_22720,N_15138,N_19343);
or U22721 (N_22721,N_18361,N_17802);
or U22722 (N_22722,N_16081,N_17901);
xor U22723 (N_22723,N_15656,N_16180);
and U22724 (N_22724,N_16141,N_16479);
and U22725 (N_22725,N_15273,N_17247);
xor U22726 (N_22726,N_16494,N_17985);
nand U22727 (N_22727,N_15948,N_19022);
or U22728 (N_22728,N_19629,N_15505);
xor U22729 (N_22729,N_18992,N_17087);
nor U22730 (N_22730,N_16124,N_17620);
nand U22731 (N_22731,N_16521,N_18862);
and U22732 (N_22732,N_17102,N_15620);
nand U22733 (N_22733,N_16298,N_17029);
xnor U22734 (N_22734,N_17151,N_18936);
and U22735 (N_22735,N_15668,N_19877);
xor U22736 (N_22736,N_15307,N_18546);
xor U22737 (N_22737,N_15863,N_16772);
nand U22738 (N_22738,N_18520,N_15926);
or U22739 (N_22739,N_16783,N_15706);
xnor U22740 (N_22740,N_18067,N_16405);
nor U22741 (N_22741,N_15284,N_19076);
nand U22742 (N_22742,N_19250,N_16530);
xor U22743 (N_22743,N_15704,N_18468);
nor U22744 (N_22744,N_17670,N_18194);
or U22745 (N_22745,N_17250,N_16343);
and U22746 (N_22746,N_18153,N_19378);
or U22747 (N_22747,N_18841,N_17647);
nor U22748 (N_22748,N_15617,N_18466);
or U22749 (N_22749,N_16944,N_17851);
or U22750 (N_22750,N_17414,N_16797);
nand U22751 (N_22751,N_17184,N_16811);
nor U22752 (N_22752,N_19883,N_19971);
xnor U22753 (N_22753,N_17444,N_16313);
nor U22754 (N_22754,N_18540,N_19853);
or U22755 (N_22755,N_17224,N_15347);
xor U22756 (N_22756,N_15781,N_19672);
nand U22757 (N_22757,N_19961,N_16757);
or U22758 (N_22758,N_15138,N_19918);
nor U22759 (N_22759,N_15304,N_15192);
nor U22760 (N_22760,N_19154,N_19814);
or U22761 (N_22761,N_19392,N_17145);
nor U22762 (N_22762,N_19488,N_15827);
or U22763 (N_22763,N_15214,N_16745);
or U22764 (N_22764,N_18873,N_19420);
xor U22765 (N_22765,N_18150,N_19717);
xor U22766 (N_22766,N_19936,N_17293);
and U22767 (N_22767,N_19884,N_18197);
or U22768 (N_22768,N_16335,N_19672);
nand U22769 (N_22769,N_19886,N_16708);
or U22770 (N_22770,N_15973,N_17773);
nor U22771 (N_22771,N_16120,N_16900);
nand U22772 (N_22772,N_19427,N_16419);
and U22773 (N_22773,N_16711,N_16810);
nand U22774 (N_22774,N_15906,N_19545);
and U22775 (N_22775,N_16504,N_16664);
and U22776 (N_22776,N_15039,N_15325);
and U22777 (N_22777,N_15404,N_18283);
or U22778 (N_22778,N_15432,N_19269);
and U22779 (N_22779,N_17658,N_18114);
xor U22780 (N_22780,N_16486,N_16485);
nor U22781 (N_22781,N_16506,N_18020);
or U22782 (N_22782,N_15010,N_17396);
and U22783 (N_22783,N_15569,N_17198);
or U22784 (N_22784,N_19199,N_16512);
and U22785 (N_22785,N_18174,N_15032);
and U22786 (N_22786,N_18947,N_17428);
xnor U22787 (N_22787,N_16568,N_18070);
nor U22788 (N_22788,N_19836,N_19799);
xnor U22789 (N_22789,N_15298,N_19986);
nor U22790 (N_22790,N_16382,N_16553);
nor U22791 (N_22791,N_15763,N_16261);
xor U22792 (N_22792,N_15290,N_17534);
and U22793 (N_22793,N_16905,N_19775);
nor U22794 (N_22794,N_15099,N_19700);
and U22795 (N_22795,N_19135,N_15756);
nor U22796 (N_22796,N_19769,N_18122);
nand U22797 (N_22797,N_15007,N_16420);
and U22798 (N_22798,N_19769,N_18534);
or U22799 (N_22799,N_15569,N_15600);
and U22800 (N_22800,N_15261,N_18270);
xnor U22801 (N_22801,N_19575,N_19302);
nor U22802 (N_22802,N_17268,N_17691);
and U22803 (N_22803,N_17242,N_18301);
xor U22804 (N_22804,N_16339,N_18896);
nand U22805 (N_22805,N_16161,N_17928);
nor U22806 (N_22806,N_15469,N_16363);
nand U22807 (N_22807,N_19765,N_15919);
or U22808 (N_22808,N_16935,N_17774);
xnor U22809 (N_22809,N_16900,N_19187);
nand U22810 (N_22810,N_15654,N_17179);
xor U22811 (N_22811,N_19044,N_19087);
xor U22812 (N_22812,N_19691,N_19481);
or U22813 (N_22813,N_19851,N_15032);
nor U22814 (N_22814,N_17319,N_19008);
nor U22815 (N_22815,N_19882,N_18374);
and U22816 (N_22816,N_19825,N_18345);
or U22817 (N_22817,N_15337,N_19071);
xor U22818 (N_22818,N_16833,N_16857);
nor U22819 (N_22819,N_17276,N_18815);
and U22820 (N_22820,N_19890,N_18193);
and U22821 (N_22821,N_15248,N_15055);
xnor U22822 (N_22822,N_19307,N_18520);
and U22823 (N_22823,N_17209,N_17662);
xor U22824 (N_22824,N_17388,N_18681);
and U22825 (N_22825,N_18460,N_15859);
xor U22826 (N_22826,N_16450,N_19136);
nor U22827 (N_22827,N_19514,N_17210);
and U22828 (N_22828,N_19099,N_15892);
nor U22829 (N_22829,N_16344,N_18649);
or U22830 (N_22830,N_16998,N_18001);
xnor U22831 (N_22831,N_18260,N_15455);
nor U22832 (N_22832,N_18211,N_17913);
nor U22833 (N_22833,N_18554,N_17813);
nand U22834 (N_22834,N_16372,N_15619);
nand U22835 (N_22835,N_19972,N_19833);
nor U22836 (N_22836,N_17416,N_19040);
and U22837 (N_22837,N_17265,N_18075);
nor U22838 (N_22838,N_15642,N_18995);
nand U22839 (N_22839,N_15921,N_18990);
or U22840 (N_22840,N_19709,N_17549);
xnor U22841 (N_22841,N_18836,N_17845);
and U22842 (N_22842,N_18635,N_18094);
and U22843 (N_22843,N_16485,N_19308);
nor U22844 (N_22844,N_16521,N_17590);
and U22845 (N_22845,N_17464,N_18170);
and U22846 (N_22846,N_18680,N_19875);
nor U22847 (N_22847,N_16182,N_19301);
and U22848 (N_22848,N_18084,N_16337);
xor U22849 (N_22849,N_15917,N_19371);
xnor U22850 (N_22850,N_18987,N_18199);
and U22851 (N_22851,N_15452,N_16512);
xor U22852 (N_22852,N_15504,N_17283);
nand U22853 (N_22853,N_15289,N_18270);
nand U22854 (N_22854,N_16353,N_19754);
xor U22855 (N_22855,N_16965,N_15565);
or U22856 (N_22856,N_16393,N_19638);
xor U22857 (N_22857,N_16193,N_16430);
and U22858 (N_22858,N_18523,N_19408);
and U22859 (N_22859,N_17856,N_19074);
nor U22860 (N_22860,N_15921,N_18489);
and U22861 (N_22861,N_18318,N_19118);
nand U22862 (N_22862,N_18322,N_18079);
xnor U22863 (N_22863,N_18900,N_17800);
or U22864 (N_22864,N_15925,N_19679);
or U22865 (N_22865,N_16550,N_18671);
nand U22866 (N_22866,N_15371,N_16103);
or U22867 (N_22867,N_19865,N_15237);
xnor U22868 (N_22868,N_18896,N_19992);
nor U22869 (N_22869,N_19493,N_17593);
xnor U22870 (N_22870,N_18482,N_17510);
xnor U22871 (N_22871,N_18163,N_16757);
nand U22872 (N_22872,N_19931,N_15410);
or U22873 (N_22873,N_16357,N_15391);
nand U22874 (N_22874,N_18840,N_15481);
nor U22875 (N_22875,N_18422,N_17823);
nor U22876 (N_22876,N_15915,N_15179);
or U22877 (N_22877,N_18334,N_16929);
xor U22878 (N_22878,N_18561,N_18065);
nor U22879 (N_22879,N_18201,N_17178);
nand U22880 (N_22880,N_19678,N_18555);
and U22881 (N_22881,N_18633,N_16298);
xor U22882 (N_22882,N_17239,N_17636);
and U22883 (N_22883,N_16788,N_18828);
and U22884 (N_22884,N_17044,N_18655);
nand U22885 (N_22885,N_16308,N_18455);
xnor U22886 (N_22886,N_18440,N_18438);
nand U22887 (N_22887,N_15012,N_19244);
and U22888 (N_22888,N_17624,N_19757);
nand U22889 (N_22889,N_19786,N_17119);
and U22890 (N_22890,N_16950,N_18030);
nand U22891 (N_22891,N_19619,N_16047);
nor U22892 (N_22892,N_19229,N_16130);
nor U22893 (N_22893,N_18386,N_18689);
or U22894 (N_22894,N_17977,N_19579);
nand U22895 (N_22895,N_15500,N_17808);
xor U22896 (N_22896,N_15786,N_16954);
or U22897 (N_22897,N_17098,N_17388);
nor U22898 (N_22898,N_15268,N_18876);
nor U22899 (N_22899,N_16264,N_18811);
or U22900 (N_22900,N_17512,N_17904);
and U22901 (N_22901,N_19561,N_19737);
and U22902 (N_22902,N_17490,N_18352);
nor U22903 (N_22903,N_19990,N_18486);
xor U22904 (N_22904,N_15861,N_17058);
or U22905 (N_22905,N_18310,N_18967);
or U22906 (N_22906,N_16599,N_18745);
or U22907 (N_22907,N_17978,N_18874);
or U22908 (N_22908,N_15796,N_19072);
and U22909 (N_22909,N_15462,N_15287);
nor U22910 (N_22910,N_18557,N_15548);
nand U22911 (N_22911,N_16355,N_15552);
nor U22912 (N_22912,N_15628,N_18561);
nor U22913 (N_22913,N_17083,N_15384);
and U22914 (N_22914,N_18602,N_19053);
nand U22915 (N_22915,N_16990,N_19017);
nor U22916 (N_22916,N_17392,N_19976);
nor U22917 (N_22917,N_16931,N_15586);
nand U22918 (N_22918,N_15833,N_19540);
or U22919 (N_22919,N_18702,N_15080);
and U22920 (N_22920,N_15865,N_17497);
xor U22921 (N_22921,N_17338,N_15817);
and U22922 (N_22922,N_19816,N_18355);
or U22923 (N_22923,N_18079,N_18171);
and U22924 (N_22924,N_15811,N_18902);
xnor U22925 (N_22925,N_16437,N_18225);
nand U22926 (N_22926,N_18306,N_15375);
nor U22927 (N_22927,N_18440,N_16459);
or U22928 (N_22928,N_18516,N_18323);
and U22929 (N_22929,N_15774,N_18399);
xor U22930 (N_22930,N_18288,N_17959);
xor U22931 (N_22931,N_15634,N_16986);
nand U22932 (N_22932,N_17379,N_18797);
nor U22933 (N_22933,N_19000,N_19871);
or U22934 (N_22934,N_17483,N_19566);
and U22935 (N_22935,N_16155,N_16136);
or U22936 (N_22936,N_18414,N_16363);
and U22937 (N_22937,N_15343,N_18345);
xnor U22938 (N_22938,N_19243,N_18431);
and U22939 (N_22939,N_19792,N_19591);
xor U22940 (N_22940,N_18536,N_16496);
xor U22941 (N_22941,N_15852,N_18101);
and U22942 (N_22942,N_15260,N_19271);
and U22943 (N_22943,N_17406,N_17233);
nand U22944 (N_22944,N_19009,N_16717);
or U22945 (N_22945,N_18714,N_19287);
nor U22946 (N_22946,N_17176,N_16757);
or U22947 (N_22947,N_15294,N_18843);
xnor U22948 (N_22948,N_17247,N_19523);
nor U22949 (N_22949,N_15610,N_19474);
xor U22950 (N_22950,N_16800,N_19574);
xnor U22951 (N_22951,N_15314,N_18261);
nor U22952 (N_22952,N_15064,N_19727);
xor U22953 (N_22953,N_17147,N_18664);
or U22954 (N_22954,N_18020,N_18087);
nand U22955 (N_22955,N_15212,N_15036);
and U22956 (N_22956,N_16633,N_16402);
and U22957 (N_22957,N_19824,N_17944);
nand U22958 (N_22958,N_19990,N_16635);
nand U22959 (N_22959,N_18358,N_17304);
xnor U22960 (N_22960,N_15443,N_19395);
nor U22961 (N_22961,N_16426,N_16387);
and U22962 (N_22962,N_17081,N_15294);
xor U22963 (N_22963,N_17262,N_15135);
and U22964 (N_22964,N_16940,N_18229);
nor U22965 (N_22965,N_16881,N_17106);
or U22966 (N_22966,N_16145,N_16172);
or U22967 (N_22967,N_17161,N_15687);
nand U22968 (N_22968,N_16540,N_17831);
and U22969 (N_22969,N_16585,N_18813);
nand U22970 (N_22970,N_16634,N_18868);
nand U22971 (N_22971,N_19337,N_16526);
and U22972 (N_22972,N_17909,N_18773);
xor U22973 (N_22973,N_16814,N_19954);
or U22974 (N_22974,N_15331,N_15185);
xnor U22975 (N_22975,N_19064,N_16906);
xnor U22976 (N_22976,N_15886,N_18176);
nand U22977 (N_22977,N_16952,N_19265);
nand U22978 (N_22978,N_15641,N_19159);
nor U22979 (N_22979,N_15016,N_18455);
and U22980 (N_22980,N_18749,N_19553);
nand U22981 (N_22981,N_16667,N_19939);
xor U22982 (N_22982,N_18243,N_19192);
nor U22983 (N_22983,N_16598,N_17704);
xnor U22984 (N_22984,N_17713,N_16690);
and U22985 (N_22985,N_15688,N_19221);
xnor U22986 (N_22986,N_17040,N_18973);
and U22987 (N_22987,N_18568,N_15148);
and U22988 (N_22988,N_17021,N_16617);
xor U22989 (N_22989,N_17555,N_19148);
nor U22990 (N_22990,N_16306,N_19168);
nand U22991 (N_22991,N_15134,N_18252);
and U22992 (N_22992,N_16351,N_16074);
and U22993 (N_22993,N_18141,N_17487);
or U22994 (N_22994,N_16464,N_18006);
nand U22995 (N_22995,N_18639,N_19719);
nand U22996 (N_22996,N_15040,N_15104);
xor U22997 (N_22997,N_15806,N_15372);
xor U22998 (N_22998,N_18396,N_17373);
or U22999 (N_22999,N_17295,N_17994);
nand U23000 (N_23000,N_19473,N_18447);
or U23001 (N_23001,N_19793,N_15323);
nand U23002 (N_23002,N_16204,N_18382);
nand U23003 (N_23003,N_18814,N_17863);
nand U23004 (N_23004,N_17018,N_18760);
xnor U23005 (N_23005,N_18172,N_16425);
nor U23006 (N_23006,N_16358,N_18463);
nand U23007 (N_23007,N_15309,N_16830);
nor U23008 (N_23008,N_18821,N_17853);
nor U23009 (N_23009,N_18372,N_18541);
and U23010 (N_23010,N_15517,N_19302);
and U23011 (N_23011,N_17526,N_18139);
or U23012 (N_23012,N_19148,N_18384);
or U23013 (N_23013,N_16180,N_19434);
nor U23014 (N_23014,N_18468,N_19996);
xor U23015 (N_23015,N_17275,N_18237);
nor U23016 (N_23016,N_16450,N_17767);
or U23017 (N_23017,N_17249,N_19816);
nand U23018 (N_23018,N_18883,N_19634);
and U23019 (N_23019,N_19042,N_15894);
nand U23020 (N_23020,N_17261,N_15184);
xnor U23021 (N_23021,N_19055,N_16129);
and U23022 (N_23022,N_15613,N_19460);
or U23023 (N_23023,N_15368,N_18140);
or U23024 (N_23024,N_15826,N_19456);
xnor U23025 (N_23025,N_16768,N_17515);
and U23026 (N_23026,N_19860,N_17290);
and U23027 (N_23027,N_17353,N_19408);
xor U23028 (N_23028,N_15663,N_19049);
and U23029 (N_23029,N_17531,N_15041);
nand U23030 (N_23030,N_16547,N_15998);
and U23031 (N_23031,N_18379,N_16942);
xor U23032 (N_23032,N_18777,N_19037);
or U23033 (N_23033,N_17216,N_16298);
nor U23034 (N_23034,N_15882,N_17059);
nor U23035 (N_23035,N_18511,N_18515);
and U23036 (N_23036,N_16808,N_19888);
or U23037 (N_23037,N_15418,N_15519);
and U23038 (N_23038,N_15594,N_16353);
nor U23039 (N_23039,N_19996,N_19600);
nor U23040 (N_23040,N_15068,N_16940);
nor U23041 (N_23041,N_15750,N_19614);
and U23042 (N_23042,N_15167,N_19486);
and U23043 (N_23043,N_16850,N_18585);
xnor U23044 (N_23044,N_18278,N_17348);
and U23045 (N_23045,N_17950,N_16413);
nor U23046 (N_23046,N_18979,N_15454);
xnor U23047 (N_23047,N_17010,N_17499);
xor U23048 (N_23048,N_16397,N_16793);
nor U23049 (N_23049,N_19640,N_17932);
or U23050 (N_23050,N_19677,N_17533);
xnor U23051 (N_23051,N_17768,N_18529);
and U23052 (N_23052,N_15228,N_15814);
and U23053 (N_23053,N_15517,N_18921);
xnor U23054 (N_23054,N_16937,N_16369);
nand U23055 (N_23055,N_19781,N_15124);
or U23056 (N_23056,N_19020,N_17478);
or U23057 (N_23057,N_19290,N_16303);
nor U23058 (N_23058,N_16888,N_19191);
or U23059 (N_23059,N_19334,N_19213);
or U23060 (N_23060,N_17940,N_19074);
nor U23061 (N_23061,N_15087,N_15259);
and U23062 (N_23062,N_18502,N_19261);
xor U23063 (N_23063,N_15317,N_18356);
or U23064 (N_23064,N_19111,N_17532);
nor U23065 (N_23065,N_15037,N_18336);
and U23066 (N_23066,N_17153,N_17090);
and U23067 (N_23067,N_15160,N_19037);
and U23068 (N_23068,N_15319,N_19100);
nand U23069 (N_23069,N_17224,N_18157);
nand U23070 (N_23070,N_18128,N_15277);
and U23071 (N_23071,N_19957,N_15973);
xnor U23072 (N_23072,N_15688,N_19504);
xnor U23073 (N_23073,N_19311,N_17488);
nor U23074 (N_23074,N_18438,N_19866);
nand U23075 (N_23075,N_16247,N_18066);
nor U23076 (N_23076,N_19078,N_15238);
or U23077 (N_23077,N_18264,N_16506);
and U23078 (N_23078,N_15947,N_18088);
nand U23079 (N_23079,N_18709,N_16914);
nor U23080 (N_23080,N_17168,N_18930);
and U23081 (N_23081,N_15622,N_16698);
and U23082 (N_23082,N_16585,N_19002);
or U23083 (N_23083,N_18881,N_18192);
and U23084 (N_23084,N_17160,N_15432);
nand U23085 (N_23085,N_17426,N_18713);
nand U23086 (N_23086,N_16795,N_15887);
xnor U23087 (N_23087,N_17715,N_18239);
nor U23088 (N_23088,N_16496,N_19489);
and U23089 (N_23089,N_17239,N_17660);
xor U23090 (N_23090,N_18524,N_16484);
or U23091 (N_23091,N_18006,N_19203);
nand U23092 (N_23092,N_19103,N_17693);
nand U23093 (N_23093,N_17459,N_17120);
xor U23094 (N_23094,N_16852,N_17244);
or U23095 (N_23095,N_16662,N_17299);
xor U23096 (N_23096,N_15885,N_15606);
nor U23097 (N_23097,N_17720,N_17480);
nor U23098 (N_23098,N_17253,N_17745);
xnor U23099 (N_23099,N_19312,N_15280);
and U23100 (N_23100,N_18111,N_18407);
nand U23101 (N_23101,N_15116,N_19026);
or U23102 (N_23102,N_18153,N_15781);
or U23103 (N_23103,N_16451,N_19863);
and U23104 (N_23104,N_19290,N_19498);
xor U23105 (N_23105,N_18835,N_19390);
nor U23106 (N_23106,N_18379,N_15587);
and U23107 (N_23107,N_16607,N_19671);
and U23108 (N_23108,N_16731,N_18103);
and U23109 (N_23109,N_16770,N_19326);
xor U23110 (N_23110,N_15455,N_19937);
nor U23111 (N_23111,N_19000,N_19845);
or U23112 (N_23112,N_16131,N_17861);
nor U23113 (N_23113,N_18318,N_19786);
and U23114 (N_23114,N_15458,N_18712);
or U23115 (N_23115,N_17436,N_17677);
nor U23116 (N_23116,N_16888,N_19841);
xnor U23117 (N_23117,N_16662,N_17259);
nor U23118 (N_23118,N_17039,N_15892);
xnor U23119 (N_23119,N_17454,N_16097);
nand U23120 (N_23120,N_16382,N_17629);
xnor U23121 (N_23121,N_18342,N_19951);
nand U23122 (N_23122,N_15692,N_18709);
or U23123 (N_23123,N_15374,N_19168);
and U23124 (N_23124,N_15196,N_19971);
or U23125 (N_23125,N_17990,N_16703);
and U23126 (N_23126,N_16313,N_15568);
and U23127 (N_23127,N_17906,N_18712);
nor U23128 (N_23128,N_16890,N_19221);
nand U23129 (N_23129,N_16173,N_15815);
nor U23130 (N_23130,N_17937,N_16824);
nand U23131 (N_23131,N_16257,N_18570);
and U23132 (N_23132,N_18384,N_15238);
and U23133 (N_23133,N_18544,N_17641);
or U23134 (N_23134,N_15679,N_16857);
nand U23135 (N_23135,N_15410,N_19729);
xor U23136 (N_23136,N_15997,N_19762);
xnor U23137 (N_23137,N_15196,N_17079);
nand U23138 (N_23138,N_18389,N_17805);
or U23139 (N_23139,N_18001,N_15470);
nand U23140 (N_23140,N_19587,N_18832);
xnor U23141 (N_23141,N_16274,N_17532);
and U23142 (N_23142,N_19187,N_15001);
and U23143 (N_23143,N_16586,N_16873);
nand U23144 (N_23144,N_17728,N_19060);
nand U23145 (N_23145,N_19138,N_15409);
and U23146 (N_23146,N_16652,N_15123);
nand U23147 (N_23147,N_15824,N_17380);
or U23148 (N_23148,N_19871,N_19069);
xor U23149 (N_23149,N_17115,N_15921);
nand U23150 (N_23150,N_15335,N_17833);
and U23151 (N_23151,N_17104,N_15733);
nor U23152 (N_23152,N_15341,N_18013);
xnor U23153 (N_23153,N_15734,N_19437);
xnor U23154 (N_23154,N_16177,N_19574);
and U23155 (N_23155,N_19552,N_17225);
or U23156 (N_23156,N_15221,N_16223);
or U23157 (N_23157,N_16778,N_15558);
nand U23158 (N_23158,N_17583,N_18566);
and U23159 (N_23159,N_17953,N_19048);
xnor U23160 (N_23160,N_17045,N_16534);
and U23161 (N_23161,N_18714,N_17823);
and U23162 (N_23162,N_17596,N_19285);
xor U23163 (N_23163,N_19120,N_17810);
and U23164 (N_23164,N_19958,N_17230);
and U23165 (N_23165,N_15182,N_18222);
nor U23166 (N_23166,N_17895,N_16815);
nand U23167 (N_23167,N_17500,N_16258);
xor U23168 (N_23168,N_17808,N_16704);
and U23169 (N_23169,N_19293,N_19313);
and U23170 (N_23170,N_19280,N_17383);
nor U23171 (N_23171,N_18228,N_15826);
nor U23172 (N_23172,N_17734,N_17650);
nor U23173 (N_23173,N_17295,N_18283);
or U23174 (N_23174,N_15926,N_17447);
nor U23175 (N_23175,N_17668,N_16671);
nand U23176 (N_23176,N_15083,N_18215);
or U23177 (N_23177,N_17688,N_15288);
xor U23178 (N_23178,N_16185,N_16626);
nor U23179 (N_23179,N_15763,N_18294);
and U23180 (N_23180,N_19144,N_18347);
nand U23181 (N_23181,N_16006,N_16214);
nor U23182 (N_23182,N_17255,N_15462);
or U23183 (N_23183,N_17890,N_15743);
nor U23184 (N_23184,N_17610,N_17975);
and U23185 (N_23185,N_16283,N_17180);
nand U23186 (N_23186,N_18095,N_18717);
xor U23187 (N_23187,N_16296,N_17223);
nor U23188 (N_23188,N_15029,N_15413);
or U23189 (N_23189,N_15629,N_18612);
xnor U23190 (N_23190,N_18032,N_16625);
nand U23191 (N_23191,N_18267,N_19478);
and U23192 (N_23192,N_17686,N_19994);
xor U23193 (N_23193,N_18252,N_15295);
or U23194 (N_23194,N_18795,N_16874);
nor U23195 (N_23195,N_19712,N_15824);
or U23196 (N_23196,N_19144,N_16843);
nor U23197 (N_23197,N_16651,N_19186);
xor U23198 (N_23198,N_16152,N_18656);
nor U23199 (N_23199,N_18592,N_19412);
nand U23200 (N_23200,N_16877,N_19427);
or U23201 (N_23201,N_15038,N_19714);
or U23202 (N_23202,N_19140,N_19862);
nand U23203 (N_23203,N_16005,N_18174);
and U23204 (N_23204,N_19788,N_15058);
and U23205 (N_23205,N_19027,N_16373);
nor U23206 (N_23206,N_16783,N_19034);
xnor U23207 (N_23207,N_18091,N_18905);
and U23208 (N_23208,N_16046,N_19189);
nand U23209 (N_23209,N_15466,N_17254);
nor U23210 (N_23210,N_16463,N_17919);
nor U23211 (N_23211,N_18868,N_18978);
and U23212 (N_23212,N_15434,N_19013);
xor U23213 (N_23213,N_17369,N_17110);
or U23214 (N_23214,N_15559,N_17450);
and U23215 (N_23215,N_15107,N_18559);
or U23216 (N_23216,N_16968,N_19386);
nor U23217 (N_23217,N_15678,N_18944);
nand U23218 (N_23218,N_17007,N_17843);
nor U23219 (N_23219,N_17679,N_18356);
nor U23220 (N_23220,N_15561,N_19456);
xor U23221 (N_23221,N_16810,N_15861);
nor U23222 (N_23222,N_19467,N_19652);
nor U23223 (N_23223,N_19104,N_16893);
or U23224 (N_23224,N_18553,N_19474);
nor U23225 (N_23225,N_18574,N_16759);
nor U23226 (N_23226,N_17107,N_16306);
nor U23227 (N_23227,N_19755,N_17496);
xnor U23228 (N_23228,N_19745,N_19056);
or U23229 (N_23229,N_17607,N_19554);
nand U23230 (N_23230,N_18726,N_16556);
or U23231 (N_23231,N_15040,N_15927);
and U23232 (N_23232,N_18263,N_16978);
nor U23233 (N_23233,N_18597,N_15104);
nand U23234 (N_23234,N_15450,N_18868);
xor U23235 (N_23235,N_19821,N_19697);
nand U23236 (N_23236,N_19088,N_16234);
and U23237 (N_23237,N_17814,N_18918);
and U23238 (N_23238,N_18096,N_16920);
nand U23239 (N_23239,N_19743,N_15736);
or U23240 (N_23240,N_17846,N_18704);
nand U23241 (N_23241,N_17660,N_19472);
or U23242 (N_23242,N_15203,N_15392);
xnor U23243 (N_23243,N_19632,N_17791);
and U23244 (N_23244,N_16548,N_16456);
nand U23245 (N_23245,N_16392,N_16265);
and U23246 (N_23246,N_19014,N_18971);
nor U23247 (N_23247,N_16338,N_16622);
nor U23248 (N_23248,N_16725,N_17452);
xor U23249 (N_23249,N_16464,N_16812);
xor U23250 (N_23250,N_19991,N_16005);
nand U23251 (N_23251,N_18460,N_18850);
nand U23252 (N_23252,N_19954,N_15322);
nand U23253 (N_23253,N_16364,N_19592);
nor U23254 (N_23254,N_18211,N_18513);
nand U23255 (N_23255,N_17366,N_17322);
and U23256 (N_23256,N_18894,N_19692);
nor U23257 (N_23257,N_19501,N_15606);
nor U23258 (N_23258,N_19236,N_15875);
and U23259 (N_23259,N_19983,N_17706);
nor U23260 (N_23260,N_15501,N_19354);
xor U23261 (N_23261,N_18517,N_16856);
nor U23262 (N_23262,N_19201,N_16356);
nand U23263 (N_23263,N_19397,N_17082);
and U23264 (N_23264,N_17925,N_17535);
nand U23265 (N_23265,N_18789,N_19988);
nor U23266 (N_23266,N_19854,N_15697);
nand U23267 (N_23267,N_18963,N_16135);
or U23268 (N_23268,N_16488,N_18633);
xor U23269 (N_23269,N_15139,N_19971);
nor U23270 (N_23270,N_18439,N_15871);
nor U23271 (N_23271,N_19701,N_15737);
xnor U23272 (N_23272,N_15739,N_17030);
or U23273 (N_23273,N_15109,N_17953);
and U23274 (N_23274,N_18550,N_15211);
nor U23275 (N_23275,N_17589,N_19176);
xor U23276 (N_23276,N_18490,N_16260);
or U23277 (N_23277,N_17225,N_18638);
and U23278 (N_23278,N_15089,N_16088);
nand U23279 (N_23279,N_16626,N_17387);
and U23280 (N_23280,N_16643,N_19632);
nor U23281 (N_23281,N_16304,N_19614);
xor U23282 (N_23282,N_16104,N_19039);
and U23283 (N_23283,N_17104,N_19035);
nand U23284 (N_23284,N_19944,N_17884);
nand U23285 (N_23285,N_16055,N_19174);
and U23286 (N_23286,N_15048,N_17901);
xor U23287 (N_23287,N_15169,N_15362);
and U23288 (N_23288,N_19630,N_15198);
xor U23289 (N_23289,N_15134,N_18802);
nor U23290 (N_23290,N_15585,N_19701);
and U23291 (N_23291,N_16585,N_16516);
nand U23292 (N_23292,N_17237,N_17294);
xor U23293 (N_23293,N_18825,N_17254);
or U23294 (N_23294,N_18594,N_17711);
nand U23295 (N_23295,N_19950,N_17616);
nor U23296 (N_23296,N_19001,N_19784);
or U23297 (N_23297,N_18611,N_17651);
or U23298 (N_23298,N_15267,N_18440);
nor U23299 (N_23299,N_16111,N_16570);
or U23300 (N_23300,N_19383,N_19462);
nand U23301 (N_23301,N_16458,N_15209);
or U23302 (N_23302,N_17714,N_15141);
and U23303 (N_23303,N_16894,N_15274);
nand U23304 (N_23304,N_19176,N_19347);
xnor U23305 (N_23305,N_18520,N_15011);
xnor U23306 (N_23306,N_19180,N_17870);
and U23307 (N_23307,N_19497,N_19222);
and U23308 (N_23308,N_18445,N_19019);
xor U23309 (N_23309,N_17234,N_17491);
and U23310 (N_23310,N_16855,N_18748);
xor U23311 (N_23311,N_18171,N_19461);
nand U23312 (N_23312,N_19438,N_19912);
nand U23313 (N_23313,N_16777,N_16146);
and U23314 (N_23314,N_18433,N_16719);
and U23315 (N_23315,N_17764,N_15404);
or U23316 (N_23316,N_16579,N_18678);
and U23317 (N_23317,N_17602,N_17767);
xor U23318 (N_23318,N_16333,N_18656);
xor U23319 (N_23319,N_19195,N_16421);
nor U23320 (N_23320,N_19931,N_19577);
nand U23321 (N_23321,N_17930,N_16475);
xnor U23322 (N_23322,N_18580,N_17959);
or U23323 (N_23323,N_19078,N_15207);
or U23324 (N_23324,N_16732,N_15580);
nor U23325 (N_23325,N_18937,N_19387);
or U23326 (N_23326,N_19163,N_18772);
xnor U23327 (N_23327,N_18927,N_15288);
xor U23328 (N_23328,N_18946,N_18006);
xor U23329 (N_23329,N_17111,N_19347);
or U23330 (N_23330,N_16727,N_19004);
nand U23331 (N_23331,N_15093,N_16797);
and U23332 (N_23332,N_19986,N_15816);
and U23333 (N_23333,N_19383,N_18851);
and U23334 (N_23334,N_19483,N_17735);
xnor U23335 (N_23335,N_17693,N_15833);
nor U23336 (N_23336,N_19732,N_18250);
and U23337 (N_23337,N_15475,N_15935);
nor U23338 (N_23338,N_18014,N_15963);
nand U23339 (N_23339,N_19838,N_18462);
nor U23340 (N_23340,N_18075,N_17289);
or U23341 (N_23341,N_18137,N_18751);
and U23342 (N_23342,N_18678,N_15357);
or U23343 (N_23343,N_17820,N_16566);
nand U23344 (N_23344,N_15635,N_15641);
and U23345 (N_23345,N_19932,N_16204);
xnor U23346 (N_23346,N_17786,N_18426);
xnor U23347 (N_23347,N_15592,N_17169);
xnor U23348 (N_23348,N_15401,N_17437);
xor U23349 (N_23349,N_17120,N_17867);
nor U23350 (N_23350,N_18385,N_17982);
xnor U23351 (N_23351,N_17919,N_19282);
or U23352 (N_23352,N_19197,N_18535);
nand U23353 (N_23353,N_16276,N_19763);
xor U23354 (N_23354,N_17947,N_17106);
or U23355 (N_23355,N_15984,N_16245);
nor U23356 (N_23356,N_16601,N_16734);
or U23357 (N_23357,N_16557,N_15668);
nor U23358 (N_23358,N_15835,N_16686);
or U23359 (N_23359,N_15238,N_15431);
and U23360 (N_23360,N_15181,N_18128);
nand U23361 (N_23361,N_16998,N_19811);
or U23362 (N_23362,N_17864,N_18720);
nor U23363 (N_23363,N_17997,N_19358);
nor U23364 (N_23364,N_16255,N_15233);
and U23365 (N_23365,N_18242,N_18355);
xor U23366 (N_23366,N_18614,N_15833);
or U23367 (N_23367,N_17729,N_17664);
nor U23368 (N_23368,N_17761,N_16258);
and U23369 (N_23369,N_17627,N_19680);
or U23370 (N_23370,N_15028,N_16681);
nand U23371 (N_23371,N_17738,N_19195);
xor U23372 (N_23372,N_18496,N_17152);
and U23373 (N_23373,N_19788,N_17390);
and U23374 (N_23374,N_19042,N_17111);
and U23375 (N_23375,N_19521,N_17305);
xor U23376 (N_23376,N_15076,N_17724);
or U23377 (N_23377,N_16827,N_16857);
xnor U23378 (N_23378,N_17664,N_17953);
nor U23379 (N_23379,N_17412,N_19108);
nor U23380 (N_23380,N_18240,N_15377);
and U23381 (N_23381,N_19106,N_19403);
nand U23382 (N_23382,N_17329,N_17660);
and U23383 (N_23383,N_17347,N_19282);
nand U23384 (N_23384,N_17740,N_17562);
nand U23385 (N_23385,N_19817,N_16743);
xor U23386 (N_23386,N_16821,N_19160);
and U23387 (N_23387,N_19561,N_15292);
nand U23388 (N_23388,N_18284,N_19821);
xor U23389 (N_23389,N_15500,N_19246);
nand U23390 (N_23390,N_19653,N_16120);
xnor U23391 (N_23391,N_19585,N_19036);
or U23392 (N_23392,N_18577,N_18213);
nor U23393 (N_23393,N_17413,N_16428);
or U23394 (N_23394,N_17337,N_17058);
and U23395 (N_23395,N_17745,N_15397);
and U23396 (N_23396,N_16351,N_18347);
and U23397 (N_23397,N_15559,N_18453);
nand U23398 (N_23398,N_15375,N_17148);
or U23399 (N_23399,N_18195,N_19530);
nand U23400 (N_23400,N_19876,N_19995);
xnor U23401 (N_23401,N_15731,N_19963);
nor U23402 (N_23402,N_17526,N_19775);
xor U23403 (N_23403,N_19542,N_16998);
xnor U23404 (N_23404,N_19698,N_16332);
xnor U23405 (N_23405,N_15054,N_18874);
xor U23406 (N_23406,N_19863,N_19512);
and U23407 (N_23407,N_19523,N_19980);
nor U23408 (N_23408,N_17639,N_17411);
and U23409 (N_23409,N_15702,N_16812);
and U23410 (N_23410,N_18514,N_15829);
or U23411 (N_23411,N_19334,N_19865);
and U23412 (N_23412,N_15652,N_19633);
xor U23413 (N_23413,N_19994,N_16884);
or U23414 (N_23414,N_16596,N_18489);
and U23415 (N_23415,N_19499,N_17708);
and U23416 (N_23416,N_17252,N_19607);
and U23417 (N_23417,N_18979,N_19105);
and U23418 (N_23418,N_15052,N_16704);
nand U23419 (N_23419,N_18425,N_15859);
and U23420 (N_23420,N_16829,N_16472);
and U23421 (N_23421,N_16108,N_17857);
and U23422 (N_23422,N_16362,N_18185);
and U23423 (N_23423,N_16846,N_17898);
nand U23424 (N_23424,N_16173,N_16174);
xnor U23425 (N_23425,N_16309,N_17063);
nor U23426 (N_23426,N_15840,N_18767);
nor U23427 (N_23427,N_15454,N_15744);
and U23428 (N_23428,N_16439,N_19727);
or U23429 (N_23429,N_19284,N_18825);
nand U23430 (N_23430,N_19031,N_17794);
xnor U23431 (N_23431,N_18302,N_19124);
nor U23432 (N_23432,N_17232,N_17259);
xor U23433 (N_23433,N_15524,N_16318);
or U23434 (N_23434,N_17059,N_15356);
and U23435 (N_23435,N_17592,N_18960);
xnor U23436 (N_23436,N_19245,N_16989);
xor U23437 (N_23437,N_18646,N_18542);
and U23438 (N_23438,N_19342,N_19531);
or U23439 (N_23439,N_18061,N_17340);
or U23440 (N_23440,N_19411,N_18339);
and U23441 (N_23441,N_16083,N_15443);
nor U23442 (N_23442,N_17582,N_19750);
nor U23443 (N_23443,N_16059,N_15103);
and U23444 (N_23444,N_18885,N_19770);
and U23445 (N_23445,N_16630,N_16976);
or U23446 (N_23446,N_17194,N_15475);
nor U23447 (N_23447,N_19914,N_17865);
or U23448 (N_23448,N_18352,N_15733);
or U23449 (N_23449,N_17631,N_15273);
xor U23450 (N_23450,N_16763,N_15052);
xnor U23451 (N_23451,N_17626,N_15613);
nand U23452 (N_23452,N_16530,N_16605);
xor U23453 (N_23453,N_17432,N_16451);
and U23454 (N_23454,N_16061,N_15919);
nand U23455 (N_23455,N_15179,N_17342);
nand U23456 (N_23456,N_17652,N_15914);
and U23457 (N_23457,N_16994,N_19644);
and U23458 (N_23458,N_17720,N_16738);
nand U23459 (N_23459,N_17958,N_19673);
and U23460 (N_23460,N_15719,N_16852);
and U23461 (N_23461,N_17501,N_15694);
nor U23462 (N_23462,N_19014,N_19804);
xnor U23463 (N_23463,N_15506,N_18705);
xor U23464 (N_23464,N_15015,N_16051);
nand U23465 (N_23465,N_18319,N_19577);
nor U23466 (N_23466,N_19237,N_17428);
or U23467 (N_23467,N_17041,N_15890);
nor U23468 (N_23468,N_17527,N_15120);
nor U23469 (N_23469,N_16643,N_18556);
nor U23470 (N_23470,N_18129,N_19952);
nand U23471 (N_23471,N_16716,N_19660);
and U23472 (N_23472,N_17636,N_15019);
nor U23473 (N_23473,N_16846,N_17206);
nand U23474 (N_23474,N_16701,N_16979);
nor U23475 (N_23475,N_15593,N_15556);
and U23476 (N_23476,N_15296,N_15024);
or U23477 (N_23477,N_18888,N_17128);
nand U23478 (N_23478,N_19490,N_16258);
xor U23479 (N_23479,N_15859,N_16243);
nor U23480 (N_23480,N_18318,N_19447);
nand U23481 (N_23481,N_17684,N_15731);
xnor U23482 (N_23482,N_19716,N_19315);
or U23483 (N_23483,N_19451,N_15550);
and U23484 (N_23484,N_18717,N_16199);
nor U23485 (N_23485,N_15986,N_19524);
xnor U23486 (N_23486,N_16060,N_17792);
xnor U23487 (N_23487,N_15297,N_16597);
or U23488 (N_23488,N_16755,N_16442);
xnor U23489 (N_23489,N_15544,N_18691);
nand U23490 (N_23490,N_17428,N_19940);
nand U23491 (N_23491,N_19147,N_18995);
xor U23492 (N_23492,N_15514,N_17784);
nand U23493 (N_23493,N_19212,N_17755);
nor U23494 (N_23494,N_16523,N_15106);
nand U23495 (N_23495,N_17323,N_18366);
nor U23496 (N_23496,N_17235,N_18666);
nand U23497 (N_23497,N_15740,N_16809);
and U23498 (N_23498,N_19247,N_17730);
or U23499 (N_23499,N_19470,N_16375);
or U23500 (N_23500,N_19682,N_16816);
xor U23501 (N_23501,N_15900,N_16321);
xnor U23502 (N_23502,N_16414,N_16697);
nand U23503 (N_23503,N_16677,N_19224);
and U23504 (N_23504,N_16568,N_17149);
nor U23505 (N_23505,N_15093,N_16423);
nor U23506 (N_23506,N_16884,N_16975);
nand U23507 (N_23507,N_17494,N_15206);
and U23508 (N_23508,N_15486,N_16534);
and U23509 (N_23509,N_15289,N_18819);
nand U23510 (N_23510,N_16859,N_16144);
and U23511 (N_23511,N_15533,N_16515);
and U23512 (N_23512,N_18587,N_15281);
and U23513 (N_23513,N_15564,N_19191);
nor U23514 (N_23514,N_19433,N_19526);
or U23515 (N_23515,N_18052,N_15050);
nand U23516 (N_23516,N_17111,N_15978);
nand U23517 (N_23517,N_16603,N_17617);
nand U23518 (N_23518,N_17666,N_17191);
or U23519 (N_23519,N_16624,N_17963);
and U23520 (N_23520,N_18738,N_17500);
nor U23521 (N_23521,N_17915,N_17406);
nor U23522 (N_23522,N_16483,N_18271);
nand U23523 (N_23523,N_18827,N_19434);
and U23524 (N_23524,N_17831,N_19208);
and U23525 (N_23525,N_15496,N_16532);
xor U23526 (N_23526,N_15167,N_15121);
xor U23527 (N_23527,N_16796,N_15243);
nand U23528 (N_23528,N_17699,N_18684);
or U23529 (N_23529,N_18381,N_19382);
nor U23530 (N_23530,N_18262,N_18798);
and U23531 (N_23531,N_17437,N_18426);
nand U23532 (N_23532,N_19055,N_19567);
xnor U23533 (N_23533,N_19802,N_16913);
nor U23534 (N_23534,N_16632,N_17567);
and U23535 (N_23535,N_16494,N_17075);
nor U23536 (N_23536,N_19113,N_15868);
xnor U23537 (N_23537,N_16032,N_16366);
nor U23538 (N_23538,N_18417,N_15613);
and U23539 (N_23539,N_18244,N_15148);
and U23540 (N_23540,N_19604,N_19159);
or U23541 (N_23541,N_19137,N_16850);
or U23542 (N_23542,N_18954,N_18425);
or U23543 (N_23543,N_18353,N_19781);
nand U23544 (N_23544,N_16859,N_16098);
nand U23545 (N_23545,N_19264,N_18931);
nor U23546 (N_23546,N_15358,N_16571);
and U23547 (N_23547,N_15355,N_18844);
or U23548 (N_23548,N_16181,N_17563);
xnor U23549 (N_23549,N_15743,N_19493);
or U23550 (N_23550,N_19135,N_19356);
and U23551 (N_23551,N_18907,N_15322);
or U23552 (N_23552,N_19970,N_15816);
and U23553 (N_23553,N_18108,N_19762);
or U23554 (N_23554,N_17249,N_15523);
xor U23555 (N_23555,N_15988,N_16438);
and U23556 (N_23556,N_16422,N_16656);
nand U23557 (N_23557,N_18281,N_17865);
xor U23558 (N_23558,N_18424,N_17988);
or U23559 (N_23559,N_15053,N_17560);
or U23560 (N_23560,N_18824,N_17493);
xor U23561 (N_23561,N_15728,N_19586);
xnor U23562 (N_23562,N_18188,N_19152);
nor U23563 (N_23563,N_19343,N_15133);
and U23564 (N_23564,N_18624,N_18961);
nand U23565 (N_23565,N_17385,N_16762);
nand U23566 (N_23566,N_15500,N_18943);
xor U23567 (N_23567,N_16528,N_15526);
nor U23568 (N_23568,N_16840,N_18776);
and U23569 (N_23569,N_19363,N_17382);
nand U23570 (N_23570,N_15482,N_18331);
nand U23571 (N_23571,N_18571,N_18729);
nor U23572 (N_23572,N_19013,N_18774);
or U23573 (N_23573,N_15513,N_17108);
xor U23574 (N_23574,N_19455,N_18231);
nor U23575 (N_23575,N_17666,N_15111);
nor U23576 (N_23576,N_16719,N_19125);
or U23577 (N_23577,N_17742,N_16796);
xor U23578 (N_23578,N_15865,N_17137);
nand U23579 (N_23579,N_18066,N_19824);
nand U23580 (N_23580,N_15953,N_17999);
nand U23581 (N_23581,N_15966,N_15561);
nand U23582 (N_23582,N_17609,N_16313);
xnor U23583 (N_23583,N_18118,N_18975);
or U23584 (N_23584,N_16046,N_18777);
or U23585 (N_23585,N_16336,N_16702);
nor U23586 (N_23586,N_15124,N_16080);
xnor U23587 (N_23587,N_16263,N_17120);
nor U23588 (N_23588,N_19899,N_17913);
xnor U23589 (N_23589,N_16085,N_15749);
xor U23590 (N_23590,N_19733,N_16872);
nand U23591 (N_23591,N_19740,N_15226);
and U23592 (N_23592,N_18146,N_16225);
nor U23593 (N_23593,N_16977,N_17751);
or U23594 (N_23594,N_15060,N_19578);
or U23595 (N_23595,N_17865,N_17548);
or U23596 (N_23596,N_16860,N_17353);
nand U23597 (N_23597,N_17701,N_19982);
xor U23598 (N_23598,N_17204,N_15803);
and U23599 (N_23599,N_17341,N_17778);
nand U23600 (N_23600,N_18664,N_19970);
or U23601 (N_23601,N_19340,N_16485);
xor U23602 (N_23602,N_18080,N_15760);
and U23603 (N_23603,N_15136,N_18747);
or U23604 (N_23604,N_19526,N_17884);
xor U23605 (N_23605,N_17997,N_19990);
nand U23606 (N_23606,N_17985,N_16586);
and U23607 (N_23607,N_18096,N_19823);
xor U23608 (N_23608,N_19680,N_17955);
nor U23609 (N_23609,N_16894,N_19220);
and U23610 (N_23610,N_16062,N_16657);
xnor U23611 (N_23611,N_19005,N_15464);
or U23612 (N_23612,N_16570,N_16523);
and U23613 (N_23613,N_18631,N_19306);
and U23614 (N_23614,N_18137,N_18632);
or U23615 (N_23615,N_19850,N_17512);
nand U23616 (N_23616,N_19593,N_16345);
and U23617 (N_23617,N_18590,N_19284);
or U23618 (N_23618,N_18633,N_19268);
and U23619 (N_23619,N_17927,N_16488);
xnor U23620 (N_23620,N_16792,N_19163);
and U23621 (N_23621,N_18490,N_16148);
and U23622 (N_23622,N_16092,N_17504);
and U23623 (N_23623,N_15667,N_17184);
nand U23624 (N_23624,N_16240,N_16183);
or U23625 (N_23625,N_15764,N_19454);
and U23626 (N_23626,N_18486,N_19830);
xnor U23627 (N_23627,N_16508,N_17120);
and U23628 (N_23628,N_16789,N_16078);
and U23629 (N_23629,N_16774,N_16513);
and U23630 (N_23630,N_16085,N_16685);
or U23631 (N_23631,N_15150,N_16566);
nor U23632 (N_23632,N_19749,N_19336);
nor U23633 (N_23633,N_15939,N_15651);
nand U23634 (N_23634,N_16178,N_19671);
and U23635 (N_23635,N_15224,N_18831);
nand U23636 (N_23636,N_16414,N_17214);
and U23637 (N_23637,N_17910,N_17043);
or U23638 (N_23638,N_19078,N_18945);
nand U23639 (N_23639,N_19022,N_19452);
nor U23640 (N_23640,N_16921,N_17627);
nor U23641 (N_23641,N_17055,N_15085);
or U23642 (N_23642,N_19883,N_16825);
nor U23643 (N_23643,N_16908,N_17986);
and U23644 (N_23644,N_19073,N_18828);
nand U23645 (N_23645,N_16153,N_17962);
nor U23646 (N_23646,N_15291,N_17038);
nor U23647 (N_23647,N_19581,N_15210);
xor U23648 (N_23648,N_17893,N_17208);
nand U23649 (N_23649,N_15092,N_19886);
or U23650 (N_23650,N_16490,N_16791);
nand U23651 (N_23651,N_16173,N_18273);
xnor U23652 (N_23652,N_19542,N_18811);
or U23653 (N_23653,N_18224,N_16652);
nor U23654 (N_23654,N_15455,N_15650);
xor U23655 (N_23655,N_19159,N_17879);
or U23656 (N_23656,N_17996,N_17708);
xnor U23657 (N_23657,N_16036,N_16864);
or U23658 (N_23658,N_17693,N_15306);
or U23659 (N_23659,N_17918,N_17127);
and U23660 (N_23660,N_15058,N_19317);
nand U23661 (N_23661,N_16608,N_17716);
xnor U23662 (N_23662,N_16453,N_15657);
nor U23663 (N_23663,N_15525,N_18171);
or U23664 (N_23664,N_15294,N_19637);
nor U23665 (N_23665,N_18614,N_19405);
nor U23666 (N_23666,N_19042,N_18274);
nand U23667 (N_23667,N_15720,N_15386);
nand U23668 (N_23668,N_19554,N_19876);
xor U23669 (N_23669,N_15776,N_17522);
or U23670 (N_23670,N_19730,N_15643);
nor U23671 (N_23671,N_17984,N_16540);
and U23672 (N_23672,N_16169,N_15736);
and U23673 (N_23673,N_16006,N_16687);
xnor U23674 (N_23674,N_19598,N_15059);
nand U23675 (N_23675,N_19625,N_16950);
nor U23676 (N_23676,N_16030,N_18212);
and U23677 (N_23677,N_16843,N_17666);
nand U23678 (N_23678,N_15171,N_17728);
or U23679 (N_23679,N_19757,N_16528);
and U23680 (N_23680,N_16955,N_19263);
xor U23681 (N_23681,N_18723,N_16442);
xnor U23682 (N_23682,N_18428,N_18616);
and U23683 (N_23683,N_18501,N_15778);
and U23684 (N_23684,N_17678,N_16537);
or U23685 (N_23685,N_15599,N_15134);
xnor U23686 (N_23686,N_17667,N_19337);
xnor U23687 (N_23687,N_19735,N_17095);
and U23688 (N_23688,N_16509,N_15004);
xnor U23689 (N_23689,N_16751,N_19430);
and U23690 (N_23690,N_17875,N_15231);
and U23691 (N_23691,N_18811,N_18968);
and U23692 (N_23692,N_17855,N_19380);
nand U23693 (N_23693,N_17359,N_15805);
or U23694 (N_23694,N_18407,N_19690);
xnor U23695 (N_23695,N_16313,N_15382);
xor U23696 (N_23696,N_15559,N_15314);
and U23697 (N_23697,N_19456,N_16922);
xor U23698 (N_23698,N_19320,N_19248);
or U23699 (N_23699,N_18249,N_18733);
nand U23700 (N_23700,N_15690,N_16046);
nand U23701 (N_23701,N_19012,N_16748);
and U23702 (N_23702,N_16469,N_16360);
and U23703 (N_23703,N_19883,N_15257);
and U23704 (N_23704,N_15561,N_15377);
and U23705 (N_23705,N_15418,N_18651);
nand U23706 (N_23706,N_17773,N_19319);
nand U23707 (N_23707,N_19891,N_16475);
nand U23708 (N_23708,N_15996,N_17979);
xnor U23709 (N_23709,N_18560,N_16113);
or U23710 (N_23710,N_19906,N_15296);
nor U23711 (N_23711,N_15239,N_18254);
or U23712 (N_23712,N_19705,N_15020);
nor U23713 (N_23713,N_19620,N_15151);
nand U23714 (N_23714,N_16590,N_19354);
nand U23715 (N_23715,N_19464,N_17463);
and U23716 (N_23716,N_19137,N_16798);
nor U23717 (N_23717,N_16973,N_18213);
or U23718 (N_23718,N_15784,N_15483);
nor U23719 (N_23719,N_19734,N_16907);
nand U23720 (N_23720,N_16212,N_15659);
nor U23721 (N_23721,N_15394,N_17985);
and U23722 (N_23722,N_19212,N_18526);
xnor U23723 (N_23723,N_17381,N_16905);
and U23724 (N_23724,N_18356,N_19430);
or U23725 (N_23725,N_19024,N_16146);
nand U23726 (N_23726,N_17836,N_19058);
and U23727 (N_23727,N_17629,N_16151);
or U23728 (N_23728,N_17473,N_15605);
xor U23729 (N_23729,N_18826,N_15451);
xor U23730 (N_23730,N_16759,N_18824);
nand U23731 (N_23731,N_17932,N_15417);
nand U23732 (N_23732,N_15070,N_15655);
xnor U23733 (N_23733,N_19872,N_19178);
nand U23734 (N_23734,N_16705,N_16608);
or U23735 (N_23735,N_17961,N_16126);
nand U23736 (N_23736,N_19039,N_16959);
or U23737 (N_23737,N_16327,N_15914);
and U23738 (N_23738,N_16660,N_18095);
nor U23739 (N_23739,N_15761,N_19934);
and U23740 (N_23740,N_19453,N_16312);
and U23741 (N_23741,N_18656,N_16605);
or U23742 (N_23742,N_17673,N_16096);
xnor U23743 (N_23743,N_18359,N_19618);
xor U23744 (N_23744,N_15082,N_18892);
nand U23745 (N_23745,N_19666,N_17777);
or U23746 (N_23746,N_17919,N_15665);
nand U23747 (N_23747,N_17951,N_19716);
and U23748 (N_23748,N_16070,N_18890);
nor U23749 (N_23749,N_15911,N_19846);
xnor U23750 (N_23750,N_19562,N_15529);
nor U23751 (N_23751,N_18274,N_19257);
or U23752 (N_23752,N_19825,N_15588);
nor U23753 (N_23753,N_16174,N_18161);
nand U23754 (N_23754,N_18510,N_17194);
and U23755 (N_23755,N_17750,N_15329);
xnor U23756 (N_23756,N_17591,N_17427);
nand U23757 (N_23757,N_19855,N_17451);
nor U23758 (N_23758,N_19611,N_15164);
and U23759 (N_23759,N_16106,N_16767);
and U23760 (N_23760,N_19053,N_15450);
nand U23761 (N_23761,N_17451,N_15761);
nand U23762 (N_23762,N_19539,N_18177);
nand U23763 (N_23763,N_15902,N_16519);
nor U23764 (N_23764,N_16849,N_15035);
xnor U23765 (N_23765,N_16753,N_17879);
nand U23766 (N_23766,N_15930,N_16957);
xnor U23767 (N_23767,N_15289,N_16938);
or U23768 (N_23768,N_16305,N_19286);
xnor U23769 (N_23769,N_17307,N_19694);
and U23770 (N_23770,N_17200,N_18640);
xor U23771 (N_23771,N_18418,N_18017);
or U23772 (N_23772,N_19880,N_16825);
nand U23773 (N_23773,N_15607,N_18763);
or U23774 (N_23774,N_17646,N_15879);
nor U23775 (N_23775,N_19103,N_19689);
xnor U23776 (N_23776,N_17511,N_19605);
nand U23777 (N_23777,N_17501,N_19053);
nor U23778 (N_23778,N_19725,N_18324);
xor U23779 (N_23779,N_18493,N_17945);
xor U23780 (N_23780,N_15698,N_16811);
nand U23781 (N_23781,N_17208,N_17143);
nand U23782 (N_23782,N_16030,N_15912);
or U23783 (N_23783,N_16817,N_17226);
and U23784 (N_23784,N_15862,N_18766);
nand U23785 (N_23785,N_18239,N_15119);
or U23786 (N_23786,N_16709,N_19782);
nand U23787 (N_23787,N_15929,N_16882);
nor U23788 (N_23788,N_19535,N_16750);
nor U23789 (N_23789,N_15270,N_18586);
nand U23790 (N_23790,N_19849,N_15131);
and U23791 (N_23791,N_19690,N_19037);
xnor U23792 (N_23792,N_18995,N_15126);
or U23793 (N_23793,N_18137,N_17796);
xnor U23794 (N_23794,N_16085,N_15186);
and U23795 (N_23795,N_18009,N_19892);
or U23796 (N_23796,N_18862,N_18909);
or U23797 (N_23797,N_17414,N_19953);
or U23798 (N_23798,N_19867,N_19317);
and U23799 (N_23799,N_15357,N_15797);
xor U23800 (N_23800,N_15066,N_19612);
nand U23801 (N_23801,N_15434,N_19747);
and U23802 (N_23802,N_19982,N_15024);
and U23803 (N_23803,N_18318,N_17299);
xnor U23804 (N_23804,N_17239,N_16889);
nor U23805 (N_23805,N_18888,N_18581);
and U23806 (N_23806,N_16503,N_15676);
nor U23807 (N_23807,N_16915,N_18315);
or U23808 (N_23808,N_18473,N_17414);
xor U23809 (N_23809,N_18800,N_17122);
nor U23810 (N_23810,N_18573,N_15848);
nand U23811 (N_23811,N_18566,N_15087);
or U23812 (N_23812,N_17363,N_19567);
xor U23813 (N_23813,N_17823,N_15488);
nor U23814 (N_23814,N_15943,N_19574);
xor U23815 (N_23815,N_18516,N_17298);
xnor U23816 (N_23816,N_19309,N_17257);
nor U23817 (N_23817,N_15541,N_16490);
xor U23818 (N_23818,N_18679,N_19885);
or U23819 (N_23819,N_17448,N_15188);
or U23820 (N_23820,N_18281,N_16357);
and U23821 (N_23821,N_16983,N_16316);
and U23822 (N_23822,N_17505,N_19857);
xnor U23823 (N_23823,N_15461,N_16712);
or U23824 (N_23824,N_15419,N_15904);
or U23825 (N_23825,N_17459,N_15197);
nand U23826 (N_23826,N_19323,N_16843);
or U23827 (N_23827,N_17655,N_17711);
nand U23828 (N_23828,N_15545,N_19420);
nor U23829 (N_23829,N_15171,N_17018);
nor U23830 (N_23830,N_15695,N_15354);
and U23831 (N_23831,N_15420,N_17840);
nand U23832 (N_23832,N_18960,N_18550);
xnor U23833 (N_23833,N_15756,N_16599);
xnor U23834 (N_23834,N_19612,N_18057);
or U23835 (N_23835,N_18488,N_18402);
and U23836 (N_23836,N_17306,N_16414);
and U23837 (N_23837,N_16002,N_19204);
and U23838 (N_23838,N_18352,N_19537);
nand U23839 (N_23839,N_16537,N_19930);
or U23840 (N_23840,N_16512,N_18830);
nor U23841 (N_23841,N_15604,N_18710);
nand U23842 (N_23842,N_17610,N_18753);
nand U23843 (N_23843,N_16729,N_16936);
nor U23844 (N_23844,N_17242,N_16487);
nor U23845 (N_23845,N_19707,N_17841);
nor U23846 (N_23846,N_18538,N_15700);
xnor U23847 (N_23847,N_17435,N_16436);
and U23848 (N_23848,N_15437,N_16664);
xnor U23849 (N_23849,N_19814,N_16691);
nand U23850 (N_23850,N_16636,N_18528);
or U23851 (N_23851,N_19151,N_18611);
or U23852 (N_23852,N_17627,N_19085);
nor U23853 (N_23853,N_15932,N_18292);
nand U23854 (N_23854,N_16417,N_15018);
or U23855 (N_23855,N_17066,N_18827);
or U23856 (N_23856,N_15213,N_17770);
or U23857 (N_23857,N_19438,N_17674);
or U23858 (N_23858,N_19154,N_19956);
and U23859 (N_23859,N_18858,N_16168);
and U23860 (N_23860,N_15949,N_17663);
nor U23861 (N_23861,N_15268,N_15201);
nand U23862 (N_23862,N_15220,N_18778);
nand U23863 (N_23863,N_15630,N_16419);
xnor U23864 (N_23864,N_17030,N_18420);
nand U23865 (N_23865,N_19873,N_16462);
nand U23866 (N_23866,N_19383,N_17015);
and U23867 (N_23867,N_15498,N_15416);
nor U23868 (N_23868,N_15930,N_16814);
nor U23869 (N_23869,N_17777,N_18198);
or U23870 (N_23870,N_15330,N_17579);
xnor U23871 (N_23871,N_16625,N_16196);
xnor U23872 (N_23872,N_16634,N_16874);
or U23873 (N_23873,N_18947,N_18167);
nor U23874 (N_23874,N_15225,N_17296);
nand U23875 (N_23875,N_18528,N_17194);
and U23876 (N_23876,N_15203,N_18640);
or U23877 (N_23877,N_16571,N_18364);
nor U23878 (N_23878,N_17092,N_17683);
nand U23879 (N_23879,N_17837,N_15632);
xnor U23880 (N_23880,N_17955,N_16074);
xor U23881 (N_23881,N_18356,N_18607);
nand U23882 (N_23882,N_17018,N_15516);
nor U23883 (N_23883,N_15535,N_19773);
and U23884 (N_23884,N_18495,N_19010);
or U23885 (N_23885,N_17882,N_18316);
nand U23886 (N_23886,N_16993,N_18239);
xnor U23887 (N_23887,N_18637,N_16913);
nor U23888 (N_23888,N_16285,N_16688);
nand U23889 (N_23889,N_17388,N_19124);
xor U23890 (N_23890,N_18134,N_19237);
nand U23891 (N_23891,N_18656,N_18062);
xnor U23892 (N_23892,N_18365,N_19063);
or U23893 (N_23893,N_17906,N_19547);
nand U23894 (N_23894,N_15604,N_15419);
or U23895 (N_23895,N_18772,N_17070);
xor U23896 (N_23896,N_16348,N_15244);
nor U23897 (N_23897,N_17078,N_19420);
and U23898 (N_23898,N_19259,N_18087);
xor U23899 (N_23899,N_19543,N_16233);
or U23900 (N_23900,N_16882,N_17681);
xnor U23901 (N_23901,N_17897,N_15094);
xor U23902 (N_23902,N_19308,N_15983);
and U23903 (N_23903,N_16157,N_17721);
nand U23904 (N_23904,N_17975,N_16409);
xor U23905 (N_23905,N_16021,N_18188);
and U23906 (N_23906,N_16919,N_15556);
nand U23907 (N_23907,N_15979,N_17164);
nor U23908 (N_23908,N_16253,N_17861);
nand U23909 (N_23909,N_18360,N_17683);
or U23910 (N_23910,N_19613,N_19924);
nor U23911 (N_23911,N_17436,N_16639);
nor U23912 (N_23912,N_19717,N_16985);
nor U23913 (N_23913,N_18887,N_16127);
xnor U23914 (N_23914,N_18366,N_18162);
nor U23915 (N_23915,N_18795,N_17638);
nand U23916 (N_23916,N_15225,N_16908);
and U23917 (N_23917,N_16961,N_17384);
or U23918 (N_23918,N_17748,N_19449);
xor U23919 (N_23919,N_18346,N_19120);
xnor U23920 (N_23920,N_18520,N_17561);
or U23921 (N_23921,N_19536,N_18414);
or U23922 (N_23922,N_18927,N_15389);
and U23923 (N_23923,N_18096,N_17655);
and U23924 (N_23924,N_19776,N_19179);
or U23925 (N_23925,N_17060,N_17502);
or U23926 (N_23926,N_18730,N_19473);
and U23927 (N_23927,N_19998,N_15970);
nand U23928 (N_23928,N_18828,N_19574);
nand U23929 (N_23929,N_15150,N_17835);
nor U23930 (N_23930,N_17004,N_17590);
and U23931 (N_23931,N_19174,N_18568);
and U23932 (N_23932,N_18350,N_16177);
nor U23933 (N_23933,N_17845,N_18828);
xor U23934 (N_23934,N_15224,N_17707);
nand U23935 (N_23935,N_19425,N_18628);
nand U23936 (N_23936,N_17075,N_17506);
nand U23937 (N_23937,N_16811,N_19962);
or U23938 (N_23938,N_18792,N_17588);
xnor U23939 (N_23939,N_17854,N_19389);
nor U23940 (N_23940,N_15577,N_15929);
and U23941 (N_23941,N_17081,N_18853);
nand U23942 (N_23942,N_15866,N_19843);
and U23943 (N_23943,N_19123,N_15546);
nand U23944 (N_23944,N_15931,N_19218);
and U23945 (N_23945,N_17587,N_15881);
or U23946 (N_23946,N_15284,N_16254);
xor U23947 (N_23947,N_16066,N_19028);
nand U23948 (N_23948,N_16944,N_18537);
nor U23949 (N_23949,N_17826,N_19915);
nor U23950 (N_23950,N_15473,N_16276);
xnor U23951 (N_23951,N_15793,N_16493);
nand U23952 (N_23952,N_15138,N_18686);
or U23953 (N_23953,N_15668,N_18296);
and U23954 (N_23954,N_18792,N_15588);
nor U23955 (N_23955,N_19429,N_17072);
or U23956 (N_23956,N_17514,N_17482);
and U23957 (N_23957,N_16599,N_15503);
and U23958 (N_23958,N_15900,N_16182);
nor U23959 (N_23959,N_16085,N_15585);
and U23960 (N_23960,N_19370,N_17880);
xor U23961 (N_23961,N_15509,N_19722);
nor U23962 (N_23962,N_19396,N_16854);
or U23963 (N_23963,N_18858,N_15099);
or U23964 (N_23964,N_16391,N_18790);
or U23965 (N_23965,N_17638,N_16720);
nand U23966 (N_23966,N_18363,N_16531);
xor U23967 (N_23967,N_18314,N_16814);
nand U23968 (N_23968,N_16700,N_15275);
and U23969 (N_23969,N_16976,N_19239);
or U23970 (N_23970,N_16676,N_18642);
nor U23971 (N_23971,N_17920,N_15058);
xor U23972 (N_23972,N_18010,N_17610);
xor U23973 (N_23973,N_15583,N_19745);
nand U23974 (N_23974,N_17213,N_16164);
and U23975 (N_23975,N_19707,N_15920);
nor U23976 (N_23976,N_18924,N_16529);
nand U23977 (N_23977,N_16967,N_16211);
or U23978 (N_23978,N_19007,N_18053);
xor U23979 (N_23979,N_15614,N_19749);
and U23980 (N_23980,N_18694,N_18159);
or U23981 (N_23981,N_19559,N_17060);
or U23982 (N_23982,N_18639,N_19181);
or U23983 (N_23983,N_17823,N_18221);
xnor U23984 (N_23984,N_16889,N_18462);
xor U23985 (N_23985,N_17559,N_15523);
or U23986 (N_23986,N_19693,N_16835);
and U23987 (N_23987,N_15314,N_15567);
and U23988 (N_23988,N_15708,N_16058);
and U23989 (N_23989,N_18373,N_18399);
and U23990 (N_23990,N_18398,N_19439);
or U23991 (N_23991,N_18648,N_18949);
or U23992 (N_23992,N_18468,N_18568);
or U23993 (N_23993,N_15050,N_19810);
xor U23994 (N_23994,N_15568,N_16206);
or U23995 (N_23995,N_19567,N_15987);
and U23996 (N_23996,N_17158,N_15664);
nand U23997 (N_23997,N_18548,N_15628);
and U23998 (N_23998,N_19544,N_15287);
nor U23999 (N_23999,N_16120,N_18260);
or U24000 (N_24000,N_18717,N_18869);
nand U24001 (N_24001,N_15134,N_15495);
or U24002 (N_24002,N_17608,N_15496);
nand U24003 (N_24003,N_18537,N_17402);
nor U24004 (N_24004,N_19112,N_18881);
nor U24005 (N_24005,N_16929,N_18810);
or U24006 (N_24006,N_19294,N_15552);
or U24007 (N_24007,N_18324,N_17179);
or U24008 (N_24008,N_18066,N_19797);
and U24009 (N_24009,N_15637,N_16003);
nor U24010 (N_24010,N_18236,N_16389);
nor U24011 (N_24011,N_17797,N_18874);
or U24012 (N_24012,N_16483,N_15344);
nand U24013 (N_24013,N_15316,N_17040);
nand U24014 (N_24014,N_17233,N_18742);
or U24015 (N_24015,N_17151,N_16234);
nand U24016 (N_24016,N_18633,N_18169);
nor U24017 (N_24017,N_19317,N_15704);
xor U24018 (N_24018,N_17388,N_16240);
nor U24019 (N_24019,N_16940,N_19779);
xnor U24020 (N_24020,N_15793,N_15741);
nor U24021 (N_24021,N_17350,N_18055);
or U24022 (N_24022,N_16675,N_19689);
xnor U24023 (N_24023,N_18535,N_18456);
nand U24024 (N_24024,N_19516,N_17932);
and U24025 (N_24025,N_19043,N_17345);
xnor U24026 (N_24026,N_19872,N_18802);
nor U24027 (N_24027,N_17323,N_18159);
nor U24028 (N_24028,N_17082,N_19955);
nand U24029 (N_24029,N_16966,N_15696);
nand U24030 (N_24030,N_19243,N_15903);
xor U24031 (N_24031,N_19607,N_18282);
xnor U24032 (N_24032,N_15529,N_19506);
or U24033 (N_24033,N_18552,N_19663);
and U24034 (N_24034,N_15516,N_16677);
and U24035 (N_24035,N_17705,N_16029);
and U24036 (N_24036,N_16399,N_15155);
nand U24037 (N_24037,N_15752,N_16793);
nor U24038 (N_24038,N_17801,N_17509);
or U24039 (N_24039,N_19064,N_17527);
xnor U24040 (N_24040,N_17910,N_16194);
nand U24041 (N_24041,N_17510,N_19424);
nand U24042 (N_24042,N_19327,N_17657);
xnor U24043 (N_24043,N_15722,N_19182);
nor U24044 (N_24044,N_19893,N_16537);
nor U24045 (N_24045,N_16581,N_15508);
and U24046 (N_24046,N_17558,N_19977);
nand U24047 (N_24047,N_19843,N_17908);
xor U24048 (N_24048,N_19391,N_18571);
xor U24049 (N_24049,N_16580,N_16865);
xnor U24050 (N_24050,N_15252,N_18508);
and U24051 (N_24051,N_15212,N_16750);
or U24052 (N_24052,N_19717,N_18901);
nor U24053 (N_24053,N_16124,N_15073);
and U24054 (N_24054,N_15987,N_16070);
nor U24055 (N_24055,N_16177,N_19228);
nand U24056 (N_24056,N_17424,N_16914);
xor U24057 (N_24057,N_15713,N_18981);
and U24058 (N_24058,N_16905,N_16659);
xnor U24059 (N_24059,N_18415,N_19465);
or U24060 (N_24060,N_15729,N_17141);
nand U24061 (N_24061,N_18472,N_19260);
or U24062 (N_24062,N_19401,N_18152);
and U24063 (N_24063,N_18260,N_19558);
nor U24064 (N_24064,N_16913,N_19119);
nor U24065 (N_24065,N_18178,N_18959);
or U24066 (N_24066,N_19448,N_18421);
nor U24067 (N_24067,N_17776,N_15114);
nor U24068 (N_24068,N_16644,N_17483);
nor U24069 (N_24069,N_15111,N_18619);
nor U24070 (N_24070,N_16610,N_18593);
and U24071 (N_24071,N_17528,N_17797);
nor U24072 (N_24072,N_15111,N_16693);
or U24073 (N_24073,N_17529,N_16030);
nor U24074 (N_24074,N_15618,N_18415);
nor U24075 (N_24075,N_15091,N_19384);
xor U24076 (N_24076,N_19267,N_18682);
or U24077 (N_24077,N_18748,N_16411);
nor U24078 (N_24078,N_19129,N_15737);
nor U24079 (N_24079,N_19633,N_16561);
xor U24080 (N_24080,N_17762,N_19174);
xnor U24081 (N_24081,N_18720,N_16214);
and U24082 (N_24082,N_17147,N_17574);
and U24083 (N_24083,N_17522,N_19096);
xor U24084 (N_24084,N_16340,N_16277);
xor U24085 (N_24085,N_16475,N_17788);
and U24086 (N_24086,N_18200,N_17433);
xor U24087 (N_24087,N_19659,N_17368);
xor U24088 (N_24088,N_17959,N_18870);
xnor U24089 (N_24089,N_15595,N_17703);
nor U24090 (N_24090,N_18609,N_16684);
nor U24091 (N_24091,N_17413,N_19650);
or U24092 (N_24092,N_15285,N_17771);
or U24093 (N_24093,N_18050,N_17310);
or U24094 (N_24094,N_17203,N_18480);
nand U24095 (N_24095,N_15724,N_18413);
nor U24096 (N_24096,N_15363,N_16989);
or U24097 (N_24097,N_16277,N_15547);
and U24098 (N_24098,N_16226,N_15397);
nand U24099 (N_24099,N_18693,N_15768);
xnor U24100 (N_24100,N_17813,N_17552);
nand U24101 (N_24101,N_19255,N_15729);
xor U24102 (N_24102,N_15169,N_18798);
nand U24103 (N_24103,N_19651,N_16322);
xor U24104 (N_24104,N_19205,N_16585);
or U24105 (N_24105,N_16224,N_19872);
xor U24106 (N_24106,N_19922,N_17269);
nand U24107 (N_24107,N_17158,N_17471);
nor U24108 (N_24108,N_16066,N_17333);
nand U24109 (N_24109,N_16461,N_19099);
and U24110 (N_24110,N_15376,N_16650);
xnor U24111 (N_24111,N_17576,N_16369);
and U24112 (N_24112,N_15806,N_18465);
or U24113 (N_24113,N_19719,N_16560);
or U24114 (N_24114,N_19210,N_18796);
nor U24115 (N_24115,N_15860,N_15934);
or U24116 (N_24116,N_15642,N_16135);
or U24117 (N_24117,N_17236,N_17294);
nand U24118 (N_24118,N_19165,N_19474);
or U24119 (N_24119,N_17763,N_19493);
nor U24120 (N_24120,N_17306,N_15190);
or U24121 (N_24121,N_15090,N_16573);
xnor U24122 (N_24122,N_15698,N_15308);
nor U24123 (N_24123,N_16382,N_17016);
and U24124 (N_24124,N_16305,N_19360);
nand U24125 (N_24125,N_15256,N_15050);
nor U24126 (N_24126,N_16003,N_17758);
or U24127 (N_24127,N_15724,N_17754);
nand U24128 (N_24128,N_17978,N_18215);
or U24129 (N_24129,N_16384,N_16077);
xor U24130 (N_24130,N_18367,N_17110);
or U24131 (N_24131,N_18304,N_19477);
or U24132 (N_24132,N_17420,N_19935);
and U24133 (N_24133,N_18381,N_19138);
nor U24134 (N_24134,N_18348,N_19734);
xor U24135 (N_24135,N_16899,N_15989);
xor U24136 (N_24136,N_17600,N_19280);
nor U24137 (N_24137,N_19703,N_17209);
or U24138 (N_24138,N_19450,N_15656);
and U24139 (N_24139,N_15637,N_17575);
nor U24140 (N_24140,N_19509,N_16278);
xnor U24141 (N_24141,N_16807,N_16216);
nand U24142 (N_24142,N_16225,N_18248);
nor U24143 (N_24143,N_16105,N_16784);
xor U24144 (N_24144,N_18816,N_19596);
nand U24145 (N_24145,N_16101,N_15404);
or U24146 (N_24146,N_16946,N_16948);
xor U24147 (N_24147,N_19973,N_16658);
nor U24148 (N_24148,N_15054,N_15261);
xor U24149 (N_24149,N_19471,N_18185);
xor U24150 (N_24150,N_18950,N_15987);
xor U24151 (N_24151,N_18059,N_17789);
or U24152 (N_24152,N_15479,N_18305);
and U24153 (N_24153,N_17918,N_17527);
nor U24154 (N_24154,N_17036,N_18481);
xnor U24155 (N_24155,N_17761,N_16174);
xnor U24156 (N_24156,N_15523,N_17485);
nand U24157 (N_24157,N_17092,N_15297);
xor U24158 (N_24158,N_15353,N_18450);
or U24159 (N_24159,N_18616,N_15698);
and U24160 (N_24160,N_15614,N_15223);
and U24161 (N_24161,N_16253,N_15637);
and U24162 (N_24162,N_19679,N_17687);
and U24163 (N_24163,N_17697,N_18076);
nand U24164 (N_24164,N_19568,N_18332);
or U24165 (N_24165,N_16606,N_19160);
nand U24166 (N_24166,N_16179,N_19624);
nand U24167 (N_24167,N_16463,N_16231);
nand U24168 (N_24168,N_19944,N_18724);
and U24169 (N_24169,N_16078,N_16228);
xnor U24170 (N_24170,N_17868,N_15141);
xnor U24171 (N_24171,N_19510,N_17354);
xor U24172 (N_24172,N_16551,N_16071);
and U24173 (N_24173,N_16975,N_15308);
nand U24174 (N_24174,N_17507,N_18604);
xnor U24175 (N_24175,N_18468,N_19994);
or U24176 (N_24176,N_17478,N_15340);
nor U24177 (N_24177,N_17813,N_17039);
xnor U24178 (N_24178,N_18131,N_19925);
nor U24179 (N_24179,N_19212,N_18219);
nor U24180 (N_24180,N_17498,N_16310);
or U24181 (N_24181,N_15119,N_19397);
and U24182 (N_24182,N_15720,N_19336);
xor U24183 (N_24183,N_15279,N_15624);
nor U24184 (N_24184,N_19854,N_18256);
nor U24185 (N_24185,N_17788,N_16589);
and U24186 (N_24186,N_19331,N_16529);
xor U24187 (N_24187,N_15239,N_16097);
nand U24188 (N_24188,N_16614,N_19935);
nor U24189 (N_24189,N_16966,N_18708);
or U24190 (N_24190,N_15108,N_18842);
xnor U24191 (N_24191,N_19262,N_16314);
or U24192 (N_24192,N_18627,N_17704);
nor U24193 (N_24193,N_17008,N_17962);
or U24194 (N_24194,N_19317,N_17767);
nand U24195 (N_24195,N_18800,N_16399);
xor U24196 (N_24196,N_18550,N_15788);
nand U24197 (N_24197,N_18373,N_17974);
xnor U24198 (N_24198,N_19766,N_15295);
nand U24199 (N_24199,N_16732,N_16748);
nor U24200 (N_24200,N_19045,N_19897);
xor U24201 (N_24201,N_19995,N_15208);
or U24202 (N_24202,N_18359,N_17619);
nor U24203 (N_24203,N_18468,N_16196);
or U24204 (N_24204,N_16305,N_19730);
nor U24205 (N_24205,N_16314,N_19800);
nor U24206 (N_24206,N_17328,N_18549);
or U24207 (N_24207,N_17451,N_18967);
or U24208 (N_24208,N_16405,N_18443);
or U24209 (N_24209,N_15960,N_18903);
nor U24210 (N_24210,N_19576,N_17320);
or U24211 (N_24211,N_19494,N_15836);
nor U24212 (N_24212,N_19615,N_19458);
and U24213 (N_24213,N_18751,N_15058);
nand U24214 (N_24214,N_16552,N_18604);
nand U24215 (N_24215,N_18382,N_15974);
nor U24216 (N_24216,N_19651,N_19162);
and U24217 (N_24217,N_15529,N_17178);
xor U24218 (N_24218,N_19592,N_15448);
xnor U24219 (N_24219,N_16514,N_18987);
or U24220 (N_24220,N_17568,N_18436);
or U24221 (N_24221,N_18428,N_16347);
xnor U24222 (N_24222,N_17081,N_16721);
xnor U24223 (N_24223,N_15388,N_18670);
nor U24224 (N_24224,N_16748,N_19719);
nor U24225 (N_24225,N_15260,N_17895);
xnor U24226 (N_24226,N_17005,N_17423);
nand U24227 (N_24227,N_18034,N_18473);
nor U24228 (N_24228,N_15154,N_19887);
nand U24229 (N_24229,N_17846,N_19239);
nor U24230 (N_24230,N_18995,N_18077);
and U24231 (N_24231,N_18163,N_15480);
or U24232 (N_24232,N_19631,N_17267);
nand U24233 (N_24233,N_16323,N_19639);
or U24234 (N_24234,N_19305,N_17528);
xor U24235 (N_24235,N_16906,N_18066);
nor U24236 (N_24236,N_18513,N_19061);
or U24237 (N_24237,N_16103,N_15247);
or U24238 (N_24238,N_17088,N_17074);
or U24239 (N_24239,N_17017,N_16908);
nor U24240 (N_24240,N_16315,N_15867);
nor U24241 (N_24241,N_18827,N_19118);
nand U24242 (N_24242,N_16258,N_17770);
nor U24243 (N_24243,N_18441,N_16427);
nand U24244 (N_24244,N_17577,N_17131);
nand U24245 (N_24245,N_16547,N_18947);
nand U24246 (N_24246,N_15790,N_16023);
nand U24247 (N_24247,N_15002,N_17422);
and U24248 (N_24248,N_15472,N_15386);
and U24249 (N_24249,N_18726,N_17634);
xnor U24250 (N_24250,N_17390,N_19221);
nand U24251 (N_24251,N_19540,N_15785);
xnor U24252 (N_24252,N_16422,N_15601);
xnor U24253 (N_24253,N_19834,N_19334);
and U24254 (N_24254,N_15091,N_15899);
xor U24255 (N_24255,N_17969,N_18232);
and U24256 (N_24256,N_15297,N_18932);
or U24257 (N_24257,N_16862,N_17741);
nand U24258 (N_24258,N_17881,N_18225);
xor U24259 (N_24259,N_16031,N_15390);
nand U24260 (N_24260,N_17083,N_16346);
and U24261 (N_24261,N_19915,N_16968);
nand U24262 (N_24262,N_18274,N_16905);
nand U24263 (N_24263,N_18414,N_19482);
nand U24264 (N_24264,N_15419,N_19394);
nor U24265 (N_24265,N_15035,N_15560);
nand U24266 (N_24266,N_16765,N_18415);
nor U24267 (N_24267,N_18400,N_15780);
nor U24268 (N_24268,N_15956,N_19466);
xor U24269 (N_24269,N_19346,N_17932);
xnor U24270 (N_24270,N_17406,N_17479);
nor U24271 (N_24271,N_19660,N_19430);
nand U24272 (N_24272,N_17077,N_19582);
nor U24273 (N_24273,N_18502,N_16353);
xnor U24274 (N_24274,N_16599,N_19162);
nor U24275 (N_24275,N_19318,N_17556);
xnor U24276 (N_24276,N_18632,N_17167);
nand U24277 (N_24277,N_16480,N_17280);
or U24278 (N_24278,N_15889,N_18763);
nand U24279 (N_24279,N_16972,N_19248);
and U24280 (N_24280,N_17175,N_16819);
nor U24281 (N_24281,N_17041,N_18318);
nor U24282 (N_24282,N_19263,N_18134);
nor U24283 (N_24283,N_19460,N_17058);
and U24284 (N_24284,N_17424,N_16143);
xor U24285 (N_24285,N_16762,N_19799);
and U24286 (N_24286,N_19323,N_16044);
or U24287 (N_24287,N_15873,N_19782);
nand U24288 (N_24288,N_19918,N_19812);
or U24289 (N_24289,N_15191,N_16434);
and U24290 (N_24290,N_18794,N_19515);
or U24291 (N_24291,N_19755,N_17947);
nand U24292 (N_24292,N_19569,N_18079);
nand U24293 (N_24293,N_15994,N_15575);
nor U24294 (N_24294,N_16332,N_16816);
or U24295 (N_24295,N_17342,N_15504);
xor U24296 (N_24296,N_19013,N_19130);
nor U24297 (N_24297,N_19984,N_15612);
or U24298 (N_24298,N_19966,N_17343);
and U24299 (N_24299,N_17285,N_19354);
nand U24300 (N_24300,N_16275,N_15127);
nand U24301 (N_24301,N_19698,N_18529);
and U24302 (N_24302,N_18650,N_18679);
xnor U24303 (N_24303,N_17769,N_19079);
xor U24304 (N_24304,N_19594,N_17035);
nor U24305 (N_24305,N_16521,N_17123);
nand U24306 (N_24306,N_17875,N_19950);
or U24307 (N_24307,N_16276,N_19114);
nor U24308 (N_24308,N_17001,N_19921);
xnor U24309 (N_24309,N_18411,N_15065);
nand U24310 (N_24310,N_15827,N_17659);
or U24311 (N_24311,N_17121,N_17746);
and U24312 (N_24312,N_16662,N_16440);
and U24313 (N_24313,N_19515,N_15587);
and U24314 (N_24314,N_15141,N_15676);
or U24315 (N_24315,N_18076,N_18552);
nand U24316 (N_24316,N_16197,N_16684);
or U24317 (N_24317,N_15788,N_17579);
nand U24318 (N_24318,N_19083,N_17026);
or U24319 (N_24319,N_15549,N_15077);
or U24320 (N_24320,N_17106,N_16192);
xor U24321 (N_24321,N_15354,N_17861);
or U24322 (N_24322,N_17192,N_17253);
xnor U24323 (N_24323,N_17747,N_18583);
and U24324 (N_24324,N_17742,N_18420);
or U24325 (N_24325,N_15166,N_19916);
nor U24326 (N_24326,N_15678,N_16883);
nand U24327 (N_24327,N_15387,N_19571);
and U24328 (N_24328,N_17130,N_19159);
or U24329 (N_24329,N_15897,N_18359);
and U24330 (N_24330,N_16456,N_19559);
nor U24331 (N_24331,N_18346,N_16158);
or U24332 (N_24332,N_15250,N_19682);
or U24333 (N_24333,N_19771,N_19124);
nand U24334 (N_24334,N_16774,N_19741);
or U24335 (N_24335,N_19388,N_18740);
or U24336 (N_24336,N_18687,N_19690);
or U24337 (N_24337,N_19200,N_18467);
nor U24338 (N_24338,N_15045,N_17946);
or U24339 (N_24339,N_19496,N_17047);
nor U24340 (N_24340,N_18233,N_17450);
and U24341 (N_24341,N_16087,N_19908);
nand U24342 (N_24342,N_16077,N_19877);
nor U24343 (N_24343,N_16688,N_19071);
nor U24344 (N_24344,N_18167,N_17479);
nor U24345 (N_24345,N_19942,N_15906);
xor U24346 (N_24346,N_19784,N_15409);
xnor U24347 (N_24347,N_15252,N_17859);
nor U24348 (N_24348,N_19322,N_17068);
or U24349 (N_24349,N_19027,N_19585);
nand U24350 (N_24350,N_19799,N_17869);
or U24351 (N_24351,N_19230,N_15133);
nor U24352 (N_24352,N_19462,N_18375);
and U24353 (N_24353,N_18863,N_18426);
nor U24354 (N_24354,N_18096,N_17738);
or U24355 (N_24355,N_15350,N_19877);
nand U24356 (N_24356,N_17148,N_16950);
nor U24357 (N_24357,N_17660,N_17601);
xnor U24358 (N_24358,N_19317,N_18655);
or U24359 (N_24359,N_15181,N_19360);
and U24360 (N_24360,N_15303,N_17005);
xor U24361 (N_24361,N_15271,N_18075);
nand U24362 (N_24362,N_19611,N_17956);
nand U24363 (N_24363,N_15401,N_17164);
nand U24364 (N_24364,N_15030,N_17046);
and U24365 (N_24365,N_19005,N_19885);
nor U24366 (N_24366,N_19462,N_15215);
nand U24367 (N_24367,N_16215,N_18854);
or U24368 (N_24368,N_16711,N_18377);
and U24369 (N_24369,N_17818,N_15988);
and U24370 (N_24370,N_19116,N_18074);
nor U24371 (N_24371,N_17521,N_18851);
or U24372 (N_24372,N_18895,N_18102);
or U24373 (N_24373,N_16063,N_18324);
or U24374 (N_24374,N_15536,N_19102);
and U24375 (N_24375,N_17958,N_19622);
or U24376 (N_24376,N_17052,N_18676);
nor U24377 (N_24377,N_15880,N_18708);
or U24378 (N_24378,N_15020,N_15390);
or U24379 (N_24379,N_19224,N_18534);
nand U24380 (N_24380,N_19963,N_18830);
nor U24381 (N_24381,N_16707,N_19341);
and U24382 (N_24382,N_16837,N_17081);
or U24383 (N_24383,N_16990,N_17334);
nand U24384 (N_24384,N_17623,N_18601);
or U24385 (N_24385,N_17362,N_18792);
nand U24386 (N_24386,N_15776,N_17322);
nand U24387 (N_24387,N_19097,N_18104);
xnor U24388 (N_24388,N_18909,N_15543);
or U24389 (N_24389,N_16047,N_16095);
nand U24390 (N_24390,N_15176,N_15735);
nand U24391 (N_24391,N_19571,N_17854);
and U24392 (N_24392,N_18977,N_18871);
and U24393 (N_24393,N_18798,N_19926);
and U24394 (N_24394,N_18677,N_15963);
nand U24395 (N_24395,N_16956,N_19125);
nor U24396 (N_24396,N_19658,N_19113);
and U24397 (N_24397,N_16900,N_19670);
xnor U24398 (N_24398,N_18760,N_18891);
and U24399 (N_24399,N_19389,N_19359);
nand U24400 (N_24400,N_19654,N_18235);
or U24401 (N_24401,N_15993,N_17634);
nand U24402 (N_24402,N_15769,N_15945);
xnor U24403 (N_24403,N_15684,N_19631);
nand U24404 (N_24404,N_16496,N_16042);
xnor U24405 (N_24405,N_17141,N_19769);
xnor U24406 (N_24406,N_18979,N_19213);
and U24407 (N_24407,N_19498,N_15208);
xnor U24408 (N_24408,N_15527,N_15963);
nor U24409 (N_24409,N_17681,N_17344);
and U24410 (N_24410,N_18338,N_18447);
or U24411 (N_24411,N_18209,N_18751);
and U24412 (N_24412,N_17904,N_17347);
and U24413 (N_24413,N_17650,N_17127);
xor U24414 (N_24414,N_19366,N_17658);
nor U24415 (N_24415,N_16004,N_18854);
nor U24416 (N_24416,N_18709,N_17123);
xor U24417 (N_24417,N_17234,N_18203);
nor U24418 (N_24418,N_15191,N_15061);
or U24419 (N_24419,N_18006,N_17402);
nor U24420 (N_24420,N_19072,N_19611);
xor U24421 (N_24421,N_19051,N_16591);
or U24422 (N_24422,N_19002,N_16152);
nand U24423 (N_24423,N_15411,N_18101);
xnor U24424 (N_24424,N_19230,N_19936);
nand U24425 (N_24425,N_16314,N_18295);
nand U24426 (N_24426,N_18227,N_17001);
and U24427 (N_24427,N_17513,N_19567);
nand U24428 (N_24428,N_15736,N_19890);
nand U24429 (N_24429,N_15904,N_16740);
nand U24430 (N_24430,N_19086,N_18372);
and U24431 (N_24431,N_18366,N_19681);
xor U24432 (N_24432,N_17675,N_15535);
nand U24433 (N_24433,N_17051,N_19336);
nor U24434 (N_24434,N_16095,N_19000);
nand U24435 (N_24435,N_18768,N_18661);
xnor U24436 (N_24436,N_15383,N_17488);
xnor U24437 (N_24437,N_17681,N_15895);
or U24438 (N_24438,N_18727,N_19119);
nand U24439 (N_24439,N_19252,N_19043);
and U24440 (N_24440,N_16448,N_19696);
and U24441 (N_24441,N_18058,N_19708);
nor U24442 (N_24442,N_19327,N_17748);
nor U24443 (N_24443,N_19656,N_15623);
or U24444 (N_24444,N_15585,N_17282);
and U24445 (N_24445,N_18274,N_15414);
and U24446 (N_24446,N_17023,N_16203);
and U24447 (N_24447,N_16100,N_19913);
nor U24448 (N_24448,N_19372,N_16777);
and U24449 (N_24449,N_17425,N_15243);
nand U24450 (N_24450,N_18534,N_19939);
or U24451 (N_24451,N_16982,N_16978);
nand U24452 (N_24452,N_17341,N_19600);
and U24453 (N_24453,N_17100,N_15064);
and U24454 (N_24454,N_18541,N_19580);
nand U24455 (N_24455,N_17214,N_19533);
nand U24456 (N_24456,N_19885,N_16253);
and U24457 (N_24457,N_16158,N_18933);
nand U24458 (N_24458,N_18645,N_16858);
and U24459 (N_24459,N_19702,N_16756);
xnor U24460 (N_24460,N_15215,N_19083);
or U24461 (N_24461,N_17567,N_15506);
xnor U24462 (N_24462,N_15970,N_17363);
and U24463 (N_24463,N_16472,N_19270);
xor U24464 (N_24464,N_18891,N_19793);
xor U24465 (N_24465,N_16581,N_17411);
nand U24466 (N_24466,N_16388,N_17096);
and U24467 (N_24467,N_17438,N_16395);
nand U24468 (N_24468,N_17220,N_15491);
xor U24469 (N_24469,N_19490,N_19372);
or U24470 (N_24470,N_19825,N_19709);
xnor U24471 (N_24471,N_18237,N_16140);
xor U24472 (N_24472,N_18406,N_16268);
or U24473 (N_24473,N_16500,N_15470);
nor U24474 (N_24474,N_19978,N_16279);
xnor U24475 (N_24475,N_15134,N_16418);
xor U24476 (N_24476,N_16289,N_19194);
nor U24477 (N_24477,N_16828,N_18656);
nor U24478 (N_24478,N_15913,N_18285);
nand U24479 (N_24479,N_17047,N_17734);
or U24480 (N_24480,N_16912,N_16789);
xnor U24481 (N_24481,N_17385,N_19753);
nand U24482 (N_24482,N_17902,N_15041);
or U24483 (N_24483,N_15890,N_18162);
nand U24484 (N_24484,N_17380,N_16439);
xnor U24485 (N_24485,N_19947,N_15264);
and U24486 (N_24486,N_19396,N_17429);
and U24487 (N_24487,N_17449,N_19255);
and U24488 (N_24488,N_17523,N_18738);
nand U24489 (N_24489,N_15753,N_19508);
nand U24490 (N_24490,N_18033,N_18292);
and U24491 (N_24491,N_17808,N_19216);
nor U24492 (N_24492,N_18197,N_15978);
nor U24493 (N_24493,N_16232,N_18945);
nand U24494 (N_24494,N_16807,N_17658);
and U24495 (N_24495,N_16821,N_16208);
nor U24496 (N_24496,N_17009,N_18722);
nor U24497 (N_24497,N_15454,N_18998);
nand U24498 (N_24498,N_16350,N_15487);
and U24499 (N_24499,N_16357,N_17654);
nand U24500 (N_24500,N_17381,N_18844);
nand U24501 (N_24501,N_18829,N_18681);
xnor U24502 (N_24502,N_18058,N_19106);
and U24503 (N_24503,N_15673,N_17377);
nor U24504 (N_24504,N_19574,N_17326);
or U24505 (N_24505,N_17382,N_16981);
nor U24506 (N_24506,N_17848,N_19238);
and U24507 (N_24507,N_15689,N_16840);
and U24508 (N_24508,N_17987,N_17716);
and U24509 (N_24509,N_16473,N_18877);
nand U24510 (N_24510,N_19105,N_17701);
nand U24511 (N_24511,N_18635,N_17784);
nand U24512 (N_24512,N_19507,N_18543);
nand U24513 (N_24513,N_16527,N_19987);
nand U24514 (N_24514,N_17421,N_15427);
nand U24515 (N_24515,N_19561,N_16419);
xor U24516 (N_24516,N_17501,N_18850);
or U24517 (N_24517,N_16691,N_15396);
xnor U24518 (N_24518,N_16387,N_16749);
xor U24519 (N_24519,N_18543,N_18388);
xor U24520 (N_24520,N_15068,N_15536);
nor U24521 (N_24521,N_17643,N_17446);
xor U24522 (N_24522,N_16392,N_19993);
and U24523 (N_24523,N_19903,N_18777);
and U24524 (N_24524,N_15817,N_18643);
nand U24525 (N_24525,N_15646,N_15968);
and U24526 (N_24526,N_19381,N_17508);
xor U24527 (N_24527,N_17177,N_16015);
xnor U24528 (N_24528,N_16719,N_19546);
nand U24529 (N_24529,N_17035,N_19669);
xor U24530 (N_24530,N_17379,N_16547);
and U24531 (N_24531,N_16599,N_19890);
nand U24532 (N_24532,N_16034,N_17517);
nand U24533 (N_24533,N_16435,N_15733);
nand U24534 (N_24534,N_15719,N_16981);
nand U24535 (N_24535,N_17244,N_15118);
or U24536 (N_24536,N_17576,N_18433);
xor U24537 (N_24537,N_17485,N_15623);
and U24538 (N_24538,N_15543,N_15894);
nor U24539 (N_24539,N_18918,N_17148);
and U24540 (N_24540,N_18224,N_18238);
and U24541 (N_24541,N_15885,N_16187);
and U24542 (N_24542,N_17941,N_18499);
xnor U24543 (N_24543,N_19242,N_16546);
nor U24544 (N_24544,N_19836,N_17045);
and U24545 (N_24545,N_16473,N_15202);
nand U24546 (N_24546,N_18408,N_18077);
and U24547 (N_24547,N_15333,N_15555);
nor U24548 (N_24548,N_19245,N_15640);
xor U24549 (N_24549,N_16544,N_17093);
xor U24550 (N_24550,N_16152,N_17893);
nand U24551 (N_24551,N_19683,N_18414);
nand U24552 (N_24552,N_16976,N_17652);
nor U24553 (N_24553,N_18733,N_17629);
and U24554 (N_24554,N_17821,N_15483);
nor U24555 (N_24555,N_18299,N_17336);
xnor U24556 (N_24556,N_18650,N_17479);
and U24557 (N_24557,N_16949,N_16093);
nand U24558 (N_24558,N_17181,N_16469);
and U24559 (N_24559,N_16813,N_18512);
nand U24560 (N_24560,N_17002,N_18418);
xnor U24561 (N_24561,N_18812,N_19399);
nand U24562 (N_24562,N_19810,N_17645);
nand U24563 (N_24563,N_17836,N_19909);
nand U24564 (N_24564,N_15738,N_15760);
or U24565 (N_24565,N_15997,N_16118);
nor U24566 (N_24566,N_18407,N_16602);
nor U24567 (N_24567,N_16950,N_19566);
nand U24568 (N_24568,N_16039,N_17472);
xnor U24569 (N_24569,N_19063,N_19824);
and U24570 (N_24570,N_18100,N_15179);
nor U24571 (N_24571,N_17501,N_19264);
xor U24572 (N_24572,N_18393,N_19517);
xnor U24573 (N_24573,N_15490,N_15868);
nor U24574 (N_24574,N_16298,N_17187);
or U24575 (N_24575,N_15669,N_19369);
nor U24576 (N_24576,N_18535,N_16315);
xnor U24577 (N_24577,N_18088,N_18568);
and U24578 (N_24578,N_18168,N_16176);
nand U24579 (N_24579,N_16841,N_15199);
and U24580 (N_24580,N_18341,N_15115);
xnor U24581 (N_24581,N_16966,N_17846);
and U24582 (N_24582,N_16992,N_18573);
nor U24583 (N_24583,N_19752,N_19221);
and U24584 (N_24584,N_17935,N_15916);
xor U24585 (N_24585,N_19848,N_18597);
and U24586 (N_24586,N_15063,N_19502);
nand U24587 (N_24587,N_17527,N_15238);
or U24588 (N_24588,N_18821,N_19151);
or U24589 (N_24589,N_17708,N_19966);
xnor U24590 (N_24590,N_19731,N_19363);
and U24591 (N_24591,N_15519,N_16974);
xor U24592 (N_24592,N_17823,N_19451);
xnor U24593 (N_24593,N_17337,N_15619);
nand U24594 (N_24594,N_18202,N_17974);
nand U24595 (N_24595,N_17061,N_16426);
and U24596 (N_24596,N_19314,N_15005);
nor U24597 (N_24597,N_17890,N_17307);
or U24598 (N_24598,N_19942,N_15449);
nand U24599 (N_24599,N_19039,N_19787);
or U24600 (N_24600,N_18451,N_19019);
or U24601 (N_24601,N_18221,N_18132);
nand U24602 (N_24602,N_17707,N_15523);
nor U24603 (N_24603,N_16071,N_16612);
and U24604 (N_24604,N_19879,N_19684);
or U24605 (N_24605,N_15248,N_17565);
or U24606 (N_24606,N_15796,N_15527);
nor U24607 (N_24607,N_19943,N_19368);
nor U24608 (N_24608,N_15696,N_19392);
nand U24609 (N_24609,N_19910,N_17400);
nor U24610 (N_24610,N_19869,N_17033);
nor U24611 (N_24611,N_17563,N_18804);
xor U24612 (N_24612,N_16413,N_15015);
or U24613 (N_24613,N_15416,N_17203);
or U24614 (N_24614,N_16144,N_16718);
or U24615 (N_24615,N_17501,N_18563);
nand U24616 (N_24616,N_17941,N_16784);
and U24617 (N_24617,N_17410,N_17094);
nand U24618 (N_24618,N_18998,N_17404);
and U24619 (N_24619,N_17304,N_19850);
nor U24620 (N_24620,N_19991,N_16363);
or U24621 (N_24621,N_15580,N_17601);
and U24622 (N_24622,N_15035,N_17502);
nand U24623 (N_24623,N_19367,N_16029);
and U24624 (N_24624,N_17235,N_18397);
nor U24625 (N_24625,N_18339,N_16159);
and U24626 (N_24626,N_16110,N_19652);
xor U24627 (N_24627,N_18138,N_18010);
nand U24628 (N_24628,N_16410,N_17809);
or U24629 (N_24629,N_19615,N_15385);
or U24630 (N_24630,N_19124,N_16705);
xnor U24631 (N_24631,N_17398,N_17609);
xnor U24632 (N_24632,N_17358,N_19186);
nor U24633 (N_24633,N_17205,N_15485);
nand U24634 (N_24634,N_19863,N_15511);
or U24635 (N_24635,N_15412,N_15507);
nor U24636 (N_24636,N_17961,N_15470);
nand U24637 (N_24637,N_17513,N_19528);
or U24638 (N_24638,N_17253,N_15729);
nor U24639 (N_24639,N_15151,N_18264);
and U24640 (N_24640,N_17721,N_18035);
nand U24641 (N_24641,N_15245,N_15052);
or U24642 (N_24642,N_16120,N_15220);
xnor U24643 (N_24643,N_18039,N_17517);
nand U24644 (N_24644,N_17171,N_15322);
xnor U24645 (N_24645,N_19189,N_15443);
nor U24646 (N_24646,N_15209,N_16043);
nand U24647 (N_24647,N_19132,N_19308);
or U24648 (N_24648,N_19597,N_18782);
nand U24649 (N_24649,N_17424,N_19448);
and U24650 (N_24650,N_15013,N_18327);
xnor U24651 (N_24651,N_18452,N_16611);
and U24652 (N_24652,N_16013,N_16557);
nand U24653 (N_24653,N_16578,N_16984);
nor U24654 (N_24654,N_18489,N_18285);
nand U24655 (N_24655,N_17931,N_19699);
or U24656 (N_24656,N_16080,N_15090);
nor U24657 (N_24657,N_16172,N_18148);
and U24658 (N_24658,N_15779,N_16366);
and U24659 (N_24659,N_17850,N_16873);
or U24660 (N_24660,N_15741,N_19051);
and U24661 (N_24661,N_15403,N_18478);
nor U24662 (N_24662,N_18053,N_17828);
and U24663 (N_24663,N_18977,N_15963);
and U24664 (N_24664,N_16696,N_17637);
xnor U24665 (N_24665,N_17912,N_16757);
and U24666 (N_24666,N_17115,N_16199);
and U24667 (N_24667,N_15186,N_19424);
xnor U24668 (N_24668,N_17222,N_17727);
nand U24669 (N_24669,N_15000,N_16199);
nor U24670 (N_24670,N_19419,N_15433);
nand U24671 (N_24671,N_17191,N_19388);
or U24672 (N_24672,N_16872,N_18787);
xnor U24673 (N_24673,N_15886,N_19361);
and U24674 (N_24674,N_17408,N_18246);
nor U24675 (N_24675,N_16943,N_19095);
or U24676 (N_24676,N_19952,N_17744);
and U24677 (N_24677,N_15538,N_15484);
or U24678 (N_24678,N_18333,N_16342);
nor U24679 (N_24679,N_18829,N_15557);
and U24680 (N_24680,N_15442,N_15075);
nand U24681 (N_24681,N_18773,N_15264);
nor U24682 (N_24682,N_17355,N_19832);
nor U24683 (N_24683,N_16954,N_18699);
or U24684 (N_24684,N_15769,N_15600);
nand U24685 (N_24685,N_15751,N_17847);
xor U24686 (N_24686,N_18075,N_17118);
xor U24687 (N_24687,N_16331,N_19349);
and U24688 (N_24688,N_15232,N_15537);
and U24689 (N_24689,N_15889,N_19294);
or U24690 (N_24690,N_16111,N_16873);
and U24691 (N_24691,N_17772,N_15831);
and U24692 (N_24692,N_18789,N_18948);
or U24693 (N_24693,N_17057,N_17429);
nand U24694 (N_24694,N_18101,N_16498);
nor U24695 (N_24695,N_17543,N_19473);
nor U24696 (N_24696,N_15037,N_16515);
or U24697 (N_24697,N_19831,N_19388);
nor U24698 (N_24698,N_16473,N_15352);
and U24699 (N_24699,N_18100,N_18619);
nand U24700 (N_24700,N_16695,N_17907);
nor U24701 (N_24701,N_17991,N_16946);
nand U24702 (N_24702,N_18900,N_16997);
nand U24703 (N_24703,N_18372,N_15759);
nor U24704 (N_24704,N_15561,N_17062);
and U24705 (N_24705,N_17320,N_16531);
nor U24706 (N_24706,N_16272,N_16925);
xor U24707 (N_24707,N_16885,N_15435);
and U24708 (N_24708,N_16403,N_17443);
xnor U24709 (N_24709,N_15645,N_16933);
nand U24710 (N_24710,N_15244,N_15438);
xor U24711 (N_24711,N_19339,N_17694);
nand U24712 (N_24712,N_17306,N_17038);
or U24713 (N_24713,N_19223,N_17748);
and U24714 (N_24714,N_15974,N_15910);
nand U24715 (N_24715,N_16457,N_15012);
and U24716 (N_24716,N_16425,N_17117);
nor U24717 (N_24717,N_15404,N_17851);
nor U24718 (N_24718,N_19192,N_19551);
or U24719 (N_24719,N_16754,N_17666);
and U24720 (N_24720,N_19323,N_18312);
nor U24721 (N_24721,N_16449,N_15290);
nand U24722 (N_24722,N_19643,N_17541);
or U24723 (N_24723,N_19714,N_16223);
nor U24724 (N_24724,N_16965,N_19259);
nand U24725 (N_24725,N_18089,N_18346);
xor U24726 (N_24726,N_15313,N_18063);
nor U24727 (N_24727,N_17455,N_15111);
or U24728 (N_24728,N_15999,N_17960);
xnor U24729 (N_24729,N_16439,N_15074);
xnor U24730 (N_24730,N_19458,N_17250);
and U24731 (N_24731,N_16760,N_15937);
or U24732 (N_24732,N_17138,N_18326);
or U24733 (N_24733,N_19404,N_19086);
nor U24734 (N_24734,N_19700,N_18050);
xor U24735 (N_24735,N_16201,N_18063);
nand U24736 (N_24736,N_15396,N_19717);
xor U24737 (N_24737,N_17568,N_15640);
xor U24738 (N_24738,N_19066,N_17231);
nor U24739 (N_24739,N_18970,N_17049);
nor U24740 (N_24740,N_18201,N_15452);
and U24741 (N_24741,N_17691,N_15762);
and U24742 (N_24742,N_15443,N_18003);
nand U24743 (N_24743,N_18228,N_16090);
xor U24744 (N_24744,N_17943,N_17011);
or U24745 (N_24745,N_16982,N_18892);
nand U24746 (N_24746,N_15869,N_18447);
xor U24747 (N_24747,N_19005,N_15310);
or U24748 (N_24748,N_19121,N_18156);
nor U24749 (N_24749,N_18328,N_17235);
xnor U24750 (N_24750,N_16050,N_15094);
and U24751 (N_24751,N_17974,N_18596);
or U24752 (N_24752,N_18514,N_15132);
nand U24753 (N_24753,N_17713,N_16541);
or U24754 (N_24754,N_15112,N_16741);
or U24755 (N_24755,N_18495,N_19681);
and U24756 (N_24756,N_19954,N_16535);
nor U24757 (N_24757,N_17348,N_18176);
xor U24758 (N_24758,N_17941,N_16992);
and U24759 (N_24759,N_19791,N_16858);
and U24760 (N_24760,N_19354,N_17607);
xnor U24761 (N_24761,N_16803,N_18443);
nand U24762 (N_24762,N_19055,N_19227);
and U24763 (N_24763,N_18778,N_18092);
nor U24764 (N_24764,N_18243,N_18352);
nand U24765 (N_24765,N_17783,N_15624);
xor U24766 (N_24766,N_17311,N_18681);
nor U24767 (N_24767,N_15889,N_18851);
xor U24768 (N_24768,N_15483,N_16338);
nand U24769 (N_24769,N_16752,N_18448);
nor U24770 (N_24770,N_15114,N_18912);
or U24771 (N_24771,N_15372,N_18586);
xnor U24772 (N_24772,N_19098,N_19810);
or U24773 (N_24773,N_15169,N_19979);
nor U24774 (N_24774,N_17864,N_19145);
or U24775 (N_24775,N_17681,N_19392);
or U24776 (N_24776,N_18335,N_19102);
or U24777 (N_24777,N_15829,N_16533);
or U24778 (N_24778,N_17403,N_16738);
nor U24779 (N_24779,N_18743,N_19733);
xor U24780 (N_24780,N_16724,N_16723);
xnor U24781 (N_24781,N_18831,N_16995);
xnor U24782 (N_24782,N_17482,N_16167);
or U24783 (N_24783,N_16847,N_18054);
xor U24784 (N_24784,N_17933,N_15257);
nand U24785 (N_24785,N_17640,N_19114);
or U24786 (N_24786,N_16015,N_18289);
nor U24787 (N_24787,N_15033,N_15051);
xor U24788 (N_24788,N_15540,N_19941);
or U24789 (N_24789,N_17655,N_16221);
nor U24790 (N_24790,N_15578,N_18829);
and U24791 (N_24791,N_16198,N_18569);
and U24792 (N_24792,N_18239,N_16547);
nor U24793 (N_24793,N_18938,N_18506);
nand U24794 (N_24794,N_16485,N_18593);
nand U24795 (N_24795,N_15216,N_17175);
nor U24796 (N_24796,N_17933,N_15184);
and U24797 (N_24797,N_17224,N_17108);
nor U24798 (N_24798,N_17685,N_16617);
and U24799 (N_24799,N_16019,N_16153);
nand U24800 (N_24800,N_17171,N_16049);
nor U24801 (N_24801,N_18518,N_18766);
or U24802 (N_24802,N_18329,N_17240);
xnor U24803 (N_24803,N_15772,N_16965);
xnor U24804 (N_24804,N_17170,N_19115);
or U24805 (N_24805,N_17571,N_18542);
nor U24806 (N_24806,N_19846,N_19580);
nor U24807 (N_24807,N_17772,N_17600);
nand U24808 (N_24808,N_17196,N_15551);
nor U24809 (N_24809,N_19175,N_19682);
nand U24810 (N_24810,N_17561,N_16376);
or U24811 (N_24811,N_16310,N_19105);
and U24812 (N_24812,N_18802,N_19135);
xnor U24813 (N_24813,N_19778,N_15730);
xnor U24814 (N_24814,N_15855,N_15345);
nor U24815 (N_24815,N_19096,N_17889);
xnor U24816 (N_24816,N_17139,N_16938);
or U24817 (N_24817,N_17459,N_15424);
nor U24818 (N_24818,N_17825,N_17393);
xor U24819 (N_24819,N_17393,N_17733);
xnor U24820 (N_24820,N_16627,N_15371);
or U24821 (N_24821,N_18848,N_16669);
nor U24822 (N_24822,N_17743,N_16513);
or U24823 (N_24823,N_18953,N_16979);
and U24824 (N_24824,N_17926,N_19969);
or U24825 (N_24825,N_17921,N_19686);
and U24826 (N_24826,N_15620,N_19156);
or U24827 (N_24827,N_18000,N_17334);
nand U24828 (N_24828,N_17402,N_18810);
or U24829 (N_24829,N_17510,N_16774);
and U24830 (N_24830,N_17315,N_19987);
nand U24831 (N_24831,N_18675,N_19565);
xnor U24832 (N_24832,N_16618,N_18067);
nand U24833 (N_24833,N_16020,N_15844);
and U24834 (N_24834,N_17700,N_16162);
and U24835 (N_24835,N_16584,N_19793);
nand U24836 (N_24836,N_17781,N_16360);
nor U24837 (N_24837,N_18872,N_19907);
nand U24838 (N_24838,N_19101,N_15950);
or U24839 (N_24839,N_18698,N_16132);
xnor U24840 (N_24840,N_19792,N_15520);
and U24841 (N_24841,N_19674,N_19351);
and U24842 (N_24842,N_19399,N_17418);
nand U24843 (N_24843,N_17459,N_15171);
or U24844 (N_24844,N_16461,N_18720);
and U24845 (N_24845,N_16937,N_16132);
xor U24846 (N_24846,N_15905,N_19990);
or U24847 (N_24847,N_17105,N_17339);
nand U24848 (N_24848,N_16150,N_17081);
xnor U24849 (N_24849,N_18122,N_19083);
and U24850 (N_24850,N_17106,N_19630);
nor U24851 (N_24851,N_16765,N_17032);
nand U24852 (N_24852,N_18120,N_15497);
xor U24853 (N_24853,N_17850,N_18593);
xnor U24854 (N_24854,N_19728,N_17348);
nand U24855 (N_24855,N_15617,N_18988);
nor U24856 (N_24856,N_18843,N_19436);
xnor U24857 (N_24857,N_18023,N_19178);
or U24858 (N_24858,N_19417,N_15617);
or U24859 (N_24859,N_15870,N_19416);
or U24860 (N_24860,N_18011,N_18016);
xnor U24861 (N_24861,N_16087,N_19599);
and U24862 (N_24862,N_16881,N_18572);
nor U24863 (N_24863,N_19419,N_19207);
nand U24864 (N_24864,N_18146,N_17815);
xnor U24865 (N_24865,N_18968,N_15129);
xor U24866 (N_24866,N_19509,N_18293);
or U24867 (N_24867,N_15433,N_15976);
nor U24868 (N_24868,N_16716,N_18119);
nand U24869 (N_24869,N_15112,N_17194);
and U24870 (N_24870,N_17219,N_16304);
xnor U24871 (N_24871,N_17026,N_16004);
nor U24872 (N_24872,N_18190,N_18041);
nand U24873 (N_24873,N_15870,N_18455);
and U24874 (N_24874,N_16749,N_16740);
and U24875 (N_24875,N_17785,N_16357);
xnor U24876 (N_24876,N_15881,N_15369);
or U24877 (N_24877,N_15515,N_16006);
xor U24878 (N_24878,N_18204,N_16648);
nand U24879 (N_24879,N_18968,N_19465);
or U24880 (N_24880,N_16729,N_19821);
xnor U24881 (N_24881,N_18189,N_16173);
nor U24882 (N_24882,N_19145,N_16759);
xnor U24883 (N_24883,N_17876,N_16808);
nor U24884 (N_24884,N_18121,N_19186);
xor U24885 (N_24885,N_19406,N_17218);
or U24886 (N_24886,N_16288,N_19737);
nor U24887 (N_24887,N_16049,N_15050);
and U24888 (N_24888,N_15536,N_17126);
nor U24889 (N_24889,N_18465,N_15019);
or U24890 (N_24890,N_19514,N_17484);
nand U24891 (N_24891,N_18522,N_15930);
nor U24892 (N_24892,N_16098,N_15095);
nor U24893 (N_24893,N_16586,N_16725);
xor U24894 (N_24894,N_16761,N_19575);
nor U24895 (N_24895,N_17120,N_17101);
or U24896 (N_24896,N_19077,N_18354);
nor U24897 (N_24897,N_16149,N_15349);
and U24898 (N_24898,N_15216,N_19643);
and U24899 (N_24899,N_15514,N_17499);
or U24900 (N_24900,N_16403,N_17519);
nand U24901 (N_24901,N_17050,N_15543);
xnor U24902 (N_24902,N_19662,N_18371);
nand U24903 (N_24903,N_18585,N_16275);
xor U24904 (N_24904,N_19126,N_16518);
or U24905 (N_24905,N_15979,N_19503);
nor U24906 (N_24906,N_16204,N_17345);
and U24907 (N_24907,N_15154,N_19823);
nand U24908 (N_24908,N_15227,N_15000);
nor U24909 (N_24909,N_17606,N_17823);
xor U24910 (N_24910,N_17103,N_16802);
nand U24911 (N_24911,N_15042,N_17200);
nand U24912 (N_24912,N_16764,N_17704);
and U24913 (N_24913,N_17458,N_19147);
or U24914 (N_24914,N_17630,N_18472);
nand U24915 (N_24915,N_17907,N_19420);
xnor U24916 (N_24916,N_17537,N_15614);
nand U24917 (N_24917,N_16255,N_17731);
or U24918 (N_24918,N_18684,N_15584);
and U24919 (N_24919,N_18809,N_17663);
xor U24920 (N_24920,N_16669,N_19973);
nor U24921 (N_24921,N_16681,N_15115);
nand U24922 (N_24922,N_16381,N_19655);
nor U24923 (N_24923,N_16961,N_15044);
nand U24924 (N_24924,N_17026,N_16972);
or U24925 (N_24925,N_18998,N_18169);
nand U24926 (N_24926,N_16181,N_16654);
and U24927 (N_24927,N_18842,N_16948);
nand U24928 (N_24928,N_19868,N_17389);
nor U24929 (N_24929,N_16314,N_16595);
and U24930 (N_24930,N_19878,N_17686);
or U24931 (N_24931,N_16678,N_15476);
nand U24932 (N_24932,N_18338,N_15237);
or U24933 (N_24933,N_18582,N_18948);
nand U24934 (N_24934,N_17325,N_18722);
or U24935 (N_24935,N_19636,N_19314);
nand U24936 (N_24936,N_18540,N_17136);
and U24937 (N_24937,N_15934,N_18608);
nor U24938 (N_24938,N_17090,N_15105);
xor U24939 (N_24939,N_17459,N_17596);
nand U24940 (N_24940,N_15358,N_17059);
xor U24941 (N_24941,N_15464,N_18341);
nand U24942 (N_24942,N_19993,N_16115);
and U24943 (N_24943,N_18123,N_15845);
and U24944 (N_24944,N_17213,N_17149);
and U24945 (N_24945,N_15940,N_18235);
nor U24946 (N_24946,N_16093,N_19808);
and U24947 (N_24947,N_17506,N_18896);
nand U24948 (N_24948,N_18837,N_19678);
xor U24949 (N_24949,N_17516,N_19463);
or U24950 (N_24950,N_17211,N_15625);
or U24951 (N_24951,N_17507,N_16389);
xor U24952 (N_24952,N_16121,N_19050);
nand U24953 (N_24953,N_15660,N_15139);
xor U24954 (N_24954,N_17235,N_18641);
xor U24955 (N_24955,N_19673,N_15741);
nor U24956 (N_24956,N_15228,N_17940);
nand U24957 (N_24957,N_17555,N_17745);
xor U24958 (N_24958,N_16225,N_17696);
nor U24959 (N_24959,N_19994,N_17607);
nand U24960 (N_24960,N_16191,N_19443);
or U24961 (N_24961,N_15128,N_15433);
nor U24962 (N_24962,N_18170,N_16108);
nand U24963 (N_24963,N_17022,N_16054);
xnor U24964 (N_24964,N_15026,N_16426);
nand U24965 (N_24965,N_18601,N_17744);
nor U24966 (N_24966,N_16901,N_15655);
nor U24967 (N_24967,N_15492,N_18254);
and U24968 (N_24968,N_19238,N_17375);
xor U24969 (N_24969,N_17216,N_16465);
or U24970 (N_24970,N_16018,N_18924);
nor U24971 (N_24971,N_19916,N_15176);
nand U24972 (N_24972,N_15164,N_16343);
and U24973 (N_24973,N_15892,N_18619);
nand U24974 (N_24974,N_19953,N_16712);
nor U24975 (N_24975,N_19485,N_17206);
nand U24976 (N_24976,N_16694,N_17997);
or U24977 (N_24977,N_17740,N_19584);
nand U24978 (N_24978,N_16550,N_16451);
xor U24979 (N_24979,N_15414,N_16002);
nor U24980 (N_24980,N_18891,N_17643);
nand U24981 (N_24981,N_16275,N_15982);
xor U24982 (N_24982,N_19222,N_18454);
or U24983 (N_24983,N_19542,N_15650);
and U24984 (N_24984,N_15309,N_19795);
and U24985 (N_24985,N_19725,N_18729);
nor U24986 (N_24986,N_17168,N_18383);
nand U24987 (N_24987,N_18671,N_17164);
nand U24988 (N_24988,N_18957,N_17769);
and U24989 (N_24989,N_19327,N_18432);
and U24990 (N_24990,N_18915,N_18315);
and U24991 (N_24991,N_17657,N_19804);
and U24992 (N_24992,N_15507,N_19117);
xnor U24993 (N_24993,N_17260,N_16284);
and U24994 (N_24994,N_16602,N_18369);
nand U24995 (N_24995,N_18151,N_15663);
xnor U24996 (N_24996,N_18678,N_16763);
and U24997 (N_24997,N_16205,N_18162);
nand U24998 (N_24998,N_17704,N_17088);
nand U24999 (N_24999,N_17363,N_17574);
or UO_0 (O_0,N_20032,N_22152);
xor UO_1 (O_1,N_23909,N_23534);
or UO_2 (O_2,N_24715,N_20542);
xnor UO_3 (O_3,N_23115,N_24274);
xnor UO_4 (O_4,N_20857,N_21623);
nand UO_5 (O_5,N_22693,N_23623);
or UO_6 (O_6,N_22493,N_22483);
or UO_7 (O_7,N_23143,N_20906);
nand UO_8 (O_8,N_24980,N_21931);
and UO_9 (O_9,N_22123,N_23283);
or UO_10 (O_10,N_20125,N_20836);
nand UO_11 (O_11,N_20081,N_20193);
and UO_12 (O_12,N_23767,N_22443);
nor UO_13 (O_13,N_20681,N_21972);
nand UO_14 (O_14,N_22830,N_21026);
or UO_15 (O_15,N_22220,N_21270);
nand UO_16 (O_16,N_20863,N_21332);
xor UO_17 (O_17,N_23768,N_20053);
and UO_18 (O_18,N_22634,N_24519);
xor UO_19 (O_19,N_22622,N_22130);
nor UO_20 (O_20,N_22743,N_21066);
or UO_21 (O_21,N_24590,N_23914);
and UO_22 (O_22,N_24101,N_20262);
nand UO_23 (O_23,N_24887,N_21017);
nand UO_24 (O_24,N_24393,N_20217);
nand UO_25 (O_25,N_21728,N_24561);
or UO_26 (O_26,N_20566,N_22770);
nand UO_27 (O_27,N_23126,N_20226);
nor UO_28 (O_28,N_21885,N_24382);
nor UO_29 (O_29,N_20517,N_24771);
or UO_30 (O_30,N_21639,N_20170);
nor UO_31 (O_31,N_21629,N_21587);
nor UO_32 (O_32,N_20908,N_23228);
nor UO_33 (O_33,N_21707,N_20143);
and UO_34 (O_34,N_23159,N_23320);
xor UO_35 (O_35,N_20813,N_23625);
or UO_36 (O_36,N_24939,N_21665);
or UO_37 (O_37,N_21459,N_24554);
xnor UO_38 (O_38,N_23619,N_24117);
and UO_39 (O_39,N_20645,N_23028);
nand UO_40 (O_40,N_24791,N_23483);
or UO_41 (O_41,N_23992,N_23217);
nor UO_42 (O_42,N_24605,N_24768);
or UO_43 (O_43,N_22313,N_22887);
nand UO_44 (O_44,N_23931,N_20151);
nand UO_45 (O_45,N_23564,N_23803);
nand UO_46 (O_46,N_20780,N_22749);
and UO_47 (O_47,N_22427,N_20690);
or UO_48 (O_48,N_24483,N_23363);
or UO_49 (O_49,N_24159,N_23955);
nand UO_50 (O_50,N_22324,N_24500);
xnor UO_51 (O_51,N_20489,N_21435);
and UO_52 (O_52,N_20460,N_24754);
and UO_53 (O_53,N_21911,N_22103);
or UO_54 (O_54,N_20046,N_21801);
nor UO_55 (O_55,N_20753,N_23740);
xor UO_56 (O_56,N_24787,N_24343);
xnor UO_57 (O_57,N_22078,N_24612);
xnor UO_58 (O_58,N_23342,N_21797);
nor UO_59 (O_59,N_21325,N_22282);
nand UO_60 (O_60,N_21679,N_20686);
and UO_61 (O_61,N_20812,N_23107);
nand UO_62 (O_62,N_21859,N_21544);
nand UO_63 (O_63,N_20253,N_21958);
xor UO_64 (O_64,N_23090,N_21499);
and UO_65 (O_65,N_23116,N_21539);
xnor UO_66 (O_66,N_22149,N_21567);
nor UO_67 (O_67,N_20414,N_22730);
nor UO_68 (O_68,N_22416,N_24462);
or UO_69 (O_69,N_21365,N_20286);
and UO_70 (O_70,N_20565,N_24060);
nand UO_71 (O_71,N_22285,N_23469);
xnor UO_72 (O_72,N_24140,N_20959);
nand UO_73 (O_73,N_21334,N_21263);
nor UO_74 (O_74,N_21526,N_21158);
or UO_75 (O_75,N_22609,N_22092);
nor UO_76 (O_76,N_20385,N_21099);
and UO_77 (O_77,N_20169,N_21530);
xnor UO_78 (O_78,N_24183,N_20149);
nor UO_79 (O_79,N_21234,N_23275);
nand UO_80 (O_80,N_21515,N_22517);
or UO_81 (O_81,N_23349,N_22806);
xnor UO_82 (O_82,N_22060,N_20982);
nor UO_83 (O_83,N_22237,N_23908);
or UO_84 (O_84,N_23950,N_23423);
xnor UO_85 (O_85,N_24824,N_20706);
xnor UO_86 (O_86,N_22071,N_24610);
and UO_87 (O_87,N_23970,N_20280);
or UO_88 (O_88,N_20096,N_20790);
and UO_89 (O_89,N_24722,N_22426);
or UO_90 (O_90,N_21032,N_21422);
and UO_91 (O_91,N_21531,N_22450);
xnor UO_92 (O_92,N_21632,N_23451);
and UO_93 (O_93,N_21177,N_20332);
xnor UO_94 (O_94,N_24852,N_23581);
or UO_95 (O_95,N_20202,N_21509);
nor UO_96 (O_96,N_22172,N_21864);
xor UO_97 (O_97,N_21252,N_22655);
xor UO_98 (O_98,N_21759,N_21602);
nand UO_99 (O_99,N_23114,N_24220);
nor UO_100 (O_100,N_20055,N_22750);
nor UO_101 (O_101,N_22341,N_23051);
nand UO_102 (O_102,N_21312,N_23954);
and UO_103 (O_103,N_21605,N_20549);
and UO_104 (O_104,N_24224,N_20709);
or UO_105 (O_105,N_20189,N_23464);
nor UO_106 (O_106,N_23396,N_23138);
or UO_107 (O_107,N_22533,N_23403);
or UO_108 (O_108,N_23073,N_21412);
and UO_109 (O_109,N_20688,N_21863);
or UO_110 (O_110,N_22320,N_21329);
or UO_111 (O_111,N_23836,N_22036);
nor UO_112 (O_112,N_20864,N_23498);
or UO_113 (O_113,N_22304,N_21411);
and UO_114 (O_114,N_20590,N_20054);
nor UO_115 (O_115,N_21829,N_23795);
or UO_116 (O_116,N_22618,N_21782);
and UO_117 (O_117,N_23134,N_24482);
and UO_118 (O_118,N_20958,N_21837);
and UO_119 (O_119,N_22265,N_22811);
nand UO_120 (O_120,N_24489,N_22175);
and UO_121 (O_121,N_24576,N_24405);
and UO_122 (O_122,N_21558,N_20601);
nand UO_123 (O_123,N_21193,N_22727);
xor UO_124 (O_124,N_21153,N_22917);
nand UO_125 (O_125,N_20713,N_20150);
and UO_126 (O_126,N_22289,N_21283);
and UO_127 (O_127,N_22291,N_20683);
nand UO_128 (O_128,N_22494,N_22751);
or UO_129 (O_129,N_23798,N_20402);
xor UO_130 (O_130,N_24777,N_20817);
nor UO_131 (O_131,N_22260,N_24734);
or UO_132 (O_132,N_23818,N_24627);
nor UO_133 (O_133,N_23250,N_21488);
nand UO_134 (O_134,N_23573,N_22512);
and UO_135 (O_135,N_22045,N_22561);
nor UO_136 (O_136,N_21615,N_20399);
nor UO_137 (O_137,N_22501,N_20341);
xor UO_138 (O_138,N_20871,N_22733);
xnor UO_139 (O_139,N_23742,N_24982);
nor UO_140 (O_140,N_20545,N_24319);
nor UO_141 (O_141,N_24935,N_23405);
nand UO_142 (O_142,N_20437,N_22183);
xor UO_143 (O_143,N_20120,N_23121);
and UO_144 (O_144,N_20249,N_23269);
nor UO_145 (O_145,N_20581,N_21890);
nor UO_146 (O_146,N_22127,N_21470);
xnor UO_147 (O_147,N_20877,N_24179);
nand UO_148 (O_148,N_21142,N_20995);
xnor UO_149 (O_149,N_20702,N_22214);
and UO_150 (O_150,N_21789,N_21727);
nand UO_151 (O_151,N_20670,N_20167);
and UO_152 (O_152,N_23639,N_20598);
nor UO_153 (O_153,N_23720,N_24602);
or UO_154 (O_154,N_21266,N_22335);
nand UO_155 (O_155,N_20388,N_22241);
or UO_156 (O_156,N_21937,N_24637);
nand UO_157 (O_157,N_24431,N_22596);
xor UO_158 (O_158,N_24424,N_24296);
or UO_159 (O_159,N_23685,N_23050);
nand UO_160 (O_160,N_20177,N_21200);
nand UO_161 (O_161,N_22467,N_23313);
nor UO_162 (O_162,N_23709,N_21658);
xnor UO_163 (O_163,N_21956,N_22570);
and UO_164 (O_164,N_22857,N_20572);
or UO_165 (O_165,N_21192,N_21477);
or UO_166 (O_166,N_23728,N_21597);
or UO_167 (O_167,N_24430,N_21216);
nor UO_168 (O_168,N_23786,N_20458);
nor UO_169 (O_169,N_20365,N_21140);
and UO_170 (O_170,N_21381,N_22620);
nor UO_171 (O_171,N_23062,N_22197);
or UO_172 (O_172,N_24732,N_20553);
or UO_173 (O_173,N_22038,N_24608);
xnor UO_174 (O_174,N_21022,N_23174);
xor UO_175 (O_175,N_21591,N_24081);
nor UO_176 (O_176,N_23177,N_22943);
nand UO_177 (O_177,N_22367,N_21380);
xnor UO_178 (O_178,N_20792,N_22336);
and UO_179 (O_179,N_23359,N_24469);
xor UO_180 (O_180,N_21982,N_20378);
and UO_181 (O_181,N_20778,N_24024);
or UO_182 (O_182,N_24166,N_22621);
xor UO_183 (O_183,N_22772,N_24978);
nor UO_184 (O_184,N_24619,N_22781);
nand UO_185 (O_185,N_22039,N_21923);
nand UO_186 (O_186,N_23086,N_23360);
and UO_187 (O_187,N_20000,N_24423);
or UO_188 (O_188,N_21028,N_20676);
xor UO_189 (O_189,N_24169,N_24510);
and UO_190 (O_190,N_24273,N_22072);
nor UO_191 (O_191,N_23297,N_24069);
nor UO_192 (O_192,N_23777,N_24257);
or UO_193 (O_193,N_24281,N_22064);
or UO_194 (O_194,N_24654,N_20219);
xnor UO_195 (O_195,N_21966,N_20756);
or UO_196 (O_196,N_20712,N_22185);
nor UO_197 (O_197,N_23976,N_20218);
nand UO_198 (O_198,N_23630,N_22852);
nand UO_199 (O_199,N_20016,N_21408);
or UO_200 (O_200,N_20939,N_22835);
and UO_201 (O_201,N_20256,N_24435);
xnor UO_202 (O_202,N_20865,N_23353);
or UO_203 (O_203,N_22745,N_23773);
xor UO_204 (O_204,N_22877,N_24243);
nor UO_205 (O_205,N_22774,N_20070);
and UO_206 (O_206,N_20154,N_24105);
xnor UO_207 (O_207,N_22980,N_21749);
nor UO_208 (O_208,N_20384,N_21571);
and UO_209 (O_209,N_23233,N_22714);
or UO_210 (O_210,N_24763,N_21869);
xnor UO_211 (O_211,N_24841,N_23856);
and UO_212 (O_212,N_23104,N_20456);
or UO_213 (O_213,N_20108,N_23435);
nand UO_214 (O_214,N_20704,N_24376);
and UO_215 (O_215,N_21154,N_23910);
xor UO_216 (O_216,N_23617,N_23157);
and UO_217 (O_217,N_24476,N_24966);
nor UO_218 (O_218,N_24641,N_22004);
and UO_219 (O_219,N_24097,N_23817);
xor UO_220 (O_220,N_23670,N_22870);
xnor UO_221 (O_221,N_22721,N_20038);
nand UO_222 (O_222,N_24156,N_23397);
or UO_223 (O_223,N_23788,N_24357);
and UO_224 (O_224,N_24956,N_24917);
or UO_225 (O_225,N_20602,N_22627);
nand UO_226 (O_226,N_23289,N_23632);
xor UO_227 (O_227,N_23301,N_20976);
nor UO_228 (O_228,N_23198,N_23354);
xnor UO_229 (O_229,N_22025,N_24538);
nand UO_230 (O_230,N_24594,N_21672);
nand UO_231 (O_231,N_24297,N_20068);
nor UO_232 (O_232,N_20354,N_22742);
nor UO_233 (O_233,N_21160,N_23013);
nand UO_234 (O_234,N_20503,N_22171);
and UO_235 (O_235,N_20749,N_22178);
nor UO_236 (O_236,N_24983,N_23902);
and UO_237 (O_237,N_21725,N_20555);
or UO_238 (O_238,N_22195,N_22272);
nor UO_239 (O_239,N_22976,N_20795);
nor UO_240 (O_240,N_23002,N_22194);
xor UO_241 (O_241,N_24968,N_24134);
xor UO_242 (O_242,N_20158,N_24813);
xor UO_243 (O_243,N_21218,N_21370);
nand UO_244 (O_244,N_22507,N_21547);
and UO_245 (O_245,N_20404,N_24672);
and UO_246 (O_246,N_23443,N_23333);
or UO_247 (O_247,N_22020,N_24525);
and UO_248 (O_248,N_21141,N_23061);
xnor UO_249 (O_249,N_22484,N_20040);
and UO_250 (O_250,N_21167,N_24713);
nand UO_251 (O_251,N_21985,N_23142);
or UO_252 (O_252,N_21290,N_24491);
xnor UO_253 (O_253,N_22221,N_21851);
or UO_254 (O_254,N_24816,N_23085);
and UO_255 (O_255,N_21085,N_23189);
xnor UO_256 (O_256,N_24304,N_23109);
xnor UO_257 (O_257,N_20396,N_20944);
and UO_258 (O_258,N_21903,N_20429);
xnor UO_259 (O_259,N_22048,N_22002);
nor UO_260 (O_260,N_23094,N_21722);
nand UO_261 (O_261,N_22170,N_20344);
and UO_262 (O_262,N_23980,N_20714);
or UO_263 (O_263,N_20299,N_20273);
or UO_264 (O_264,N_20515,N_23937);
nor UO_265 (O_265,N_20692,N_23430);
nor UO_266 (O_266,N_20471,N_20094);
nand UO_267 (O_267,N_23668,N_22334);
nor UO_268 (O_268,N_22584,N_22710);
or UO_269 (O_269,N_23848,N_20392);
nor UO_270 (O_270,N_20201,N_22018);
and UO_271 (O_271,N_20236,N_24679);
nor UO_272 (O_272,N_21950,N_21814);
or UO_273 (O_273,N_24905,N_20754);
nand UO_274 (O_274,N_20058,N_24217);
nand UO_275 (O_275,N_24401,N_23338);
xor UO_276 (O_276,N_22227,N_24616);
nand UO_277 (O_277,N_21399,N_20381);
nand UO_278 (O_278,N_23277,N_21720);
and UO_279 (O_279,N_22274,N_21339);
nor UO_280 (O_280,N_20786,N_22053);
nor UO_281 (O_281,N_21278,N_24687);
and UO_282 (O_282,N_22496,N_20905);
nor UO_283 (O_283,N_22682,N_21304);
xor UO_284 (O_284,N_22856,N_24459);
and UO_285 (O_285,N_24830,N_23305);
nor UO_286 (O_286,N_21005,N_22906);
xnor UO_287 (O_287,N_21616,N_21137);
xor UO_288 (O_288,N_23854,N_20793);
xor UO_289 (O_289,N_22791,N_22793);
and UO_290 (O_290,N_21425,N_20333);
or UO_291 (O_291,N_22333,N_24766);
nand UO_292 (O_292,N_20057,N_24667);
or UO_293 (O_293,N_21319,N_23330);
and UO_294 (O_294,N_24969,N_24542);
nor UO_295 (O_295,N_22563,N_24829);
xor UO_296 (O_296,N_20407,N_21996);
xnor UO_297 (O_297,N_24848,N_24564);
xnor UO_298 (O_298,N_21806,N_24248);
xnor UO_299 (O_299,N_21166,N_21913);
nor UO_300 (O_300,N_23102,N_21008);
and UO_301 (O_301,N_23234,N_20675);
nor UO_302 (O_302,N_23493,N_21702);
and UO_303 (O_303,N_23331,N_23997);
or UO_304 (O_304,N_24014,N_21767);
or UO_305 (O_305,N_23745,N_24827);
nand UO_306 (O_306,N_22753,N_21293);
and UO_307 (O_307,N_21264,N_24575);
nand UO_308 (O_308,N_23473,N_24515);
nor UO_309 (O_309,N_21036,N_21955);
xnor UO_310 (O_310,N_24936,N_20853);
or UO_311 (O_311,N_22595,N_23667);
or UO_312 (O_312,N_24387,N_23064);
nand UO_313 (O_313,N_23302,N_20530);
nand UO_314 (O_314,N_22641,N_24316);
nor UO_315 (O_315,N_23265,N_23928);
nor UO_316 (O_316,N_24417,N_21345);
nor UO_317 (O_317,N_21687,N_22810);
or UO_318 (O_318,N_24571,N_24863);
nor UO_319 (O_319,N_20575,N_20708);
and UO_320 (O_320,N_22046,N_20130);
nand UO_321 (O_321,N_23763,N_22579);
and UO_322 (O_322,N_24184,N_23059);
nand UO_323 (O_323,N_22514,N_21900);
xnor UO_324 (O_324,N_22700,N_20584);
nor UO_325 (O_325,N_22722,N_23465);
nand UO_326 (O_326,N_21667,N_20508);
xnor UO_327 (O_327,N_20470,N_23514);
xnor UO_328 (O_328,N_24632,N_21841);
xor UO_329 (O_329,N_23551,N_24262);
nand UO_330 (O_330,N_21635,N_20020);
nand UO_331 (O_331,N_21291,N_23404);
and UO_332 (O_332,N_21506,N_20306);
and UO_333 (O_333,N_21272,N_21092);
and UO_334 (O_334,N_22407,N_22669);
nand UO_335 (O_335,N_22628,N_21211);
and UO_336 (O_336,N_23318,N_20535);
xnor UO_337 (O_337,N_24981,N_20629);
nand UO_338 (O_338,N_24256,N_24651);
or UO_339 (O_339,N_20486,N_20611);
xnor UO_340 (O_340,N_20736,N_24840);
and UO_341 (O_341,N_23470,N_23251);
and UO_342 (O_342,N_21152,N_20438);
or UO_343 (O_343,N_21525,N_22182);
nor UO_344 (O_344,N_23167,N_21397);
nand UO_345 (O_345,N_23634,N_24909);
xor UO_346 (O_346,N_20375,N_21052);
nor UO_347 (O_347,N_22115,N_21756);
xnor UO_348 (O_348,N_24931,N_20896);
and UO_349 (O_349,N_23292,N_23022);
or UO_350 (O_350,N_24778,N_23647);
or UO_351 (O_351,N_21277,N_21976);
or UO_352 (O_352,N_22586,N_21532);
nor UO_353 (O_353,N_22937,N_23799);
or UO_354 (O_354,N_22211,N_24349);
and UO_355 (O_355,N_23585,N_20580);
and UO_356 (O_356,N_20539,N_24261);
or UO_357 (O_357,N_23247,N_21812);
or UO_358 (O_358,N_24924,N_23479);
xnor UO_359 (O_359,N_24037,N_21969);
xnor UO_360 (O_360,N_20035,N_21289);
xnor UO_361 (O_361,N_22396,N_23590);
xnor UO_362 (O_362,N_21427,N_22112);
xnor UO_363 (O_363,N_21201,N_23426);
xor UO_364 (O_364,N_24109,N_23760);
or UO_365 (O_365,N_21241,N_23546);
and UO_366 (O_366,N_20664,N_20967);
and UO_367 (O_367,N_24888,N_23052);
and UO_368 (O_368,N_23152,N_24221);
xor UO_369 (O_369,N_22399,N_24422);
and UO_370 (O_370,N_24186,N_23759);
nand UO_371 (O_371,N_22853,N_24048);
xor UO_372 (O_372,N_24884,N_21731);
nor UO_373 (O_373,N_22633,N_23082);
or UO_374 (O_374,N_22219,N_20796);
or UO_375 (O_375,N_20705,N_23171);
and UO_376 (O_376,N_20911,N_21057);
and UO_377 (O_377,N_21125,N_23593);
nand UO_378 (O_378,N_22932,N_22780);
xor UO_379 (O_379,N_22264,N_21527);
or UO_380 (O_380,N_23723,N_24825);
nand UO_381 (O_381,N_20733,N_20671);
xor UO_382 (O_382,N_20182,N_21671);
nand UO_383 (O_383,N_23312,N_22307);
and UO_384 (O_384,N_21643,N_21195);
or UO_385 (O_385,N_24959,N_21744);
nor UO_386 (O_386,N_20100,N_23600);
nand UO_387 (O_387,N_21686,N_21986);
nor UO_388 (O_388,N_24901,N_20157);
and UO_389 (O_389,N_21033,N_23232);
nor UO_390 (O_390,N_20131,N_24769);
xnor UO_391 (O_391,N_21662,N_24633);
xor UO_392 (O_392,N_21748,N_23778);
nand UO_393 (O_393,N_20222,N_24514);
nor UO_394 (O_394,N_20400,N_23537);
nor UO_395 (O_395,N_20593,N_24736);
and UO_396 (O_396,N_22992,N_21575);
and UO_397 (O_397,N_20710,N_20875);
and UO_398 (O_398,N_22342,N_21684);
and UO_399 (O_399,N_23553,N_21354);
xnor UO_400 (O_400,N_22097,N_21764);
nand UO_401 (O_401,N_22548,N_24383);
or UO_402 (O_402,N_21469,N_22421);
nand UO_403 (O_403,N_21367,N_23398);
xnor UO_404 (O_404,N_24533,N_20265);
nand UO_405 (O_405,N_24219,N_20652);
and UO_406 (O_406,N_20806,N_24027);
and UO_407 (O_407,N_22317,N_21834);
nand UO_408 (O_408,N_22650,N_23438);
xnor UO_409 (O_409,N_20631,N_24870);
xnor UO_410 (O_410,N_21997,N_24091);
xor UO_411 (O_411,N_23088,N_20428);
nor UO_412 (O_412,N_24820,N_24366);
nand UO_413 (O_413,N_20113,N_23821);
xnor UO_414 (O_414,N_22143,N_21657);
and UO_415 (O_415,N_24615,N_20604);
nor UO_416 (O_416,N_24192,N_21472);
nor UO_417 (O_417,N_20041,N_22480);
or UO_418 (O_418,N_22716,N_24876);
nor UO_419 (O_419,N_23660,N_24558);
nor UO_420 (O_420,N_23717,N_21693);
nand UO_421 (O_421,N_23603,N_24860);
or UO_422 (O_422,N_22973,N_24020);
xor UO_423 (O_423,N_20283,N_22222);
and UO_424 (O_424,N_22569,N_22818);
xnor UO_425 (O_425,N_21134,N_23644);
xnor UO_426 (O_426,N_24292,N_21984);
xnor UO_427 (O_427,N_20453,N_24804);
nor UO_428 (O_428,N_24157,N_23948);
and UO_429 (O_429,N_22922,N_21924);
or UO_430 (O_430,N_22638,N_22134);
xnor UO_431 (O_431,N_20326,N_22804);
nand UO_432 (O_432,N_24851,N_20981);
nand UO_433 (O_433,N_22165,N_23032);
and UO_434 (O_434,N_21016,N_20129);
xnor UO_435 (O_435,N_22829,N_24765);
xor UO_436 (O_436,N_23458,N_22371);
nor UO_437 (O_437,N_20651,N_20888);
and UO_438 (O_438,N_20480,N_24495);
and UO_439 (O_439,N_20866,N_23755);
and UO_440 (O_440,N_20243,N_22217);
and UO_441 (O_441,N_21854,N_21729);
nand UO_442 (O_442,N_20882,N_21096);
or UO_443 (O_443,N_23505,N_21557);
nor UO_444 (O_444,N_22677,N_22147);
and UO_445 (O_445,N_24927,N_22985);
or UO_446 (O_446,N_24923,N_24314);
xor UO_447 (O_447,N_23662,N_22604);
and UO_448 (O_448,N_24552,N_20919);
and UO_449 (O_449,N_20304,N_22258);
nor UO_450 (O_450,N_23393,N_20948);
nand UO_451 (O_451,N_21636,N_21645);
nor UO_452 (O_452,N_22453,N_22910);
xnor UO_453 (O_453,N_23422,N_20314);
xnor UO_454 (O_454,N_21059,N_22111);
or UO_455 (O_455,N_23154,N_22715);
nand UO_456 (O_456,N_21828,N_24180);
or UO_457 (O_457,N_24639,N_20893);
and UO_458 (O_458,N_22827,N_22539);
or UO_459 (O_459,N_23144,N_20779);
xnor UO_460 (O_460,N_20634,N_23300);
xnor UO_461 (O_461,N_20738,N_22543);
nor UO_462 (O_462,N_24606,N_22381);
xnor UO_463 (O_463,N_22571,N_21441);
xnor UO_464 (O_464,N_22209,N_22245);
and UO_465 (O_465,N_23370,N_21184);
and UO_466 (O_466,N_24295,N_22890);
nor UO_467 (O_467,N_24227,N_20596);
nor UO_468 (O_468,N_23047,N_24229);
and UO_469 (O_469,N_22576,N_20327);
and UO_470 (O_470,N_21190,N_21240);
xnor UO_471 (O_471,N_23038,N_24812);
nor UO_472 (O_472,N_20628,N_20606);
nor UO_473 (O_473,N_23737,N_20952);
xnor UO_474 (O_474,N_23368,N_23865);
and UO_475 (O_475,N_23796,N_21971);
nand UO_476 (O_476,N_24474,N_22357);
nand UO_477 (O_477,N_23210,N_21536);
nand UO_478 (O_478,N_23476,N_22204);
or UO_479 (O_479,N_24042,N_24467);
or UO_480 (O_480,N_22343,N_21872);
and UO_481 (O_481,N_23099,N_23389);
nand UO_482 (O_482,N_24463,N_21151);
xnor UO_483 (O_483,N_24864,N_24572);
or UO_484 (O_484,N_23833,N_24494);
or UO_485 (O_485,N_22549,N_23775);
nor UO_486 (O_486,N_23314,N_20678);
and UO_487 (O_487,N_21480,N_20469);
nand UO_488 (O_488,N_24313,N_24776);
nor UO_489 (O_489,N_21051,N_22713);
or UO_490 (O_490,N_24664,N_21675);
nand UO_491 (O_491,N_20649,N_22814);
xor UO_492 (O_492,N_20984,N_21598);
and UO_493 (O_493,N_22212,N_20874);
or UO_494 (O_494,N_24078,N_23640);
or UO_495 (O_495,N_20443,N_20669);
nor UO_496 (O_496,N_21884,N_23220);
or UO_497 (O_497,N_20275,N_22744);
nor UO_498 (O_498,N_22177,N_20610);
nand UO_499 (O_499,N_23373,N_21337);
or UO_500 (O_500,N_21973,N_21604);
or UO_501 (O_501,N_23194,N_23148);
xor UO_502 (O_502,N_24280,N_20042);
xor UO_503 (O_503,N_20173,N_23684);
nor UO_504 (O_504,N_20444,N_22905);
or UO_505 (O_505,N_20014,N_23046);
or UO_506 (O_506,N_20107,N_21100);
nand UO_507 (O_507,N_24468,N_22613);
and UO_508 (O_508,N_21622,N_21495);
xnor UO_509 (O_509,N_22659,N_21095);
xor UO_510 (O_510,N_22229,N_24622);
nand UO_511 (O_511,N_21186,N_23621);
or UO_512 (O_512,N_21174,N_23358);
nand UO_513 (O_513,N_24591,N_22951);
or UO_514 (O_514,N_24836,N_22649);
or UO_515 (O_515,N_24333,N_20913);
or UO_516 (O_516,N_24547,N_21056);
or UO_517 (O_517,N_24151,N_24324);
nand UO_518 (O_518,N_23307,N_23023);
nor UO_519 (O_519,N_21940,N_23904);
and UO_520 (O_520,N_20357,N_20499);
xor UO_521 (O_521,N_23690,N_23872);
or UO_522 (O_522,N_20717,N_24411);
and UO_523 (O_523,N_23453,N_22950);
and UO_524 (O_524,N_21541,N_20746);
xor UO_525 (O_525,N_24076,N_22228);
or UO_526 (O_526,N_24753,N_24167);
and UO_527 (O_527,N_21564,N_21389);
nand UO_528 (O_528,N_20536,N_20413);
nand UO_529 (O_529,N_22664,N_22662);
or UO_530 (O_530,N_24045,N_22947);
and UO_531 (O_531,N_20358,N_24861);
nor UO_532 (O_532,N_24949,N_21120);
and UO_533 (O_533,N_21431,N_20804);
or UO_534 (O_534,N_20680,N_20901);
and UO_535 (O_535,N_22760,N_21723);
xnor UO_536 (O_536,N_24344,N_24397);
and UO_537 (O_537,N_24388,N_21080);
and UO_538 (O_538,N_20697,N_21231);
nand UO_539 (O_539,N_21701,N_22881);
or UO_540 (O_540,N_23739,N_20869);
xnor UO_541 (O_541,N_23448,N_20331);
xnor UO_542 (O_542,N_23408,N_20230);
nand UO_543 (O_543,N_23826,N_22235);
or UO_544 (O_544,N_20511,N_21330);
and UO_545 (O_545,N_21914,N_23158);
nand UO_546 (O_546,N_24970,N_20516);
nor UO_547 (O_547,N_21742,N_20238);
nor UO_548 (O_548,N_21554,N_21978);
nor UO_549 (O_549,N_24697,N_22889);
or UO_550 (O_550,N_20077,N_21690);
and UO_551 (O_551,N_21660,N_23984);
nor UO_552 (O_552,N_22159,N_23119);
and UO_553 (O_553,N_21089,N_21612);
nor UO_554 (O_554,N_24279,N_21437);
nor UO_555 (O_555,N_23284,N_24242);
nand UO_556 (O_556,N_24793,N_24260);
and UO_557 (O_557,N_22001,N_20512);
and UO_558 (O_558,N_20582,N_21053);
xor UO_559 (O_559,N_22757,N_22090);
and UO_560 (O_560,N_24979,N_23783);
xor UO_561 (O_561,N_20386,N_20186);
or UO_562 (O_562,N_21521,N_22775);
nand UO_563 (O_563,N_24206,N_21642);
or UO_564 (O_564,N_20393,N_21114);
xnor UO_565 (O_565,N_20497,N_20294);
or UO_566 (O_566,N_23238,N_22139);
or UO_567 (O_567,N_22156,N_21434);
nor UO_568 (O_568,N_20420,N_20632);
xor UO_569 (O_569,N_22658,N_20026);
xnor UO_570 (O_570,N_20899,N_20531);
nor UO_571 (O_571,N_20592,N_21156);
and UO_572 (O_572,N_20963,N_20319);
nand UO_573 (O_573,N_23926,N_24683);
nor UO_574 (O_574,N_23563,N_22273);
nor UO_575 (O_575,N_21073,N_24057);
nand UO_576 (O_576,N_22361,N_24798);
nand UO_577 (O_577,N_21581,N_22671);
nor UO_578 (O_578,N_24744,N_20320);
nor UO_579 (O_579,N_23766,N_23156);
nor UO_580 (O_580,N_20969,N_23496);
nor UO_581 (O_581,N_20783,N_21316);
nand UO_582 (O_582,N_23575,N_24385);
xnor UO_583 (O_583,N_20050,N_22699);
xor UO_584 (O_584,N_22711,N_21196);
or UO_585 (O_585,N_24805,N_23164);
and UO_586 (O_586,N_20086,N_22766);
nor UO_587 (O_587,N_21583,N_21268);
nor UO_588 (O_588,N_20270,N_21214);
and UO_589 (O_589,N_21979,N_21466);
nor UO_590 (O_590,N_22884,N_21220);
or UO_591 (O_591,N_22295,N_24361);
nor UO_592 (O_592,N_23362,N_21990);
and UO_593 (O_593,N_22537,N_23927);
nor UO_594 (O_594,N_22011,N_24904);
and UO_595 (O_595,N_22848,N_23477);
xnor UO_596 (O_596,N_24223,N_20760);
and UO_597 (O_597,N_22612,N_22878);
and UO_598 (O_598,N_22602,N_22226);
nor UO_599 (O_599,N_22841,N_23568);
nand UO_600 (O_600,N_20524,N_24880);
xnor UO_601 (O_601,N_23687,N_24721);
nand UO_602 (O_602,N_23382,N_20723);
nand UO_603 (O_603,N_20936,N_24738);
and UO_604 (O_604,N_20481,N_20347);
xor UO_605 (O_605,N_22174,N_24922);
xnor UO_606 (O_606,N_23919,N_21935);
and UO_607 (O_607,N_20965,N_23010);
or UO_608 (O_608,N_23983,N_24675);
or UO_609 (O_609,N_22203,N_23308);
nor UO_610 (O_610,N_20496,N_23981);
and UO_611 (O_611,N_24298,N_21585);
nor UO_612 (O_612,N_24908,N_20623);
and UO_613 (O_613,N_23609,N_23880);
and UO_614 (O_614,N_20595,N_22995);
nor UO_615 (O_615,N_21444,N_24077);
and UO_616 (O_616,N_21776,N_23956);
nor UO_617 (O_617,N_20289,N_20134);
nor UO_618 (O_618,N_23622,N_22849);
or UO_619 (O_619,N_22940,N_21249);
and UO_620 (O_620,N_22872,N_23348);
or UO_621 (O_621,N_24600,N_22459);
nand UO_622 (O_622,N_21013,N_22865);
and UO_623 (O_623,N_21607,N_23097);
nor UO_624 (O_624,N_22084,N_21208);
and UO_625 (O_625,N_21105,N_22173);
xor UO_626 (O_626,N_22276,N_23492);
xor UO_627 (O_627,N_22325,N_20145);
or UO_628 (O_628,N_20759,N_20532);
and UO_629 (O_629,N_20638,N_20599);
and UO_630 (O_630,N_22712,N_23392);
or UO_631 (O_631,N_24278,N_20183);
or UO_632 (O_632,N_24267,N_24250);
or UO_633 (O_633,N_23649,N_22386);
nand UO_634 (O_634,N_22434,N_23530);
or UO_635 (O_635,N_22967,N_22094);
or UO_636 (O_636,N_24788,N_24512);
and UO_637 (O_637,N_23957,N_22629);
nand UO_638 (O_638,N_23907,N_20339);
and UO_639 (O_639,N_21520,N_20647);
nor UO_640 (O_640,N_24399,N_20904);
nand UO_641 (O_641,N_20255,N_21235);
nor UO_642 (O_642,N_22394,N_20841);
nand UO_643 (O_643,N_22499,N_22452);
nor UO_644 (O_644,N_21191,N_22966);
nand UO_645 (O_645,N_20910,N_23840);
and UO_646 (O_646,N_22929,N_22765);
nand UO_647 (O_647,N_20476,N_23794);
nand UO_648 (O_648,N_23129,N_22803);
or UO_649 (O_649,N_20179,N_22312);
or UO_650 (O_650,N_23884,N_23419);
nor UO_651 (O_651,N_22986,N_22224);
nand UO_652 (O_652,N_24036,N_24019);
nor UO_653 (O_653,N_20729,N_21775);
nor UO_654 (O_654,N_24285,N_24130);
and UO_655 (O_655,N_23557,N_23306);
nor UO_656 (O_656,N_24729,N_20104);
nand UO_657 (O_657,N_22925,N_23169);
nand UO_658 (O_658,N_23106,N_22836);
xor UO_659 (O_659,N_22702,N_22557);
xnor UO_660 (O_660,N_20544,N_23689);
or UO_661 (O_661,N_22391,N_23003);
nand UO_662 (O_662,N_24643,N_24065);
xnor UO_663 (O_663,N_22474,N_22102);
nand UO_664 (O_664,N_24869,N_23704);
nor UO_665 (O_665,N_21377,N_20194);
xor UO_666 (O_666,N_24269,N_21705);
and UO_667 (O_667,N_21394,N_23385);
or UO_668 (O_668,N_21164,N_20854);
and UO_669 (O_669,N_20626,N_22318);
or UO_670 (O_670,N_24182,N_22593);
or UO_671 (O_671,N_23978,N_23791);
xor UO_672 (O_672,N_24653,N_23117);
or UO_673 (O_673,N_20335,N_23989);
and UO_674 (O_674,N_23245,N_22420);
or UO_675 (O_675,N_23386,N_22234);
nand UO_676 (O_676,N_23587,N_20269);
xor UO_677 (O_677,N_20288,N_23676);
xor UO_678 (O_678,N_23123,N_21802);
nand UO_679 (O_679,N_20642,N_23439);
xor UO_680 (O_680,N_23166,N_22787);
nand UO_681 (O_681,N_22454,N_20209);
or UO_682 (O_682,N_24258,N_20787);
or UO_683 (O_683,N_22373,N_23658);
or UO_684 (O_684,N_24123,N_22074);
xnor UO_685 (O_685,N_24508,N_21529);
or UO_686 (O_686,N_21439,N_22070);
nor UO_687 (O_687,N_20491,N_22068);
xnor UO_688 (O_688,N_24677,N_22137);
nor UO_689 (O_689,N_24976,N_21093);
nand UO_690 (O_690,N_23214,N_24255);
xnor UO_691 (O_691,N_20221,N_21548);
nand UO_692 (O_692,N_21628,N_23524);
nand UO_693 (O_693,N_21373,N_23825);
nor UO_694 (O_694,N_20724,N_21951);
or UO_695 (O_695,N_22329,N_24682);
nand UO_696 (O_696,N_24034,N_24689);
nand UO_697 (O_697,N_24972,N_24562);
nand UO_698 (O_698,N_20242,N_21750);
nand UO_699 (O_699,N_24249,N_23643);
nand UO_700 (O_700,N_23641,N_23578);
and UO_701 (O_701,N_20887,N_22128);
and UO_702 (O_702,N_24504,N_22476);
and UO_703 (O_703,N_20802,N_24412);
and UO_704 (O_704,N_20559,N_23490);
xnor UO_705 (O_705,N_22051,N_20060);
or UO_706 (O_706,N_20494,N_22695);
and UO_707 (O_707,N_20791,N_21355);
nand UO_708 (O_708,N_22897,N_21880);
xnor UO_709 (O_709,N_21887,N_23661);
xor UO_710 (O_710,N_24874,N_21387);
nand UO_711 (O_711,N_24009,N_20684);
or UO_712 (O_712,N_20052,N_22470);
or UO_713 (O_713,N_21351,N_24535);
nand UO_714 (O_714,N_22734,N_24106);
xnor UO_715 (O_715,N_23018,N_20165);
xnor UO_716 (O_716,N_24671,N_21771);
nor UO_717 (O_717,N_23033,N_21910);
nor UO_718 (O_718,N_20362,N_21849);
nand UO_719 (O_719,N_22843,N_24457);
and UO_720 (O_720,N_24526,N_24944);
xnor UO_721 (O_721,N_24453,N_20916);
and UO_722 (O_722,N_21883,N_24364);
and UO_723 (O_723,N_22968,N_20278);
nor UO_724 (O_724,N_23484,N_21682);
xor UO_725 (O_725,N_23900,N_20425);
and UO_726 (O_726,N_21540,N_23725);
xor UO_727 (O_727,N_22444,N_21960);
xor UO_728 (O_728,N_21625,N_20636);
or UO_729 (O_729,N_21428,N_20007);
xor UO_730 (O_730,N_22081,N_23633);
xnor UO_731 (O_731,N_20674,N_22624);
xor UO_732 (O_732,N_22900,N_23135);
or UO_733 (O_733,N_23224,N_23665);
nor UO_734 (O_734,N_20352,N_21823);
nor UO_735 (O_735,N_22169,N_22508);
and UO_736 (O_736,N_24802,N_22223);
nor UO_737 (O_737,N_21415,N_21907);
nor UO_738 (O_738,N_24565,N_24135);
xor UO_739 (O_739,N_23168,N_20488);
and UO_740 (O_740,N_24465,N_22587);
or UO_741 (O_741,N_22298,N_24475);
or UO_742 (O_742,N_21139,N_20142);
nand UO_743 (O_743,N_24681,N_21281);
xnor UO_744 (O_744,N_23591,N_20317);
nor UO_745 (O_745,N_23409,N_21609);
nand UO_746 (O_746,N_20338,N_23730);
xnor UO_747 (O_747,N_22953,N_22777);
nor UO_748 (O_748,N_20835,N_20608);
xor UO_749 (O_749,N_21533,N_23582);
nor UO_750 (O_750,N_21522,N_22520);
nand UO_751 (O_751,N_21916,N_24201);
nand UO_752 (O_752,N_24998,N_22225);
xnor UO_753 (O_753,N_23994,N_22954);
or UO_754 (O_754,N_20303,N_22580);
and UO_755 (O_755,N_21656,N_21905);
or UO_756 (O_756,N_23845,N_21825);
or UO_757 (O_757,N_22351,N_21696);
nand UO_758 (O_758,N_24374,N_24001);
and UO_759 (O_759,N_21651,N_20526);
xor UO_760 (O_760,N_21157,N_20988);
xnor UO_761 (O_761,N_20589,N_20406);
nand UO_762 (O_762,N_24767,N_21968);
and UO_763 (O_763,N_21580,N_22984);
or UO_764 (O_764,N_24821,N_22661);
nor UO_765 (O_765,N_22955,N_22790);
and UO_766 (O_766,N_24194,N_20518);
nand UO_767 (O_767,N_23828,N_22475);
nor UO_768 (O_768,N_22086,N_20842);
and UO_769 (O_769,N_24110,N_22277);
and UO_770 (O_770,N_22080,N_23290);
nand UO_771 (O_771,N_22635,N_21282);
nor UO_772 (O_772,N_24530,N_22614);
or UO_773 (O_773,N_21484,N_23356);
xor UO_774 (O_774,N_21998,N_23929);
or UO_775 (O_775,N_23651,N_20409);
nand UO_776 (O_776,N_21260,N_22417);
nor UO_777 (O_777,N_22585,N_23427);
nand UO_778 (O_778,N_21245,N_22875);
nor UO_779 (O_779,N_22736,N_21225);
or UO_780 (O_780,N_22492,N_24093);
nand UO_781 (O_781,N_22903,N_24174);
xor UO_782 (O_782,N_24846,N_21407);
nand UO_783 (O_783,N_20561,N_24900);
nor UO_784 (O_784,N_21614,N_21899);
nor UO_785 (O_785,N_22254,N_21647);
or UO_786 (O_786,N_23962,N_20140);
or UO_787 (O_787,N_23377,N_24035);
and UO_788 (O_788,N_20773,N_23287);
xnor UO_789 (O_789,N_21857,N_21840);
or UO_790 (O_790,N_24127,N_24124);
or UO_791 (O_791,N_24085,N_23024);
xor UO_792 (O_792,N_21418,N_20231);
nor UO_793 (O_793,N_24740,N_21816);
or UO_794 (O_794,N_21386,N_22164);
nor UO_795 (O_795,N_22141,N_20844);
xor UO_796 (O_796,N_23754,N_24073);
nor UO_797 (O_797,N_24363,N_23100);
and UO_798 (O_798,N_21432,N_21098);
nor UO_799 (O_799,N_24254,N_21794);
and UO_800 (O_800,N_22449,N_23225);
and UO_801 (O_801,N_22240,N_22368);
nand UO_802 (O_802,N_24718,N_24370);
nand UO_803 (O_803,N_20290,N_23998);
or UO_804 (O_804,N_21819,N_21213);
and UO_805 (O_805,N_23172,N_20639);
nor UO_806 (O_806,N_21949,N_21975);
nor UO_807 (O_807,N_22033,N_24329);
nor UO_808 (O_808,N_22413,N_21170);
nor UO_809 (O_809,N_20285,N_24277);
and UO_810 (O_810,N_23674,N_24178);
and UO_811 (O_811,N_22560,N_20928);
nor UO_812 (O_812,N_24583,N_21826);
nor UO_813 (O_813,N_24287,N_20220);
nor UO_814 (O_814,N_20445,N_21537);
or UO_815 (O_815,N_22842,N_21491);
nor UO_816 (O_816,N_20987,N_20301);
nor UO_817 (O_817,N_24375,N_22619);
nor UO_818 (O_818,N_21634,N_21001);
nand UO_819 (O_819,N_20721,N_24756);
nor UO_820 (O_820,N_23724,N_23672);
and UO_821 (O_821,N_23482,N_23554);
and UO_822 (O_822,N_24875,N_22121);
nand UO_823 (O_823,N_20293,N_22683);
nor UO_824 (O_824,N_23437,N_20695);
nand UO_825 (O_825,N_23057,N_20281);
and UO_826 (O_826,N_23075,N_21390);
xnor UO_827 (O_827,N_23433,N_20924);
nand UO_828 (O_828,N_23635,N_24799);
and UO_829 (O_829,N_20163,N_20788);
and UO_830 (O_830,N_24236,N_24480);
or UO_831 (O_831,N_20851,N_24773);
xor UO_832 (O_832,N_21391,N_23750);
and UO_833 (O_833,N_20560,N_22979);
xnor UO_834 (O_834,N_24118,N_22541);
or UO_835 (O_835,N_21516,N_22489);
xnor UO_836 (O_836,N_23388,N_21344);
and UO_837 (O_837,N_23832,N_23733);
nand UO_838 (O_838,N_21076,N_24038);
xor UO_839 (O_839,N_21364,N_24894);
nor UO_840 (O_840,N_21429,N_22832);
xnor UO_841 (O_841,N_21577,N_20401);
nand UO_842 (O_842,N_22406,N_23528);
or UO_843 (O_843,N_20095,N_21123);
and UO_844 (O_844,N_20977,N_24541);
or UO_845 (O_845,N_21831,N_22293);
nand UO_846 (O_846,N_24745,N_24149);
or UO_847 (O_847,N_22687,N_24492);
and UO_848 (O_848,N_22564,N_22100);
xnor UO_849 (O_849,N_23912,N_22663);
xnor UO_850 (O_850,N_24028,N_24056);
and UO_851 (O_851,N_24104,N_23208);
or UO_852 (O_852,N_22845,N_24568);
nor UO_853 (O_853,N_23636,N_22989);
or UO_854 (O_854,N_24461,N_23547);
nand UO_855 (O_855,N_24282,N_24945);
nor UO_856 (O_856,N_21463,N_23758);
xnor UO_857 (O_857,N_20800,N_22113);
xnor UO_858 (O_858,N_23229,N_22024);
xor UO_859 (O_859,N_23916,N_23711);
and UO_860 (O_860,N_20761,N_24580);
and UO_861 (O_861,N_21210,N_24185);
or UO_862 (O_862,N_21423,N_22935);
xor UO_863 (O_863,N_23542,N_21844);
and UO_864 (O_864,N_24321,N_21925);
nand UO_865 (O_865,N_22676,N_21159);
nor UO_866 (O_866,N_22756,N_22384);
xnor UO_867 (O_867,N_22741,N_23244);
nand UO_868 (O_868,N_23874,N_21461);
nand UO_869 (O_869,N_21983,N_20794);
xnor UO_870 (O_870,N_22270,N_21223);
or UO_871 (O_871,N_22908,N_22725);
nor UO_872 (O_872,N_24699,N_21113);
nor UO_873 (O_873,N_24083,N_21375);
and UO_874 (O_874,N_23527,N_22527);
nor UO_875 (O_875,N_23941,N_22200);
xor UO_876 (O_876,N_23436,N_24822);
or UO_877 (O_877,N_23922,N_22644);
or UO_878 (O_878,N_23958,N_21079);
nor UO_879 (O_879,N_21405,N_21867);
xnor UO_880 (O_880,N_23867,N_22202);
or UO_881 (O_881,N_23004,N_20975);
xor UO_882 (O_882,N_21395,N_21791);
or UO_883 (O_883,N_22383,N_24534);
xnor UO_884 (O_884,N_21821,N_24003);
nand UO_885 (O_885,N_21809,N_23416);
xor UO_886 (O_886,N_23604,N_20198);
xnor UO_887 (O_887,N_21269,N_22180);
nand UO_888 (O_888,N_24177,N_21161);
nor UO_889 (O_889,N_23700,N_20941);
nor UO_890 (O_890,N_24731,N_23103);
and UO_891 (O_891,N_21296,N_23049);
nor UO_892 (O_892,N_22198,N_20258);
and UO_893 (O_893,N_20935,N_22688);
and UO_894 (O_894,N_23536,N_24933);
or UO_895 (O_895,N_22647,N_23237);
xnor UO_896 (O_896,N_20945,N_21740);
and UO_897 (O_897,N_22697,N_24749);
nand UO_898 (O_898,N_21086,N_23176);
and UO_899 (O_899,N_20147,N_20943);
nor UO_900 (O_900,N_22703,N_20360);
nor UO_901 (O_901,N_23764,N_24111);
nand UO_902 (O_902,N_20679,N_23255);
xor UO_903 (O_903,N_24570,N_23611);
and UO_904 (O_904,N_24578,N_23021);
nor UO_905 (O_905,N_20477,N_23346);
nand UO_906 (O_906,N_20363,N_22083);
nor UO_907 (O_907,N_20124,N_22439);
and UO_908 (O_908,N_22962,N_20677);
nor UO_909 (O_909,N_21894,N_23535);
xor UO_910 (O_910,N_21845,N_20955);
and UO_911 (O_911,N_22047,N_24665);
nand UO_912 (O_912,N_20487,N_23471);
xor UO_913 (O_913,N_20522,N_22691);
nand UO_914 (O_914,N_24121,N_23657);
nor UO_915 (O_915,N_22681,N_24010);
or UO_916 (O_916,N_23337,N_20062);
nor UO_917 (O_917,N_23446,N_22555);
and UO_918 (O_918,N_21524,N_20564);
nor UO_919 (O_919,N_22904,N_24283);
and UO_920 (O_920,N_21568,N_22776);
nand UO_921 (O_921,N_20164,N_22389);
nor UO_922 (O_922,N_22901,N_20066);
or UO_923 (O_923,N_22869,N_21739);
and UO_924 (O_924,N_20546,N_24473);
or UO_925 (O_925,N_20315,N_22551);
xor UO_926 (O_926,N_24355,N_20308);
xnor UO_927 (O_927,N_24963,N_23526);
or UO_928 (O_928,N_24241,N_21865);
nand UO_929 (O_929,N_20199,N_22794);
xnor UO_930 (O_930,N_23495,N_21818);
nor UO_931 (O_931,N_23183,N_22161);
nor UO_932 (O_932,N_22106,N_21805);
or UO_933 (O_933,N_24302,N_23340);
and UO_934 (O_934,N_23533,N_20620);
xnor UO_935 (O_935,N_23413,N_24603);
xor UO_936 (O_936,N_23136,N_21668);
and UO_937 (O_937,N_20426,N_23812);
xnor UO_938 (O_938,N_22566,N_21343);
nor UO_939 (O_939,N_22238,N_24112);
and UO_940 (O_940,N_22882,N_23811);
nor UO_941 (O_941,N_21654,N_24507);
nand UO_942 (O_942,N_21328,N_21691);
nand UO_943 (O_943,N_22597,N_23653);
xor UO_944 (O_944,N_21401,N_23838);
and UO_945 (O_945,N_23366,N_21545);
nand UO_946 (O_946,N_22388,N_22353);
and UO_947 (O_947,N_21822,N_22031);
and UO_948 (O_948,N_23899,N_20440);
or UO_949 (O_949,N_20873,N_21265);
or UO_950 (O_950,N_21414,N_22617);
or UO_951 (O_951,N_24566,N_23620);
nor UO_952 (O_952,N_21574,N_24730);
nor UO_953 (O_953,N_22888,N_24717);
nand UO_954 (O_954,N_22409,N_22321);
nor UO_955 (O_955,N_23800,N_21518);
nand UO_956 (O_956,N_24506,N_22674);
nor UO_957 (O_957,N_21772,N_20627);
and UO_958 (O_958,N_21915,N_23181);
nor UO_959 (O_959,N_22589,N_20820);
and UO_960 (O_960,N_23084,N_23060);
and UO_961 (O_961,N_23953,N_24247);
xor UO_962 (O_962,N_21462,N_22511);
or UO_963 (O_963,N_24501,N_21436);
nor UO_964 (O_964,N_23445,N_21176);
and UO_965 (O_965,N_23428,N_23231);
and UO_966 (O_966,N_21046,N_20616);
nor UO_967 (O_967,N_24339,N_20123);
or UO_968 (O_968,N_21523,N_23209);
nand UO_969 (O_969,N_21374,N_20550);
nand UO_970 (O_970,N_20954,N_22588);
or UO_971 (O_971,N_21035,N_20382);
xor UO_972 (O_972,N_22941,N_21257);
or UO_973 (O_973,N_24707,N_21255);
and UO_974 (O_974,N_23571,N_24511);
xor UO_975 (O_975,N_23150,N_20744);
or UO_976 (O_976,N_20644,N_23805);
and UO_977 (O_977,N_23043,N_23459);
and UO_978 (O_978,N_23520,N_22921);
nor UO_979 (O_979,N_23036,N_22591);
nand UO_980 (O_980,N_20417,N_20380);
xnor UO_981 (O_981,N_22779,N_24997);
or UO_982 (O_982,N_20398,N_24914);
nand UO_983 (O_983,N_24803,N_22981);
or UO_984 (O_984,N_22358,N_20359);
nand UO_985 (O_985,N_23424,N_23015);
nor UO_986 (O_986,N_20442,N_23932);
or UO_987 (O_987,N_23722,N_23877);
nor UO_988 (O_988,N_22855,N_24597);
nand UO_989 (O_989,N_20284,N_20892);
and UO_990 (O_990,N_22208,N_22352);
or UO_991 (O_991,N_24712,N_23572);
nand UO_992 (O_992,N_24896,N_23815);
nand UO_993 (O_993,N_21295,N_20903);
nand UO_994 (O_994,N_23849,N_20266);
nand UO_995 (O_995,N_23381,N_21736);
nand UO_996 (O_996,N_20031,N_24834);
and UO_997 (O_997,N_24347,N_23947);
or UO_998 (O_998,N_20933,N_20994);
nor UO_999 (O_999,N_23153,N_20091);
nor UO_1000 (O_1000,N_22518,N_24921);
nand UO_1001 (O_1001,N_21963,N_20464);
and UO_1002 (O_1002,N_24903,N_24806);
nand UO_1003 (O_1003,N_23971,N_20022);
and UO_1004 (O_1004,N_22643,N_22839);
and UO_1005 (O_1005,N_20106,N_23918);
nand UO_1006 (O_1006,N_23548,N_24434);
nor UO_1007 (O_1007,N_24895,N_22945);
and UO_1008 (O_1008,N_22288,N_22920);
and UO_1009 (O_1009,N_21735,N_23638);
nor UO_1010 (O_1010,N_20971,N_20657);
xor UO_1011 (O_1011,N_20537,N_20412);
or UO_1012 (O_1012,N_20251,N_23844);
nand UO_1013 (O_1013,N_21048,N_21122);
nor UO_1014 (O_1014,N_23506,N_20478);
xnor UO_1015 (O_1015,N_20461,N_23646);
or UO_1016 (O_1016,N_23336,N_22438);
xnor UO_1017 (O_1017,N_20785,N_21835);
nor UO_1018 (O_1018,N_20370,N_21710);
nand UO_1019 (O_1019,N_21130,N_24133);
and UO_1020 (O_1020,N_21458,N_21694);
nand UO_1021 (O_1021,N_22861,N_21559);
and UO_1022 (O_1022,N_23248,N_22800);
and UO_1023 (O_1023,N_21594,N_24954);
or UO_1024 (O_1024,N_22694,N_24380);
nor UO_1025 (O_1025,N_21109,N_22665);
nor UO_1026 (O_1026,N_20436,N_24191);
xnor UO_1027 (O_1027,N_20776,N_23195);
and UO_1028 (O_1028,N_21007,N_20144);
nor UO_1029 (O_1029,N_20137,N_22574);
nand UO_1030 (O_1030,N_23048,N_21148);
nand UO_1031 (O_1031,N_24371,N_21455);
xor UO_1032 (O_1032,N_20211,N_22021);
nand UO_1033 (O_1033,N_22746,N_22310);
nand UO_1034 (O_1034,N_21600,N_22319);
xor UO_1035 (O_1035,N_22041,N_23782);
or UO_1036 (O_1036,N_20960,N_20543);
nor UO_1037 (O_1037,N_22306,N_22076);
nor UO_1038 (O_1038,N_22085,N_24061);
xnor UO_1039 (O_1039,N_24557,N_23655);
xnor UO_1040 (O_1040,N_23781,N_23242);
nor UO_1041 (O_1041,N_23326,N_20774);
or UO_1042 (O_1042,N_23940,N_24710);
or UO_1043 (O_1043,N_20907,N_24584);
nor UO_1044 (O_1044,N_21504,N_20506);
nand UO_1045 (O_1045,N_23964,N_21041);
nand UO_1046 (O_1046,N_23911,N_21027);
nand UO_1047 (O_1047,N_22191,N_20828);
nor UO_1048 (O_1048,N_20161,N_24832);
nor UO_1049 (O_1049,N_23365,N_20138);
and UO_1050 (O_1050,N_21502,N_22073);
and UO_1051 (O_1051,N_24008,N_22356);
nor UO_1052 (O_1052,N_24993,N_21737);
nand UO_1053 (O_1053,N_20940,N_22435);
or UO_1054 (O_1054,N_21212,N_21261);
nor UO_1055 (O_1055,N_23588,N_23125);
and UO_1056 (O_1056,N_22886,N_20126);
or UO_1057 (O_1057,N_21465,N_22581);
and UO_1058 (O_1058,N_22871,N_23529);
nor UO_1059 (O_1059,N_20345,N_23830);
and UO_1060 (O_1060,N_22926,N_24481);
xor UO_1061 (O_1061,N_22758,N_23400);
nor UO_1062 (O_1062,N_24335,N_24625);
nor UO_1063 (O_1063,N_23543,N_22490);
nor UO_1064 (O_1064,N_23335,N_21149);
nor UO_1065 (O_1065,N_21875,N_21314);
xor UO_1066 (O_1066,N_23831,N_23985);
or UO_1067 (O_1067,N_22846,N_21785);
xor UO_1068 (O_1068,N_23017,N_22326);
or UO_1069 (O_1069,N_22050,N_24833);
nand UO_1070 (O_1070,N_21896,N_23037);
and UO_1071 (O_1071,N_20547,N_21006);
xor UO_1072 (O_1072,N_21596,N_21464);
xor UO_1073 (O_1073,N_22346,N_23406);
xor UO_1074 (O_1074,N_21021,N_21070);
and UO_1075 (O_1075,N_23853,N_24416);
or UO_1076 (O_1076,N_21538,N_22054);
or UO_1077 (O_1077,N_23675,N_22187);
nand UO_1078 (O_1078,N_21649,N_21570);
xor UO_1079 (O_1079,N_20176,N_21226);
or UO_1080 (O_1080,N_20313,N_24070);
and UO_1081 (O_1081,N_22639,N_23560);
nor UO_1082 (O_1082,N_21417,N_22837);
xnor UO_1083 (O_1083,N_23776,N_22625);
or UO_1084 (O_1084,N_20886,N_22257);
xnor UO_1085 (O_1085,N_24974,N_21698);
xor UO_1086 (O_1086,N_22419,N_21081);
or UO_1087 (O_1087,N_24030,N_21920);
and UO_1088 (O_1088,N_20208,N_21063);
nand UO_1089 (O_1089,N_21783,N_22314);
or UO_1090 (O_1090,N_21147,N_22640);
or UO_1091 (O_1091,N_23139,N_23039);
or UO_1092 (O_1092,N_24369,N_24691);
nand UO_1093 (O_1093,N_23507,N_21758);
nand UO_1094 (O_1094,N_20459,N_22971);
xnor UO_1095 (O_1095,N_24011,N_22028);
and UO_1096 (O_1096,N_22813,N_23576);
nor UO_1097 (O_1097,N_23669,N_21681);
nor UO_1098 (O_1098,N_22190,N_23652);
and UO_1099 (O_1099,N_21376,N_24661);
nand UO_1100 (O_1100,N_23025,N_24725);
xor UO_1101 (O_1101,N_21090,N_24796);
or UO_1102 (O_1102,N_24337,N_21689);
or UO_1103 (O_1103,N_22799,N_21549);
nand UO_1104 (O_1104,N_22151,N_24636);
and UO_1105 (O_1105,N_21534,N_20180);
and UO_1106 (O_1106,N_21019,N_20951);
nand UO_1107 (O_1107,N_22268,N_20085);
nand UO_1108 (O_1108,N_23969,N_24487);
nand UO_1109 (O_1109,N_24384,N_24141);
nand UO_1110 (O_1110,N_20973,N_22034);
and UO_1111 (O_1111,N_24449,N_24154);
nand UO_1112 (O_1112,N_20500,N_20112);
nand UO_1113 (O_1113,N_23264,N_24847);
and UO_1114 (O_1114,N_23807,N_23185);
and UO_1115 (O_1115,N_24850,N_21838);
xor UO_1116 (O_1116,N_22087,N_21877);
and UO_1117 (O_1117,N_21309,N_21321);
nand UO_1118 (O_1118,N_22652,N_20900);
xor UO_1119 (O_1119,N_20246,N_24628);
xor UO_1120 (O_1120,N_23321,N_22912);
or UO_1121 (O_1121,N_22565,N_20084);
nor UO_1122 (O_1122,N_20646,N_24811);
or UO_1123 (O_1123,N_24240,N_24026);
or UO_1124 (O_1124,N_20661,N_24726);
nor UO_1125 (O_1125,N_21034,N_20902);
nand UO_1126 (O_1126,N_22729,N_20870);
nand UO_1127 (O_1127,N_22376,N_24907);
or UO_1128 (O_1128,N_22675,N_23772);
or UO_1129 (O_1129,N_22398,N_21251);
and UO_1130 (O_1130,N_23875,N_22783);
nor UO_1131 (O_1131,N_23866,N_20855);
xnor UO_1132 (O_1132,N_22479,N_21115);
nand UO_1133 (O_1133,N_23618,N_24521);
and UO_1134 (O_1134,N_22471,N_24662);
or UO_1135 (O_1135,N_21565,N_20576);
or UO_1136 (O_1136,N_20594,N_24211);
xnor UO_1137 (O_1137,N_20203,N_20613);
and UO_1138 (O_1138,N_22215,N_23076);
nor UO_1139 (O_1139,N_24873,N_21350);
xnor UO_1140 (O_1140,N_22880,N_21361);
and UO_1141 (O_1141,N_21517,N_24648);
nand UO_1142 (O_1142,N_24524,N_23412);
nor UO_1143 (O_1143,N_20098,N_21886);
and UO_1144 (O_1144,N_20340,N_23190);
xnor UO_1145 (O_1145,N_23574,N_24598);
nand UO_1146 (O_1146,N_24402,N_22280);
nand UO_1147 (O_1147,N_23512,N_22509);
and UO_1148 (O_1148,N_24017,N_20263);
xor UO_1149 (O_1149,N_23011,N_22303);
xnor UO_1150 (O_1150,N_24739,N_21652);
and UO_1151 (O_1151,N_20768,N_24356);
xor UO_1152 (O_1152,N_23485,N_24747);
nand UO_1153 (O_1153,N_22411,N_21769);
or UO_1154 (O_1154,N_20316,N_20116);
nor UO_1155 (O_1155,N_21362,N_24582);
and UO_1156 (O_1156,N_22503,N_23058);
xor UO_1157 (O_1157,N_24971,N_22281);
or UO_1158 (O_1158,N_22762,N_20653);
xnor UO_1159 (O_1159,N_22899,N_23350);
or UO_1160 (O_1160,N_21155,N_24391);
nand UO_1161 (O_1161,N_22065,N_21118);
nand UO_1162 (O_1162,N_20722,N_24669);
or UO_1163 (O_1163,N_23990,N_20394);
nand UO_1164 (O_1164,N_22162,N_20329);
xnor UO_1165 (O_1165,N_22755,N_22466);
or UO_1166 (O_1166,N_20071,N_22465);
nand UO_1167 (O_1167,N_22014,N_20730);
xor UO_1168 (O_1168,N_23466,N_23613);
xnor UO_1169 (O_1169,N_23411,N_20986);
xnor UO_1170 (O_1170,N_24623,N_22487);
or UO_1171 (O_1171,N_21800,N_21994);
nor UO_1172 (O_1172,N_21677,N_20001);
nor UO_1173 (O_1173,N_20034,N_21116);
nor UO_1174 (O_1174,N_22363,N_20297);
xor UO_1175 (O_1175,N_24173,N_21578);
nand UO_1176 (O_1176,N_23721,N_20737);
nor UO_1177 (O_1177,N_24054,N_21023);
or UO_1178 (O_1178,N_23606,N_24937);
or UO_1179 (O_1179,N_24735,N_24325);
xor UO_1180 (O_1180,N_24757,N_22553);
xnor UO_1181 (O_1181,N_24529,N_20139);
xor UO_1182 (O_1182,N_23170,N_24737);
and UO_1183 (O_1183,N_24116,N_24276);
xor UO_1184 (O_1184,N_23421,N_20968);
nand UO_1185 (O_1185,N_20740,N_20452);
or UO_1186 (O_1186,N_23303,N_23222);
nand UO_1187 (O_1187,N_22255,N_21000);
xnor UO_1188 (O_1188,N_22286,N_20972);
and UO_1189 (O_1189,N_23212,N_20244);
and UO_1190 (O_1190,N_21106,N_20397);
xnor UO_1191 (O_1191,N_24646,N_20259);
nand UO_1192 (O_1192,N_21338,N_21817);
and UO_1193 (O_1193,N_23789,N_24551);
nor UO_1194 (O_1194,N_23707,N_21301);
xnor UO_1195 (O_1195,N_24230,N_22994);
and UO_1196 (O_1196,N_20731,N_21964);
or UO_1197 (O_1197,N_20846,N_24751);
nor UO_1198 (O_1198,N_21306,N_24666);
nor UO_1199 (O_1199,N_20287,N_20711);
nor UO_1200 (O_1200,N_23608,N_21850);
nor UO_1201 (O_1201,N_20716,N_21175);
nand UO_1202 (O_1202,N_20367,N_22440);
nand UO_1203 (O_1203,N_24838,N_21603);
and UO_1204 (O_1204,N_22308,N_21669);
and UO_1205 (O_1205,N_23127,N_21552);
xnor UO_1206 (O_1206,N_23235,N_23878);
xnor UO_1207 (O_1207,N_20087,N_20282);
or UO_1208 (O_1208,N_21644,N_23935);
nand UO_1209 (O_1209,N_23005,N_22302);
nand UO_1210 (O_1210,N_20814,N_22016);
xor UO_1211 (O_1211,N_21010,N_20334);
xnor UO_1212 (O_1212,N_21496,N_24814);
nand UO_1213 (O_1213,N_21941,N_21550);
or UO_1214 (O_1214,N_20097,N_20867);
nor UO_1215 (O_1215,N_24496,N_22347);
nor UO_1216 (O_1216,N_21413,N_21655);
nor UO_1217 (O_1217,N_24532,N_21124);
xor UO_1218 (O_1218,N_23343,N_23494);
nor UO_1219 (O_1219,N_23083,N_24992);
and UO_1220 (O_1220,N_21999,N_21258);
xnor UO_1221 (O_1221,N_23822,N_22510);
or UO_1222 (O_1222,N_22253,N_21133);
nand UO_1223 (O_1223,N_22350,N_20188);
and UO_1224 (O_1224,N_21453,N_23434);
xnor UO_1225 (O_1225,N_21018,N_22027);
or UO_1226 (O_1226,N_24858,N_22529);
nand UO_1227 (O_1227,N_20523,N_23650);
or UO_1228 (O_1228,N_21452,N_21711);
or UO_1229 (O_1229,N_20343,N_22481);
and UO_1230 (O_1230,N_20878,N_22408);
nand UO_1231 (O_1231,N_22797,N_21074);
and UO_1232 (O_1232,N_20133,N_24484);
xor UO_1233 (O_1233,N_22359,N_22696);
or UO_1234 (O_1234,N_21847,N_23161);
nand UO_1235 (O_1235,N_20563,N_24145);
nand UO_1236 (O_1236,N_20880,N_21832);
nand UO_1237 (O_1237,N_24548,N_22500);
or UO_1238 (O_1238,N_23311,N_22422);
and UO_1239 (O_1239,N_23925,N_23175);
nor UO_1240 (O_1240,N_20660,N_24994);
xnor UO_1241 (O_1241,N_22249,N_24443);
xnor UO_1242 (O_1242,N_24147,N_24693);
nand UO_1243 (O_1243,N_21948,N_20305);
xnor UO_1244 (O_1244,N_20696,N_22124);
nor UO_1245 (O_1245,N_21637,N_22247);
xnor UO_1246 (O_1246,N_23040,N_21989);
and UO_1247 (O_1247,N_21861,N_20408);
and UO_1248 (O_1248,N_21037,N_24452);
nand UO_1249 (O_1249,N_23594,N_21908);
nor UO_1250 (O_1250,N_20548,N_24390);
xor UO_1251 (O_1251,N_20748,N_23488);
or UO_1252 (O_1252,N_22472,N_24163);
and UO_1253 (O_1253,N_23734,N_20296);
and UO_1254 (O_1254,N_22558,N_24244);
xnor UO_1255 (O_1255,N_20743,N_23999);
and UO_1256 (O_1256,N_22893,N_23254);
nand UO_1257 (O_1257,N_21627,N_23199);
xnor UO_1258 (O_1258,N_22140,N_23612);
or UO_1259 (O_1259,N_24792,N_21945);
and UO_1260 (O_1260,N_21893,N_23133);
or UO_1261 (O_1261,N_24807,N_23204);
or UO_1262 (O_1262,N_20336,N_20463);
nand UO_1263 (O_1263,N_23327,N_20699);
and UO_1264 (O_1264,N_22425,N_20551);
nor UO_1265 (O_1265,N_21528,N_21573);
nand UO_1266 (O_1266,N_22885,N_22497);
nand UO_1267 (O_1267,N_23355,N_21511);
nor UO_1268 (O_1268,N_21824,N_20762);
xnor UO_1269 (O_1269,N_24698,N_22136);
nor UO_1270 (O_1270,N_21680,N_21315);
nand UO_1271 (O_1271,N_24372,N_21846);
nand UO_1272 (O_1272,N_20200,N_22327);
xnor UO_1273 (O_1273,N_24866,N_24522);
nor UO_1274 (O_1274,N_24055,N_23200);
xnor UO_1275 (O_1275,N_22874,N_22231);
and UO_1276 (O_1276,N_23774,N_21162);
xor UO_1277 (O_1277,N_20603,N_23562);
xnor UO_1278 (O_1278,N_20023,N_20691);
and UO_1279 (O_1279,N_21194,N_23080);
or UO_1280 (O_1280,N_24006,N_24210);
nand UO_1281 (O_1281,N_21708,N_24784);
or UO_1282 (O_1282,N_23415,N_23503);
xor UO_1283 (O_1283,N_21617,N_24479);
or UO_1284 (O_1284,N_21810,N_23770);
nor UO_1285 (O_1285,N_22263,N_24062);
xnor UO_1286 (O_1286,N_23187,N_23938);
nor UO_1287 (O_1287,N_24340,N_22022);
nand UO_1288 (O_1288,N_24426,N_24831);
nand UO_1289 (O_1289,N_21279,N_20069);
or UO_1290 (O_1290,N_24268,N_23101);
and UO_1291 (O_1291,N_24216,N_24879);
xnor UO_1292 (O_1292,N_22970,N_22847);
or UO_1293 (O_1293,N_20311,N_22401);
and UO_1294 (O_1294,N_22656,N_20122);
xor UO_1295 (O_1295,N_24429,N_20036);
xor UO_1296 (O_1296,N_23677,N_20387);
and UO_1297 (O_1297,N_24585,N_24162);
nand UO_1298 (O_1298,N_20726,N_23615);
nand UO_1299 (O_1299,N_24742,N_21143);
xor UO_1300 (O_1300,N_24464,N_20755);
xnor UO_1301 (O_1301,N_20961,N_22456);
or UO_1302 (O_1302,N_21248,N_21237);
nor UO_1303 (O_1303,N_22093,N_24826);
nand UO_1304 (O_1304,N_21065,N_24604);
nand UO_1305 (O_1305,N_23793,N_23995);
or UO_1306 (O_1306,N_23680,N_21202);
or UO_1307 (O_1307,N_20368,N_21974);
nand UO_1308 (O_1308,N_20845,N_20240);
and UO_1309 (O_1309,N_21188,N_22505);
xor UO_1310 (O_1310,N_24129,N_22339);
nand UO_1311 (O_1311,N_22798,N_22393);
nor UO_1312 (O_1312,N_23624,N_24999);
nor UO_1313 (O_1313,N_24214,N_20021);
nand UO_1314 (O_1314,N_23583,N_22667);
xor UO_1315 (O_1315,N_21371,N_20930);
nor UO_1316 (O_1316,N_24089,N_24595);
xor UO_1317 (O_1317,N_23160,N_23197);
or UO_1318 (O_1318,N_24264,N_23236);
or UO_1319 (O_1319,N_20947,N_24000);
nor UO_1320 (O_1320,N_21784,N_24063);
xor UO_1321 (O_1321,N_21317,N_21962);
and UO_1322 (O_1322,N_22292,N_22330);
xnor UO_1323 (O_1323,N_24082,N_22125);
and UO_1324 (O_1324,N_22961,N_22322);
nor UO_1325 (O_1325,N_22859,N_20043);
or UO_1326 (O_1326,N_22948,N_22075);
or UO_1327 (O_1327,N_21250,N_24913);
or UO_1328 (O_1328,N_21882,N_20859);
or UO_1329 (O_1329,N_24950,N_24952);
or UO_1330 (O_1330,N_23966,N_24609);
and UO_1331 (O_1331,N_20991,N_20166);
or UO_1332 (O_1332,N_22495,N_22860);
and UO_1333 (O_1333,N_24043,N_21943);
xor UO_1334 (O_1334,N_22771,N_20856);
nand UO_1335 (O_1335,N_22199,N_20654);
and UO_1336 (O_1336,N_22611,N_23944);
or UO_1337 (O_1337,N_24447,N_24263);
and UO_1338 (O_1338,N_22718,N_21762);
nor UO_1339 (O_1339,N_20997,N_24553);
nand UO_1340 (O_1340,N_22982,N_24286);
nor UO_1341 (O_1341,N_22206,N_24087);
nand UO_1342 (O_1342,N_23888,N_22256);
and UO_1343 (O_1343,N_21918,N_24235);
xor UO_1344 (O_1344,N_23806,N_24634);
xnor UO_1345 (O_1345,N_22556,N_22323);
nand UO_1346 (O_1346,N_20789,N_24058);
nor UO_1347 (O_1347,N_22239,N_24002);
and UO_1348 (O_1348,N_22542,N_20992);
or UO_1349 (O_1349,N_21286,N_20815);
or UO_1350 (O_1350,N_22546,N_23891);
nor UO_1351 (O_1351,N_23539,N_22952);
and UO_1352 (O_1352,N_24345,N_21487);
xor UO_1353 (O_1353,N_21403,N_21590);
and UO_1354 (O_1354,N_20840,N_22991);
nand UO_1355 (O_1355,N_20554,N_20088);
nand UO_1356 (O_1356,N_24138,N_23525);
nand UO_1357 (O_1357,N_22506,N_20049);
nand UO_1358 (O_1358,N_24930,N_22328);
and UO_1359 (O_1359,N_22717,N_21476);
and UO_1360 (O_1360,N_22332,N_20931);
nand UO_1361 (O_1361,N_21555,N_21576);
nand UO_1362 (O_1362,N_20538,N_21556);
and UO_1363 (O_1363,N_21163,N_24190);
nand UO_1364 (O_1364,N_23569,N_24559);
nand UO_1365 (O_1365,N_20728,N_23801);
and UO_1366 (O_1366,N_22919,N_22761);
and UO_1367 (O_1367,N_20568,N_24701);
nor UO_1368 (O_1368,N_22451,N_21150);
nand UO_1369 (O_1369,N_22724,N_23341);
nand UO_1370 (O_1370,N_20513,N_22993);
and UO_1371 (O_1371,N_20082,N_22965);
nor UO_1372 (O_1372,N_20002,N_24493);
nand UO_1373 (O_1373,N_22942,N_22387);
and UO_1374 (O_1374,N_24033,N_20156);
xor UO_1375 (O_1375,N_23771,N_22969);
or UO_1376 (O_1376,N_21136,N_20037);
or UO_1377 (O_1377,N_23111,N_22259);
nand UO_1378 (O_1378,N_21274,N_24898);
or UO_1379 (O_1379,N_20672,N_22812);
nand UO_1380 (O_1380,N_24991,N_21341);
or UO_1381 (O_1381,N_21126,N_20912);
xnor UO_1382 (O_1382,N_21873,N_21620);
nor UO_1383 (O_1383,N_21372,N_22271);
nand UO_1384 (O_1384,N_24270,N_20641);
and UO_1385 (O_1385,N_21097,N_22464);
and UO_1386 (O_1386,N_23497,N_23328);
xnor UO_1387 (O_1387,N_21513,N_21336);
or UO_1388 (O_1388,N_23027,N_21075);
nor UO_1389 (O_1389,N_24882,N_23420);
xnor UO_1390 (O_1390,N_22990,N_23193);
nand UO_1391 (O_1391,N_20318,N_24588);
xor UO_1392 (O_1392,N_23602,N_22526);
and UO_1393 (O_1393,N_20028,N_22375);
or UO_1394 (O_1394,N_23184,N_24790);
or UO_1395 (O_1395,N_23876,N_20277);
nor UO_1396 (O_1396,N_22821,N_21613);
and UO_1397 (O_1397,N_21275,N_21014);
or UO_1398 (O_1398,N_23837,N_23491);
nor UO_1399 (O_1399,N_21440,N_20065);
or UO_1400 (O_1400,N_21173,N_24783);
nand UO_1401 (O_1401,N_24353,N_22142);
nor UO_1402 (O_1402,N_22568,N_24195);
and UO_1403 (O_1403,N_21566,N_23996);
nor UO_1404 (O_1404,N_22768,N_21936);
or UO_1405 (O_1405,N_22802,N_24132);
and UO_1406 (O_1406,N_21718,N_20727);
and UO_1407 (O_1407,N_21360,N_20769);
nand UO_1408 (O_1408,N_20964,N_21648);
or UO_1409 (O_1409,N_20237,N_20205);
and UO_1410 (O_1410,N_22851,N_23871);
nand UO_1411 (O_1411,N_22894,N_20617);
xnor UO_1412 (O_1412,N_24303,N_23296);
or UO_1413 (O_1413,N_21827,N_22469);
nand UO_1414 (O_1414,N_20662,N_24478);
or UO_1415 (O_1415,N_20715,N_21247);
xnor UO_1416 (O_1416,N_24929,N_21128);
and UO_1417 (O_1417,N_22207,N_20914);
xor UO_1418 (O_1418,N_20822,N_21204);
xnor UO_1419 (O_1419,N_21262,N_22868);
nand UO_1420 (O_1420,N_21182,N_21203);
xor UO_1421 (O_1421,N_21207,N_20770);
nor UO_1422 (O_1422,N_20342,N_20279);
or UO_1423 (O_1423,N_23293,N_24016);
xor UO_1424 (O_1424,N_24358,N_22201);
nand UO_1425 (O_1425,N_23748,N_21284);
nor UO_1426 (O_1426,N_23827,N_23936);
or UO_1427 (O_1427,N_22157,N_24961);
and UO_1428 (O_1428,N_23345,N_22876);
xor UO_1429 (O_1429,N_23417,N_23091);
xnor UO_1430 (O_1430,N_24218,N_20192);
nand UO_1431 (O_1431,N_22315,N_23589);
nor UO_1432 (O_1432,N_24102,N_22442);
or UO_1433 (O_1433,N_24007,N_24943);
or UO_1434 (O_1434,N_21991,N_24171);
or UO_1435 (O_1435,N_22759,N_21505);
or UO_1436 (O_1436,N_22232,N_21664);
nand UO_1437 (O_1437,N_24160,N_24203);
and UO_1438 (O_1438,N_22754,N_21443);
or UO_1439 (O_1439,N_21938,N_22340);
xor UO_1440 (O_1440,N_24649,N_24331);
or UO_1441 (O_1441,N_23682,N_20195);
or UO_1442 (O_1442,N_21363,N_20235);
and UO_1443 (O_1443,N_22354,N_22987);
nand UO_1444 (O_1444,N_23029,N_21119);
nor UO_1445 (O_1445,N_22432,N_23243);
xor UO_1446 (O_1446,N_24440,N_21601);
xor UO_1447 (O_1447,N_24770,N_24338);
or UO_1448 (O_1448,N_24237,N_21287);
nand UO_1449 (O_1449,N_20215,N_22365);
or UO_1450 (O_1450,N_20881,N_20004);
xor UO_1451 (O_1451,N_22653,N_23716);
nand UO_1452 (O_1452,N_23079,N_22410);
and UO_1453 (O_1453,N_24022,N_21752);
and UO_1454 (O_1454,N_21562,N_24647);
nor UO_1455 (O_1455,N_24906,N_20155);
and UO_1456 (O_1456,N_24631,N_22244);
and UO_1457 (O_1457,N_20742,N_21259);
nor UO_1458 (O_1458,N_24013,N_22109);
nor UO_1459 (O_1459,N_22988,N_24587);
nor UO_1460 (O_1460,N_24621,N_24546);
and UO_1461 (O_1461,N_23291,N_20767);
xnor UO_1462 (O_1462,N_24673,N_22430);
nand UO_1463 (O_1463,N_23726,N_21878);
nand UO_1464 (O_1464,N_24759,N_23213);
xnor UO_1465 (O_1465,N_22132,N_21790);
or UO_1466 (O_1466,N_23951,N_21305);
nor UO_1467 (O_1467,N_24107,N_22107);
or UO_1468 (O_1468,N_23278,N_21830);
nand UO_1469 (O_1469,N_20083,N_22956);
nand UO_1470 (O_1470,N_20295,N_20337);
or UO_1471 (O_1471,N_20920,N_24072);
nor UO_1472 (O_1472,N_21535,N_24114);
nand UO_1473 (O_1473,N_24317,N_20424);
and UO_1474 (O_1474,N_24362,N_21003);
xor UO_1475 (O_1475,N_20821,N_20751);
or UO_1476 (O_1476,N_24915,N_24023);
nor UO_1477 (O_1477,N_22748,N_22654);
nand UO_1478 (O_1478,N_23894,N_22689);
nand UO_1479 (O_1479,N_24360,N_20693);
or UO_1480 (O_1480,N_21897,N_21384);
and UO_1481 (O_1481,N_20260,N_20816);
nand UO_1482 (O_1482,N_21619,N_20766);
and UO_1483 (O_1483,N_21038,N_22300);
nand UO_1484 (O_1484,N_21714,N_21560);
nor UO_1485 (O_1485,N_22218,N_24092);
or UO_1486 (O_1486,N_21015,N_24394);
and UO_1487 (O_1487,N_21447,N_20578);
nand UO_1488 (O_1488,N_23991,N_20527);
nor UO_1489 (O_1489,N_22246,N_23035);
or UO_1490 (O_1490,N_24232,N_23280);
nand UO_1491 (O_1491,N_23402,N_24446);
xnor UO_1492 (O_1492,N_22058,N_21060);
and UO_1493 (O_1493,N_23532,N_23819);
xnor UO_1494 (O_1494,N_23942,N_21569);
nor UO_1495 (O_1495,N_20832,N_22844);
nand UO_1496 (O_1496,N_21424,N_22362);
xor UO_1497 (O_1497,N_23070,N_22544);
nor UO_1498 (O_1498,N_20018,N_23173);
or UO_1499 (O_1499,N_22862,N_23889);
nand UO_1500 (O_1500,N_20127,N_21981);
nor UO_1501 (O_1501,N_24079,N_23298);
or UO_1502 (O_1502,N_22337,N_21855);
nor UO_1503 (O_1503,N_23645,N_22405);
xor UO_1504 (O_1504,N_21695,N_20372);
or UO_1505 (O_1505,N_23504,N_20241);
and UO_1506 (O_1506,N_22099,N_24450);
xor UO_1507 (O_1507,N_22684,N_23475);
nor UO_1508 (O_1508,N_23761,N_24890);
and UO_1509 (O_1509,N_20735,N_24499);
xnor UO_1510 (O_1510,N_20540,N_24052);
nand UO_1511 (O_1511,N_20942,N_20185);
and UO_1512 (O_1512,N_21970,N_21747);
nor UO_1513 (O_1513,N_21024,N_21482);
and UO_1514 (O_1514,N_21303,N_24556);
nand UO_1515 (O_1515,N_20807,N_23357);
nand UO_1516 (O_1516,N_23500,N_22578);
and UO_1517 (O_1517,N_23149,N_23816);
or UO_1518 (O_1518,N_20441,N_20276);
and UO_1519 (O_1519,N_20419,N_24346);
nand UO_1520 (O_1520,N_21489,N_22594);
nand UO_1521 (O_1521,N_21406,N_20946);
xnor UO_1522 (O_1522,N_22252,N_20369);
xnor UO_1523 (O_1523,N_23887,N_22911);
nor UO_1524 (O_1524,N_24988,N_22642);
nor UO_1525 (O_1525,N_22606,N_21298);
nand UO_1526 (O_1526,N_20504,N_24407);
nor UO_1527 (O_1527,N_21876,N_20468);
and UO_1528 (O_1528,N_23260,N_20110);
and UO_1529 (O_1529,N_22883,N_22460);
nor UO_1530 (O_1530,N_20114,N_22101);
and UO_1531 (O_1531,N_22801,N_24404);
or UO_1532 (O_1532,N_20493,N_21874);
and UO_1533 (O_1533,N_24115,N_20045);
or UO_1534 (O_1534,N_22530,N_21404);
xor UO_1535 (O_1535,N_22287,N_21927);
nor UO_1536 (O_1536,N_22666,N_20798);
nand UO_1537 (O_1537,N_22133,N_21324);
or UO_1538 (O_1538,N_24413,N_23226);
xnor UO_1539 (O_1539,N_21606,N_24238);
or UO_1540 (O_1540,N_20826,N_22516);
xor UO_1541 (O_1541,N_24442,N_20379);
or UO_1542 (O_1542,N_21448,N_24251);
and UO_1543 (O_1543,N_23414,N_23686);
or UO_1544 (O_1544,N_20884,N_22243);
xor UO_1545 (O_1545,N_22296,N_24403);
nor UO_1546 (O_1546,N_22600,N_22554);
nand UO_1547 (O_1547,N_24694,N_20148);
or UO_1548 (O_1548,N_20909,N_24574);
and UO_1549 (O_1549,N_20415,N_22077);
and UO_1550 (O_1550,N_23960,N_21901);
xnor UO_1551 (O_1551,N_20080,N_21145);
nand UO_1552 (O_1552,N_22283,N_24733);
nand UO_1553 (O_1553,N_22680,N_20213);
and UO_1554 (O_1554,N_23965,N_22150);
xnor UO_1555 (O_1555,N_21755,N_24354);
nand UO_1556 (O_1556,N_24322,N_22262);
or UO_1557 (O_1557,N_21456,N_23518);
xor UO_1558 (O_1558,N_20225,N_24299);
nor UO_1559 (O_1559,N_24131,N_21799);
nor UO_1560 (O_1560,N_21773,N_21839);
xnor UO_1561 (O_1561,N_24477,N_20819);
nand UO_1562 (O_1562,N_24928,N_20229);
nor UO_1563 (O_1563,N_20567,N_21546);
nor UO_1564 (O_1564,N_20643,N_24490);
nor UO_1565 (O_1565,N_23917,N_23429);
nand UO_1566 (O_1566,N_23654,N_22615);
nor UO_1567 (O_1567,N_22773,N_23299);
and UO_1568 (O_1568,N_22457,N_24748);
and UO_1569 (O_1569,N_24318,N_23270);
and UO_1570 (O_1570,N_24188,N_23785);
and UO_1571 (O_1571,N_21697,N_23659);
and UO_1572 (O_1572,N_24743,N_21930);
nand UO_1573 (O_1573,N_23274,N_21357);
xor UO_1574 (O_1574,N_20609,N_22404);
xor UO_1575 (O_1575,N_21650,N_24503);
nor UO_1576 (O_1576,N_23467,N_24015);
xor UO_1577 (O_1577,N_23901,N_22502);
nor UO_1578 (O_1578,N_24472,N_20117);
nand UO_1579 (O_1579,N_23946,N_23120);
and UO_1580 (O_1580,N_20569,N_21009);
or UO_1581 (O_1581,N_23253,N_20003);
nor UO_1582 (O_1582,N_22369,N_20989);
nor UO_1583 (O_1583,N_21442,N_22577);
nand UO_1584 (O_1584,N_22701,N_20272);
nor UO_1585 (O_1585,N_23294,N_23110);
or UO_1586 (O_1586,N_20625,N_21392);
or UO_1587 (O_1587,N_24823,N_24049);
nor UO_1588 (O_1588,N_23949,N_22559);
nand UO_1589 (O_1589,N_24307,N_22891);
and UO_1590 (O_1590,N_24951,N_23738);
nand UO_1591 (O_1591,N_21011,N_24990);
and UO_1592 (O_1592,N_20934,N_20089);
nor UO_1593 (O_1593,N_24193,N_23561);
nand UO_1594 (O_1594,N_22023,N_22461);
xor UO_1595 (O_1595,N_20389,N_24142);
or UO_1596 (O_1596,N_24050,N_24046);
nor UO_1597 (O_1597,N_24310,N_22468);
nand UO_1598 (O_1598,N_21050,N_20698);
nor UO_1599 (O_1599,N_24323,N_24432);
and UO_1600 (O_1600,N_20624,N_20395);
nand UO_1601 (O_1601,N_20450,N_22902);
nand UO_1602 (O_1602,N_24774,N_22763);
nand UO_1603 (O_1603,N_22436,N_21766);
nand UO_1604 (O_1604,N_22916,N_24985);
nand UO_1605 (O_1605,N_22879,N_23895);
nand UO_1606 (O_1606,N_20824,N_21895);
nor UO_1607 (O_1607,N_23903,N_23480);
nand UO_1608 (O_1608,N_23276,N_23870);
or UO_1609 (O_1609,N_23779,N_21586);
and UO_1610 (O_1610,N_23095,N_22747);
or UO_1611 (O_1611,N_20239,N_22540);
nand UO_1612 (O_1612,N_24856,N_21025);
nor UO_1613 (O_1613,N_21256,N_21318);
or UO_1614 (O_1614,N_24164,N_23258);
nand UO_1615 (O_1615,N_24068,N_21743);
and UO_1616 (O_1616,N_23879,N_20894);
xor UO_1617 (O_1617,N_22963,N_22895);
nand UO_1618 (O_1618,N_23701,N_20128);
xor UO_1619 (O_1619,N_23472,N_24855);
or UO_1620 (O_1620,N_20025,N_20996);
nor UO_1621 (O_1621,N_20300,N_20577);
xor UO_1622 (O_1622,N_24517,N_23702);
nand UO_1623 (O_1623,N_23614,N_24128);
and UO_1624 (O_1624,N_22958,N_20483);
and UO_1625 (O_1625,N_24294,N_22767);
and UO_1626 (O_1626,N_24161,N_21888);
nand UO_1627 (O_1627,N_22477,N_21663);
nand UO_1628 (O_1628,N_22019,N_22445);
or UO_1629 (O_1629,N_20013,N_23939);
and UO_1630 (O_1630,N_21733,N_23952);
nand UO_1631 (O_1631,N_24607,N_23732);
xnor UO_1632 (O_1632,N_22397,N_20446);
xor UO_1633 (O_1633,N_24709,N_22163);
and UO_1634 (O_1634,N_24392,N_24271);
and UO_1635 (O_1635,N_22864,N_22907);
or UO_1636 (O_1636,N_21871,N_21514);
nand UO_1637 (O_1637,N_23077,N_20184);
or UO_1638 (O_1638,N_23399,N_22670);
or UO_1639 (O_1639,N_24986,N_24488);
and UO_1640 (O_1640,N_23128,N_20187);
xor UO_1641 (O_1641,N_24122,N_21219);
nor UO_1642 (O_1642,N_24962,N_24657);
and UO_1643 (O_1643,N_22913,N_21471);
nor UO_1644 (O_1644,N_22061,N_21091);
and UO_1645 (O_1645,N_23481,N_22944);
nand UO_1646 (O_1646,N_24175,N_21967);
nor UO_1647 (O_1647,N_20985,N_20268);
xnor UO_1648 (O_1648,N_23369,N_24205);
or UO_1649 (O_1649,N_23580,N_20374);
nand UO_1650 (O_1650,N_24854,N_24086);
or UO_1651 (O_1651,N_23478,N_23205);
and UO_1652 (O_1652,N_20586,N_23239);
nand UO_1653 (O_1653,N_23262,N_24599);
or UO_1654 (O_1654,N_24674,N_21042);
nor UO_1655 (O_1655,N_22145,N_20764);
nand UO_1656 (O_1656,N_22366,N_20090);
xnor UO_1657 (O_1657,N_22003,N_23432);
nand UO_1658 (O_1658,N_24797,N_21366);
and UO_1659 (O_1659,N_22909,N_23055);
xnor UO_1660 (O_1660,N_21595,N_20782);
xnor UO_1661 (O_1661,N_23387,N_23376);
nor UO_1662 (O_1662,N_23113,N_22278);
nand UO_1663 (O_1663,N_24995,N_24139);
nand UO_1664 (O_1664,N_23933,N_23797);
or UO_1665 (O_1665,N_23592,N_21121);
xnor UO_1666 (O_1666,N_24758,N_20234);
xnor UO_1667 (O_1667,N_22196,N_24964);
nand UO_1668 (O_1668,N_22924,N_21054);
and UO_1669 (O_1669,N_24794,N_22562);
nand UO_1670 (O_1670,N_23044,N_24098);
nand UO_1671 (O_1671,N_24741,N_20694);
nor UO_1672 (O_1672,N_23474,N_21795);
and UO_1673 (O_1673,N_21700,N_23555);
nor UO_1674 (O_1674,N_24004,N_23455);
nor UO_1675 (O_1675,N_23869,N_20978);
nor UO_1676 (O_1676,N_20072,N_21178);
or UO_1677 (O_1677,N_20825,N_23703);
xor UO_1678 (O_1678,N_20585,N_20421);
or UO_1679 (O_1679,N_20949,N_22402);
xnor UO_1680 (O_1680,N_22498,N_22822);
or UO_1681 (O_1681,N_22949,N_22590);
nor UO_1682 (O_1682,N_21803,N_24987);
xnor UO_1683 (O_1683,N_21254,N_21299);
nand UO_1684 (O_1684,N_23523,N_22108);
nand UO_1685 (O_1685,N_24716,N_24789);
nor UO_1686 (O_1686,N_24523,N_20257);
or UO_1687 (O_1687,N_23923,N_23155);
xnor UO_1688 (O_1688,N_21144,N_20451);
xor UO_1689 (O_1689,N_22364,N_23851);
xor UO_1690 (O_1690,N_24644,N_22236);
nand UO_1691 (O_1691,N_23810,N_20519);
nand UO_1692 (O_1692,N_24327,N_24989);
xor UO_1693 (O_1693,N_20895,N_24196);
nor UO_1694 (O_1694,N_24592,N_20505);
nor UO_1695 (O_1695,N_20758,N_24960);
or UO_1696 (O_1696,N_23924,N_24700);
nor UO_1697 (O_1697,N_21842,N_22415);
xnor UO_1698 (O_1698,N_22414,N_24892);
and UO_1699 (O_1699,N_21088,N_20248);
xnor UO_1700 (O_1700,N_24659,N_21944);
nor UO_1701 (O_1701,N_20482,N_23697);
or UO_1702 (O_1702,N_21012,N_23007);
nor UO_1703 (O_1703,N_22088,N_24074);
nand UO_1704 (O_1704,N_23014,N_24531);
nor UO_1705 (O_1705,N_22116,N_22248);
nand UO_1706 (O_1706,N_21421,N_20223);
nand UO_1707 (O_1707,N_22189,N_24719);
and UO_1708 (O_1708,N_20974,N_20621);
and UO_1709 (O_1709,N_20732,N_21127);
and UO_1710 (O_1710,N_20775,N_23892);
xnor UO_1711 (O_1711,N_22815,N_20622);
nor UO_1712 (O_1712,N_20918,N_22605);
and UO_1713 (O_1713,N_20010,N_24957);
nand UO_1714 (O_1714,N_22996,N_23579);
nor UO_1715 (O_1715,N_23316,N_22032);
xor UO_1716 (O_1716,N_23975,N_24642);
or UO_1717 (O_1717,N_22778,N_22817);
and UO_1718 (O_1718,N_20435,N_21706);
xor UO_1719 (O_1719,N_24200,N_20784);
nor UO_1720 (O_1720,N_20423,N_21904);
nand UO_1721 (O_1721,N_20741,N_23078);
nand UO_1722 (O_1722,N_24520,N_20687);
or UO_1723 (O_1723,N_20591,N_20917);
nand UO_1724 (O_1724,N_24539,N_23374);
nor UO_1725 (O_1725,N_20862,N_22052);
or UO_1726 (O_1726,N_23710,N_23841);
nand UO_1727 (O_1727,N_23631,N_24253);
or UO_1728 (O_1728,N_24579,N_22915);
or UO_1729 (O_1729,N_23813,N_24680);
nand UO_1730 (O_1730,N_21206,N_24334);
and UO_1731 (O_1731,N_23001,N_22013);
and UO_1732 (O_1732,N_20390,N_21485);
xnor UO_1733 (O_1733,N_20640,N_24828);
nor UO_1734 (O_1734,N_22737,N_21181);
and UO_1735 (O_1735,N_21879,N_20510);
or UO_1736 (O_1736,N_21292,N_23271);
nor UO_1737 (O_1737,N_22017,N_20663);
nor UO_1738 (O_1738,N_21020,N_20190);
nand UO_1739 (O_1739,N_20837,N_20416);
and UO_1740 (O_1740,N_20298,N_22458);
xnor UO_1741 (O_1741,N_20890,N_22535);
and UO_1742 (O_1742,N_21276,N_24581);
nand UO_1743 (O_1743,N_22607,N_23390);
or UO_1744 (O_1744,N_23272,N_21917);
nand UO_1745 (O_1745,N_20701,N_20074);
and UO_1746 (O_1746,N_24381,N_24809);
or UO_1747 (O_1747,N_24445,N_21308);
xnor UO_1748 (O_1748,N_22205,N_24398);
or UO_1749 (O_1749,N_20757,N_21777);
nor UO_1750 (O_1750,N_23463,N_24245);
and UO_1751 (O_1751,N_20141,N_21852);
xor UO_1752 (O_1752,N_20829,N_20925);
xnor UO_1753 (O_1753,N_20181,N_24919);
nand UO_1754 (O_1754,N_24032,N_23146);
and UO_1755 (O_1755,N_21064,N_24406);
or UO_1756 (O_1756,N_20271,N_23751);
and UO_1757 (O_1757,N_20745,N_20431);
and UO_1758 (O_1758,N_23122,N_23034);
nor UO_1759 (O_1759,N_24513,N_23596);
nor UO_1760 (O_1760,N_20810,N_24153);
xnor UO_1761 (O_1761,N_24835,N_22686);
or UO_1762 (O_1762,N_23263,N_23787);
and UO_1763 (O_1763,N_23440,N_20607);
xnor UO_1764 (O_1764,N_22040,N_24670);
or UO_1765 (O_1765,N_22592,N_24152);
nand UO_1766 (O_1766,N_23556,N_20966);
or UO_1767 (O_1767,N_23843,N_22035);
nand UO_1768 (O_1768,N_21713,N_22630);
nand UO_1769 (O_1769,N_20105,N_21947);
xor UO_1770 (O_1770,N_20619,N_24301);
nand UO_1771 (O_1771,N_23637,N_23809);
nand UO_1772 (O_1772,N_20455,N_23510);
nand UO_1773 (O_1773,N_22374,N_22131);
nand UO_1774 (O_1774,N_21760,N_23747);
or UO_1775 (O_1775,N_24658,N_22626);
nand UO_1776 (O_1776,N_24544,N_21703);
and UO_1777 (O_1777,N_24408,N_23261);
or UO_1778 (O_1778,N_21780,N_22429);
or UO_1779 (O_1779,N_23391,N_21954);
nor UO_1780 (O_1780,N_22646,N_20132);
or UO_1781 (O_1781,N_20418,N_23673);
nand UO_1782 (O_1782,N_24348,N_23699);
or UO_1783 (O_1783,N_22059,N_23375);
and UO_1784 (O_1784,N_22063,N_23006);
and UO_1785 (O_1785,N_20152,N_23223);
xnor UO_1786 (O_1786,N_20501,N_21519);
xor UO_1787 (O_1787,N_23545,N_22455);
nor UO_1788 (O_1788,N_22043,N_21246);
nor UO_1789 (O_1789,N_24940,N_23319);
xnor UO_1790 (O_1790,N_24005,N_22598);
nor UO_1791 (O_1791,N_21498,N_21039);
nand UO_1792 (O_1792,N_20999,N_21881);
nand UO_1793 (O_1793,N_21232,N_22977);
or UO_1794 (O_1794,N_24225,N_22608);
xor UO_1795 (O_1795,N_22345,N_23323);
xor UO_1796 (O_1796,N_20719,N_24021);
or UO_1797 (O_1797,N_21638,N_20739);
nand UO_1798 (O_1798,N_23124,N_20073);
nand UO_1799 (O_1799,N_22668,N_20876);
nor UO_1800 (O_1800,N_20267,N_20953);
and UO_1801 (O_1801,N_20115,N_20860);
nand UO_1802 (O_1802,N_21798,N_23511);
xor UO_1803 (O_1803,N_23986,N_22305);
nand UO_1804 (O_1804,N_23285,N_21870);
nand UO_1805 (O_1805,N_23112,N_21676);
nand UO_1806 (O_1806,N_23487,N_21811);
nand UO_1807 (O_1807,N_23814,N_24228);
nand UO_1808 (O_1808,N_21630,N_20162);
nor UO_1809 (O_1809,N_23108,N_24883);
xor UO_1810 (O_1810,N_22155,N_21486);
and UO_1811 (O_1811,N_21331,N_20614);
nor UO_1812 (O_1812,N_21692,N_23823);
nor UO_1813 (O_1813,N_20027,N_24433);
nand UO_1814 (O_1814,N_23762,N_23257);
xor UO_1815 (O_1815,N_24859,N_20980);
or UO_1816 (O_1816,N_21433,N_23988);
nand UO_1817 (O_1817,N_20597,N_24031);
xnor UO_1818 (O_1818,N_20534,N_21934);
nor UO_1819 (O_1819,N_22673,N_24095);
nand UO_1820 (O_1820,N_23227,N_22349);
and UO_1821 (O_1821,N_20008,N_22933);
or UO_1822 (O_1822,N_24044,N_20848);
and UO_1823 (O_1823,N_23395,N_24067);
nand UO_1824 (O_1824,N_22138,N_24640);
nand UO_1825 (O_1825,N_23756,N_24265);
nand UO_1826 (O_1826,N_22250,N_24293);
nand UO_1827 (O_1827,N_20366,N_21659);
nor UO_1828 (O_1828,N_23731,N_22983);
xor UO_1829 (O_1829,N_21132,N_23769);
nor UO_1830 (O_1830,N_22786,N_23883);
and UO_1831 (O_1831,N_22441,N_24320);
xnor UO_1832 (O_1832,N_23230,N_24916);
or UO_1833 (O_1833,N_24018,N_22936);
or UO_1834 (O_1834,N_21683,N_23286);
or UO_1835 (O_1835,N_24308,N_24486);
and UO_1836 (O_1836,N_20849,N_21230);
xnor UO_1837 (O_1837,N_23698,N_22931);
nor UO_1838 (O_1838,N_24624,N_23718);
or UO_1839 (O_1839,N_24213,N_22186);
xor UO_1840 (O_1840,N_20439,N_24684);
or UO_1841 (O_1841,N_23691,N_24137);
nor UO_1842 (O_1842,N_21853,N_22521);
nor UO_1843 (O_1843,N_24352,N_20763);
or UO_1844 (O_1844,N_22379,N_21953);
nor UO_1845 (O_1845,N_21813,N_21451);
and UO_1846 (O_1846,N_24096,N_20212);
nor UO_1847 (O_1847,N_20250,N_21902);
or UO_1848 (O_1848,N_21346,N_20252);
and UO_1849 (O_1849,N_20932,N_22030);
nor UO_1850 (O_1850,N_21224,N_24233);
and UO_1851 (O_1851,N_23913,N_23859);
and UO_1852 (O_1852,N_23753,N_24291);
and UO_1853 (O_1853,N_20376,N_24720);
nand UO_1854 (O_1854,N_21926,N_23627);
xnor UO_1855 (O_1855,N_24696,N_21474);
and UO_1856 (O_1856,N_21068,N_21340);
nand UO_1857 (O_1857,N_24099,N_24586);
and UO_1858 (O_1858,N_22491,N_24620);
or UO_1859 (O_1859,N_24688,N_20174);
nand UO_1860 (O_1860,N_21479,N_22978);
or UO_1861 (O_1861,N_23019,N_23570);
nor UO_1862 (O_1862,N_24146,N_21796);
nor UO_1863 (O_1863,N_20574,N_21957);
xor UO_1864 (O_1864,N_21239,N_20227);
and UO_1865 (O_1865,N_24144,N_22708);
xnor UO_1866 (O_1866,N_24378,N_23069);
xnor UO_1867 (O_1867,N_24678,N_24212);
xnor UO_1868 (O_1868,N_21030,N_23671);
or UO_1869 (O_1869,N_24762,N_23616);
and UO_1870 (O_1870,N_21741,N_20348);
nand UO_1871 (O_1871,N_23394,N_24912);
xnor UO_1872 (O_1872,N_20048,N_24029);
nand UO_1873 (O_1873,N_20861,N_23371);
nand UO_1874 (O_1874,N_22403,N_20983);
or UO_1875 (O_1875,N_21416,N_24365);
and UO_1876 (O_1876,N_23930,N_22463);
nand UO_1877 (O_1877,N_24108,N_21862);
and UO_1878 (O_1878,N_21631,N_20361);
xnor UO_1879 (O_1879,N_21029,N_23215);
nand UO_1880 (O_1880,N_24839,N_20650);
or UO_1881 (O_1881,N_21185,N_21045);
and UO_1882 (O_1882,N_21952,N_21922);
xor UO_1883 (O_1883,N_24458,N_24239);
xor UO_1884 (O_1884,N_23746,N_22385);
xor UO_1885 (O_1885,N_24170,N_21083);
xnor UO_1886 (O_1886,N_20111,N_23137);
and UO_1887 (O_1887,N_23945,N_23705);
nor UO_1888 (O_1888,N_23752,N_21921);
xnor UO_1889 (O_1889,N_21189,N_24702);
nand UO_1890 (O_1890,N_21793,N_23628);
nor UO_1891 (O_1891,N_20472,N_22117);
and UO_1892 (O_1892,N_22892,N_21704);
nor UO_1893 (O_1893,N_24656,N_22290);
xnor UO_1894 (O_1894,N_20771,N_20498);
nor UO_1895 (O_1895,N_23162,N_20206);
and UO_1896 (O_1896,N_21044,N_20447);
xor UO_1897 (O_1897,N_22946,N_23339);
xnor UO_1898 (O_1898,N_24080,N_20970);
nor UO_1899 (O_1899,N_22601,N_23864);
and UO_1900 (O_1900,N_22610,N_20029);
nand UO_1901 (O_1901,N_20291,N_23132);
and UO_1902 (O_1902,N_24252,N_24760);
and UO_1903 (O_1903,N_23544,N_23855);
and UO_1904 (O_1904,N_21792,N_20637);
nand UO_1905 (O_1905,N_21087,N_24727);
nand UO_1906 (O_1906,N_23808,N_23735);
and UO_1907 (O_1907,N_20033,N_20302);
or UO_1908 (O_1908,N_23334,N_20633);
nor UO_1909 (O_1909,N_22637,N_20015);
and UO_1910 (O_1910,N_20520,N_23000);
or UO_1911 (O_1911,N_23383,N_24090);
or UO_1912 (O_1912,N_23460,N_22230);
nor UO_1913 (O_1913,N_21608,N_23249);
xor UO_1914 (O_1914,N_20321,N_21673);
and UO_1915 (O_1915,N_21685,N_21313);
nand UO_1916 (O_1916,N_21348,N_24690);
and UO_1917 (O_1917,N_22057,N_21858);
nor UO_1918 (O_1918,N_20307,N_20915);
xor UO_1919 (O_1919,N_23256,N_22789);
or UO_1920 (O_1920,N_20502,N_24418);
or UO_1921 (O_1921,N_20309,N_23626);
and UO_1922 (O_1922,N_22370,N_21102);
or UO_1923 (O_1923,N_20349,N_23045);
nor UO_1924 (O_1924,N_22538,N_20801);
nand UO_1925 (O_1925,N_22437,N_24518);
and UO_1926 (O_1926,N_21302,N_22863);
nor UO_1927 (O_1927,N_24780,N_21856);
nand UO_1928 (O_1928,N_23577,N_24881);
and UO_1929 (O_1929,N_23461,N_21131);
or UO_1930 (O_1930,N_23741,N_24910);
nand UO_1931 (O_1931,N_24289,N_23384);
and UO_1932 (O_1932,N_23281,N_21205);
nand UO_1933 (O_1933,N_20885,N_22672);
nand UO_1934 (O_1934,N_24655,N_20630);
and UO_1935 (O_1935,N_20011,N_23041);
and UO_1936 (O_1936,N_23165,N_22213);
nor UO_1937 (O_1937,N_22805,N_24614);
nand UO_1938 (O_1938,N_24920,N_23030);
xor UO_1939 (O_1939,N_23540,N_20655);
nand UO_1940 (O_1940,N_23141,N_24485);
nand UO_1941 (O_1941,N_20204,N_21624);
nor UO_1942 (O_1942,N_24663,N_21165);
xnor UO_1943 (O_1943,N_24275,N_24810);
nor UO_1944 (O_1944,N_20044,N_22188);
nor UO_1945 (O_1945,N_21135,N_20175);
nand UO_1946 (O_1946,N_20079,N_22930);
and UO_1947 (O_1947,N_20462,N_23489);
nand UO_1948 (O_1948,N_22807,N_21221);
nor UO_1949 (O_1949,N_22522,N_23074);
or UO_1950 (O_1950,N_21294,N_24025);
nand UO_1951 (O_1951,N_20689,N_24942);
nand UO_1952 (O_1952,N_21618,N_22792);
and UO_1953 (O_1953,N_20216,N_22482);
and UO_1954 (O_1954,N_22424,N_24630);
nand UO_1955 (O_1955,N_22331,N_23468);
nor UO_1956 (O_1956,N_21072,N_21751);
or UO_1957 (O_1957,N_22181,N_22709);
xor UO_1958 (O_1958,N_22042,N_23087);
and UO_1959 (O_1959,N_20618,N_22645);
xor UO_1960 (O_1960,N_21347,N_22154);
or UO_1961 (O_1961,N_21457,N_24867);
nor UO_1962 (O_1962,N_20573,N_22826);
and UO_1963 (O_1963,N_22055,N_20017);
and UO_1964 (O_1964,N_21763,N_23780);
or UO_1965 (O_1965,N_23147,N_22193);
nor UO_1966 (O_1966,N_21335,N_24801);
or UO_1967 (O_1967,N_21993,N_23860);
nor UO_1968 (O_1968,N_20377,N_20587);
nand UO_1969 (O_1969,N_20765,N_22294);
xnor UO_1970 (O_1970,N_22532,N_24451);
or UO_1971 (O_1971,N_21678,N_22833);
xnor UO_1972 (O_1972,N_21110,N_21393);
xnor UO_1973 (O_1973,N_24865,N_20673);
or UO_1974 (O_1974,N_21493,N_20067);
and UO_1975 (O_1975,N_21323,N_21860);
and UO_1976 (O_1976,N_23538,N_23898);
and UO_1977 (O_1977,N_20521,N_20410);
nor UO_1978 (O_1978,N_21995,N_23541);
xor UO_1979 (O_1979,N_24208,N_20562);
xor UO_1980 (O_1980,N_24782,N_24714);
nand UO_1981 (O_1981,N_21715,N_21699);
nand UO_1982 (O_1982,N_21481,N_21300);
nor UO_1983 (O_1983,N_21716,N_21243);
and UO_1984 (O_1984,N_22850,N_22167);
or UO_1985 (O_1985,N_23656,N_21067);
nand UO_1986 (O_1986,N_23559,N_24889);
nand UO_1987 (O_1987,N_22377,N_22648);
and UO_1988 (O_1988,N_21988,N_23031);
nor UO_1989 (O_1989,N_24053,N_23151);
xnor UO_1990 (O_1990,N_23522,N_21754);
xor UO_1991 (O_1991,N_22934,N_21310);
and UO_1992 (O_1992,N_22418,N_23324);
or UO_1993 (O_1993,N_23678,N_20734);
xnor UO_1994 (O_1994,N_24454,N_23372);
or UO_1995 (O_1995,N_20355,N_20883);
nand UO_1996 (O_1996,N_22972,N_24941);
nor UO_1997 (O_1997,N_23882,N_24934);
or UO_1998 (O_1998,N_21670,N_20852);
nor UO_1999 (O_1999,N_20274,N_20528);
nor UO_2000 (O_2000,N_24728,N_24750);
or UO_2001 (O_2001,N_20889,N_24437);
xnor UO_2002 (O_2002,N_20797,N_21187);
nor UO_2003 (O_2003,N_24222,N_22939);
nor UO_2004 (O_2004,N_21483,N_24764);
xnor UO_2005 (O_2005,N_20937,N_20346);
and UO_2006 (O_2006,N_23317,N_22534);
or UO_2007 (O_2007,N_24100,N_22000);
or UO_2008 (O_2008,N_22918,N_21450);
nor UO_2009 (O_2009,N_24819,N_23897);
xnor UO_2010 (O_2010,N_23835,N_23401);
nand UO_2011 (O_2011,N_23790,N_22462);
or UO_2012 (O_2012,N_21807,N_23972);
xnor UO_2013 (O_2013,N_24088,N_23499);
nor UO_2014 (O_2014,N_23240,N_20064);
xor UO_2015 (O_2015,N_20956,N_22858);
or UO_2016 (O_2016,N_24084,N_24039);
or UO_2017 (O_2017,N_23868,N_21961);
and UO_2018 (O_2018,N_21919,N_21788);
xnor UO_2019 (O_2019,N_24946,N_24231);
xor UO_2020 (O_2020,N_22118,N_20818);
or UO_2021 (O_2021,N_22690,N_21327);
nor UO_2022 (O_2022,N_22486,N_24779);
nor UO_2023 (O_2023,N_22528,N_24958);
nor UO_2024 (O_2024,N_20466,N_20479);
xor UO_2025 (O_2025,N_24368,N_23182);
and UO_2026 (O_2026,N_24330,N_20051);
xnor UO_2027 (O_2027,N_20364,N_23890);
xnor UO_2028 (O_2028,N_20119,N_24886);
or UO_2029 (O_2029,N_22012,N_21094);
nand UO_2030 (O_2030,N_20703,N_21236);
and UO_2031 (O_2031,N_22008,N_20059);
or UO_2032 (O_2032,N_23456,N_22957);
xnor UO_2033 (O_2033,N_22616,N_20685);
or UO_2034 (O_2034,N_21709,N_20159);
or UO_2035 (O_2035,N_23873,N_22583);
nor UO_2036 (O_2036,N_23509,N_21445);
nand UO_2037 (O_2037,N_22523,N_24341);
nor UO_2038 (O_2038,N_21572,N_24386);
nand UO_2039 (O_2039,N_24460,N_20750);
xor UO_2040 (O_2040,N_21543,N_24189);
nor UO_2041 (O_2041,N_23839,N_21987);
nor UO_2042 (O_2042,N_22005,N_20056);
xor UO_2043 (O_2043,N_22110,N_24284);
xor UO_2044 (O_2044,N_22964,N_22166);
nor UO_2045 (O_2045,N_20718,N_21503);
xor UO_2046 (O_2046,N_20254,N_22015);
nand UO_2047 (O_2047,N_21342,N_21734);
and UO_2048 (O_2048,N_24817,N_23729);
or UO_2049 (O_2049,N_23847,N_23042);
or UO_2050 (O_2050,N_23216,N_20172);
and UO_2051 (O_2051,N_22998,N_22769);
or UO_2052 (O_2052,N_21633,N_21593);
xor UO_2053 (O_2053,N_20475,N_24871);
or UO_2054 (O_2054,N_21356,N_22297);
and UO_2055 (O_2055,N_23517,N_24126);
nand UO_2056 (O_2056,N_23056,N_22788);
and UO_2057 (O_2057,N_21460,N_24438);
nor UO_2058 (O_2058,N_24305,N_22572);
nor UO_2059 (O_2059,N_20146,N_24911);
nor UO_2060 (O_2060,N_24545,N_20772);
or UO_2061 (O_2061,N_22433,N_23802);
nand UO_2062 (O_2062,N_20615,N_22079);
xor UO_2063 (O_2063,N_23915,N_24555);
xnor UO_2064 (O_2064,N_24444,N_22651);
nor UO_2065 (O_2065,N_23266,N_21333);
or UO_2066 (O_2066,N_24075,N_23558);
and UO_2067 (O_2067,N_24761,N_24176);
and UO_2068 (O_2068,N_24885,N_22698);
nor UO_2069 (O_2069,N_20514,N_22158);
or UO_2070 (O_2070,N_22210,N_21992);
or UO_2071 (O_2071,N_23063,N_23241);
and UO_2072 (O_2072,N_23325,N_20811);
nand UO_2073 (O_2073,N_21244,N_20383);
and UO_2074 (O_2074,N_20330,N_21848);
and UO_2075 (O_2075,N_24168,N_24414);
and UO_2076 (O_2076,N_24342,N_24868);
nand UO_2077 (O_2077,N_22428,N_24849);
xnor UO_2078 (O_2078,N_21610,N_24396);
and UO_2079 (O_2079,N_23378,N_22867);
nand UO_2080 (O_2080,N_21368,N_21369);
or UO_2081 (O_2081,N_20006,N_24373);
or UO_2082 (O_2082,N_23629,N_21661);
nand UO_2083 (O_2083,N_24300,N_20405);
and UO_2084 (O_2084,N_24567,N_22067);
xnor UO_2085 (O_2085,N_21359,N_23886);
nor UO_2086 (O_2086,N_24695,N_20030);
and UO_2087 (O_2087,N_20495,N_23664);
nor UO_2088 (O_2088,N_23550,N_21320);
nor UO_2089 (O_2089,N_20725,N_23066);
and UO_2090 (O_2090,N_24288,N_24938);
xnor UO_2091 (O_2091,N_20720,N_22390);
nand UO_2092 (O_2092,N_22706,N_24420);
xor UO_2093 (O_2093,N_24439,N_23804);
nand UO_2094 (O_2094,N_23757,N_23009);
nor UO_2095 (O_2095,N_22828,N_24926);
and UO_2096 (O_2096,N_24676,N_22029);
and UO_2097 (O_2097,N_23920,N_20850);
nor UO_2098 (O_2098,N_23347,N_24638);
nand UO_2099 (O_2099,N_23020,N_22056);
xor UO_2100 (O_2100,N_24844,N_20324);
nor UO_2101 (O_2101,N_21396,N_21738);
nor UO_2102 (O_2102,N_24148,N_22959);
xnor UO_2103 (O_2103,N_23367,N_24577);
and UO_2104 (O_2104,N_21222,N_20136);
nor UO_2105 (O_2105,N_24918,N_24155);
or UO_2106 (O_2106,N_22338,N_23963);
nand UO_2107 (O_2107,N_24818,N_23344);
nand UO_2108 (O_2108,N_20109,N_23310);
or UO_2109 (O_2109,N_23065,N_23846);
xor UO_2110 (O_2110,N_20245,N_20485);
xor UO_2111 (O_2111,N_22567,N_23858);
nor UO_2112 (O_2112,N_23196,N_20834);
xnor UO_2113 (O_2113,N_20579,N_21589);
or UO_2114 (O_2114,N_21626,N_22823);
nor UO_2115 (O_2115,N_21410,N_21674);
nor UO_2116 (O_2116,N_24509,N_23595);
xor UO_2117 (O_2117,N_22752,N_22146);
xnor UO_2118 (O_2118,N_20465,N_24560);
nor UO_2119 (O_2119,N_22873,N_20666);
or UO_2120 (O_2120,N_20351,N_24528);
xnor UO_2121 (O_2121,N_23072,N_22599);
and UO_2122 (O_2122,N_23696,N_23715);
nand UO_2123 (O_2123,N_22344,N_24618);
nor UO_2124 (O_2124,N_21311,N_22573);
or UO_2125 (O_2125,N_24290,N_20588);
or UO_2126 (O_2126,N_22267,N_20467);
nand UO_2127 (O_2127,N_21786,N_21500);
or UO_2128 (O_2128,N_20507,N_22037);
nor UO_2129 (O_2129,N_23315,N_22400);
and UO_2130 (O_2130,N_21420,N_22923);
and UO_2131 (O_2131,N_23712,N_23861);
xor UO_2132 (O_2132,N_24199,N_22819);
and UO_2133 (O_2133,N_23206,N_24965);
xnor UO_2134 (O_2134,N_23267,N_22135);
and UO_2135 (O_2135,N_21774,N_23219);
and UO_2136 (O_2136,N_22938,N_20558);
nand UO_2137 (O_2137,N_23607,N_21611);
nand UO_2138 (O_2138,N_22006,N_22705);
xor UO_2139 (O_2139,N_20808,N_23893);
and UO_2140 (O_2140,N_20092,N_22707);
and UO_2141 (O_2141,N_24502,N_23693);
nor UO_2142 (O_2142,N_21419,N_24872);
nor UO_2143 (O_2143,N_24601,N_22316);
or UO_2144 (O_2144,N_21768,N_21449);
nor UO_2145 (O_2145,N_23714,N_23068);
and UO_2146 (O_2146,N_22355,N_24311);
nor UO_2147 (O_2147,N_21322,N_24611);
nor UO_2148 (O_2148,N_22825,N_21765);
and UO_2149 (O_2149,N_22105,N_23418);
and UO_2150 (O_2150,N_23462,N_21326);
or UO_2151 (O_2151,N_20099,N_22066);
or UO_2152 (O_2152,N_24755,N_24550);
and UO_2153 (O_2153,N_24593,N_23508);
nor UO_2154 (O_2154,N_23857,N_20830);
nand UO_2155 (O_2155,N_23252,N_20926);
or UO_2156 (O_2156,N_24505,N_24703);
xor UO_2157 (O_2157,N_21168,N_21717);
or UO_2158 (O_2158,N_21061,N_20938);
nand UO_2159 (O_2159,N_21808,N_24573);
nand UO_2160 (O_2160,N_24409,N_21349);
or UO_2161 (O_2161,N_20839,N_23850);
xor UO_2162 (O_2162,N_24421,N_21385);
or UO_2163 (O_2163,N_22720,N_21253);
nor UO_2164 (O_2164,N_21965,N_24808);
nor UO_2165 (O_2165,N_21719,N_22974);
and UO_2166 (O_2166,N_20879,N_20422);
or UO_2167 (O_2167,N_23268,N_22524);
or UO_2168 (O_2168,N_20207,N_20525);
and UO_2169 (O_2169,N_24652,N_23092);
and UO_2170 (O_2170,N_22525,N_21217);
and UO_2171 (O_2171,N_23706,N_23140);
or UO_2172 (O_2172,N_20261,N_24332);
nor UO_2173 (O_2173,N_24051,N_23708);
and UO_2174 (O_2174,N_20557,N_20093);
xnor UO_2175 (O_2175,N_24119,N_22657);
xnor UO_2176 (O_2176,N_20454,N_21787);
or UO_2177 (O_2177,N_21959,N_20659);
nor UO_2178 (O_2178,N_24143,N_23566);
and UO_2179 (O_2179,N_22448,N_22026);
and UO_2180 (O_2180,N_21179,N_22513);
nor UO_2181 (O_2181,N_22044,N_24425);
nand UO_2182 (O_2182,N_22007,N_20019);
and UO_2183 (O_2183,N_23361,N_24540);
and UO_2184 (O_2184,N_21833,N_21229);
nor UO_2185 (O_2185,N_22372,N_21512);
nand UO_2186 (O_2186,N_21815,N_21497);
xor UO_2187 (O_2187,N_20135,N_22261);
and UO_2188 (O_2188,N_24953,N_20707);
nor UO_2189 (O_2189,N_21031,N_24752);
nor UO_2190 (O_2190,N_20605,N_22728);
xor UO_2191 (O_2191,N_21929,N_21866);
nand UO_2192 (O_2192,N_24746,N_22120);
xnor UO_2193 (O_2193,N_22192,N_24893);
and UO_2194 (O_2194,N_22914,N_24549);
nand UO_2195 (O_2195,N_24704,N_23351);
and UO_2196 (O_2196,N_22184,N_21977);
or UO_2197 (O_2197,N_20047,N_23130);
nor UO_2198 (O_2198,N_22284,N_22069);
and UO_2199 (O_2199,N_21409,N_23974);
nor UO_2200 (O_2200,N_24359,N_24877);
and UO_2201 (O_2201,N_21197,N_24967);
nand UO_2202 (O_2202,N_24226,N_24207);
xnor UO_2203 (O_2203,N_21501,N_21507);
or UO_2204 (O_2204,N_24415,N_21946);
and UO_2205 (O_2205,N_22796,N_20682);
nand UO_2206 (O_2206,N_24012,N_22685);
or UO_2207 (O_2207,N_24891,N_20635);
nor UO_2208 (O_2208,N_21288,N_23842);
or UO_2209 (O_2209,N_23163,N_20153);
nor UO_2210 (O_2210,N_21383,N_22446);
or UO_2211 (O_2211,N_23449,N_23521);
and UO_2212 (O_2212,N_20667,N_21640);
nor UO_2213 (O_2213,N_24047,N_24596);
nand UO_2214 (O_2214,N_20061,N_20473);
nand UO_2215 (O_2215,N_20449,N_24466);
nand UO_2216 (O_2216,N_21104,N_24204);
and UO_2217 (O_2217,N_21778,N_24660);
or UO_2218 (O_2218,N_20990,N_22096);
or UO_2219 (O_2219,N_23192,N_24692);
xnor UO_2220 (O_2220,N_21402,N_21077);
xnor UO_2221 (O_2221,N_20427,N_23863);
or UO_2222 (O_2222,N_24436,N_20898);
xor UO_2223 (O_2223,N_22784,N_24419);
nor UO_2224 (O_2224,N_24379,N_22840);
xor UO_2225 (O_2225,N_22395,N_24686);
and UO_2226 (O_2226,N_21273,N_21378);
and UO_2227 (O_2227,N_22782,N_23973);
or UO_2228 (O_2228,N_24613,N_22731);
nor UO_2229 (O_2229,N_21352,N_20197);
xor UO_2230 (O_2230,N_24645,N_20323);
nor UO_2231 (O_2231,N_21551,N_20264);
nand UO_2232 (O_2232,N_21473,N_21745);
and UO_2233 (O_2233,N_24120,N_21233);
xor UO_2234 (O_2234,N_23431,N_24948);
nand UO_2235 (O_2235,N_21069,N_23516);
and UO_2236 (O_2236,N_24336,N_24902);
and UO_2237 (O_2237,N_23442,N_23663);
nor UO_2238 (O_2238,N_24569,N_23273);
and UO_2239 (O_2239,N_21868,N_20328);
or UO_2240 (O_2240,N_20823,N_24094);
or UO_2241 (O_2241,N_23502,N_24071);
nor UO_2242 (O_2242,N_22623,N_24996);
nor UO_2243 (O_2243,N_23959,N_22216);
xnor UO_2244 (O_2244,N_21280,N_22447);
nand UO_2245 (O_2245,N_24785,N_23934);
or UO_2246 (O_2246,N_23447,N_21138);
nand UO_2247 (O_2247,N_20118,N_22547);
xor UO_2248 (O_2248,N_21107,N_21078);
or UO_2249 (O_2249,N_22423,N_22179);
or UO_2250 (O_2250,N_23309,N_22808);
xor UO_2251 (O_2251,N_23993,N_22631);
and UO_2252 (O_2252,N_22485,N_23295);
and UO_2253 (O_2253,N_22723,N_20371);
nor UO_2254 (O_2254,N_21646,N_22738);
and UO_2255 (O_2255,N_21761,N_24471);
and UO_2256 (O_2256,N_21468,N_24113);
nand UO_2257 (O_2257,N_23688,N_21781);
nand UO_2258 (O_2258,N_24862,N_23501);
xnor UO_2259 (O_2259,N_24040,N_20612);
and UO_2260 (O_2260,N_20102,N_22062);
and UO_2261 (O_2261,N_24842,N_21238);
nor UO_2262 (O_2262,N_20448,N_20929);
and UO_2263 (O_2263,N_22242,N_20950);
nand UO_2264 (O_2264,N_21712,N_20656);
or UO_2265 (O_2265,N_20432,N_24635);
xor UO_2266 (O_2266,N_20411,N_24266);
xor UO_2267 (O_2267,N_24103,N_21297);
nand UO_2268 (O_2268,N_24781,N_20843);
xor UO_2269 (O_2269,N_21285,N_24723);
xor UO_2270 (O_2270,N_24815,N_23093);
nand UO_2271 (O_2271,N_21271,N_21047);
nor UO_2272 (O_2272,N_23681,N_20325);
nand UO_2273 (O_2273,N_24066,N_21721);
xnor UO_2274 (O_2274,N_24536,N_20570);
xor UO_2275 (O_2275,N_21002,N_20831);
or UO_2276 (O_2276,N_21426,N_23067);
xor UO_2277 (O_2277,N_21049,N_21172);
nor UO_2278 (O_2278,N_21379,N_20552);
or UO_2279 (O_2279,N_23211,N_21071);
xnor UO_2280 (O_2280,N_20373,N_24389);
nand UO_2281 (O_2281,N_23642,N_21732);
nand UO_2282 (O_2282,N_22153,N_24215);
nand UO_2283 (O_2283,N_21804,N_22095);
nand UO_2284 (O_2284,N_21653,N_22678);
nand UO_2285 (O_2285,N_24795,N_21084);
nor UO_2286 (O_2286,N_20350,N_24309);
and UO_2287 (O_2287,N_22816,N_22632);
or UO_2288 (O_2288,N_23565,N_24800);
xnor UO_2289 (O_2289,N_24306,N_22660);
or UO_2290 (O_2290,N_23098,N_22764);
and UO_2291 (O_2291,N_21454,N_24272);
nor UO_2292 (O_2292,N_22301,N_24786);
xnor UO_2293 (O_2293,N_23605,N_22091);
or UO_2294 (O_2294,N_21928,N_21836);
nand UO_2295 (O_2295,N_24470,N_23679);
nor UO_2296 (O_2296,N_22049,N_21980);
xor UO_2297 (O_2297,N_20160,N_22719);
nand UO_2298 (O_2298,N_22740,N_23203);
nor UO_2299 (O_2299,N_23186,N_20232);
nor UO_2300 (O_2300,N_24685,N_23694);
xnor UO_2301 (O_2301,N_22473,N_23695);
xor UO_2302 (O_2302,N_20312,N_23118);
nand UO_2303 (O_2303,N_23648,N_24172);
or UO_2304 (O_2304,N_22148,N_22785);
nor UO_2305 (O_2305,N_22488,N_24626);
nor UO_2306 (O_2306,N_24955,N_20474);
nor UO_2307 (O_2307,N_24136,N_21666);
nor UO_2308 (O_2308,N_23352,N_22519);
xor UO_2309 (O_2309,N_23885,N_20805);
nand UO_2310 (O_2310,N_21906,N_22960);
and UO_2311 (O_2311,N_23598,N_22089);
xnor UO_2312 (O_2312,N_24158,N_20228);
and UO_2313 (O_2313,N_23105,N_21641);
xnor UO_2314 (O_2314,N_24312,N_24516);
nor UO_2315 (O_2315,N_23089,N_20490);
nor UO_2316 (O_2316,N_21358,N_22732);
nor UO_2317 (O_2317,N_23178,N_22898);
nor UO_2318 (O_2318,N_24150,N_21561);
xor UO_2319 (O_2319,N_23968,N_23719);
xor UO_2320 (O_2320,N_21267,N_21584);
or UO_2321 (O_2321,N_24377,N_22834);
and UO_2322 (O_2322,N_24977,N_23486);
and UO_2323 (O_2323,N_20039,N_21726);
or UO_2324 (O_2324,N_22378,N_20492);
nor UO_2325 (O_2325,N_21592,N_22010);
xnor UO_2326 (O_2326,N_22478,N_22552);
nand UO_2327 (O_2327,N_21542,N_20927);
xor UO_2328 (O_2328,N_23967,N_23441);
xnor UO_2329 (O_2329,N_21909,N_20847);
and UO_2330 (O_2330,N_21553,N_24629);
xnor UO_2331 (O_2331,N_20752,N_24708);
nor UO_2332 (O_2332,N_23749,N_22360);
or UO_2333 (O_2333,N_20356,N_24350);
or UO_2334 (O_2334,N_21724,N_24202);
nand UO_2335 (O_2335,N_24527,N_24897);
and UO_2336 (O_2336,N_22824,N_21492);
nor UO_2337 (O_2337,N_21215,N_23552);
nand UO_2338 (O_2338,N_24455,N_22269);
nand UO_2339 (O_2339,N_23601,N_24537);
nand UO_2340 (O_2340,N_21730,N_21171);
or UO_2341 (O_2341,N_23567,N_22896);
nand UO_2342 (O_2342,N_20196,N_23145);
nand UO_2343 (O_2343,N_23513,N_22382);
xnor UO_2344 (O_2344,N_21933,N_23054);
nand UO_2345 (O_2345,N_21621,N_23820);
nand UO_2346 (O_2346,N_23218,N_23380);
and UO_2347 (O_2347,N_24947,N_23862);
xor UO_2348 (O_2348,N_24975,N_21398);
or UO_2349 (O_2349,N_20484,N_21430);
or UO_2350 (O_2350,N_22726,N_21242);
nor UO_2351 (O_2351,N_24563,N_23304);
or UO_2352 (O_2352,N_22999,N_21111);
xor UO_2353 (O_2353,N_24772,N_24246);
or UO_2354 (O_2354,N_23692,N_24326);
nor UO_2355 (O_2355,N_23191,N_21599);
nor UO_2356 (O_2356,N_21129,N_20541);
and UO_2357 (O_2357,N_22412,N_21475);
and UO_2358 (O_2358,N_24617,N_20178);
and UO_2359 (O_2359,N_21478,N_23407);
and UO_2360 (O_2360,N_22380,N_21198);
or UO_2361 (O_2361,N_20075,N_20665);
nand UO_2362 (O_2362,N_20012,N_20434);
or UO_2363 (O_2363,N_23961,N_24410);
or UO_2364 (O_2364,N_20224,N_23096);
or UO_2365 (O_2365,N_22309,N_20838);
or UO_2366 (O_2366,N_20063,N_20322);
nor UO_2367 (O_2367,N_20998,N_23179);
nor UO_2368 (O_2368,N_21117,N_20005);
or UO_2369 (O_2369,N_21939,N_23379);
nand UO_2370 (O_2370,N_23202,N_21183);
nand UO_2371 (O_2371,N_21307,N_23452);
nand UO_2372 (O_2372,N_20009,N_24367);
or UO_2373 (O_2373,N_22119,N_20457);
and UO_2374 (O_2374,N_21101,N_23201);
nand UO_2375 (O_2375,N_24724,N_21146);
xor UO_2376 (O_2376,N_22927,N_20509);
nand UO_2377 (O_2377,N_20310,N_21942);
or UO_2378 (O_2378,N_23454,N_21494);
xor UO_2379 (O_2379,N_20101,N_23288);
xnor UO_2380 (O_2380,N_24843,N_20233);
xor UO_2381 (O_2381,N_23221,N_23834);
or UO_2382 (O_2382,N_21180,N_23943);
nand UO_2383 (O_2383,N_22739,N_20247);
or UO_2384 (O_2384,N_24234,N_23410);
xor UO_2385 (O_2385,N_23982,N_21891);
nor UO_2386 (O_2386,N_21112,N_24351);
xnor UO_2387 (O_2387,N_21082,N_23332);
nand UO_2388 (O_2388,N_23599,N_22104);
nand UO_2389 (O_2389,N_23792,N_21753);
nor UO_2390 (O_2390,N_21209,N_20433);
or UO_2391 (O_2391,N_23180,N_24197);
and UO_2392 (O_2392,N_20833,N_24973);
xnor UO_2393 (O_2393,N_23016,N_23279);
nand UO_2394 (O_2394,N_21438,N_20872);
or UO_2395 (O_2395,N_24209,N_22160);
or UO_2396 (O_2396,N_22854,N_21820);
and UO_2397 (O_2397,N_23905,N_22279);
and UO_2398 (O_2398,N_23519,N_20921);
nor UO_2399 (O_2399,N_24041,N_20897);
or UO_2400 (O_2400,N_20868,N_22129);
or UO_2401 (O_2401,N_23457,N_22735);
nand UO_2402 (O_2402,N_22176,N_21582);
nand UO_2403 (O_2403,N_20809,N_22679);
xor UO_2404 (O_2404,N_23012,N_24984);
nor UO_2405 (O_2405,N_21040,N_24428);
and UO_2406 (O_2406,N_24165,N_24198);
nor UO_2407 (O_2407,N_21400,N_20781);
xnor UO_2408 (O_2408,N_22603,N_22504);
nor UO_2409 (O_2409,N_23282,N_20529);
or UO_2410 (O_2410,N_21510,N_21103);
nand UO_2411 (O_2411,N_23246,N_24706);
nand UO_2412 (O_2412,N_20700,N_20777);
nand UO_2413 (O_2413,N_24328,N_22545);
nor UO_2414 (O_2414,N_22009,N_24668);
xor UO_2415 (O_2415,N_22531,N_21446);
nand UO_2416 (O_2416,N_22168,N_22928);
xor UO_2417 (O_2417,N_23597,N_23829);
nand UO_2418 (O_2418,N_20076,N_21688);
nand UO_2419 (O_2419,N_24878,N_21508);
xnor UO_2420 (O_2420,N_20979,N_22838);
nand UO_2421 (O_2421,N_24181,N_23906);
or UO_2422 (O_2422,N_22311,N_22126);
nand UO_2423 (O_2423,N_24837,N_21563);
and UO_2424 (O_2424,N_22114,N_23784);
xor UO_2425 (O_2425,N_24259,N_23549);
nand UO_2426 (O_2426,N_20210,N_23683);
and UO_2427 (O_2427,N_23979,N_23364);
xnor UO_2428 (O_2428,N_21382,N_21757);
xnor UO_2429 (O_2429,N_23727,N_24315);
nand UO_2430 (O_2430,N_22348,N_22082);
and UO_2431 (O_2431,N_20430,N_20191);
nand UO_2432 (O_2432,N_22575,N_20993);
or UO_2433 (O_2433,N_23736,N_23131);
xor UO_2434 (O_2434,N_23008,N_23425);
nor UO_2435 (O_2435,N_21353,N_20168);
xor UO_2436 (O_2436,N_23765,N_24456);
and UO_2437 (O_2437,N_23188,N_24064);
or UO_2438 (O_2438,N_23450,N_22809);
and UO_2439 (O_2439,N_21388,N_24845);
nor UO_2440 (O_2440,N_24441,N_20403);
nor UO_2441 (O_2441,N_20923,N_21108);
nor UO_2442 (O_2442,N_23207,N_23026);
and UO_2443 (O_2443,N_21892,N_22431);
xor UO_2444 (O_2444,N_21912,N_23515);
xnor UO_2445 (O_2445,N_22636,N_23329);
xnor UO_2446 (O_2446,N_20121,N_20648);
xnor UO_2447 (O_2447,N_20827,N_23852);
and UO_2448 (O_2448,N_20571,N_22582);
xnor UO_2449 (O_2449,N_24448,N_20600);
nor UO_2450 (O_2450,N_23081,N_20103);
and UO_2451 (O_2451,N_20024,N_23666);
and UO_2452 (O_2452,N_21932,N_21062);
or UO_2453 (O_2453,N_22831,N_23881);
nand UO_2454 (O_2454,N_20583,N_20556);
nand UO_2455 (O_2455,N_24395,N_20957);
nor UO_2456 (O_2456,N_22866,N_21058);
nand UO_2457 (O_2457,N_20668,N_22122);
xnor UO_2458 (O_2458,N_20533,N_22275);
xor UO_2459 (O_2459,N_23896,N_24498);
nand UO_2460 (O_2460,N_21228,N_23071);
xor UO_2461 (O_2461,N_24650,N_21055);
or UO_2462 (O_2462,N_22997,N_22704);
xnor UO_2463 (O_2463,N_20803,N_21490);
xnor UO_2464 (O_2464,N_22550,N_21169);
nor UO_2465 (O_2465,N_24899,N_22392);
or UO_2466 (O_2466,N_24925,N_22975);
and UO_2467 (O_2467,N_21779,N_22251);
nor UO_2468 (O_2468,N_20922,N_23987);
or UO_2469 (O_2469,N_23824,N_23713);
xor UO_2470 (O_2470,N_24589,N_23584);
and UO_2471 (O_2471,N_24125,N_22233);
nor UO_2472 (O_2472,N_24497,N_23610);
nor UO_2473 (O_2473,N_21199,N_24427);
nor UO_2474 (O_2474,N_24543,N_23744);
and UO_2475 (O_2475,N_23743,N_23259);
xor UO_2476 (O_2476,N_22515,N_21843);
nand UO_2477 (O_2477,N_21588,N_22144);
and UO_2478 (O_2478,N_24400,N_20078);
nand UO_2479 (O_2479,N_20391,N_23977);
or UO_2480 (O_2480,N_23322,N_24857);
xor UO_2481 (O_2481,N_22098,N_20747);
or UO_2482 (O_2482,N_21579,N_23444);
xnor UO_2483 (O_2483,N_24705,N_20658);
and UO_2484 (O_2484,N_23921,N_22266);
or UO_2485 (O_2485,N_21043,N_23586);
or UO_2486 (O_2486,N_20171,N_20891);
or UO_2487 (O_2487,N_21770,N_20858);
xor UO_2488 (O_2488,N_20214,N_21889);
nor UO_2489 (O_2489,N_22299,N_20292);
nor UO_2490 (O_2490,N_22795,N_24775);
and UO_2491 (O_2491,N_21898,N_24711);
and UO_2492 (O_2492,N_24932,N_24059);
xnor UO_2493 (O_2493,N_22692,N_20353);
and UO_2494 (O_2494,N_21227,N_21004);
nor UO_2495 (O_2495,N_20962,N_24187);
or UO_2496 (O_2496,N_23531,N_23053);
nand UO_2497 (O_2497,N_24853,N_21746);
or UO_2498 (O_2498,N_22536,N_20799);
nand UO_2499 (O_2499,N_21467,N_22820);
nand UO_2500 (O_2500,N_20463,N_24884);
or UO_2501 (O_2501,N_21090,N_20317);
and UO_2502 (O_2502,N_23201,N_21102);
nor UO_2503 (O_2503,N_22084,N_21922);
xor UO_2504 (O_2504,N_22808,N_20029);
and UO_2505 (O_2505,N_21421,N_22704);
nand UO_2506 (O_2506,N_23791,N_22831);
xnor UO_2507 (O_2507,N_24695,N_24269);
nand UO_2508 (O_2508,N_21818,N_23464);
xor UO_2509 (O_2509,N_21190,N_24929);
and UO_2510 (O_2510,N_20524,N_24342);
nand UO_2511 (O_2511,N_22554,N_22254);
nor UO_2512 (O_2512,N_22532,N_22625);
xor UO_2513 (O_2513,N_23093,N_21328);
or UO_2514 (O_2514,N_22272,N_22409);
xor UO_2515 (O_2515,N_20977,N_22990);
nor UO_2516 (O_2516,N_21643,N_22747);
xor UO_2517 (O_2517,N_21502,N_24354);
or UO_2518 (O_2518,N_22843,N_22179);
nand UO_2519 (O_2519,N_21927,N_24270);
xor UO_2520 (O_2520,N_21926,N_22655);
nand UO_2521 (O_2521,N_22476,N_20031);
nor UO_2522 (O_2522,N_24973,N_23248);
nand UO_2523 (O_2523,N_24304,N_24390);
nand UO_2524 (O_2524,N_22029,N_23267);
and UO_2525 (O_2525,N_20179,N_22994);
and UO_2526 (O_2526,N_21048,N_24628);
nand UO_2527 (O_2527,N_20837,N_20354);
or UO_2528 (O_2528,N_23260,N_23864);
nor UO_2529 (O_2529,N_20423,N_24153);
xor UO_2530 (O_2530,N_23734,N_21491);
nor UO_2531 (O_2531,N_22374,N_23500);
nand UO_2532 (O_2532,N_20933,N_24233);
and UO_2533 (O_2533,N_22083,N_23777);
xnor UO_2534 (O_2534,N_20617,N_21734);
nor UO_2535 (O_2535,N_22043,N_23803);
or UO_2536 (O_2536,N_20887,N_24587);
nand UO_2537 (O_2537,N_24938,N_20245);
nor UO_2538 (O_2538,N_23848,N_22774);
or UO_2539 (O_2539,N_24198,N_24221);
xor UO_2540 (O_2540,N_24017,N_21428);
nand UO_2541 (O_2541,N_21995,N_23933);
nor UO_2542 (O_2542,N_21173,N_21820);
or UO_2543 (O_2543,N_22004,N_20398);
nor UO_2544 (O_2544,N_23913,N_22758);
and UO_2545 (O_2545,N_21967,N_23421);
nand UO_2546 (O_2546,N_21512,N_24122);
xnor UO_2547 (O_2547,N_23360,N_22212);
xor UO_2548 (O_2548,N_20270,N_24835);
nand UO_2549 (O_2549,N_24872,N_22678);
nand UO_2550 (O_2550,N_23151,N_21471);
or UO_2551 (O_2551,N_22988,N_22742);
nand UO_2552 (O_2552,N_23549,N_21063);
nor UO_2553 (O_2553,N_21001,N_21224);
or UO_2554 (O_2554,N_23652,N_22256);
or UO_2555 (O_2555,N_20604,N_22778);
and UO_2556 (O_2556,N_21640,N_24057);
and UO_2557 (O_2557,N_24631,N_22143);
nor UO_2558 (O_2558,N_23261,N_24355);
xor UO_2559 (O_2559,N_20681,N_20461);
nor UO_2560 (O_2560,N_21812,N_21511);
xnor UO_2561 (O_2561,N_24025,N_20700);
xnor UO_2562 (O_2562,N_20326,N_21649);
nor UO_2563 (O_2563,N_21661,N_20269);
nand UO_2564 (O_2564,N_22596,N_22035);
nor UO_2565 (O_2565,N_21799,N_22996);
or UO_2566 (O_2566,N_20312,N_22345);
xor UO_2567 (O_2567,N_20359,N_22143);
nor UO_2568 (O_2568,N_24421,N_24137);
or UO_2569 (O_2569,N_22534,N_23523);
and UO_2570 (O_2570,N_24072,N_23474);
and UO_2571 (O_2571,N_21710,N_24364);
xor UO_2572 (O_2572,N_20585,N_24435);
nand UO_2573 (O_2573,N_23147,N_24251);
and UO_2574 (O_2574,N_24311,N_20587);
or UO_2575 (O_2575,N_22431,N_24410);
or UO_2576 (O_2576,N_24962,N_22167);
xor UO_2577 (O_2577,N_20013,N_24530);
or UO_2578 (O_2578,N_22778,N_23587);
and UO_2579 (O_2579,N_23593,N_22224);
nand UO_2580 (O_2580,N_20005,N_20185);
xor UO_2581 (O_2581,N_20042,N_21556);
and UO_2582 (O_2582,N_20177,N_23637);
xnor UO_2583 (O_2583,N_24725,N_20714);
xnor UO_2584 (O_2584,N_24433,N_22826);
nor UO_2585 (O_2585,N_20749,N_21136);
nor UO_2586 (O_2586,N_21913,N_23221);
xor UO_2587 (O_2587,N_24877,N_24655);
xor UO_2588 (O_2588,N_23638,N_20300);
or UO_2589 (O_2589,N_24181,N_22239);
xnor UO_2590 (O_2590,N_20249,N_24549);
nor UO_2591 (O_2591,N_22673,N_24651);
nand UO_2592 (O_2592,N_23007,N_21334);
or UO_2593 (O_2593,N_21701,N_23843);
nand UO_2594 (O_2594,N_21931,N_22906);
and UO_2595 (O_2595,N_20910,N_23489);
xor UO_2596 (O_2596,N_24043,N_24505);
or UO_2597 (O_2597,N_24719,N_22660);
nor UO_2598 (O_2598,N_20784,N_20781);
nor UO_2599 (O_2599,N_23696,N_20916);
or UO_2600 (O_2600,N_22961,N_22679);
nand UO_2601 (O_2601,N_21065,N_21359);
and UO_2602 (O_2602,N_21234,N_20044);
and UO_2603 (O_2603,N_20567,N_22267);
or UO_2604 (O_2604,N_22085,N_20924);
nor UO_2605 (O_2605,N_22706,N_24952);
or UO_2606 (O_2606,N_23444,N_23424);
nand UO_2607 (O_2607,N_20838,N_22356);
nor UO_2608 (O_2608,N_21892,N_20406);
or UO_2609 (O_2609,N_24577,N_22058);
xor UO_2610 (O_2610,N_20705,N_22100);
nand UO_2611 (O_2611,N_24257,N_20288);
nand UO_2612 (O_2612,N_24582,N_24992);
or UO_2613 (O_2613,N_23376,N_24017);
xnor UO_2614 (O_2614,N_23980,N_23440);
xnor UO_2615 (O_2615,N_20782,N_20142);
nor UO_2616 (O_2616,N_24810,N_20352);
nor UO_2617 (O_2617,N_23991,N_21728);
xor UO_2618 (O_2618,N_20179,N_20187);
nor UO_2619 (O_2619,N_23531,N_20429);
nand UO_2620 (O_2620,N_20642,N_24018);
nand UO_2621 (O_2621,N_21327,N_20597);
or UO_2622 (O_2622,N_22651,N_24423);
or UO_2623 (O_2623,N_21992,N_22252);
or UO_2624 (O_2624,N_21992,N_23122);
nor UO_2625 (O_2625,N_21505,N_22824);
nand UO_2626 (O_2626,N_20747,N_20539);
nor UO_2627 (O_2627,N_24130,N_23689);
and UO_2628 (O_2628,N_21521,N_21191);
nor UO_2629 (O_2629,N_20234,N_21993);
xor UO_2630 (O_2630,N_24801,N_24266);
nand UO_2631 (O_2631,N_21105,N_20447);
nand UO_2632 (O_2632,N_24087,N_20861);
xor UO_2633 (O_2633,N_20344,N_21228);
nand UO_2634 (O_2634,N_23831,N_20803);
or UO_2635 (O_2635,N_20877,N_20547);
nor UO_2636 (O_2636,N_22478,N_22124);
xor UO_2637 (O_2637,N_21312,N_20149);
xor UO_2638 (O_2638,N_23181,N_23737);
or UO_2639 (O_2639,N_23782,N_22298);
nor UO_2640 (O_2640,N_20098,N_24135);
or UO_2641 (O_2641,N_20469,N_20062);
xnor UO_2642 (O_2642,N_22931,N_23977);
xnor UO_2643 (O_2643,N_24600,N_24711);
nand UO_2644 (O_2644,N_22136,N_23884);
or UO_2645 (O_2645,N_24775,N_23012);
or UO_2646 (O_2646,N_24388,N_24462);
and UO_2647 (O_2647,N_21956,N_21463);
xor UO_2648 (O_2648,N_24902,N_21606);
nor UO_2649 (O_2649,N_20058,N_22431);
or UO_2650 (O_2650,N_22810,N_21072);
nand UO_2651 (O_2651,N_24062,N_22105);
or UO_2652 (O_2652,N_20901,N_20827);
nand UO_2653 (O_2653,N_22864,N_22268);
nand UO_2654 (O_2654,N_20713,N_22514);
or UO_2655 (O_2655,N_23476,N_23023);
or UO_2656 (O_2656,N_21913,N_22502);
nand UO_2657 (O_2657,N_22270,N_23853);
nor UO_2658 (O_2658,N_20878,N_21042);
nor UO_2659 (O_2659,N_22341,N_22419);
nor UO_2660 (O_2660,N_20024,N_22331);
nor UO_2661 (O_2661,N_20806,N_20538);
or UO_2662 (O_2662,N_23021,N_23209);
xnor UO_2663 (O_2663,N_20669,N_22792);
nand UO_2664 (O_2664,N_23366,N_20196);
nor UO_2665 (O_2665,N_21915,N_22584);
or UO_2666 (O_2666,N_24790,N_22852);
nand UO_2667 (O_2667,N_21715,N_24151);
or UO_2668 (O_2668,N_20608,N_20179);
xnor UO_2669 (O_2669,N_24961,N_21250);
and UO_2670 (O_2670,N_24093,N_21240);
and UO_2671 (O_2671,N_21144,N_22399);
xnor UO_2672 (O_2672,N_24211,N_21829);
xnor UO_2673 (O_2673,N_22201,N_22192);
and UO_2674 (O_2674,N_23538,N_21623);
xnor UO_2675 (O_2675,N_24287,N_21272);
nand UO_2676 (O_2676,N_22049,N_23899);
or UO_2677 (O_2677,N_23306,N_20408);
and UO_2678 (O_2678,N_20895,N_21657);
or UO_2679 (O_2679,N_22546,N_21631);
xor UO_2680 (O_2680,N_21752,N_24440);
nor UO_2681 (O_2681,N_23345,N_21197);
or UO_2682 (O_2682,N_21816,N_24151);
nand UO_2683 (O_2683,N_20269,N_23996);
xor UO_2684 (O_2684,N_23252,N_21609);
xnor UO_2685 (O_2685,N_21129,N_23773);
or UO_2686 (O_2686,N_23482,N_21200);
xnor UO_2687 (O_2687,N_22531,N_22359);
nand UO_2688 (O_2688,N_23482,N_22190);
and UO_2689 (O_2689,N_20012,N_24912);
xnor UO_2690 (O_2690,N_22029,N_23298);
nand UO_2691 (O_2691,N_23638,N_20604);
and UO_2692 (O_2692,N_21257,N_20710);
and UO_2693 (O_2693,N_23820,N_22849);
nand UO_2694 (O_2694,N_24034,N_23692);
xor UO_2695 (O_2695,N_20142,N_20733);
nand UO_2696 (O_2696,N_23291,N_24884);
and UO_2697 (O_2697,N_21797,N_22339);
nand UO_2698 (O_2698,N_22063,N_21482);
or UO_2699 (O_2699,N_24409,N_23463);
nand UO_2700 (O_2700,N_21441,N_21277);
nand UO_2701 (O_2701,N_24849,N_23233);
nand UO_2702 (O_2702,N_23815,N_21230);
or UO_2703 (O_2703,N_21390,N_22863);
nand UO_2704 (O_2704,N_20454,N_22548);
nor UO_2705 (O_2705,N_24014,N_20966);
nor UO_2706 (O_2706,N_20299,N_24823);
and UO_2707 (O_2707,N_21138,N_24903);
or UO_2708 (O_2708,N_22209,N_24166);
xor UO_2709 (O_2709,N_22532,N_20029);
nor UO_2710 (O_2710,N_20130,N_22795);
xor UO_2711 (O_2711,N_22512,N_22352);
xor UO_2712 (O_2712,N_21945,N_21476);
and UO_2713 (O_2713,N_23294,N_23793);
nand UO_2714 (O_2714,N_20549,N_23881);
and UO_2715 (O_2715,N_21984,N_20396);
or UO_2716 (O_2716,N_24461,N_23861);
and UO_2717 (O_2717,N_21669,N_23273);
or UO_2718 (O_2718,N_24208,N_20593);
nor UO_2719 (O_2719,N_22910,N_20381);
xor UO_2720 (O_2720,N_21804,N_23338);
or UO_2721 (O_2721,N_23315,N_21100);
and UO_2722 (O_2722,N_20413,N_22560);
and UO_2723 (O_2723,N_24173,N_20636);
or UO_2724 (O_2724,N_21166,N_23857);
or UO_2725 (O_2725,N_20676,N_22880);
and UO_2726 (O_2726,N_22292,N_22037);
nand UO_2727 (O_2727,N_20595,N_22223);
and UO_2728 (O_2728,N_20536,N_21929);
or UO_2729 (O_2729,N_24201,N_20948);
or UO_2730 (O_2730,N_24530,N_20963);
xor UO_2731 (O_2731,N_24828,N_24817);
and UO_2732 (O_2732,N_21741,N_21924);
xnor UO_2733 (O_2733,N_20406,N_21445);
nor UO_2734 (O_2734,N_23803,N_24834);
and UO_2735 (O_2735,N_20441,N_22544);
nor UO_2736 (O_2736,N_24058,N_23175);
nor UO_2737 (O_2737,N_21523,N_20318);
or UO_2738 (O_2738,N_22812,N_21261);
nand UO_2739 (O_2739,N_24103,N_21300);
or UO_2740 (O_2740,N_22422,N_23128);
or UO_2741 (O_2741,N_24493,N_23431);
nor UO_2742 (O_2742,N_20782,N_24423);
or UO_2743 (O_2743,N_20282,N_22358);
nor UO_2744 (O_2744,N_21005,N_22226);
and UO_2745 (O_2745,N_24426,N_24468);
and UO_2746 (O_2746,N_20264,N_23437);
xor UO_2747 (O_2747,N_22469,N_23129);
nand UO_2748 (O_2748,N_23368,N_23638);
xor UO_2749 (O_2749,N_20842,N_22920);
or UO_2750 (O_2750,N_22598,N_20729);
xor UO_2751 (O_2751,N_21600,N_22949);
or UO_2752 (O_2752,N_20477,N_20104);
xnor UO_2753 (O_2753,N_23778,N_22560);
or UO_2754 (O_2754,N_24024,N_24300);
nand UO_2755 (O_2755,N_22600,N_20275);
nand UO_2756 (O_2756,N_20258,N_21755);
nand UO_2757 (O_2757,N_22776,N_24657);
and UO_2758 (O_2758,N_20656,N_24347);
xnor UO_2759 (O_2759,N_23188,N_21547);
nor UO_2760 (O_2760,N_22650,N_20089);
xor UO_2761 (O_2761,N_21940,N_23796);
and UO_2762 (O_2762,N_22299,N_23199);
and UO_2763 (O_2763,N_21169,N_23667);
nand UO_2764 (O_2764,N_24788,N_21840);
nand UO_2765 (O_2765,N_22056,N_20560);
nand UO_2766 (O_2766,N_23604,N_24838);
nand UO_2767 (O_2767,N_21027,N_23151);
or UO_2768 (O_2768,N_22184,N_20720);
and UO_2769 (O_2769,N_24457,N_23347);
nor UO_2770 (O_2770,N_20891,N_21446);
nand UO_2771 (O_2771,N_22878,N_22503);
xnor UO_2772 (O_2772,N_20980,N_23843);
nor UO_2773 (O_2773,N_21483,N_20448);
nor UO_2774 (O_2774,N_23747,N_24202);
and UO_2775 (O_2775,N_22822,N_21218);
nor UO_2776 (O_2776,N_22453,N_21917);
and UO_2777 (O_2777,N_24138,N_21597);
nand UO_2778 (O_2778,N_20898,N_23458);
xnor UO_2779 (O_2779,N_24086,N_24690);
nand UO_2780 (O_2780,N_22568,N_21849);
or UO_2781 (O_2781,N_23649,N_24934);
nor UO_2782 (O_2782,N_24618,N_21609);
nor UO_2783 (O_2783,N_24044,N_21385);
xnor UO_2784 (O_2784,N_24158,N_23513);
nor UO_2785 (O_2785,N_21021,N_23458);
and UO_2786 (O_2786,N_23982,N_22763);
nand UO_2787 (O_2787,N_21958,N_20278);
nor UO_2788 (O_2788,N_21684,N_24976);
and UO_2789 (O_2789,N_22446,N_21956);
nand UO_2790 (O_2790,N_22866,N_21646);
xor UO_2791 (O_2791,N_22512,N_21122);
nand UO_2792 (O_2792,N_21692,N_22272);
nor UO_2793 (O_2793,N_20705,N_20892);
nor UO_2794 (O_2794,N_22468,N_23267);
or UO_2795 (O_2795,N_22150,N_24872);
nand UO_2796 (O_2796,N_20907,N_20614);
and UO_2797 (O_2797,N_20232,N_20020);
nor UO_2798 (O_2798,N_20855,N_21810);
xnor UO_2799 (O_2799,N_24543,N_21578);
xnor UO_2800 (O_2800,N_24568,N_20160);
and UO_2801 (O_2801,N_22604,N_23807);
nand UO_2802 (O_2802,N_20357,N_23889);
xor UO_2803 (O_2803,N_22198,N_24305);
or UO_2804 (O_2804,N_23838,N_21146);
and UO_2805 (O_2805,N_24519,N_24236);
nand UO_2806 (O_2806,N_20435,N_21116);
nor UO_2807 (O_2807,N_23421,N_22683);
and UO_2808 (O_2808,N_21795,N_22635);
and UO_2809 (O_2809,N_24100,N_20615);
xor UO_2810 (O_2810,N_21307,N_20228);
and UO_2811 (O_2811,N_24005,N_21526);
and UO_2812 (O_2812,N_22565,N_24704);
or UO_2813 (O_2813,N_24785,N_22740);
and UO_2814 (O_2814,N_22036,N_22254);
nor UO_2815 (O_2815,N_23014,N_24548);
nor UO_2816 (O_2816,N_21422,N_21759);
nor UO_2817 (O_2817,N_22922,N_24084);
xor UO_2818 (O_2818,N_21664,N_21336);
or UO_2819 (O_2819,N_24211,N_24845);
xnor UO_2820 (O_2820,N_21812,N_22401);
and UO_2821 (O_2821,N_20126,N_22492);
nor UO_2822 (O_2822,N_23034,N_22354);
xnor UO_2823 (O_2823,N_21177,N_22252);
or UO_2824 (O_2824,N_23884,N_21469);
or UO_2825 (O_2825,N_21790,N_24611);
nor UO_2826 (O_2826,N_24370,N_20138);
nor UO_2827 (O_2827,N_23149,N_23773);
and UO_2828 (O_2828,N_24420,N_21777);
xor UO_2829 (O_2829,N_22401,N_24172);
or UO_2830 (O_2830,N_20151,N_23325);
nor UO_2831 (O_2831,N_24733,N_22665);
nor UO_2832 (O_2832,N_21604,N_24338);
or UO_2833 (O_2833,N_23939,N_24099);
and UO_2834 (O_2834,N_20122,N_24469);
nand UO_2835 (O_2835,N_21246,N_21410);
nor UO_2836 (O_2836,N_24692,N_24017);
xnor UO_2837 (O_2837,N_22594,N_20040);
xor UO_2838 (O_2838,N_20360,N_21060);
or UO_2839 (O_2839,N_21501,N_24776);
nand UO_2840 (O_2840,N_21941,N_20543);
or UO_2841 (O_2841,N_21445,N_21998);
or UO_2842 (O_2842,N_23740,N_22443);
xor UO_2843 (O_2843,N_22557,N_24799);
or UO_2844 (O_2844,N_22712,N_24759);
and UO_2845 (O_2845,N_23550,N_23205);
or UO_2846 (O_2846,N_24185,N_22128);
xor UO_2847 (O_2847,N_22681,N_24112);
or UO_2848 (O_2848,N_20380,N_20246);
nand UO_2849 (O_2849,N_22202,N_21459);
or UO_2850 (O_2850,N_21298,N_24542);
and UO_2851 (O_2851,N_24668,N_22947);
xor UO_2852 (O_2852,N_22676,N_24128);
nor UO_2853 (O_2853,N_22346,N_21515);
and UO_2854 (O_2854,N_23586,N_21686);
xor UO_2855 (O_2855,N_23259,N_22760);
and UO_2856 (O_2856,N_24046,N_24300);
nand UO_2857 (O_2857,N_24009,N_22203);
or UO_2858 (O_2858,N_23027,N_20080);
nor UO_2859 (O_2859,N_21044,N_24843);
or UO_2860 (O_2860,N_22228,N_24336);
or UO_2861 (O_2861,N_21088,N_23495);
and UO_2862 (O_2862,N_21063,N_20271);
or UO_2863 (O_2863,N_20027,N_21340);
or UO_2864 (O_2864,N_20086,N_22418);
nor UO_2865 (O_2865,N_22502,N_24567);
nor UO_2866 (O_2866,N_22304,N_21521);
nand UO_2867 (O_2867,N_24248,N_23325);
nand UO_2868 (O_2868,N_23657,N_20893);
xnor UO_2869 (O_2869,N_22243,N_22371);
or UO_2870 (O_2870,N_23369,N_24158);
nand UO_2871 (O_2871,N_21304,N_22525);
xnor UO_2872 (O_2872,N_24746,N_23778);
nor UO_2873 (O_2873,N_23879,N_24215);
nand UO_2874 (O_2874,N_23735,N_22116);
or UO_2875 (O_2875,N_20009,N_20164);
nand UO_2876 (O_2876,N_23987,N_24335);
or UO_2877 (O_2877,N_20673,N_24782);
xor UO_2878 (O_2878,N_23318,N_20949);
nand UO_2879 (O_2879,N_24119,N_22047);
nand UO_2880 (O_2880,N_22850,N_20091);
or UO_2881 (O_2881,N_20667,N_21249);
nor UO_2882 (O_2882,N_20072,N_21548);
or UO_2883 (O_2883,N_20749,N_23284);
nor UO_2884 (O_2884,N_21964,N_20345);
nand UO_2885 (O_2885,N_20068,N_22309);
nor UO_2886 (O_2886,N_24417,N_23802);
nand UO_2887 (O_2887,N_23274,N_20366);
or UO_2888 (O_2888,N_22316,N_21847);
nand UO_2889 (O_2889,N_23844,N_23865);
nor UO_2890 (O_2890,N_23077,N_20250);
xnor UO_2891 (O_2891,N_24142,N_24230);
nand UO_2892 (O_2892,N_23396,N_24064);
xnor UO_2893 (O_2893,N_20972,N_23584);
nor UO_2894 (O_2894,N_22306,N_24830);
nand UO_2895 (O_2895,N_20772,N_24860);
and UO_2896 (O_2896,N_24136,N_22579);
nor UO_2897 (O_2897,N_21596,N_21391);
nor UO_2898 (O_2898,N_24570,N_24314);
nor UO_2899 (O_2899,N_20224,N_21186);
xnor UO_2900 (O_2900,N_20473,N_20245);
nor UO_2901 (O_2901,N_20399,N_22551);
xnor UO_2902 (O_2902,N_22288,N_24091);
nor UO_2903 (O_2903,N_23231,N_23281);
or UO_2904 (O_2904,N_22040,N_23537);
nor UO_2905 (O_2905,N_22273,N_23005);
nor UO_2906 (O_2906,N_24476,N_20667);
or UO_2907 (O_2907,N_23051,N_24026);
nand UO_2908 (O_2908,N_22025,N_21130);
nand UO_2909 (O_2909,N_21604,N_21475);
xor UO_2910 (O_2910,N_20201,N_23868);
nand UO_2911 (O_2911,N_24853,N_21866);
nand UO_2912 (O_2912,N_20519,N_23117);
nand UO_2913 (O_2913,N_22444,N_23041);
xnor UO_2914 (O_2914,N_24749,N_21518);
nor UO_2915 (O_2915,N_22026,N_20724);
and UO_2916 (O_2916,N_22274,N_22071);
nor UO_2917 (O_2917,N_20588,N_22116);
nand UO_2918 (O_2918,N_21390,N_23357);
and UO_2919 (O_2919,N_20686,N_22934);
and UO_2920 (O_2920,N_23555,N_23736);
xnor UO_2921 (O_2921,N_20332,N_21710);
and UO_2922 (O_2922,N_24987,N_22880);
xor UO_2923 (O_2923,N_21242,N_23954);
and UO_2924 (O_2924,N_21101,N_20210);
xor UO_2925 (O_2925,N_21192,N_23331);
or UO_2926 (O_2926,N_22818,N_23850);
nor UO_2927 (O_2927,N_24559,N_20307);
xor UO_2928 (O_2928,N_21511,N_23370);
or UO_2929 (O_2929,N_23273,N_20805);
or UO_2930 (O_2930,N_22164,N_21328);
and UO_2931 (O_2931,N_22445,N_21803);
nand UO_2932 (O_2932,N_22222,N_22812);
xor UO_2933 (O_2933,N_22435,N_24308);
xnor UO_2934 (O_2934,N_22381,N_20100);
xor UO_2935 (O_2935,N_23512,N_21242);
nand UO_2936 (O_2936,N_23637,N_24659);
xor UO_2937 (O_2937,N_20491,N_21925);
xnor UO_2938 (O_2938,N_20526,N_24474);
and UO_2939 (O_2939,N_22259,N_23177);
or UO_2940 (O_2940,N_21894,N_22380);
xnor UO_2941 (O_2941,N_23407,N_24054);
and UO_2942 (O_2942,N_20281,N_20153);
xor UO_2943 (O_2943,N_20294,N_20083);
and UO_2944 (O_2944,N_21858,N_23955);
and UO_2945 (O_2945,N_22508,N_21221);
or UO_2946 (O_2946,N_22110,N_21501);
and UO_2947 (O_2947,N_20679,N_22306);
and UO_2948 (O_2948,N_24643,N_20977);
xnor UO_2949 (O_2949,N_23670,N_20939);
or UO_2950 (O_2950,N_23917,N_20404);
or UO_2951 (O_2951,N_21375,N_24108);
or UO_2952 (O_2952,N_23036,N_21192);
nor UO_2953 (O_2953,N_21046,N_23044);
nand UO_2954 (O_2954,N_23127,N_23436);
and UO_2955 (O_2955,N_24997,N_20462);
nand UO_2956 (O_2956,N_24519,N_20749);
nor UO_2957 (O_2957,N_24775,N_23484);
or UO_2958 (O_2958,N_23177,N_20346);
or UO_2959 (O_2959,N_24781,N_22501);
nor UO_2960 (O_2960,N_23759,N_21809);
and UO_2961 (O_2961,N_22560,N_22648);
or UO_2962 (O_2962,N_24149,N_20890);
or UO_2963 (O_2963,N_22281,N_20372);
or UO_2964 (O_2964,N_23712,N_23340);
nor UO_2965 (O_2965,N_22693,N_20535);
xnor UO_2966 (O_2966,N_24967,N_23215);
and UO_2967 (O_2967,N_24535,N_22156);
xnor UO_2968 (O_2968,N_22788,N_23379);
nand UO_2969 (O_2969,N_21099,N_20943);
and UO_2970 (O_2970,N_23984,N_24916);
nand UO_2971 (O_2971,N_23017,N_22451);
and UO_2972 (O_2972,N_22694,N_23388);
and UO_2973 (O_2973,N_22319,N_20600);
and UO_2974 (O_2974,N_24809,N_23654);
xor UO_2975 (O_2975,N_24166,N_21105);
xnor UO_2976 (O_2976,N_22873,N_21936);
nor UO_2977 (O_2977,N_23402,N_22723);
and UO_2978 (O_2978,N_21483,N_21424);
nand UO_2979 (O_2979,N_20789,N_21356);
nor UO_2980 (O_2980,N_24329,N_20904);
nand UO_2981 (O_2981,N_20387,N_21846);
nand UO_2982 (O_2982,N_23183,N_22192);
nand UO_2983 (O_2983,N_24505,N_21157);
xnor UO_2984 (O_2984,N_24669,N_22555);
nor UO_2985 (O_2985,N_23474,N_22720);
xnor UO_2986 (O_2986,N_22550,N_21916);
nor UO_2987 (O_2987,N_24336,N_20774);
or UO_2988 (O_2988,N_22093,N_22489);
and UO_2989 (O_2989,N_22039,N_21052);
xor UO_2990 (O_2990,N_21941,N_20796);
xnor UO_2991 (O_2991,N_24055,N_22848);
or UO_2992 (O_2992,N_23901,N_20879);
xor UO_2993 (O_2993,N_24226,N_21386);
nand UO_2994 (O_2994,N_20217,N_24855);
and UO_2995 (O_2995,N_21021,N_20720);
nor UO_2996 (O_2996,N_21213,N_21970);
or UO_2997 (O_2997,N_23791,N_24214);
nand UO_2998 (O_2998,N_22828,N_24650);
and UO_2999 (O_2999,N_20051,N_21841);
endmodule