module basic_500_3000_500_50_levels_1xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_132,In_478);
or U1 (N_1,In_368,In_36);
and U2 (N_2,In_48,In_471);
nand U3 (N_3,In_474,In_339);
or U4 (N_4,In_145,In_21);
nand U5 (N_5,In_114,In_196);
nor U6 (N_6,In_483,In_260);
nand U7 (N_7,In_4,In_460);
or U8 (N_8,In_51,In_288);
and U9 (N_9,In_447,In_61);
nand U10 (N_10,In_23,In_292);
nor U11 (N_11,In_46,In_231);
nand U12 (N_12,In_58,In_286);
nor U13 (N_13,In_420,In_381);
or U14 (N_14,In_446,In_392);
nor U15 (N_15,In_477,In_246);
and U16 (N_16,In_52,In_130);
and U17 (N_17,In_80,In_302);
nand U18 (N_18,In_82,In_230);
or U19 (N_19,In_265,In_121);
or U20 (N_20,In_140,In_393);
or U21 (N_21,In_15,In_306);
and U22 (N_22,In_427,In_489);
nand U23 (N_23,In_285,In_225);
nor U24 (N_24,In_150,In_300);
nor U25 (N_25,In_390,In_401);
nor U26 (N_26,In_104,In_139);
and U27 (N_27,In_45,In_269);
xnor U28 (N_28,In_487,In_350);
nand U29 (N_29,In_181,In_55);
or U30 (N_30,In_463,In_490);
nand U31 (N_31,In_253,In_450);
nor U32 (N_32,In_404,In_206);
or U33 (N_33,In_14,In_195);
xor U34 (N_34,In_391,In_372);
nand U35 (N_35,In_448,In_492);
and U36 (N_36,In_12,In_256);
nor U37 (N_37,In_277,In_374);
and U38 (N_38,In_220,In_214);
nor U39 (N_39,In_77,In_408);
nand U40 (N_40,In_428,In_112);
nor U41 (N_41,In_356,In_464);
and U42 (N_42,In_168,In_326);
nor U43 (N_43,In_74,In_352);
nand U44 (N_44,In_63,In_67);
nor U45 (N_45,In_336,In_396);
nand U46 (N_46,In_353,In_304);
or U47 (N_47,In_432,In_403);
or U48 (N_48,In_482,In_346);
or U49 (N_49,In_355,In_362);
nand U50 (N_50,In_19,In_60);
nor U51 (N_51,In_115,In_197);
and U52 (N_52,In_186,In_238);
and U53 (N_53,In_227,In_129);
nand U54 (N_54,In_81,In_125);
and U55 (N_55,In_154,In_223);
or U56 (N_56,In_496,In_436);
or U57 (N_57,In_272,In_117);
nand U58 (N_58,In_116,In_365);
or U59 (N_59,In_177,In_134);
nor U60 (N_60,In_271,In_449);
and U61 (N_61,In_59,In_205);
and U62 (N_62,In_409,In_191);
and U63 (N_63,In_194,In_152);
and U64 (N_64,In_417,In_491);
or U65 (N_65,In_166,In_466);
nand U66 (N_66,In_314,In_6);
or U67 (N_67,In_252,In_171);
nand U68 (N_68,In_210,In_493);
nor U69 (N_69,In_249,N_22);
and U70 (N_70,N_9,In_78);
or U71 (N_71,In_42,In_273);
and U72 (N_72,In_451,In_142);
nor U73 (N_73,In_192,In_416);
nor U74 (N_74,In_293,In_377);
and U75 (N_75,In_0,In_439);
and U76 (N_76,In_308,In_50);
and U77 (N_77,In_16,In_88);
nand U78 (N_78,In_65,In_280);
nand U79 (N_79,In_208,In_101);
nand U80 (N_80,In_454,In_481);
or U81 (N_81,In_226,In_85);
nand U82 (N_82,In_324,In_367);
or U83 (N_83,In_479,N_52);
nor U84 (N_84,In_27,In_160);
and U85 (N_85,In_30,N_12);
nor U86 (N_86,In_187,In_334);
nand U87 (N_87,In_289,In_146);
nand U88 (N_88,In_320,In_128);
or U89 (N_89,In_297,In_384);
nor U90 (N_90,N_33,In_433);
or U91 (N_91,In_5,N_23);
nand U92 (N_92,In_494,In_322);
and U93 (N_93,In_375,In_109);
or U94 (N_94,In_266,In_354);
and U95 (N_95,In_475,In_26);
nand U96 (N_96,N_38,In_107);
or U97 (N_97,In_268,In_440);
and U98 (N_98,N_18,In_175);
and U99 (N_99,In_411,In_202);
nand U100 (N_100,In_189,In_207);
or U101 (N_101,N_30,In_119);
and U102 (N_102,N_13,In_102);
and U103 (N_103,In_243,In_113);
nand U104 (N_104,In_453,In_96);
or U105 (N_105,In_437,In_216);
or U106 (N_106,In_472,In_485);
nor U107 (N_107,N_0,In_167);
or U108 (N_108,In_105,In_28);
nand U109 (N_109,In_159,N_34);
or U110 (N_110,In_127,In_183);
or U111 (N_111,In_120,N_24);
and U112 (N_112,In_307,In_338);
or U113 (N_113,In_376,In_301);
and U114 (N_114,In_124,In_203);
nor U115 (N_115,N_55,N_56);
nand U116 (N_116,In_332,In_126);
nor U117 (N_117,In_278,In_330);
or U118 (N_118,In_349,In_274);
and U119 (N_119,In_443,In_283);
nor U120 (N_120,In_32,In_122);
and U121 (N_121,In_18,In_499);
nand U122 (N_122,In_182,N_4);
nand U123 (N_123,In_295,N_112);
nand U124 (N_124,In_158,In_262);
and U125 (N_125,In_62,N_7);
nor U126 (N_126,N_54,In_184);
xnor U127 (N_127,In_76,N_84);
and U128 (N_128,N_57,N_76);
nor U129 (N_129,In_402,In_198);
nor U130 (N_130,In_370,N_39);
nand U131 (N_131,In_110,In_235);
and U132 (N_132,In_413,In_357);
nor U133 (N_133,In_73,N_27);
nand U134 (N_134,In_53,N_6);
or U135 (N_135,In_318,In_213);
and U136 (N_136,In_83,In_284);
or U137 (N_137,N_36,In_406);
nor U138 (N_138,In_219,In_398);
xnor U139 (N_139,In_294,In_407);
or U140 (N_140,In_310,N_16);
nor U141 (N_141,N_35,In_399);
or U142 (N_142,In_465,N_41);
nand U143 (N_143,In_379,In_261);
nand U144 (N_144,In_250,In_305);
or U145 (N_145,In_147,In_144);
nand U146 (N_146,In_9,N_59);
and U147 (N_147,In_106,N_99);
nand U148 (N_148,In_426,N_44);
nor U149 (N_149,In_345,In_70);
and U150 (N_150,N_100,N_51);
nand U151 (N_151,In_228,N_50);
or U152 (N_152,In_133,N_96);
and U153 (N_153,In_363,In_25);
nand U154 (N_154,N_89,In_169);
or U155 (N_155,N_115,N_43);
nor U156 (N_156,In_342,N_11);
nor U157 (N_157,N_110,N_113);
nand U158 (N_158,In_108,N_60);
or U159 (N_159,In_329,In_364);
and U160 (N_160,In_344,In_43);
or U161 (N_161,In_244,In_369);
nor U162 (N_162,N_14,In_313);
nand U163 (N_163,N_117,In_199);
or U164 (N_164,In_452,In_291);
or U165 (N_165,In_149,In_118);
and U166 (N_166,N_82,In_87);
nand U167 (N_167,In_495,In_211);
nand U168 (N_168,N_66,In_3);
and U169 (N_169,In_240,In_173);
and U170 (N_170,N_29,In_31);
and U171 (N_171,In_431,In_204);
or U172 (N_172,In_461,In_455);
nor U173 (N_173,N_91,In_395);
and U174 (N_174,N_46,N_65);
nor U175 (N_175,In_424,In_361);
or U176 (N_176,In_312,In_131);
nor U177 (N_177,N_25,In_212);
nor U178 (N_178,N_85,N_119);
nor U179 (N_179,In_69,In_20);
and U180 (N_180,In_237,In_234);
or U181 (N_181,In_34,In_341);
nor U182 (N_182,N_179,N_10);
nand U183 (N_183,In_366,N_160);
or U184 (N_184,In_467,In_303);
or U185 (N_185,In_57,N_105);
or U186 (N_186,In_236,In_488);
nand U187 (N_187,In_434,In_41);
and U188 (N_188,In_425,In_111);
nand U189 (N_189,In_84,In_279);
nor U190 (N_190,N_68,In_97);
nand U191 (N_191,N_8,In_233);
nand U192 (N_192,N_144,In_90);
xnor U193 (N_193,N_37,In_13);
nor U194 (N_194,N_107,In_299);
nand U195 (N_195,N_75,In_296);
and U196 (N_196,N_31,N_106);
nand U197 (N_197,In_165,In_75);
or U198 (N_198,N_125,N_162);
or U199 (N_199,N_19,N_72);
or U200 (N_200,In_281,N_95);
nand U201 (N_201,N_93,In_72);
nor U202 (N_202,In_98,In_480);
nor U203 (N_203,In_347,N_170);
nand U204 (N_204,N_80,In_323);
nand U205 (N_205,In_360,N_135);
nor U206 (N_206,In_333,N_94);
nor U207 (N_207,In_54,In_242);
nand U208 (N_208,In_358,In_456);
or U209 (N_209,In_351,N_127);
nand U210 (N_210,In_422,N_158);
nor U211 (N_211,In_429,In_359);
and U212 (N_212,N_118,N_143);
nand U213 (N_213,N_155,In_270);
or U214 (N_214,In_135,In_143);
and U215 (N_215,N_92,In_185);
nor U216 (N_216,In_64,N_150);
and U217 (N_217,N_3,In_259);
and U218 (N_218,In_2,In_412);
nand U219 (N_219,In_8,In_190);
or U220 (N_220,In_441,N_167);
and U221 (N_221,In_335,In_340);
or U222 (N_222,N_42,In_17);
nand U223 (N_223,In_331,N_97);
xnor U224 (N_224,N_78,N_28);
nor U225 (N_225,N_21,N_98);
nand U226 (N_226,In_394,In_193);
nand U227 (N_227,N_176,N_147);
nor U228 (N_228,In_290,N_40);
nand U229 (N_229,In_287,N_109);
and U230 (N_230,N_70,In_275);
nand U231 (N_231,N_53,In_248);
and U232 (N_232,N_169,In_405);
nor U233 (N_233,N_108,In_321);
or U234 (N_234,In_180,In_24);
nor U235 (N_235,N_67,N_141);
nand U236 (N_236,In_430,N_145);
and U237 (N_237,N_142,In_267);
and U238 (N_238,In_457,In_47);
or U239 (N_239,In_319,In_497);
nor U240 (N_240,N_165,N_177);
and U241 (N_241,In_100,N_219);
and U242 (N_242,N_184,In_387);
and U243 (N_243,N_83,N_171);
nor U244 (N_244,N_213,N_178);
nand U245 (N_245,N_227,N_196);
nor U246 (N_246,In_201,In_151);
or U247 (N_247,In_317,In_311);
nor U248 (N_248,N_77,N_104);
nand U249 (N_249,N_202,N_32);
nor U250 (N_250,N_189,In_282);
nor U251 (N_251,N_199,N_86);
and U252 (N_252,In_161,In_241);
or U253 (N_253,In_385,N_223);
or U254 (N_254,N_207,N_5);
or U255 (N_255,N_215,In_445);
or U256 (N_256,N_197,N_128);
nand U257 (N_257,In_33,N_222);
nor U258 (N_258,In_7,N_88);
and U259 (N_259,In_157,N_237);
and U260 (N_260,In_136,N_140);
and U261 (N_261,N_126,In_163);
nand U262 (N_262,N_15,In_419);
or U263 (N_263,In_92,N_63);
and U264 (N_264,In_217,In_221);
and U265 (N_265,N_190,In_325);
or U266 (N_266,In_470,N_116);
nor U267 (N_267,N_182,N_208);
or U268 (N_268,In_473,N_48);
nand U269 (N_269,N_180,N_209);
nand U270 (N_270,N_203,N_111);
and U271 (N_271,In_298,N_101);
or U272 (N_272,In_1,N_232);
and U273 (N_273,In_141,N_225);
or U274 (N_274,In_484,N_216);
and U275 (N_275,N_164,N_73);
or U276 (N_276,N_212,N_156);
nor U277 (N_277,In_99,N_149);
or U278 (N_278,N_175,In_418);
or U279 (N_279,In_435,N_131);
nor U280 (N_280,N_62,N_120);
nand U281 (N_281,N_186,N_195);
nor U282 (N_282,In_486,In_258);
nand U283 (N_283,In_468,In_257);
nor U284 (N_284,N_218,In_380);
or U285 (N_285,N_123,N_69);
nand U286 (N_286,N_168,N_2);
or U287 (N_287,In_254,N_81);
nor U288 (N_288,N_228,In_378);
nand U289 (N_289,N_214,In_383);
nand U290 (N_290,N_198,N_45);
nand U291 (N_291,N_230,In_328);
and U292 (N_292,N_205,In_476);
nor U293 (N_293,In_44,N_166);
nor U294 (N_294,N_157,N_136);
and U295 (N_295,In_93,In_400);
nand U296 (N_296,In_38,In_232);
or U297 (N_297,In_200,N_192);
and U298 (N_298,In_11,In_164);
or U299 (N_299,N_26,In_458);
and U300 (N_300,In_276,N_181);
and U301 (N_301,N_172,N_152);
or U302 (N_302,In_224,In_397);
or U303 (N_303,N_235,N_286);
or U304 (N_304,In_170,N_295);
or U305 (N_305,In_153,N_244);
and U306 (N_306,In_388,N_20);
or U307 (N_307,N_259,In_421);
nor U308 (N_308,N_248,N_234);
or U309 (N_309,N_292,In_382);
and U310 (N_310,N_211,N_262);
nand U311 (N_311,N_138,N_267);
or U312 (N_312,In_247,In_155);
nand U313 (N_313,N_194,N_266);
and U314 (N_314,N_139,N_283);
nand U315 (N_315,In_218,N_246);
and U316 (N_316,N_71,In_179);
nor U317 (N_317,N_298,N_121);
nand U318 (N_318,In_327,In_79);
or U319 (N_319,N_261,In_22);
nand U320 (N_320,In_86,N_255);
nand U321 (N_321,N_217,N_284);
nand U322 (N_322,In_138,N_133);
nand U323 (N_323,N_294,N_49);
and U324 (N_324,N_224,In_71);
nor U325 (N_325,N_17,N_245);
nor U326 (N_326,N_270,N_191);
nand U327 (N_327,In_35,In_371);
or U328 (N_328,N_233,N_240);
and U329 (N_329,In_459,In_264);
or U330 (N_330,N_279,In_239);
and U331 (N_331,In_10,N_183);
nand U332 (N_332,In_373,N_282);
nor U333 (N_333,N_154,In_442);
and U334 (N_334,In_172,N_87);
nor U335 (N_335,In_337,N_200);
or U336 (N_336,In_444,N_204);
or U337 (N_337,N_220,N_229);
nor U338 (N_338,N_206,In_176);
and U339 (N_339,N_260,N_146);
or U340 (N_340,N_231,In_410);
or U341 (N_341,N_250,In_29);
and U342 (N_342,In_37,N_226);
nand U343 (N_343,N_272,N_124);
and U344 (N_344,N_241,N_174);
and U345 (N_345,N_290,In_162);
nor U346 (N_346,N_275,N_159);
or U347 (N_347,N_287,N_79);
nand U348 (N_348,In_49,N_243);
nor U349 (N_349,In_316,N_277);
nor U350 (N_350,In_315,N_193);
or U351 (N_351,N_265,N_274);
nor U352 (N_352,In_56,N_161);
and U353 (N_353,N_281,In_68);
and U354 (N_354,N_132,In_137);
nand U355 (N_355,In_414,N_254);
nor U356 (N_356,In_123,N_242);
nor U357 (N_357,In_309,In_95);
nand U358 (N_358,N_288,N_247);
nand U359 (N_359,N_278,N_251);
and U360 (N_360,N_185,In_498);
nand U361 (N_361,N_103,N_258);
or U362 (N_362,N_345,In_156);
or U363 (N_363,N_355,In_255);
nor U364 (N_364,In_89,N_299);
and U365 (N_365,N_289,N_151);
and U366 (N_366,N_291,N_349);
or U367 (N_367,N_306,N_359);
nand U368 (N_368,N_352,In_39);
nand U369 (N_369,N_354,In_94);
or U370 (N_370,N_336,N_102);
or U371 (N_371,N_269,N_339);
nand U372 (N_372,N_153,In_348);
and U373 (N_373,N_305,N_256);
or U374 (N_374,N_302,N_337);
nor U375 (N_375,N_307,N_356);
and U376 (N_376,N_328,N_114);
nor U377 (N_377,N_329,N_342);
or U378 (N_378,N_271,N_173);
nor U379 (N_379,N_319,N_313);
or U380 (N_380,N_163,N_61);
nor U381 (N_381,In_40,In_103);
or U382 (N_382,In_389,N_325);
or U383 (N_383,N_344,In_386);
nor U384 (N_384,N_249,N_326);
nor U385 (N_385,N_348,In_251);
and U386 (N_386,N_353,In_245);
nand U387 (N_387,N_358,N_334);
nor U388 (N_388,N_347,N_285);
nand U389 (N_389,In_174,N_323);
and U390 (N_390,N_310,N_350);
or U391 (N_391,N_303,N_312);
nand U392 (N_392,N_239,N_322);
nand U393 (N_393,N_148,N_357);
nor U394 (N_394,N_324,N_280);
and U395 (N_395,In_91,N_273);
or U396 (N_396,N_346,N_264);
or U397 (N_397,In_343,N_221);
nand U398 (N_398,N_276,N_122);
nor U399 (N_399,N_343,In_229);
or U400 (N_400,N_304,N_318);
nand U401 (N_401,In_263,N_327);
and U402 (N_402,In_188,In_415);
or U403 (N_403,N_257,N_309);
nand U404 (N_404,N_58,N_253);
and U405 (N_405,In_222,N_130);
nor U406 (N_406,N_333,N_316);
nor U407 (N_407,N_201,N_297);
and U408 (N_408,N_236,N_308);
or U409 (N_409,N_134,N_293);
or U410 (N_410,N_332,N_210);
or U411 (N_411,N_1,In_178);
and U412 (N_412,N_330,N_311);
nor U413 (N_413,N_129,N_331);
or U414 (N_414,In_423,N_263);
nand U415 (N_415,In_438,N_335);
nor U416 (N_416,N_320,In_66);
nor U417 (N_417,N_321,In_469);
and U418 (N_418,In_209,N_90);
or U419 (N_419,N_74,N_238);
nand U420 (N_420,N_408,N_381);
or U421 (N_421,N_341,N_399);
nor U422 (N_422,N_409,N_315);
nand U423 (N_423,N_372,N_366);
and U424 (N_424,N_401,N_400);
and U425 (N_425,N_338,N_407);
nor U426 (N_426,N_317,N_351);
and U427 (N_427,N_403,N_418);
nand U428 (N_428,N_187,N_379);
or U429 (N_429,N_374,N_402);
nand U430 (N_430,N_414,N_404);
nand U431 (N_431,N_361,N_367);
nand U432 (N_432,N_388,N_380);
and U433 (N_433,N_268,N_396);
and U434 (N_434,N_419,In_215);
and U435 (N_435,N_413,N_301);
nand U436 (N_436,N_398,N_394);
nor U437 (N_437,N_252,N_64);
or U438 (N_438,N_340,N_376);
or U439 (N_439,N_385,N_415);
nand U440 (N_440,N_370,N_397);
nor U441 (N_441,N_417,N_300);
and U442 (N_442,N_405,N_395);
and U443 (N_443,N_47,N_378);
nor U444 (N_444,N_412,N_373);
and U445 (N_445,In_462,N_365);
or U446 (N_446,N_389,N_188);
xor U447 (N_447,N_371,N_410);
or U448 (N_448,N_386,N_392);
nor U449 (N_449,N_362,N_382);
and U450 (N_450,N_384,N_369);
or U451 (N_451,N_360,N_368);
or U452 (N_452,N_416,N_363);
nand U453 (N_453,N_391,N_375);
or U454 (N_454,N_406,N_390);
nor U455 (N_455,In_148,N_137);
nor U456 (N_456,N_364,N_314);
nand U457 (N_457,N_393,N_411);
nand U458 (N_458,N_296,N_387);
or U459 (N_459,N_377,N_383);
or U460 (N_460,N_394,N_406);
and U461 (N_461,N_137,N_384);
nand U462 (N_462,N_367,N_407);
or U463 (N_463,N_377,N_396);
nand U464 (N_464,N_377,N_374);
and U465 (N_465,N_296,N_388);
xor U466 (N_466,N_405,N_315);
or U467 (N_467,N_368,N_296);
and U468 (N_468,N_407,N_360);
nor U469 (N_469,N_340,N_365);
nand U470 (N_470,N_414,N_386);
nand U471 (N_471,N_377,N_188);
and U472 (N_472,N_187,N_373);
nand U473 (N_473,N_314,N_296);
nand U474 (N_474,N_385,N_387);
nand U475 (N_475,N_314,N_399);
nor U476 (N_476,N_391,N_390);
nand U477 (N_477,N_383,N_366);
nor U478 (N_478,N_370,In_148);
nor U479 (N_479,N_363,N_409);
or U480 (N_480,N_442,N_473);
nand U481 (N_481,N_455,N_475);
and U482 (N_482,N_468,N_428);
or U483 (N_483,N_433,N_454);
nor U484 (N_484,N_453,N_466);
and U485 (N_485,N_447,N_427);
nor U486 (N_486,N_439,N_448);
or U487 (N_487,N_429,N_426);
nand U488 (N_488,N_425,N_471);
nand U489 (N_489,N_470,N_436);
or U490 (N_490,N_440,N_432);
and U491 (N_491,N_452,N_467);
or U492 (N_492,N_479,N_476);
and U493 (N_493,N_464,N_445);
nor U494 (N_494,N_451,N_424);
or U495 (N_495,N_469,N_430);
or U496 (N_496,N_441,N_458);
nand U497 (N_497,N_463,N_431);
and U498 (N_498,N_421,N_457);
or U499 (N_499,N_444,N_446);
and U500 (N_500,N_474,N_478);
and U501 (N_501,N_437,N_460);
nand U502 (N_502,N_477,N_435);
nor U503 (N_503,N_438,N_443);
and U504 (N_504,N_472,N_434);
xnor U505 (N_505,N_423,N_420);
or U506 (N_506,N_422,N_465);
or U507 (N_507,N_461,N_459);
and U508 (N_508,N_449,N_450);
and U509 (N_509,N_456,N_462);
nor U510 (N_510,N_472,N_443);
or U511 (N_511,N_476,N_432);
and U512 (N_512,N_477,N_459);
and U513 (N_513,N_450,N_425);
nand U514 (N_514,N_445,N_457);
xor U515 (N_515,N_453,N_469);
or U516 (N_516,N_473,N_479);
nand U517 (N_517,N_431,N_430);
nor U518 (N_518,N_436,N_471);
nor U519 (N_519,N_435,N_474);
or U520 (N_520,N_424,N_440);
and U521 (N_521,N_469,N_427);
and U522 (N_522,N_432,N_425);
and U523 (N_523,N_452,N_436);
nand U524 (N_524,N_434,N_465);
and U525 (N_525,N_451,N_471);
or U526 (N_526,N_465,N_460);
nand U527 (N_527,N_459,N_456);
and U528 (N_528,N_425,N_434);
or U529 (N_529,N_461,N_440);
or U530 (N_530,N_472,N_437);
nand U531 (N_531,N_479,N_449);
and U532 (N_532,N_470,N_444);
and U533 (N_533,N_427,N_443);
and U534 (N_534,N_479,N_475);
and U535 (N_535,N_478,N_453);
or U536 (N_536,N_479,N_471);
nand U537 (N_537,N_435,N_459);
and U538 (N_538,N_467,N_479);
and U539 (N_539,N_423,N_445);
nor U540 (N_540,N_480,N_511);
or U541 (N_541,N_529,N_514);
or U542 (N_542,N_506,N_499);
nand U543 (N_543,N_522,N_491);
and U544 (N_544,N_508,N_496);
and U545 (N_545,N_535,N_482);
or U546 (N_546,N_505,N_483);
nor U547 (N_547,N_489,N_523);
and U548 (N_548,N_520,N_502);
and U549 (N_549,N_527,N_534);
and U550 (N_550,N_526,N_485);
xor U551 (N_551,N_516,N_492);
and U552 (N_552,N_536,N_513);
and U553 (N_553,N_500,N_490);
and U554 (N_554,N_493,N_532);
nor U555 (N_555,N_481,N_501);
or U556 (N_556,N_488,N_486);
and U557 (N_557,N_521,N_504);
nor U558 (N_558,N_515,N_537);
nand U559 (N_559,N_487,N_509);
or U560 (N_560,N_538,N_484);
and U561 (N_561,N_494,N_531);
and U562 (N_562,N_524,N_497);
or U563 (N_563,N_512,N_519);
or U564 (N_564,N_517,N_533);
and U565 (N_565,N_530,N_510);
or U566 (N_566,N_518,N_525);
nand U567 (N_567,N_495,N_503);
nand U568 (N_568,N_528,N_539);
nor U569 (N_569,N_507,N_498);
or U570 (N_570,N_490,N_517);
nand U571 (N_571,N_515,N_489);
nor U572 (N_572,N_505,N_507);
or U573 (N_573,N_524,N_508);
or U574 (N_574,N_521,N_528);
or U575 (N_575,N_509,N_528);
nor U576 (N_576,N_490,N_538);
or U577 (N_577,N_538,N_488);
nor U578 (N_578,N_495,N_529);
nor U579 (N_579,N_522,N_508);
and U580 (N_580,N_499,N_531);
nor U581 (N_581,N_538,N_521);
nand U582 (N_582,N_519,N_486);
nor U583 (N_583,N_525,N_515);
nand U584 (N_584,N_483,N_534);
or U585 (N_585,N_491,N_499);
nor U586 (N_586,N_536,N_510);
nor U587 (N_587,N_484,N_492);
nor U588 (N_588,N_521,N_513);
or U589 (N_589,N_505,N_536);
nand U590 (N_590,N_535,N_503);
nand U591 (N_591,N_495,N_502);
and U592 (N_592,N_484,N_517);
nor U593 (N_593,N_515,N_480);
nor U594 (N_594,N_506,N_519);
nand U595 (N_595,N_506,N_500);
or U596 (N_596,N_490,N_537);
nor U597 (N_597,N_532,N_529);
nor U598 (N_598,N_539,N_513);
nor U599 (N_599,N_482,N_485);
nand U600 (N_600,N_553,N_556);
nor U601 (N_601,N_557,N_591);
or U602 (N_602,N_578,N_570);
and U603 (N_603,N_574,N_568);
nand U604 (N_604,N_566,N_549);
nor U605 (N_605,N_592,N_565);
nor U606 (N_606,N_582,N_590);
and U607 (N_607,N_597,N_552);
or U608 (N_608,N_575,N_551);
nor U609 (N_609,N_554,N_548);
and U610 (N_610,N_585,N_598);
or U611 (N_611,N_546,N_544);
and U612 (N_612,N_560,N_586);
nand U613 (N_613,N_577,N_569);
nand U614 (N_614,N_561,N_588);
or U615 (N_615,N_572,N_580);
or U616 (N_616,N_581,N_559);
or U617 (N_617,N_593,N_579);
and U618 (N_618,N_555,N_543);
and U619 (N_619,N_584,N_563);
or U620 (N_620,N_567,N_564);
nand U621 (N_621,N_595,N_594);
nor U622 (N_622,N_589,N_550);
nand U623 (N_623,N_587,N_571);
and U624 (N_624,N_547,N_542);
or U625 (N_625,N_545,N_576);
nand U626 (N_626,N_562,N_573);
nand U627 (N_627,N_599,N_596);
or U628 (N_628,N_541,N_558);
and U629 (N_629,N_540,N_583);
nand U630 (N_630,N_575,N_594);
nor U631 (N_631,N_564,N_549);
nor U632 (N_632,N_594,N_563);
nand U633 (N_633,N_597,N_576);
and U634 (N_634,N_566,N_595);
nor U635 (N_635,N_561,N_562);
nor U636 (N_636,N_598,N_573);
and U637 (N_637,N_570,N_596);
nor U638 (N_638,N_599,N_541);
nand U639 (N_639,N_568,N_557);
or U640 (N_640,N_598,N_584);
nand U641 (N_641,N_540,N_588);
nand U642 (N_642,N_552,N_588);
nor U643 (N_643,N_542,N_575);
or U644 (N_644,N_558,N_549);
and U645 (N_645,N_573,N_550);
nand U646 (N_646,N_552,N_568);
nor U647 (N_647,N_551,N_547);
and U648 (N_648,N_580,N_588);
or U649 (N_649,N_555,N_574);
and U650 (N_650,N_543,N_561);
or U651 (N_651,N_547,N_552);
nor U652 (N_652,N_575,N_550);
nand U653 (N_653,N_545,N_575);
or U654 (N_654,N_595,N_564);
nor U655 (N_655,N_541,N_578);
xor U656 (N_656,N_558,N_580);
or U657 (N_657,N_554,N_571);
and U658 (N_658,N_545,N_555);
and U659 (N_659,N_557,N_578);
and U660 (N_660,N_628,N_651);
nand U661 (N_661,N_627,N_637);
and U662 (N_662,N_641,N_623);
nand U663 (N_663,N_625,N_646);
nor U664 (N_664,N_603,N_631);
or U665 (N_665,N_642,N_634);
and U666 (N_666,N_656,N_601);
and U667 (N_667,N_604,N_619);
nor U668 (N_668,N_653,N_632);
or U669 (N_669,N_629,N_639);
or U670 (N_670,N_622,N_657);
or U671 (N_671,N_621,N_606);
nand U672 (N_672,N_611,N_654);
nand U673 (N_673,N_638,N_643);
nand U674 (N_674,N_655,N_607);
and U675 (N_675,N_626,N_630);
nand U676 (N_676,N_612,N_618);
and U677 (N_677,N_652,N_608);
or U678 (N_678,N_613,N_659);
nor U679 (N_679,N_610,N_645);
and U680 (N_680,N_620,N_640);
and U681 (N_681,N_602,N_648);
nand U682 (N_682,N_647,N_644);
or U683 (N_683,N_649,N_658);
and U684 (N_684,N_614,N_609);
or U685 (N_685,N_615,N_605);
nand U686 (N_686,N_635,N_600);
nand U687 (N_687,N_633,N_617);
nand U688 (N_688,N_616,N_624);
or U689 (N_689,N_636,N_650);
nand U690 (N_690,N_618,N_628);
nor U691 (N_691,N_615,N_651);
nor U692 (N_692,N_612,N_636);
and U693 (N_693,N_651,N_643);
and U694 (N_694,N_617,N_626);
or U695 (N_695,N_633,N_604);
nand U696 (N_696,N_635,N_650);
nand U697 (N_697,N_622,N_602);
or U698 (N_698,N_636,N_633);
and U699 (N_699,N_632,N_633);
nor U700 (N_700,N_639,N_649);
or U701 (N_701,N_632,N_639);
or U702 (N_702,N_655,N_656);
nand U703 (N_703,N_648,N_603);
or U704 (N_704,N_640,N_610);
or U705 (N_705,N_624,N_656);
nand U706 (N_706,N_622,N_653);
nand U707 (N_707,N_633,N_656);
or U708 (N_708,N_613,N_623);
and U709 (N_709,N_607,N_657);
nand U710 (N_710,N_612,N_659);
and U711 (N_711,N_655,N_644);
nor U712 (N_712,N_633,N_627);
nor U713 (N_713,N_638,N_628);
nor U714 (N_714,N_620,N_635);
or U715 (N_715,N_649,N_619);
and U716 (N_716,N_619,N_648);
nand U717 (N_717,N_655,N_651);
xnor U718 (N_718,N_636,N_618);
nand U719 (N_719,N_657,N_604);
nor U720 (N_720,N_676,N_690);
or U721 (N_721,N_668,N_663);
or U722 (N_722,N_679,N_675);
nor U723 (N_723,N_673,N_678);
or U724 (N_724,N_706,N_688);
and U725 (N_725,N_704,N_713);
or U726 (N_726,N_710,N_702);
nand U727 (N_727,N_677,N_689);
or U728 (N_728,N_674,N_666);
and U729 (N_729,N_703,N_715);
nor U730 (N_730,N_664,N_694);
nand U731 (N_731,N_692,N_709);
nor U732 (N_732,N_699,N_707);
nor U733 (N_733,N_671,N_719);
nor U734 (N_734,N_708,N_683);
xor U735 (N_735,N_682,N_667);
nand U736 (N_736,N_684,N_705);
nand U737 (N_737,N_686,N_712);
and U738 (N_738,N_680,N_698);
nor U739 (N_739,N_697,N_687);
and U740 (N_740,N_670,N_695);
nor U741 (N_741,N_661,N_711);
nand U742 (N_742,N_691,N_700);
nor U743 (N_743,N_660,N_669);
and U744 (N_744,N_685,N_696);
nand U745 (N_745,N_701,N_718);
nand U746 (N_746,N_672,N_681);
or U747 (N_747,N_665,N_716);
and U748 (N_748,N_714,N_717);
nor U749 (N_749,N_662,N_693);
and U750 (N_750,N_719,N_662);
nand U751 (N_751,N_661,N_671);
nand U752 (N_752,N_715,N_677);
and U753 (N_753,N_701,N_662);
nor U754 (N_754,N_673,N_689);
nand U755 (N_755,N_670,N_709);
nor U756 (N_756,N_712,N_692);
nand U757 (N_757,N_703,N_712);
and U758 (N_758,N_669,N_706);
or U759 (N_759,N_711,N_694);
nor U760 (N_760,N_704,N_661);
or U761 (N_761,N_694,N_707);
and U762 (N_762,N_691,N_682);
and U763 (N_763,N_669,N_698);
nor U764 (N_764,N_690,N_703);
and U765 (N_765,N_696,N_717);
nor U766 (N_766,N_687,N_678);
nor U767 (N_767,N_703,N_693);
nand U768 (N_768,N_696,N_671);
nand U769 (N_769,N_666,N_715);
nor U770 (N_770,N_690,N_714);
nand U771 (N_771,N_716,N_670);
nor U772 (N_772,N_673,N_695);
nor U773 (N_773,N_706,N_693);
and U774 (N_774,N_702,N_688);
or U775 (N_775,N_662,N_699);
and U776 (N_776,N_673,N_675);
nand U777 (N_777,N_683,N_686);
or U778 (N_778,N_676,N_702);
nand U779 (N_779,N_699,N_701);
or U780 (N_780,N_740,N_750);
nor U781 (N_781,N_755,N_775);
nor U782 (N_782,N_765,N_772);
nor U783 (N_783,N_766,N_728);
nor U784 (N_784,N_730,N_749);
and U785 (N_785,N_744,N_769);
nor U786 (N_786,N_767,N_758);
and U787 (N_787,N_720,N_751);
or U788 (N_788,N_770,N_753);
and U789 (N_789,N_736,N_761);
nand U790 (N_790,N_757,N_721);
or U791 (N_791,N_742,N_754);
nand U792 (N_792,N_732,N_726);
nand U793 (N_793,N_748,N_779);
and U794 (N_794,N_737,N_762);
nor U795 (N_795,N_735,N_724);
and U796 (N_796,N_745,N_727);
nor U797 (N_797,N_778,N_752);
and U798 (N_798,N_771,N_760);
nor U799 (N_799,N_773,N_733);
or U800 (N_800,N_723,N_768);
or U801 (N_801,N_747,N_763);
nor U802 (N_802,N_741,N_759);
and U803 (N_803,N_777,N_739);
nor U804 (N_804,N_776,N_729);
and U805 (N_805,N_743,N_756);
nand U806 (N_806,N_725,N_774);
or U807 (N_807,N_746,N_722);
or U808 (N_808,N_738,N_734);
and U809 (N_809,N_764,N_731);
or U810 (N_810,N_744,N_776);
and U811 (N_811,N_766,N_755);
nand U812 (N_812,N_765,N_747);
or U813 (N_813,N_779,N_762);
nor U814 (N_814,N_751,N_745);
or U815 (N_815,N_727,N_721);
nor U816 (N_816,N_777,N_723);
nand U817 (N_817,N_773,N_772);
or U818 (N_818,N_752,N_722);
or U819 (N_819,N_747,N_772);
nand U820 (N_820,N_771,N_750);
xor U821 (N_821,N_738,N_762);
or U822 (N_822,N_720,N_776);
nand U823 (N_823,N_751,N_772);
nor U824 (N_824,N_722,N_729);
and U825 (N_825,N_764,N_761);
and U826 (N_826,N_776,N_741);
or U827 (N_827,N_777,N_745);
nand U828 (N_828,N_740,N_747);
nor U829 (N_829,N_772,N_720);
nor U830 (N_830,N_731,N_745);
or U831 (N_831,N_745,N_746);
and U832 (N_832,N_728,N_721);
nor U833 (N_833,N_751,N_726);
and U834 (N_834,N_722,N_777);
and U835 (N_835,N_747,N_726);
nand U836 (N_836,N_767,N_742);
or U837 (N_837,N_721,N_746);
nand U838 (N_838,N_772,N_758);
nand U839 (N_839,N_748,N_777);
and U840 (N_840,N_830,N_810);
or U841 (N_841,N_838,N_833);
nand U842 (N_842,N_818,N_780);
nand U843 (N_843,N_781,N_814);
nand U844 (N_844,N_836,N_820);
nand U845 (N_845,N_794,N_784);
or U846 (N_846,N_806,N_832);
nor U847 (N_847,N_783,N_812);
and U848 (N_848,N_787,N_785);
and U849 (N_849,N_828,N_807);
nor U850 (N_850,N_802,N_801);
nand U851 (N_851,N_813,N_823);
or U852 (N_852,N_800,N_793);
and U853 (N_853,N_835,N_824);
and U854 (N_854,N_786,N_831);
nor U855 (N_855,N_837,N_811);
or U856 (N_856,N_826,N_809);
nand U857 (N_857,N_808,N_817);
nand U858 (N_858,N_822,N_791);
nor U859 (N_859,N_827,N_816);
nand U860 (N_860,N_825,N_790);
and U861 (N_861,N_797,N_815);
nor U862 (N_862,N_829,N_798);
and U863 (N_863,N_799,N_839);
or U864 (N_864,N_805,N_821);
and U865 (N_865,N_788,N_782);
nand U866 (N_866,N_789,N_803);
and U867 (N_867,N_819,N_792);
and U868 (N_868,N_834,N_804);
nor U869 (N_869,N_796,N_795);
nand U870 (N_870,N_830,N_784);
or U871 (N_871,N_791,N_815);
or U872 (N_872,N_793,N_812);
nand U873 (N_873,N_824,N_807);
nor U874 (N_874,N_817,N_805);
nor U875 (N_875,N_807,N_832);
nand U876 (N_876,N_795,N_837);
nand U877 (N_877,N_828,N_805);
and U878 (N_878,N_806,N_801);
nor U879 (N_879,N_804,N_833);
and U880 (N_880,N_839,N_822);
nand U881 (N_881,N_819,N_817);
or U882 (N_882,N_793,N_835);
and U883 (N_883,N_815,N_814);
and U884 (N_884,N_790,N_810);
nor U885 (N_885,N_824,N_808);
nand U886 (N_886,N_829,N_834);
nand U887 (N_887,N_811,N_787);
or U888 (N_888,N_815,N_800);
and U889 (N_889,N_795,N_790);
nand U890 (N_890,N_789,N_822);
and U891 (N_891,N_781,N_811);
and U892 (N_892,N_783,N_794);
nor U893 (N_893,N_821,N_822);
or U894 (N_894,N_823,N_800);
and U895 (N_895,N_836,N_808);
and U896 (N_896,N_825,N_817);
or U897 (N_897,N_819,N_836);
xnor U898 (N_898,N_793,N_794);
xnor U899 (N_899,N_838,N_796);
and U900 (N_900,N_898,N_879);
nor U901 (N_901,N_880,N_886);
nand U902 (N_902,N_857,N_854);
nor U903 (N_903,N_896,N_878);
or U904 (N_904,N_861,N_847);
and U905 (N_905,N_842,N_862);
nor U906 (N_906,N_892,N_889);
nand U907 (N_907,N_881,N_875);
nand U908 (N_908,N_883,N_899);
nor U909 (N_909,N_845,N_849);
nand U910 (N_910,N_858,N_884);
or U911 (N_911,N_882,N_851);
nand U912 (N_912,N_895,N_846);
nand U913 (N_913,N_843,N_856);
or U914 (N_914,N_877,N_885);
or U915 (N_915,N_876,N_841);
nor U916 (N_916,N_865,N_891);
nor U917 (N_917,N_897,N_873);
nor U918 (N_918,N_869,N_866);
nand U919 (N_919,N_852,N_853);
nand U920 (N_920,N_874,N_872);
nand U921 (N_921,N_844,N_894);
or U922 (N_922,N_870,N_855);
nor U923 (N_923,N_840,N_848);
or U924 (N_924,N_864,N_890);
and U925 (N_925,N_867,N_868);
nor U926 (N_926,N_863,N_871);
and U927 (N_927,N_859,N_893);
nor U928 (N_928,N_860,N_850);
nor U929 (N_929,N_887,N_888);
and U930 (N_930,N_854,N_860);
or U931 (N_931,N_882,N_887);
or U932 (N_932,N_892,N_873);
or U933 (N_933,N_878,N_870);
or U934 (N_934,N_893,N_882);
and U935 (N_935,N_853,N_856);
nor U936 (N_936,N_865,N_889);
or U937 (N_937,N_854,N_874);
nand U938 (N_938,N_862,N_878);
nand U939 (N_939,N_877,N_888);
and U940 (N_940,N_886,N_859);
and U941 (N_941,N_871,N_840);
or U942 (N_942,N_840,N_858);
nor U943 (N_943,N_894,N_854);
nor U944 (N_944,N_847,N_863);
nor U945 (N_945,N_848,N_860);
and U946 (N_946,N_876,N_855);
and U947 (N_947,N_840,N_883);
and U948 (N_948,N_853,N_857);
nand U949 (N_949,N_866,N_889);
and U950 (N_950,N_890,N_846);
xor U951 (N_951,N_889,N_856);
nor U952 (N_952,N_861,N_844);
nor U953 (N_953,N_855,N_840);
nor U954 (N_954,N_861,N_859);
and U955 (N_955,N_850,N_863);
or U956 (N_956,N_846,N_865);
or U957 (N_957,N_842,N_872);
nor U958 (N_958,N_857,N_885);
or U959 (N_959,N_886,N_854);
nand U960 (N_960,N_904,N_941);
nand U961 (N_961,N_958,N_928);
and U962 (N_962,N_913,N_944);
nand U963 (N_963,N_949,N_945);
nor U964 (N_964,N_940,N_932);
or U965 (N_965,N_915,N_936);
or U966 (N_966,N_905,N_946);
or U967 (N_967,N_923,N_902);
or U968 (N_968,N_957,N_937);
nand U969 (N_969,N_956,N_909);
or U970 (N_970,N_939,N_959);
and U971 (N_971,N_903,N_916);
or U972 (N_972,N_950,N_907);
or U973 (N_973,N_931,N_906);
or U974 (N_974,N_942,N_908);
nand U975 (N_975,N_918,N_925);
or U976 (N_976,N_900,N_924);
nand U977 (N_977,N_927,N_954);
or U978 (N_978,N_947,N_934);
nand U979 (N_979,N_922,N_901);
nand U980 (N_980,N_951,N_920);
nor U981 (N_981,N_921,N_930);
and U982 (N_982,N_929,N_952);
nand U983 (N_983,N_911,N_919);
nand U984 (N_984,N_914,N_943);
nor U985 (N_985,N_933,N_953);
or U986 (N_986,N_938,N_912);
or U987 (N_987,N_910,N_926);
and U988 (N_988,N_935,N_948);
nand U989 (N_989,N_917,N_955);
nand U990 (N_990,N_904,N_937);
and U991 (N_991,N_914,N_911);
and U992 (N_992,N_940,N_955);
and U993 (N_993,N_936,N_957);
and U994 (N_994,N_913,N_942);
nand U995 (N_995,N_930,N_933);
nand U996 (N_996,N_927,N_933);
nor U997 (N_997,N_937,N_922);
and U998 (N_998,N_929,N_934);
xor U999 (N_999,N_938,N_914);
and U1000 (N_1000,N_920,N_955);
nand U1001 (N_1001,N_921,N_912);
and U1002 (N_1002,N_922,N_907);
or U1003 (N_1003,N_918,N_943);
nand U1004 (N_1004,N_903,N_935);
or U1005 (N_1005,N_906,N_914);
nor U1006 (N_1006,N_926,N_920);
and U1007 (N_1007,N_938,N_942);
nand U1008 (N_1008,N_928,N_902);
and U1009 (N_1009,N_904,N_910);
or U1010 (N_1010,N_941,N_959);
nand U1011 (N_1011,N_948,N_943);
nor U1012 (N_1012,N_954,N_904);
nor U1013 (N_1013,N_920,N_928);
nand U1014 (N_1014,N_917,N_950);
nor U1015 (N_1015,N_956,N_923);
nand U1016 (N_1016,N_952,N_944);
nor U1017 (N_1017,N_902,N_920);
nand U1018 (N_1018,N_912,N_920);
and U1019 (N_1019,N_943,N_959);
or U1020 (N_1020,N_968,N_989);
or U1021 (N_1021,N_1004,N_1003);
nor U1022 (N_1022,N_971,N_984);
nand U1023 (N_1023,N_980,N_1000);
nand U1024 (N_1024,N_1013,N_966);
nand U1025 (N_1025,N_1017,N_1016);
nand U1026 (N_1026,N_999,N_969);
xor U1027 (N_1027,N_1014,N_986);
nand U1028 (N_1028,N_983,N_992);
nand U1029 (N_1029,N_961,N_1018);
nand U1030 (N_1030,N_991,N_1008);
or U1031 (N_1031,N_990,N_965);
or U1032 (N_1032,N_978,N_977);
xnor U1033 (N_1033,N_964,N_976);
or U1034 (N_1034,N_1010,N_960);
and U1035 (N_1035,N_979,N_995);
or U1036 (N_1036,N_1011,N_1009);
and U1037 (N_1037,N_985,N_973);
nor U1038 (N_1038,N_975,N_974);
nor U1039 (N_1039,N_962,N_1002);
nor U1040 (N_1040,N_972,N_993);
nand U1041 (N_1041,N_998,N_1015);
and U1042 (N_1042,N_994,N_987);
nor U1043 (N_1043,N_967,N_1001);
and U1044 (N_1044,N_970,N_981);
nand U1045 (N_1045,N_997,N_996);
and U1046 (N_1046,N_982,N_1005);
nor U1047 (N_1047,N_1012,N_1019);
and U1048 (N_1048,N_1007,N_963);
nor U1049 (N_1049,N_1006,N_988);
xor U1050 (N_1050,N_988,N_981);
and U1051 (N_1051,N_994,N_967);
nand U1052 (N_1052,N_1019,N_985);
and U1053 (N_1053,N_975,N_1002);
nor U1054 (N_1054,N_980,N_1013);
and U1055 (N_1055,N_978,N_1003);
nor U1056 (N_1056,N_989,N_1012);
and U1057 (N_1057,N_993,N_1013);
or U1058 (N_1058,N_960,N_964);
and U1059 (N_1059,N_1011,N_989);
and U1060 (N_1060,N_1002,N_991);
nor U1061 (N_1061,N_972,N_984);
nor U1062 (N_1062,N_989,N_967);
or U1063 (N_1063,N_967,N_1008);
and U1064 (N_1064,N_1009,N_980);
or U1065 (N_1065,N_971,N_1014);
or U1066 (N_1066,N_1001,N_979);
nand U1067 (N_1067,N_979,N_1011);
nand U1068 (N_1068,N_1019,N_996);
xnor U1069 (N_1069,N_966,N_986);
nor U1070 (N_1070,N_1019,N_987);
nor U1071 (N_1071,N_970,N_1017);
and U1072 (N_1072,N_970,N_1008);
nand U1073 (N_1073,N_985,N_1002);
nand U1074 (N_1074,N_968,N_974);
and U1075 (N_1075,N_1002,N_1012);
or U1076 (N_1076,N_963,N_994);
and U1077 (N_1077,N_997,N_981);
nand U1078 (N_1078,N_991,N_977);
and U1079 (N_1079,N_1004,N_963);
or U1080 (N_1080,N_1023,N_1037);
or U1081 (N_1081,N_1025,N_1033);
nor U1082 (N_1082,N_1055,N_1046);
nand U1083 (N_1083,N_1031,N_1052);
nor U1084 (N_1084,N_1029,N_1054);
nor U1085 (N_1085,N_1042,N_1056);
nor U1086 (N_1086,N_1067,N_1059);
nand U1087 (N_1087,N_1065,N_1063);
nand U1088 (N_1088,N_1071,N_1024);
or U1089 (N_1089,N_1069,N_1053);
and U1090 (N_1090,N_1061,N_1066);
and U1091 (N_1091,N_1064,N_1078);
nand U1092 (N_1092,N_1040,N_1075);
and U1093 (N_1093,N_1047,N_1068);
nand U1094 (N_1094,N_1070,N_1062);
nand U1095 (N_1095,N_1032,N_1022);
nor U1096 (N_1096,N_1045,N_1044);
or U1097 (N_1097,N_1060,N_1076);
nand U1098 (N_1098,N_1026,N_1074);
xnor U1099 (N_1099,N_1048,N_1038);
nor U1100 (N_1100,N_1077,N_1043);
and U1101 (N_1101,N_1039,N_1057);
and U1102 (N_1102,N_1020,N_1051);
nand U1103 (N_1103,N_1049,N_1034);
and U1104 (N_1104,N_1027,N_1030);
or U1105 (N_1105,N_1035,N_1079);
and U1106 (N_1106,N_1072,N_1041);
and U1107 (N_1107,N_1021,N_1050);
nor U1108 (N_1108,N_1073,N_1058);
or U1109 (N_1109,N_1036,N_1028);
and U1110 (N_1110,N_1047,N_1025);
and U1111 (N_1111,N_1044,N_1066);
or U1112 (N_1112,N_1027,N_1076);
or U1113 (N_1113,N_1033,N_1057);
or U1114 (N_1114,N_1033,N_1023);
nor U1115 (N_1115,N_1053,N_1076);
nand U1116 (N_1116,N_1059,N_1026);
nand U1117 (N_1117,N_1025,N_1053);
or U1118 (N_1118,N_1062,N_1037);
nand U1119 (N_1119,N_1060,N_1070);
nand U1120 (N_1120,N_1035,N_1052);
nand U1121 (N_1121,N_1028,N_1066);
nand U1122 (N_1122,N_1040,N_1068);
and U1123 (N_1123,N_1063,N_1058);
nand U1124 (N_1124,N_1046,N_1049);
or U1125 (N_1125,N_1036,N_1041);
nand U1126 (N_1126,N_1074,N_1043);
nor U1127 (N_1127,N_1066,N_1046);
and U1128 (N_1128,N_1074,N_1068);
and U1129 (N_1129,N_1065,N_1069);
nor U1130 (N_1130,N_1029,N_1021);
nor U1131 (N_1131,N_1021,N_1057);
or U1132 (N_1132,N_1058,N_1038);
nand U1133 (N_1133,N_1021,N_1040);
or U1134 (N_1134,N_1046,N_1024);
nand U1135 (N_1135,N_1042,N_1065);
and U1136 (N_1136,N_1029,N_1042);
xor U1137 (N_1137,N_1069,N_1023);
and U1138 (N_1138,N_1033,N_1045);
or U1139 (N_1139,N_1060,N_1043);
nor U1140 (N_1140,N_1088,N_1089);
and U1141 (N_1141,N_1124,N_1094);
and U1142 (N_1142,N_1100,N_1121);
or U1143 (N_1143,N_1139,N_1098);
or U1144 (N_1144,N_1103,N_1102);
nand U1145 (N_1145,N_1120,N_1118);
or U1146 (N_1146,N_1134,N_1137);
nor U1147 (N_1147,N_1091,N_1081);
and U1148 (N_1148,N_1095,N_1101);
or U1149 (N_1149,N_1122,N_1130);
and U1150 (N_1150,N_1114,N_1126);
nand U1151 (N_1151,N_1099,N_1112);
nand U1152 (N_1152,N_1132,N_1136);
nand U1153 (N_1153,N_1129,N_1119);
or U1154 (N_1154,N_1084,N_1110);
nand U1155 (N_1155,N_1080,N_1117);
nor U1156 (N_1156,N_1093,N_1113);
and U1157 (N_1157,N_1092,N_1090);
nor U1158 (N_1158,N_1105,N_1115);
or U1159 (N_1159,N_1087,N_1131);
and U1160 (N_1160,N_1125,N_1106);
nor U1161 (N_1161,N_1097,N_1123);
nor U1162 (N_1162,N_1108,N_1116);
nand U1163 (N_1163,N_1085,N_1082);
and U1164 (N_1164,N_1138,N_1127);
and U1165 (N_1165,N_1128,N_1086);
or U1166 (N_1166,N_1083,N_1135);
xnor U1167 (N_1167,N_1133,N_1104);
nand U1168 (N_1168,N_1096,N_1109);
nor U1169 (N_1169,N_1111,N_1107);
nor U1170 (N_1170,N_1090,N_1136);
nand U1171 (N_1171,N_1124,N_1104);
nor U1172 (N_1172,N_1087,N_1122);
or U1173 (N_1173,N_1093,N_1102);
nor U1174 (N_1174,N_1127,N_1081);
or U1175 (N_1175,N_1128,N_1108);
nand U1176 (N_1176,N_1087,N_1110);
nor U1177 (N_1177,N_1124,N_1111);
and U1178 (N_1178,N_1099,N_1118);
and U1179 (N_1179,N_1134,N_1123);
or U1180 (N_1180,N_1084,N_1129);
or U1181 (N_1181,N_1103,N_1134);
and U1182 (N_1182,N_1122,N_1115);
and U1183 (N_1183,N_1120,N_1090);
and U1184 (N_1184,N_1118,N_1102);
or U1185 (N_1185,N_1106,N_1095);
and U1186 (N_1186,N_1095,N_1124);
nand U1187 (N_1187,N_1131,N_1114);
nand U1188 (N_1188,N_1096,N_1087);
and U1189 (N_1189,N_1106,N_1090);
nor U1190 (N_1190,N_1122,N_1121);
or U1191 (N_1191,N_1127,N_1109);
or U1192 (N_1192,N_1103,N_1090);
nor U1193 (N_1193,N_1132,N_1109);
nor U1194 (N_1194,N_1129,N_1113);
nand U1195 (N_1195,N_1085,N_1138);
nor U1196 (N_1196,N_1106,N_1110);
nand U1197 (N_1197,N_1087,N_1102);
and U1198 (N_1198,N_1080,N_1136);
and U1199 (N_1199,N_1101,N_1133);
nor U1200 (N_1200,N_1174,N_1176);
nand U1201 (N_1201,N_1144,N_1142);
nand U1202 (N_1202,N_1167,N_1146);
and U1203 (N_1203,N_1158,N_1169);
nor U1204 (N_1204,N_1185,N_1175);
nand U1205 (N_1205,N_1152,N_1172);
nor U1206 (N_1206,N_1155,N_1179);
and U1207 (N_1207,N_1140,N_1166);
nand U1208 (N_1208,N_1196,N_1153);
nor U1209 (N_1209,N_1143,N_1150);
nor U1210 (N_1210,N_1187,N_1164);
and U1211 (N_1211,N_1178,N_1190);
and U1212 (N_1212,N_1186,N_1168);
and U1213 (N_1213,N_1160,N_1195);
or U1214 (N_1214,N_1171,N_1156);
nand U1215 (N_1215,N_1192,N_1165);
nor U1216 (N_1216,N_1191,N_1159);
nand U1217 (N_1217,N_1177,N_1162);
nand U1218 (N_1218,N_1170,N_1151);
nand U1219 (N_1219,N_1182,N_1154);
or U1220 (N_1220,N_1188,N_1189);
and U1221 (N_1221,N_1157,N_1194);
nor U1222 (N_1222,N_1147,N_1141);
nor U1223 (N_1223,N_1184,N_1173);
nor U1224 (N_1224,N_1161,N_1183);
nor U1225 (N_1225,N_1180,N_1145);
nand U1226 (N_1226,N_1149,N_1198);
and U1227 (N_1227,N_1199,N_1197);
or U1228 (N_1228,N_1181,N_1193);
or U1229 (N_1229,N_1163,N_1148);
nand U1230 (N_1230,N_1162,N_1196);
nand U1231 (N_1231,N_1181,N_1170);
or U1232 (N_1232,N_1158,N_1145);
and U1233 (N_1233,N_1167,N_1171);
or U1234 (N_1234,N_1141,N_1163);
nor U1235 (N_1235,N_1197,N_1151);
or U1236 (N_1236,N_1191,N_1152);
nor U1237 (N_1237,N_1142,N_1161);
nor U1238 (N_1238,N_1197,N_1196);
and U1239 (N_1239,N_1194,N_1160);
or U1240 (N_1240,N_1153,N_1195);
and U1241 (N_1241,N_1180,N_1144);
nor U1242 (N_1242,N_1141,N_1162);
nor U1243 (N_1243,N_1165,N_1163);
nand U1244 (N_1244,N_1152,N_1173);
nor U1245 (N_1245,N_1168,N_1163);
and U1246 (N_1246,N_1199,N_1184);
and U1247 (N_1247,N_1167,N_1168);
or U1248 (N_1248,N_1187,N_1143);
nand U1249 (N_1249,N_1172,N_1146);
and U1250 (N_1250,N_1143,N_1171);
nor U1251 (N_1251,N_1192,N_1149);
and U1252 (N_1252,N_1144,N_1161);
nand U1253 (N_1253,N_1164,N_1192);
or U1254 (N_1254,N_1153,N_1141);
xnor U1255 (N_1255,N_1167,N_1157);
and U1256 (N_1256,N_1178,N_1189);
nor U1257 (N_1257,N_1189,N_1197);
nor U1258 (N_1258,N_1150,N_1172);
and U1259 (N_1259,N_1163,N_1157);
nand U1260 (N_1260,N_1244,N_1221);
or U1261 (N_1261,N_1235,N_1214);
nand U1262 (N_1262,N_1218,N_1200);
and U1263 (N_1263,N_1239,N_1237);
or U1264 (N_1264,N_1228,N_1217);
nand U1265 (N_1265,N_1203,N_1256);
and U1266 (N_1266,N_1232,N_1234);
nor U1267 (N_1267,N_1258,N_1249);
or U1268 (N_1268,N_1250,N_1230);
and U1269 (N_1269,N_1252,N_1253);
nand U1270 (N_1270,N_1255,N_1247);
nand U1271 (N_1271,N_1204,N_1205);
and U1272 (N_1272,N_1248,N_1211);
and U1273 (N_1273,N_1220,N_1225);
and U1274 (N_1274,N_1229,N_1257);
nand U1275 (N_1275,N_1206,N_1216);
or U1276 (N_1276,N_1246,N_1233);
or U1277 (N_1277,N_1242,N_1251);
nor U1278 (N_1278,N_1212,N_1224);
or U1279 (N_1279,N_1213,N_1226);
nand U1280 (N_1280,N_1238,N_1231);
nand U1281 (N_1281,N_1227,N_1259);
or U1282 (N_1282,N_1236,N_1215);
and U1283 (N_1283,N_1219,N_1209);
and U1284 (N_1284,N_1202,N_1222);
and U1285 (N_1285,N_1254,N_1245);
nand U1286 (N_1286,N_1243,N_1207);
nor U1287 (N_1287,N_1208,N_1240);
nand U1288 (N_1288,N_1241,N_1210);
or U1289 (N_1289,N_1201,N_1223);
nor U1290 (N_1290,N_1257,N_1201);
and U1291 (N_1291,N_1205,N_1255);
or U1292 (N_1292,N_1200,N_1230);
nor U1293 (N_1293,N_1213,N_1212);
xor U1294 (N_1294,N_1213,N_1210);
nand U1295 (N_1295,N_1223,N_1247);
nand U1296 (N_1296,N_1214,N_1205);
nor U1297 (N_1297,N_1258,N_1251);
and U1298 (N_1298,N_1218,N_1214);
nor U1299 (N_1299,N_1212,N_1230);
nor U1300 (N_1300,N_1247,N_1200);
xor U1301 (N_1301,N_1251,N_1223);
xor U1302 (N_1302,N_1214,N_1227);
and U1303 (N_1303,N_1203,N_1227);
nand U1304 (N_1304,N_1239,N_1225);
or U1305 (N_1305,N_1233,N_1235);
nor U1306 (N_1306,N_1208,N_1200);
nor U1307 (N_1307,N_1218,N_1242);
and U1308 (N_1308,N_1256,N_1255);
and U1309 (N_1309,N_1241,N_1227);
or U1310 (N_1310,N_1212,N_1217);
and U1311 (N_1311,N_1212,N_1210);
nand U1312 (N_1312,N_1237,N_1238);
and U1313 (N_1313,N_1244,N_1216);
and U1314 (N_1314,N_1249,N_1243);
nand U1315 (N_1315,N_1204,N_1213);
nand U1316 (N_1316,N_1246,N_1240);
nor U1317 (N_1317,N_1217,N_1249);
nand U1318 (N_1318,N_1209,N_1202);
nor U1319 (N_1319,N_1236,N_1202);
nor U1320 (N_1320,N_1272,N_1263);
or U1321 (N_1321,N_1282,N_1313);
nor U1322 (N_1322,N_1315,N_1281);
or U1323 (N_1323,N_1309,N_1308);
nand U1324 (N_1324,N_1290,N_1285);
nand U1325 (N_1325,N_1260,N_1318);
or U1326 (N_1326,N_1261,N_1298);
or U1327 (N_1327,N_1311,N_1304);
or U1328 (N_1328,N_1288,N_1264);
and U1329 (N_1329,N_1284,N_1294);
and U1330 (N_1330,N_1303,N_1317);
or U1331 (N_1331,N_1277,N_1278);
and U1332 (N_1332,N_1275,N_1283);
nor U1333 (N_1333,N_1269,N_1287);
nand U1334 (N_1334,N_1297,N_1301);
nand U1335 (N_1335,N_1268,N_1302);
and U1336 (N_1336,N_1271,N_1310);
and U1337 (N_1337,N_1274,N_1312);
nand U1338 (N_1338,N_1279,N_1295);
nor U1339 (N_1339,N_1280,N_1292);
nand U1340 (N_1340,N_1296,N_1299);
and U1341 (N_1341,N_1289,N_1276);
nor U1342 (N_1342,N_1306,N_1305);
or U1343 (N_1343,N_1273,N_1316);
nor U1344 (N_1344,N_1286,N_1319);
and U1345 (N_1345,N_1291,N_1266);
nor U1346 (N_1346,N_1314,N_1270);
nor U1347 (N_1347,N_1267,N_1265);
nand U1348 (N_1348,N_1300,N_1307);
and U1349 (N_1349,N_1293,N_1262);
and U1350 (N_1350,N_1260,N_1310);
or U1351 (N_1351,N_1303,N_1275);
or U1352 (N_1352,N_1281,N_1285);
nand U1353 (N_1353,N_1295,N_1280);
nand U1354 (N_1354,N_1284,N_1267);
nand U1355 (N_1355,N_1311,N_1276);
nor U1356 (N_1356,N_1290,N_1264);
nand U1357 (N_1357,N_1280,N_1310);
and U1358 (N_1358,N_1295,N_1260);
nand U1359 (N_1359,N_1308,N_1275);
or U1360 (N_1360,N_1296,N_1304);
nand U1361 (N_1361,N_1295,N_1275);
nand U1362 (N_1362,N_1260,N_1282);
nand U1363 (N_1363,N_1296,N_1267);
nor U1364 (N_1364,N_1274,N_1277);
nand U1365 (N_1365,N_1307,N_1260);
or U1366 (N_1366,N_1297,N_1282);
nor U1367 (N_1367,N_1289,N_1307);
nand U1368 (N_1368,N_1283,N_1291);
or U1369 (N_1369,N_1317,N_1280);
nand U1370 (N_1370,N_1266,N_1316);
nor U1371 (N_1371,N_1315,N_1294);
and U1372 (N_1372,N_1289,N_1300);
or U1373 (N_1373,N_1286,N_1312);
or U1374 (N_1374,N_1318,N_1287);
or U1375 (N_1375,N_1265,N_1311);
and U1376 (N_1376,N_1260,N_1268);
xnor U1377 (N_1377,N_1307,N_1275);
nor U1378 (N_1378,N_1306,N_1275);
nand U1379 (N_1379,N_1289,N_1297);
nand U1380 (N_1380,N_1322,N_1336);
nor U1381 (N_1381,N_1373,N_1356);
or U1382 (N_1382,N_1321,N_1370);
and U1383 (N_1383,N_1371,N_1330);
nand U1384 (N_1384,N_1365,N_1329);
nor U1385 (N_1385,N_1372,N_1337);
and U1386 (N_1386,N_1328,N_1362);
nor U1387 (N_1387,N_1351,N_1376);
nor U1388 (N_1388,N_1338,N_1353);
or U1389 (N_1389,N_1320,N_1345);
nor U1390 (N_1390,N_1377,N_1346);
nand U1391 (N_1391,N_1333,N_1368);
or U1392 (N_1392,N_1361,N_1375);
and U1393 (N_1393,N_1359,N_1360);
or U1394 (N_1394,N_1323,N_1378);
nor U1395 (N_1395,N_1364,N_1354);
nor U1396 (N_1396,N_1357,N_1342);
nor U1397 (N_1397,N_1340,N_1349);
nor U1398 (N_1398,N_1369,N_1326);
and U1399 (N_1399,N_1355,N_1348);
and U1400 (N_1400,N_1344,N_1339);
nor U1401 (N_1401,N_1341,N_1367);
or U1402 (N_1402,N_1343,N_1324);
nand U1403 (N_1403,N_1366,N_1327);
and U1404 (N_1404,N_1363,N_1374);
or U1405 (N_1405,N_1335,N_1350);
nand U1406 (N_1406,N_1352,N_1379);
and U1407 (N_1407,N_1358,N_1347);
or U1408 (N_1408,N_1331,N_1334);
and U1409 (N_1409,N_1332,N_1325);
or U1410 (N_1410,N_1366,N_1360);
nor U1411 (N_1411,N_1321,N_1331);
and U1412 (N_1412,N_1320,N_1370);
and U1413 (N_1413,N_1333,N_1326);
and U1414 (N_1414,N_1370,N_1337);
or U1415 (N_1415,N_1333,N_1377);
and U1416 (N_1416,N_1366,N_1353);
and U1417 (N_1417,N_1369,N_1348);
xnor U1418 (N_1418,N_1339,N_1355);
nor U1419 (N_1419,N_1375,N_1322);
and U1420 (N_1420,N_1321,N_1376);
or U1421 (N_1421,N_1326,N_1321);
nand U1422 (N_1422,N_1368,N_1369);
and U1423 (N_1423,N_1340,N_1323);
nand U1424 (N_1424,N_1377,N_1353);
nand U1425 (N_1425,N_1326,N_1352);
or U1426 (N_1426,N_1371,N_1362);
and U1427 (N_1427,N_1320,N_1321);
or U1428 (N_1428,N_1349,N_1343);
or U1429 (N_1429,N_1372,N_1340);
nand U1430 (N_1430,N_1358,N_1333);
or U1431 (N_1431,N_1371,N_1370);
nand U1432 (N_1432,N_1353,N_1341);
nor U1433 (N_1433,N_1339,N_1333);
nand U1434 (N_1434,N_1331,N_1376);
nand U1435 (N_1435,N_1348,N_1332);
and U1436 (N_1436,N_1345,N_1330);
nor U1437 (N_1437,N_1340,N_1337);
nor U1438 (N_1438,N_1365,N_1324);
nand U1439 (N_1439,N_1369,N_1358);
nor U1440 (N_1440,N_1393,N_1430);
nor U1441 (N_1441,N_1403,N_1406);
or U1442 (N_1442,N_1410,N_1391);
or U1443 (N_1443,N_1383,N_1436);
or U1444 (N_1444,N_1419,N_1392);
nor U1445 (N_1445,N_1427,N_1416);
and U1446 (N_1446,N_1401,N_1396);
and U1447 (N_1447,N_1380,N_1404);
and U1448 (N_1448,N_1386,N_1424);
and U1449 (N_1449,N_1429,N_1397);
and U1450 (N_1450,N_1411,N_1390);
and U1451 (N_1451,N_1435,N_1382);
xnor U1452 (N_1452,N_1398,N_1413);
and U1453 (N_1453,N_1431,N_1414);
nand U1454 (N_1454,N_1417,N_1438);
nor U1455 (N_1455,N_1409,N_1415);
nor U1456 (N_1456,N_1408,N_1381);
nor U1457 (N_1457,N_1400,N_1420);
nor U1458 (N_1458,N_1402,N_1388);
and U1459 (N_1459,N_1394,N_1422);
and U1460 (N_1460,N_1425,N_1426);
and U1461 (N_1461,N_1433,N_1421);
or U1462 (N_1462,N_1405,N_1395);
or U1463 (N_1463,N_1423,N_1439);
nand U1464 (N_1464,N_1399,N_1437);
or U1465 (N_1465,N_1418,N_1412);
nand U1466 (N_1466,N_1432,N_1389);
or U1467 (N_1467,N_1428,N_1385);
nor U1468 (N_1468,N_1407,N_1384);
and U1469 (N_1469,N_1434,N_1387);
nand U1470 (N_1470,N_1385,N_1409);
nand U1471 (N_1471,N_1427,N_1437);
nor U1472 (N_1472,N_1424,N_1402);
nor U1473 (N_1473,N_1406,N_1426);
or U1474 (N_1474,N_1402,N_1414);
and U1475 (N_1475,N_1411,N_1429);
or U1476 (N_1476,N_1431,N_1401);
or U1477 (N_1477,N_1411,N_1384);
and U1478 (N_1478,N_1388,N_1436);
or U1479 (N_1479,N_1401,N_1382);
nor U1480 (N_1480,N_1435,N_1390);
and U1481 (N_1481,N_1407,N_1393);
or U1482 (N_1482,N_1383,N_1426);
nor U1483 (N_1483,N_1403,N_1388);
and U1484 (N_1484,N_1412,N_1385);
or U1485 (N_1485,N_1436,N_1429);
or U1486 (N_1486,N_1385,N_1433);
nand U1487 (N_1487,N_1402,N_1438);
nand U1488 (N_1488,N_1402,N_1423);
or U1489 (N_1489,N_1417,N_1428);
and U1490 (N_1490,N_1422,N_1390);
or U1491 (N_1491,N_1383,N_1384);
or U1492 (N_1492,N_1431,N_1426);
nand U1493 (N_1493,N_1419,N_1383);
and U1494 (N_1494,N_1409,N_1425);
nand U1495 (N_1495,N_1431,N_1404);
nor U1496 (N_1496,N_1437,N_1438);
nor U1497 (N_1497,N_1389,N_1422);
and U1498 (N_1498,N_1403,N_1381);
nor U1499 (N_1499,N_1403,N_1382);
or U1500 (N_1500,N_1446,N_1463);
or U1501 (N_1501,N_1491,N_1449);
and U1502 (N_1502,N_1483,N_1471);
or U1503 (N_1503,N_1440,N_1473);
and U1504 (N_1504,N_1482,N_1445);
and U1505 (N_1505,N_1443,N_1499);
or U1506 (N_1506,N_1472,N_1464);
nand U1507 (N_1507,N_1496,N_1469);
or U1508 (N_1508,N_1451,N_1455);
and U1509 (N_1509,N_1476,N_1470);
nand U1510 (N_1510,N_1460,N_1494);
or U1511 (N_1511,N_1484,N_1444);
nor U1512 (N_1512,N_1493,N_1467);
nor U1513 (N_1513,N_1480,N_1450);
nor U1514 (N_1514,N_1497,N_1490);
nor U1515 (N_1515,N_1452,N_1475);
or U1516 (N_1516,N_1489,N_1454);
nor U1517 (N_1517,N_1461,N_1481);
or U1518 (N_1518,N_1457,N_1459);
nor U1519 (N_1519,N_1453,N_1486);
nor U1520 (N_1520,N_1442,N_1487);
or U1521 (N_1521,N_1441,N_1492);
and U1522 (N_1522,N_1498,N_1485);
and U1523 (N_1523,N_1479,N_1462);
or U1524 (N_1524,N_1456,N_1488);
or U1525 (N_1525,N_1465,N_1448);
and U1526 (N_1526,N_1447,N_1466);
nor U1527 (N_1527,N_1495,N_1458);
and U1528 (N_1528,N_1477,N_1468);
nand U1529 (N_1529,N_1474,N_1478);
or U1530 (N_1530,N_1476,N_1469);
nor U1531 (N_1531,N_1452,N_1488);
or U1532 (N_1532,N_1444,N_1459);
nor U1533 (N_1533,N_1445,N_1492);
or U1534 (N_1534,N_1445,N_1476);
nor U1535 (N_1535,N_1447,N_1491);
nor U1536 (N_1536,N_1472,N_1473);
nand U1537 (N_1537,N_1486,N_1493);
nor U1538 (N_1538,N_1459,N_1470);
nor U1539 (N_1539,N_1490,N_1441);
nor U1540 (N_1540,N_1464,N_1467);
nor U1541 (N_1541,N_1496,N_1471);
nor U1542 (N_1542,N_1448,N_1482);
or U1543 (N_1543,N_1462,N_1483);
and U1544 (N_1544,N_1496,N_1458);
and U1545 (N_1545,N_1472,N_1444);
and U1546 (N_1546,N_1452,N_1494);
or U1547 (N_1547,N_1463,N_1493);
nor U1548 (N_1548,N_1460,N_1468);
or U1549 (N_1549,N_1468,N_1464);
and U1550 (N_1550,N_1466,N_1455);
nand U1551 (N_1551,N_1460,N_1463);
nand U1552 (N_1552,N_1481,N_1456);
nor U1553 (N_1553,N_1485,N_1461);
nor U1554 (N_1554,N_1443,N_1446);
or U1555 (N_1555,N_1495,N_1453);
and U1556 (N_1556,N_1451,N_1476);
nor U1557 (N_1557,N_1489,N_1452);
and U1558 (N_1558,N_1456,N_1468);
nor U1559 (N_1559,N_1499,N_1457);
and U1560 (N_1560,N_1514,N_1545);
and U1561 (N_1561,N_1526,N_1551);
or U1562 (N_1562,N_1516,N_1555);
nand U1563 (N_1563,N_1559,N_1506);
nor U1564 (N_1564,N_1517,N_1557);
nor U1565 (N_1565,N_1501,N_1534);
nand U1566 (N_1566,N_1513,N_1548);
nor U1567 (N_1567,N_1547,N_1535);
and U1568 (N_1568,N_1509,N_1500);
and U1569 (N_1569,N_1524,N_1540);
or U1570 (N_1570,N_1556,N_1515);
nand U1571 (N_1571,N_1537,N_1507);
or U1572 (N_1572,N_1508,N_1522);
nor U1573 (N_1573,N_1532,N_1527);
nor U1574 (N_1574,N_1530,N_1546);
nand U1575 (N_1575,N_1531,N_1519);
or U1576 (N_1576,N_1521,N_1505);
nand U1577 (N_1577,N_1549,N_1533);
and U1578 (N_1578,N_1511,N_1529);
or U1579 (N_1579,N_1503,N_1512);
nand U1580 (N_1580,N_1542,N_1525);
nor U1581 (N_1581,N_1536,N_1554);
and U1582 (N_1582,N_1550,N_1504);
nor U1583 (N_1583,N_1510,N_1543);
or U1584 (N_1584,N_1502,N_1541);
or U1585 (N_1585,N_1539,N_1544);
nand U1586 (N_1586,N_1528,N_1518);
or U1587 (N_1587,N_1538,N_1520);
nor U1588 (N_1588,N_1523,N_1552);
or U1589 (N_1589,N_1553,N_1558);
nand U1590 (N_1590,N_1516,N_1532);
and U1591 (N_1591,N_1527,N_1551);
and U1592 (N_1592,N_1533,N_1532);
and U1593 (N_1593,N_1521,N_1500);
and U1594 (N_1594,N_1525,N_1535);
and U1595 (N_1595,N_1540,N_1518);
and U1596 (N_1596,N_1532,N_1534);
or U1597 (N_1597,N_1519,N_1557);
or U1598 (N_1598,N_1510,N_1523);
nand U1599 (N_1599,N_1547,N_1537);
nor U1600 (N_1600,N_1550,N_1548);
and U1601 (N_1601,N_1505,N_1523);
nor U1602 (N_1602,N_1508,N_1550);
or U1603 (N_1603,N_1558,N_1529);
nor U1604 (N_1604,N_1556,N_1501);
and U1605 (N_1605,N_1514,N_1532);
or U1606 (N_1606,N_1532,N_1501);
nand U1607 (N_1607,N_1545,N_1546);
nor U1608 (N_1608,N_1526,N_1505);
nand U1609 (N_1609,N_1526,N_1544);
nand U1610 (N_1610,N_1536,N_1548);
or U1611 (N_1611,N_1524,N_1539);
or U1612 (N_1612,N_1529,N_1512);
or U1613 (N_1613,N_1524,N_1559);
nor U1614 (N_1614,N_1537,N_1503);
or U1615 (N_1615,N_1507,N_1540);
and U1616 (N_1616,N_1516,N_1551);
and U1617 (N_1617,N_1559,N_1550);
nor U1618 (N_1618,N_1558,N_1544);
and U1619 (N_1619,N_1556,N_1502);
and U1620 (N_1620,N_1584,N_1601);
nand U1621 (N_1621,N_1609,N_1565);
or U1622 (N_1622,N_1599,N_1572);
nand U1623 (N_1623,N_1593,N_1588);
nand U1624 (N_1624,N_1560,N_1606);
nand U1625 (N_1625,N_1610,N_1573);
or U1626 (N_1626,N_1583,N_1585);
nand U1627 (N_1627,N_1600,N_1611);
or U1628 (N_1628,N_1619,N_1587);
nand U1629 (N_1629,N_1581,N_1578);
or U1630 (N_1630,N_1608,N_1597);
nand U1631 (N_1631,N_1615,N_1566);
nand U1632 (N_1632,N_1614,N_1579);
and U1633 (N_1633,N_1595,N_1604);
nand U1634 (N_1634,N_1602,N_1562);
or U1635 (N_1635,N_1591,N_1603);
and U1636 (N_1636,N_1577,N_1612);
xnor U1637 (N_1637,N_1605,N_1618);
nand U1638 (N_1638,N_1567,N_1613);
nor U1639 (N_1639,N_1568,N_1589);
and U1640 (N_1640,N_1576,N_1586);
nor U1641 (N_1641,N_1582,N_1570);
nand U1642 (N_1642,N_1594,N_1575);
or U1643 (N_1643,N_1580,N_1571);
nand U1644 (N_1644,N_1592,N_1616);
nor U1645 (N_1645,N_1569,N_1617);
or U1646 (N_1646,N_1596,N_1590);
nand U1647 (N_1647,N_1598,N_1561);
nor U1648 (N_1648,N_1564,N_1607);
nand U1649 (N_1649,N_1574,N_1563);
and U1650 (N_1650,N_1614,N_1561);
nand U1651 (N_1651,N_1563,N_1576);
xor U1652 (N_1652,N_1618,N_1606);
and U1653 (N_1653,N_1607,N_1619);
nor U1654 (N_1654,N_1567,N_1592);
and U1655 (N_1655,N_1590,N_1595);
and U1656 (N_1656,N_1596,N_1589);
xnor U1657 (N_1657,N_1561,N_1584);
or U1658 (N_1658,N_1578,N_1590);
and U1659 (N_1659,N_1603,N_1576);
and U1660 (N_1660,N_1581,N_1592);
and U1661 (N_1661,N_1568,N_1619);
and U1662 (N_1662,N_1567,N_1590);
or U1663 (N_1663,N_1565,N_1589);
nor U1664 (N_1664,N_1618,N_1573);
or U1665 (N_1665,N_1582,N_1599);
nand U1666 (N_1666,N_1618,N_1569);
nand U1667 (N_1667,N_1589,N_1582);
nand U1668 (N_1668,N_1615,N_1613);
and U1669 (N_1669,N_1570,N_1564);
nand U1670 (N_1670,N_1585,N_1606);
or U1671 (N_1671,N_1607,N_1585);
nor U1672 (N_1672,N_1563,N_1590);
and U1673 (N_1673,N_1580,N_1605);
nand U1674 (N_1674,N_1614,N_1598);
nor U1675 (N_1675,N_1616,N_1564);
nand U1676 (N_1676,N_1597,N_1615);
or U1677 (N_1677,N_1570,N_1602);
nand U1678 (N_1678,N_1574,N_1568);
nand U1679 (N_1679,N_1605,N_1598);
nand U1680 (N_1680,N_1656,N_1620);
nand U1681 (N_1681,N_1643,N_1634);
nand U1682 (N_1682,N_1631,N_1653);
or U1683 (N_1683,N_1677,N_1622);
and U1684 (N_1684,N_1675,N_1669);
nand U1685 (N_1685,N_1654,N_1674);
or U1686 (N_1686,N_1660,N_1679);
or U1687 (N_1687,N_1666,N_1647);
or U1688 (N_1688,N_1630,N_1645);
nor U1689 (N_1689,N_1649,N_1662);
nor U1690 (N_1690,N_1627,N_1667);
or U1691 (N_1691,N_1638,N_1658);
nor U1692 (N_1692,N_1624,N_1642);
and U1693 (N_1693,N_1621,N_1663);
xnor U1694 (N_1694,N_1668,N_1665);
or U1695 (N_1695,N_1637,N_1646);
nor U1696 (N_1696,N_1661,N_1664);
nand U1697 (N_1697,N_1671,N_1676);
and U1698 (N_1698,N_1648,N_1639);
nor U1699 (N_1699,N_1623,N_1626);
and U1700 (N_1700,N_1628,N_1629);
nor U1701 (N_1701,N_1672,N_1673);
nand U1702 (N_1702,N_1657,N_1633);
nor U1703 (N_1703,N_1651,N_1655);
xnor U1704 (N_1704,N_1625,N_1644);
or U1705 (N_1705,N_1670,N_1636);
or U1706 (N_1706,N_1640,N_1650);
nand U1707 (N_1707,N_1641,N_1678);
or U1708 (N_1708,N_1632,N_1659);
and U1709 (N_1709,N_1652,N_1635);
nand U1710 (N_1710,N_1653,N_1637);
or U1711 (N_1711,N_1663,N_1674);
and U1712 (N_1712,N_1652,N_1632);
and U1713 (N_1713,N_1646,N_1664);
and U1714 (N_1714,N_1630,N_1662);
nand U1715 (N_1715,N_1656,N_1647);
nand U1716 (N_1716,N_1672,N_1634);
nand U1717 (N_1717,N_1677,N_1672);
and U1718 (N_1718,N_1670,N_1668);
nand U1719 (N_1719,N_1633,N_1647);
nand U1720 (N_1720,N_1661,N_1632);
or U1721 (N_1721,N_1674,N_1643);
or U1722 (N_1722,N_1666,N_1658);
and U1723 (N_1723,N_1643,N_1657);
and U1724 (N_1724,N_1647,N_1645);
or U1725 (N_1725,N_1669,N_1679);
and U1726 (N_1726,N_1665,N_1621);
nor U1727 (N_1727,N_1648,N_1678);
or U1728 (N_1728,N_1668,N_1633);
and U1729 (N_1729,N_1666,N_1664);
nor U1730 (N_1730,N_1658,N_1663);
nand U1731 (N_1731,N_1640,N_1635);
and U1732 (N_1732,N_1672,N_1642);
or U1733 (N_1733,N_1661,N_1628);
or U1734 (N_1734,N_1674,N_1679);
nor U1735 (N_1735,N_1652,N_1671);
nand U1736 (N_1736,N_1677,N_1663);
and U1737 (N_1737,N_1645,N_1644);
nand U1738 (N_1738,N_1674,N_1676);
or U1739 (N_1739,N_1655,N_1671);
nand U1740 (N_1740,N_1736,N_1691);
nand U1741 (N_1741,N_1715,N_1725);
nor U1742 (N_1742,N_1732,N_1720);
nand U1743 (N_1743,N_1684,N_1738);
and U1744 (N_1744,N_1708,N_1681);
nand U1745 (N_1745,N_1717,N_1710);
or U1746 (N_1746,N_1734,N_1707);
or U1747 (N_1747,N_1711,N_1696);
and U1748 (N_1748,N_1689,N_1705);
and U1749 (N_1749,N_1735,N_1694);
and U1750 (N_1750,N_1698,N_1730);
nor U1751 (N_1751,N_1739,N_1712);
nor U1752 (N_1752,N_1722,N_1695);
nor U1753 (N_1753,N_1693,N_1702);
nand U1754 (N_1754,N_1718,N_1729);
nand U1755 (N_1755,N_1706,N_1703);
and U1756 (N_1756,N_1716,N_1680);
nand U1757 (N_1757,N_1688,N_1713);
or U1758 (N_1758,N_1683,N_1701);
nor U1759 (N_1759,N_1686,N_1733);
nand U1760 (N_1760,N_1731,N_1699);
nor U1761 (N_1761,N_1709,N_1687);
nor U1762 (N_1762,N_1690,N_1728);
nand U1763 (N_1763,N_1723,N_1714);
and U1764 (N_1764,N_1685,N_1737);
and U1765 (N_1765,N_1704,N_1700);
or U1766 (N_1766,N_1726,N_1724);
xor U1767 (N_1767,N_1727,N_1697);
and U1768 (N_1768,N_1692,N_1721);
nand U1769 (N_1769,N_1719,N_1682);
nand U1770 (N_1770,N_1730,N_1727);
or U1771 (N_1771,N_1682,N_1721);
or U1772 (N_1772,N_1729,N_1736);
nand U1773 (N_1773,N_1730,N_1687);
or U1774 (N_1774,N_1726,N_1704);
and U1775 (N_1775,N_1689,N_1723);
xor U1776 (N_1776,N_1712,N_1727);
or U1777 (N_1777,N_1684,N_1734);
or U1778 (N_1778,N_1704,N_1718);
and U1779 (N_1779,N_1708,N_1720);
and U1780 (N_1780,N_1698,N_1734);
and U1781 (N_1781,N_1724,N_1692);
and U1782 (N_1782,N_1726,N_1733);
and U1783 (N_1783,N_1728,N_1703);
nand U1784 (N_1784,N_1722,N_1731);
and U1785 (N_1785,N_1722,N_1703);
nor U1786 (N_1786,N_1696,N_1701);
nor U1787 (N_1787,N_1697,N_1724);
or U1788 (N_1788,N_1731,N_1700);
xnor U1789 (N_1789,N_1695,N_1714);
and U1790 (N_1790,N_1720,N_1731);
nand U1791 (N_1791,N_1715,N_1739);
nor U1792 (N_1792,N_1726,N_1700);
xor U1793 (N_1793,N_1724,N_1737);
nor U1794 (N_1794,N_1716,N_1682);
nor U1795 (N_1795,N_1736,N_1697);
nor U1796 (N_1796,N_1711,N_1695);
nor U1797 (N_1797,N_1711,N_1697);
nand U1798 (N_1798,N_1699,N_1681);
and U1799 (N_1799,N_1681,N_1716);
or U1800 (N_1800,N_1779,N_1786);
xnor U1801 (N_1801,N_1798,N_1754);
and U1802 (N_1802,N_1796,N_1764);
nand U1803 (N_1803,N_1768,N_1771);
nand U1804 (N_1804,N_1741,N_1746);
and U1805 (N_1805,N_1763,N_1769);
or U1806 (N_1806,N_1776,N_1783);
or U1807 (N_1807,N_1756,N_1793);
nand U1808 (N_1808,N_1745,N_1753);
nand U1809 (N_1809,N_1792,N_1789);
and U1810 (N_1810,N_1770,N_1759);
nand U1811 (N_1811,N_1740,N_1766);
nand U1812 (N_1812,N_1784,N_1790);
nand U1813 (N_1813,N_1744,N_1762);
nor U1814 (N_1814,N_1765,N_1760);
nor U1815 (N_1815,N_1794,N_1799);
nor U1816 (N_1816,N_1747,N_1780);
nor U1817 (N_1817,N_1772,N_1787);
and U1818 (N_1818,N_1755,N_1775);
nand U1819 (N_1819,N_1742,N_1797);
and U1820 (N_1820,N_1752,N_1750);
or U1821 (N_1821,N_1761,N_1743);
or U1822 (N_1822,N_1785,N_1767);
and U1823 (N_1823,N_1774,N_1751);
nor U1824 (N_1824,N_1773,N_1757);
nor U1825 (N_1825,N_1777,N_1749);
and U1826 (N_1826,N_1758,N_1781);
nor U1827 (N_1827,N_1782,N_1748);
or U1828 (N_1828,N_1778,N_1795);
and U1829 (N_1829,N_1791,N_1788);
nor U1830 (N_1830,N_1773,N_1793);
nor U1831 (N_1831,N_1782,N_1774);
nand U1832 (N_1832,N_1764,N_1772);
nor U1833 (N_1833,N_1779,N_1798);
nand U1834 (N_1834,N_1775,N_1778);
and U1835 (N_1835,N_1790,N_1797);
or U1836 (N_1836,N_1777,N_1791);
and U1837 (N_1837,N_1788,N_1771);
nand U1838 (N_1838,N_1774,N_1797);
or U1839 (N_1839,N_1768,N_1794);
nor U1840 (N_1840,N_1768,N_1753);
and U1841 (N_1841,N_1750,N_1757);
nor U1842 (N_1842,N_1785,N_1793);
or U1843 (N_1843,N_1799,N_1796);
nand U1844 (N_1844,N_1780,N_1764);
nor U1845 (N_1845,N_1798,N_1780);
or U1846 (N_1846,N_1748,N_1757);
nand U1847 (N_1847,N_1789,N_1797);
or U1848 (N_1848,N_1768,N_1750);
or U1849 (N_1849,N_1778,N_1787);
nor U1850 (N_1850,N_1776,N_1782);
nor U1851 (N_1851,N_1797,N_1747);
and U1852 (N_1852,N_1788,N_1754);
nor U1853 (N_1853,N_1751,N_1783);
nor U1854 (N_1854,N_1789,N_1793);
nand U1855 (N_1855,N_1747,N_1783);
and U1856 (N_1856,N_1769,N_1743);
nor U1857 (N_1857,N_1765,N_1751);
or U1858 (N_1858,N_1763,N_1742);
nand U1859 (N_1859,N_1748,N_1761);
nand U1860 (N_1860,N_1839,N_1818);
or U1861 (N_1861,N_1808,N_1851);
nand U1862 (N_1862,N_1829,N_1809);
and U1863 (N_1863,N_1811,N_1859);
and U1864 (N_1864,N_1823,N_1837);
nor U1865 (N_1865,N_1845,N_1848);
nand U1866 (N_1866,N_1831,N_1840);
nor U1867 (N_1867,N_1803,N_1801);
nand U1868 (N_1868,N_1821,N_1826);
or U1869 (N_1869,N_1853,N_1836);
or U1870 (N_1870,N_1832,N_1856);
xnor U1871 (N_1871,N_1835,N_1838);
and U1872 (N_1872,N_1842,N_1804);
or U1873 (N_1873,N_1820,N_1841);
and U1874 (N_1874,N_1817,N_1858);
and U1875 (N_1875,N_1852,N_1815);
or U1876 (N_1876,N_1847,N_1844);
and U1877 (N_1877,N_1800,N_1816);
nand U1878 (N_1878,N_1843,N_1830);
nor U1879 (N_1879,N_1805,N_1806);
or U1880 (N_1880,N_1850,N_1834);
nor U1881 (N_1881,N_1828,N_1812);
xor U1882 (N_1882,N_1822,N_1846);
nand U1883 (N_1883,N_1827,N_1824);
nand U1884 (N_1884,N_1807,N_1825);
nand U1885 (N_1885,N_1854,N_1814);
nand U1886 (N_1886,N_1819,N_1802);
or U1887 (N_1887,N_1857,N_1813);
and U1888 (N_1888,N_1849,N_1810);
nand U1889 (N_1889,N_1833,N_1855);
nor U1890 (N_1890,N_1801,N_1808);
or U1891 (N_1891,N_1842,N_1807);
or U1892 (N_1892,N_1833,N_1847);
and U1893 (N_1893,N_1830,N_1804);
or U1894 (N_1894,N_1838,N_1811);
nor U1895 (N_1895,N_1803,N_1826);
or U1896 (N_1896,N_1852,N_1818);
or U1897 (N_1897,N_1804,N_1858);
nor U1898 (N_1898,N_1857,N_1846);
nand U1899 (N_1899,N_1825,N_1814);
nand U1900 (N_1900,N_1852,N_1830);
nand U1901 (N_1901,N_1820,N_1840);
or U1902 (N_1902,N_1835,N_1855);
and U1903 (N_1903,N_1853,N_1848);
and U1904 (N_1904,N_1809,N_1812);
nand U1905 (N_1905,N_1824,N_1832);
xnor U1906 (N_1906,N_1859,N_1808);
nand U1907 (N_1907,N_1835,N_1841);
or U1908 (N_1908,N_1800,N_1826);
and U1909 (N_1909,N_1828,N_1843);
nand U1910 (N_1910,N_1800,N_1810);
and U1911 (N_1911,N_1828,N_1824);
and U1912 (N_1912,N_1812,N_1831);
nor U1913 (N_1913,N_1820,N_1817);
or U1914 (N_1914,N_1846,N_1807);
and U1915 (N_1915,N_1832,N_1815);
or U1916 (N_1916,N_1846,N_1808);
or U1917 (N_1917,N_1815,N_1828);
nor U1918 (N_1918,N_1804,N_1854);
nor U1919 (N_1919,N_1828,N_1836);
or U1920 (N_1920,N_1916,N_1875);
nor U1921 (N_1921,N_1880,N_1897);
or U1922 (N_1922,N_1877,N_1884);
and U1923 (N_1923,N_1870,N_1905);
and U1924 (N_1924,N_1886,N_1900);
and U1925 (N_1925,N_1919,N_1908);
or U1926 (N_1926,N_1878,N_1874);
and U1927 (N_1927,N_1862,N_1860);
nand U1928 (N_1928,N_1881,N_1868);
and U1929 (N_1929,N_1901,N_1918);
and U1930 (N_1930,N_1912,N_1914);
and U1931 (N_1931,N_1873,N_1865);
nand U1932 (N_1932,N_1896,N_1871);
or U1933 (N_1933,N_1885,N_1893);
nor U1934 (N_1934,N_1890,N_1902);
and U1935 (N_1935,N_1913,N_1904);
nor U1936 (N_1936,N_1907,N_1869);
and U1937 (N_1937,N_1888,N_1899);
nor U1938 (N_1938,N_1887,N_1898);
and U1939 (N_1939,N_1867,N_1872);
or U1940 (N_1940,N_1889,N_1861);
and U1941 (N_1941,N_1894,N_1917);
nand U1942 (N_1942,N_1882,N_1891);
nand U1943 (N_1943,N_1864,N_1909);
nand U1944 (N_1944,N_1915,N_1876);
or U1945 (N_1945,N_1863,N_1906);
or U1946 (N_1946,N_1911,N_1879);
or U1947 (N_1947,N_1903,N_1866);
nand U1948 (N_1948,N_1892,N_1883);
nor U1949 (N_1949,N_1895,N_1910);
nand U1950 (N_1950,N_1893,N_1918);
and U1951 (N_1951,N_1889,N_1860);
nor U1952 (N_1952,N_1913,N_1865);
nor U1953 (N_1953,N_1892,N_1865);
and U1954 (N_1954,N_1866,N_1874);
nor U1955 (N_1955,N_1919,N_1879);
or U1956 (N_1956,N_1889,N_1919);
nor U1957 (N_1957,N_1914,N_1902);
and U1958 (N_1958,N_1889,N_1870);
nor U1959 (N_1959,N_1904,N_1860);
or U1960 (N_1960,N_1891,N_1902);
nand U1961 (N_1961,N_1878,N_1877);
nor U1962 (N_1962,N_1899,N_1866);
or U1963 (N_1963,N_1894,N_1878);
and U1964 (N_1964,N_1874,N_1865);
nor U1965 (N_1965,N_1902,N_1893);
and U1966 (N_1966,N_1875,N_1912);
and U1967 (N_1967,N_1907,N_1888);
nand U1968 (N_1968,N_1863,N_1882);
and U1969 (N_1969,N_1914,N_1898);
or U1970 (N_1970,N_1889,N_1904);
nand U1971 (N_1971,N_1888,N_1904);
nand U1972 (N_1972,N_1916,N_1890);
xnor U1973 (N_1973,N_1876,N_1880);
and U1974 (N_1974,N_1891,N_1899);
nor U1975 (N_1975,N_1861,N_1886);
and U1976 (N_1976,N_1873,N_1877);
nand U1977 (N_1977,N_1883,N_1917);
nor U1978 (N_1978,N_1894,N_1914);
or U1979 (N_1979,N_1896,N_1865);
nor U1980 (N_1980,N_1979,N_1921);
nor U1981 (N_1981,N_1932,N_1956);
and U1982 (N_1982,N_1952,N_1945);
and U1983 (N_1983,N_1939,N_1947);
and U1984 (N_1984,N_1976,N_1964);
and U1985 (N_1985,N_1963,N_1924);
nor U1986 (N_1986,N_1977,N_1950);
nand U1987 (N_1987,N_1955,N_1958);
nor U1988 (N_1988,N_1975,N_1936);
and U1989 (N_1989,N_1941,N_1974);
nand U1990 (N_1990,N_1920,N_1929);
nand U1991 (N_1991,N_1962,N_1930);
nor U1992 (N_1992,N_1967,N_1948);
nand U1993 (N_1993,N_1938,N_1926);
nand U1994 (N_1994,N_1933,N_1953);
or U1995 (N_1995,N_1934,N_1925);
nand U1996 (N_1996,N_1970,N_1972);
nand U1997 (N_1997,N_1943,N_1968);
nand U1998 (N_1998,N_1935,N_1960);
or U1999 (N_1999,N_1942,N_1922);
nor U2000 (N_2000,N_1951,N_1965);
nand U2001 (N_2001,N_1928,N_1966);
or U2002 (N_2002,N_1931,N_1954);
nor U2003 (N_2003,N_1971,N_1937);
and U2004 (N_2004,N_1944,N_1949);
and U2005 (N_2005,N_1946,N_1973);
and U2006 (N_2006,N_1969,N_1978);
nor U2007 (N_2007,N_1957,N_1940);
and U2008 (N_2008,N_1959,N_1927);
or U2009 (N_2009,N_1961,N_1923);
nor U2010 (N_2010,N_1953,N_1937);
nor U2011 (N_2011,N_1964,N_1968);
nand U2012 (N_2012,N_1920,N_1931);
and U2013 (N_2013,N_1920,N_1955);
nand U2014 (N_2014,N_1955,N_1952);
and U2015 (N_2015,N_1944,N_1927);
and U2016 (N_2016,N_1942,N_1964);
and U2017 (N_2017,N_1928,N_1962);
or U2018 (N_2018,N_1951,N_1963);
or U2019 (N_2019,N_1965,N_1968);
or U2020 (N_2020,N_1952,N_1933);
or U2021 (N_2021,N_1944,N_1971);
nand U2022 (N_2022,N_1972,N_1950);
or U2023 (N_2023,N_1946,N_1935);
and U2024 (N_2024,N_1929,N_1973);
nor U2025 (N_2025,N_1943,N_1947);
nor U2026 (N_2026,N_1973,N_1922);
or U2027 (N_2027,N_1942,N_1969);
and U2028 (N_2028,N_1951,N_1944);
nand U2029 (N_2029,N_1969,N_1946);
and U2030 (N_2030,N_1927,N_1967);
nor U2031 (N_2031,N_1926,N_1923);
nor U2032 (N_2032,N_1965,N_1957);
or U2033 (N_2033,N_1947,N_1951);
nand U2034 (N_2034,N_1972,N_1946);
nand U2035 (N_2035,N_1935,N_1955);
nor U2036 (N_2036,N_1964,N_1959);
nand U2037 (N_2037,N_1943,N_1960);
or U2038 (N_2038,N_1978,N_1925);
nand U2039 (N_2039,N_1938,N_1922);
nor U2040 (N_2040,N_2015,N_1999);
nor U2041 (N_2041,N_1998,N_1990);
nor U2042 (N_2042,N_2007,N_2038);
or U2043 (N_2043,N_1983,N_2000);
and U2044 (N_2044,N_2035,N_2011);
or U2045 (N_2045,N_2031,N_1988);
nor U2046 (N_2046,N_1992,N_2023);
nand U2047 (N_2047,N_2018,N_2032);
and U2048 (N_2048,N_2012,N_2022);
or U2049 (N_2049,N_1987,N_1991);
xnor U2050 (N_2050,N_2008,N_1994);
nand U2051 (N_2051,N_2034,N_1981);
nand U2052 (N_2052,N_2014,N_2001);
or U2053 (N_2053,N_2021,N_1984);
nor U2054 (N_2054,N_2027,N_1980);
and U2055 (N_2055,N_2025,N_1989);
nand U2056 (N_2056,N_1997,N_1996);
or U2057 (N_2057,N_2006,N_1995);
or U2058 (N_2058,N_2004,N_2002);
nand U2059 (N_2059,N_1986,N_1993);
or U2060 (N_2060,N_2010,N_2030);
or U2061 (N_2061,N_2036,N_2024);
nor U2062 (N_2062,N_2037,N_2017);
and U2063 (N_2063,N_2033,N_2028);
or U2064 (N_2064,N_2016,N_2003);
nand U2065 (N_2065,N_2009,N_2020);
nor U2066 (N_2066,N_2019,N_2026);
nand U2067 (N_2067,N_1985,N_2039);
nor U2068 (N_2068,N_2005,N_2029);
nor U2069 (N_2069,N_2013,N_1982);
xor U2070 (N_2070,N_2032,N_2033);
nor U2071 (N_2071,N_2000,N_2002);
nor U2072 (N_2072,N_2020,N_2035);
nand U2073 (N_2073,N_2029,N_2026);
or U2074 (N_2074,N_2016,N_2010);
and U2075 (N_2075,N_2017,N_2034);
nand U2076 (N_2076,N_2039,N_2027);
and U2077 (N_2077,N_2016,N_2009);
or U2078 (N_2078,N_1991,N_1983);
and U2079 (N_2079,N_2008,N_2038);
nand U2080 (N_2080,N_2016,N_2026);
nor U2081 (N_2081,N_2006,N_2023);
nor U2082 (N_2082,N_1990,N_2013);
nor U2083 (N_2083,N_1986,N_1999);
nor U2084 (N_2084,N_2000,N_2021);
xnor U2085 (N_2085,N_2022,N_2004);
nand U2086 (N_2086,N_1985,N_1986);
nor U2087 (N_2087,N_2014,N_2000);
xor U2088 (N_2088,N_2027,N_1994);
or U2089 (N_2089,N_2002,N_2021);
nor U2090 (N_2090,N_2031,N_2002);
xor U2091 (N_2091,N_1989,N_2027);
and U2092 (N_2092,N_2036,N_2025);
nor U2093 (N_2093,N_2037,N_2022);
or U2094 (N_2094,N_1980,N_1990);
nor U2095 (N_2095,N_2033,N_1980);
nor U2096 (N_2096,N_1992,N_2020);
or U2097 (N_2097,N_1999,N_1984);
nor U2098 (N_2098,N_2009,N_1985);
and U2099 (N_2099,N_2028,N_2039);
nor U2100 (N_2100,N_2077,N_2087);
nand U2101 (N_2101,N_2070,N_2093);
nor U2102 (N_2102,N_2076,N_2080);
or U2103 (N_2103,N_2074,N_2046);
nand U2104 (N_2104,N_2053,N_2083);
nand U2105 (N_2105,N_2085,N_2065);
nand U2106 (N_2106,N_2049,N_2061);
nand U2107 (N_2107,N_2059,N_2055);
nor U2108 (N_2108,N_2060,N_2096);
nand U2109 (N_2109,N_2079,N_2047);
nand U2110 (N_2110,N_2082,N_2078);
or U2111 (N_2111,N_2041,N_2098);
and U2112 (N_2112,N_2051,N_2094);
nand U2113 (N_2113,N_2073,N_2040);
or U2114 (N_2114,N_2091,N_2063);
nor U2115 (N_2115,N_2057,N_2050);
or U2116 (N_2116,N_2092,N_2068);
or U2117 (N_2117,N_2043,N_2052);
nor U2118 (N_2118,N_2056,N_2081);
and U2119 (N_2119,N_2045,N_2090);
or U2120 (N_2120,N_2097,N_2071);
and U2121 (N_2121,N_2044,N_2075);
nand U2122 (N_2122,N_2067,N_2084);
nand U2123 (N_2123,N_2048,N_2062);
or U2124 (N_2124,N_2088,N_2069);
or U2125 (N_2125,N_2042,N_2086);
nand U2126 (N_2126,N_2099,N_2095);
nand U2127 (N_2127,N_2072,N_2089);
nor U2128 (N_2128,N_2064,N_2054);
and U2129 (N_2129,N_2066,N_2058);
nand U2130 (N_2130,N_2095,N_2094);
nand U2131 (N_2131,N_2095,N_2069);
or U2132 (N_2132,N_2090,N_2043);
nand U2133 (N_2133,N_2044,N_2099);
or U2134 (N_2134,N_2087,N_2049);
nand U2135 (N_2135,N_2080,N_2096);
nand U2136 (N_2136,N_2093,N_2055);
or U2137 (N_2137,N_2063,N_2086);
nand U2138 (N_2138,N_2072,N_2040);
nand U2139 (N_2139,N_2069,N_2043);
nand U2140 (N_2140,N_2057,N_2080);
or U2141 (N_2141,N_2043,N_2055);
and U2142 (N_2142,N_2071,N_2086);
or U2143 (N_2143,N_2062,N_2061);
and U2144 (N_2144,N_2094,N_2050);
or U2145 (N_2145,N_2080,N_2098);
or U2146 (N_2146,N_2080,N_2079);
or U2147 (N_2147,N_2045,N_2060);
or U2148 (N_2148,N_2092,N_2089);
or U2149 (N_2149,N_2087,N_2047);
nand U2150 (N_2150,N_2063,N_2057);
and U2151 (N_2151,N_2067,N_2063);
nor U2152 (N_2152,N_2051,N_2089);
nand U2153 (N_2153,N_2061,N_2072);
or U2154 (N_2154,N_2065,N_2045);
nor U2155 (N_2155,N_2083,N_2049);
and U2156 (N_2156,N_2092,N_2074);
and U2157 (N_2157,N_2084,N_2076);
or U2158 (N_2158,N_2060,N_2069);
or U2159 (N_2159,N_2083,N_2047);
and U2160 (N_2160,N_2124,N_2125);
nor U2161 (N_2161,N_2108,N_2121);
and U2162 (N_2162,N_2128,N_2137);
or U2163 (N_2163,N_2157,N_2141);
or U2164 (N_2164,N_2113,N_2120);
nor U2165 (N_2165,N_2119,N_2104);
or U2166 (N_2166,N_2144,N_2159);
or U2167 (N_2167,N_2148,N_2103);
nand U2168 (N_2168,N_2118,N_2134);
and U2169 (N_2169,N_2111,N_2100);
and U2170 (N_2170,N_2139,N_2147);
or U2171 (N_2171,N_2117,N_2133);
or U2172 (N_2172,N_2131,N_2126);
nor U2173 (N_2173,N_2149,N_2101);
nand U2174 (N_2174,N_2142,N_2153);
nor U2175 (N_2175,N_2138,N_2106);
nand U2176 (N_2176,N_2132,N_2158);
or U2177 (N_2177,N_2154,N_2146);
and U2178 (N_2178,N_2122,N_2112);
or U2179 (N_2179,N_2116,N_2102);
or U2180 (N_2180,N_2155,N_2135);
and U2181 (N_2181,N_2105,N_2130);
xor U2182 (N_2182,N_2127,N_2150);
and U2183 (N_2183,N_2110,N_2143);
or U2184 (N_2184,N_2123,N_2145);
nor U2185 (N_2185,N_2156,N_2152);
nand U2186 (N_2186,N_2136,N_2115);
nand U2187 (N_2187,N_2129,N_2107);
nor U2188 (N_2188,N_2114,N_2140);
or U2189 (N_2189,N_2109,N_2151);
nor U2190 (N_2190,N_2137,N_2126);
and U2191 (N_2191,N_2114,N_2137);
nand U2192 (N_2192,N_2159,N_2146);
nand U2193 (N_2193,N_2101,N_2113);
or U2194 (N_2194,N_2154,N_2102);
nor U2195 (N_2195,N_2129,N_2154);
nand U2196 (N_2196,N_2127,N_2133);
or U2197 (N_2197,N_2139,N_2157);
or U2198 (N_2198,N_2129,N_2138);
or U2199 (N_2199,N_2138,N_2120);
or U2200 (N_2200,N_2140,N_2137);
nor U2201 (N_2201,N_2146,N_2143);
nand U2202 (N_2202,N_2105,N_2116);
nor U2203 (N_2203,N_2157,N_2116);
or U2204 (N_2204,N_2155,N_2130);
nand U2205 (N_2205,N_2116,N_2138);
or U2206 (N_2206,N_2158,N_2125);
nor U2207 (N_2207,N_2146,N_2104);
nor U2208 (N_2208,N_2103,N_2102);
nor U2209 (N_2209,N_2136,N_2106);
nand U2210 (N_2210,N_2138,N_2153);
nor U2211 (N_2211,N_2125,N_2111);
and U2212 (N_2212,N_2146,N_2155);
and U2213 (N_2213,N_2105,N_2109);
nand U2214 (N_2214,N_2141,N_2151);
nand U2215 (N_2215,N_2113,N_2111);
and U2216 (N_2216,N_2119,N_2103);
and U2217 (N_2217,N_2127,N_2144);
or U2218 (N_2218,N_2127,N_2148);
or U2219 (N_2219,N_2109,N_2115);
or U2220 (N_2220,N_2187,N_2160);
or U2221 (N_2221,N_2202,N_2176);
or U2222 (N_2222,N_2181,N_2196);
and U2223 (N_2223,N_2201,N_2192);
nor U2224 (N_2224,N_2170,N_2195);
and U2225 (N_2225,N_2219,N_2169);
or U2226 (N_2226,N_2164,N_2165);
and U2227 (N_2227,N_2167,N_2216);
or U2228 (N_2228,N_2206,N_2174);
or U2229 (N_2229,N_2199,N_2194);
nor U2230 (N_2230,N_2197,N_2209);
or U2231 (N_2231,N_2175,N_2204);
or U2232 (N_2232,N_2177,N_2212);
or U2233 (N_2233,N_2186,N_2198);
nand U2234 (N_2234,N_2217,N_2207);
nor U2235 (N_2235,N_2168,N_2203);
nand U2236 (N_2236,N_2171,N_2162);
or U2237 (N_2237,N_2210,N_2211);
nand U2238 (N_2238,N_2214,N_2193);
nor U2239 (N_2239,N_2179,N_2205);
nand U2240 (N_2240,N_2184,N_2218);
nor U2241 (N_2241,N_2173,N_2213);
nand U2242 (N_2242,N_2161,N_2180);
nand U2243 (N_2243,N_2178,N_2183);
and U2244 (N_2244,N_2189,N_2191);
nor U2245 (N_2245,N_2190,N_2182);
and U2246 (N_2246,N_2188,N_2163);
and U2247 (N_2247,N_2215,N_2166);
xnor U2248 (N_2248,N_2208,N_2200);
or U2249 (N_2249,N_2185,N_2172);
nand U2250 (N_2250,N_2161,N_2169);
and U2251 (N_2251,N_2205,N_2216);
nand U2252 (N_2252,N_2179,N_2161);
or U2253 (N_2253,N_2193,N_2187);
or U2254 (N_2254,N_2192,N_2203);
nand U2255 (N_2255,N_2217,N_2202);
and U2256 (N_2256,N_2218,N_2209);
nand U2257 (N_2257,N_2218,N_2203);
and U2258 (N_2258,N_2165,N_2187);
nor U2259 (N_2259,N_2203,N_2167);
nor U2260 (N_2260,N_2207,N_2162);
and U2261 (N_2261,N_2212,N_2198);
and U2262 (N_2262,N_2168,N_2205);
nor U2263 (N_2263,N_2214,N_2204);
nand U2264 (N_2264,N_2172,N_2173);
or U2265 (N_2265,N_2173,N_2219);
or U2266 (N_2266,N_2218,N_2178);
nor U2267 (N_2267,N_2169,N_2203);
and U2268 (N_2268,N_2171,N_2195);
or U2269 (N_2269,N_2182,N_2198);
nand U2270 (N_2270,N_2175,N_2208);
nand U2271 (N_2271,N_2178,N_2161);
nor U2272 (N_2272,N_2169,N_2162);
nand U2273 (N_2273,N_2167,N_2180);
or U2274 (N_2274,N_2206,N_2179);
nor U2275 (N_2275,N_2171,N_2189);
nor U2276 (N_2276,N_2169,N_2175);
nand U2277 (N_2277,N_2165,N_2173);
or U2278 (N_2278,N_2162,N_2198);
nand U2279 (N_2279,N_2180,N_2196);
or U2280 (N_2280,N_2248,N_2253);
and U2281 (N_2281,N_2244,N_2260);
nor U2282 (N_2282,N_2268,N_2277);
nand U2283 (N_2283,N_2257,N_2236);
nor U2284 (N_2284,N_2251,N_2274);
nor U2285 (N_2285,N_2229,N_2232);
or U2286 (N_2286,N_2238,N_2259);
nor U2287 (N_2287,N_2275,N_2269);
or U2288 (N_2288,N_2231,N_2225);
and U2289 (N_2289,N_2247,N_2245);
nand U2290 (N_2290,N_2235,N_2272);
and U2291 (N_2291,N_2240,N_2249);
and U2292 (N_2292,N_2254,N_2220);
and U2293 (N_2293,N_2228,N_2241);
and U2294 (N_2294,N_2246,N_2271);
nand U2295 (N_2295,N_2243,N_2258);
or U2296 (N_2296,N_2223,N_2239);
and U2297 (N_2297,N_2252,N_2278);
or U2298 (N_2298,N_2256,N_2276);
nand U2299 (N_2299,N_2237,N_2273);
nand U2300 (N_2300,N_2267,N_2266);
nor U2301 (N_2301,N_2222,N_2242);
and U2302 (N_2302,N_2234,N_2261);
and U2303 (N_2303,N_2226,N_2230);
and U2304 (N_2304,N_2279,N_2265);
nand U2305 (N_2305,N_2255,N_2270);
nand U2306 (N_2306,N_2233,N_2262);
nand U2307 (N_2307,N_2264,N_2224);
nor U2308 (N_2308,N_2263,N_2250);
nand U2309 (N_2309,N_2221,N_2227);
nand U2310 (N_2310,N_2278,N_2273);
or U2311 (N_2311,N_2240,N_2224);
nand U2312 (N_2312,N_2257,N_2241);
nor U2313 (N_2313,N_2233,N_2250);
nor U2314 (N_2314,N_2270,N_2279);
or U2315 (N_2315,N_2231,N_2250);
or U2316 (N_2316,N_2276,N_2253);
or U2317 (N_2317,N_2279,N_2246);
and U2318 (N_2318,N_2277,N_2243);
or U2319 (N_2319,N_2253,N_2240);
and U2320 (N_2320,N_2266,N_2261);
nand U2321 (N_2321,N_2273,N_2264);
nor U2322 (N_2322,N_2225,N_2258);
or U2323 (N_2323,N_2251,N_2227);
nor U2324 (N_2324,N_2272,N_2276);
and U2325 (N_2325,N_2268,N_2274);
and U2326 (N_2326,N_2225,N_2254);
nor U2327 (N_2327,N_2237,N_2229);
and U2328 (N_2328,N_2274,N_2270);
and U2329 (N_2329,N_2247,N_2232);
or U2330 (N_2330,N_2269,N_2243);
nand U2331 (N_2331,N_2265,N_2254);
or U2332 (N_2332,N_2239,N_2241);
nand U2333 (N_2333,N_2254,N_2249);
or U2334 (N_2334,N_2227,N_2246);
nand U2335 (N_2335,N_2222,N_2265);
nand U2336 (N_2336,N_2279,N_2241);
nand U2337 (N_2337,N_2227,N_2266);
or U2338 (N_2338,N_2242,N_2264);
nor U2339 (N_2339,N_2259,N_2274);
or U2340 (N_2340,N_2282,N_2326);
nand U2341 (N_2341,N_2285,N_2298);
and U2342 (N_2342,N_2315,N_2317);
nor U2343 (N_2343,N_2283,N_2311);
or U2344 (N_2344,N_2328,N_2325);
nor U2345 (N_2345,N_2289,N_2290);
nor U2346 (N_2346,N_2304,N_2318);
or U2347 (N_2347,N_2324,N_2314);
or U2348 (N_2348,N_2312,N_2296);
nor U2349 (N_2349,N_2302,N_2332);
nor U2350 (N_2350,N_2339,N_2280);
and U2351 (N_2351,N_2281,N_2330);
nand U2352 (N_2352,N_2333,N_2291);
nand U2353 (N_2353,N_2295,N_2319);
nor U2354 (N_2354,N_2288,N_2308);
nor U2355 (N_2355,N_2297,N_2322);
or U2356 (N_2356,N_2286,N_2309);
and U2357 (N_2357,N_2292,N_2284);
nor U2358 (N_2358,N_2307,N_2293);
and U2359 (N_2359,N_2320,N_2316);
or U2360 (N_2360,N_2338,N_2306);
nand U2361 (N_2361,N_2321,N_2335);
and U2362 (N_2362,N_2327,N_2334);
or U2363 (N_2363,N_2313,N_2310);
nand U2364 (N_2364,N_2331,N_2299);
nor U2365 (N_2365,N_2303,N_2287);
nand U2366 (N_2366,N_2300,N_2337);
or U2367 (N_2367,N_2336,N_2329);
nand U2368 (N_2368,N_2294,N_2301);
nor U2369 (N_2369,N_2305,N_2323);
or U2370 (N_2370,N_2287,N_2283);
or U2371 (N_2371,N_2308,N_2323);
nand U2372 (N_2372,N_2282,N_2309);
or U2373 (N_2373,N_2320,N_2336);
nor U2374 (N_2374,N_2334,N_2328);
and U2375 (N_2375,N_2282,N_2285);
nand U2376 (N_2376,N_2298,N_2308);
nor U2377 (N_2377,N_2330,N_2328);
and U2378 (N_2378,N_2287,N_2304);
or U2379 (N_2379,N_2296,N_2326);
and U2380 (N_2380,N_2323,N_2285);
or U2381 (N_2381,N_2286,N_2291);
nand U2382 (N_2382,N_2302,N_2310);
nand U2383 (N_2383,N_2282,N_2311);
and U2384 (N_2384,N_2309,N_2316);
nand U2385 (N_2385,N_2297,N_2325);
nor U2386 (N_2386,N_2292,N_2334);
nand U2387 (N_2387,N_2303,N_2317);
nor U2388 (N_2388,N_2314,N_2310);
nand U2389 (N_2389,N_2337,N_2328);
or U2390 (N_2390,N_2313,N_2332);
and U2391 (N_2391,N_2333,N_2286);
and U2392 (N_2392,N_2284,N_2295);
and U2393 (N_2393,N_2286,N_2332);
nor U2394 (N_2394,N_2318,N_2322);
nor U2395 (N_2395,N_2331,N_2313);
and U2396 (N_2396,N_2287,N_2307);
or U2397 (N_2397,N_2303,N_2327);
nand U2398 (N_2398,N_2284,N_2285);
nor U2399 (N_2399,N_2321,N_2333);
and U2400 (N_2400,N_2359,N_2357);
or U2401 (N_2401,N_2372,N_2389);
or U2402 (N_2402,N_2392,N_2347);
nor U2403 (N_2403,N_2340,N_2366);
nor U2404 (N_2404,N_2374,N_2386);
nor U2405 (N_2405,N_2384,N_2367);
nand U2406 (N_2406,N_2387,N_2399);
nand U2407 (N_2407,N_2379,N_2360);
or U2408 (N_2408,N_2348,N_2377);
or U2409 (N_2409,N_2371,N_2380);
or U2410 (N_2410,N_2365,N_2373);
or U2411 (N_2411,N_2368,N_2358);
nand U2412 (N_2412,N_2382,N_2351);
nor U2413 (N_2413,N_2355,N_2341);
or U2414 (N_2414,N_2390,N_2345);
nor U2415 (N_2415,N_2349,N_2363);
nand U2416 (N_2416,N_2378,N_2362);
or U2417 (N_2417,N_2397,N_2342);
nor U2418 (N_2418,N_2388,N_2394);
or U2419 (N_2419,N_2370,N_2344);
and U2420 (N_2420,N_2395,N_2383);
or U2421 (N_2421,N_2354,N_2396);
or U2422 (N_2422,N_2346,N_2356);
nand U2423 (N_2423,N_2343,N_2391);
or U2424 (N_2424,N_2353,N_2361);
and U2425 (N_2425,N_2393,N_2385);
and U2426 (N_2426,N_2352,N_2350);
nor U2427 (N_2427,N_2375,N_2376);
nor U2428 (N_2428,N_2369,N_2364);
nand U2429 (N_2429,N_2398,N_2381);
or U2430 (N_2430,N_2386,N_2359);
nor U2431 (N_2431,N_2351,N_2353);
nor U2432 (N_2432,N_2392,N_2378);
nor U2433 (N_2433,N_2395,N_2355);
nand U2434 (N_2434,N_2379,N_2384);
or U2435 (N_2435,N_2387,N_2351);
or U2436 (N_2436,N_2368,N_2391);
nor U2437 (N_2437,N_2395,N_2394);
or U2438 (N_2438,N_2346,N_2354);
or U2439 (N_2439,N_2352,N_2354);
and U2440 (N_2440,N_2367,N_2369);
nor U2441 (N_2441,N_2363,N_2380);
and U2442 (N_2442,N_2390,N_2369);
xor U2443 (N_2443,N_2376,N_2347);
and U2444 (N_2444,N_2359,N_2362);
nor U2445 (N_2445,N_2381,N_2393);
nand U2446 (N_2446,N_2393,N_2377);
nor U2447 (N_2447,N_2399,N_2369);
nand U2448 (N_2448,N_2360,N_2393);
nor U2449 (N_2449,N_2377,N_2342);
and U2450 (N_2450,N_2347,N_2373);
and U2451 (N_2451,N_2344,N_2380);
nor U2452 (N_2452,N_2392,N_2353);
and U2453 (N_2453,N_2386,N_2376);
and U2454 (N_2454,N_2392,N_2376);
and U2455 (N_2455,N_2394,N_2376);
or U2456 (N_2456,N_2352,N_2398);
or U2457 (N_2457,N_2362,N_2392);
and U2458 (N_2458,N_2398,N_2341);
and U2459 (N_2459,N_2345,N_2397);
and U2460 (N_2460,N_2443,N_2459);
and U2461 (N_2461,N_2449,N_2407);
and U2462 (N_2462,N_2408,N_2435);
or U2463 (N_2463,N_2418,N_2409);
or U2464 (N_2464,N_2414,N_2440);
or U2465 (N_2465,N_2400,N_2411);
nor U2466 (N_2466,N_2441,N_2434);
or U2467 (N_2467,N_2447,N_2427);
or U2468 (N_2468,N_2439,N_2403);
nand U2469 (N_2469,N_2426,N_2448);
or U2470 (N_2470,N_2456,N_2429);
or U2471 (N_2471,N_2420,N_2451);
and U2472 (N_2472,N_2452,N_2454);
and U2473 (N_2473,N_2431,N_2453);
nor U2474 (N_2474,N_2446,N_2438);
nor U2475 (N_2475,N_2424,N_2455);
nor U2476 (N_2476,N_2442,N_2444);
or U2477 (N_2477,N_2402,N_2401);
and U2478 (N_2478,N_2458,N_2415);
nor U2479 (N_2479,N_2432,N_2436);
nor U2480 (N_2480,N_2425,N_2419);
nand U2481 (N_2481,N_2457,N_2416);
nand U2482 (N_2482,N_2417,N_2428);
or U2483 (N_2483,N_2433,N_2421);
xor U2484 (N_2484,N_2450,N_2406);
nor U2485 (N_2485,N_2410,N_2422);
nand U2486 (N_2486,N_2430,N_2412);
nor U2487 (N_2487,N_2423,N_2413);
or U2488 (N_2488,N_2405,N_2437);
nor U2489 (N_2489,N_2404,N_2445);
nand U2490 (N_2490,N_2439,N_2422);
or U2491 (N_2491,N_2402,N_2451);
nand U2492 (N_2492,N_2428,N_2424);
nand U2493 (N_2493,N_2408,N_2419);
and U2494 (N_2494,N_2403,N_2401);
nor U2495 (N_2495,N_2407,N_2411);
nand U2496 (N_2496,N_2414,N_2424);
nor U2497 (N_2497,N_2454,N_2411);
nor U2498 (N_2498,N_2447,N_2458);
or U2499 (N_2499,N_2450,N_2413);
nand U2500 (N_2500,N_2453,N_2413);
nand U2501 (N_2501,N_2438,N_2424);
or U2502 (N_2502,N_2426,N_2434);
nand U2503 (N_2503,N_2450,N_2424);
nor U2504 (N_2504,N_2432,N_2430);
and U2505 (N_2505,N_2411,N_2445);
nor U2506 (N_2506,N_2428,N_2402);
and U2507 (N_2507,N_2402,N_2424);
and U2508 (N_2508,N_2429,N_2408);
nand U2509 (N_2509,N_2440,N_2429);
nor U2510 (N_2510,N_2434,N_2456);
nor U2511 (N_2511,N_2456,N_2401);
nand U2512 (N_2512,N_2456,N_2436);
or U2513 (N_2513,N_2412,N_2431);
or U2514 (N_2514,N_2417,N_2416);
or U2515 (N_2515,N_2415,N_2404);
nand U2516 (N_2516,N_2418,N_2425);
or U2517 (N_2517,N_2456,N_2428);
and U2518 (N_2518,N_2404,N_2411);
nor U2519 (N_2519,N_2415,N_2450);
and U2520 (N_2520,N_2483,N_2467);
nand U2521 (N_2521,N_2499,N_2515);
nand U2522 (N_2522,N_2490,N_2481);
nand U2523 (N_2523,N_2465,N_2461);
and U2524 (N_2524,N_2488,N_2510);
nor U2525 (N_2525,N_2497,N_2472);
or U2526 (N_2526,N_2469,N_2463);
and U2527 (N_2527,N_2505,N_2517);
and U2528 (N_2528,N_2477,N_2476);
nor U2529 (N_2529,N_2501,N_2485);
and U2530 (N_2530,N_2466,N_2516);
nor U2531 (N_2531,N_2484,N_2519);
and U2532 (N_2532,N_2513,N_2495);
or U2533 (N_2533,N_2474,N_2482);
nor U2534 (N_2534,N_2473,N_2468);
and U2535 (N_2535,N_2475,N_2491);
and U2536 (N_2536,N_2496,N_2500);
nand U2537 (N_2537,N_2460,N_2506);
nand U2538 (N_2538,N_2486,N_2511);
nand U2539 (N_2539,N_2493,N_2479);
or U2540 (N_2540,N_2508,N_2514);
or U2541 (N_2541,N_2462,N_2504);
nor U2542 (N_2542,N_2518,N_2480);
and U2543 (N_2543,N_2487,N_2470);
or U2544 (N_2544,N_2471,N_2478);
and U2545 (N_2545,N_2502,N_2492);
or U2546 (N_2546,N_2494,N_2464);
and U2547 (N_2547,N_2507,N_2509);
and U2548 (N_2548,N_2503,N_2489);
nand U2549 (N_2549,N_2512,N_2498);
nand U2550 (N_2550,N_2493,N_2465);
or U2551 (N_2551,N_2480,N_2465);
and U2552 (N_2552,N_2468,N_2467);
nor U2553 (N_2553,N_2472,N_2513);
nand U2554 (N_2554,N_2486,N_2502);
and U2555 (N_2555,N_2516,N_2473);
and U2556 (N_2556,N_2477,N_2467);
nor U2557 (N_2557,N_2473,N_2502);
nand U2558 (N_2558,N_2461,N_2515);
or U2559 (N_2559,N_2509,N_2508);
nor U2560 (N_2560,N_2500,N_2476);
nor U2561 (N_2561,N_2514,N_2477);
or U2562 (N_2562,N_2466,N_2506);
nand U2563 (N_2563,N_2495,N_2512);
nor U2564 (N_2564,N_2460,N_2509);
nand U2565 (N_2565,N_2512,N_2486);
or U2566 (N_2566,N_2474,N_2464);
nor U2567 (N_2567,N_2488,N_2498);
and U2568 (N_2568,N_2460,N_2461);
nand U2569 (N_2569,N_2484,N_2513);
and U2570 (N_2570,N_2491,N_2460);
or U2571 (N_2571,N_2468,N_2502);
or U2572 (N_2572,N_2519,N_2501);
and U2573 (N_2573,N_2473,N_2519);
and U2574 (N_2574,N_2502,N_2496);
nand U2575 (N_2575,N_2470,N_2481);
nand U2576 (N_2576,N_2489,N_2483);
nand U2577 (N_2577,N_2469,N_2513);
or U2578 (N_2578,N_2468,N_2505);
or U2579 (N_2579,N_2518,N_2470);
nand U2580 (N_2580,N_2529,N_2539);
and U2581 (N_2581,N_2534,N_2568);
or U2582 (N_2582,N_2560,N_2555);
nand U2583 (N_2583,N_2558,N_2547);
nor U2584 (N_2584,N_2565,N_2542);
nor U2585 (N_2585,N_2557,N_2549);
or U2586 (N_2586,N_2527,N_2562);
or U2587 (N_2587,N_2531,N_2575);
and U2588 (N_2588,N_2573,N_2541);
nor U2589 (N_2589,N_2528,N_2540);
nand U2590 (N_2590,N_2543,N_2566);
and U2591 (N_2591,N_2523,N_2570);
or U2592 (N_2592,N_2574,N_2567);
nor U2593 (N_2593,N_2576,N_2545);
nor U2594 (N_2594,N_2561,N_2525);
and U2595 (N_2595,N_2544,N_2520);
nand U2596 (N_2596,N_2522,N_2521);
or U2597 (N_2597,N_2537,N_2556);
nand U2598 (N_2598,N_2538,N_2548);
nand U2599 (N_2599,N_2551,N_2546);
nand U2600 (N_2600,N_2533,N_2563);
xnor U2601 (N_2601,N_2552,N_2530);
nor U2602 (N_2602,N_2526,N_2559);
nand U2603 (N_2603,N_2532,N_2578);
or U2604 (N_2604,N_2571,N_2553);
nor U2605 (N_2605,N_2579,N_2554);
or U2606 (N_2606,N_2572,N_2536);
nor U2607 (N_2607,N_2524,N_2550);
nor U2608 (N_2608,N_2564,N_2577);
nor U2609 (N_2609,N_2535,N_2569);
nand U2610 (N_2610,N_2539,N_2562);
and U2611 (N_2611,N_2543,N_2562);
or U2612 (N_2612,N_2527,N_2526);
nand U2613 (N_2613,N_2559,N_2548);
nand U2614 (N_2614,N_2570,N_2569);
nand U2615 (N_2615,N_2521,N_2533);
nor U2616 (N_2616,N_2530,N_2549);
and U2617 (N_2617,N_2567,N_2566);
and U2618 (N_2618,N_2526,N_2563);
and U2619 (N_2619,N_2524,N_2571);
or U2620 (N_2620,N_2543,N_2529);
and U2621 (N_2621,N_2575,N_2533);
nand U2622 (N_2622,N_2531,N_2521);
nand U2623 (N_2623,N_2570,N_2560);
and U2624 (N_2624,N_2571,N_2532);
nand U2625 (N_2625,N_2568,N_2558);
nor U2626 (N_2626,N_2561,N_2547);
xnor U2627 (N_2627,N_2561,N_2551);
or U2628 (N_2628,N_2563,N_2551);
or U2629 (N_2629,N_2538,N_2521);
and U2630 (N_2630,N_2560,N_2535);
or U2631 (N_2631,N_2536,N_2533);
or U2632 (N_2632,N_2565,N_2558);
nor U2633 (N_2633,N_2575,N_2526);
nand U2634 (N_2634,N_2531,N_2522);
nand U2635 (N_2635,N_2538,N_2523);
and U2636 (N_2636,N_2556,N_2523);
nand U2637 (N_2637,N_2539,N_2549);
and U2638 (N_2638,N_2542,N_2532);
nand U2639 (N_2639,N_2527,N_2524);
nand U2640 (N_2640,N_2632,N_2624);
nor U2641 (N_2641,N_2593,N_2588);
and U2642 (N_2642,N_2636,N_2612);
nor U2643 (N_2643,N_2596,N_2587);
nor U2644 (N_2644,N_2625,N_2620);
nor U2645 (N_2645,N_2582,N_2630);
and U2646 (N_2646,N_2606,N_2591);
nand U2647 (N_2647,N_2594,N_2599);
nor U2648 (N_2648,N_2585,N_2617);
or U2649 (N_2649,N_2631,N_2609);
nand U2650 (N_2650,N_2613,N_2602);
and U2651 (N_2651,N_2615,N_2597);
or U2652 (N_2652,N_2627,N_2622);
nand U2653 (N_2653,N_2600,N_2618);
nand U2654 (N_2654,N_2603,N_2628);
nand U2655 (N_2655,N_2583,N_2607);
or U2656 (N_2656,N_2635,N_2580);
and U2657 (N_2657,N_2581,N_2616);
nand U2658 (N_2658,N_2598,N_2605);
and U2659 (N_2659,N_2610,N_2611);
or U2660 (N_2660,N_2608,N_2604);
and U2661 (N_2661,N_2629,N_2638);
nor U2662 (N_2662,N_2623,N_2633);
nor U2663 (N_2663,N_2637,N_2584);
or U2664 (N_2664,N_2586,N_2619);
nand U2665 (N_2665,N_2634,N_2589);
nand U2666 (N_2666,N_2626,N_2614);
and U2667 (N_2667,N_2601,N_2621);
nor U2668 (N_2668,N_2590,N_2595);
nand U2669 (N_2669,N_2639,N_2592);
xnor U2670 (N_2670,N_2621,N_2627);
nor U2671 (N_2671,N_2609,N_2627);
nand U2672 (N_2672,N_2634,N_2582);
or U2673 (N_2673,N_2591,N_2585);
nor U2674 (N_2674,N_2586,N_2608);
and U2675 (N_2675,N_2582,N_2598);
nor U2676 (N_2676,N_2626,N_2616);
and U2677 (N_2677,N_2611,N_2628);
nand U2678 (N_2678,N_2637,N_2620);
nor U2679 (N_2679,N_2627,N_2583);
nor U2680 (N_2680,N_2637,N_2639);
and U2681 (N_2681,N_2587,N_2602);
and U2682 (N_2682,N_2624,N_2595);
nor U2683 (N_2683,N_2586,N_2611);
nand U2684 (N_2684,N_2612,N_2614);
or U2685 (N_2685,N_2629,N_2592);
nand U2686 (N_2686,N_2582,N_2632);
nand U2687 (N_2687,N_2632,N_2618);
nor U2688 (N_2688,N_2586,N_2635);
and U2689 (N_2689,N_2614,N_2615);
nand U2690 (N_2690,N_2635,N_2615);
or U2691 (N_2691,N_2636,N_2601);
nand U2692 (N_2692,N_2620,N_2584);
nand U2693 (N_2693,N_2627,N_2600);
or U2694 (N_2694,N_2639,N_2638);
or U2695 (N_2695,N_2633,N_2604);
nor U2696 (N_2696,N_2586,N_2624);
and U2697 (N_2697,N_2630,N_2608);
nor U2698 (N_2698,N_2599,N_2590);
nand U2699 (N_2699,N_2582,N_2586);
nand U2700 (N_2700,N_2663,N_2697);
or U2701 (N_2701,N_2673,N_2688);
nor U2702 (N_2702,N_2659,N_2670);
or U2703 (N_2703,N_2684,N_2648);
and U2704 (N_2704,N_2667,N_2696);
or U2705 (N_2705,N_2671,N_2650);
or U2706 (N_2706,N_2678,N_2644);
nor U2707 (N_2707,N_2645,N_2643);
xor U2708 (N_2708,N_2680,N_2656);
or U2709 (N_2709,N_2642,N_2641);
nor U2710 (N_2710,N_2664,N_2661);
and U2711 (N_2711,N_2654,N_2665);
nand U2712 (N_2712,N_2640,N_2690);
and U2713 (N_2713,N_2686,N_2653);
nor U2714 (N_2714,N_2655,N_2675);
and U2715 (N_2715,N_2651,N_2666);
nand U2716 (N_2716,N_2658,N_2672);
and U2717 (N_2717,N_2677,N_2681);
nor U2718 (N_2718,N_2699,N_2660);
xnor U2719 (N_2719,N_2689,N_2649);
nand U2720 (N_2720,N_2682,N_2652);
nand U2721 (N_2721,N_2693,N_2698);
and U2722 (N_2722,N_2683,N_2685);
xnor U2723 (N_2723,N_2674,N_2687);
and U2724 (N_2724,N_2692,N_2657);
or U2725 (N_2725,N_2668,N_2647);
nor U2726 (N_2726,N_2679,N_2662);
nand U2727 (N_2727,N_2695,N_2691);
nand U2728 (N_2728,N_2694,N_2669);
nor U2729 (N_2729,N_2646,N_2676);
xnor U2730 (N_2730,N_2656,N_2663);
nand U2731 (N_2731,N_2682,N_2692);
and U2732 (N_2732,N_2668,N_2684);
nor U2733 (N_2733,N_2657,N_2646);
nor U2734 (N_2734,N_2687,N_2698);
and U2735 (N_2735,N_2681,N_2649);
nand U2736 (N_2736,N_2686,N_2660);
or U2737 (N_2737,N_2664,N_2676);
and U2738 (N_2738,N_2642,N_2648);
nand U2739 (N_2739,N_2667,N_2646);
nand U2740 (N_2740,N_2697,N_2653);
nor U2741 (N_2741,N_2672,N_2650);
or U2742 (N_2742,N_2679,N_2674);
and U2743 (N_2743,N_2644,N_2673);
or U2744 (N_2744,N_2672,N_2682);
and U2745 (N_2745,N_2681,N_2670);
nor U2746 (N_2746,N_2690,N_2674);
nand U2747 (N_2747,N_2661,N_2693);
nor U2748 (N_2748,N_2659,N_2678);
nand U2749 (N_2749,N_2665,N_2656);
nand U2750 (N_2750,N_2669,N_2645);
and U2751 (N_2751,N_2689,N_2656);
nand U2752 (N_2752,N_2657,N_2650);
nand U2753 (N_2753,N_2647,N_2678);
nand U2754 (N_2754,N_2679,N_2683);
nor U2755 (N_2755,N_2642,N_2654);
and U2756 (N_2756,N_2691,N_2688);
and U2757 (N_2757,N_2660,N_2646);
nand U2758 (N_2758,N_2692,N_2673);
or U2759 (N_2759,N_2665,N_2698);
nor U2760 (N_2760,N_2728,N_2716);
and U2761 (N_2761,N_2704,N_2742);
nand U2762 (N_2762,N_2732,N_2755);
or U2763 (N_2763,N_2754,N_2756);
nor U2764 (N_2764,N_2736,N_2709);
and U2765 (N_2765,N_2737,N_2734);
or U2766 (N_2766,N_2725,N_2740);
nor U2767 (N_2767,N_2730,N_2744);
and U2768 (N_2768,N_2733,N_2719);
nor U2769 (N_2769,N_2702,N_2749);
and U2770 (N_2770,N_2714,N_2706);
or U2771 (N_2771,N_2757,N_2724);
and U2772 (N_2772,N_2721,N_2729);
or U2773 (N_2773,N_2711,N_2735);
nand U2774 (N_2774,N_2758,N_2750);
nand U2775 (N_2775,N_2741,N_2748);
nor U2776 (N_2776,N_2752,N_2739);
or U2777 (N_2777,N_2759,N_2705);
and U2778 (N_2778,N_2751,N_2708);
nor U2779 (N_2779,N_2727,N_2723);
and U2780 (N_2780,N_2701,N_2703);
and U2781 (N_2781,N_2720,N_2745);
nand U2782 (N_2782,N_2753,N_2712);
and U2783 (N_2783,N_2717,N_2722);
nor U2784 (N_2784,N_2715,N_2707);
nor U2785 (N_2785,N_2713,N_2731);
and U2786 (N_2786,N_2743,N_2700);
nand U2787 (N_2787,N_2746,N_2710);
and U2788 (N_2788,N_2747,N_2718);
nand U2789 (N_2789,N_2738,N_2726);
nand U2790 (N_2790,N_2735,N_2758);
nand U2791 (N_2791,N_2740,N_2739);
or U2792 (N_2792,N_2739,N_2711);
or U2793 (N_2793,N_2722,N_2753);
and U2794 (N_2794,N_2714,N_2725);
nand U2795 (N_2795,N_2733,N_2758);
nor U2796 (N_2796,N_2742,N_2746);
nand U2797 (N_2797,N_2701,N_2702);
nand U2798 (N_2798,N_2738,N_2712);
or U2799 (N_2799,N_2736,N_2742);
and U2800 (N_2800,N_2700,N_2705);
nor U2801 (N_2801,N_2721,N_2728);
nand U2802 (N_2802,N_2724,N_2720);
or U2803 (N_2803,N_2744,N_2706);
nand U2804 (N_2804,N_2731,N_2752);
nand U2805 (N_2805,N_2715,N_2719);
nor U2806 (N_2806,N_2705,N_2738);
nor U2807 (N_2807,N_2755,N_2749);
or U2808 (N_2808,N_2743,N_2756);
or U2809 (N_2809,N_2721,N_2730);
and U2810 (N_2810,N_2710,N_2703);
or U2811 (N_2811,N_2719,N_2745);
or U2812 (N_2812,N_2711,N_2747);
nand U2813 (N_2813,N_2730,N_2737);
nor U2814 (N_2814,N_2700,N_2713);
and U2815 (N_2815,N_2703,N_2732);
or U2816 (N_2816,N_2710,N_2730);
nand U2817 (N_2817,N_2735,N_2721);
nand U2818 (N_2818,N_2737,N_2750);
or U2819 (N_2819,N_2744,N_2741);
nand U2820 (N_2820,N_2794,N_2787);
and U2821 (N_2821,N_2799,N_2765);
and U2822 (N_2822,N_2813,N_2793);
or U2823 (N_2823,N_2776,N_2786);
or U2824 (N_2824,N_2807,N_2777);
and U2825 (N_2825,N_2805,N_2769);
or U2826 (N_2826,N_2780,N_2797);
xnor U2827 (N_2827,N_2803,N_2768);
and U2828 (N_2828,N_2811,N_2814);
nor U2829 (N_2829,N_2764,N_2818);
nor U2830 (N_2830,N_2788,N_2785);
and U2831 (N_2831,N_2783,N_2798);
or U2832 (N_2832,N_2779,N_2775);
xnor U2833 (N_2833,N_2763,N_2781);
and U2834 (N_2834,N_2760,N_2801);
nand U2835 (N_2835,N_2791,N_2778);
nor U2836 (N_2836,N_2762,N_2817);
or U2837 (N_2837,N_2810,N_2767);
or U2838 (N_2838,N_2790,N_2761);
nor U2839 (N_2839,N_2802,N_2772);
nand U2840 (N_2840,N_2796,N_2770);
and U2841 (N_2841,N_2809,N_2812);
or U2842 (N_2842,N_2808,N_2806);
and U2843 (N_2843,N_2774,N_2782);
or U2844 (N_2844,N_2771,N_2819);
or U2845 (N_2845,N_2816,N_2789);
nand U2846 (N_2846,N_2795,N_2792);
nand U2847 (N_2847,N_2815,N_2784);
nand U2848 (N_2848,N_2800,N_2766);
nand U2849 (N_2849,N_2804,N_2773);
and U2850 (N_2850,N_2808,N_2772);
or U2851 (N_2851,N_2787,N_2769);
and U2852 (N_2852,N_2811,N_2800);
and U2853 (N_2853,N_2816,N_2788);
nor U2854 (N_2854,N_2771,N_2780);
and U2855 (N_2855,N_2815,N_2777);
nand U2856 (N_2856,N_2781,N_2805);
and U2857 (N_2857,N_2790,N_2779);
nor U2858 (N_2858,N_2799,N_2784);
or U2859 (N_2859,N_2776,N_2777);
or U2860 (N_2860,N_2794,N_2769);
and U2861 (N_2861,N_2777,N_2779);
and U2862 (N_2862,N_2801,N_2765);
nand U2863 (N_2863,N_2773,N_2795);
and U2864 (N_2864,N_2817,N_2785);
nand U2865 (N_2865,N_2769,N_2795);
nor U2866 (N_2866,N_2799,N_2809);
or U2867 (N_2867,N_2764,N_2811);
nand U2868 (N_2868,N_2789,N_2762);
and U2869 (N_2869,N_2811,N_2819);
nor U2870 (N_2870,N_2776,N_2814);
and U2871 (N_2871,N_2802,N_2776);
and U2872 (N_2872,N_2810,N_2771);
and U2873 (N_2873,N_2760,N_2802);
and U2874 (N_2874,N_2776,N_2762);
nor U2875 (N_2875,N_2791,N_2816);
nand U2876 (N_2876,N_2807,N_2793);
nor U2877 (N_2877,N_2780,N_2773);
nor U2878 (N_2878,N_2768,N_2767);
and U2879 (N_2879,N_2765,N_2770);
nor U2880 (N_2880,N_2869,N_2877);
nor U2881 (N_2881,N_2852,N_2873);
and U2882 (N_2882,N_2851,N_2874);
nand U2883 (N_2883,N_2843,N_2865);
nand U2884 (N_2884,N_2879,N_2844);
or U2885 (N_2885,N_2825,N_2845);
nor U2886 (N_2886,N_2876,N_2868);
nand U2887 (N_2887,N_2826,N_2860);
and U2888 (N_2888,N_2863,N_2850);
nor U2889 (N_2889,N_2847,N_2853);
nor U2890 (N_2890,N_2828,N_2822);
nor U2891 (N_2891,N_2872,N_2862);
nor U2892 (N_2892,N_2854,N_2837);
and U2893 (N_2893,N_2841,N_2857);
or U2894 (N_2894,N_2823,N_2859);
and U2895 (N_2895,N_2824,N_2820);
or U2896 (N_2896,N_2835,N_2878);
nor U2897 (N_2897,N_2834,N_2829);
nor U2898 (N_2898,N_2866,N_2864);
and U2899 (N_2899,N_2832,N_2821);
and U2900 (N_2900,N_2870,N_2855);
nor U2901 (N_2901,N_2846,N_2861);
and U2902 (N_2902,N_2856,N_2842);
nor U2903 (N_2903,N_2858,N_2839);
or U2904 (N_2904,N_2875,N_2871);
or U2905 (N_2905,N_2827,N_2838);
xor U2906 (N_2906,N_2840,N_2867);
and U2907 (N_2907,N_2848,N_2833);
nand U2908 (N_2908,N_2849,N_2836);
and U2909 (N_2909,N_2831,N_2830);
nand U2910 (N_2910,N_2824,N_2845);
nor U2911 (N_2911,N_2875,N_2851);
nand U2912 (N_2912,N_2834,N_2859);
or U2913 (N_2913,N_2872,N_2853);
nor U2914 (N_2914,N_2830,N_2834);
and U2915 (N_2915,N_2820,N_2865);
or U2916 (N_2916,N_2843,N_2861);
xnor U2917 (N_2917,N_2869,N_2830);
nor U2918 (N_2918,N_2827,N_2835);
nand U2919 (N_2919,N_2857,N_2850);
nand U2920 (N_2920,N_2864,N_2828);
or U2921 (N_2921,N_2840,N_2875);
or U2922 (N_2922,N_2829,N_2869);
nor U2923 (N_2923,N_2873,N_2827);
nand U2924 (N_2924,N_2838,N_2851);
nor U2925 (N_2925,N_2877,N_2872);
nand U2926 (N_2926,N_2835,N_2871);
nand U2927 (N_2927,N_2854,N_2853);
xnor U2928 (N_2928,N_2824,N_2853);
or U2929 (N_2929,N_2849,N_2847);
nand U2930 (N_2930,N_2853,N_2842);
or U2931 (N_2931,N_2864,N_2876);
or U2932 (N_2932,N_2849,N_2842);
and U2933 (N_2933,N_2830,N_2821);
nor U2934 (N_2934,N_2856,N_2878);
nor U2935 (N_2935,N_2844,N_2858);
and U2936 (N_2936,N_2834,N_2861);
or U2937 (N_2937,N_2858,N_2874);
or U2938 (N_2938,N_2849,N_2874);
and U2939 (N_2939,N_2860,N_2835);
nor U2940 (N_2940,N_2933,N_2902);
nor U2941 (N_2941,N_2935,N_2920);
nand U2942 (N_2942,N_2937,N_2899);
nor U2943 (N_2943,N_2900,N_2918);
nand U2944 (N_2944,N_2910,N_2898);
nor U2945 (N_2945,N_2886,N_2883);
nor U2946 (N_2946,N_2885,N_2890);
nor U2947 (N_2947,N_2930,N_2911);
xnor U2948 (N_2948,N_2914,N_2889);
nand U2949 (N_2949,N_2906,N_2931);
nand U2950 (N_2950,N_2922,N_2925);
nor U2951 (N_2951,N_2887,N_2905);
and U2952 (N_2952,N_2891,N_2907);
nand U2953 (N_2953,N_2897,N_2904);
nand U2954 (N_2954,N_2896,N_2908);
nand U2955 (N_2955,N_2916,N_2884);
and U2956 (N_2956,N_2939,N_2926);
nor U2957 (N_2957,N_2880,N_2919);
nand U2958 (N_2958,N_2915,N_2938);
and U2959 (N_2959,N_2936,N_2903);
nand U2960 (N_2960,N_2934,N_2921);
or U2961 (N_2961,N_2924,N_2917);
nor U2962 (N_2962,N_2895,N_2929);
nor U2963 (N_2963,N_2882,N_2913);
or U2964 (N_2964,N_2894,N_2932);
nand U2965 (N_2965,N_2923,N_2909);
nand U2966 (N_2966,N_2928,N_2912);
and U2967 (N_2967,N_2888,N_2901);
and U2968 (N_2968,N_2927,N_2892);
xnor U2969 (N_2969,N_2881,N_2893);
or U2970 (N_2970,N_2897,N_2923);
or U2971 (N_2971,N_2929,N_2920);
or U2972 (N_2972,N_2932,N_2914);
nand U2973 (N_2973,N_2926,N_2921);
or U2974 (N_2974,N_2903,N_2893);
nor U2975 (N_2975,N_2887,N_2935);
nor U2976 (N_2976,N_2929,N_2921);
and U2977 (N_2977,N_2893,N_2920);
nor U2978 (N_2978,N_2934,N_2938);
or U2979 (N_2979,N_2893,N_2890);
nand U2980 (N_2980,N_2932,N_2930);
and U2981 (N_2981,N_2894,N_2935);
or U2982 (N_2982,N_2910,N_2917);
nand U2983 (N_2983,N_2938,N_2905);
nor U2984 (N_2984,N_2928,N_2890);
or U2985 (N_2985,N_2928,N_2888);
nor U2986 (N_2986,N_2918,N_2906);
and U2987 (N_2987,N_2896,N_2901);
or U2988 (N_2988,N_2922,N_2923);
xor U2989 (N_2989,N_2888,N_2916);
nor U2990 (N_2990,N_2925,N_2892);
and U2991 (N_2991,N_2912,N_2936);
and U2992 (N_2992,N_2889,N_2912);
or U2993 (N_2993,N_2883,N_2892);
or U2994 (N_2994,N_2902,N_2937);
and U2995 (N_2995,N_2890,N_2912);
and U2996 (N_2996,N_2914,N_2885);
or U2997 (N_2997,N_2912,N_2903);
or U2998 (N_2998,N_2891,N_2913);
nor U2999 (N_2999,N_2913,N_2901);
and UO_0 (O_0,N_2940,N_2958);
and UO_1 (O_1,N_2980,N_2962);
nor UO_2 (O_2,N_2944,N_2943);
nor UO_3 (O_3,N_2975,N_2990);
nand UO_4 (O_4,N_2967,N_2965);
and UO_5 (O_5,N_2970,N_2954);
and UO_6 (O_6,N_2966,N_2978);
nand UO_7 (O_7,N_2953,N_2963);
nor UO_8 (O_8,N_2957,N_2985);
or UO_9 (O_9,N_2952,N_2960);
nand UO_10 (O_10,N_2988,N_2947);
or UO_11 (O_11,N_2989,N_2976);
nand UO_12 (O_12,N_2997,N_2959);
and UO_13 (O_13,N_2992,N_2948);
nand UO_14 (O_14,N_2961,N_2986);
nor UO_15 (O_15,N_2968,N_2955);
nand UO_16 (O_16,N_2983,N_2977);
nand UO_17 (O_17,N_2971,N_2969);
and UO_18 (O_18,N_2941,N_2979);
or UO_19 (O_19,N_2995,N_2996);
nor UO_20 (O_20,N_2945,N_2942);
or UO_21 (O_21,N_2964,N_2956);
and UO_22 (O_22,N_2946,N_2972);
or UO_23 (O_23,N_2974,N_2987);
and UO_24 (O_24,N_2984,N_2994);
or UO_25 (O_25,N_2950,N_2999);
and UO_26 (O_26,N_2949,N_2998);
nor UO_27 (O_27,N_2991,N_2993);
and UO_28 (O_28,N_2973,N_2951);
nor UO_29 (O_29,N_2982,N_2981);
nand UO_30 (O_30,N_2976,N_2984);
or UO_31 (O_31,N_2957,N_2964);
or UO_32 (O_32,N_2983,N_2965);
nor UO_33 (O_33,N_2947,N_2986);
nand UO_34 (O_34,N_2971,N_2983);
nand UO_35 (O_35,N_2950,N_2974);
or UO_36 (O_36,N_2954,N_2973);
nor UO_37 (O_37,N_2957,N_2975);
nor UO_38 (O_38,N_2978,N_2952);
or UO_39 (O_39,N_2972,N_2966);
nand UO_40 (O_40,N_2954,N_2949);
nor UO_41 (O_41,N_2941,N_2993);
and UO_42 (O_42,N_2989,N_2992);
nor UO_43 (O_43,N_2969,N_2946);
nor UO_44 (O_44,N_2943,N_2958);
nand UO_45 (O_45,N_2989,N_2998);
or UO_46 (O_46,N_2973,N_2940);
and UO_47 (O_47,N_2990,N_2999);
or UO_48 (O_48,N_2943,N_2953);
nand UO_49 (O_49,N_2953,N_2955);
nor UO_50 (O_50,N_2941,N_2943);
nand UO_51 (O_51,N_2952,N_2986);
or UO_52 (O_52,N_2958,N_2971);
or UO_53 (O_53,N_2965,N_2976);
nor UO_54 (O_54,N_2969,N_2959);
nor UO_55 (O_55,N_2985,N_2952);
or UO_56 (O_56,N_2969,N_2955);
or UO_57 (O_57,N_2997,N_2981);
and UO_58 (O_58,N_2984,N_2942);
nand UO_59 (O_59,N_2987,N_2994);
or UO_60 (O_60,N_2961,N_2949);
nor UO_61 (O_61,N_2965,N_2990);
nor UO_62 (O_62,N_2972,N_2965);
and UO_63 (O_63,N_2972,N_2974);
or UO_64 (O_64,N_2974,N_2947);
nand UO_65 (O_65,N_2948,N_2977);
nand UO_66 (O_66,N_2945,N_2956);
or UO_67 (O_67,N_2986,N_2993);
nand UO_68 (O_68,N_2991,N_2955);
and UO_69 (O_69,N_2960,N_2954);
and UO_70 (O_70,N_2951,N_2995);
and UO_71 (O_71,N_2998,N_2945);
or UO_72 (O_72,N_2967,N_2984);
nor UO_73 (O_73,N_2950,N_2956);
and UO_74 (O_74,N_2962,N_2955);
and UO_75 (O_75,N_2973,N_2968);
and UO_76 (O_76,N_2971,N_2986);
or UO_77 (O_77,N_2943,N_2996);
or UO_78 (O_78,N_2992,N_2978);
nand UO_79 (O_79,N_2993,N_2988);
nand UO_80 (O_80,N_2946,N_2993);
nor UO_81 (O_81,N_2966,N_2961);
and UO_82 (O_82,N_2963,N_2987);
nand UO_83 (O_83,N_2969,N_2980);
nor UO_84 (O_84,N_2946,N_2986);
nand UO_85 (O_85,N_2992,N_2963);
nor UO_86 (O_86,N_2978,N_2993);
nand UO_87 (O_87,N_2980,N_2998);
nor UO_88 (O_88,N_2969,N_2985);
or UO_89 (O_89,N_2954,N_2966);
and UO_90 (O_90,N_2981,N_2964);
or UO_91 (O_91,N_2983,N_2989);
nand UO_92 (O_92,N_2943,N_2947);
nand UO_93 (O_93,N_2982,N_2974);
nand UO_94 (O_94,N_2996,N_2980);
and UO_95 (O_95,N_2966,N_2982);
nand UO_96 (O_96,N_2998,N_2992);
or UO_97 (O_97,N_2990,N_2988);
or UO_98 (O_98,N_2940,N_2990);
or UO_99 (O_99,N_2960,N_2979);
nand UO_100 (O_100,N_2940,N_2965);
nand UO_101 (O_101,N_2988,N_2958);
nor UO_102 (O_102,N_2981,N_2992);
and UO_103 (O_103,N_2981,N_2959);
nor UO_104 (O_104,N_2984,N_2954);
or UO_105 (O_105,N_2963,N_2985);
nor UO_106 (O_106,N_2955,N_2978);
nor UO_107 (O_107,N_2986,N_2974);
and UO_108 (O_108,N_2957,N_2965);
nor UO_109 (O_109,N_2966,N_2949);
nor UO_110 (O_110,N_2948,N_2946);
nor UO_111 (O_111,N_2964,N_2992);
nand UO_112 (O_112,N_2975,N_2949);
and UO_113 (O_113,N_2984,N_2949);
or UO_114 (O_114,N_2986,N_2948);
and UO_115 (O_115,N_2967,N_2972);
and UO_116 (O_116,N_2949,N_2979);
and UO_117 (O_117,N_2943,N_2946);
or UO_118 (O_118,N_2970,N_2984);
or UO_119 (O_119,N_2953,N_2996);
nor UO_120 (O_120,N_2986,N_2999);
and UO_121 (O_121,N_2954,N_2946);
and UO_122 (O_122,N_2973,N_2975);
or UO_123 (O_123,N_2996,N_2977);
nor UO_124 (O_124,N_2998,N_2966);
nand UO_125 (O_125,N_2987,N_2990);
nand UO_126 (O_126,N_2986,N_2953);
or UO_127 (O_127,N_2941,N_2973);
nor UO_128 (O_128,N_2943,N_2992);
nand UO_129 (O_129,N_2972,N_2970);
or UO_130 (O_130,N_2972,N_2994);
and UO_131 (O_131,N_2968,N_2947);
nand UO_132 (O_132,N_2976,N_2963);
and UO_133 (O_133,N_2992,N_2980);
nor UO_134 (O_134,N_2941,N_2991);
nand UO_135 (O_135,N_2990,N_2971);
and UO_136 (O_136,N_2999,N_2974);
and UO_137 (O_137,N_2942,N_2992);
nor UO_138 (O_138,N_2958,N_2982);
nor UO_139 (O_139,N_2941,N_2965);
and UO_140 (O_140,N_2947,N_2994);
and UO_141 (O_141,N_2944,N_2986);
and UO_142 (O_142,N_2958,N_2962);
or UO_143 (O_143,N_2990,N_2959);
and UO_144 (O_144,N_2964,N_2944);
nor UO_145 (O_145,N_2956,N_2991);
nand UO_146 (O_146,N_2945,N_2951);
or UO_147 (O_147,N_2985,N_2974);
and UO_148 (O_148,N_2960,N_2950);
nor UO_149 (O_149,N_2954,N_2944);
or UO_150 (O_150,N_2953,N_2972);
nor UO_151 (O_151,N_2940,N_2976);
nor UO_152 (O_152,N_2951,N_2965);
and UO_153 (O_153,N_2987,N_2950);
nor UO_154 (O_154,N_2971,N_2981);
or UO_155 (O_155,N_2977,N_2973);
nand UO_156 (O_156,N_2955,N_2948);
nand UO_157 (O_157,N_2959,N_2995);
and UO_158 (O_158,N_2971,N_2952);
nand UO_159 (O_159,N_2970,N_2979);
and UO_160 (O_160,N_2945,N_2941);
or UO_161 (O_161,N_2972,N_2951);
nor UO_162 (O_162,N_2974,N_2994);
nand UO_163 (O_163,N_2957,N_2978);
or UO_164 (O_164,N_2965,N_2955);
nand UO_165 (O_165,N_2947,N_2951);
and UO_166 (O_166,N_2945,N_2994);
nor UO_167 (O_167,N_2989,N_2956);
or UO_168 (O_168,N_2950,N_2958);
nor UO_169 (O_169,N_2959,N_2967);
nand UO_170 (O_170,N_2944,N_2961);
or UO_171 (O_171,N_2979,N_2958);
nor UO_172 (O_172,N_2983,N_2998);
nor UO_173 (O_173,N_2961,N_2975);
or UO_174 (O_174,N_2959,N_2955);
and UO_175 (O_175,N_2941,N_2958);
or UO_176 (O_176,N_2979,N_2995);
nor UO_177 (O_177,N_2994,N_2940);
nand UO_178 (O_178,N_2994,N_2955);
nand UO_179 (O_179,N_2947,N_2956);
or UO_180 (O_180,N_2946,N_2966);
nand UO_181 (O_181,N_2946,N_2999);
nor UO_182 (O_182,N_2960,N_2982);
and UO_183 (O_183,N_2946,N_2960);
and UO_184 (O_184,N_2954,N_2995);
and UO_185 (O_185,N_2987,N_2980);
nor UO_186 (O_186,N_2941,N_2969);
and UO_187 (O_187,N_2941,N_2948);
nand UO_188 (O_188,N_2947,N_2970);
or UO_189 (O_189,N_2987,N_2993);
and UO_190 (O_190,N_2996,N_2969);
and UO_191 (O_191,N_2967,N_2961);
and UO_192 (O_192,N_2951,N_2952);
or UO_193 (O_193,N_2992,N_2951);
nand UO_194 (O_194,N_2981,N_2960);
or UO_195 (O_195,N_2987,N_2968);
and UO_196 (O_196,N_2977,N_2945);
and UO_197 (O_197,N_2953,N_2976);
and UO_198 (O_198,N_2961,N_2997);
and UO_199 (O_199,N_2946,N_2944);
and UO_200 (O_200,N_2940,N_2983);
nand UO_201 (O_201,N_2952,N_2942);
and UO_202 (O_202,N_2984,N_2953);
and UO_203 (O_203,N_2982,N_2998);
and UO_204 (O_204,N_2940,N_2956);
nor UO_205 (O_205,N_2969,N_2992);
or UO_206 (O_206,N_2988,N_2991);
nor UO_207 (O_207,N_2972,N_2957);
or UO_208 (O_208,N_2967,N_2962);
nor UO_209 (O_209,N_2987,N_2959);
or UO_210 (O_210,N_2975,N_2940);
and UO_211 (O_211,N_2952,N_2984);
or UO_212 (O_212,N_2949,N_2994);
nor UO_213 (O_213,N_2970,N_2953);
or UO_214 (O_214,N_2982,N_2962);
or UO_215 (O_215,N_2941,N_2989);
nor UO_216 (O_216,N_2987,N_2978);
and UO_217 (O_217,N_2949,N_2976);
nor UO_218 (O_218,N_2961,N_2940);
nand UO_219 (O_219,N_2981,N_2940);
nand UO_220 (O_220,N_2969,N_2950);
nand UO_221 (O_221,N_2962,N_2945);
and UO_222 (O_222,N_2951,N_2956);
nor UO_223 (O_223,N_2956,N_2965);
and UO_224 (O_224,N_2944,N_2948);
and UO_225 (O_225,N_2960,N_2985);
nor UO_226 (O_226,N_2993,N_2949);
nand UO_227 (O_227,N_2999,N_2944);
or UO_228 (O_228,N_2985,N_2955);
or UO_229 (O_229,N_2970,N_2992);
or UO_230 (O_230,N_2979,N_2975);
or UO_231 (O_231,N_2965,N_2964);
and UO_232 (O_232,N_2987,N_2979);
nor UO_233 (O_233,N_2957,N_2983);
or UO_234 (O_234,N_2998,N_2981);
nor UO_235 (O_235,N_2985,N_2951);
and UO_236 (O_236,N_2993,N_2967);
or UO_237 (O_237,N_2977,N_2967);
or UO_238 (O_238,N_2962,N_2949);
and UO_239 (O_239,N_2983,N_2987);
nand UO_240 (O_240,N_2991,N_2945);
nor UO_241 (O_241,N_2999,N_2976);
and UO_242 (O_242,N_2946,N_2985);
and UO_243 (O_243,N_2963,N_2984);
or UO_244 (O_244,N_2940,N_2946);
nor UO_245 (O_245,N_2978,N_2963);
or UO_246 (O_246,N_2942,N_2996);
nor UO_247 (O_247,N_2949,N_2956);
and UO_248 (O_248,N_2976,N_2982);
nor UO_249 (O_249,N_2989,N_2953);
nand UO_250 (O_250,N_2945,N_2981);
and UO_251 (O_251,N_2962,N_2971);
nand UO_252 (O_252,N_2967,N_2956);
nand UO_253 (O_253,N_2999,N_2943);
nor UO_254 (O_254,N_2949,N_2970);
and UO_255 (O_255,N_2949,N_2951);
and UO_256 (O_256,N_2940,N_2954);
nand UO_257 (O_257,N_2947,N_2991);
nor UO_258 (O_258,N_2943,N_2986);
or UO_259 (O_259,N_2958,N_2992);
or UO_260 (O_260,N_2993,N_2960);
nor UO_261 (O_261,N_2956,N_2954);
nor UO_262 (O_262,N_2980,N_2958);
nor UO_263 (O_263,N_2989,N_2990);
nand UO_264 (O_264,N_2986,N_2957);
nand UO_265 (O_265,N_2997,N_2994);
and UO_266 (O_266,N_2941,N_2985);
nor UO_267 (O_267,N_2957,N_2979);
nand UO_268 (O_268,N_2984,N_2978);
nor UO_269 (O_269,N_2999,N_2965);
nor UO_270 (O_270,N_2945,N_2992);
nor UO_271 (O_271,N_2950,N_2986);
or UO_272 (O_272,N_2956,N_2993);
and UO_273 (O_273,N_2983,N_2985);
nand UO_274 (O_274,N_2956,N_2946);
nor UO_275 (O_275,N_2978,N_2956);
or UO_276 (O_276,N_2949,N_2960);
nand UO_277 (O_277,N_2988,N_2981);
and UO_278 (O_278,N_2970,N_2950);
nand UO_279 (O_279,N_2973,N_2972);
or UO_280 (O_280,N_2973,N_2947);
or UO_281 (O_281,N_2950,N_2985);
and UO_282 (O_282,N_2941,N_2964);
nor UO_283 (O_283,N_2990,N_2941);
nand UO_284 (O_284,N_2971,N_2988);
nor UO_285 (O_285,N_2982,N_2951);
nor UO_286 (O_286,N_2983,N_2967);
and UO_287 (O_287,N_2942,N_2997);
nand UO_288 (O_288,N_2965,N_2973);
nor UO_289 (O_289,N_2950,N_2964);
and UO_290 (O_290,N_2941,N_2963);
and UO_291 (O_291,N_2946,N_2996);
or UO_292 (O_292,N_2999,N_2977);
nand UO_293 (O_293,N_2953,N_2979);
nor UO_294 (O_294,N_2965,N_2966);
nor UO_295 (O_295,N_2989,N_2980);
nand UO_296 (O_296,N_2996,N_2993);
or UO_297 (O_297,N_2998,N_2946);
nand UO_298 (O_298,N_2991,N_2952);
or UO_299 (O_299,N_2949,N_2971);
nor UO_300 (O_300,N_2972,N_2999);
or UO_301 (O_301,N_2972,N_2996);
nor UO_302 (O_302,N_2970,N_2998);
or UO_303 (O_303,N_2942,N_2960);
or UO_304 (O_304,N_2987,N_2995);
nand UO_305 (O_305,N_2967,N_2948);
nor UO_306 (O_306,N_2948,N_2975);
nor UO_307 (O_307,N_2945,N_2961);
and UO_308 (O_308,N_2991,N_2981);
nor UO_309 (O_309,N_2957,N_2963);
xnor UO_310 (O_310,N_2980,N_2967);
nand UO_311 (O_311,N_2982,N_2961);
or UO_312 (O_312,N_2944,N_2974);
and UO_313 (O_313,N_2997,N_2996);
or UO_314 (O_314,N_2967,N_2994);
nor UO_315 (O_315,N_2944,N_2951);
nor UO_316 (O_316,N_2998,N_2953);
nand UO_317 (O_317,N_2967,N_2958);
or UO_318 (O_318,N_2941,N_2974);
and UO_319 (O_319,N_2964,N_2982);
nand UO_320 (O_320,N_2978,N_2946);
nand UO_321 (O_321,N_2950,N_2955);
nor UO_322 (O_322,N_2974,N_2979);
and UO_323 (O_323,N_2981,N_2948);
or UO_324 (O_324,N_2967,N_2952);
and UO_325 (O_325,N_2995,N_2992);
or UO_326 (O_326,N_2966,N_2956);
and UO_327 (O_327,N_2955,N_2980);
nand UO_328 (O_328,N_2978,N_2948);
nand UO_329 (O_329,N_2953,N_2987);
or UO_330 (O_330,N_2961,N_2990);
nor UO_331 (O_331,N_2964,N_2961);
and UO_332 (O_332,N_2951,N_2975);
nand UO_333 (O_333,N_2971,N_2980);
nor UO_334 (O_334,N_2970,N_2971);
and UO_335 (O_335,N_2949,N_2945);
nor UO_336 (O_336,N_2947,N_2950);
or UO_337 (O_337,N_2965,N_2998);
and UO_338 (O_338,N_2984,N_2955);
nor UO_339 (O_339,N_2963,N_2964);
xor UO_340 (O_340,N_2992,N_2941);
and UO_341 (O_341,N_2982,N_2940);
or UO_342 (O_342,N_2945,N_2943);
nand UO_343 (O_343,N_2957,N_2974);
nor UO_344 (O_344,N_2954,N_2993);
and UO_345 (O_345,N_2973,N_2963);
nor UO_346 (O_346,N_2991,N_2944);
nor UO_347 (O_347,N_2968,N_2942);
nand UO_348 (O_348,N_2997,N_2948);
or UO_349 (O_349,N_2970,N_2974);
nor UO_350 (O_350,N_2946,N_2990);
and UO_351 (O_351,N_2943,N_2942);
nor UO_352 (O_352,N_2992,N_2944);
or UO_353 (O_353,N_2978,N_2981);
and UO_354 (O_354,N_2981,N_2975);
and UO_355 (O_355,N_2993,N_2958);
or UO_356 (O_356,N_2962,N_2990);
nand UO_357 (O_357,N_2950,N_2972);
nor UO_358 (O_358,N_2941,N_2953);
nand UO_359 (O_359,N_2945,N_2984);
nand UO_360 (O_360,N_2951,N_2941);
nand UO_361 (O_361,N_2977,N_2981);
or UO_362 (O_362,N_2952,N_2974);
and UO_363 (O_363,N_2955,N_2945);
nand UO_364 (O_364,N_2978,N_2941);
xnor UO_365 (O_365,N_2964,N_2958);
or UO_366 (O_366,N_2967,N_2976);
or UO_367 (O_367,N_2972,N_2956);
nor UO_368 (O_368,N_2974,N_2969);
nor UO_369 (O_369,N_2952,N_2989);
or UO_370 (O_370,N_2996,N_2998);
and UO_371 (O_371,N_2979,N_2965);
nor UO_372 (O_372,N_2999,N_2958);
nand UO_373 (O_373,N_2999,N_2985);
nand UO_374 (O_374,N_2941,N_2983);
and UO_375 (O_375,N_2989,N_2964);
nor UO_376 (O_376,N_2995,N_2999);
nor UO_377 (O_377,N_2942,N_2954);
nor UO_378 (O_378,N_2992,N_2955);
or UO_379 (O_379,N_2989,N_2949);
or UO_380 (O_380,N_2952,N_2953);
nor UO_381 (O_381,N_2966,N_2967);
or UO_382 (O_382,N_2976,N_2980);
nor UO_383 (O_383,N_2990,N_2974);
nand UO_384 (O_384,N_2962,N_2963);
and UO_385 (O_385,N_2964,N_2980);
and UO_386 (O_386,N_2951,N_2940);
and UO_387 (O_387,N_2947,N_2993);
and UO_388 (O_388,N_2987,N_2955);
or UO_389 (O_389,N_2975,N_2992);
nor UO_390 (O_390,N_2981,N_2965);
nor UO_391 (O_391,N_2991,N_2967);
nor UO_392 (O_392,N_2972,N_2959);
nor UO_393 (O_393,N_2971,N_2987);
or UO_394 (O_394,N_2971,N_2978);
or UO_395 (O_395,N_2947,N_2980);
nand UO_396 (O_396,N_2970,N_2967);
nor UO_397 (O_397,N_2960,N_2983);
and UO_398 (O_398,N_2990,N_2942);
nor UO_399 (O_399,N_2993,N_2979);
and UO_400 (O_400,N_2959,N_2979);
and UO_401 (O_401,N_2974,N_2995);
or UO_402 (O_402,N_2955,N_2961);
nor UO_403 (O_403,N_2999,N_2973);
nor UO_404 (O_404,N_2961,N_2995);
or UO_405 (O_405,N_2979,N_2998);
or UO_406 (O_406,N_2990,N_2997);
or UO_407 (O_407,N_2988,N_2996);
nor UO_408 (O_408,N_2997,N_2943);
or UO_409 (O_409,N_2991,N_2960);
nor UO_410 (O_410,N_2964,N_2952);
and UO_411 (O_411,N_2984,N_2977);
nand UO_412 (O_412,N_2961,N_2968);
and UO_413 (O_413,N_2955,N_2946);
nor UO_414 (O_414,N_2973,N_2981);
nor UO_415 (O_415,N_2973,N_2996);
xnor UO_416 (O_416,N_2990,N_2954);
or UO_417 (O_417,N_2974,N_2943);
nor UO_418 (O_418,N_2959,N_2991);
nand UO_419 (O_419,N_2950,N_2961);
or UO_420 (O_420,N_2978,N_2986);
and UO_421 (O_421,N_2962,N_2994);
or UO_422 (O_422,N_2954,N_2998);
nand UO_423 (O_423,N_2964,N_2953);
nor UO_424 (O_424,N_2972,N_2942);
or UO_425 (O_425,N_2945,N_2953);
or UO_426 (O_426,N_2982,N_2955);
and UO_427 (O_427,N_2955,N_2966);
nor UO_428 (O_428,N_2980,N_2986);
nand UO_429 (O_429,N_2950,N_2995);
and UO_430 (O_430,N_2998,N_2961);
nor UO_431 (O_431,N_2985,N_2966);
or UO_432 (O_432,N_2982,N_2948);
and UO_433 (O_433,N_2966,N_2984);
nand UO_434 (O_434,N_2970,N_2993);
or UO_435 (O_435,N_2943,N_2948);
nand UO_436 (O_436,N_2982,N_2972);
nand UO_437 (O_437,N_2978,N_2999);
nand UO_438 (O_438,N_2945,N_2980);
nand UO_439 (O_439,N_2942,N_2986);
and UO_440 (O_440,N_2984,N_2985);
and UO_441 (O_441,N_2983,N_2979);
and UO_442 (O_442,N_2995,N_2997);
nor UO_443 (O_443,N_2972,N_2961);
or UO_444 (O_444,N_2947,N_2996);
or UO_445 (O_445,N_2988,N_2968);
nor UO_446 (O_446,N_2964,N_2960);
and UO_447 (O_447,N_2972,N_2962);
nor UO_448 (O_448,N_2977,N_2993);
and UO_449 (O_449,N_2970,N_2997);
and UO_450 (O_450,N_2942,N_2961);
nor UO_451 (O_451,N_2943,N_2956);
nor UO_452 (O_452,N_2968,N_2978);
nor UO_453 (O_453,N_2986,N_2966);
nor UO_454 (O_454,N_2955,N_2976);
nand UO_455 (O_455,N_2999,N_2957);
or UO_456 (O_456,N_2977,N_2961);
nand UO_457 (O_457,N_2980,N_2990);
or UO_458 (O_458,N_2966,N_2941);
nand UO_459 (O_459,N_2962,N_2954);
nand UO_460 (O_460,N_2947,N_2990);
and UO_461 (O_461,N_2947,N_2997);
nor UO_462 (O_462,N_2949,N_2942);
or UO_463 (O_463,N_2957,N_2977);
nand UO_464 (O_464,N_2986,N_2956);
nand UO_465 (O_465,N_2982,N_2977);
nor UO_466 (O_466,N_2989,N_2999);
or UO_467 (O_467,N_2970,N_2948);
or UO_468 (O_468,N_2960,N_2961);
nor UO_469 (O_469,N_2983,N_2975);
and UO_470 (O_470,N_2946,N_2979);
nor UO_471 (O_471,N_2994,N_2943);
nor UO_472 (O_472,N_2968,N_2990);
nor UO_473 (O_473,N_2992,N_2967);
nor UO_474 (O_474,N_2954,N_2961);
nand UO_475 (O_475,N_2948,N_2990);
nor UO_476 (O_476,N_2993,N_2959);
or UO_477 (O_477,N_2975,N_2997);
or UO_478 (O_478,N_2998,N_2960);
nor UO_479 (O_479,N_2986,N_2982);
or UO_480 (O_480,N_2967,N_2971);
and UO_481 (O_481,N_2954,N_2977);
nor UO_482 (O_482,N_2985,N_2954);
or UO_483 (O_483,N_2955,N_2979);
nand UO_484 (O_484,N_2983,N_2992);
nor UO_485 (O_485,N_2976,N_2987);
or UO_486 (O_486,N_2971,N_2950);
xor UO_487 (O_487,N_2945,N_2963);
nor UO_488 (O_488,N_2970,N_2988);
and UO_489 (O_489,N_2989,N_2961);
or UO_490 (O_490,N_2970,N_2982);
xor UO_491 (O_491,N_2958,N_2944);
nand UO_492 (O_492,N_2985,N_2942);
nor UO_493 (O_493,N_2960,N_2972);
nor UO_494 (O_494,N_2978,N_2983);
nor UO_495 (O_495,N_2954,N_2972);
nor UO_496 (O_496,N_2980,N_2994);
or UO_497 (O_497,N_2986,N_2940);
nor UO_498 (O_498,N_2951,N_2966);
nand UO_499 (O_499,N_2943,N_2961);
endmodule