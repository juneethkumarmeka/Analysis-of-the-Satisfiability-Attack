module basic_500_3000_500_60_levels_1xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_158,In_476);
or U1 (N_1,In_141,In_401);
nor U2 (N_2,In_102,In_246);
nor U3 (N_3,In_277,In_486);
and U4 (N_4,In_441,In_323);
nand U5 (N_5,In_87,In_301);
nor U6 (N_6,In_25,In_260);
or U7 (N_7,In_494,In_342);
or U8 (N_8,In_411,In_1);
nand U9 (N_9,In_393,In_202);
nor U10 (N_10,In_49,In_495);
and U11 (N_11,In_354,In_251);
or U12 (N_12,In_20,In_402);
nor U13 (N_13,In_430,In_168);
nor U14 (N_14,In_465,In_250);
nand U15 (N_15,In_57,In_155);
nor U16 (N_16,In_304,In_24);
and U17 (N_17,In_473,In_311);
or U18 (N_18,In_159,In_103);
nor U19 (N_19,In_109,In_409);
nand U20 (N_20,In_172,In_468);
or U21 (N_21,In_435,In_208);
or U22 (N_22,In_429,In_188);
nor U23 (N_23,In_197,In_222);
or U24 (N_24,In_252,In_330);
nand U25 (N_25,In_297,In_193);
or U26 (N_26,In_77,In_366);
nand U27 (N_27,In_329,In_167);
nor U28 (N_28,In_205,In_358);
nand U29 (N_29,In_387,In_209);
and U30 (N_30,In_313,In_198);
nor U31 (N_31,In_258,In_477);
nor U32 (N_32,In_284,In_433);
nand U33 (N_33,In_51,In_458);
or U34 (N_34,In_32,In_471);
and U35 (N_35,In_307,In_444);
and U36 (N_36,In_448,In_418);
nor U37 (N_37,In_230,In_177);
or U38 (N_38,In_162,In_244);
nand U39 (N_39,In_12,In_455);
nor U40 (N_40,In_275,In_247);
nor U41 (N_41,In_175,In_136);
nor U42 (N_42,In_64,In_82);
nand U43 (N_43,In_83,In_100);
nor U44 (N_44,In_176,In_427);
or U45 (N_45,In_368,In_319);
nor U46 (N_46,In_178,In_376);
nor U47 (N_47,In_219,In_68);
nor U48 (N_48,In_104,In_55);
nor U49 (N_49,In_273,In_328);
and U50 (N_50,In_333,In_43);
nor U51 (N_51,In_388,In_496);
nor U52 (N_52,In_443,In_10);
nand U53 (N_53,In_90,In_293);
xor U54 (N_54,In_254,In_460);
nand U55 (N_55,In_54,In_279);
or U56 (N_56,N_41,In_417);
nand U57 (N_57,N_25,N_4);
nand U58 (N_58,In_271,In_361);
nor U59 (N_59,In_152,In_288);
nor U60 (N_60,N_49,In_404);
nor U61 (N_61,In_78,In_351);
nand U62 (N_62,In_299,In_239);
or U63 (N_63,In_373,In_144);
or U64 (N_64,In_28,In_326);
nand U65 (N_65,In_223,N_32);
and U66 (N_66,In_154,N_28);
and U67 (N_67,In_370,In_186);
and U68 (N_68,In_105,N_5);
or U69 (N_69,In_332,In_220);
nand U70 (N_70,In_436,In_62);
or U71 (N_71,N_35,In_462);
nor U72 (N_72,In_470,In_201);
and U73 (N_73,In_353,In_286);
or U74 (N_74,In_298,In_335);
nor U75 (N_75,N_8,In_425);
nand U76 (N_76,In_497,In_243);
nand U77 (N_77,In_121,In_189);
and U78 (N_78,In_161,In_337);
nor U79 (N_79,N_34,In_467);
or U80 (N_80,In_253,In_327);
nor U81 (N_81,In_117,In_280);
and U82 (N_82,In_127,In_97);
nand U83 (N_83,In_445,In_287);
nor U84 (N_84,In_157,In_18);
and U85 (N_85,In_461,In_169);
nor U86 (N_86,In_142,In_281);
nand U87 (N_87,In_384,In_389);
or U88 (N_88,In_80,In_40);
nor U89 (N_89,In_416,N_27);
or U90 (N_90,In_67,In_428);
and U91 (N_91,In_15,In_295);
and U92 (N_92,In_400,In_475);
nor U93 (N_93,In_75,N_17);
nor U94 (N_94,In_382,In_99);
or U95 (N_95,In_65,In_122);
nor U96 (N_96,In_283,In_89);
or U97 (N_97,In_94,In_480);
nand U98 (N_98,In_294,N_0);
xor U99 (N_99,In_211,In_124);
and U100 (N_100,In_199,In_255);
nand U101 (N_101,In_360,In_414);
nand U102 (N_102,In_282,N_96);
and U103 (N_103,In_432,N_86);
or U104 (N_104,In_215,In_14);
nor U105 (N_105,N_18,In_196);
nand U106 (N_106,In_314,In_58);
nor U107 (N_107,In_482,In_276);
or U108 (N_108,In_133,In_101);
nand U109 (N_109,In_146,In_268);
and U110 (N_110,In_320,In_372);
nand U111 (N_111,In_344,In_108);
or U112 (N_112,In_35,N_2);
or U113 (N_113,N_57,In_61);
nor U114 (N_114,N_75,In_120);
or U115 (N_115,In_9,In_347);
and U116 (N_116,N_7,In_406);
nand U117 (N_117,N_11,In_262);
and U118 (N_118,In_21,In_138);
or U119 (N_119,N_58,In_378);
and U120 (N_120,N_40,In_363);
nand U121 (N_121,In_207,In_11);
nor U122 (N_122,N_38,In_278);
and U123 (N_123,In_259,In_221);
and U124 (N_124,In_70,In_339);
or U125 (N_125,In_464,In_424);
nand U126 (N_126,In_426,In_180);
or U127 (N_127,In_86,N_39);
or U128 (N_128,In_466,In_390);
and U129 (N_129,In_423,In_463);
nand U130 (N_130,N_92,In_257);
or U131 (N_131,In_130,N_94);
nor U132 (N_132,In_371,N_22);
nor U133 (N_133,N_30,In_8);
xnor U134 (N_134,In_148,In_179);
nor U135 (N_135,In_302,In_398);
nor U136 (N_136,In_274,N_14);
nand U137 (N_137,In_454,In_79);
nor U138 (N_138,In_194,In_449);
nor U139 (N_139,N_47,N_19);
nor U140 (N_140,In_397,N_9);
or U141 (N_141,In_47,In_212);
nand U142 (N_142,N_62,In_334);
and U143 (N_143,N_81,In_153);
and U144 (N_144,In_434,In_399);
nand U145 (N_145,In_410,In_217);
nor U146 (N_146,In_362,N_54);
or U147 (N_147,In_93,N_44);
nor U148 (N_148,In_116,In_234);
and U149 (N_149,In_340,N_66);
nor U150 (N_150,N_84,N_97);
and U151 (N_151,In_45,N_6);
and U152 (N_152,In_22,In_156);
nor U153 (N_153,In_149,N_144);
nand U154 (N_154,In_346,N_99);
nand U155 (N_155,In_30,In_349);
nor U156 (N_156,In_171,In_487);
or U157 (N_157,In_27,In_377);
nor U158 (N_158,In_63,In_266);
nor U159 (N_159,In_126,N_69);
nand U160 (N_160,N_53,N_24);
nand U161 (N_161,N_149,In_488);
and U162 (N_162,In_394,In_160);
nor U163 (N_163,In_345,N_109);
nand U164 (N_164,In_137,In_383);
nand U165 (N_165,In_73,In_492);
or U166 (N_166,N_141,In_272);
or U167 (N_167,N_67,N_107);
and U168 (N_168,In_364,In_413);
or U169 (N_169,In_439,N_10);
nand U170 (N_170,In_147,In_42);
nor U171 (N_171,N_63,In_5);
nor U172 (N_172,In_34,N_77);
or U173 (N_173,In_249,In_459);
nor U174 (N_174,In_264,N_126);
nand U175 (N_175,N_88,N_89);
nand U176 (N_176,In_483,N_76);
or U177 (N_177,In_407,N_115);
nand U178 (N_178,N_122,In_195);
nor U179 (N_179,N_143,In_485);
nand U180 (N_180,N_105,N_79);
and U181 (N_181,In_318,In_131);
and U182 (N_182,In_292,In_107);
or U183 (N_183,In_269,In_182);
nand U184 (N_184,In_392,In_60);
nand U185 (N_185,N_106,In_452);
and U186 (N_186,N_145,In_412);
nand U187 (N_187,In_421,In_106);
or U188 (N_188,In_395,N_93);
or U189 (N_189,In_469,In_74);
nand U190 (N_190,In_232,In_96);
and U191 (N_191,N_100,In_484);
nand U192 (N_192,In_355,In_491);
nand U193 (N_193,In_237,In_256);
nor U194 (N_194,In_479,N_56);
nor U195 (N_195,In_343,In_151);
nor U196 (N_196,In_490,N_139);
nor U197 (N_197,In_129,N_20);
nand U198 (N_198,In_300,In_396);
nor U199 (N_199,In_312,N_131);
or U200 (N_200,In_405,N_52);
nand U201 (N_201,N_192,In_38);
and U202 (N_202,N_29,In_69);
nand U203 (N_203,In_350,In_308);
and U204 (N_204,In_306,In_84);
nand U205 (N_205,In_218,N_199);
nor U206 (N_206,N_110,In_325);
or U207 (N_207,In_71,In_123);
or U208 (N_208,N_26,N_135);
nor U209 (N_209,In_270,N_64);
or U210 (N_210,N_162,N_48);
nand U211 (N_211,In_29,In_164);
nor U212 (N_212,N_118,N_158);
and U213 (N_213,In_446,N_65);
nor U214 (N_214,In_310,In_191);
or U215 (N_215,N_154,N_113);
nand U216 (N_216,N_151,In_39);
and U217 (N_217,N_159,N_71);
or U218 (N_218,In_375,In_303);
or U219 (N_219,In_145,In_26);
nor U220 (N_220,In_98,In_231);
and U221 (N_221,N_168,In_111);
nor U222 (N_222,In_50,In_37);
or U223 (N_223,In_419,In_324);
or U224 (N_224,N_187,In_224);
nand U225 (N_225,In_381,In_7);
and U226 (N_226,N_129,N_70);
or U227 (N_227,In_489,In_2);
nor U228 (N_228,In_115,N_166);
nor U229 (N_229,N_55,N_3);
and U230 (N_230,In_261,In_163);
nand U231 (N_231,N_156,In_336);
nor U232 (N_232,In_17,In_72);
nor U233 (N_233,In_296,In_369);
and U234 (N_234,N_23,In_357);
nand U235 (N_235,In_13,N_175);
nand U236 (N_236,N_37,In_309);
and U237 (N_237,N_147,In_19);
or U238 (N_238,In_236,In_190);
nand U239 (N_239,N_13,N_108);
nand U240 (N_240,N_153,In_499);
nor U241 (N_241,In_474,N_138);
nand U242 (N_242,In_331,N_160);
nor U243 (N_243,N_87,In_213);
and U244 (N_244,In_315,In_379);
nand U245 (N_245,In_216,N_82);
and U246 (N_246,In_134,In_173);
and U247 (N_247,In_265,N_102);
or U248 (N_248,In_235,N_190);
or U249 (N_249,N_152,In_317);
or U250 (N_250,N_228,N_136);
nand U251 (N_251,N_121,N_123);
nand U252 (N_252,In_385,N_91);
nand U253 (N_253,In_359,N_200);
nor U254 (N_254,N_111,N_165);
nor U255 (N_255,In_227,N_161);
nor U256 (N_256,N_197,N_220);
nor U257 (N_257,N_193,In_132);
and U258 (N_258,N_134,In_91);
or U259 (N_259,In_348,In_457);
nand U260 (N_260,N_98,N_195);
nor U261 (N_261,In_316,N_172);
nor U262 (N_262,In_31,In_447);
and U263 (N_263,N_120,In_187);
nor U264 (N_264,N_60,N_246);
or U265 (N_265,In_66,In_85);
nand U266 (N_266,In_181,N_185);
nand U267 (N_267,N_191,In_263);
nand U268 (N_268,N_217,N_244);
nand U269 (N_269,N_101,N_21);
and U270 (N_270,In_165,N_51);
nand U271 (N_271,In_143,N_61);
nand U272 (N_272,In_23,N_237);
nor U273 (N_273,N_177,In_192);
nand U274 (N_274,N_178,In_472);
nand U275 (N_275,N_181,N_157);
nor U276 (N_276,N_95,In_226);
nor U277 (N_277,N_208,In_33);
nor U278 (N_278,In_140,N_203);
or U279 (N_279,N_132,N_125);
nor U280 (N_280,N_194,N_234);
nand U281 (N_281,In_498,In_185);
nor U282 (N_282,N_229,N_31);
or U283 (N_283,In_174,In_380);
nor U284 (N_284,N_206,In_59);
nand U285 (N_285,N_249,In_95);
or U286 (N_286,N_179,N_73);
nor U287 (N_287,In_135,N_45);
and U288 (N_288,In_440,In_241);
or U289 (N_289,N_128,In_238);
nand U290 (N_290,N_50,N_242);
nand U291 (N_291,In_3,In_233);
and U292 (N_292,N_72,N_198);
nand U293 (N_293,In_119,N_146);
or U294 (N_294,N_16,N_224);
nor U295 (N_295,In_48,N_245);
nor U296 (N_296,N_116,N_189);
or U297 (N_297,In_92,In_403);
and U298 (N_298,N_12,N_186);
and U299 (N_299,N_114,N_80);
nor U300 (N_300,N_119,In_184);
or U301 (N_301,N_280,N_238);
nand U302 (N_302,N_222,In_112);
and U303 (N_303,N_216,In_41);
nand U304 (N_304,In_150,N_271);
nor U305 (N_305,In_166,N_276);
or U306 (N_306,In_46,In_170);
nand U307 (N_307,N_140,N_205);
and U308 (N_308,N_15,N_137);
and U309 (N_309,In_4,N_293);
nand U310 (N_310,In_352,In_305);
nor U311 (N_311,In_229,In_114);
nor U312 (N_312,In_415,N_174);
nor U313 (N_313,In_242,N_256);
or U314 (N_314,N_207,N_223);
and U315 (N_315,In_53,N_142);
and U316 (N_316,In_289,N_42);
nand U317 (N_317,In_110,In_128);
nand U318 (N_318,In_125,N_171);
or U319 (N_319,N_215,N_270);
or U320 (N_320,N_167,In_442);
nand U321 (N_321,In_391,N_133);
nor U322 (N_322,In_88,In_36);
or U323 (N_323,N_74,N_210);
or U324 (N_324,N_279,In_374);
or U325 (N_325,N_112,N_231);
and U326 (N_326,N_204,N_252);
or U327 (N_327,N_267,N_46);
or U328 (N_328,N_201,N_265);
nor U329 (N_329,N_188,In_408);
or U330 (N_330,N_212,N_291);
nand U331 (N_331,In_245,N_1);
nor U332 (N_332,N_273,In_214);
nand U333 (N_333,N_281,In_450);
xnor U334 (N_334,N_184,In_200);
or U335 (N_335,N_127,N_227);
nor U336 (N_336,N_258,N_247);
nor U337 (N_337,In_285,In_56);
and U338 (N_338,In_322,N_278);
nor U339 (N_339,N_43,N_248);
or U340 (N_340,N_274,N_68);
or U341 (N_341,In_16,N_298);
and U342 (N_342,N_148,In_118);
nor U343 (N_343,In_210,N_36);
nor U344 (N_344,N_103,N_226);
nand U345 (N_345,N_290,N_173);
or U346 (N_346,In_6,N_272);
and U347 (N_347,N_183,N_176);
and U348 (N_348,In_356,N_251);
or U349 (N_349,In_481,N_236);
nor U350 (N_350,N_318,In_321);
nand U351 (N_351,N_232,N_235);
nor U352 (N_352,N_240,N_196);
and U353 (N_353,N_329,In_206);
nand U354 (N_354,N_346,N_301);
nor U355 (N_355,In_183,N_338);
nand U356 (N_356,N_297,N_317);
or U357 (N_357,N_349,N_259);
nor U358 (N_358,N_241,N_261);
nand U359 (N_359,In_113,N_283);
and U360 (N_360,In_76,In_456);
and U361 (N_361,In_453,N_221);
or U362 (N_362,N_250,N_330);
nor U363 (N_363,N_322,N_150);
nand U364 (N_364,N_257,In_52);
or U365 (N_365,N_343,N_263);
xor U366 (N_366,N_305,N_341);
and U367 (N_367,N_255,N_304);
nor U368 (N_368,In_291,N_308);
nand U369 (N_369,In_267,N_312);
nor U370 (N_370,In_248,N_243);
nor U371 (N_371,In_367,N_316);
and U372 (N_372,N_287,In_203);
nand U373 (N_373,N_307,N_83);
nor U374 (N_374,In_451,N_294);
and U375 (N_375,N_170,N_269);
nor U376 (N_376,N_306,In_493);
nor U377 (N_377,N_117,N_296);
or U378 (N_378,In_338,In_81);
nand U379 (N_379,N_59,N_299);
and U380 (N_380,N_285,In_139);
nor U381 (N_381,N_303,N_85);
nand U382 (N_382,N_319,N_275);
nor U383 (N_383,N_321,N_347);
or U384 (N_384,N_302,N_180);
nor U385 (N_385,N_230,N_218);
nor U386 (N_386,N_345,N_337);
nand U387 (N_387,N_164,N_155);
or U388 (N_388,N_266,N_326);
or U389 (N_389,N_264,N_311);
nand U390 (N_390,N_325,N_292);
and U391 (N_391,N_277,In_44);
nor U392 (N_392,In_0,N_348);
nor U393 (N_393,N_334,N_233);
nor U394 (N_394,N_104,N_90);
nor U395 (N_395,N_323,N_284);
nand U396 (N_396,N_310,In_438);
and U397 (N_397,N_288,N_328);
or U398 (N_398,In_225,In_240);
or U399 (N_399,N_219,N_331);
or U400 (N_400,N_351,N_390);
or U401 (N_401,N_327,N_182);
nand U402 (N_402,N_253,N_225);
and U403 (N_403,N_356,N_391);
nand U404 (N_404,N_239,N_363);
nor U405 (N_405,N_361,N_362);
or U406 (N_406,In_341,N_209);
and U407 (N_407,N_397,N_392);
and U408 (N_408,N_377,N_369);
nand U409 (N_409,N_262,In_365);
and U410 (N_410,N_395,In_431);
nor U411 (N_411,N_324,N_352);
nor U412 (N_412,N_371,N_211);
and U413 (N_413,N_393,N_332);
xor U414 (N_414,N_344,N_385);
nor U415 (N_415,N_295,N_376);
nand U416 (N_416,N_214,N_260);
or U417 (N_417,N_357,N_124);
nor U418 (N_418,N_358,N_309);
nor U419 (N_419,N_374,N_388);
nand U420 (N_420,N_289,N_384);
nor U421 (N_421,N_370,N_339);
and U422 (N_422,N_396,N_314);
nor U423 (N_423,N_336,N_386);
nor U424 (N_424,In_290,N_383);
nor U425 (N_425,N_202,N_367);
or U426 (N_426,In_437,N_333);
and U427 (N_427,N_300,In_204);
or U428 (N_428,N_342,N_373);
nor U429 (N_429,N_254,N_213);
nor U430 (N_430,N_335,In_228);
nand U431 (N_431,N_387,N_372);
nor U432 (N_432,N_375,N_380);
xnor U433 (N_433,In_478,N_398);
and U434 (N_434,N_354,N_389);
or U435 (N_435,N_394,N_268);
or U436 (N_436,N_33,N_366);
nand U437 (N_437,N_315,N_282);
and U438 (N_438,N_163,N_399);
nand U439 (N_439,N_78,N_130);
nand U440 (N_440,N_364,N_340);
and U441 (N_441,N_169,In_420);
nor U442 (N_442,N_379,N_353);
and U443 (N_443,N_313,N_360);
nand U444 (N_444,N_365,N_359);
and U445 (N_445,N_350,N_378);
and U446 (N_446,In_422,N_355);
nand U447 (N_447,N_381,In_386);
nor U448 (N_448,N_382,N_286);
or U449 (N_449,N_320,N_368);
nand U450 (N_450,N_409,N_404);
nand U451 (N_451,N_445,N_426);
nand U452 (N_452,N_408,N_420);
nand U453 (N_453,N_405,N_438);
or U454 (N_454,N_434,N_430);
nor U455 (N_455,N_435,N_441);
or U456 (N_456,N_436,N_444);
and U457 (N_457,N_412,N_414);
nand U458 (N_458,N_433,N_400);
or U459 (N_459,N_440,N_402);
nand U460 (N_460,N_417,N_421);
or U461 (N_461,N_422,N_428);
and U462 (N_462,N_447,N_429);
nand U463 (N_463,N_427,N_415);
and U464 (N_464,N_411,N_437);
nand U465 (N_465,N_439,N_443);
nor U466 (N_466,N_401,N_403);
nand U467 (N_467,N_442,N_449);
nand U468 (N_468,N_431,N_425);
or U469 (N_469,N_448,N_406);
and U470 (N_470,N_423,N_413);
nand U471 (N_471,N_419,N_416);
and U472 (N_472,N_410,N_446);
nor U473 (N_473,N_432,N_418);
nand U474 (N_474,N_424,N_407);
or U475 (N_475,N_445,N_432);
nor U476 (N_476,N_447,N_441);
and U477 (N_477,N_406,N_415);
nor U478 (N_478,N_444,N_418);
nor U479 (N_479,N_415,N_426);
nor U480 (N_480,N_438,N_404);
nor U481 (N_481,N_437,N_443);
or U482 (N_482,N_405,N_443);
and U483 (N_483,N_414,N_400);
nor U484 (N_484,N_428,N_443);
or U485 (N_485,N_412,N_426);
nand U486 (N_486,N_411,N_443);
nor U487 (N_487,N_409,N_438);
or U488 (N_488,N_428,N_411);
or U489 (N_489,N_439,N_400);
or U490 (N_490,N_409,N_423);
or U491 (N_491,N_439,N_420);
nor U492 (N_492,N_419,N_413);
and U493 (N_493,N_429,N_424);
or U494 (N_494,N_435,N_417);
or U495 (N_495,N_402,N_414);
nor U496 (N_496,N_404,N_447);
nor U497 (N_497,N_431,N_443);
and U498 (N_498,N_446,N_414);
nand U499 (N_499,N_400,N_412);
and U500 (N_500,N_493,N_483);
or U501 (N_501,N_491,N_481);
and U502 (N_502,N_466,N_474);
nand U503 (N_503,N_470,N_475);
xnor U504 (N_504,N_486,N_488);
nor U505 (N_505,N_487,N_465);
or U506 (N_506,N_456,N_479);
nand U507 (N_507,N_496,N_460);
or U508 (N_508,N_477,N_469);
nor U509 (N_509,N_499,N_482);
nand U510 (N_510,N_492,N_476);
or U511 (N_511,N_478,N_457);
or U512 (N_512,N_480,N_472);
and U513 (N_513,N_497,N_468);
or U514 (N_514,N_452,N_495);
and U515 (N_515,N_494,N_485);
and U516 (N_516,N_467,N_463);
or U517 (N_517,N_473,N_489);
nor U518 (N_518,N_459,N_484);
nor U519 (N_519,N_450,N_454);
nand U520 (N_520,N_462,N_451);
and U521 (N_521,N_458,N_490);
or U522 (N_522,N_471,N_498);
nand U523 (N_523,N_461,N_453);
and U524 (N_524,N_464,N_455);
nand U525 (N_525,N_480,N_483);
nand U526 (N_526,N_496,N_451);
nor U527 (N_527,N_481,N_475);
and U528 (N_528,N_496,N_475);
or U529 (N_529,N_450,N_480);
nor U530 (N_530,N_454,N_469);
nand U531 (N_531,N_481,N_452);
nor U532 (N_532,N_498,N_454);
nor U533 (N_533,N_483,N_472);
nor U534 (N_534,N_465,N_481);
nand U535 (N_535,N_489,N_488);
nor U536 (N_536,N_485,N_450);
nand U537 (N_537,N_490,N_470);
and U538 (N_538,N_482,N_466);
nand U539 (N_539,N_458,N_468);
or U540 (N_540,N_492,N_472);
or U541 (N_541,N_498,N_452);
nor U542 (N_542,N_455,N_454);
nand U543 (N_543,N_497,N_477);
or U544 (N_544,N_485,N_483);
or U545 (N_545,N_456,N_485);
or U546 (N_546,N_469,N_451);
and U547 (N_547,N_457,N_490);
and U548 (N_548,N_471,N_476);
and U549 (N_549,N_456,N_481);
nor U550 (N_550,N_525,N_530);
or U551 (N_551,N_502,N_526);
nor U552 (N_552,N_528,N_518);
nor U553 (N_553,N_542,N_515);
and U554 (N_554,N_521,N_523);
and U555 (N_555,N_503,N_514);
nor U556 (N_556,N_541,N_548);
nand U557 (N_557,N_533,N_504);
and U558 (N_558,N_511,N_501);
xor U559 (N_559,N_507,N_546);
or U560 (N_560,N_538,N_520);
or U561 (N_561,N_519,N_539);
nand U562 (N_562,N_506,N_505);
and U563 (N_563,N_508,N_522);
nor U564 (N_564,N_537,N_549);
nand U565 (N_565,N_527,N_531);
and U566 (N_566,N_544,N_524);
or U567 (N_567,N_536,N_500);
or U568 (N_568,N_540,N_510);
nor U569 (N_569,N_532,N_545);
and U570 (N_570,N_516,N_535);
nand U571 (N_571,N_534,N_517);
and U572 (N_572,N_529,N_513);
nand U573 (N_573,N_543,N_509);
nand U574 (N_574,N_547,N_512);
nand U575 (N_575,N_537,N_535);
nand U576 (N_576,N_542,N_545);
and U577 (N_577,N_509,N_540);
and U578 (N_578,N_528,N_530);
nand U579 (N_579,N_526,N_549);
nand U580 (N_580,N_543,N_544);
nand U581 (N_581,N_504,N_508);
and U582 (N_582,N_519,N_517);
nor U583 (N_583,N_547,N_549);
or U584 (N_584,N_509,N_539);
or U585 (N_585,N_501,N_532);
nor U586 (N_586,N_531,N_522);
nand U587 (N_587,N_510,N_547);
nor U588 (N_588,N_528,N_516);
nor U589 (N_589,N_505,N_508);
or U590 (N_590,N_512,N_513);
nor U591 (N_591,N_528,N_510);
and U592 (N_592,N_500,N_541);
or U593 (N_593,N_502,N_541);
nand U594 (N_594,N_527,N_540);
nand U595 (N_595,N_549,N_511);
or U596 (N_596,N_510,N_541);
nor U597 (N_597,N_545,N_526);
or U598 (N_598,N_548,N_529);
nand U599 (N_599,N_507,N_510);
or U600 (N_600,N_577,N_558);
or U601 (N_601,N_578,N_586);
or U602 (N_602,N_593,N_582);
nor U603 (N_603,N_599,N_560);
and U604 (N_604,N_567,N_557);
and U605 (N_605,N_581,N_565);
or U606 (N_606,N_573,N_563);
and U607 (N_607,N_597,N_564);
nor U608 (N_608,N_595,N_590);
and U609 (N_609,N_580,N_575);
or U610 (N_610,N_589,N_550);
nand U611 (N_611,N_562,N_587);
or U612 (N_612,N_584,N_556);
and U613 (N_613,N_588,N_561);
and U614 (N_614,N_574,N_583);
nand U615 (N_615,N_570,N_572);
and U616 (N_616,N_553,N_568);
nand U617 (N_617,N_585,N_551);
nor U618 (N_618,N_594,N_576);
or U619 (N_619,N_579,N_591);
nand U620 (N_620,N_571,N_566);
nand U621 (N_621,N_592,N_552);
nor U622 (N_622,N_598,N_569);
or U623 (N_623,N_596,N_555);
nor U624 (N_624,N_554,N_559);
and U625 (N_625,N_559,N_561);
or U626 (N_626,N_558,N_598);
and U627 (N_627,N_584,N_593);
nand U628 (N_628,N_577,N_551);
and U629 (N_629,N_574,N_563);
and U630 (N_630,N_578,N_580);
and U631 (N_631,N_572,N_557);
xor U632 (N_632,N_554,N_585);
and U633 (N_633,N_595,N_567);
nand U634 (N_634,N_572,N_565);
and U635 (N_635,N_564,N_563);
or U636 (N_636,N_575,N_552);
or U637 (N_637,N_588,N_581);
nor U638 (N_638,N_598,N_571);
nor U639 (N_639,N_595,N_579);
and U640 (N_640,N_595,N_583);
or U641 (N_641,N_557,N_582);
or U642 (N_642,N_560,N_589);
or U643 (N_643,N_554,N_577);
nand U644 (N_644,N_559,N_597);
or U645 (N_645,N_567,N_586);
nor U646 (N_646,N_588,N_559);
and U647 (N_647,N_584,N_580);
nor U648 (N_648,N_592,N_562);
and U649 (N_649,N_580,N_587);
and U650 (N_650,N_626,N_630);
nand U651 (N_651,N_647,N_612);
nand U652 (N_652,N_638,N_646);
and U653 (N_653,N_640,N_604);
or U654 (N_654,N_643,N_605);
nand U655 (N_655,N_642,N_618);
nand U656 (N_656,N_617,N_641);
nor U657 (N_657,N_609,N_615);
or U658 (N_658,N_623,N_625);
and U659 (N_659,N_619,N_634);
or U660 (N_660,N_644,N_635);
nor U661 (N_661,N_620,N_616);
nand U662 (N_662,N_628,N_622);
nor U663 (N_663,N_613,N_614);
nand U664 (N_664,N_649,N_645);
nand U665 (N_665,N_624,N_600);
and U666 (N_666,N_621,N_648);
and U667 (N_667,N_601,N_607);
nand U668 (N_668,N_611,N_629);
nor U669 (N_669,N_603,N_631);
nor U670 (N_670,N_633,N_627);
or U671 (N_671,N_608,N_610);
and U672 (N_672,N_636,N_632);
nand U673 (N_673,N_606,N_639);
or U674 (N_674,N_637,N_602);
nor U675 (N_675,N_646,N_625);
or U676 (N_676,N_624,N_609);
nand U677 (N_677,N_613,N_616);
and U678 (N_678,N_606,N_635);
or U679 (N_679,N_614,N_620);
nand U680 (N_680,N_606,N_645);
and U681 (N_681,N_632,N_635);
and U682 (N_682,N_611,N_644);
nor U683 (N_683,N_608,N_642);
and U684 (N_684,N_612,N_634);
or U685 (N_685,N_643,N_602);
nor U686 (N_686,N_639,N_641);
nand U687 (N_687,N_639,N_646);
nor U688 (N_688,N_622,N_605);
nand U689 (N_689,N_637,N_646);
or U690 (N_690,N_633,N_614);
nand U691 (N_691,N_628,N_637);
and U692 (N_692,N_613,N_611);
nor U693 (N_693,N_643,N_618);
nor U694 (N_694,N_639,N_603);
nor U695 (N_695,N_616,N_618);
or U696 (N_696,N_601,N_640);
nor U697 (N_697,N_641,N_615);
nor U698 (N_698,N_641,N_608);
nor U699 (N_699,N_606,N_641);
and U700 (N_700,N_652,N_659);
nor U701 (N_701,N_693,N_671);
nor U702 (N_702,N_670,N_686);
or U703 (N_703,N_657,N_667);
and U704 (N_704,N_684,N_675);
and U705 (N_705,N_651,N_685);
nor U706 (N_706,N_666,N_680);
nor U707 (N_707,N_689,N_672);
nor U708 (N_708,N_673,N_692);
and U709 (N_709,N_699,N_665);
or U710 (N_710,N_655,N_679);
nor U711 (N_711,N_677,N_688);
nor U712 (N_712,N_683,N_687);
and U713 (N_713,N_668,N_656);
nand U714 (N_714,N_682,N_678);
nor U715 (N_715,N_690,N_661);
nand U716 (N_716,N_662,N_658);
or U717 (N_717,N_650,N_676);
nor U718 (N_718,N_698,N_694);
and U719 (N_719,N_664,N_669);
or U720 (N_720,N_695,N_674);
nand U721 (N_721,N_663,N_660);
and U722 (N_722,N_697,N_696);
or U723 (N_723,N_681,N_654);
nor U724 (N_724,N_691,N_653);
and U725 (N_725,N_664,N_698);
xor U726 (N_726,N_696,N_699);
nor U727 (N_727,N_651,N_666);
xor U728 (N_728,N_698,N_667);
nand U729 (N_729,N_680,N_665);
nor U730 (N_730,N_692,N_691);
or U731 (N_731,N_657,N_651);
nand U732 (N_732,N_651,N_692);
and U733 (N_733,N_688,N_661);
nor U734 (N_734,N_665,N_682);
nand U735 (N_735,N_680,N_682);
nor U736 (N_736,N_688,N_682);
nand U737 (N_737,N_697,N_694);
nand U738 (N_738,N_677,N_652);
xor U739 (N_739,N_671,N_662);
or U740 (N_740,N_651,N_673);
and U741 (N_741,N_650,N_696);
and U742 (N_742,N_660,N_680);
and U743 (N_743,N_675,N_677);
nand U744 (N_744,N_684,N_674);
nor U745 (N_745,N_674,N_687);
and U746 (N_746,N_674,N_675);
and U747 (N_747,N_658,N_669);
or U748 (N_748,N_687,N_685);
nor U749 (N_749,N_673,N_661);
nand U750 (N_750,N_744,N_726);
nor U751 (N_751,N_716,N_745);
nand U752 (N_752,N_712,N_711);
nor U753 (N_753,N_708,N_701);
and U754 (N_754,N_718,N_709);
nor U755 (N_755,N_715,N_730);
nor U756 (N_756,N_714,N_732);
and U757 (N_757,N_742,N_734);
and U758 (N_758,N_738,N_748);
or U759 (N_759,N_707,N_749);
or U760 (N_760,N_741,N_729);
nor U761 (N_761,N_743,N_747);
nand U762 (N_762,N_733,N_725);
or U763 (N_763,N_704,N_737);
nor U764 (N_764,N_735,N_700);
nand U765 (N_765,N_721,N_723);
or U766 (N_766,N_719,N_702);
and U767 (N_767,N_731,N_710);
or U768 (N_768,N_713,N_746);
nand U769 (N_769,N_724,N_703);
nand U770 (N_770,N_717,N_736);
or U771 (N_771,N_720,N_705);
or U772 (N_772,N_706,N_727);
and U773 (N_773,N_728,N_739);
or U774 (N_774,N_740,N_722);
nand U775 (N_775,N_733,N_706);
nand U776 (N_776,N_715,N_736);
nor U777 (N_777,N_725,N_736);
or U778 (N_778,N_747,N_715);
nor U779 (N_779,N_718,N_732);
xnor U780 (N_780,N_733,N_726);
and U781 (N_781,N_706,N_730);
nor U782 (N_782,N_731,N_702);
xor U783 (N_783,N_705,N_746);
or U784 (N_784,N_744,N_705);
and U785 (N_785,N_729,N_718);
nand U786 (N_786,N_743,N_714);
or U787 (N_787,N_741,N_725);
or U788 (N_788,N_724,N_746);
or U789 (N_789,N_705,N_717);
and U790 (N_790,N_742,N_745);
and U791 (N_791,N_728,N_737);
and U792 (N_792,N_702,N_700);
and U793 (N_793,N_729,N_739);
and U794 (N_794,N_718,N_712);
nand U795 (N_795,N_703,N_719);
and U796 (N_796,N_720,N_726);
and U797 (N_797,N_721,N_717);
nor U798 (N_798,N_718,N_737);
or U799 (N_799,N_745,N_711);
or U800 (N_800,N_799,N_775);
or U801 (N_801,N_773,N_759);
nand U802 (N_802,N_753,N_798);
nand U803 (N_803,N_765,N_763);
nand U804 (N_804,N_796,N_752);
or U805 (N_805,N_779,N_787);
nor U806 (N_806,N_751,N_767);
nand U807 (N_807,N_795,N_760);
and U808 (N_808,N_781,N_776);
and U809 (N_809,N_770,N_755);
and U810 (N_810,N_778,N_792);
nand U811 (N_811,N_774,N_782);
and U812 (N_812,N_750,N_764);
nand U813 (N_813,N_754,N_786);
nor U814 (N_814,N_780,N_788);
and U815 (N_815,N_784,N_772);
or U816 (N_816,N_766,N_794);
or U817 (N_817,N_790,N_768);
nor U818 (N_818,N_793,N_771);
nor U819 (N_819,N_791,N_761);
or U820 (N_820,N_769,N_758);
nand U821 (N_821,N_756,N_789);
nor U822 (N_822,N_762,N_757);
nor U823 (N_823,N_783,N_797);
or U824 (N_824,N_785,N_777);
and U825 (N_825,N_762,N_753);
nand U826 (N_826,N_772,N_767);
nor U827 (N_827,N_754,N_766);
and U828 (N_828,N_782,N_797);
xnor U829 (N_829,N_774,N_756);
and U830 (N_830,N_776,N_765);
nor U831 (N_831,N_755,N_795);
or U832 (N_832,N_785,N_772);
and U833 (N_833,N_789,N_784);
nand U834 (N_834,N_778,N_752);
nand U835 (N_835,N_759,N_782);
nor U836 (N_836,N_795,N_787);
nor U837 (N_837,N_777,N_763);
nand U838 (N_838,N_765,N_791);
nor U839 (N_839,N_792,N_789);
nor U840 (N_840,N_780,N_787);
or U841 (N_841,N_754,N_768);
nor U842 (N_842,N_761,N_775);
nand U843 (N_843,N_757,N_761);
nor U844 (N_844,N_799,N_783);
nand U845 (N_845,N_794,N_750);
nor U846 (N_846,N_753,N_772);
or U847 (N_847,N_759,N_751);
nand U848 (N_848,N_753,N_781);
nor U849 (N_849,N_754,N_787);
nand U850 (N_850,N_837,N_835);
nor U851 (N_851,N_825,N_810);
xnor U852 (N_852,N_829,N_840);
nand U853 (N_853,N_819,N_839);
nand U854 (N_854,N_817,N_812);
and U855 (N_855,N_830,N_806);
xor U856 (N_856,N_834,N_826);
nor U857 (N_857,N_816,N_821);
and U858 (N_858,N_805,N_804);
or U859 (N_859,N_843,N_844);
or U860 (N_860,N_849,N_841);
and U861 (N_861,N_809,N_824);
or U862 (N_862,N_831,N_800);
nor U863 (N_863,N_820,N_814);
nor U864 (N_864,N_842,N_813);
nand U865 (N_865,N_811,N_801);
and U866 (N_866,N_833,N_846);
nand U867 (N_867,N_823,N_827);
and U868 (N_868,N_828,N_818);
or U869 (N_869,N_807,N_815);
or U870 (N_870,N_803,N_832);
and U871 (N_871,N_848,N_847);
nor U872 (N_872,N_845,N_822);
and U873 (N_873,N_836,N_802);
nor U874 (N_874,N_838,N_808);
nor U875 (N_875,N_800,N_837);
or U876 (N_876,N_814,N_819);
and U877 (N_877,N_812,N_840);
and U878 (N_878,N_823,N_848);
nand U879 (N_879,N_836,N_845);
and U880 (N_880,N_844,N_813);
nor U881 (N_881,N_827,N_833);
or U882 (N_882,N_819,N_803);
or U883 (N_883,N_837,N_848);
nand U884 (N_884,N_825,N_844);
nor U885 (N_885,N_846,N_809);
nor U886 (N_886,N_841,N_806);
nor U887 (N_887,N_808,N_846);
or U888 (N_888,N_813,N_806);
xnor U889 (N_889,N_825,N_826);
nor U890 (N_890,N_839,N_829);
and U891 (N_891,N_813,N_839);
and U892 (N_892,N_821,N_844);
nor U893 (N_893,N_843,N_828);
nand U894 (N_894,N_837,N_826);
nor U895 (N_895,N_835,N_800);
nand U896 (N_896,N_806,N_843);
and U897 (N_897,N_806,N_833);
or U898 (N_898,N_815,N_832);
and U899 (N_899,N_815,N_844);
nand U900 (N_900,N_856,N_891);
and U901 (N_901,N_879,N_877);
nor U902 (N_902,N_889,N_855);
and U903 (N_903,N_887,N_899);
or U904 (N_904,N_866,N_860);
or U905 (N_905,N_884,N_870);
or U906 (N_906,N_890,N_864);
and U907 (N_907,N_896,N_859);
nand U908 (N_908,N_862,N_869);
and U909 (N_909,N_878,N_893);
and U910 (N_910,N_867,N_880);
or U911 (N_911,N_876,N_868);
and U912 (N_912,N_854,N_872);
nor U913 (N_913,N_886,N_881);
nand U914 (N_914,N_865,N_853);
nand U915 (N_915,N_858,N_883);
and U916 (N_916,N_898,N_851);
and U917 (N_917,N_897,N_871);
and U918 (N_918,N_892,N_895);
and U919 (N_919,N_885,N_874);
and U920 (N_920,N_888,N_875);
nor U921 (N_921,N_850,N_873);
and U922 (N_922,N_857,N_861);
nor U923 (N_923,N_863,N_852);
or U924 (N_924,N_882,N_894);
nand U925 (N_925,N_891,N_858);
nor U926 (N_926,N_856,N_858);
nor U927 (N_927,N_851,N_850);
nor U928 (N_928,N_889,N_893);
nand U929 (N_929,N_894,N_878);
or U930 (N_930,N_895,N_875);
nor U931 (N_931,N_859,N_889);
and U932 (N_932,N_879,N_862);
or U933 (N_933,N_884,N_862);
nand U934 (N_934,N_853,N_871);
nor U935 (N_935,N_851,N_860);
nor U936 (N_936,N_852,N_887);
or U937 (N_937,N_872,N_873);
nor U938 (N_938,N_894,N_851);
and U939 (N_939,N_852,N_858);
or U940 (N_940,N_867,N_875);
or U941 (N_941,N_892,N_874);
or U942 (N_942,N_850,N_877);
nor U943 (N_943,N_892,N_858);
or U944 (N_944,N_875,N_891);
nand U945 (N_945,N_853,N_858);
and U946 (N_946,N_865,N_871);
and U947 (N_947,N_890,N_894);
or U948 (N_948,N_876,N_889);
nand U949 (N_949,N_881,N_870);
or U950 (N_950,N_932,N_938);
and U951 (N_951,N_916,N_933);
nor U952 (N_952,N_923,N_934);
or U953 (N_953,N_905,N_919);
nand U954 (N_954,N_914,N_910);
or U955 (N_955,N_920,N_917);
nor U956 (N_956,N_939,N_931);
or U957 (N_957,N_915,N_900);
nand U958 (N_958,N_949,N_903);
nor U959 (N_959,N_922,N_921);
nor U960 (N_960,N_925,N_927);
or U961 (N_961,N_904,N_947);
nand U962 (N_962,N_906,N_946);
and U963 (N_963,N_945,N_918);
and U964 (N_964,N_937,N_948);
or U965 (N_965,N_940,N_928);
and U966 (N_966,N_929,N_936);
or U967 (N_967,N_941,N_930);
nor U968 (N_968,N_902,N_926);
or U969 (N_969,N_942,N_913);
nor U970 (N_970,N_909,N_907);
nand U971 (N_971,N_912,N_908);
or U972 (N_972,N_901,N_943);
nand U973 (N_973,N_924,N_911);
and U974 (N_974,N_944,N_935);
nand U975 (N_975,N_937,N_906);
nor U976 (N_976,N_910,N_920);
nor U977 (N_977,N_907,N_943);
and U978 (N_978,N_902,N_905);
and U979 (N_979,N_941,N_912);
or U980 (N_980,N_939,N_924);
nor U981 (N_981,N_910,N_944);
nor U982 (N_982,N_905,N_927);
nor U983 (N_983,N_929,N_949);
nand U984 (N_984,N_917,N_935);
nor U985 (N_985,N_906,N_901);
or U986 (N_986,N_944,N_938);
nand U987 (N_987,N_922,N_944);
nor U988 (N_988,N_910,N_931);
and U989 (N_989,N_907,N_935);
and U990 (N_990,N_937,N_927);
and U991 (N_991,N_901,N_922);
nor U992 (N_992,N_906,N_913);
and U993 (N_993,N_919,N_901);
nor U994 (N_994,N_903,N_908);
or U995 (N_995,N_929,N_922);
and U996 (N_996,N_900,N_947);
or U997 (N_997,N_917,N_918);
nand U998 (N_998,N_949,N_905);
nor U999 (N_999,N_915,N_919);
nand U1000 (N_1000,N_964,N_995);
or U1001 (N_1001,N_973,N_996);
nand U1002 (N_1002,N_988,N_959);
or U1003 (N_1003,N_972,N_967);
and U1004 (N_1004,N_986,N_977);
or U1005 (N_1005,N_966,N_963);
nor U1006 (N_1006,N_960,N_990);
nand U1007 (N_1007,N_979,N_950);
nor U1008 (N_1008,N_952,N_970);
or U1009 (N_1009,N_981,N_992);
nor U1010 (N_1010,N_951,N_971);
or U1011 (N_1011,N_974,N_989);
nand U1012 (N_1012,N_954,N_999);
and U1013 (N_1013,N_953,N_962);
nor U1014 (N_1014,N_968,N_998);
nand U1015 (N_1015,N_985,N_991);
and U1016 (N_1016,N_957,N_956);
or U1017 (N_1017,N_983,N_975);
nor U1018 (N_1018,N_994,N_978);
and U1019 (N_1019,N_955,N_987);
nor U1020 (N_1020,N_969,N_982);
nand U1021 (N_1021,N_961,N_980);
and U1022 (N_1022,N_993,N_997);
nand U1023 (N_1023,N_984,N_976);
or U1024 (N_1024,N_958,N_965);
or U1025 (N_1025,N_987,N_991);
nand U1026 (N_1026,N_964,N_952);
or U1027 (N_1027,N_958,N_991);
and U1028 (N_1028,N_970,N_961);
or U1029 (N_1029,N_988,N_955);
nand U1030 (N_1030,N_966,N_996);
nor U1031 (N_1031,N_955,N_998);
nand U1032 (N_1032,N_953,N_994);
and U1033 (N_1033,N_982,N_993);
and U1034 (N_1034,N_972,N_996);
nand U1035 (N_1035,N_982,N_980);
nor U1036 (N_1036,N_956,N_973);
or U1037 (N_1037,N_991,N_993);
nor U1038 (N_1038,N_975,N_978);
nand U1039 (N_1039,N_993,N_983);
nor U1040 (N_1040,N_996,N_967);
or U1041 (N_1041,N_991,N_957);
nor U1042 (N_1042,N_998,N_981);
nor U1043 (N_1043,N_956,N_992);
and U1044 (N_1044,N_992,N_973);
and U1045 (N_1045,N_986,N_995);
xnor U1046 (N_1046,N_977,N_983);
nor U1047 (N_1047,N_958,N_959);
nor U1048 (N_1048,N_950,N_995);
or U1049 (N_1049,N_983,N_955);
or U1050 (N_1050,N_1008,N_1018);
and U1051 (N_1051,N_1005,N_1004);
or U1052 (N_1052,N_1029,N_1033);
and U1053 (N_1053,N_1041,N_1028);
or U1054 (N_1054,N_1002,N_1020);
nor U1055 (N_1055,N_1044,N_1030);
and U1056 (N_1056,N_1023,N_1000);
and U1057 (N_1057,N_1034,N_1024);
and U1058 (N_1058,N_1043,N_1013);
nor U1059 (N_1059,N_1006,N_1015);
nor U1060 (N_1060,N_1039,N_1009);
nor U1061 (N_1061,N_1049,N_1027);
and U1062 (N_1062,N_1010,N_1037);
and U1063 (N_1063,N_1007,N_1021);
and U1064 (N_1064,N_1038,N_1011);
xor U1065 (N_1065,N_1040,N_1012);
or U1066 (N_1066,N_1047,N_1042);
or U1067 (N_1067,N_1025,N_1045);
nor U1068 (N_1068,N_1017,N_1046);
or U1069 (N_1069,N_1032,N_1019);
and U1070 (N_1070,N_1036,N_1035);
nand U1071 (N_1071,N_1022,N_1016);
or U1072 (N_1072,N_1048,N_1031);
nand U1073 (N_1073,N_1003,N_1001);
and U1074 (N_1074,N_1014,N_1026);
or U1075 (N_1075,N_1002,N_1027);
nand U1076 (N_1076,N_1023,N_1006);
nand U1077 (N_1077,N_1036,N_1027);
nand U1078 (N_1078,N_1033,N_1008);
and U1079 (N_1079,N_1015,N_1041);
nand U1080 (N_1080,N_1006,N_1017);
and U1081 (N_1081,N_1028,N_1019);
nor U1082 (N_1082,N_1029,N_1014);
nand U1083 (N_1083,N_1002,N_1046);
or U1084 (N_1084,N_1003,N_1014);
nand U1085 (N_1085,N_1008,N_1036);
nor U1086 (N_1086,N_1028,N_1036);
or U1087 (N_1087,N_1032,N_1038);
and U1088 (N_1088,N_1007,N_1044);
and U1089 (N_1089,N_1022,N_1036);
and U1090 (N_1090,N_1046,N_1032);
and U1091 (N_1091,N_1023,N_1041);
nand U1092 (N_1092,N_1006,N_1018);
or U1093 (N_1093,N_1015,N_1020);
and U1094 (N_1094,N_1034,N_1013);
and U1095 (N_1095,N_1020,N_1036);
nand U1096 (N_1096,N_1026,N_1049);
nor U1097 (N_1097,N_1024,N_1015);
and U1098 (N_1098,N_1023,N_1020);
nor U1099 (N_1099,N_1006,N_1036);
and U1100 (N_1100,N_1099,N_1052);
and U1101 (N_1101,N_1081,N_1056);
nand U1102 (N_1102,N_1095,N_1083);
nand U1103 (N_1103,N_1067,N_1086);
or U1104 (N_1104,N_1058,N_1054);
nand U1105 (N_1105,N_1088,N_1094);
nand U1106 (N_1106,N_1070,N_1055);
or U1107 (N_1107,N_1065,N_1061);
nor U1108 (N_1108,N_1073,N_1078);
or U1109 (N_1109,N_1077,N_1069);
and U1110 (N_1110,N_1071,N_1090);
and U1111 (N_1111,N_1074,N_1084);
or U1112 (N_1112,N_1089,N_1050);
nand U1113 (N_1113,N_1064,N_1092);
or U1114 (N_1114,N_1066,N_1087);
or U1115 (N_1115,N_1082,N_1057);
and U1116 (N_1116,N_1075,N_1093);
nor U1117 (N_1117,N_1059,N_1076);
nand U1118 (N_1118,N_1085,N_1080);
xnor U1119 (N_1119,N_1079,N_1098);
nor U1120 (N_1120,N_1063,N_1072);
nor U1121 (N_1121,N_1091,N_1051);
nand U1122 (N_1122,N_1097,N_1068);
and U1123 (N_1123,N_1062,N_1096);
or U1124 (N_1124,N_1053,N_1060);
nor U1125 (N_1125,N_1055,N_1074);
nor U1126 (N_1126,N_1096,N_1085);
nor U1127 (N_1127,N_1053,N_1064);
nand U1128 (N_1128,N_1080,N_1064);
or U1129 (N_1129,N_1072,N_1098);
or U1130 (N_1130,N_1062,N_1090);
and U1131 (N_1131,N_1070,N_1093);
or U1132 (N_1132,N_1065,N_1082);
or U1133 (N_1133,N_1094,N_1096);
and U1134 (N_1134,N_1093,N_1090);
or U1135 (N_1135,N_1094,N_1050);
or U1136 (N_1136,N_1092,N_1056);
nand U1137 (N_1137,N_1067,N_1081);
and U1138 (N_1138,N_1093,N_1057);
and U1139 (N_1139,N_1070,N_1051);
and U1140 (N_1140,N_1095,N_1067);
and U1141 (N_1141,N_1089,N_1056);
and U1142 (N_1142,N_1095,N_1080);
nand U1143 (N_1143,N_1089,N_1077);
nor U1144 (N_1144,N_1062,N_1094);
nor U1145 (N_1145,N_1072,N_1094);
and U1146 (N_1146,N_1065,N_1088);
or U1147 (N_1147,N_1081,N_1057);
xnor U1148 (N_1148,N_1052,N_1089);
nor U1149 (N_1149,N_1096,N_1081);
or U1150 (N_1150,N_1104,N_1109);
or U1151 (N_1151,N_1119,N_1130);
nand U1152 (N_1152,N_1149,N_1123);
nand U1153 (N_1153,N_1103,N_1105);
and U1154 (N_1154,N_1125,N_1143);
or U1155 (N_1155,N_1137,N_1121);
or U1156 (N_1156,N_1114,N_1136);
or U1157 (N_1157,N_1146,N_1138);
and U1158 (N_1158,N_1145,N_1101);
nor U1159 (N_1159,N_1129,N_1118);
and U1160 (N_1160,N_1100,N_1113);
and U1161 (N_1161,N_1107,N_1124);
or U1162 (N_1162,N_1134,N_1127);
nor U1163 (N_1163,N_1128,N_1142);
or U1164 (N_1164,N_1139,N_1120);
and U1165 (N_1165,N_1106,N_1147);
nand U1166 (N_1166,N_1133,N_1140);
or U1167 (N_1167,N_1135,N_1112);
and U1168 (N_1168,N_1144,N_1131);
nand U1169 (N_1169,N_1115,N_1117);
or U1170 (N_1170,N_1122,N_1126);
and U1171 (N_1171,N_1148,N_1110);
nand U1172 (N_1172,N_1132,N_1108);
nand U1173 (N_1173,N_1111,N_1102);
nand U1174 (N_1174,N_1116,N_1141);
nand U1175 (N_1175,N_1114,N_1127);
nand U1176 (N_1176,N_1113,N_1127);
nor U1177 (N_1177,N_1105,N_1107);
nand U1178 (N_1178,N_1123,N_1111);
nor U1179 (N_1179,N_1120,N_1104);
nand U1180 (N_1180,N_1127,N_1128);
or U1181 (N_1181,N_1101,N_1121);
and U1182 (N_1182,N_1136,N_1127);
nor U1183 (N_1183,N_1107,N_1104);
xor U1184 (N_1184,N_1146,N_1109);
nor U1185 (N_1185,N_1102,N_1112);
or U1186 (N_1186,N_1125,N_1142);
nor U1187 (N_1187,N_1129,N_1115);
and U1188 (N_1188,N_1124,N_1100);
nand U1189 (N_1189,N_1134,N_1111);
nor U1190 (N_1190,N_1127,N_1146);
nand U1191 (N_1191,N_1149,N_1114);
nor U1192 (N_1192,N_1132,N_1145);
and U1193 (N_1193,N_1104,N_1135);
nor U1194 (N_1194,N_1114,N_1143);
nor U1195 (N_1195,N_1141,N_1144);
xnor U1196 (N_1196,N_1136,N_1105);
or U1197 (N_1197,N_1113,N_1149);
and U1198 (N_1198,N_1135,N_1102);
nand U1199 (N_1199,N_1143,N_1116);
nor U1200 (N_1200,N_1189,N_1185);
nor U1201 (N_1201,N_1175,N_1178);
or U1202 (N_1202,N_1157,N_1198);
or U1203 (N_1203,N_1168,N_1176);
nand U1204 (N_1204,N_1164,N_1195);
and U1205 (N_1205,N_1151,N_1154);
nand U1206 (N_1206,N_1187,N_1167);
nand U1207 (N_1207,N_1180,N_1199);
nand U1208 (N_1208,N_1159,N_1153);
and U1209 (N_1209,N_1194,N_1161);
or U1210 (N_1210,N_1155,N_1182);
nand U1211 (N_1211,N_1173,N_1170);
nor U1212 (N_1212,N_1162,N_1196);
or U1213 (N_1213,N_1184,N_1158);
nand U1214 (N_1214,N_1188,N_1183);
and U1215 (N_1215,N_1165,N_1152);
and U1216 (N_1216,N_1174,N_1190);
or U1217 (N_1217,N_1191,N_1169);
nor U1218 (N_1218,N_1193,N_1177);
nor U1219 (N_1219,N_1150,N_1186);
nor U1220 (N_1220,N_1160,N_1192);
and U1221 (N_1221,N_1197,N_1163);
nor U1222 (N_1222,N_1171,N_1179);
or U1223 (N_1223,N_1166,N_1181);
nand U1224 (N_1224,N_1172,N_1156);
and U1225 (N_1225,N_1168,N_1172);
nand U1226 (N_1226,N_1174,N_1184);
nor U1227 (N_1227,N_1177,N_1156);
and U1228 (N_1228,N_1192,N_1159);
and U1229 (N_1229,N_1174,N_1188);
nand U1230 (N_1230,N_1161,N_1181);
nor U1231 (N_1231,N_1163,N_1176);
and U1232 (N_1232,N_1173,N_1187);
nand U1233 (N_1233,N_1190,N_1177);
nand U1234 (N_1234,N_1164,N_1150);
and U1235 (N_1235,N_1158,N_1164);
or U1236 (N_1236,N_1165,N_1170);
nand U1237 (N_1237,N_1177,N_1162);
nor U1238 (N_1238,N_1190,N_1158);
nand U1239 (N_1239,N_1160,N_1174);
nand U1240 (N_1240,N_1185,N_1184);
nand U1241 (N_1241,N_1188,N_1175);
and U1242 (N_1242,N_1164,N_1159);
or U1243 (N_1243,N_1155,N_1199);
nor U1244 (N_1244,N_1152,N_1192);
nor U1245 (N_1245,N_1180,N_1160);
or U1246 (N_1246,N_1158,N_1159);
nand U1247 (N_1247,N_1197,N_1164);
or U1248 (N_1248,N_1150,N_1160);
and U1249 (N_1249,N_1167,N_1177);
or U1250 (N_1250,N_1246,N_1211);
nand U1251 (N_1251,N_1223,N_1216);
or U1252 (N_1252,N_1248,N_1210);
nor U1253 (N_1253,N_1225,N_1217);
and U1254 (N_1254,N_1224,N_1236);
and U1255 (N_1255,N_1233,N_1240);
nor U1256 (N_1256,N_1242,N_1237);
nor U1257 (N_1257,N_1208,N_1232);
nor U1258 (N_1258,N_1228,N_1230);
nor U1259 (N_1259,N_1243,N_1226);
or U1260 (N_1260,N_1241,N_1203);
or U1261 (N_1261,N_1201,N_1204);
nor U1262 (N_1262,N_1213,N_1235);
nor U1263 (N_1263,N_1244,N_1207);
and U1264 (N_1264,N_1221,N_1200);
nor U1265 (N_1265,N_1220,N_1218);
nand U1266 (N_1266,N_1234,N_1249);
or U1267 (N_1267,N_1209,N_1229);
xnor U1268 (N_1268,N_1222,N_1247);
nand U1269 (N_1269,N_1227,N_1245);
or U1270 (N_1270,N_1231,N_1212);
xor U1271 (N_1271,N_1219,N_1206);
nand U1272 (N_1272,N_1239,N_1202);
and U1273 (N_1273,N_1214,N_1215);
nor U1274 (N_1274,N_1238,N_1205);
or U1275 (N_1275,N_1231,N_1217);
or U1276 (N_1276,N_1231,N_1245);
and U1277 (N_1277,N_1220,N_1221);
or U1278 (N_1278,N_1228,N_1232);
nor U1279 (N_1279,N_1231,N_1218);
or U1280 (N_1280,N_1235,N_1239);
nor U1281 (N_1281,N_1231,N_1228);
or U1282 (N_1282,N_1219,N_1248);
nand U1283 (N_1283,N_1247,N_1209);
nor U1284 (N_1284,N_1231,N_1203);
and U1285 (N_1285,N_1247,N_1238);
nand U1286 (N_1286,N_1203,N_1208);
and U1287 (N_1287,N_1208,N_1202);
and U1288 (N_1288,N_1221,N_1235);
nor U1289 (N_1289,N_1233,N_1203);
nand U1290 (N_1290,N_1246,N_1205);
and U1291 (N_1291,N_1208,N_1234);
or U1292 (N_1292,N_1230,N_1222);
nand U1293 (N_1293,N_1226,N_1211);
and U1294 (N_1294,N_1229,N_1237);
nor U1295 (N_1295,N_1206,N_1215);
or U1296 (N_1296,N_1221,N_1247);
xor U1297 (N_1297,N_1244,N_1218);
and U1298 (N_1298,N_1240,N_1225);
nand U1299 (N_1299,N_1222,N_1229);
xnor U1300 (N_1300,N_1294,N_1278);
or U1301 (N_1301,N_1258,N_1299);
nand U1302 (N_1302,N_1256,N_1271);
or U1303 (N_1303,N_1270,N_1250);
nand U1304 (N_1304,N_1267,N_1260);
nor U1305 (N_1305,N_1287,N_1289);
and U1306 (N_1306,N_1286,N_1295);
nand U1307 (N_1307,N_1251,N_1254);
or U1308 (N_1308,N_1264,N_1263);
nor U1309 (N_1309,N_1297,N_1280);
or U1310 (N_1310,N_1293,N_1272);
nor U1311 (N_1311,N_1290,N_1291);
and U1312 (N_1312,N_1262,N_1284);
or U1313 (N_1313,N_1255,N_1259);
nand U1314 (N_1314,N_1282,N_1274);
nor U1315 (N_1315,N_1253,N_1268);
and U1316 (N_1316,N_1285,N_1292);
nor U1317 (N_1317,N_1281,N_1252);
nor U1318 (N_1318,N_1275,N_1265);
or U1319 (N_1319,N_1298,N_1296);
or U1320 (N_1320,N_1288,N_1273);
nand U1321 (N_1321,N_1276,N_1266);
or U1322 (N_1322,N_1279,N_1283);
or U1323 (N_1323,N_1257,N_1269);
and U1324 (N_1324,N_1261,N_1277);
nand U1325 (N_1325,N_1295,N_1257);
and U1326 (N_1326,N_1286,N_1273);
nor U1327 (N_1327,N_1296,N_1255);
nor U1328 (N_1328,N_1267,N_1287);
and U1329 (N_1329,N_1260,N_1262);
or U1330 (N_1330,N_1257,N_1281);
nor U1331 (N_1331,N_1299,N_1251);
nor U1332 (N_1332,N_1268,N_1270);
or U1333 (N_1333,N_1265,N_1293);
or U1334 (N_1334,N_1275,N_1292);
xor U1335 (N_1335,N_1257,N_1251);
nor U1336 (N_1336,N_1291,N_1292);
and U1337 (N_1337,N_1298,N_1286);
nand U1338 (N_1338,N_1271,N_1262);
nand U1339 (N_1339,N_1256,N_1297);
nand U1340 (N_1340,N_1283,N_1280);
nand U1341 (N_1341,N_1279,N_1270);
or U1342 (N_1342,N_1276,N_1263);
and U1343 (N_1343,N_1275,N_1272);
nand U1344 (N_1344,N_1293,N_1254);
nand U1345 (N_1345,N_1285,N_1250);
and U1346 (N_1346,N_1260,N_1286);
nor U1347 (N_1347,N_1251,N_1279);
and U1348 (N_1348,N_1288,N_1299);
nor U1349 (N_1349,N_1250,N_1256);
nand U1350 (N_1350,N_1301,N_1328);
nand U1351 (N_1351,N_1343,N_1300);
and U1352 (N_1352,N_1308,N_1338);
or U1353 (N_1353,N_1335,N_1320);
nor U1354 (N_1354,N_1345,N_1329);
or U1355 (N_1355,N_1323,N_1324);
nor U1356 (N_1356,N_1342,N_1302);
or U1357 (N_1357,N_1314,N_1304);
and U1358 (N_1358,N_1318,N_1307);
nand U1359 (N_1359,N_1319,N_1341);
nor U1360 (N_1360,N_1330,N_1325);
or U1361 (N_1361,N_1305,N_1336);
or U1362 (N_1362,N_1348,N_1316);
and U1363 (N_1363,N_1306,N_1327);
and U1364 (N_1364,N_1347,N_1346);
or U1365 (N_1365,N_1334,N_1333);
or U1366 (N_1366,N_1313,N_1311);
and U1367 (N_1367,N_1315,N_1322);
and U1368 (N_1368,N_1332,N_1310);
or U1369 (N_1369,N_1326,N_1317);
nor U1370 (N_1370,N_1349,N_1331);
or U1371 (N_1371,N_1309,N_1321);
nor U1372 (N_1372,N_1337,N_1312);
and U1373 (N_1373,N_1339,N_1344);
nand U1374 (N_1374,N_1340,N_1303);
nand U1375 (N_1375,N_1301,N_1326);
and U1376 (N_1376,N_1328,N_1348);
nand U1377 (N_1377,N_1303,N_1332);
nor U1378 (N_1378,N_1306,N_1313);
nand U1379 (N_1379,N_1320,N_1334);
nand U1380 (N_1380,N_1307,N_1336);
or U1381 (N_1381,N_1317,N_1348);
and U1382 (N_1382,N_1339,N_1348);
nand U1383 (N_1383,N_1341,N_1309);
or U1384 (N_1384,N_1333,N_1347);
or U1385 (N_1385,N_1323,N_1311);
and U1386 (N_1386,N_1344,N_1313);
or U1387 (N_1387,N_1338,N_1310);
or U1388 (N_1388,N_1319,N_1315);
nand U1389 (N_1389,N_1327,N_1315);
or U1390 (N_1390,N_1316,N_1311);
or U1391 (N_1391,N_1317,N_1336);
or U1392 (N_1392,N_1334,N_1310);
nor U1393 (N_1393,N_1335,N_1301);
nand U1394 (N_1394,N_1317,N_1323);
nand U1395 (N_1395,N_1325,N_1341);
and U1396 (N_1396,N_1310,N_1322);
or U1397 (N_1397,N_1332,N_1325);
nand U1398 (N_1398,N_1338,N_1326);
and U1399 (N_1399,N_1309,N_1303);
xnor U1400 (N_1400,N_1357,N_1389);
and U1401 (N_1401,N_1395,N_1358);
or U1402 (N_1402,N_1356,N_1370);
nand U1403 (N_1403,N_1386,N_1388);
and U1404 (N_1404,N_1379,N_1368);
or U1405 (N_1405,N_1363,N_1393);
or U1406 (N_1406,N_1355,N_1352);
and U1407 (N_1407,N_1387,N_1366);
nor U1408 (N_1408,N_1372,N_1375);
and U1409 (N_1409,N_1382,N_1380);
nand U1410 (N_1410,N_1364,N_1381);
nor U1411 (N_1411,N_1353,N_1396);
nor U1412 (N_1412,N_1394,N_1354);
nand U1413 (N_1413,N_1374,N_1359);
nor U1414 (N_1414,N_1371,N_1383);
or U1415 (N_1415,N_1385,N_1392);
nand U1416 (N_1416,N_1367,N_1377);
nor U1417 (N_1417,N_1373,N_1378);
nor U1418 (N_1418,N_1362,N_1398);
nor U1419 (N_1419,N_1384,N_1390);
nor U1420 (N_1420,N_1399,N_1391);
or U1421 (N_1421,N_1350,N_1351);
nor U1422 (N_1422,N_1397,N_1365);
nand U1423 (N_1423,N_1369,N_1361);
xor U1424 (N_1424,N_1376,N_1360);
and U1425 (N_1425,N_1390,N_1359);
and U1426 (N_1426,N_1365,N_1370);
and U1427 (N_1427,N_1358,N_1394);
or U1428 (N_1428,N_1379,N_1369);
nand U1429 (N_1429,N_1394,N_1376);
nor U1430 (N_1430,N_1351,N_1394);
and U1431 (N_1431,N_1361,N_1358);
nand U1432 (N_1432,N_1377,N_1354);
or U1433 (N_1433,N_1399,N_1362);
and U1434 (N_1434,N_1364,N_1372);
nor U1435 (N_1435,N_1383,N_1378);
nor U1436 (N_1436,N_1388,N_1350);
nand U1437 (N_1437,N_1356,N_1352);
and U1438 (N_1438,N_1386,N_1382);
nor U1439 (N_1439,N_1378,N_1350);
or U1440 (N_1440,N_1387,N_1395);
nor U1441 (N_1441,N_1374,N_1382);
nor U1442 (N_1442,N_1357,N_1367);
or U1443 (N_1443,N_1354,N_1352);
nor U1444 (N_1444,N_1367,N_1362);
nand U1445 (N_1445,N_1392,N_1388);
nand U1446 (N_1446,N_1392,N_1355);
nand U1447 (N_1447,N_1381,N_1389);
nand U1448 (N_1448,N_1383,N_1381);
and U1449 (N_1449,N_1377,N_1394);
nor U1450 (N_1450,N_1418,N_1427);
or U1451 (N_1451,N_1422,N_1432);
nand U1452 (N_1452,N_1406,N_1412);
nor U1453 (N_1453,N_1434,N_1413);
or U1454 (N_1454,N_1435,N_1438);
or U1455 (N_1455,N_1416,N_1400);
or U1456 (N_1456,N_1409,N_1403);
nand U1457 (N_1457,N_1404,N_1402);
nand U1458 (N_1458,N_1401,N_1430);
or U1459 (N_1459,N_1440,N_1419);
and U1460 (N_1460,N_1442,N_1429);
and U1461 (N_1461,N_1444,N_1407);
nand U1462 (N_1462,N_1443,N_1447);
nor U1463 (N_1463,N_1431,N_1421);
nand U1464 (N_1464,N_1446,N_1428);
and U1465 (N_1465,N_1437,N_1414);
nor U1466 (N_1466,N_1449,N_1436);
and U1467 (N_1467,N_1410,N_1408);
nor U1468 (N_1468,N_1433,N_1439);
or U1469 (N_1469,N_1423,N_1417);
nand U1470 (N_1470,N_1426,N_1441);
and U1471 (N_1471,N_1448,N_1420);
and U1472 (N_1472,N_1415,N_1424);
or U1473 (N_1473,N_1411,N_1445);
nor U1474 (N_1474,N_1405,N_1425);
or U1475 (N_1475,N_1443,N_1402);
nand U1476 (N_1476,N_1412,N_1422);
nor U1477 (N_1477,N_1449,N_1437);
and U1478 (N_1478,N_1416,N_1440);
nand U1479 (N_1479,N_1401,N_1403);
nor U1480 (N_1480,N_1423,N_1411);
and U1481 (N_1481,N_1436,N_1419);
nor U1482 (N_1482,N_1419,N_1404);
nor U1483 (N_1483,N_1433,N_1417);
nand U1484 (N_1484,N_1401,N_1405);
and U1485 (N_1485,N_1432,N_1429);
nor U1486 (N_1486,N_1411,N_1415);
or U1487 (N_1487,N_1407,N_1411);
and U1488 (N_1488,N_1425,N_1443);
or U1489 (N_1489,N_1413,N_1421);
nor U1490 (N_1490,N_1404,N_1401);
or U1491 (N_1491,N_1445,N_1412);
and U1492 (N_1492,N_1433,N_1432);
nand U1493 (N_1493,N_1430,N_1404);
nor U1494 (N_1494,N_1433,N_1411);
and U1495 (N_1495,N_1418,N_1422);
nand U1496 (N_1496,N_1420,N_1440);
or U1497 (N_1497,N_1448,N_1402);
and U1498 (N_1498,N_1449,N_1426);
nor U1499 (N_1499,N_1447,N_1439);
nor U1500 (N_1500,N_1454,N_1476);
nand U1501 (N_1501,N_1485,N_1477);
or U1502 (N_1502,N_1462,N_1481);
or U1503 (N_1503,N_1465,N_1457);
xnor U1504 (N_1504,N_1464,N_1480);
or U1505 (N_1505,N_1483,N_1488);
and U1506 (N_1506,N_1470,N_1498);
or U1507 (N_1507,N_1452,N_1463);
nor U1508 (N_1508,N_1479,N_1455);
nor U1509 (N_1509,N_1490,N_1499);
or U1510 (N_1510,N_1466,N_1475);
or U1511 (N_1511,N_1494,N_1461);
nor U1512 (N_1512,N_1493,N_1468);
nand U1513 (N_1513,N_1487,N_1458);
nand U1514 (N_1514,N_1486,N_1467);
nor U1515 (N_1515,N_1456,N_1472);
or U1516 (N_1516,N_1474,N_1453);
nand U1517 (N_1517,N_1471,N_1478);
and U1518 (N_1518,N_1473,N_1459);
nand U1519 (N_1519,N_1450,N_1469);
nand U1520 (N_1520,N_1482,N_1495);
nand U1521 (N_1521,N_1484,N_1491);
nor U1522 (N_1522,N_1496,N_1492);
or U1523 (N_1523,N_1489,N_1497);
or U1524 (N_1524,N_1451,N_1460);
nand U1525 (N_1525,N_1498,N_1490);
xor U1526 (N_1526,N_1460,N_1494);
nor U1527 (N_1527,N_1469,N_1485);
and U1528 (N_1528,N_1454,N_1461);
or U1529 (N_1529,N_1455,N_1466);
or U1530 (N_1530,N_1487,N_1466);
or U1531 (N_1531,N_1452,N_1451);
nand U1532 (N_1532,N_1477,N_1494);
or U1533 (N_1533,N_1499,N_1460);
nand U1534 (N_1534,N_1484,N_1450);
or U1535 (N_1535,N_1470,N_1488);
nand U1536 (N_1536,N_1477,N_1493);
nand U1537 (N_1537,N_1481,N_1465);
or U1538 (N_1538,N_1474,N_1466);
and U1539 (N_1539,N_1492,N_1481);
and U1540 (N_1540,N_1451,N_1494);
nor U1541 (N_1541,N_1492,N_1488);
and U1542 (N_1542,N_1489,N_1487);
nor U1543 (N_1543,N_1486,N_1466);
or U1544 (N_1544,N_1464,N_1460);
or U1545 (N_1545,N_1474,N_1497);
nand U1546 (N_1546,N_1492,N_1477);
nand U1547 (N_1547,N_1458,N_1456);
nand U1548 (N_1548,N_1481,N_1480);
nor U1549 (N_1549,N_1498,N_1467);
and U1550 (N_1550,N_1543,N_1537);
nand U1551 (N_1551,N_1545,N_1546);
nor U1552 (N_1552,N_1538,N_1523);
nor U1553 (N_1553,N_1506,N_1549);
and U1554 (N_1554,N_1547,N_1524);
and U1555 (N_1555,N_1528,N_1520);
nand U1556 (N_1556,N_1534,N_1525);
nand U1557 (N_1557,N_1516,N_1517);
and U1558 (N_1558,N_1542,N_1504);
nand U1559 (N_1559,N_1539,N_1527);
nand U1560 (N_1560,N_1502,N_1521);
nand U1561 (N_1561,N_1501,N_1540);
nand U1562 (N_1562,N_1515,N_1532);
nand U1563 (N_1563,N_1518,N_1512);
nor U1564 (N_1564,N_1541,N_1513);
or U1565 (N_1565,N_1507,N_1533);
nor U1566 (N_1566,N_1500,N_1505);
or U1567 (N_1567,N_1510,N_1548);
and U1568 (N_1568,N_1536,N_1526);
nor U1569 (N_1569,N_1535,N_1511);
nor U1570 (N_1570,N_1508,N_1514);
nor U1571 (N_1571,N_1531,N_1522);
or U1572 (N_1572,N_1503,N_1529);
nand U1573 (N_1573,N_1530,N_1509);
or U1574 (N_1574,N_1544,N_1519);
or U1575 (N_1575,N_1540,N_1505);
and U1576 (N_1576,N_1545,N_1540);
nor U1577 (N_1577,N_1538,N_1521);
and U1578 (N_1578,N_1513,N_1547);
nor U1579 (N_1579,N_1546,N_1540);
and U1580 (N_1580,N_1548,N_1526);
nand U1581 (N_1581,N_1516,N_1547);
or U1582 (N_1582,N_1504,N_1526);
or U1583 (N_1583,N_1527,N_1519);
nor U1584 (N_1584,N_1501,N_1526);
and U1585 (N_1585,N_1503,N_1536);
and U1586 (N_1586,N_1548,N_1533);
nand U1587 (N_1587,N_1526,N_1520);
nand U1588 (N_1588,N_1524,N_1538);
nand U1589 (N_1589,N_1531,N_1512);
or U1590 (N_1590,N_1535,N_1531);
nor U1591 (N_1591,N_1503,N_1523);
and U1592 (N_1592,N_1510,N_1508);
or U1593 (N_1593,N_1505,N_1542);
or U1594 (N_1594,N_1547,N_1521);
or U1595 (N_1595,N_1508,N_1512);
nor U1596 (N_1596,N_1510,N_1534);
nand U1597 (N_1597,N_1545,N_1503);
or U1598 (N_1598,N_1543,N_1534);
nor U1599 (N_1599,N_1542,N_1508);
or U1600 (N_1600,N_1561,N_1565);
or U1601 (N_1601,N_1574,N_1595);
nand U1602 (N_1602,N_1553,N_1564);
or U1603 (N_1603,N_1550,N_1569);
and U1604 (N_1604,N_1552,N_1576);
or U1605 (N_1605,N_1556,N_1585);
nor U1606 (N_1606,N_1579,N_1596);
and U1607 (N_1607,N_1597,N_1586);
nor U1608 (N_1608,N_1591,N_1583);
xnor U1609 (N_1609,N_1566,N_1582);
nand U1610 (N_1610,N_1568,N_1567);
or U1611 (N_1611,N_1577,N_1571);
nor U1612 (N_1612,N_1589,N_1578);
and U1613 (N_1613,N_1584,N_1555);
nand U1614 (N_1614,N_1598,N_1588);
xor U1615 (N_1615,N_1594,N_1581);
nand U1616 (N_1616,N_1554,N_1560);
xor U1617 (N_1617,N_1593,N_1563);
nor U1618 (N_1618,N_1599,N_1572);
nor U1619 (N_1619,N_1559,N_1558);
or U1620 (N_1620,N_1557,N_1551);
and U1621 (N_1621,N_1587,N_1562);
or U1622 (N_1622,N_1580,N_1570);
or U1623 (N_1623,N_1573,N_1592);
and U1624 (N_1624,N_1575,N_1590);
and U1625 (N_1625,N_1596,N_1552);
or U1626 (N_1626,N_1573,N_1550);
nand U1627 (N_1627,N_1580,N_1577);
or U1628 (N_1628,N_1574,N_1594);
nand U1629 (N_1629,N_1583,N_1568);
nor U1630 (N_1630,N_1585,N_1576);
nor U1631 (N_1631,N_1597,N_1582);
and U1632 (N_1632,N_1557,N_1597);
nand U1633 (N_1633,N_1560,N_1580);
or U1634 (N_1634,N_1576,N_1588);
and U1635 (N_1635,N_1556,N_1588);
or U1636 (N_1636,N_1592,N_1554);
nand U1637 (N_1637,N_1563,N_1575);
and U1638 (N_1638,N_1557,N_1586);
or U1639 (N_1639,N_1551,N_1568);
or U1640 (N_1640,N_1574,N_1588);
and U1641 (N_1641,N_1560,N_1559);
nand U1642 (N_1642,N_1565,N_1596);
nor U1643 (N_1643,N_1574,N_1561);
or U1644 (N_1644,N_1590,N_1576);
nand U1645 (N_1645,N_1599,N_1597);
nand U1646 (N_1646,N_1599,N_1568);
nand U1647 (N_1647,N_1574,N_1585);
and U1648 (N_1648,N_1592,N_1565);
nor U1649 (N_1649,N_1555,N_1553);
nand U1650 (N_1650,N_1639,N_1604);
or U1651 (N_1651,N_1641,N_1612);
or U1652 (N_1652,N_1611,N_1618);
nand U1653 (N_1653,N_1628,N_1608);
and U1654 (N_1654,N_1636,N_1624);
nor U1655 (N_1655,N_1647,N_1643);
nand U1656 (N_1656,N_1600,N_1642);
nand U1657 (N_1657,N_1638,N_1619);
nand U1658 (N_1658,N_1626,N_1615);
nor U1659 (N_1659,N_1606,N_1622);
nand U1660 (N_1660,N_1610,N_1634);
nand U1661 (N_1661,N_1614,N_1603);
or U1662 (N_1662,N_1602,N_1630);
nand U1663 (N_1663,N_1635,N_1648);
or U1664 (N_1664,N_1640,N_1637);
nand U1665 (N_1665,N_1623,N_1616);
and U1666 (N_1666,N_1617,N_1605);
and U1667 (N_1667,N_1607,N_1625);
or U1668 (N_1668,N_1609,N_1631);
or U1669 (N_1669,N_1629,N_1633);
nor U1670 (N_1670,N_1649,N_1646);
and U1671 (N_1671,N_1644,N_1645);
nand U1672 (N_1672,N_1601,N_1632);
and U1673 (N_1673,N_1621,N_1620);
and U1674 (N_1674,N_1627,N_1613);
nor U1675 (N_1675,N_1602,N_1606);
nor U1676 (N_1676,N_1619,N_1635);
nand U1677 (N_1677,N_1610,N_1611);
or U1678 (N_1678,N_1649,N_1622);
or U1679 (N_1679,N_1626,N_1632);
nand U1680 (N_1680,N_1612,N_1622);
or U1681 (N_1681,N_1622,N_1613);
or U1682 (N_1682,N_1602,N_1604);
or U1683 (N_1683,N_1626,N_1631);
and U1684 (N_1684,N_1602,N_1642);
or U1685 (N_1685,N_1640,N_1645);
and U1686 (N_1686,N_1628,N_1630);
or U1687 (N_1687,N_1624,N_1617);
nand U1688 (N_1688,N_1613,N_1600);
nor U1689 (N_1689,N_1648,N_1619);
or U1690 (N_1690,N_1646,N_1622);
or U1691 (N_1691,N_1603,N_1639);
and U1692 (N_1692,N_1605,N_1613);
and U1693 (N_1693,N_1648,N_1623);
nand U1694 (N_1694,N_1616,N_1612);
nand U1695 (N_1695,N_1609,N_1610);
nand U1696 (N_1696,N_1613,N_1649);
nor U1697 (N_1697,N_1631,N_1616);
and U1698 (N_1698,N_1604,N_1614);
nor U1699 (N_1699,N_1616,N_1635);
nand U1700 (N_1700,N_1677,N_1683);
and U1701 (N_1701,N_1684,N_1676);
and U1702 (N_1702,N_1697,N_1681);
nand U1703 (N_1703,N_1680,N_1658);
nand U1704 (N_1704,N_1664,N_1674);
or U1705 (N_1705,N_1659,N_1661);
or U1706 (N_1706,N_1670,N_1671);
or U1707 (N_1707,N_1653,N_1679);
nor U1708 (N_1708,N_1689,N_1690);
or U1709 (N_1709,N_1694,N_1687);
nor U1710 (N_1710,N_1652,N_1654);
nand U1711 (N_1711,N_1665,N_1666);
nor U1712 (N_1712,N_1685,N_1650);
or U1713 (N_1713,N_1660,N_1693);
nor U1714 (N_1714,N_1663,N_1657);
and U1715 (N_1715,N_1662,N_1651);
or U1716 (N_1716,N_1669,N_1667);
nor U1717 (N_1717,N_1695,N_1691);
and U1718 (N_1718,N_1688,N_1692);
nand U1719 (N_1719,N_1699,N_1675);
nor U1720 (N_1720,N_1672,N_1678);
nand U1721 (N_1721,N_1655,N_1668);
or U1722 (N_1722,N_1682,N_1698);
and U1723 (N_1723,N_1696,N_1686);
or U1724 (N_1724,N_1656,N_1673);
or U1725 (N_1725,N_1676,N_1657);
and U1726 (N_1726,N_1696,N_1679);
or U1727 (N_1727,N_1695,N_1674);
nor U1728 (N_1728,N_1662,N_1670);
nand U1729 (N_1729,N_1651,N_1653);
and U1730 (N_1730,N_1682,N_1694);
and U1731 (N_1731,N_1680,N_1687);
and U1732 (N_1732,N_1653,N_1656);
and U1733 (N_1733,N_1695,N_1690);
or U1734 (N_1734,N_1675,N_1687);
or U1735 (N_1735,N_1655,N_1684);
and U1736 (N_1736,N_1672,N_1650);
or U1737 (N_1737,N_1658,N_1674);
or U1738 (N_1738,N_1675,N_1667);
nor U1739 (N_1739,N_1653,N_1681);
nor U1740 (N_1740,N_1694,N_1658);
nand U1741 (N_1741,N_1676,N_1672);
nand U1742 (N_1742,N_1691,N_1674);
and U1743 (N_1743,N_1694,N_1699);
nor U1744 (N_1744,N_1689,N_1669);
nor U1745 (N_1745,N_1682,N_1651);
or U1746 (N_1746,N_1665,N_1685);
or U1747 (N_1747,N_1650,N_1686);
and U1748 (N_1748,N_1653,N_1696);
and U1749 (N_1749,N_1680,N_1695);
or U1750 (N_1750,N_1735,N_1724);
and U1751 (N_1751,N_1742,N_1725);
and U1752 (N_1752,N_1731,N_1711);
or U1753 (N_1753,N_1706,N_1743);
and U1754 (N_1754,N_1730,N_1729);
nor U1755 (N_1755,N_1716,N_1748);
and U1756 (N_1756,N_1736,N_1726);
or U1757 (N_1757,N_1728,N_1718);
and U1758 (N_1758,N_1715,N_1737);
or U1759 (N_1759,N_1712,N_1713);
nor U1760 (N_1760,N_1700,N_1727);
nand U1761 (N_1761,N_1705,N_1703);
or U1762 (N_1762,N_1704,N_1702);
nor U1763 (N_1763,N_1733,N_1749);
nor U1764 (N_1764,N_1722,N_1719);
and U1765 (N_1765,N_1744,N_1747);
nand U1766 (N_1766,N_1746,N_1709);
or U1767 (N_1767,N_1741,N_1714);
nand U1768 (N_1768,N_1721,N_1734);
or U1769 (N_1769,N_1732,N_1739);
or U1770 (N_1770,N_1701,N_1717);
and U1771 (N_1771,N_1740,N_1720);
xnor U1772 (N_1772,N_1723,N_1708);
or U1773 (N_1773,N_1707,N_1710);
nand U1774 (N_1774,N_1738,N_1745);
and U1775 (N_1775,N_1701,N_1719);
and U1776 (N_1776,N_1704,N_1735);
and U1777 (N_1777,N_1747,N_1715);
and U1778 (N_1778,N_1708,N_1714);
nor U1779 (N_1779,N_1743,N_1729);
nor U1780 (N_1780,N_1710,N_1733);
and U1781 (N_1781,N_1746,N_1723);
nor U1782 (N_1782,N_1713,N_1728);
and U1783 (N_1783,N_1703,N_1730);
nand U1784 (N_1784,N_1735,N_1740);
and U1785 (N_1785,N_1701,N_1743);
and U1786 (N_1786,N_1719,N_1732);
and U1787 (N_1787,N_1715,N_1702);
and U1788 (N_1788,N_1710,N_1749);
nand U1789 (N_1789,N_1725,N_1741);
and U1790 (N_1790,N_1709,N_1721);
and U1791 (N_1791,N_1744,N_1703);
or U1792 (N_1792,N_1721,N_1712);
or U1793 (N_1793,N_1712,N_1704);
nor U1794 (N_1794,N_1712,N_1729);
nand U1795 (N_1795,N_1709,N_1729);
or U1796 (N_1796,N_1749,N_1716);
or U1797 (N_1797,N_1720,N_1716);
and U1798 (N_1798,N_1717,N_1700);
and U1799 (N_1799,N_1727,N_1738);
or U1800 (N_1800,N_1787,N_1756);
or U1801 (N_1801,N_1770,N_1752);
or U1802 (N_1802,N_1786,N_1750);
nor U1803 (N_1803,N_1760,N_1791);
nand U1804 (N_1804,N_1755,N_1767);
and U1805 (N_1805,N_1769,N_1792);
and U1806 (N_1806,N_1796,N_1766);
nand U1807 (N_1807,N_1768,N_1795);
nand U1808 (N_1808,N_1778,N_1782);
nand U1809 (N_1809,N_1789,N_1771);
nand U1810 (N_1810,N_1757,N_1763);
nand U1811 (N_1811,N_1784,N_1777);
nand U1812 (N_1812,N_1762,N_1775);
nand U1813 (N_1813,N_1759,N_1776);
nand U1814 (N_1814,N_1785,N_1797);
and U1815 (N_1815,N_1798,N_1764);
or U1816 (N_1816,N_1793,N_1765);
nand U1817 (N_1817,N_1799,N_1758);
nor U1818 (N_1818,N_1753,N_1794);
or U1819 (N_1819,N_1772,N_1781);
nand U1820 (N_1820,N_1774,N_1751);
and U1821 (N_1821,N_1779,N_1754);
or U1822 (N_1822,N_1783,N_1790);
or U1823 (N_1823,N_1780,N_1761);
nor U1824 (N_1824,N_1773,N_1788);
nor U1825 (N_1825,N_1763,N_1791);
or U1826 (N_1826,N_1751,N_1755);
nor U1827 (N_1827,N_1774,N_1763);
and U1828 (N_1828,N_1786,N_1778);
nor U1829 (N_1829,N_1762,N_1752);
and U1830 (N_1830,N_1761,N_1763);
nand U1831 (N_1831,N_1769,N_1755);
nand U1832 (N_1832,N_1753,N_1755);
nor U1833 (N_1833,N_1782,N_1783);
or U1834 (N_1834,N_1792,N_1757);
nand U1835 (N_1835,N_1766,N_1751);
nand U1836 (N_1836,N_1791,N_1751);
or U1837 (N_1837,N_1761,N_1776);
and U1838 (N_1838,N_1750,N_1763);
nand U1839 (N_1839,N_1762,N_1768);
nand U1840 (N_1840,N_1791,N_1783);
nor U1841 (N_1841,N_1773,N_1755);
and U1842 (N_1842,N_1770,N_1795);
nand U1843 (N_1843,N_1756,N_1765);
xnor U1844 (N_1844,N_1768,N_1763);
and U1845 (N_1845,N_1771,N_1781);
and U1846 (N_1846,N_1796,N_1767);
and U1847 (N_1847,N_1765,N_1782);
nand U1848 (N_1848,N_1763,N_1786);
or U1849 (N_1849,N_1783,N_1758);
or U1850 (N_1850,N_1822,N_1832);
or U1851 (N_1851,N_1813,N_1804);
or U1852 (N_1852,N_1830,N_1844);
and U1853 (N_1853,N_1824,N_1826);
nand U1854 (N_1854,N_1840,N_1842);
nor U1855 (N_1855,N_1810,N_1808);
and U1856 (N_1856,N_1841,N_1819);
and U1857 (N_1857,N_1833,N_1828);
nand U1858 (N_1858,N_1848,N_1837);
nand U1859 (N_1859,N_1825,N_1821);
or U1860 (N_1860,N_1812,N_1849);
nand U1861 (N_1861,N_1820,N_1811);
and U1862 (N_1862,N_1802,N_1817);
or U1863 (N_1863,N_1827,N_1823);
nor U1864 (N_1864,N_1800,N_1839);
nand U1865 (N_1865,N_1807,N_1834);
xnor U1866 (N_1866,N_1809,N_1831);
nand U1867 (N_1867,N_1847,N_1814);
nand U1868 (N_1868,N_1846,N_1843);
or U1869 (N_1869,N_1806,N_1803);
or U1870 (N_1870,N_1805,N_1816);
nor U1871 (N_1871,N_1815,N_1836);
nor U1872 (N_1872,N_1801,N_1838);
or U1873 (N_1873,N_1835,N_1818);
nand U1874 (N_1874,N_1829,N_1845);
nand U1875 (N_1875,N_1831,N_1829);
nor U1876 (N_1876,N_1809,N_1818);
or U1877 (N_1877,N_1802,N_1827);
nor U1878 (N_1878,N_1830,N_1818);
nor U1879 (N_1879,N_1838,N_1832);
and U1880 (N_1880,N_1810,N_1804);
nor U1881 (N_1881,N_1806,N_1844);
nor U1882 (N_1882,N_1810,N_1844);
or U1883 (N_1883,N_1807,N_1828);
and U1884 (N_1884,N_1819,N_1830);
and U1885 (N_1885,N_1837,N_1820);
nor U1886 (N_1886,N_1840,N_1806);
or U1887 (N_1887,N_1848,N_1822);
nor U1888 (N_1888,N_1820,N_1801);
nand U1889 (N_1889,N_1847,N_1828);
or U1890 (N_1890,N_1820,N_1835);
nand U1891 (N_1891,N_1829,N_1847);
nor U1892 (N_1892,N_1822,N_1840);
nor U1893 (N_1893,N_1840,N_1807);
and U1894 (N_1894,N_1814,N_1827);
and U1895 (N_1895,N_1810,N_1823);
or U1896 (N_1896,N_1814,N_1845);
or U1897 (N_1897,N_1819,N_1834);
and U1898 (N_1898,N_1808,N_1823);
nand U1899 (N_1899,N_1807,N_1816);
nor U1900 (N_1900,N_1854,N_1889);
nand U1901 (N_1901,N_1861,N_1873);
and U1902 (N_1902,N_1859,N_1858);
nand U1903 (N_1903,N_1881,N_1894);
and U1904 (N_1904,N_1857,N_1877);
nand U1905 (N_1905,N_1874,N_1876);
and U1906 (N_1906,N_1864,N_1856);
nand U1907 (N_1907,N_1879,N_1896);
and U1908 (N_1908,N_1890,N_1892);
or U1909 (N_1909,N_1850,N_1887);
xor U1910 (N_1910,N_1872,N_1885);
and U1911 (N_1911,N_1868,N_1882);
nor U1912 (N_1912,N_1865,N_1897);
and U1913 (N_1913,N_1898,N_1862);
nor U1914 (N_1914,N_1895,N_1869);
and U1915 (N_1915,N_1888,N_1899);
and U1916 (N_1916,N_1866,N_1893);
nand U1917 (N_1917,N_1878,N_1851);
nor U1918 (N_1918,N_1886,N_1884);
or U1919 (N_1919,N_1883,N_1867);
or U1920 (N_1920,N_1855,N_1863);
and U1921 (N_1921,N_1875,N_1860);
nor U1922 (N_1922,N_1871,N_1870);
nor U1923 (N_1923,N_1880,N_1853);
nand U1924 (N_1924,N_1891,N_1852);
nand U1925 (N_1925,N_1856,N_1854);
nor U1926 (N_1926,N_1869,N_1860);
or U1927 (N_1927,N_1850,N_1884);
or U1928 (N_1928,N_1851,N_1868);
nand U1929 (N_1929,N_1882,N_1885);
nand U1930 (N_1930,N_1853,N_1887);
and U1931 (N_1931,N_1881,N_1859);
and U1932 (N_1932,N_1850,N_1874);
nor U1933 (N_1933,N_1850,N_1899);
nand U1934 (N_1934,N_1886,N_1882);
or U1935 (N_1935,N_1878,N_1887);
or U1936 (N_1936,N_1863,N_1857);
nor U1937 (N_1937,N_1862,N_1887);
nor U1938 (N_1938,N_1851,N_1893);
nand U1939 (N_1939,N_1871,N_1868);
or U1940 (N_1940,N_1860,N_1887);
nor U1941 (N_1941,N_1861,N_1887);
and U1942 (N_1942,N_1895,N_1864);
nand U1943 (N_1943,N_1859,N_1850);
nor U1944 (N_1944,N_1856,N_1874);
or U1945 (N_1945,N_1851,N_1862);
or U1946 (N_1946,N_1875,N_1881);
or U1947 (N_1947,N_1858,N_1893);
or U1948 (N_1948,N_1885,N_1854);
and U1949 (N_1949,N_1852,N_1855);
and U1950 (N_1950,N_1929,N_1919);
and U1951 (N_1951,N_1902,N_1917);
nor U1952 (N_1952,N_1912,N_1910);
and U1953 (N_1953,N_1949,N_1944);
nor U1954 (N_1954,N_1922,N_1911);
nor U1955 (N_1955,N_1939,N_1947);
or U1956 (N_1956,N_1930,N_1937);
nor U1957 (N_1957,N_1907,N_1936);
nor U1958 (N_1958,N_1928,N_1914);
and U1959 (N_1959,N_1945,N_1940);
nor U1960 (N_1960,N_1943,N_1942);
nor U1961 (N_1961,N_1904,N_1903);
and U1962 (N_1962,N_1941,N_1901);
nand U1963 (N_1963,N_1932,N_1918);
or U1964 (N_1964,N_1933,N_1905);
nor U1965 (N_1965,N_1935,N_1900);
and U1966 (N_1966,N_1946,N_1916);
or U1967 (N_1967,N_1906,N_1948);
or U1968 (N_1968,N_1908,N_1923);
xor U1969 (N_1969,N_1921,N_1931);
and U1970 (N_1970,N_1938,N_1915);
nor U1971 (N_1971,N_1913,N_1920);
nand U1972 (N_1972,N_1924,N_1909);
or U1973 (N_1973,N_1927,N_1934);
or U1974 (N_1974,N_1926,N_1925);
or U1975 (N_1975,N_1942,N_1941);
and U1976 (N_1976,N_1930,N_1917);
nor U1977 (N_1977,N_1917,N_1907);
and U1978 (N_1978,N_1902,N_1923);
and U1979 (N_1979,N_1944,N_1901);
xor U1980 (N_1980,N_1919,N_1914);
or U1981 (N_1981,N_1942,N_1913);
nand U1982 (N_1982,N_1916,N_1935);
nand U1983 (N_1983,N_1939,N_1929);
or U1984 (N_1984,N_1949,N_1904);
nor U1985 (N_1985,N_1909,N_1938);
nand U1986 (N_1986,N_1946,N_1921);
nand U1987 (N_1987,N_1913,N_1906);
and U1988 (N_1988,N_1901,N_1929);
or U1989 (N_1989,N_1923,N_1942);
nand U1990 (N_1990,N_1928,N_1902);
nor U1991 (N_1991,N_1908,N_1904);
nor U1992 (N_1992,N_1925,N_1915);
nor U1993 (N_1993,N_1910,N_1916);
nor U1994 (N_1994,N_1945,N_1909);
nor U1995 (N_1995,N_1917,N_1908);
nor U1996 (N_1996,N_1946,N_1944);
and U1997 (N_1997,N_1943,N_1926);
or U1998 (N_1998,N_1919,N_1908);
nor U1999 (N_1999,N_1925,N_1910);
and U2000 (N_2000,N_1972,N_1951);
nor U2001 (N_2001,N_1975,N_1977);
nor U2002 (N_2002,N_1996,N_1969);
nand U2003 (N_2003,N_1993,N_1981);
or U2004 (N_2004,N_1960,N_1999);
or U2005 (N_2005,N_1978,N_1998);
nor U2006 (N_2006,N_1959,N_1964);
nand U2007 (N_2007,N_1965,N_1955);
or U2008 (N_2008,N_1961,N_1962);
nor U2009 (N_2009,N_1992,N_1957);
and U2010 (N_2010,N_1987,N_1963);
and U2011 (N_2011,N_1994,N_1967);
and U2012 (N_2012,N_1988,N_1995);
or U2013 (N_2013,N_1953,N_1984);
nor U2014 (N_2014,N_1971,N_1986);
nand U2015 (N_2015,N_1983,N_1985);
nand U2016 (N_2016,N_1991,N_1950);
or U2017 (N_2017,N_1954,N_1952);
and U2018 (N_2018,N_1956,N_1958);
and U2019 (N_2019,N_1970,N_1982);
nor U2020 (N_2020,N_1980,N_1976);
or U2021 (N_2021,N_1973,N_1968);
nor U2022 (N_2022,N_1974,N_1989);
nand U2023 (N_2023,N_1966,N_1990);
nor U2024 (N_2024,N_1997,N_1979);
nor U2025 (N_2025,N_1952,N_1998);
nor U2026 (N_2026,N_1982,N_1961);
nand U2027 (N_2027,N_1987,N_1981);
or U2028 (N_2028,N_1956,N_1990);
and U2029 (N_2029,N_1992,N_1961);
nor U2030 (N_2030,N_1969,N_1979);
nand U2031 (N_2031,N_1994,N_1956);
nor U2032 (N_2032,N_1958,N_1955);
and U2033 (N_2033,N_1992,N_1987);
nor U2034 (N_2034,N_1978,N_1991);
nand U2035 (N_2035,N_1978,N_1970);
nand U2036 (N_2036,N_1968,N_1985);
xor U2037 (N_2037,N_1965,N_1976);
or U2038 (N_2038,N_1972,N_1970);
or U2039 (N_2039,N_1990,N_1957);
nor U2040 (N_2040,N_1997,N_1967);
or U2041 (N_2041,N_1980,N_1950);
or U2042 (N_2042,N_1960,N_1981);
or U2043 (N_2043,N_1960,N_1994);
nor U2044 (N_2044,N_1959,N_1957);
nand U2045 (N_2045,N_1960,N_1975);
nor U2046 (N_2046,N_1958,N_1971);
or U2047 (N_2047,N_1984,N_1969);
and U2048 (N_2048,N_1951,N_1982);
nor U2049 (N_2049,N_1992,N_1954);
and U2050 (N_2050,N_2010,N_2027);
nor U2051 (N_2051,N_2015,N_2008);
nand U2052 (N_2052,N_2040,N_2032);
and U2053 (N_2053,N_2000,N_2030);
and U2054 (N_2054,N_2014,N_2049);
nor U2055 (N_2055,N_2047,N_2005);
nand U2056 (N_2056,N_2013,N_2004);
nor U2057 (N_2057,N_2035,N_2011);
or U2058 (N_2058,N_2017,N_2006);
and U2059 (N_2059,N_2020,N_2016);
nand U2060 (N_2060,N_2048,N_2026);
and U2061 (N_2061,N_2002,N_2037);
and U2062 (N_2062,N_2012,N_2046);
or U2063 (N_2063,N_2034,N_2003);
nor U2064 (N_2064,N_2033,N_2038);
or U2065 (N_2065,N_2043,N_2019);
nor U2066 (N_2066,N_2018,N_2022);
and U2067 (N_2067,N_2009,N_2023);
or U2068 (N_2068,N_2041,N_2045);
and U2069 (N_2069,N_2036,N_2029);
nor U2070 (N_2070,N_2021,N_2025);
nand U2071 (N_2071,N_2024,N_2028);
nor U2072 (N_2072,N_2031,N_2007);
or U2073 (N_2073,N_2001,N_2044);
or U2074 (N_2074,N_2039,N_2042);
and U2075 (N_2075,N_2005,N_2040);
and U2076 (N_2076,N_2004,N_2008);
and U2077 (N_2077,N_2032,N_2016);
and U2078 (N_2078,N_2030,N_2002);
and U2079 (N_2079,N_2015,N_2012);
and U2080 (N_2080,N_2011,N_2023);
nand U2081 (N_2081,N_2025,N_2041);
and U2082 (N_2082,N_2025,N_2024);
nand U2083 (N_2083,N_2046,N_2024);
and U2084 (N_2084,N_2044,N_2035);
or U2085 (N_2085,N_2024,N_2006);
nand U2086 (N_2086,N_2035,N_2020);
xor U2087 (N_2087,N_2020,N_2045);
and U2088 (N_2088,N_2046,N_2026);
nand U2089 (N_2089,N_2048,N_2017);
nand U2090 (N_2090,N_2019,N_2008);
nor U2091 (N_2091,N_2010,N_2035);
nand U2092 (N_2092,N_2034,N_2000);
nand U2093 (N_2093,N_2023,N_2041);
nand U2094 (N_2094,N_2023,N_2046);
and U2095 (N_2095,N_2031,N_2011);
nand U2096 (N_2096,N_2007,N_2003);
or U2097 (N_2097,N_2001,N_2008);
or U2098 (N_2098,N_2033,N_2047);
and U2099 (N_2099,N_2013,N_2040);
nor U2100 (N_2100,N_2066,N_2059);
and U2101 (N_2101,N_2068,N_2095);
nand U2102 (N_2102,N_2064,N_2070);
nand U2103 (N_2103,N_2094,N_2053);
nand U2104 (N_2104,N_2075,N_2085);
nor U2105 (N_2105,N_2051,N_2081);
nor U2106 (N_2106,N_2074,N_2077);
nand U2107 (N_2107,N_2055,N_2080);
and U2108 (N_2108,N_2061,N_2054);
and U2109 (N_2109,N_2088,N_2097);
or U2110 (N_2110,N_2083,N_2057);
nand U2111 (N_2111,N_2087,N_2079);
and U2112 (N_2112,N_2096,N_2093);
or U2113 (N_2113,N_2082,N_2091);
or U2114 (N_2114,N_2086,N_2090);
or U2115 (N_2115,N_2052,N_2072);
nand U2116 (N_2116,N_2073,N_2065);
or U2117 (N_2117,N_2098,N_2050);
or U2118 (N_2118,N_2092,N_2067);
nor U2119 (N_2119,N_2078,N_2099);
and U2120 (N_2120,N_2071,N_2084);
nand U2121 (N_2121,N_2069,N_2076);
nand U2122 (N_2122,N_2063,N_2056);
nor U2123 (N_2123,N_2058,N_2062);
nor U2124 (N_2124,N_2089,N_2060);
or U2125 (N_2125,N_2060,N_2081);
and U2126 (N_2126,N_2082,N_2071);
or U2127 (N_2127,N_2051,N_2096);
nor U2128 (N_2128,N_2067,N_2083);
nand U2129 (N_2129,N_2084,N_2081);
nand U2130 (N_2130,N_2097,N_2071);
nor U2131 (N_2131,N_2093,N_2090);
and U2132 (N_2132,N_2051,N_2058);
nor U2133 (N_2133,N_2062,N_2089);
or U2134 (N_2134,N_2073,N_2078);
nor U2135 (N_2135,N_2062,N_2085);
nor U2136 (N_2136,N_2069,N_2099);
nand U2137 (N_2137,N_2091,N_2068);
or U2138 (N_2138,N_2069,N_2071);
nor U2139 (N_2139,N_2089,N_2079);
or U2140 (N_2140,N_2081,N_2092);
nand U2141 (N_2141,N_2050,N_2063);
nand U2142 (N_2142,N_2084,N_2089);
or U2143 (N_2143,N_2075,N_2067);
nand U2144 (N_2144,N_2080,N_2076);
or U2145 (N_2145,N_2066,N_2050);
nand U2146 (N_2146,N_2079,N_2078);
nor U2147 (N_2147,N_2099,N_2054);
nor U2148 (N_2148,N_2074,N_2054);
nor U2149 (N_2149,N_2053,N_2089);
nor U2150 (N_2150,N_2103,N_2121);
and U2151 (N_2151,N_2115,N_2111);
and U2152 (N_2152,N_2132,N_2146);
nor U2153 (N_2153,N_2117,N_2104);
nor U2154 (N_2154,N_2140,N_2102);
nor U2155 (N_2155,N_2137,N_2113);
or U2156 (N_2156,N_2141,N_2126);
and U2157 (N_2157,N_2129,N_2145);
nor U2158 (N_2158,N_2131,N_2101);
nand U2159 (N_2159,N_2127,N_2133);
nand U2160 (N_2160,N_2106,N_2139);
or U2161 (N_2161,N_2124,N_2144);
nand U2162 (N_2162,N_2149,N_2123);
nor U2163 (N_2163,N_2107,N_2120);
and U2164 (N_2164,N_2105,N_2134);
and U2165 (N_2165,N_2136,N_2119);
nor U2166 (N_2166,N_2142,N_2128);
nand U2167 (N_2167,N_2122,N_2148);
or U2168 (N_2168,N_2100,N_2108);
nand U2169 (N_2169,N_2147,N_2143);
or U2170 (N_2170,N_2109,N_2118);
nor U2171 (N_2171,N_2138,N_2110);
and U2172 (N_2172,N_2125,N_2112);
or U2173 (N_2173,N_2135,N_2114);
nand U2174 (N_2174,N_2116,N_2130);
and U2175 (N_2175,N_2100,N_2106);
or U2176 (N_2176,N_2129,N_2126);
and U2177 (N_2177,N_2101,N_2133);
nor U2178 (N_2178,N_2141,N_2109);
nor U2179 (N_2179,N_2120,N_2140);
nand U2180 (N_2180,N_2111,N_2147);
nand U2181 (N_2181,N_2139,N_2126);
or U2182 (N_2182,N_2105,N_2126);
nand U2183 (N_2183,N_2109,N_2115);
or U2184 (N_2184,N_2132,N_2115);
or U2185 (N_2185,N_2138,N_2147);
nand U2186 (N_2186,N_2113,N_2140);
and U2187 (N_2187,N_2123,N_2132);
or U2188 (N_2188,N_2106,N_2109);
nand U2189 (N_2189,N_2139,N_2117);
or U2190 (N_2190,N_2106,N_2113);
nor U2191 (N_2191,N_2116,N_2119);
and U2192 (N_2192,N_2116,N_2145);
nand U2193 (N_2193,N_2146,N_2130);
nand U2194 (N_2194,N_2126,N_2111);
nand U2195 (N_2195,N_2100,N_2132);
and U2196 (N_2196,N_2141,N_2146);
nand U2197 (N_2197,N_2137,N_2114);
nor U2198 (N_2198,N_2144,N_2115);
or U2199 (N_2199,N_2105,N_2115);
and U2200 (N_2200,N_2157,N_2186);
nor U2201 (N_2201,N_2154,N_2171);
or U2202 (N_2202,N_2175,N_2178);
nor U2203 (N_2203,N_2170,N_2165);
or U2204 (N_2204,N_2191,N_2176);
nand U2205 (N_2205,N_2156,N_2177);
nand U2206 (N_2206,N_2185,N_2174);
nand U2207 (N_2207,N_2166,N_2196);
nor U2208 (N_2208,N_2190,N_2195);
nand U2209 (N_2209,N_2188,N_2181);
nand U2210 (N_2210,N_2151,N_2180);
nand U2211 (N_2211,N_2162,N_2193);
or U2212 (N_2212,N_2158,N_2164);
nor U2213 (N_2213,N_2150,N_2155);
or U2214 (N_2214,N_2153,N_2167);
nor U2215 (N_2215,N_2192,N_2183);
or U2216 (N_2216,N_2159,N_2198);
or U2217 (N_2217,N_2194,N_2160);
or U2218 (N_2218,N_2189,N_2172);
and U2219 (N_2219,N_2197,N_2182);
or U2220 (N_2220,N_2169,N_2184);
nor U2221 (N_2221,N_2179,N_2168);
nand U2222 (N_2222,N_2199,N_2187);
or U2223 (N_2223,N_2163,N_2173);
nand U2224 (N_2224,N_2161,N_2152);
and U2225 (N_2225,N_2170,N_2157);
or U2226 (N_2226,N_2191,N_2184);
nand U2227 (N_2227,N_2161,N_2192);
and U2228 (N_2228,N_2166,N_2187);
or U2229 (N_2229,N_2172,N_2156);
nor U2230 (N_2230,N_2164,N_2174);
nor U2231 (N_2231,N_2173,N_2175);
nand U2232 (N_2232,N_2158,N_2179);
and U2233 (N_2233,N_2170,N_2193);
and U2234 (N_2234,N_2177,N_2176);
and U2235 (N_2235,N_2166,N_2170);
nor U2236 (N_2236,N_2164,N_2154);
nor U2237 (N_2237,N_2166,N_2181);
or U2238 (N_2238,N_2183,N_2176);
or U2239 (N_2239,N_2171,N_2159);
nand U2240 (N_2240,N_2160,N_2170);
or U2241 (N_2241,N_2153,N_2185);
or U2242 (N_2242,N_2194,N_2184);
nor U2243 (N_2243,N_2182,N_2188);
xor U2244 (N_2244,N_2186,N_2173);
nand U2245 (N_2245,N_2188,N_2190);
nand U2246 (N_2246,N_2199,N_2167);
nor U2247 (N_2247,N_2186,N_2160);
nor U2248 (N_2248,N_2181,N_2161);
or U2249 (N_2249,N_2177,N_2167);
nand U2250 (N_2250,N_2217,N_2220);
nor U2251 (N_2251,N_2247,N_2239);
or U2252 (N_2252,N_2212,N_2230);
and U2253 (N_2253,N_2238,N_2203);
and U2254 (N_2254,N_2222,N_2246);
nor U2255 (N_2255,N_2229,N_2202);
and U2256 (N_2256,N_2232,N_2245);
and U2257 (N_2257,N_2228,N_2216);
and U2258 (N_2258,N_2209,N_2201);
nor U2259 (N_2259,N_2249,N_2241);
nor U2260 (N_2260,N_2211,N_2208);
nand U2261 (N_2261,N_2200,N_2223);
and U2262 (N_2262,N_2206,N_2210);
nor U2263 (N_2263,N_2234,N_2226);
or U2264 (N_2264,N_2244,N_2243);
nor U2265 (N_2265,N_2231,N_2224);
and U2266 (N_2266,N_2205,N_2219);
nor U2267 (N_2267,N_2207,N_2214);
and U2268 (N_2268,N_2215,N_2237);
and U2269 (N_2269,N_2235,N_2221);
or U2270 (N_2270,N_2218,N_2236);
or U2271 (N_2271,N_2213,N_2204);
or U2272 (N_2272,N_2248,N_2225);
and U2273 (N_2273,N_2227,N_2242);
nand U2274 (N_2274,N_2233,N_2240);
nand U2275 (N_2275,N_2226,N_2203);
xor U2276 (N_2276,N_2230,N_2219);
and U2277 (N_2277,N_2204,N_2206);
nor U2278 (N_2278,N_2243,N_2238);
nor U2279 (N_2279,N_2200,N_2222);
or U2280 (N_2280,N_2236,N_2220);
nor U2281 (N_2281,N_2224,N_2215);
nor U2282 (N_2282,N_2206,N_2216);
and U2283 (N_2283,N_2240,N_2214);
nand U2284 (N_2284,N_2218,N_2219);
and U2285 (N_2285,N_2223,N_2245);
nand U2286 (N_2286,N_2200,N_2213);
xor U2287 (N_2287,N_2206,N_2223);
or U2288 (N_2288,N_2226,N_2225);
xnor U2289 (N_2289,N_2236,N_2240);
and U2290 (N_2290,N_2201,N_2202);
and U2291 (N_2291,N_2237,N_2223);
nand U2292 (N_2292,N_2223,N_2241);
nor U2293 (N_2293,N_2208,N_2216);
nor U2294 (N_2294,N_2238,N_2200);
or U2295 (N_2295,N_2248,N_2208);
and U2296 (N_2296,N_2206,N_2219);
nand U2297 (N_2297,N_2231,N_2227);
nor U2298 (N_2298,N_2249,N_2221);
or U2299 (N_2299,N_2215,N_2234);
or U2300 (N_2300,N_2288,N_2261);
nor U2301 (N_2301,N_2290,N_2268);
or U2302 (N_2302,N_2275,N_2278);
or U2303 (N_2303,N_2296,N_2283);
nor U2304 (N_2304,N_2291,N_2265);
nand U2305 (N_2305,N_2251,N_2273);
nor U2306 (N_2306,N_2298,N_2258);
and U2307 (N_2307,N_2297,N_2271);
and U2308 (N_2308,N_2257,N_2295);
or U2309 (N_2309,N_2293,N_2286);
or U2310 (N_2310,N_2266,N_2277);
or U2311 (N_2311,N_2299,N_2255);
and U2312 (N_2312,N_2254,N_2280);
nand U2313 (N_2313,N_2284,N_2282);
and U2314 (N_2314,N_2287,N_2272);
or U2315 (N_2315,N_2289,N_2264);
xor U2316 (N_2316,N_2294,N_2292);
or U2317 (N_2317,N_2269,N_2250);
and U2318 (N_2318,N_2285,N_2253);
nand U2319 (N_2319,N_2252,N_2281);
or U2320 (N_2320,N_2279,N_2259);
or U2321 (N_2321,N_2274,N_2262);
nor U2322 (N_2322,N_2260,N_2270);
nand U2323 (N_2323,N_2256,N_2267);
nor U2324 (N_2324,N_2276,N_2263);
or U2325 (N_2325,N_2251,N_2286);
nor U2326 (N_2326,N_2270,N_2293);
nor U2327 (N_2327,N_2282,N_2293);
and U2328 (N_2328,N_2281,N_2263);
or U2329 (N_2329,N_2278,N_2260);
or U2330 (N_2330,N_2251,N_2285);
and U2331 (N_2331,N_2264,N_2267);
xnor U2332 (N_2332,N_2260,N_2263);
and U2333 (N_2333,N_2293,N_2276);
or U2334 (N_2334,N_2293,N_2257);
nand U2335 (N_2335,N_2263,N_2261);
and U2336 (N_2336,N_2285,N_2257);
and U2337 (N_2337,N_2274,N_2282);
and U2338 (N_2338,N_2293,N_2252);
and U2339 (N_2339,N_2292,N_2279);
or U2340 (N_2340,N_2271,N_2263);
nand U2341 (N_2341,N_2269,N_2257);
and U2342 (N_2342,N_2277,N_2259);
nand U2343 (N_2343,N_2276,N_2270);
or U2344 (N_2344,N_2292,N_2297);
nand U2345 (N_2345,N_2295,N_2293);
nand U2346 (N_2346,N_2292,N_2272);
nand U2347 (N_2347,N_2287,N_2280);
nand U2348 (N_2348,N_2264,N_2270);
nand U2349 (N_2349,N_2273,N_2257);
xor U2350 (N_2350,N_2347,N_2323);
nand U2351 (N_2351,N_2340,N_2313);
and U2352 (N_2352,N_2309,N_2322);
nand U2353 (N_2353,N_2319,N_2348);
nand U2354 (N_2354,N_2317,N_2332);
or U2355 (N_2355,N_2331,N_2304);
or U2356 (N_2356,N_2330,N_2302);
or U2357 (N_2357,N_2315,N_2301);
or U2358 (N_2358,N_2329,N_2349);
or U2359 (N_2359,N_2310,N_2316);
or U2360 (N_2360,N_2321,N_2325);
or U2361 (N_2361,N_2311,N_2314);
nor U2362 (N_2362,N_2333,N_2318);
or U2363 (N_2363,N_2324,N_2305);
nor U2364 (N_2364,N_2339,N_2320);
nand U2365 (N_2365,N_2338,N_2327);
nand U2366 (N_2366,N_2342,N_2344);
or U2367 (N_2367,N_2300,N_2335);
nand U2368 (N_2368,N_2308,N_2326);
and U2369 (N_2369,N_2307,N_2341);
and U2370 (N_2370,N_2345,N_2306);
and U2371 (N_2371,N_2343,N_2328);
nor U2372 (N_2372,N_2303,N_2334);
nand U2373 (N_2373,N_2337,N_2336);
nor U2374 (N_2374,N_2346,N_2312);
nand U2375 (N_2375,N_2307,N_2346);
and U2376 (N_2376,N_2339,N_2328);
and U2377 (N_2377,N_2346,N_2343);
nand U2378 (N_2378,N_2317,N_2304);
and U2379 (N_2379,N_2308,N_2309);
or U2380 (N_2380,N_2317,N_2331);
or U2381 (N_2381,N_2329,N_2339);
or U2382 (N_2382,N_2319,N_2335);
or U2383 (N_2383,N_2303,N_2310);
or U2384 (N_2384,N_2308,N_2314);
nand U2385 (N_2385,N_2331,N_2329);
nor U2386 (N_2386,N_2317,N_2347);
nand U2387 (N_2387,N_2332,N_2337);
and U2388 (N_2388,N_2326,N_2333);
and U2389 (N_2389,N_2310,N_2330);
nor U2390 (N_2390,N_2327,N_2303);
nand U2391 (N_2391,N_2349,N_2301);
or U2392 (N_2392,N_2324,N_2331);
nand U2393 (N_2393,N_2309,N_2348);
or U2394 (N_2394,N_2311,N_2331);
and U2395 (N_2395,N_2302,N_2309);
nand U2396 (N_2396,N_2331,N_2328);
nand U2397 (N_2397,N_2346,N_2310);
or U2398 (N_2398,N_2324,N_2329);
nand U2399 (N_2399,N_2345,N_2318);
nand U2400 (N_2400,N_2392,N_2389);
nand U2401 (N_2401,N_2393,N_2372);
and U2402 (N_2402,N_2357,N_2364);
nor U2403 (N_2403,N_2368,N_2378);
or U2404 (N_2404,N_2377,N_2380);
nor U2405 (N_2405,N_2369,N_2366);
and U2406 (N_2406,N_2353,N_2397);
and U2407 (N_2407,N_2386,N_2398);
or U2408 (N_2408,N_2354,N_2387);
nand U2409 (N_2409,N_2356,N_2388);
nor U2410 (N_2410,N_2355,N_2374);
nor U2411 (N_2411,N_2395,N_2376);
nor U2412 (N_2412,N_2351,N_2370);
and U2413 (N_2413,N_2399,N_2382);
nand U2414 (N_2414,N_2358,N_2383);
or U2415 (N_2415,N_2394,N_2381);
and U2416 (N_2416,N_2363,N_2371);
nor U2417 (N_2417,N_2375,N_2384);
nor U2418 (N_2418,N_2367,N_2360);
and U2419 (N_2419,N_2359,N_2361);
nor U2420 (N_2420,N_2390,N_2373);
nand U2421 (N_2421,N_2365,N_2362);
nor U2422 (N_2422,N_2391,N_2396);
or U2423 (N_2423,N_2350,N_2379);
nand U2424 (N_2424,N_2352,N_2385);
nor U2425 (N_2425,N_2375,N_2362);
nor U2426 (N_2426,N_2370,N_2369);
and U2427 (N_2427,N_2393,N_2380);
or U2428 (N_2428,N_2360,N_2374);
nand U2429 (N_2429,N_2357,N_2385);
nand U2430 (N_2430,N_2381,N_2372);
or U2431 (N_2431,N_2353,N_2393);
nand U2432 (N_2432,N_2358,N_2376);
or U2433 (N_2433,N_2372,N_2383);
or U2434 (N_2434,N_2396,N_2357);
or U2435 (N_2435,N_2398,N_2397);
or U2436 (N_2436,N_2381,N_2398);
or U2437 (N_2437,N_2377,N_2351);
or U2438 (N_2438,N_2351,N_2388);
nand U2439 (N_2439,N_2365,N_2369);
or U2440 (N_2440,N_2398,N_2359);
nand U2441 (N_2441,N_2384,N_2380);
nor U2442 (N_2442,N_2399,N_2365);
and U2443 (N_2443,N_2391,N_2398);
nor U2444 (N_2444,N_2359,N_2386);
or U2445 (N_2445,N_2367,N_2397);
nor U2446 (N_2446,N_2387,N_2390);
and U2447 (N_2447,N_2371,N_2359);
nand U2448 (N_2448,N_2366,N_2378);
nor U2449 (N_2449,N_2372,N_2384);
and U2450 (N_2450,N_2445,N_2416);
nand U2451 (N_2451,N_2421,N_2443);
or U2452 (N_2452,N_2405,N_2420);
nand U2453 (N_2453,N_2404,N_2402);
or U2454 (N_2454,N_2424,N_2407);
or U2455 (N_2455,N_2446,N_2444);
nand U2456 (N_2456,N_2403,N_2406);
nor U2457 (N_2457,N_2410,N_2438);
nand U2458 (N_2458,N_2417,N_2440);
xor U2459 (N_2459,N_2447,N_2401);
and U2460 (N_2460,N_2429,N_2433);
nand U2461 (N_2461,N_2423,N_2430);
and U2462 (N_2462,N_2441,N_2400);
or U2463 (N_2463,N_2449,N_2442);
nand U2464 (N_2464,N_2411,N_2415);
or U2465 (N_2465,N_2419,N_2439);
and U2466 (N_2466,N_2409,N_2418);
and U2467 (N_2467,N_2426,N_2435);
nor U2468 (N_2468,N_2414,N_2408);
nand U2469 (N_2469,N_2434,N_2428);
or U2470 (N_2470,N_2422,N_2436);
xnor U2471 (N_2471,N_2432,N_2437);
and U2472 (N_2472,N_2413,N_2427);
nor U2473 (N_2473,N_2448,N_2425);
nand U2474 (N_2474,N_2431,N_2412);
nor U2475 (N_2475,N_2410,N_2439);
nor U2476 (N_2476,N_2415,N_2427);
nand U2477 (N_2477,N_2446,N_2418);
or U2478 (N_2478,N_2440,N_2408);
nor U2479 (N_2479,N_2414,N_2439);
and U2480 (N_2480,N_2408,N_2405);
nand U2481 (N_2481,N_2420,N_2430);
and U2482 (N_2482,N_2412,N_2421);
nand U2483 (N_2483,N_2430,N_2422);
and U2484 (N_2484,N_2443,N_2428);
nor U2485 (N_2485,N_2405,N_2434);
xnor U2486 (N_2486,N_2407,N_2405);
and U2487 (N_2487,N_2448,N_2419);
nor U2488 (N_2488,N_2428,N_2423);
and U2489 (N_2489,N_2412,N_2414);
or U2490 (N_2490,N_2404,N_2434);
or U2491 (N_2491,N_2428,N_2425);
nand U2492 (N_2492,N_2418,N_2438);
or U2493 (N_2493,N_2417,N_2419);
nand U2494 (N_2494,N_2400,N_2439);
and U2495 (N_2495,N_2448,N_2415);
or U2496 (N_2496,N_2433,N_2431);
or U2497 (N_2497,N_2430,N_2402);
or U2498 (N_2498,N_2413,N_2449);
and U2499 (N_2499,N_2437,N_2446);
and U2500 (N_2500,N_2455,N_2498);
nor U2501 (N_2501,N_2456,N_2491);
or U2502 (N_2502,N_2450,N_2475);
or U2503 (N_2503,N_2458,N_2473);
and U2504 (N_2504,N_2468,N_2485);
xnor U2505 (N_2505,N_2484,N_2452);
or U2506 (N_2506,N_2460,N_2487);
or U2507 (N_2507,N_2494,N_2495);
and U2508 (N_2508,N_2479,N_2478);
nand U2509 (N_2509,N_2492,N_2481);
or U2510 (N_2510,N_2477,N_2464);
or U2511 (N_2511,N_2471,N_2490);
and U2512 (N_2512,N_2457,N_2480);
nor U2513 (N_2513,N_2499,N_2472);
nand U2514 (N_2514,N_2459,N_2454);
and U2515 (N_2515,N_2451,N_2474);
or U2516 (N_2516,N_2470,N_2465);
nand U2517 (N_2517,N_2482,N_2488);
or U2518 (N_2518,N_2497,N_2467);
nand U2519 (N_2519,N_2486,N_2476);
nand U2520 (N_2520,N_2469,N_2462);
nand U2521 (N_2521,N_2461,N_2489);
nor U2522 (N_2522,N_2496,N_2483);
nor U2523 (N_2523,N_2463,N_2466);
or U2524 (N_2524,N_2453,N_2493);
nand U2525 (N_2525,N_2494,N_2457);
and U2526 (N_2526,N_2465,N_2484);
nand U2527 (N_2527,N_2478,N_2482);
and U2528 (N_2528,N_2469,N_2474);
nor U2529 (N_2529,N_2490,N_2480);
nor U2530 (N_2530,N_2495,N_2453);
or U2531 (N_2531,N_2462,N_2467);
or U2532 (N_2532,N_2466,N_2450);
or U2533 (N_2533,N_2455,N_2472);
and U2534 (N_2534,N_2498,N_2491);
nor U2535 (N_2535,N_2465,N_2455);
xor U2536 (N_2536,N_2493,N_2489);
or U2537 (N_2537,N_2469,N_2463);
and U2538 (N_2538,N_2496,N_2497);
nor U2539 (N_2539,N_2495,N_2499);
and U2540 (N_2540,N_2481,N_2491);
nand U2541 (N_2541,N_2456,N_2464);
or U2542 (N_2542,N_2471,N_2488);
and U2543 (N_2543,N_2462,N_2475);
nor U2544 (N_2544,N_2461,N_2468);
nor U2545 (N_2545,N_2472,N_2484);
nor U2546 (N_2546,N_2481,N_2472);
nor U2547 (N_2547,N_2477,N_2470);
nand U2548 (N_2548,N_2456,N_2457);
and U2549 (N_2549,N_2458,N_2468);
xnor U2550 (N_2550,N_2548,N_2509);
nor U2551 (N_2551,N_2510,N_2522);
or U2552 (N_2552,N_2526,N_2547);
nor U2553 (N_2553,N_2532,N_2516);
and U2554 (N_2554,N_2549,N_2542);
or U2555 (N_2555,N_2546,N_2541);
or U2556 (N_2556,N_2543,N_2540);
or U2557 (N_2557,N_2530,N_2511);
nand U2558 (N_2558,N_2518,N_2528);
nor U2559 (N_2559,N_2520,N_2504);
and U2560 (N_2560,N_2508,N_2535);
or U2561 (N_2561,N_2523,N_2527);
and U2562 (N_2562,N_2515,N_2531);
nor U2563 (N_2563,N_2539,N_2536);
nand U2564 (N_2564,N_2505,N_2545);
nand U2565 (N_2565,N_2529,N_2500);
and U2566 (N_2566,N_2503,N_2514);
or U2567 (N_2567,N_2521,N_2517);
nor U2568 (N_2568,N_2534,N_2513);
or U2569 (N_2569,N_2537,N_2507);
nand U2570 (N_2570,N_2533,N_2506);
or U2571 (N_2571,N_2524,N_2525);
and U2572 (N_2572,N_2512,N_2538);
or U2573 (N_2573,N_2544,N_2502);
and U2574 (N_2574,N_2501,N_2519);
or U2575 (N_2575,N_2524,N_2505);
or U2576 (N_2576,N_2536,N_2501);
or U2577 (N_2577,N_2504,N_2522);
and U2578 (N_2578,N_2533,N_2526);
or U2579 (N_2579,N_2516,N_2522);
or U2580 (N_2580,N_2530,N_2510);
and U2581 (N_2581,N_2548,N_2513);
or U2582 (N_2582,N_2501,N_2537);
or U2583 (N_2583,N_2545,N_2519);
or U2584 (N_2584,N_2521,N_2540);
nand U2585 (N_2585,N_2524,N_2539);
and U2586 (N_2586,N_2529,N_2516);
or U2587 (N_2587,N_2537,N_2545);
nor U2588 (N_2588,N_2519,N_2548);
and U2589 (N_2589,N_2526,N_2504);
nor U2590 (N_2590,N_2517,N_2528);
or U2591 (N_2591,N_2521,N_2504);
and U2592 (N_2592,N_2512,N_2540);
nor U2593 (N_2593,N_2510,N_2514);
nor U2594 (N_2594,N_2534,N_2541);
nor U2595 (N_2595,N_2527,N_2537);
nand U2596 (N_2596,N_2508,N_2530);
and U2597 (N_2597,N_2541,N_2531);
and U2598 (N_2598,N_2521,N_2509);
nand U2599 (N_2599,N_2506,N_2517);
nand U2600 (N_2600,N_2550,N_2583);
nor U2601 (N_2601,N_2558,N_2587);
and U2602 (N_2602,N_2575,N_2556);
nor U2603 (N_2603,N_2570,N_2596);
or U2604 (N_2604,N_2562,N_2573);
nor U2605 (N_2605,N_2590,N_2564);
nor U2606 (N_2606,N_2579,N_2574);
nand U2607 (N_2607,N_2593,N_2585);
nand U2608 (N_2608,N_2576,N_2595);
and U2609 (N_2609,N_2552,N_2559);
nand U2610 (N_2610,N_2572,N_2568);
nor U2611 (N_2611,N_2551,N_2599);
or U2612 (N_2612,N_2598,N_2577);
or U2613 (N_2613,N_2584,N_2569);
and U2614 (N_2614,N_2563,N_2571);
nand U2615 (N_2615,N_2594,N_2561);
nor U2616 (N_2616,N_2567,N_2586);
nor U2617 (N_2617,N_2578,N_2589);
nand U2618 (N_2618,N_2565,N_2555);
nor U2619 (N_2619,N_2588,N_2553);
or U2620 (N_2620,N_2581,N_2592);
nand U2621 (N_2621,N_2554,N_2582);
nor U2622 (N_2622,N_2597,N_2557);
nor U2623 (N_2623,N_2591,N_2580);
or U2624 (N_2624,N_2560,N_2566);
nor U2625 (N_2625,N_2561,N_2556);
nor U2626 (N_2626,N_2579,N_2569);
nand U2627 (N_2627,N_2597,N_2565);
and U2628 (N_2628,N_2575,N_2598);
nand U2629 (N_2629,N_2551,N_2576);
nor U2630 (N_2630,N_2551,N_2555);
and U2631 (N_2631,N_2588,N_2599);
or U2632 (N_2632,N_2554,N_2552);
and U2633 (N_2633,N_2587,N_2575);
nand U2634 (N_2634,N_2569,N_2563);
or U2635 (N_2635,N_2592,N_2578);
and U2636 (N_2636,N_2570,N_2577);
and U2637 (N_2637,N_2596,N_2550);
nand U2638 (N_2638,N_2559,N_2589);
nand U2639 (N_2639,N_2584,N_2580);
nor U2640 (N_2640,N_2586,N_2560);
nand U2641 (N_2641,N_2575,N_2594);
nor U2642 (N_2642,N_2590,N_2595);
nand U2643 (N_2643,N_2573,N_2579);
or U2644 (N_2644,N_2578,N_2570);
nand U2645 (N_2645,N_2593,N_2598);
and U2646 (N_2646,N_2588,N_2570);
and U2647 (N_2647,N_2552,N_2580);
nor U2648 (N_2648,N_2563,N_2579);
nor U2649 (N_2649,N_2566,N_2595);
and U2650 (N_2650,N_2614,N_2641);
nand U2651 (N_2651,N_2637,N_2608);
or U2652 (N_2652,N_2615,N_2618);
or U2653 (N_2653,N_2632,N_2627);
or U2654 (N_2654,N_2612,N_2626);
and U2655 (N_2655,N_2635,N_2619);
nand U2656 (N_2656,N_2605,N_2620);
nor U2657 (N_2657,N_2639,N_2631);
and U2658 (N_2658,N_2642,N_2617);
or U2659 (N_2659,N_2604,N_2611);
nand U2660 (N_2660,N_2616,N_2607);
nor U2661 (N_2661,N_2649,N_2602);
nor U2662 (N_2662,N_2623,N_2648);
nand U2663 (N_2663,N_2638,N_2646);
or U2664 (N_2664,N_2603,N_2600);
and U2665 (N_2665,N_2636,N_2609);
or U2666 (N_2666,N_2645,N_2622);
and U2667 (N_2667,N_2613,N_2628);
xor U2668 (N_2668,N_2624,N_2630);
nand U2669 (N_2669,N_2610,N_2644);
xor U2670 (N_2670,N_2647,N_2625);
nor U2671 (N_2671,N_2643,N_2606);
nor U2672 (N_2672,N_2633,N_2629);
nor U2673 (N_2673,N_2601,N_2634);
and U2674 (N_2674,N_2621,N_2640);
nand U2675 (N_2675,N_2630,N_2607);
nor U2676 (N_2676,N_2629,N_2627);
or U2677 (N_2677,N_2614,N_2642);
nor U2678 (N_2678,N_2634,N_2604);
nand U2679 (N_2679,N_2607,N_2637);
nor U2680 (N_2680,N_2606,N_2603);
or U2681 (N_2681,N_2600,N_2612);
or U2682 (N_2682,N_2636,N_2619);
nor U2683 (N_2683,N_2623,N_2606);
or U2684 (N_2684,N_2600,N_2643);
and U2685 (N_2685,N_2625,N_2636);
nor U2686 (N_2686,N_2631,N_2630);
nor U2687 (N_2687,N_2622,N_2629);
or U2688 (N_2688,N_2642,N_2603);
and U2689 (N_2689,N_2623,N_2626);
or U2690 (N_2690,N_2602,N_2604);
or U2691 (N_2691,N_2606,N_2637);
and U2692 (N_2692,N_2628,N_2623);
and U2693 (N_2693,N_2631,N_2628);
nor U2694 (N_2694,N_2602,N_2641);
nor U2695 (N_2695,N_2639,N_2635);
nand U2696 (N_2696,N_2604,N_2629);
or U2697 (N_2697,N_2628,N_2647);
nor U2698 (N_2698,N_2642,N_2637);
or U2699 (N_2699,N_2605,N_2614);
nand U2700 (N_2700,N_2675,N_2691);
or U2701 (N_2701,N_2694,N_2657);
nand U2702 (N_2702,N_2695,N_2692);
nand U2703 (N_2703,N_2658,N_2678);
nor U2704 (N_2704,N_2689,N_2697);
nor U2705 (N_2705,N_2685,N_2690);
nand U2706 (N_2706,N_2655,N_2687);
and U2707 (N_2707,N_2673,N_2669);
and U2708 (N_2708,N_2696,N_2653);
nand U2709 (N_2709,N_2656,N_2665);
nor U2710 (N_2710,N_2684,N_2671);
nor U2711 (N_2711,N_2662,N_2670);
nand U2712 (N_2712,N_2680,N_2698);
nor U2713 (N_2713,N_2672,N_2650);
nor U2714 (N_2714,N_2677,N_2674);
nor U2715 (N_2715,N_2682,N_2667);
nor U2716 (N_2716,N_2686,N_2663);
nand U2717 (N_2717,N_2652,N_2683);
or U2718 (N_2718,N_2666,N_2693);
nor U2719 (N_2719,N_2688,N_2654);
nor U2720 (N_2720,N_2668,N_2651);
nand U2721 (N_2721,N_2681,N_2659);
and U2722 (N_2722,N_2664,N_2660);
and U2723 (N_2723,N_2699,N_2661);
nor U2724 (N_2724,N_2676,N_2679);
and U2725 (N_2725,N_2657,N_2676);
nand U2726 (N_2726,N_2666,N_2670);
and U2727 (N_2727,N_2660,N_2683);
nor U2728 (N_2728,N_2687,N_2679);
nor U2729 (N_2729,N_2695,N_2665);
and U2730 (N_2730,N_2675,N_2658);
or U2731 (N_2731,N_2684,N_2699);
or U2732 (N_2732,N_2656,N_2688);
or U2733 (N_2733,N_2679,N_2650);
nand U2734 (N_2734,N_2661,N_2679);
or U2735 (N_2735,N_2658,N_2682);
nor U2736 (N_2736,N_2683,N_2672);
nand U2737 (N_2737,N_2697,N_2680);
and U2738 (N_2738,N_2677,N_2690);
and U2739 (N_2739,N_2670,N_2674);
nor U2740 (N_2740,N_2688,N_2673);
or U2741 (N_2741,N_2666,N_2650);
and U2742 (N_2742,N_2685,N_2679);
or U2743 (N_2743,N_2686,N_2658);
or U2744 (N_2744,N_2679,N_2696);
or U2745 (N_2745,N_2692,N_2676);
nand U2746 (N_2746,N_2698,N_2665);
or U2747 (N_2747,N_2680,N_2663);
and U2748 (N_2748,N_2689,N_2692);
or U2749 (N_2749,N_2692,N_2687);
nor U2750 (N_2750,N_2721,N_2714);
and U2751 (N_2751,N_2731,N_2707);
nand U2752 (N_2752,N_2738,N_2716);
and U2753 (N_2753,N_2701,N_2742);
nor U2754 (N_2754,N_2747,N_2718);
nor U2755 (N_2755,N_2746,N_2740);
nor U2756 (N_2756,N_2749,N_2744);
nand U2757 (N_2757,N_2709,N_2732);
and U2758 (N_2758,N_2727,N_2748);
nand U2759 (N_2759,N_2705,N_2723);
xnor U2760 (N_2760,N_2730,N_2708);
or U2761 (N_2761,N_2743,N_2722);
nand U2762 (N_2762,N_2713,N_2710);
nor U2763 (N_2763,N_2717,N_2733);
nand U2764 (N_2764,N_2703,N_2725);
nand U2765 (N_2765,N_2706,N_2715);
xor U2766 (N_2766,N_2729,N_2720);
nor U2767 (N_2767,N_2726,N_2736);
or U2768 (N_2768,N_2737,N_2739);
or U2769 (N_2769,N_2700,N_2711);
and U2770 (N_2770,N_2734,N_2735);
and U2771 (N_2771,N_2745,N_2724);
nand U2772 (N_2772,N_2719,N_2704);
nor U2773 (N_2773,N_2728,N_2741);
and U2774 (N_2774,N_2712,N_2702);
nor U2775 (N_2775,N_2718,N_2728);
nand U2776 (N_2776,N_2700,N_2749);
nor U2777 (N_2777,N_2742,N_2735);
or U2778 (N_2778,N_2724,N_2712);
or U2779 (N_2779,N_2744,N_2737);
nor U2780 (N_2780,N_2741,N_2743);
and U2781 (N_2781,N_2744,N_2729);
nor U2782 (N_2782,N_2716,N_2735);
and U2783 (N_2783,N_2705,N_2724);
or U2784 (N_2784,N_2733,N_2711);
nand U2785 (N_2785,N_2706,N_2730);
nand U2786 (N_2786,N_2712,N_2713);
or U2787 (N_2787,N_2713,N_2706);
nand U2788 (N_2788,N_2713,N_2701);
nor U2789 (N_2789,N_2728,N_2710);
nor U2790 (N_2790,N_2714,N_2749);
nand U2791 (N_2791,N_2707,N_2723);
nand U2792 (N_2792,N_2720,N_2735);
nand U2793 (N_2793,N_2737,N_2736);
nor U2794 (N_2794,N_2749,N_2742);
nor U2795 (N_2795,N_2713,N_2716);
nor U2796 (N_2796,N_2729,N_2735);
and U2797 (N_2797,N_2728,N_2730);
or U2798 (N_2798,N_2723,N_2725);
nand U2799 (N_2799,N_2720,N_2740);
nand U2800 (N_2800,N_2758,N_2787);
nand U2801 (N_2801,N_2785,N_2754);
nor U2802 (N_2802,N_2793,N_2789);
and U2803 (N_2803,N_2786,N_2788);
or U2804 (N_2804,N_2765,N_2784);
or U2805 (N_2805,N_2771,N_2796);
and U2806 (N_2806,N_2797,N_2782);
nor U2807 (N_2807,N_2775,N_2778);
nor U2808 (N_2808,N_2780,N_2772);
nor U2809 (N_2809,N_2774,N_2790);
nand U2810 (N_2810,N_2799,N_2798);
nor U2811 (N_2811,N_2794,N_2791);
nor U2812 (N_2812,N_2760,N_2763);
and U2813 (N_2813,N_2762,N_2770);
nand U2814 (N_2814,N_2768,N_2767);
nand U2815 (N_2815,N_2752,N_2766);
or U2816 (N_2816,N_2755,N_2759);
nand U2817 (N_2817,N_2753,N_2764);
nor U2818 (N_2818,N_2792,N_2769);
nand U2819 (N_2819,N_2761,N_2779);
or U2820 (N_2820,N_2756,N_2773);
nand U2821 (N_2821,N_2777,N_2757);
nor U2822 (N_2822,N_2783,N_2750);
or U2823 (N_2823,N_2776,N_2751);
or U2824 (N_2824,N_2795,N_2781);
and U2825 (N_2825,N_2798,N_2780);
nand U2826 (N_2826,N_2759,N_2767);
nand U2827 (N_2827,N_2757,N_2778);
or U2828 (N_2828,N_2798,N_2772);
or U2829 (N_2829,N_2781,N_2788);
and U2830 (N_2830,N_2799,N_2767);
nand U2831 (N_2831,N_2772,N_2786);
and U2832 (N_2832,N_2783,N_2796);
nand U2833 (N_2833,N_2787,N_2785);
or U2834 (N_2834,N_2790,N_2795);
and U2835 (N_2835,N_2796,N_2786);
nand U2836 (N_2836,N_2781,N_2786);
nor U2837 (N_2837,N_2777,N_2762);
nand U2838 (N_2838,N_2764,N_2752);
nand U2839 (N_2839,N_2797,N_2766);
nand U2840 (N_2840,N_2784,N_2763);
or U2841 (N_2841,N_2763,N_2753);
and U2842 (N_2842,N_2764,N_2798);
and U2843 (N_2843,N_2786,N_2764);
nand U2844 (N_2844,N_2767,N_2775);
or U2845 (N_2845,N_2794,N_2766);
nor U2846 (N_2846,N_2786,N_2766);
or U2847 (N_2847,N_2776,N_2753);
nor U2848 (N_2848,N_2761,N_2799);
nor U2849 (N_2849,N_2754,N_2766);
nand U2850 (N_2850,N_2802,N_2833);
nand U2851 (N_2851,N_2842,N_2815);
and U2852 (N_2852,N_2828,N_2829);
or U2853 (N_2853,N_2844,N_2805);
and U2854 (N_2854,N_2837,N_2835);
and U2855 (N_2855,N_2807,N_2831);
or U2856 (N_2856,N_2813,N_2808);
nand U2857 (N_2857,N_2832,N_2830);
nor U2858 (N_2858,N_2848,N_2800);
and U2859 (N_2859,N_2801,N_2817);
or U2860 (N_2860,N_2804,N_2824);
or U2861 (N_2861,N_2819,N_2843);
nor U2862 (N_2862,N_2809,N_2838);
or U2863 (N_2863,N_2812,N_2847);
nor U2864 (N_2864,N_2834,N_2818);
nand U2865 (N_2865,N_2849,N_2839);
nor U2866 (N_2866,N_2820,N_2822);
nand U2867 (N_2867,N_2827,N_2825);
and U2868 (N_2868,N_2823,N_2826);
and U2869 (N_2869,N_2836,N_2821);
and U2870 (N_2870,N_2803,N_2845);
and U2871 (N_2871,N_2846,N_2814);
and U2872 (N_2872,N_2811,N_2810);
or U2873 (N_2873,N_2841,N_2840);
nand U2874 (N_2874,N_2816,N_2806);
and U2875 (N_2875,N_2832,N_2840);
nor U2876 (N_2876,N_2810,N_2822);
nor U2877 (N_2877,N_2811,N_2801);
nand U2878 (N_2878,N_2832,N_2826);
or U2879 (N_2879,N_2848,N_2820);
nand U2880 (N_2880,N_2845,N_2824);
nor U2881 (N_2881,N_2811,N_2821);
nand U2882 (N_2882,N_2806,N_2810);
nor U2883 (N_2883,N_2838,N_2817);
or U2884 (N_2884,N_2847,N_2818);
nor U2885 (N_2885,N_2803,N_2835);
and U2886 (N_2886,N_2833,N_2804);
nor U2887 (N_2887,N_2824,N_2801);
and U2888 (N_2888,N_2842,N_2803);
and U2889 (N_2889,N_2846,N_2818);
nor U2890 (N_2890,N_2802,N_2821);
nor U2891 (N_2891,N_2807,N_2819);
or U2892 (N_2892,N_2826,N_2839);
or U2893 (N_2893,N_2813,N_2835);
nor U2894 (N_2894,N_2846,N_2824);
or U2895 (N_2895,N_2823,N_2803);
and U2896 (N_2896,N_2823,N_2822);
and U2897 (N_2897,N_2810,N_2809);
or U2898 (N_2898,N_2808,N_2841);
and U2899 (N_2899,N_2820,N_2819);
nor U2900 (N_2900,N_2885,N_2886);
nand U2901 (N_2901,N_2893,N_2889);
nand U2902 (N_2902,N_2867,N_2879);
nor U2903 (N_2903,N_2873,N_2875);
nand U2904 (N_2904,N_2850,N_2877);
and U2905 (N_2905,N_2895,N_2878);
and U2906 (N_2906,N_2899,N_2896);
nand U2907 (N_2907,N_2861,N_2862);
nor U2908 (N_2908,N_2892,N_2872);
nor U2909 (N_2909,N_2881,N_2870);
and U2910 (N_2910,N_2883,N_2866);
and U2911 (N_2911,N_2852,N_2859);
or U2912 (N_2912,N_2891,N_2871);
and U2913 (N_2913,N_2856,N_2884);
nor U2914 (N_2914,N_2865,N_2854);
nor U2915 (N_2915,N_2897,N_2855);
or U2916 (N_2916,N_2868,N_2860);
or U2917 (N_2917,N_2882,N_2858);
and U2918 (N_2918,N_2864,N_2863);
nand U2919 (N_2919,N_2869,N_2853);
or U2920 (N_2920,N_2851,N_2894);
or U2921 (N_2921,N_2857,N_2887);
nor U2922 (N_2922,N_2888,N_2898);
nor U2923 (N_2923,N_2890,N_2876);
nand U2924 (N_2924,N_2874,N_2880);
or U2925 (N_2925,N_2865,N_2876);
and U2926 (N_2926,N_2884,N_2881);
or U2927 (N_2927,N_2899,N_2867);
nand U2928 (N_2928,N_2891,N_2853);
nor U2929 (N_2929,N_2867,N_2866);
and U2930 (N_2930,N_2877,N_2897);
or U2931 (N_2931,N_2898,N_2872);
and U2932 (N_2932,N_2893,N_2868);
and U2933 (N_2933,N_2880,N_2870);
nor U2934 (N_2934,N_2887,N_2867);
nor U2935 (N_2935,N_2852,N_2892);
or U2936 (N_2936,N_2875,N_2891);
and U2937 (N_2937,N_2851,N_2858);
nor U2938 (N_2938,N_2872,N_2852);
nor U2939 (N_2939,N_2856,N_2869);
nand U2940 (N_2940,N_2854,N_2893);
or U2941 (N_2941,N_2899,N_2862);
nand U2942 (N_2942,N_2879,N_2854);
and U2943 (N_2943,N_2883,N_2872);
nand U2944 (N_2944,N_2899,N_2888);
nand U2945 (N_2945,N_2880,N_2878);
and U2946 (N_2946,N_2850,N_2851);
or U2947 (N_2947,N_2866,N_2891);
nor U2948 (N_2948,N_2861,N_2865);
and U2949 (N_2949,N_2869,N_2867);
or U2950 (N_2950,N_2943,N_2900);
nand U2951 (N_2951,N_2927,N_2902);
and U2952 (N_2952,N_2918,N_2912);
nor U2953 (N_2953,N_2944,N_2909);
nand U2954 (N_2954,N_2920,N_2901);
and U2955 (N_2955,N_2946,N_2911);
nand U2956 (N_2956,N_2921,N_2941);
and U2957 (N_2957,N_2907,N_2948);
and U2958 (N_2958,N_2906,N_2942);
or U2959 (N_2959,N_2914,N_2945);
or U2960 (N_2960,N_2947,N_2919);
nand U2961 (N_2961,N_2933,N_2926);
nor U2962 (N_2962,N_2939,N_2923);
and U2963 (N_2963,N_2937,N_2904);
nor U2964 (N_2964,N_2932,N_2931);
nand U2965 (N_2965,N_2930,N_2903);
and U2966 (N_2966,N_2929,N_2915);
nand U2967 (N_2967,N_2922,N_2917);
nor U2968 (N_2968,N_2908,N_2925);
or U2969 (N_2969,N_2928,N_2924);
and U2970 (N_2970,N_2935,N_2938);
and U2971 (N_2971,N_2916,N_2934);
or U2972 (N_2972,N_2913,N_2949);
nor U2973 (N_2973,N_2905,N_2936);
and U2974 (N_2974,N_2940,N_2910);
and U2975 (N_2975,N_2935,N_2947);
nor U2976 (N_2976,N_2946,N_2902);
or U2977 (N_2977,N_2925,N_2919);
and U2978 (N_2978,N_2947,N_2911);
nor U2979 (N_2979,N_2943,N_2949);
and U2980 (N_2980,N_2904,N_2902);
and U2981 (N_2981,N_2907,N_2921);
and U2982 (N_2982,N_2916,N_2929);
and U2983 (N_2983,N_2900,N_2935);
and U2984 (N_2984,N_2919,N_2949);
nand U2985 (N_2985,N_2928,N_2926);
nor U2986 (N_2986,N_2902,N_2910);
or U2987 (N_2987,N_2912,N_2943);
nor U2988 (N_2988,N_2927,N_2922);
and U2989 (N_2989,N_2902,N_2920);
or U2990 (N_2990,N_2915,N_2925);
or U2991 (N_2991,N_2928,N_2908);
nor U2992 (N_2992,N_2922,N_2930);
nor U2993 (N_2993,N_2908,N_2949);
and U2994 (N_2994,N_2937,N_2941);
nor U2995 (N_2995,N_2938,N_2917);
nor U2996 (N_2996,N_2920,N_2933);
nand U2997 (N_2997,N_2901,N_2944);
or U2998 (N_2998,N_2948,N_2942);
and U2999 (N_2999,N_2916,N_2942);
nand UO_0 (O_0,N_2952,N_2978);
nor UO_1 (O_1,N_2959,N_2982);
or UO_2 (O_2,N_2998,N_2975);
or UO_3 (O_3,N_2981,N_2954);
or UO_4 (O_4,N_2955,N_2994);
nor UO_5 (O_5,N_2969,N_2951);
nor UO_6 (O_6,N_2960,N_2950);
nand UO_7 (O_7,N_2958,N_2963);
or UO_8 (O_8,N_2983,N_2990);
and UO_9 (O_9,N_2999,N_2984);
nor UO_10 (O_10,N_2989,N_2966);
nor UO_11 (O_11,N_2973,N_2956);
nand UO_12 (O_12,N_2957,N_2961);
nor UO_13 (O_13,N_2992,N_2977);
or UO_14 (O_14,N_2991,N_2967);
nand UO_15 (O_15,N_2979,N_2988);
and UO_16 (O_16,N_2980,N_2968);
or UO_17 (O_17,N_2965,N_2987);
nor UO_18 (O_18,N_2953,N_2993);
nand UO_19 (O_19,N_2962,N_2985);
or UO_20 (O_20,N_2964,N_2971);
nor UO_21 (O_21,N_2974,N_2995);
and UO_22 (O_22,N_2986,N_2976);
nor UO_23 (O_23,N_2972,N_2996);
or UO_24 (O_24,N_2997,N_2970);
or UO_25 (O_25,N_2975,N_2977);
and UO_26 (O_26,N_2951,N_2954);
nor UO_27 (O_27,N_2962,N_2967);
nand UO_28 (O_28,N_2981,N_2994);
nand UO_29 (O_29,N_2952,N_2951);
and UO_30 (O_30,N_2976,N_2977);
or UO_31 (O_31,N_2994,N_2997);
nand UO_32 (O_32,N_2963,N_2994);
nand UO_33 (O_33,N_2979,N_2950);
nand UO_34 (O_34,N_2996,N_2967);
and UO_35 (O_35,N_2963,N_2977);
and UO_36 (O_36,N_2978,N_2984);
nor UO_37 (O_37,N_2983,N_2991);
and UO_38 (O_38,N_2953,N_2975);
nand UO_39 (O_39,N_2989,N_2994);
nand UO_40 (O_40,N_2980,N_2999);
nand UO_41 (O_41,N_2992,N_2987);
or UO_42 (O_42,N_2985,N_2968);
or UO_43 (O_43,N_2958,N_2977);
xnor UO_44 (O_44,N_2952,N_2968);
and UO_45 (O_45,N_2970,N_2966);
nand UO_46 (O_46,N_2970,N_2968);
nor UO_47 (O_47,N_2977,N_2952);
nand UO_48 (O_48,N_2995,N_2961);
or UO_49 (O_49,N_2992,N_2978);
and UO_50 (O_50,N_2993,N_2973);
or UO_51 (O_51,N_2980,N_2972);
nand UO_52 (O_52,N_2973,N_2985);
nand UO_53 (O_53,N_2953,N_2960);
nand UO_54 (O_54,N_2974,N_2960);
and UO_55 (O_55,N_2953,N_2985);
nand UO_56 (O_56,N_2970,N_2972);
nor UO_57 (O_57,N_2996,N_2966);
or UO_58 (O_58,N_2986,N_2956);
and UO_59 (O_59,N_2960,N_2954);
nor UO_60 (O_60,N_2970,N_2996);
nor UO_61 (O_61,N_2980,N_2996);
nor UO_62 (O_62,N_2969,N_2971);
nand UO_63 (O_63,N_2965,N_2982);
nor UO_64 (O_64,N_2961,N_2951);
and UO_65 (O_65,N_2972,N_2954);
and UO_66 (O_66,N_2963,N_2982);
or UO_67 (O_67,N_2996,N_2974);
nand UO_68 (O_68,N_2959,N_2971);
and UO_69 (O_69,N_2976,N_2993);
and UO_70 (O_70,N_2980,N_2991);
nor UO_71 (O_71,N_2992,N_2976);
nor UO_72 (O_72,N_2984,N_2957);
and UO_73 (O_73,N_2971,N_2997);
and UO_74 (O_74,N_2997,N_2962);
xor UO_75 (O_75,N_2990,N_2977);
or UO_76 (O_76,N_2982,N_2968);
nor UO_77 (O_77,N_2955,N_2970);
nand UO_78 (O_78,N_2975,N_2964);
nor UO_79 (O_79,N_2957,N_2960);
or UO_80 (O_80,N_2983,N_2982);
or UO_81 (O_81,N_2986,N_2954);
nor UO_82 (O_82,N_2957,N_2987);
nor UO_83 (O_83,N_2987,N_2959);
nand UO_84 (O_84,N_2998,N_2952);
nand UO_85 (O_85,N_2984,N_2954);
and UO_86 (O_86,N_2963,N_2974);
nand UO_87 (O_87,N_2962,N_2969);
nand UO_88 (O_88,N_2963,N_2953);
or UO_89 (O_89,N_2956,N_2955);
nor UO_90 (O_90,N_2975,N_2989);
and UO_91 (O_91,N_2970,N_2957);
and UO_92 (O_92,N_2953,N_2961);
and UO_93 (O_93,N_2996,N_2954);
nor UO_94 (O_94,N_2950,N_2991);
or UO_95 (O_95,N_2955,N_2964);
nand UO_96 (O_96,N_2955,N_2967);
nor UO_97 (O_97,N_2999,N_2974);
or UO_98 (O_98,N_2987,N_2986);
nor UO_99 (O_99,N_2984,N_2970);
and UO_100 (O_100,N_2991,N_2993);
or UO_101 (O_101,N_2963,N_2992);
nand UO_102 (O_102,N_2971,N_2966);
or UO_103 (O_103,N_2971,N_2998);
nand UO_104 (O_104,N_2974,N_2979);
and UO_105 (O_105,N_2958,N_2976);
nor UO_106 (O_106,N_2981,N_2968);
or UO_107 (O_107,N_2965,N_2958);
nand UO_108 (O_108,N_2965,N_2972);
nand UO_109 (O_109,N_2973,N_2978);
and UO_110 (O_110,N_2993,N_2969);
nor UO_111 (O_111,N_2961,N_2965);
and UO_112 (O_112,N_2972,N_2973);
and UO_113 (O_113,N_2978,N_2987);
nor UO_114 (O_114,N_2972,N_2977);
nand UO_115 (O_115,N_2986,N_2984);
or UO_116 (O_116,N_2963,N_2964);
nor UO_117 (O_117,N_2973,N_2984);
and UO_118 (O_118,N_2974,N_2953);
nand UO_119 (O_119,N_2984,N_2961);
or UO_120 (O_120,N_2986,N_2983);
nor UO_121 (O_121,N_2954,N_2955);
nor UO_122 (O_122,N_2966,N_2997);
nor UO_123 (O_123,N_2971,N_2950);
nand UO_124 (O_124,N_2988,N_2993);
or UO_125 (O_125,N_2953,N_2969);
nand UO_126 (O_126,N_2982,N_2961);
and UO_127 (O_127,N_2990,N_2979);
or UO_128 (O_128,N_2976,N_2973);
or UO_129 (O_129,N_2997,N_2961);
nand UO_130 (O_130,N_2984,N_2952);
nor UO_131 (O_131,N_2998,N_2950);
or UO_132 (O_132,N_2976,N_2995);
nand UO_133 (O_133,N_2997,N_2951);
nor UO_134 (O_134,N_2968,N_2988);
xnor UO_135 (O_135,N_2980,N_2997);
nor UO_136 (O_136,N_2990,N_2950);
or UO_137 (O_137,N_2984,N_2976);
nand UO_138 (O_138,N_2981,N_2999);
or UO_139 (O_139,N_2987,N_2990);
and UO_140 (O_140,N_2989,N_2952);
and UO_141 (O_141,N_2988,N_2977);
or UO_142 (O_142,N_2989,N_2981);
or UO_143 (O_143,N_2963,N_2965);
and UO_144 (O_144,N_2996,N_2993);
and UO_145 (O_145,N_2963,N_2976);
or UO_146 (O_146,N_2991,N_2982);
nand UO_147 (O_147,N_2993,N_2997);
and UO_148 (O_148,N_2957,N_2977);
or UO_149 (O_149,N_2967,N_2976);
nand UO_150 (O_150,N_2967,N_2986);
nand UO_151 (O_151,N_2996,N_2977);
or UO_152 (O_152,N_2994,N_2970);
and UO_153 (O_153,N_2961,N_2979);
or UO_154 (O_154,N_2956,N_2974);
nand UO_155 (O_155,N_2973,N_2961);
nand UO_156 (O_156,N_2978,N_2997);
xnor UO_157 (O_157,N_2977,N_2980);
or UO_158 (O_158,N_2957,N_2953);
nor UO_159 (O_159,N_2959,N_2962);
or UO_160 (O_160,N_2972,N_2978);
nor UO_161 (O_161,N_2993,N_2978);
and UO_162 (O_162,N_2951,N_2992);
or UO_163 (O_163,N_2981,N_2961);
nor UO_164 (O_164,N_2953,N_2999);
or UO_165 (O_165,N_2984,N_2951);
nand UO_166 (O_166,N_2968,N_2996);
or UO_167 (O_167,N_2986,N_2998);
nand UO_168 (O_168,N_2956,N_2977);
nor UO_169 (O_169,N_2969,N_2982);
nor UO_170 (O_170,N_2955,N_2975);
nand UO_171 (O_171,N_2954,N_2950);
or UO_172 (O_172,N_2967,N_2963);
or UO_173 (O_173,N_2966,N_2950);
nand UO_174 (O_174,N_2981,N_2957);
or UO_175 (O_175,N_2974,N_2998);
or UO_176 (O_176,N_2955,N_2976);
nand UO_177 (O_177,N_2987,N_2998);
or UO_178 (O_178,N_2987,N_2973);
or UO_179 (O_179,N_2953,N_2992);
or UO_180 (O_180,N_2984,N_2962);
or UO_181 (O_181,N_2972,N_2983);
nand UO_182 (O_182,N_2980,N_2953);
and UO_183 (O_183,N_2975,N_2992);
or UO_184 (O_184,N_2963,N_2954);
or UO_185 (O_185,N_2988,N_2990);
nor UO_186 (O_186,N_2998,N_2957);
nor UO_187 (O_187,N_2985,N_2988);
and UO_188 (O_188,N_2987,N_2956);
or UO_189 (O_189,N_2999,N_2987);
or UO_190 (O_190,N_2964,N_2983);
nand UO_191 (O_191,N_2995,N_2951);
or UO_192 (O_192,N_2961,N_2954);
and UO_193 (O_193,N_2989,N_2985);
or UO_194 (O_194,N_2997,N_2996);
or UO_195 (O_195,N_2983,N_2995);
nand UO_196 (O_196,N_2971,N_2965);
or UO_197 (O_197,N_2983,N_2996);
nor UO_198 (O_198,N_2981,N_2951);
or UO_199 (O_199,N_2960,N_2978);
nor UO_200 (O_200,N_2966,N_2976);
or UO_201 (O_201,N_2976,N_2989);
or UO_202 (O_202,N_2994,N_2967);
nor UO_203 (O_203,N_2959,N_2958);
nor UO_204 (O_204,N_2994,N_2961);
nor UO_205 (O_205,N_2977,N_2966);
or UO_206 (O_206,N_2997,N_2960);
and UO_207 (O_207,N_2991,N_2984);
and UO_208 (O_208,N_2990,N_2958);
or UO_209 (O_209,N_2986,N_2995);
or UO_210 (O_210,N_2983,N_2950);
nand UO_211 (O_211,N_2951,N_2973);
or UO_212 (O_212,N_2992,N_2967);
and UO_213 (O_213,N_2951,N_2982);
and UO_214 (O_214,N_2951,N_2956);
and UO_215 (O_215,N_2952,N_2992);
nand UO_216 (O_216,N_2959,N_2990);
xnor UO_217 (O_217,N_2963,N_2989);
and UO_218 (O_218,N_2969,N_2978);
or UO_219 (O_219,N_2970,N_2981);
or UO_220 (O_220,N_2980,N_2966);
or UO_221 (O_221,N_2993,N_2960);
and UO_222 (O_222,N_2990,N_2975);
and UO_223 (O_223,N_2995,N_2960);
xor UO_224 (O_224,N_2958,N_2971);
and UO_225 (O_225,N_2976,N_2965);
nand UO_226 (O_226,N_2990,N_2970);
or UO_227 (O_227,N_2986,N_2992);
and UO_228 (O_228,N_2958,N_2966);
and UO_229 (O_229,N_2962,N_2998);
nand UO_230 (O_230,N_2980,N_2989);
nor UO_231 (O_231,N_2990,N_2973);
or UO_232 (O_232,N_2976,N_2974);
nand UO_233 (O_233,N_2971,N_2990);
xor UO_234 (O_234,N_2976,N_2991);
nand UO_235 (O_235,N_2998,N_2999);
or UO_236 (O_236,N_2968,N_2958);
or UO_237 (O_237,N_2996,N_2988);
nand UO_238 (O_238,N_2970,N_2954);
nand UO_239 (O_239,N_2998,N_2981);
nand UO_240 (O_240,N_2986,N_2981);
nand UO_241 (O_241,N_2959,N_2989);
nand UO_242 (O_242,N_2953,N_2964);
and UO_243 (O_243,N_2957,N_2993);
nor UO_244 (O_244,N_2970,N_2956);
nor UO_245 (O_245,N_2971,N_2987);
and UO_246 (O_246,N_2972,N_2955);
nand UO_247 (O_247,N_2977,N_2960);
nor UO_248 (O_248,N_2959,N_2976);
and UO_249 (O_249,N_2964,N_2995);
or UO_250 (O_250,N_2957,N_2969);
or UO_251 (O_251,N_2956,N_2989);
or UO_252 (O_252,N_2953,N_2958);
or UO_253 (O_253,N_2987,N_2993);
and UO_254 (O_254,N_2990,N_2996);
and UO_255 (O_255,N_2972,N_2979);
and UO_256 (O_256,N_2955,N_2960);
nand UO_257 (O_257,N_2968,N_2951);
or UO_258 (O_258,N_2997,N_2981);
or UO_259 (O_259,N_2989,N_2979);
or UO_260 (O_260,N_2953,N_2955);
nand UO_261 (O_261,N_2963,N_2985);
and UO_262 (O_262,N_2991,N_2966);
nor UO_263 (O_263,N_2963,N_2995);
or UO_264 (O_264,N_2993,N_2990);
xnor UO_265 (O_265,N_2965,N_2975);
and UO_266 (O_266,N_2972,N_2997);
and UO_267 (O_267,N_2990,N_2965);
nand UO_268 (O_268,N_2994,N_2993);
nand UO_269 (O_269,N_2996,N_2962);
and UO_270 (O_270,N_2999,N_2986);
and UO_271 (O_271,N_2978,N_2991);
or UO_272 (O_272,N_2999,N_2950);
and UO_273 (O_273,N_2985,N_2983);
nand UO_274 (O_274,N_2991,N_2996);
nand UO_275 (O_275,N_2966,N_2995);
nor UO_276 (O_276,N_2950,N_2995);
and UO_277 (O_277,N_2990,N_2981);
nand UO_278 (O_278,N_2985,N_2994);
or UO_279 (O_279,N_2988,N_2997);
nand UO_280 (O_280,N_2955,N_2951);
nor UO_281 (O_281,N_2993,N_2979);
and UO_282 (O_282,N_2950,N_2988);
nand UO_283 (O_283,N_2990,N_2966);
and UO_284 (O_284,N_2987,N_2958);
and UO_285 (O_285,N_2994,N_2991);
or UO_286 (O_286,N_2993,N_2962);
or UO_287 (O_287,N_2980,N_2964);
nor UO_288 (O_288,N_2979,N_2992);
or UO_289 (O_289,N_2983,N_2957);
nand UO_290 (O_290,N_2955,N_2985);
or UO_291 (O_291,N_2977,N_2959);
or UO_292 (O_292,N_2992,N_2960);
and UO_293 (O_293,N_2965,N_2983);
nor UO_294 (O_294,N_2952,N_2980);
nor UO_295 (O_295,N_2965,N_2980);
or UO_296 (O_296,N_2981,N_2950);
nand UO_297 (O_297,N_2985,N_2970);
or UO_298 (O_298,N_2951,N_2993);
and UO_299 (O_299,N_2981,N_2974);
nand UO_300 (O_300,N_2953,N_2997);
or UO_301 (O_301,N_2974,N_2954);
nor UO_302 (O_302,N_2956,N_2992);
nor UO_303 (O_303,N_2959,N_2961);
and UO_304 (O_304,N_2985,N_2995);
or UO_305 (O_305,N_2964,N_2990);
or UO_306 (O_306,N_2953,N_2996);
or UO_307 (O_307,N_2957,N_2990);
nand UO_308 (O_308,N_2969,N_2981);
and UO_309 (O_309,N_2952,N_2991);
and UO_310 (O_310,N_2994,N_2999);
or UO_311 (O_311,N_2972,N_2986);
and UO_312 (O_312,N_2974,N_2983);
and UO_313 (O_313,N_2955,N_2968);
or UO_314 (O_314,N_2989,N_2960);
or UO_315 (O_315,N_2952,N_2995);
nand UO_316 (O_316,N_2983,N_2968);
nor UO_317 (O_317,N_2975,N_2987);
nor UO_318 (O_318,N_2992,N_2974);
nor UO_319 (O_319,N_2991,N_2977);
or UO_320 (O_320,N_2970,N_2950);
and UO_321 (O_321,N_2965,N_2986);
or UO_322 (O_322,N_2998,N_2961);
and UO_323 (O_323,N_2989,N_2954);
nand UO_324 (O_324,N_2956,N_2968);
or UO_325 (O_325,N_2980,N_2984);
nor UO_326 (O_326,N_2987,N_2967);
and UO_327 (O_327,N_2999,N_2955);
and UO_328 (O_328,N_2961,N_2983);
nor UO_329 (O_329,N_2964,N_2989);
nor UO_330 (O_330,N_2955,N_2979);
or UO_331 (O_331,N_2990,N_2978);
or UO_332 (O_332,N_2988,N_2952);
or UO_333 (O_333,N_2990,N_2997);
nor UO_334 (O_334,N_2955,N_2982);
and UO_335 (O_335,N_2976,N_2999);
and UO_336 (O_336,N_2997,N_2959);
and UO_337 (O_337,N_2971,N_2960);
nand UO_338 (O_338,N_2969,N_2992);
nor UO_339 (O_339,N_2999,N_2973);
and UO_340 (O_340,N_2973,N_2991);
and UO_341 (O_341,N_2996,N_2975);
nor UO_342 (O_342,N_2984,N_2964);
or UO_343 (O_343,N_2965,N_2998);
and UO_344 (O_344,N_2976,N_2950);
and UO_345 (O_345,N_2976,N_2961);
or UO_346 (O_346,N_2975,N_2957);
and UO_347 (O_347,N_2978,N_2995);
and UO_348 (O_348,N_2957,N_2982);
and UO_349 (O_349,N_2980,N_2978);
nor UO_350 (O_350,N_2992,N_2973);
or UO_351 (O_351,N_2967,N_2951);
or UO_352 (O_352,N_2985,N_2950);
nor UO_353 (O_353,N_2960,N_2969);
nor UO_354 (O_354,N_2989,N_2997);
and UO_355 (O_355,N_2976,N_2956);
or UO_356 (O_356,N_2956,N_2960);
or UO_357 (O_357,N_2985,N_2979);
or UO_358 (O_358,N_2995,N_2959);
nor UO_359 (O_359,N_2972,N_2951);
and UO_360 (O_360,N_2988,N_2960);
nand UO_361 (O_361,N_2968,N_2975);
and UO_362 (O_362,N_2986,N_2971);
nand UO_363 (O_363,N_2958,N_2970);
nand UO_364 (O_364,N_2979,N_2960);
and UO_365 (O_365,N_2956,N_2953);
nor UO_366 (O_366,N_2978,N_2965);
and UO_367 (O_367,N_2969,N_2984);
nand UO_368 (O_368,N_2975,N_2988);
nor UO_369 (O_369,N_2950,N_2968);
and UO_370 (O_370,N_2967,N_2954);
and UO_371 (O_371,N_2951,N_2950);
nand UO_372 (O_372,N_2961,N_2963);
or UO_373 (O_373,N_2993,N_2971);
nor UO_374 (O_374,N_2989,N_2992);
and UO_375 (O_375,N_2952,N_2969);
nor UO_376 (O_376,N_2966,N_2959);
and UO_377 (O_377,N_2972,N_2950);
nand UO_378 (O_378,N_2991,N_2957);
and UO_379 (O_379,N_2995,N_2971);
or UO_380 (O_380,N_2954,N_2976);
or UO_381 (O_381,N_2967,N_2971);
and UO_382 (O_382,N_2976,N_2972);
and UO_383 (O_383,N_2971,N_2983);
and UO_384 (O_384,N_2966,N_2955);
and UO_385 (O_385,N_2969,N_2967);
or UO_386 (O_386,N_2985,N_2998);
nor UO_387 (O_387,N_2991,N_2961);
and UO_388 (O_388,N_2970,N_2998);
and UO_389 (O_389,N_2968,N_2977);
nor UO_390 (O_390,N_2972,N_2968);
nor UO_391 (O_391,N_2984,N_2993);
nand UO_392 (O_392,N_2986,N_2952);
or UO_393 (O_393,N_2994,N_2973);
nor UO_394 (O_394,N_2980,N_2971);
nand UO_395 (O_395,N_2954,N_2977);
or UO_396 (O_396,N_2985,N_2975);
or UO_397 (O_397,N_2989,N_2971);
or UO_398 (O_398,N_2994,N_2951);
and UO_399 (O_399,N_2989,N_2984);
or UO_400 (O_400,N_2957,N_2986);
or UO_401 (O_401,N_2959,N_2950);
or UO_402 (O_402,N_2993,N_2975);
and UO_403 (O_403,N_2961,N_2980);
or UO_404 (O_404,N_2968,N_2957);
and UO_405 (O_405,N_2970,N_2991);
or UO_406 (O_406,N_2972,N_2975);
or UO_407 (O_407,N_2979,N_2991);
nand UO_408 (O_408,N_2968,N_2984);
and UO_409 (O_409,N_2995,N_2977);
and UO_410 (O_410,N_2962,N_2957);
nand UO_411 (O_411,N_2982,N_2993);
or UO_412 (O_412,N_2982,N_2967);
and UO_413 (O_413,N_2967,N_2965);
and UO_414 (O_414,N_2991,N_2962);
nor UO_415 (O_415,N_2968,N_2999);
nand UO_416 (O_416,N_2979,N_2999);
and UO_417 (O_417,N_2953,N_2988);
or UO_418 (O_418,N_2958,N_2995);
and UO_419 (O_419,N_2991,N_2985);
and UO_420 (O_420,N_2970,N_2986);
nor UO_421 (O_421,N_2976,N_2953);
nor UO_422 (O_422,N_2963,N_2975);
or UO_423 (O_423,N_2951,N_2965);
and UO_424 (O_424,N_2974,N_2950);
or UO_425 (O_425,N_2977,N_2982);
and UO_426 (O_426,N_2981,N_2996);
nand UO_427 (O_427,N_2961,N_2989);
nand UO_428 (O_428,N_2953,N_2959);
and UO_429 (O_429,N_2990,N_2956);
and UO_430 (O_430,N_2990,N_2969);
and UO_431 (O_431,N_2992,N_2982);
and UO_432 (O_432,N_2956,N_2964);
nor UO_433 (O_433,N_2991,N_2974);
and UO_434 (O_434,N_2965,N_2995);
and UO_435 (O_435,N_2950,N_2969);
xnor UO_436 (O_436,N_2994,N_2952);
and UO_437 (O_437,N_2976,N_2981);
nor UO_438 (O_438,N_2967,N_2956);
nand UO_439 (O_439,N_2987,N_2977);
or UO_440 (O_440,N_2995,N_2970);
or UO_441 (O_441,N_2979,N_2957);
xor UO_442 (O_442,N_2966,N_2953);
or UO_443 (O_443,N_2987,N_2961);
or UO_444 (O_444,N_2972,N_2963);
nor UO_445 (O_445,N_2999,N_2972);
and UO_446 (O_446,N_2983,N_2987);
or UO_447 (O_447,N_2959,N_2970);
and UO_448 (O_448,N_2964,N_2993);
or UO_449 (O_449,N_2968,N_2966);
nand UO_450 (O_450,N_2959,N_2965);
or UO_451 (O_451,N_2988,N_2971);
nand UO_452 (O_452,N_2964,N_2967);
nand UO_453 (O_453,N_2965,N_2974);
or UO_454 (O_454,N_2985,N_2980);
and UO_455 (O_455,N_2971,N_2975);
and UO_456 (O_456,N_2990,N_2980);
nand UO_457 (O_457,N_2970,N_2977);
nor UO_458 (O_458,N_2954,N_2987);
nand UO_459 (O_459,N_2957,N_2994);
or UO_460 (O_460,N_2960,N_2998);
nand UO_461 (O_461,N_2996,N_2963);
or UO_462 (O_462,N_2981,N_2952);
nor UO_463 (O_463,N_2999,N_2962);
and UO_464 (O_464,N_2988,N_2992);
nor UO_465 (O_465,N_2984,N_2982);
nand UO_466 (O_466,N_2957,N_2951);
and UO_467 (O_467,N_2955,N_2981);
nand UO_468 (O_468,N_2984,N_2990);
nor UO_469 (O_469,N_2994,N_2978);
nor UO_470 (O_470,N_2968,N_2990);
nor UO_471 (O_471,N_2963,N_2959);
nor UO_472 (O_472,N_2990,N_2995);
and UO_473 (O_473,N_2994,N_2968);
nor UO_474 (O_474,N_2956,N_2950);
or UO_475 (O_475,N_2958,N_2961);
nor UO_476 (O_476,N_2969,N_2958);
and UO_477 (O_477,N_2972,N_2964);
xnor UO_478 (O_478,N_2989,N_2993);
and UO_479 (O_479,N_2967,N_2966);
nor UO_480 (O_480,N_2952,N_2961);
and UO_481 (O_481,N_2980,N_2973);
or UO_482 (O_482,N_2996,N_2961);
and UO_483 (O_483,N_2978,N_2989);
nand UO_484 (O_484,N_2968,N_2973);
or UO_485 (O_485,N_2952,N_2958);
nor UO_486 (O_486,N_2954,N_2997);
and UO_487 (O_487,N_2981,N_2988);
or UO_488 (O_488,N_2973,N_2981);
nand UO_489 (O_489,N_2987,N_2976);
nand UO_490 (O_490,N_2967,N_2984);
nor UO_491 (O_491,N_2955,N_2957);
or UO_492 (O_492,N_2975,N_2961);
and UO_493 (O_493,N_2965,N_2950);
and UO_494 (O_494,N_2963,N_2984);
or UO_495 (O_495,N_2970,N_2980);
and UO_496 (O_496,N_2970,N_2971);
and UO_497 (O_497,N_2983,N_2952);
nand UO_498 (O_498,N_2974,N_2990);
nand UO_499 (O_499,N_2989,N_2967);
endmodule