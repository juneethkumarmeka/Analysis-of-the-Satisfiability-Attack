module basic_1500_15000_2000_5_levels_10xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
nand U0 (N_0,In_98,In_950);
xnor U1 (N_1,In_1377,In_824);
nand U2 (N_2,In_242,In_794);
and U3 (N_3,In_1476,In_403);
nor U4 (N_4,In_84,In_9);
or U5 (N_5,In_838,In_1398);
nand U6 (N_6,In_1175,In_879);
xor U7 (N_7,In_1164,In_268);
nand U8 (N_8,In_72,In_478);
or U9 (N_9,In_487,In_407);
nor U10 (N_10,In_789,In_336);
nor U11 (N_11,In_833,In_469);
xnor U12 (N_12,In_1029,In_714);
nor U13 (N_13,In_992,In_1305);
nand U14 (N_14,In_607,In_1117);
nand U15 (N_15,In_720,In_920);
and U16 (N_16,In_539,In_708);
and U17 (N_17,In_322,In_1044);
or U18 (N_18,In_1439,In_370);
and U19 (N_19,In_381,In_1201);
nand U20 (N_20,In_145,In_776);
nand U21 (N_21,In_1437,In_1079);
nand U22 (N_22,In_1453,In_1276);
and U23 (N_23,In_673,In_740);
nand U24 (N_24,In_626,In_25);
nor U25 (N_25,In_1241,In_1351);
nand U26 (N_26,In_1093,In_812);
nor U27 (N_27,In_1180,In_817);
xor U28 (N_28,In_951,In_1422);
nor U29 (N_29,In_560,In_259);
or U30 (N_30,In_520,In_1178);
xor U31 (N_31,In_711,In_877);
xnor U32 (N_32,In_994,In_411);
xor U33 (N_33,In_173,In_266);
or U34 (N_34,In_1378,In_65);
nor U35 (N_35,In_77,In_479);
nor U36 (N_36,In_86,In_1361);
and U37 (N_37,In_438,In_21);
or U38 (N_38,In_1163,In_335);
nor U39 (N_39,In_839,In_495);
or U40 (N_40,In_1233,In_346);
and U41 (N_41,In_953,In_409);
or U42 (N_42,In_429,In_1033);
xor U43 (N_43,In_1129,In_451);
or U44 (N_44,In_784,In_1100);
nor U45 (N_45,In_822,In_538);
nor U46 (N_46,In_739,In_929);
nor U47 (N_47,In_219,In_301);
or U48 (N_48,In_884,In_428);
nand U49 (N_49,In_496,In_730);
nand U50 (N_50,In_800,In_97);
or U51 (N_51,In_1206,In_375);
or U52 (N_52,In_27,In_1463);
xnor U53 (N_53,In_589,In_347);
or U54 (N_54,In_30,In_926);
and U55 (N_55,In_1282,In_666);
xnor U56 (N_56,In_1401,In_1457);
or U57 (N_57,In_417,In_1096);
xnor U58 (N_58,In_540,In_1406);
xor U59 (N_59,In_1389,In_2);
or U60 (N_60,In_113,In_1462);
nor U61 (N_61,In_1022,In_1386);
or U62 (N_62,In_1006,In_224);
nor U63 (N_63,In_1298,In_1034);
or U64 (N_64,In_859,In_352);
nand U65 (N_65,In_1396,In_1397);
xor U66 (N_66,In_803,In_401);
nor U67 (N_67,In_677,In_1458);
and U68 (N_68,In_296,In_15);
or U69 (N_69,In_881,In_94);
xnor U70 (N_70,In_531,In_311);
xnor U71 (N_71,In_191,In_826);
nand U72 (N_72,In_661,In_1204);
nand U73 (N_73,In_1465,In_781);
nor U74 (N_74,In_1092,In_362);
nor U75 (N_75,In_549,In_155);
and U76 (N_76,In_1318,In_737);
or U77 (N_77,In_547,In_842);
and U78 (N_78,In_1207,In_984);
or U79 (N_79,In_111,In_947);
nor U80 (N_80,In_1359,In_138);
nor U81 (N_81,In_265,In_535);
nand U82 (N_82,In_1292,In_100);
nand U83 (N_83,In_351,In_218);
xnor U84 (N_84,In_328,In_1496);
and U85 (N_85,In_184,In_384);
nor U86 (N_86,In_1407,In_485);
and U87 (N_87,In_1139,In_456);
nor U88 (N_88,In_277,In_1347);
nand U89 (N_89,In_90,In_1340);
and U90 (N_90,In_443,In_169);
nor U91 (N_91,In_371,In_543);
or U92 (N_92,In_503,In_735);
or U93 (N_93,In_69,In_732);
or U94 (N_94,In_857,In_189);
nor U95 (N_95,In_1057,In_1333);
nor U96 (N_96,In_132,In_193);
nand U97 (N_97,In_837,In_1294);
nand U98 (N_98,In_1098,In_147);
xnor U99 (N_99,In_596,In_629);
or U100 (N_100,In_1099,In_287);
nor U101 (N_101,In_576,In_57);
or U102 (N_102,In_572,In_960);
xnor U103 (N_103,In_70,In_868);
xor U104 (N_104,In_562,In_1144);
xnor U105 (N_105,In_742,In_1425);
nor U106 (N_106,In_280,In_378);
xor U107 (N_107,In_1337,In_778);
or U108 (N_108,In_813,In_671);
nand U109 (N_109,In_913,In_1312);
nor U110 (N_110,In_302,In_1162);
nor U111 (N_111,In_315,In_1459);
nor U112 (N_112,In_324,In_927);
and U113 (N_113,In_1372,In_873);
xor U114 (N_114,In_1274,In_472);
or U115 (N_115,In_627,In_849);
xor U116 (N_116,In_208,In_13);
or U117 (N_117,In_1370,In_1141);
xor U118 (N_118,In_1393,In_751);
nand U119 (N_119,In_1332,In_1160);
or U120 (N_120,In_1106,In_1125);
nor U121 (N_121,In_633,In_88);
or U122 (N_122,In_1155,In_151);
nand U123 (N_123,In_886,In_1188);
nand U124 (N_124,In_1364,In_710);
nand U125 (N_125,In_554,In_441);
nor U126 (N_126,In_507,In_1115);
xnor U127 (N_127,In_1183,In_119);
or U128 (N_128,In_187,In_582);
xor U129 (N_129,In_1421,In_665);
xnor U130 (N_130,In_148,In_488);
xnor U131 (N_131,In_1140,In_103);
nand U132 (N_132,In_1086,In_439);
and U133 (N_133,In_1105,In_1260);
or U134 (N_134,In_772,In_230);
or U135 (N_135,In_284,In_660);
xnor U136 (N_136,In_593,In_83);
and U137 (N_137,In_1071,In_166);
nor U138 (N_138,In_618,In_917);
nand U139 (N_139,In_275,In_434);
nand U140 (N_140,In_934,In_75);
or U141 (N_141,In_963,In_1084);
xnor U142 (N_142,In_855,In_762);
xnor U143 (N_143,In_1280,In_449);
or U144 (N_144,In_271,In_1);
nand U145 (N_145,In_413,In_1018);
nor U146 (N_146,In_1247,In_274);
and U147 (N_147,In_47,In_1296);
xor U148 (N_148,In_484,In_1134);
and U149 (N_149,In_700,In_217);
nand U150 (N_150,In_1443,In_44);
xor U151 (N_151,In_68,In_149);
nand U152 (N_152,In_143,In_717);
or U153 (N_153,In_1118,In_432);
nand U154 (N_154,In_421,In_911);
nand U155 (N_155,In_1268,In_1264);
and U156 (N_156,In_175,In_255);
xor U157 (N_157,In_1366,In_983);
nor U158 (N_158,In_1263,In_771);
nor U159 (N_159,In_499,In_896);
nor U160 (N_160,In_402,In_999);
nand U161 (N_161,In_1246,In_1423);
and U162 (N_162,In_1116,In_508);
nand U163 (N_163,In_718,In_606);
and U164 (N_164,In_865,In_486);
or U165 (N_165,In_802,In_501);
or U166 (N_166,In_1248,In_519);
or U167 (N_167,In_621,In_204);
nor U168 (N_168,In_1197,In_634);
nor U169 (N_169,In_1266,In_974);
nor U170 (N_170,In_1059,In_131);
or U171 (N_171,In_1066,In_971);
nand U172 (N_172,In_815,In_1227);
xor U173 (N_173,In_548,In_400);
nand U174 (N_174,In_1104,In_801);
nand U175 (N_175,In_1323,In_1403);
xnor U176 (N_176,In_885,In_787);
and U177 (N_177,In_565,In_1343);
or U178 (N_178,In_1039,In_1480);
and U179 (N_179,In_910,In_105);
or U180 (N_180,In_197,In_1238);
nor U181 (N_181,In_939,In_205);
or U182 (N_182,In_91,In_723);
nand U183 (N_183,In_161,In_87);
nand U184 (N_184,In_680,In_600);
or U185 (N_185,In_141,In_74);
and U186 (N_186,In_1110,In_733);
nand U187 (N_187,In_1433,In_1293);
nor U188 (N_188,In_987,In_990);
and U189 (N_189,In_581,In_1286);
or U190 (N_190,In_142,In_36);
or U191 (N_191,In_1460,In_869);
and U192 (N_192,In_190,In_258);
nand U193 (N_193,In_566,In_1489);
xor U194 (N_194,In_1408,In_1005);
xnor U195 (N_195,In_1085,In_1038);
or U196 (N_196,In_42,In_851);
nand U197 (N_197,In_1113,In_1035);
xnor U198 (N_198,In_11,In_1017);
or U199 (N_199,In_412,In_769);
nor U200 (N_200,In_1265,In_89);
xnor U201 (N_201,In_1424,In_73);
nand U202 (N_202,In_1003,In_31);
xor U203 (N_203,In_1479,In_152);
nor U204 (N_204,In_290,In_158);
and U205 (N_205,In_110,In_599);
and U206 (N_206,In_609,In_1102);
or U207 (N_207,In_1076,In_342);
xor U208 (N_208,In_1136,In_905);
xor U209 (N_209,In_1448,In_1015);
xor U210 (N_210,In_256,In_764);
nand U211 (N_211,In_466,In_355);
nand U212 (N_212,In_32,In_1184);
nand U213 (N_213,In_808,In_343);
nand U214 (N_214,In_1088,In_631);
nand U215 (N_215,In_321,In_180);
xnor U216 (N_216,In_361,In_919);
or U217 (N_217,In_1069,In_819);
nor U218 (N_218,In_1077,In_28);
or U219 (N_219,In_1349,In_1491);
and U220 (N_220,In_1215,In_1150);
xor U221 (N_221,In_891,In_288);
nand U222 (N_222,In_592,In_1157);
nor U223 (N_223,In_1357,In_374);
nor U224 (N_224,In_568,In_1036);
and U225 (N_225,In_648,In_1000);
xnor U226 (N_226,In_688,In_796);
or U227 (N_227,In_45,In_1171);
or U228 (N_228,In_270,In_890);
xor U229 (N_229,In_1225,In_308);
nor U230 (N_230,In_1295,In_64);
or U231 (N_231,In_1189,In_492);
or U232 (N_232,In_498,In_664);
or U233 (N_233,In_745,In_228);
and U234 (N_234,In_1475,In_468);
and U235 (N_235,In_1212,In_1048);
nand U236 (N_236,In_973,In_728);
xnor U237 (N_237,In_883,In_59);
or U238 (N_238,In_852,In_127);
nor U239 (N_239,In_450,In_1242);
and U240 (N_240,In_840,In_404);
nand U241 (N_241,In_1346,In_137);
or U242 (N_242,In_1485,In_1195);
and U243 (N_243,In_1329,In_1159);
nand U244 (N_244,In_1154,In_1445);
nor U245 (N_245,In_1047,In_1056);
nor U246 (N_246,In_689,In_1254);
nand U247 (N_247,In_364,In_941);
or U248 (N_248,In_961,In_603);
nand U249 (N_249,In_367,In_620);
nand U250 (N_250,In_570,In_1371);
nor U251 (N_251,In_1373,In_853);
or U252 (N_252,In_712,In_1245);
or U253 (N_253,In_1091,In_1101);
or U254 (N_254,In_610,In_329);
or U255 (N_255,In_1031,In_1331);
and U256 (N_256,In_1146,In_139);
nor U257 (N_257,In_1257,In_989);
nor U258 (N_258,In_649,In_932);
nor U259 (N_259,In_194,In_1374);
nand U260 (N_260,In_1446,In_251);
nand U261 (N_261,In_536,In_1199);
nand U262 (N_262,In_1187,In_19);
nand U263 (N_263,In_475,In_653);
xnor U264 (N_264,In_528,In_426);
xnor U265 (N_265,In_10,In_995);
nor U266 (N_266,In_157,In_605);
nor U267 (N_267,In_53,In_415);
nand U268 (N_268,In_798,In_1275);
and U269 (N_269,In_332,In_0);
nor U270 (N_270,In_445,In_1094);
or U271 (N_271,In_870,In_1449);
nor U272 (N_272,In_1179,In_656);
nor U273 (N_273,In_368,In_1137);
and U274 (N_274,In_1114,In_1469);
or U275 (N_275,In_117,In_514);
xnor U276 (N_276,In_1481,In_588);
or U277 (N_277,In_1313,In_1454);
xor U278 (N_278,In_888,In_1440);
or U279 (N_279,In_765,In_1284);
nor U280 (N_280,In_211,In_192);
nor U281 (N_281,In_312,In_897);
xor U282 (N_282,In_976,In_1027);
xnor U283 (N_283,In_159,In_483);
or U284 (N_284,In_38,In_1169);
xnor U285 (N_285,In_325,In_965);
nor U286 (N_286,In_170,In_667);
or U287 (N_287,In_1339,In_1132);
nor U288 (N_288,In_1097,In_880);
or U289 (N_289,In_858,In_390);
nor U290 (N_290,In_1484,In_76);
nand U291 (N_291,In_1172,In_617);
and U292 (N_292,In_386,In_571);
or U293 (N_293,In_318,In_247);
nor U294 (N_294,In_510,In_383);
and U295 (N_295,In_1336,In_1367);
or U296 (N_296,In_1306,In_24);
and U297 (N_297,In_654,In_699);
xnor U298 (N_298,In_267,In_243);
nand U299 (N_299,In_1353,In_226);
and U300 (N_300,In_894,In_597);
or U301 (N_301,In_703,In_1095);
nor U302 (N_302,In_882,In_54);
nand U303 (N_303,In_422,In_1495);
nor U304 (N_304,In_624,In_210);
nand U305 (N_305,In_273,In_986);
nor U306 (N_306,In_458,In_1494);
and U307 (N_307,In_537,In_753);
nor U308 (N_308,In_970,In_788);
and U309 (N_309,In_552,In_1431);
nor U310 (N_310,In_71,In_1324);
and U311 (N_311,In_1067,In_497);
xor U312 (N_312,In_534,In_757);
xor U313 (N_313,In_731,In_1130);
xor U314 (N_314,In_254,In_467);
or U315 (N_315,In_300,In_1252);
nor U316 (N_316,In_1289,In_1391);
xnor U317 (N_317,In_202,In_1072);
xnor U318 (N_318,In_440,In_830);
and U319 (N_319,In_854,In_1123);
xor U320 (N_320,In_129,In_904);
nor U321 (N_321,In_845,In_774);
nand U322 (N_322,In_921,In_177);
nand U323 (N_323,In_200,In_188);
nor U324 (N_324,In_823,In_435);
or U325 (N_325,In_214,In_922);
and U326 (N_326,In_1471,In_602);
xnor U327 (N_327,In_293,In_783);
and U328 (N_328,In_135,In_1040);
nand U329 (N_329,In_637,In_1028);
nand U330 (N_330,In_305,In_782);
or U331 (N_331,In_178,In_282);
xnor U332 (N_332,In_1281,In_234);
or U333 (N_333,In_1277,In_835);
nor U334 (N_334,In_1412,In_1411);
nor U335 (N_335,In_662,In_348);
and U336 (N_336,In_1488,In_222);
and U337 (N_337,In_442,In_291);
nor U338 (N_338,In_517,In_1191);
and U339 (N_339,In_1490,In_697);
and U340 (N_340,In_1107,In_736);
nor U341 (N_341,In_1001,In_744);
or U342 (N_342,In_500,In_93);
and U343 (N_343,In_556,In_1473);
xor U344 (N_344,In_481,In_471);
nand U345 (N_345,In_907,In_299);
xor U346 (N_346,In_727,In_459);
xnor U347 (N_347,In_1392,In_201);
or U348 (N_348,In_345,In_1244);
nand U349 (N_349,In_12,In_542);
nor U350 (N_350,In_1236,In_1417);
nor U351 (N_351,In_1045,In_1243);
and U352 (N_352,In_793,In_559);
nor U353 (N_353,In_521,In_902);
nor U354 (N_354,In_925,In_333);
and U355 (N_355,In_220,In_1138);
xnor U356 (N_356,In_1111,In_16);
and U357 (N_357,In_779,In_674);
and U358 (N_358,In_1404,In_1438);
and U359 (N_359,In_687,In_1325);
and U360 (N_360,In_993,In_250);
and U361 (N_361,In_1258,In_692);
xnor U362 (N_362,In_1012,In_860);
and U363 (N_363,In_309,In_1149);
nor U364 (N_364,In_227,In_509);
xor U365 (N_365,In_1365,In_590);
nand U366 (N_366,In_62,In_385);
nor U367 (N_367,In_1388,In_1004);
and U368 (N_368,In_975,In_327);
and U369 (N_369,In_758,In_23);
xor U370 (N_370,In_1309,In_652);
xnor U371 (N_371,In_229,In_338);
xor U372 (N_372,In_946,In_1319);
and U373 (N_373,In_635,In_20);
nand U374 (N_374,In_636,In_901);
nor U375 (N_375,In_396,In_645);
and U376 (N_376,In_1251,In_199);
nor U377 (N_377,In_847,In_1025);
nor U378 (N_378,In_454,In_307);
and U379 (N_379,In_678,In_1315);
nand U380 (N_380,In_770,In_186);
or U381 (N_381,In_116,In_231);
xnor U382 (N_382,In_1350,In_1482);
or U383 (N_383,In_56,In_806);
nand U384 (N_384,In_625,In_1335);
and U385 (N_385,In_213,In_153);
nand U386 (N_386,In_1226,In_283);
nand U387 (N_387,In_1120,In_433);
nor U388 (N_388,In_460,In_1250);
xnor U389 (N_389,In_1083,In_795);
nor U390 (N_390,In_1415,In_330);
and U391 (N_391,In_1213,In_1121);
nor U392 (N_392,In_1043,In_33);
and U393 (N_393,In_1320,In_825);
or U394 (N_394,In_1153,In_1341);
and U395 (N_395,In_405,In_1052);
or U396 (N_396,In_414,In_874);
or U397 (N_397,In_1026,In_320);
or U398 (N_398,In_900,In_644);
nor U399 (N_399,In_829,In_780);
nor U400 (N_400,In_1426,In_423);
nand U401 (N_401,In_358,In_940);
nor U402 (N_402,In_353,In_246);
and U403 (N_403,In_1427,In_1429);
xnor U404 (N_404,In_1253,In_585);
nor U405 (N_405,In_1065,In_836);
and U406 (N_406,In_1483,In_285);
and U407 (N_407,In_1249,In_968);
or U408 (N_408,In_269,In_115);
xor U409 (N_409,In_908,In_1234);
and U410 (N_410,In_1222,In_1186);
and U411 (N_411,In_679,In_1259);
xnor U412 (N_412,In_264,In_512);
nand U413 (N_413,In_756,In_1152);
xor U414 (N_414,In_1127,In_365);
nor U415 (N_415,In_1413,In_1087);
xnor U416 (N_416,In_643,In_446);
nor U417 (N_417,In_6,In_1109);
and U418 (N_418,In_1230,In_875);
and U419 (N_419,In_1390,In_959);
or U420 (N_420,In_944,In_1419);
or U421 (N_421,In_638,In_1054);
xor U422 (N_422,In_1418,In_1356);
nor U423 (N_423,In_1135,In_40);
xor U424 (N_424,In_713,In_672);
and U425 (N_425,In_408,In_958);
and U426 (N_426,In_935,In_359);
xor U427 (N_427,In_575,In_457);
nand U428 (N_428,In_790,In_695);
nand U429 (N_429,In_533,In_1414);
nand U430 (N_430,In_489,In_930);
nor U431 (N_431,In_1394,In_1255);
nor U432 (N_432,In_1158,In_864);
or U433 (N_433,In_1002,In_912);
and U434 (N_434,In_448,In_719);
xor U435 (N_435,In_614,In_1308);
nor U436 (N_436,In_79,In_393);
nor U437 (N_437,In_1317,In_1384);
nand U438 (N_438,In_350,In_122);
and U439 (N_439,In_260,In_957);
nand U440 (N_440,In_257,In_867);
nand U441 (N_441,In_558,In_1273);
nand U442 (N_442,In_130,In_1478);
and U443 (N_443,In_1420,In_998);
nand U444 (N_444,In_474,In_761);
nand U445 (N_445,In_591,In_372);
and U446 (N_446,In_586,In_1291);
nand U447 (N_447,In_1217,In_1352);
xnor U448 (N_448,In_455,In_326);
and U449 (N_449,In_1181,In_646);
or U450 (N_450,In_1272,In_5);
xor U451 (N_451,In_235,In_430);
and U452 (N_452,In_124,In_1147);
nor U453 (N_453,In_1262,In_1058);
xnor U454 (N_454,In_373,In_918);
xor U455 (N_455,In_1030,In_453);
and U456 (N_456,In_48,In_357);
nor U457 (N_457,In_544,In_1409);
nand U458 (N_458,In_419,In_954);
and U459 (N_459,In_382,In_1148);
xor U460 (N_460,In_248,In_1124);
nand U461 (N_461,In_425,In_647);
nand U462 (N_462,In_755,In_1128);
nor U463 (N_463,In_967,In_574);
and U464 (N_464,In_1368,In_766);
nor U465 (N_465,In_55,In_1287);
and U466 (N_466,In_245,In_871);
or U467 (N_467,In_1301,In_1405);
or U468 (N_468,In_17,In_655);
or U469 (N_469,In_1185,In_1435);
nand U470 (N_470,In_948,In_239);
xor U471 (N_471,In_563,In_1170);
and U472 (N_472,In_1467,In_1279);
and U473 (N_473,In_613,In_1078);
and U474 (N_474,In_601,In_792);
or U475 (N_475,In_410,In_741);
nand U476 (N_476,In_734,In_50);
or U477 (N_477,In_690,In_377);
or U478 (N_478,In_1300,In_1432);
or U479 (N_479,In_1299,In_682);
xor U480 (N_480,In_811,In_933);
nand U481 (N_481,In_337,In_1165);
xnor U482 (N_482,In_172,In_804);
xnor U483 (N_483,In_1362,In_102);
and U484 (N_484,In_1235,In_167);
or U485 (N_485,In_786,In_1070);
xor U486 (N_486,In_1049,In_462);
xnor U487 (N_487,In_1103,In_580);
nand U488 (N_488,In_1342,In_515);
xor U489 (N_489,In_759,In_144);
nor U490 (N_490,In_982,In_1174);
or U491 (N_491,In_964,In_340);
nand U492 (N_492,In_319,In_814);
xor U493 (N_493,In_505,In_196);
or U494 (N_494,In_195,In_223);
and U495 (N_495,In_686,In_476);
or U496 (N_496,In_876,In_567);
xor U497 (N_497,In_225,In_569);
and U498 (N_498,In_58,In_1383);
nor U499 (N_499,In_545,In_991);
and U500 (N_500,In_1399,In_810);
nand U501 (N_501,In_834,In_715);
nand U502 (N_502,In_1307,In_578);
or U503 (N_503,In_1327,In_1231);
or U504 (N_504,In_316,In_709);
or U505 (N_505,In_356,In_1470);
or U506 (N_506,In_1283,In_612);
and U507 (N_507,In_694,In_221);
or U508 (N_508,In_82,In_81);
nand U509 (N_509,In_506,In_1355);
and U510 (N_510,In_388,In_154);
or U511 (N_511,In_163,In_43);
nor U512 (N_512,In_1219,In_583);
nor U513 (N_513,In_1321,In_1074);
xnor U514 (N_514,In_996,In_1173);
nand U515 (N_515,In_125,In_1024);
and U516 (N_516,In_1239,In_1486);
nand U517 (N_517,In_164,In_1014);
or U518 (N_518,In_639,In_304);
nand U519 (N_519,In_831,In_821);
or U520 (N_520,In_1211,In_640);
nor U521 (N_521,In_165,In_693);
or U522 (N_522,In_1311,In_1009);
or U523 (N_523,In_1089,In_668);
or U524 (N_524,In_121,In_705);
nand U525 (N_525,In_915,In_4);
nand U526 (N_526,In_313,In_1064);
or U527 (N_527,In_1081,In_1334);
nor U528 (N_528,In_750,In_1041);
nand U529 (N_529,In_1161,In_289);
and U530 (N_530,In_889,In_168);
and U531 (N_531,In_18,In_1063);
or U532 (N_532,In_701,In_841);
nand U533 (N_533,In_706,In_1208);
nor U534 (N_534,In_928,In_1228);
nand U535 (N_535,In_611,In_878);
nand U536 (N_536,In_1376,In_206);
nor U537 (N_537,In_936,In_615);
or U538 (N_538,In_1493,In_1011);
and U539 (N_539,In_1082,In_369);
xnor U540 (N_540,In_1382,In_1387);
nor U541 (N_541,In_397,In_395);
xor U542 (N_542,In_1013,In_791);
nor U543 (N_543,In_37,In_262);
xor U544 (N_544,In_244,In_1060);
or U545 (N_545,In_1133,In_1330);
nor U546 (N_546,In_272,In_1108);
or U547 (N_547,In_716,In_1345);
or U548 (N_548,In_518,In_1326);
and U549 (N_549,In_323,In_938);
nor U550 (N_550,In_1338,In_1073);
or U551 (N_551,In_494,In_1271);
nand U552 (N_552,In_1020,In_216);
or U553 (N_553,In_743,In_1497);
and U554 (N_554,In_238,In_773);
and U555 (N_555,In_1303,In_760);
xnor U556 (N_556,In_863,In_832);
or U557 (N_557,In_641,In_156);
xor U558 (N_558,In_241,In_1278);
nand U559 (N_559,In_525,In_314);
nand U560 (N_560,In_557,In_1410);
and U561 (N_561,In_1177,In_746);
nand U562 (N_562,In_721,In_1182);
nand U563 (N_563,In_632,In_41);
xor U564 (N_564,In_294,In_317);
nand U565 (N_565,In_988,In_140);
nor U566 (N_566,In_630,In_555);
and U567 (N_567,In_292,In_1075);
or U568 (N_568,In_887,In_777);
and U569 (N_569,In_1037,In_1285);
nor U570 (N_570,In_61,In_604);
nor U571 (N_571,In_490,In_112);
and U572 (N_572,In_1464,In_1156);
or U573 (N_573,In_1344,In_1232);
and U574 (N_574,In_797,In_1468);
nor U575 (N_575,In_980,In_34);
and U576 (N_576,In_685,In_1142);
xnor U577 (N_577,In_1267,In_1472);
nor U578 (N_578,In_1126,In_1395);
nand U579 (N_579,In_650,In_747);
and U580 (N_580,In_491,In_1050);
nor U581 (N_581,In_424,In_702);
nor U582 (N_582,In_1090,In_249);
nor U583 (N_583,In_573,In_587);
nand U584 (N_584,In_738,In_1348);
nand U585 (N_585,In_962,In_331);
or U586 (N_586,In_67,In_1112);
xnor U587 (N_587,In_843,In_844);
and U588 (N_588,In_1381,In_1270);
and U589 (N_589,In_684,In_171);
xor U590 (N_590,In_966,In_807);
nor U591 (N_591,In_399,In_14);
nand U592 (N_592,In_895,In_237);
xor U593 (N_593,In_943,In_26);
xor U594 (N_594,In_898,In_303);
and U595 (N_595,In_1198,In_704);
xnor U596 (N_596,In_502,In_848);
and U597 (N_597,In_866,In_550);
and U598 (N_598,In_376,In_1205);
or U599 (N_599,In_1354,In_146);
nand U600 (N_600,In_1256,In_1168);
xnor U601 (N_601,In_49,In_846);
nor U602 (N_602,In_985,In_516);
nor U603 (N_603,In_1229,In_561);
and U604 (N_604,In_676,In_1032);
nand U605 (N_605,In_349,In_949);
nand U606 (N_606,In_1209,In_1385);
nand U607 (N_607,In_1428,In_240);
nor U608 (N_608,In_828,In_176);
nand U609 (N_609,In_276,In_1499);
and U610 (N_610,In_181,In_80);
nor U611 (N_611,In_387,In_341);
nand U612 (N_612,In_1062,In_903);
and U613 (N_613,In_394,In_114);
nand U614 (N_614,In_447,In_598);
or U615 (N_615,In_278,In_1456);
xnor U616 (N_616,In_1216,In_752);
or U617 (N_617,In_1166,In_1042);
nor U618 (N_618,In_1498,In_1288);
or U619 (N_619,In_1360,In_945);
nor U620 (N_620,In_136,In_916);
and U621 (N_621,In_101,In_1190);
nand U622 (N_622,In_1193,In_334);
and U623 (N_623,In_51,In_546);
nand U624 (N_624,In_748,In_437);
nand U625 (N_625,In_233,In_698);
and U626 (N_626,In_109,In_452);
or U627 (N_627,In_1302,In_809);
xor U628 (N_628,In_252,In_66);
nor U629 (N_629,In_670,In_551);
or U630 (N_630,In_92,In_1466);
nand U631 (N_631,In_529,In_691);
nand U632 (N_632,In_1046,In_297);
or U633 (N_633,In_179,In_1167);
and U634 (N_634,In_579,In_1297);
xnor U635 (N_635,In_526,In_464);
xnor U636 (N_636,In_1202,In_763);
nor U637 (N_637,In_969,In_363);
or U638 (N_638,In_1008,In_1214);
xnor U639 (N_639,In_584,In_107);
or U640 (N_640,In_133,In_1363);
xor U641 (N_641,In_203,In_310);
xnor U642 (N_642,In_1218,In_1007);
xor U643 (N_643,In_937,In_981);
nor U644 (N_644,In_1444,In_420);
nand U645 (N_645,In_85,In_63);
nand U646 (N_646,In_482,In_675);
nor U647 (N_647,In_52,In_1080);
or U648 (N_648,In_924,In_398);
nand U649 (N_649,In_118,In_972);
or U650 (N_650,In_22,In_997);
and U651 (N_651,In_978,In_8);
nor U652 (N_652,In_511,In_1021);
and U653 (N_653,In_622,In_663);
nor U654 (N_654,In_389,In_1143);
or U655 (N_655,In_722,In_1379);
nand U656 (N_656,In_1261,In_295);
xor U657 (N_657,In_279,In_1369);
and U658 (N_658,In_183,In_162);
or U659 (N_659,In_150,In_1131);
nor U660 (N_660,In_391,In_1492);
or U661 (N_661,In_3,In_1224);
and U662 (N_662,In_1194,In_1461);
nand U663 (N_663,In_1203,In_522);
xnor U664 (N_664,In_174,In_726);
nor U665 (N_665,In_29,In_1122);
xor U666 (N_666,In_1455,In_470);
nor U667 (N_667,In_281,In_120);
or U668 (N_668,In_785,In_339);
nor U669 (N_669,In_1447,In_553);
xor U670 (N_670,In_493,In_354);
nor U671 (N_671,In_209,In_463);
xnor U672 (N_672,In_564,In_616);
or U673 (N_673,In_1316,In_1290);
or U674 (N_674,In_1061,In_906);
nand U675 (N_675,In_95,In_263);
or U676 (N_676,In_1051,In_1328);
nand U677 (N_677,In_977,In_856);
xnor U678 (N_678,In_504,In_527);
and U679 (N_679,In_380,In_893);
xnor U680 (N_680,In_657,In_530);
nand U681 (N_681,In_942,In_1474);
or U682 (N_682,In_1322,In_253);
nor U683 (N_683,In_123,In_775);
or U684 (N_684,In_1068,In_1416);
nand U685 (N_685,In_215,In_108);
or U686 (N_686,In_749,In_1221);
nor U687 (N_687,In_182,In_1019);
nand U688 (N_688,In_1442,In_1452);
nor U689 (N_689,In_768,In_444);
nand U690 (N_690,In_1487,In_754);
or U691 (N_691,In_126,In_524);
or U692 (N_692,In_594,In_78);
nand U693 (N_693,In_1269,In_952);
nor U694 (N_694,In_185,In_366);
nor U695 (N_695,In_1314,In_659);
nand U696 (N_696,In_1210,In_923);
and U697 (N_697,In_669,In_899);
nand U698 (N_698,In_1176,In_1010);
nor U699 (N_699,In_861,In_236);
nor U700 (N_700,In_1310,In_160);
or U701 (N_701,In_1402,In_431);
nor U702 (N_702,In_956,In_306);
nor U703 (N_703,In_1119,In_46);
and U704 (N_704,In_979,In_1237);
xor U705 (N_705,In_207,In_707);
nor U706 (N_706,In_104,In_1223);
and U707 (N_707,In_1053,In_805);
xor U708 (N_708,In_1016,In_931);
and U709 (N_709,In_827,In_724);
nor U710 (N_710,In_1375,In_477);
nor U711 (N_711,In_696,In_60);
nand U712 (N_712,In_1380,In_642);
nand U713 (N_713,In_725,In_595);
nor U714 (N_714,In_513,In_344);
nand U715 (N_715,In_577,In_914);
nand U716 (N_716,In_651,In_1196);
nor U717 (N_717,In_1400,In_128);
xnor U718 (N_718,In_1436,In_541);
and U719 (N_719,In_1200,In_1055);
or U720 (N_720,In_955,In_1220);
xnor U721 (N_721,In_1145,In_480);
xnor U722 (N_722,In_683,In_623);
or U723 (N_723,In_1430,In_106);
nor U724 (N_724,In_523,In_212);
nand U725 (N_725,In_619,In_850);
and U726 (N_726,In_96,In_1441);
nand U727 (N_727,In_628,In_360);
xnor U728 (N_728,In_1451,In_35);
and U729 (N_729,In_1240,In_909);
nand U730 (N_730,In_461,In_392);
nor U731 (N_731,In_820,In_298);
or U732 (N_732,In_1358,In_436);
or U733 (N_733,In_1304,In_799);
nor U734 (N_734,In_286,In_198);
xnor U735 (N_735,In_818,In_1023);
or U736 (N_736,In_816,In_7);
xor U737 (N_737,In_261,In_892);
or U738 (N_738,In_608,In_767);
nand U739 (N_739,In_729,In_39);
xor U740 (N_740,In_379,In_681);
xnor U741 (N_741,In_416,In_1477);
nand U742 (N_742,In_1450,In_134);
nand U743 (N_743,In_862,In_1192);
nand U744 (N_744,In_473,In_872);
nor U745 (N_745,In_427,In_1151);
and U746 (N_746,In_1434,In_658);
nand U747 (N_747,In_418,In_99);
or U748 (N_748,In_406,In_532);
or U749 (N_749,In_232,In_465);
and U750 (N_750,In_631,In_1077);
nor U751 (N_751,In_1338,In_157);
nor U752 (N_752,In_596,In_473);
xor U753 (N_753,In_13,In_1199);
and U754 (N_754,In_201,In_442);
xnor U755 (N_755,In_84,In_299);
and U756 (N_756,In_1495,In_315);
xnor U757 (N_757,In_832,In_899);
or U758 (N_758,In_1087,In_336);
nor U759 (N_759,In_588,In_1446);
and U760 (N_760,In_1330,In_763);
nand U761 (N_761,In_1112,In_937);
and U762 (N_762,In_1337,In_52);
nand U763 (N_763,In_911,In_561);
xor U764 (N_764,In_1264,In_299);
and U765 (N_765,In_618,In_51);
nor U766 (N_766,In_206,In_1369);
or U767 (N_767,In_645,In_1421);
nand U768 (N_768,In_501,In_1466);
nor U769 (N_769,In_1343,In_151);
and U770 (N_770,In_832,In_1304);
nand U771 (N_771,In_1225,In_433);
and U772 (N_772,In_1032,In_1405);
nand U773 (N_773,In_233,In_1228);
nor U774 (N_774,In_950,In_580);
nand U775 (N_775,In_233,In_1444);
nand U776 (N_776,In_1260,In_163);
or U777 (N_777,In_335,In_332);
or U778 (N_778,In_877,In_855);
nor U779 (N_779,In_1180,In_789);
and U780 (N_780,In_1267,In_708);
nand U781 (N_781,In_464,In_834);
and U782 (N_782,In_725,In_242);
and U783 (N_783,In_1475,In_1192);
nand U784 (N_784,In_1280,In_767);
xor U785 (N_785,In_1148,In_369);
xor U786 (N_786,In_53,In_616);
nand U787 (N_787,In_270,In_989);
and U788 (N_788,In_841,In_1494);
nand U789 (N_789,In_617,In_1104);
xnor U790 (N_790,In_624,In_1224);
nor U791 (N_791,In_82,In_1132);
or U792 (N_792,In_1088,In_218);
xnor U793 (N_793,In_1495,In_1034);
and U794 (N_794,In_1499,In_907);
xnor U795 (N_795,In_1360,In_1133);
nand U796 (N_796,In_96,In_411);
xor U797 (N_797,In_1468,In_87);
and U798 (N_798,In_640,In_859);
xnor U799 (N_799,In_888,In_503);
or U800 (N_800,In_195,In_530);
and U801 (N_801,In_213,In_644);
and U802 (N_802,In_40,In_1015);
nor U803 (N_803,In_327,In_844);
or U804 (N_804,In_1146,In_925);
nand U805 (N_805,In_584,In_1271);
nor U806 (N_806,In_1124,In_1084);
and U807 (N_807,In_1133,In_191);
or U808 (N_808,In_1212,In_977);
and U809 (N_809,In_1349,In_1226);
xor U810 (N_810,In_1037,In_1492);
xnor U811 (N_811,In_1101,In_789);
or U812 (N_812,In_1434,In_454);
nor U813 (N_813,In_1067,In_1123);
and U814 (N_814,In_860,In_1354);
xor U815 (N_815,In_230,In_662);
xnor U816 (N_816,In_379,In_945);
nor U817 (N_817,In_172,In_434);
xnor U818 (N_818,In_565,In_977);
or U819 (N_819,In_411,In_465);
xnor U820 (N_820,In_501,In_481);
and U821 (N_821,In_508,In_954);
xor U822 (N_822,In_1068,In_1490);
nand U823 (N_823,In_500,In_1320);
nor U824 (N_824,In_488,In_873);
nor U825 (N_825,In_1100,In_618);
nor U826 (N_826,In_528,In_876);
xnor U827 (N_827,In_598,In_308);
and U828 (N_828,In_743,In_103);
and U829 (N_829,In_84,In_1349);
xor U830 (N_830,In_987,In_788);
nand U831 (N_831,In_544,In_739);
xor U832 (N_832,In_515,In_1286);
xor U833 (N_833,In_83,In_1495);
or U834 (N_834,In_1402,In_510);
or U835 (N_835,In_537,In_997);
and U836 (N_836,In_1175,In_1287);
and U837 (N_837,In_1322,In_1223);
nor U838 (N_838,In_683,In_357);
nand U839 (N_839,In_984,In_1456);
and U840 (N_840,In_735,In_673);
nand U841 (N_841,In_689,In_1473);
nor U842 (N_842,In_284,In_294);
nand U843 (N_843,In_1184,In_754);
xor U844 (N_844,In_396,In_130);
and U845 (N_845,In_163,In_565);
xor U846 (N_846,In_429,In_109);
and U847 (N_847,In_437,In_1077);
and U848 (N_848,In_501,In_752);
nand U849 (N_849,In_699,In_405);
nand U850 (N_850,In_1185,In_1482);
nand U851 (N_851,In_13,In_1310);
xor U852 (N_852,In_67,In_347);
nor U853 (N_853,In_458,In_412);
nor U854 (N_854,In_970,In_911);
nor U855 (N_855,In_101,In_434);
xor U856 (N_856,In_1430,In_1088);
or U857 (N_857,In_1229,In_1131);
xnor U858 (N_858,In_1275,In_897);
nor U859 (N_859,In_110,In_104);
xor U860 (N_860,In_924,In_68);
or U861 (N_861,In_1118,In_500);
nor U862 (N_862,In_215,In_256);
nor U863 (N_863,In_1240,In_1052);
or U864 (N_864,In_274,In_742);
nor U865 (N_865,In_250,In_513);
nand U866 (N_866,In_4,In_325);
and U867 (N_867,In_1042,In_874);
and U868 (N_868,In_895,In_1080);
nor U869 (N_869,In_1293,In_1270);
nor U870 (N_870,In_232,In_1325);
and U871 (N_871,In_256,In_589);
and U872 (N_872,In_107,In_822);
xor U873 (N_873,In_1099,In_859);
and U874 (N_874,In_69,In_343);
nand U875 (N_875,In_374,In_468);
or U876 (N_876,In_870,In_1156);
xor U877 (N_877,In_1410,In_361);
xnor U878 (N_878,In_1102,In_1230);
xnor U879 (N_879,In_1349,In_1043);
and U880 (N_880,In_408,In_952);
or U881 (N_881,In_1194,In_670);
nand U882 (N_882,In_680,In_1403);
xor U883 (N_883,In_977,In_1033);
nor U884 (N_884,In_804,In_1486);
nand U885 (N_885,In_131,In_524);
nor U886 (N_886,In_1390,In_176);
or U887 (N_887,In_722,In_1048);
xnor U888 (N_888,In_1334,In_592);
and U889 (N_889,In_1479,In_1457);
nand U890 (N_890,In_968,In_842);
nand U891 (N_891,In_1286,In_1202);
nor U892 (N_892,In_682,In_1156);
nand U893 (N_893,In_1014,In_88);
or U894 (N_894,In_1439,In_1161);
xor U895 (N_895,In_695,In_943);
nor U896 (N_896,In_1305,In_185);
nand U897 (N_897,In_861,In_1168);
or U898 (N_898,In_1151,In_1281);
or U899 (N_899,In_1336,In_120);
nor U900 (N_900,In_1248,In_1279);
nor U901 (N_901,In_539,In_118);
nor U902 (N_902,In_1439,In_257);
xor U903 (N_903,In_1308,In_1490);
xor U904 (N_904,In_649,In_714);
and U905 (N_905,In_1148,In_1459);
and U906 (N_906,In_1481,In_520);
and U907 (N_907,In_747,In_932);
nor U908 (N_908,In_855,In_25);
nand U909 (N_909,In_738,In_463);
and U910 (N_910,In_7,In_633);
and U911 (N_911,In_274,In_811);
or U912 (N_912,In_1253,In_527);
and U913 (N_913,In_19,In_838);
or U914 (N_914,In_1413,In_1417);
or U915 (N_915,In_157,In_654);
or U916 (N_916,In_397,In_692);
nor U917 (N_917,In_372,In_72);
nor U918 (N_918,In_1401,In_518);
or U919 (N_919,In_720,In_943);
nand U920 (N_920,In_1434,In_361);
xor U921 (N_921,In_1021,In_1298);
or U922 (N_922,In_657,In_1284);
nor U923 (N_923,In_1381,In_9);
nor U924 (N_924,In_761,In_1425);
and U925 (N_925,In_57,In_1158);
xnor U926 (N_926,In_260,In_236);
nand U927 (N_927,In_39,In_423);
xnor U928 (N_928,In_1354,In_344);
xnor U929 (N_929,In_1388,In_841);
xnor U930 (N_930,In_1236,In_523);
or U931 (N_931,In_510,In_1456);
nor U932 (N_932,In_1048,In_1056);
and U933 (N_933,In_997,In_1264);
nand U934 (N_934,In_1040,In_1165);
xnor U935 (N_935,In_308,In_260);
xnor U936 (N_936,In_17,In_1116);
nand U937 (N_937,In_199,In_985);
nand U938 (N_938,In_957,In_295);
nand U939 (N_939,In_644,In_276);
nand U940 (N_940,In_955,In_1493);
and U941 (N_941,In_1097,In_504);
nor U942 (N_942,In_1294,In_470);
and U943 (N_943,In_841,In_1225);
xnor U944 (N_944,In_1353,In_699);
and U945 (N_945,In_221,In_1142);
nor U946 (N_946,In_609,In_1052);
or U947 (N_947,In_419,In_568);
nand U948 (N_948,In_1369,In_907);
or U949 (N_949,In_193,In_108);
xnor U950 (N_950,In_1180,In_827);
nor U951 (N_951,In_1070,In_190);
nor U952 (N_952,In_886,In_114);
xor U953 (N_953,In_348,In_773);
nor U954 (N_954,In_954,In_1264);
xor U955 (N_955,In_244,In_892);
or U956 (N_956,In_819,In_1090);
nor U957 (N_957,In_357,In_304);
or U958 (N_958,In_928,In_725);
or U959 (N_959,In_262,In_1362);
xor U960 (N_960,In_956,In_871);
xnor U961 (N_961,In_1052,In_1492);
xnor U962 (N_962,In_1351,In_985);
xor U963 (N_963,In_497,In_1273);
nand U964 (N_964,In_916,In_261);
nand U965 (N_965,In_453,In_332);
and U966 (N_966,In_599,In_1230);
nand U967 (N_967,In_746,In_260);
or U968 (N_968,In_254,In_266);
and U969 (N_969,In_522,In_279);
xor U970 (N_970,In_1173,In_946);
nor U971 (N_971,In_1322,In_578);
nand U972 (N_972,In_553,In_251);
or U973 (N_973,In_580,In_1316);
nor U974 (N_974,In_666,In_588);
and U975 (N_975,In_1317,In_131);
xor U976 (N_976,In_613,In_136);
nand U977 (N_977,In_706,In_916);
nand U978 (N_978,In_117,In_531);
or U979 (N_979,In_996,In_935);
or U980 (N_980,In_519,In_1396);
or U981 (N_981,In_1271,In_1077);
xor U982 (N_982,In_935,In_553);
nand U983 (N_983,In_1231,In_169);
nand U984 (N_984,In_78,In_81);
nor U985 (N_985,In_311,In_744);
and U986 (N_986,In_623,In_810);
and U987 (N_987,In_1035,In_829);
or U988 (N_988,In_736,In_20);
or U989 (N_989,In_194,In_1356);
nand U990 (N_990,In_1279,In_550);
nand U991 (N_991,In_1209,In_842);
or U992 (N_992,In_209,In_995);
nand U993 (N_993,In_356,In_1061);
nor U994 (N_994,In_617,In_148);
or U995 (N_995,In_666,In_962);
or U996 (N_996,In_930,In_1409);
nor U997 (N_997,In_1455,In_456);
nand U998 (N_998,In_1302,In_1070);
xnor U999 (N_999,In_1151,In_537);
and U1000 (N_1000,In_187,In_623);
or U1001 (N_1001,In_1021,In_1153);
nor U1002 (N_1002,In_382,In_136);
and U1003 (N_1003,In_406,In_40);
xor U1004 (N_1004,In_1029,In_175);
xnor U1005 (N_1005,In_193,In_1316);
or U1006 (N_1006,In_1282,In_654);
nand U1007 (N_1007,In_714,In_735);
nand U1008 (N_1008,In_537,In_905);
and U1009 (N_1009,In_926,In_726);
xor U1010 (N_1010,In_12,In_281);
nand U1011 (N_1011,In_995,In_910);
and U1012 (N_1012,In_1158,In_852);
nor U1013 (N_1013,In_781,In_780);
and U1014 (N_1014,In_894,In_1261);
xnor U1015 (N_1015,In_817,In_1394);
xnor U1016 (N_1016,In_124,In_151);
and U1017 (N_1017,In_127,In_842);
and U1018 (N_1018,In_1200,In_987);
and U1019 (N_1019,In_885,In_1189);
nand U1020 (N_1020,In_601,In_941);
xnor U1021 (N_1021,In_86,In_614);
or U1022 (N_1022,In_418,In_1318);
and U1023 (N_1023,In_181,In_885);
and U1024 (N_1024,In_293,In_847);
xor U1025 (N_1025,In_277,In_1087);
nor U1026 (N_1026,In_1094,In_74);
and U1027 (N_1027,In_708,In_883);
xnor U1028 (N_1028,In_154,In_299);
nand U1029 (N_1029,In_1175,In_164);
nand U1030 (N_1030,In_570,In_1396);
xnor U1031 (N_1031,In_571,In_481);
nand U1032 (N_1032,In_898,In_739);
or U1033 (N_1033,In_749,In_579);
nor U1034 (N_1034,In_1253,In_875);
and U1035 (N_1035,In_301,In_1131);
or U1036 (N_1036,In_720,In_85);
and U1037 (N_1037,In_904,In_1388);
nor U1038 (N_1038,In_543,In_1020);
and U1039 (N_1039,In_1090,In_1038);
and U1040 (N_1040,In_293,In_472);
nor U1041 (N_1041,In_1497,In_1155);
nand U1042 (N_1042,In_130,In_1031);
nand U1043 (N_1043,In_556,In_1392);
nor U1044 (N_1044,In_1011,In_10);
xnor U1045 (N_1045,In_352,In_1275);
and U1046 (N_1046,In_977,In_119);
nor U1047 (N_1047,In_894,In_747);
nand U1048 (N_1048,In_928,In_918);
and U1049 (N_1049,In_627,In_1090);
and U1050 (N_1050,In_963,In_1150);
xnor U1051 (N_1051,In_649,In_192);
nand U1052 (N_1052,In_791,In_140);
nand U1053 (N_1053,In_101,In_1165);
xnor U1054 (N_1054,In_1101,In_910);
and U1055 (N_1055,In_1366,In_460);
nor U1056 (N_1056,In_166,In_277);
or U1057 (N_1057,In_362,In_150);
and U1058 (N_1058,In_264,In_424);
xnor U1059 (N_1059,In_325,In_456);
xnor U1060 (N_1060,In_198,In_1331);
xor U1061 (N_1061,In_173,In_431);
nand U1062 (N_1062,In_1440,In_303);
nor U1063 (N_1063,In_1351,In_741);
or U1064 (N_1064,In_162,In_1345);
nor U1065 (N_1065,In_455,In_761);
xnor U1066 (N_1066,In_1021,In_309);
or U1067 (N_1067,In_1017,In_625);
or U1068 (N_1068,In_963,In_1130);
xnor U1069 (N_1069,In_333,In_708);
nor U1070 (N_1070,In_495,In_1401);
xor U1071 (N_1071,In_1479,In_155);
nand U1072 (N_1072,In_426,In_1489);
or U1073 (N_1073,In_1149,In_1006);
xnor U1074 (N_1074,In_71,In_190);
and U1075 (N_1075,In_994,In_495);
nor U1076 (N_1076,In_46,In_987);
nand U1077 (N_1077,In_848,In_1437);
nor U1078 (N_1078,In_1392,In_1191);
xor U1079 (N_1079,In_109,In_1119);
nand U1080 (N_1080,In_481,In_1291);
or U1081 (N_1081,In_503,In_302);
nand U1082 (N_1082,In_1236,In_1487);
nor U1083 (N_1083,In_1399,In_1404);
xnor U1084 (N_1084,In_466,In_272);
nand U1085 (N_1085,In_341,In_762);
xor U1086 (N_1086,In_1465,In_1164);
nand U1087 (N_1087,In_42,In_1378);
and U1088 (N_1088,In_1461,In_893);
nand U1089 (N_1089,In_1054,In_297);
nand U1090 (N_1090,In_819,In_563);
nor U1091 (N_1091,In_816,In_574);
and U1092 (N_1092,In_632,In_1312);
nand U1093 (N_1093,In_818,In_205);
and U1094 (N_1094,In_1309,In_1222);
nor U1095 (N_1095,In_1285,In_694);
nand U1096 (N_1096,In_1122,In_968);
or U1097 (N_1097,In_1158,In_439);
and U1098 (N_1098,In_565,In_1295);
xnor U1099 (N_1099,In_923,In_1020);
or U1100 (N_1100,In_383,In_1001);
nor U1101 (N_1101,In_1332,In_499);
nor U1102 (N_1102,In_910,In_1265);
and U1103 (N_1103,In_579,In_1309);
nor U1104 (N_1104,In_251,In_823);
and U1105 (N_1105,In_483,In_921);
or U1106 (N_1106,In_886,In_1163);
or U1107 (N_1107,In_1160,In_364);
nor U1108 (N_1108,In_1361,In_896);
and U1109 (N_1109,In_764,In_952);
nor U1110 (N_1110,In_290,In_160);
and U1111 (N_1111,In_1062,In_421);
or U1112 (N_1112,In_1240,In_352);
nor U1113 (N_1113,In_1050,In_966);
or U1114 (N_1114,In_273,In_1110);
and U1115 (N_1115,In_870,In_900);
and U1116 (N_1116,In_1036,In_685);
xor U1117 (N_1117,In_916,In_1240);
nor U1118 (N_1118,In_333,In_1274);
xnor U1119 (N_1119,In_194,In_926);
nor U1120 (N_1120,In_1101,In_510);
and U1121 (N_1121,In_934,In_1035);
or U1122 (N_1122,In_1080,In_476);
nor U1123 (N_1123,In_1052,In_895);
xnor U1124 (N_1124,In_1410,In_818);
nand U1125 (N_1125,In_1489,In_733);
and U1126 (N_1126,In_1014,In_1042);
and U1127 (N_1127,In_136,In_1197);
nand U1128 (N_1128,In_831,In_1150);
nand U1129 (N_1129,In_611,In_953);
or U1130 (N_1130,In_263,In_1069);
and U1131 (N_1131,In_435,In_1286);
nand U1132 (N_1132,In_1300,In_1366);
xnor U1133 (N_1133,In_511,In_353);
nor U1134 (N_1134,In_1292,In_1498);
and U1135 (N_1135,In_1025,In_677);
nand U1136 (N_1136,In_457,In_1376);
xnor U1137 (N_1137,In_582,In_1035);
nand U1138 (N_1138,In_741,In_862);
and U1139 (N_1139,In_1061,In_661);
or U1140 (N_1140,In_416,In_1156);
and U1141 (N_1141,In_838,In_1120);
nor U1142 (N_1142,In_1357,In_366);
xnor U1143 (N_1143,In_373,In_1384);
nor U1144 (N_1144,In_671,In_788);
nor U1145 (N_1145,In_1459,In_388);
xor U1146 (N_1146,In_1477,In_663);
nor U1147 (N_1147,In_572,In_1401);
nand U1148 (N_1148,In_226,In_1118);
nand U1149 (N_1149,In_1387,In_17);
nor U1150 (N_1150,In_330,In_970);
xnor U1151 (N_1151,In_612,In_999);
nor U1152 (N_1152,In_901,In_1261);
and U1153 (N_1153,In_377,In_1029);
xor U1154 (N_1154,In_917,In_395);
nand U1155 (N_1155,In_1212,In_406);
nor U1156 (N_1156,In_44,In_1214);
or U1157 (N_1157,In_605,In_384);
and U1158 (N_1158,In_1095,In_270);
xnor U1159 (N_1159,In_1442,In_378);
or U1160 (N_1160,In_483,In_1082);
nor U1161 (N_1161,In_486,In_134);
or U1162 (N_1162,In_970,In_985);
or U1163 (N_1163,In_138,In_724);
and U1164 (N_1164,In_322,In_399);
nor U1165 (N_1165,In_1210,In_73);
or U1166 (N_1166,In_743,In_910);
or U1167 (N_1167,In_516,In_286);
or U1168 (N_1168,In_173,In_669);
and U1169 (N_1169,In_1486,In_395);
nand U1170 (N_1170,In_849,In_614);
nor U1171 (N_1171,In_1479,In_434);
nor U1172 (N_1172,In_327,In_692);
xor U1173 (N_1173,In_840,In_204);
or U1174 (N_1174,In_1476,In_448);
nand U1175 (N_1175,In_442,In_1063);
nand U1176 (N_1176,In_1419,In_219);
nand U1177 (N_1177,In_1106,In_427);
and U1178 (N_1178,In_5,In_1373);
nor U1179 (N_1179,In_1339,In_816);
and U1180 (N_1180,In_331,In_619);
and U1181 (N_1181,In_746,In_809);
nand U1182 (N_1182,In_494,In_412);
xnor U1183 (N_1183,In_1238,In_1225);
or U1184 (N_1184,In_246,In_1424);
nand U1185 (N_1185,In_727,In_1383);
xnor U1186 (N_1186,In_209,In_90);
or U1187 (N_1187,In_47,In_1295);
nand U1188 (N_1188,In_13,In_334);
nor U1189 (N_1189,In_1364,In_849);
nand U1190 (N_1190,In_493,In_903);
nand U1191 (N_1191,In_842,In_338);
or U1192 (N_1192,In_412,In_159);
and U1193 (N_1193,In_69,In_1366);
or U1194 (N_1194,In_956,In_1377);
nand U1195 (N_1195,In_716,In_280);
nand U1196 (N_1196,In_787,In_955);
or U1197 (N_1197,In_806,In_1182);
nor U1198 (N_1198,In_625,In_334);
nor U1199 (N_1199,In_1323,In_1418);
or U1200 (N_1200,In_381,In_13);
or U1201 (N_1201,In_1316,In_332);
xnor U1202 (N_1202,In_1484,In_1055);
nor U1203 (N_1203,In_1134,In_876);
xor U1204 (N_1204,In_1288,In_1021);
nand U1205 (N_1205,In_1408,In_1092);
or U1206 (N_1206,In_264,In_965);
nand U1207 (N_1207,In_1133,In_226);
and U1208 (N_1208,In_384,In_1109);
and U1209 (N_1209,In_1390,In_253);
nand U1210 (N_1210,In_525,In_839);
nand U1211 (N_1211,In_1202,In_1278);
nand U1212 (N_1212,In_1364,In_489);
and U1213 (N_1213,In_1243,In_801);
nand U1214 (N_1214,In_349,In_1427);
nor U1215 (N_1215,In_476,In_1114);
and U1216 (N_1216,In_706,In_276);
nand U1217 (N_1217,In_345,In_658);
xnor U1218 (N_1218,In_1312,In_943);
or U1219 (N_1219,In_1118,In_1262);
xnor U1220 (N_1220,In_929,In_1270);
and U1221 (N_1221,In_618,In_650);
nor U1222 (N_1222,In_933,In_808);
nor U1223 (N_1223,In_1269,In_546);
nor U1224 (N_1224,In_1277,In_1341);
or U1225 (N_1225,In_727,In_35);
and U1226 (N_1226,In_351,In_593);
or U1227 (N_1227,In_1154,In_580);
and U1228 (N_1228,In_133,In_600);
nand U1229 (N_1229,In_467,In_786);
nand U1230 (N_1230,In_978,In_1397);
nand U1231 (N_1231,In_58,In_983);
nor U1232 (N_1232,In_1303,In_140);
nor U1233 (N_1233,In_1490,In_1043);
nand U1234 (N_1234,In_803,In_330);
nand U1235 (N_1235,In_1178,In_1327);
xor U1236 (N_1236,In_21,In_250);
nand U1237 (N_1237,In_1284,In_814);
nor U1238 (N_1238,In_1450,In_230);
xnor U1239 (N_1239,In_1079,In_1360);
nand U1240 (N_1240,In_716,In_759);
and U1241 (N_1241,In_302,In_358);
nor U1242 (N_1242,In_54,In_611);
nor U1243 (N_1243,In_955,In_1060);
or U1244 (N_1244,In_1448,In_1119);
or U1245 (N_1245,In_1197,In_662);
xor U1246 (N_1246,In_223,In_863);
xnor U1247 (N_1247,In_412,In_605);
or U1248 (N_1248,In_572,In_486);
and U1249 (N_1249,In_1466,In_370);
nor U1250 (N_1250,In_242,In_944);
xnor U1251 (N_1251,In_46,In_1437);
and U1252 (N_1252,In_882,In_1434);
or U1253 (N_1253,In_655,In_1023);
and U1254 (N_1254,In_780,In_130);
or U1255 (N_1255,In_428,In_914);
nand U1256 (N_1256,In_1233,In_753);
and U1257 (N_1257,In_4,In_384);
or U1258 (N_1258,In_939,In_1163);
xor U1259 (N_1259,In_478,In_587);
and U1260 (N_1260,In_639,In_638);
and U1261 (N_1261,In_499,In_69);
and U1262 (N_1262,In_868,In_1363);
nor U1263 (N_1263,In_545,In_1070);
nand U1264 (N_1264,In_833,In_451);
and U1265 (N_1265,In_1246,In_1378);
nor U1266 (N_1266,In_705,In_1239);
and U1267 (N_1267,In_43,In_1039);
xor U1268 (N_1268,In_1191,In_781);
nand U1269 (N_1269,In_231,In_259);
xor U1270 (N_1270,In_1213,In_520);
nand U1271 (N_1271,In_578,In_436);
and U1272 (N_1272,In_640,In_1363);
and U1273 (N_1273,In_1168,In_545);
nand U1274 (N_1274,In_539,In_1427);
nand U1275 (N_1275,In_1211,In_1443);
and U1276 (N_1276,In_693,In_344);
nand U1277 (N_1277,In_807,In_1320);
nand U1278 (N_1278,In_344,In_1011);
xor U1279 (N_1279,In_631,In_230);
or U1280 (N_1280,In_961,In_467);
nand U1281 (N_1281,In_12,In_1343);
or U1282 (N_1282,In_864,In_911);
nor U1283 (N_1283,In_735,In_1121);
or U1284 (N_1284,In_80,In_91);
and U1285 (N_1285,In_1371,In_1088);
or U1286 (N_1286,In_1342,In_587);
nor U1287 (N_1287,In_110,In_218);
xnor U1288 (N_1288,In_81,In_1412);
nor U1289 (N_1289,In_370,In_302);
or U1290 (N_1290,In_797,In_909);
xnor U1291 (N_1291,In_964,In_248);
and U1292 (N_1292,In_1008,In_248);
nand U1293 (N_1293,In_1403,In_630);
or U1294 (N_1294,In_399,In_1144);
or U1295 (N_1295,In_1172,In_1418);
nand U1296 (N_1296,In_1286,In_191);
or U1297 (N_1297,In_1107,In_260);
or U1298 (N_1298,In_1233,In_691);
nand U1299 (N_1299,In_1111,In_768);
or U1300 (N_1300,In_683,In_1335);
or U1301 (N_1301,In_1175,In_394);
and U1302 (N_1302,In_1218,In_291);
nand U1303 (N_1303,In_465,In_1032);
nand U1304 (N_1304,In_617,In_72);
nand U1305 (N_1305,In_606,In_1405);
or U1306 (N_1306,In_1286,In_1101);
xor U1307 (N_1307,In_1060,In_1355);
nand U1308 (N_1308,In_2,In_1017);
nor U1309 (N_1309,In_116,In_1441);
xor U1310 (N_1310,In_1056,In_387);
nand U1311 (N_1311,In_1431,In_218);
nand U1312 (N_1312,In_443,In_1010);
nand U1313 (N_1313,In_474,In_1294);
or U1314 (N_1314,In_918,In_947);
nor U1315 (N_1315,In_1389,In_617);
nor U1316 (N_1316,In_1397,In_711);
or U1317 (N_1317,In_440,In_509);
or U1318 (N_1318,In_1082,In_1481);
nor U1319 (N_1319,In_80,In_613);
xnor U1320 (N_1320,In_165,In_784);
nand U1321 (N_1321,In_108,In_727);
or U1322 (N_1322,In_726,In_1469);
nand U1323 (N_1323,In_326,In_67);
and U1324 (N_1324,In_427,In_112);
nor U1325 (N_1325,In_331,In_1007);
nor U1326 (N_1326,In_231,In_1358);
or U1327 (N_1327,In_984,In_766);
nand U1328 (N_1328,In_671,In_549);
or U1329 (N_1329,In_1393,In_658);
xnor U1330 (N_1330,In_1203,In_1192);
nand U1331 (N_1331,In_908,In_1060);
xor U1332 (N_1332,In_1018,In_599);
or U1333 (N_1333,In_986,In_1015);
and U1334 (N_1334,In_161,In_822);
and U1335 (N_1335,In_821,In_387);
or U1336 (N_1336,In_625,In_1254);
nand U1337 (N_1337,In_1087,In_36);
xnor U1338 (N_1338,In_1015,In_137);
xor U1339 (N_1339,In_1404,In_219);
xnor U1340 (N_1340,In_25,In_997);
and U1341 (N_1341,In_1075,In_121);
nor U1342 (N_1342,In_152,In_1060);
nor U1343 (N_1343,In_205,In_765);
nor U1344 (N_1344,In_1300,In_786);
and U1345 (N_1345,In_371,In_1394);
nand U1346 (N_1346,In_105,In_1465);
nand U1347 (N_1347,In_344,In_749);
nand U1348 (N_1348,In_823,In_1219);
or U1349 (N_1349,In_718,In_582);
or U1350 (N_1350,In_693,In_411);
xor U1351 (N_1351,In_581,In_553);
or U1352 (N_1352,In_859,In_1093);
nand U1353 (N_1353,In_610,In_574);
nor U1354 (N_1354,In_60,In_717);
xor U1355 (N_1355,In_186,In_99);
nor U1356 (N_1356,In_1204,In_1181);
or U1357 (N_1357,In_1133,In_243);
or U1358 (N_1358,In_341,In_1469);
xnor U1359 (N_1359,In_224,In_1046);
xnor U1360 (N_1360,In_231,In_577);
nor U1361 (N_1361,In_825,In_160);
and U1362 (N_1362,In_483,In_268);
xor U1363 (N_1363,In_1057,In_1432);
or U1364 (N_1364,In_1382,In_1003);
nand U1365 (N_1365,In_515,In_1070);
and U1366 (N_1366,In_246,In_491);
xnor U1367 (N_1367,In_886,In_1197);
nand U1368 (N_1368,In_1075,In_1148);
nor U1369 (N_1369,In_1180,In_972);
nor U1370 (N_1370,In_228,In_1361);
and U1371 (N_1371,In_1,In_59);
and U1372 (N_1372,In_446,In_609);
xor U1373 (N_1373,In_552,In_5);
nand U1374 (N_1374,In_1490,In_1145);
or U1375 (N_1375,In_396,In_362);
xnor U1376 (N_1376,In_641,In_306);
and U1377 (N_1377,In_1191,In_1240);
nand U1378 (N_1378,In_659,In_1426);
nand U1379 (N_1379,In_1475,In_1217);
nor U1380 (N_1380,In_373,In_826);
or U1381 (N_1381,In_1354,In_1428);
nand U1382 (N_1382,In_399,In_23);
nor U1383 (N_1383,In_918,In_1148);
xor U1384 (N_1384,In_1330,In_550);
nor U1385 (N_1385,In_359,In_518);
or U1386 (N_1386,In_1175,In_130);
nand U1387 (N_1387,In_1460,In_521);
nor U1388 (N_1388,In_163,In_1176);
nand U1389 (N_1389,In_287,In_694);
nand U1390 (N_1390,In_137,In_1072);
and U1391 (N_1391,In_1468,In_1313);
xnor U1392 (N_1392,In_1119,In_1098);
nand U1393 (N_1393,In_10,In_528);
nand U1394 (N_1394,In_5,In_794);
nand U1395 (N_1395,In_717,In_639);
nor U1396 (N_1396,In_169,In_183);
or U1397 (N_1397,In_977,In_1020);
nor U1398 (N_1398,In_645,In_1104);
or U1399 (N_1399,In_264,In_683);
xnor U1400 (N_1400,In_304,In_385);
and U1401 (N_1401,In_1181,In_739);
xnor U1402 (N_1402,In_443,In_375);
nand U1403 (N_1403,In_718,In_1273);
nor U1404 (N_1404,In_32,In_1209);
and U1405 (N_1405,In_375,In_126);
nand U1406 (N_1406,In_1011,In_692);
nor U1407 (N_1407,In_1299,In_387);
or U1408 (N_1408,In_977,In_712);
xnor U1409 (N_1409,In_445,In_371);
and U1410 (N_1410,In_1369,In_57);
nand U1411 (N_1411,In_1214,In_894);
nor U1412 (N_1412,In_1196,In_367);
nand U1413 (N_1413,In_141,In_972);
xnor U1414 (N_1414,In_941,In_423);
nand U1415 (N_1415,In_553,In_812);
nor U1416 (N_1416,In_1428,In_1424);
or U1417 (N_1417,In_1070,In_1447);
nor U1418 (N_1418,In_1183,In_602);
nand U1419 (N_1419,In_997,In_787);
nand U1420 (N_1420,In_540,In_1282);
and U1421 (N_1421,In_967,In_71);
nor U1422 (N_1422,In_156,In_786);
or U1423 (N_1423,In_1332,In_1317);
and U1424 (N_1424,In_1048,In_1141);
and U1425 (N_1425,In_291,In_1316);
and U1426 (N_1426,In_858,In_1065);
xnor U1427 (N_1427,In_221,In_998);
or U1428 (N_1428,In_994,In_1012);
nand U1429 (N_1429,In_283,In_347);
or U1430 (N_1430,In_1231,In_232);
or U1431 (N_1431,In_1023,In_806);
nand U1432 (N_1432,In_704,In_1286);
xnor U1433 (N_1433,In_1154,In_1343);
or U1434 (N_1434,In_1455,In_706);
nand U1435 (N_1435,In_413,In_848);
nor U1436 (N_1436,In_406,In_1400);
nand U1437 (N_1437,In_1021,In_134);
xor U1438 (N_1438,In_976,In_15);
nor U1439 (N_1439,In_447,In_915);
nand U1440 (N_1440,In_1161,In_578);
nand U1441 (N_1441,In_73,In_158);
or U1442 (N_1442,In_1477,In_686);
or U1443 (N_1443,In_397,In_151);
or U1444 (N_1444,In_580,In_1203);
xor U1445 (N_1445,In_986,In_430);
or U1446 (N_1446,In_835,In_1088);
and U1447 (N_1447,In_570,In_1248);
and U1448 (N_1448,In_418,In_681);
xnor U1449 (N_1449,In_1152,In_104);
nand U1450 (N_1450,In_746,In_1475);
or U1451 (N_1451,In_494,In_194);
nand U1452 (N_1452,In_944,In_1114);
and U1453 (N_1453,In_820,In_1155);
and U1454 (N_1454,In_501,In_160);
nand U1455 (N_1455,In_861,In_381);
nand U1456 (N_1456,In_1066,In_860);
or U1457 (N_1457,In_504,In_1286);
xor U1458 (N_1458,In_236,In_1355);
nor U1459 (N_1459,In_674,In_1458);
and U1460 (N_1460,In_892,In_458);
nor U1461 (N_1461,In_912,In_1251);
nor U1462 (N_1462,In_247,In_666);
or U1463 (N_1463,In_1336,In_960);
or U1464 (N_1464,In_202,In_989);
and U1465 (N_1465,In_569,In_991);
and U1466 (N_1466,In_286,In_688);
and U1467 (N_1467,In_1449,In_1308);
xor U1468 (N_1468,In_920,In_648);
nor U1469 (N_1469,In_1050,In_146);
nor U1470 (N_1470,In_432,In_752);
nand U1471 (N_1471,In_786,In_937);
nand U1472 (N_1472,In_1248,In_198);
nand U1473 (N_1473,In_523,In_454);
nand U1474 (N_1474,In_1086,In_1178);
xor U1475 (N_1475,In_1173,In_1409);
or U1476 (N_1476,In_1200,In_171);
xor U1477 (N_1477,In_159,In_1397);
nor U1478 (N_1478,In_605,In_1268);
and U1479 (N_1479,In_1341,In_704);
nor U1480 (N_1480,In_800,In_264);
or U1481 (N_1481,In_1231,In_1414);
nor U1482 (N_1482,In_835,In_299);
nor U1483 (N_1483,In_452,In_665);
nor U1484 (N_1484,In_459,In_377);
xor U1485 (N_1485,In_949,In_283);
and U1486 (N_1486,In_502,In_45);
and U1487 (N_1487,In_398,In_535);
nand U1488 (N_1488,In_1264,In_1398);
nand U1489 (N_1489,In_201,In_502);
or U1490 (N_1490,In_439,In_528);
xnor U1491 (N_1491,In_341,In_922);
and U1492 (N_1492,In_775,In_1372);
nor U1493 (N_1493,In_1463,In_792);
and U1494 (N_1494,In_1195,In_388);
xnor U1495 (N_1495,In_291,In_961);
xor U1496 (N_1496,In_38,In_1363);
xor U1497 (N_1497,In_1072,In_427);
and U1498 (N_1498,In_1032,In_627);
and U1499 (N_1499,In_853,In_116);
and U1500 (N_1500,In_278,In_214);
nor U1501 (N_1501,In_279,In_1479);
nand U1502 (N_1502,In_655,In_1483);
and U1503 (N_1503,In_860,In_123);
nand U1504 (N_1504,In_926,In_847);
xnor U1505 (N_1505,In_52,In_729);
and U1506 (N_1506,In_118,In_913);
xnor U1507 (N_1507,In_514,In_336);
or U1508 (N_1508,In_341,In_236);
or U1509 (N_1509,In_602,In_516);
nand U1510 (N_1510,In_1464,In_528);
and U1511 (N_1511,In_1218,In_259);
and U1512 (N_1512,In_1389,In_1142);
nand U1513 (N_1513,In_611,In_1190);
or U1514 (N_1514,In_1285,In_22);
xor U1515 (N_1515,In_457,In_202);
and U1516 (N_1516,In_574,In_1447);
xnor U1517 (N_1517,In_1268,In_584);
nor U1518 (N_1518,In_339,In_984);
nand U1519 (N_1519,In_631,In_860);
or U1520 (N_1520,In_1378,In_821);
nor U1521 (N_1521,In_737,In_971);
nand U1522 (N_1522,In_607,In_1444);
xor U1523 (N_1523,In_1482,In_629);
xnor U1524 (N_1524,In_388,In_1131);
xnor U1525 (N_1525,In_1348,In_1295);
or U1526 (N_1526,In_1467,In_900);
or U1527 (N_1527,In_1298,In_803);
nor U1528 (N_1528,In_621,In_1138);
xnor U1529 (N_1529,In_1377,In_1025);
or U1530 (N_1530,In_765,In_410);
and U1531 (N_1531,In_210,In_1129);
nor U1532 (N_1532,In_904,In_811);
nor U1533 (N_1533,In_7,In_275);
nand U1534 (N_1534,In_1447,In_658);
or U1535 (N_1535,In_1275,In_1073);
nand U1536 (N_1536,In_1016,In_1138);
and U1537 (N_1537,In_330,In_943);
or U1538 (N_1538,In_814,In_1381);
xnor U1539 (N_1539,In_1210,In_1385);
nor U1540 (N_1540,In_765,In_1294);
xnor U1541 (N_1541,In_1426,In_923);
xor U1542 (N_1542,In_572,In_624);
nand U1543 (N_1543,In_570,In_771);
nor U1544 (N_1544,In_21,In_691);
and U1545 (N_1545,In_766,In_1424);
or U1546 (N_1546,In_1112,In_1199);
and U1547 (N_1547,In_388,In_503);
xnor U1548 (N_1548,In_1420,In_749);
nand U1549 (N_1549,In_740,In_306);
nor U1550 (N_1550,In_1375,In_411);
and U1551 (N_1551,In_73,In_1415);
and U1552 (N_1552,In_1079,In_768);
nor U1553 (N_1553,In_1488,In_234);
nand U1554 (N_1554,In_502,In_13);
nor U1555 (N_1555,In_629,In_1080);
or U1556 (N_1556,In_623,In_1387);
xor U1557 (N_1557,In_1179,In_266);
or U1558 (N_1558,In_427,In_1232);
nor U1559 (N_1559,In_1307,In_1390);
nor U1560 (N_1560,In_304,In_746);
and U1561 (N_1561,In_835,In_1118);
xnor U1562 (N_1562,In_695,In_38);
nand U1563 (N_1563,In_244,In_1017);
nor U1564 (N_1564,In_46,In_1456);
and U1565 (N_1565,In_826,In_1284);
nand U1566 (N_1566,In_828,In_1216);
nor U1567 (N_1567,In_115,In_199);
and U1568 (N_1568,In_759,In_802);
or U1569 (N_1569,In_1410,In_625);
and U1570 (N_1570,In_339,In_1238);
or U1571 (N_1571,In_662,In_890);
xnor U1572 (N_1572,In_653,In_773);
nand U1573 (N_1573,In_991,In_332);
or U1574 (N_1574,In_1203,In_1153);
and U1575 (N_1575,In_258,In_1199);
nor U1576 (N_1576,In_488,In_368);
or U1577 (N_1577,In_456,In_793);
and U1578 (N_1578,In_7,In_711);
nand U1579 (N_1579,In_487,In_1459);
nand U1580 (N_1580,In_397,In_773);
nand U1581 (N_1581,In_65,In_146);
or U1582 (N_1582,In_1356,In_500);
nor U1583 (N_1583,In_899,In_1272);
xor U1584 (N_1584,In_915,In_1200);
and U1585 (N_1585,In_494,In_391);
xor U1586 (N_1586,In_1197,In_46);
nand U1587 (N_1587,In_811,In_97);
nor U1588 (N_1588,In_1118,In_2);
and U1589 (N_1589,In_1392,In_1091);
nand U1590 (N_1590,In_814,In_1081);
or U1591 (N_1591,In_1024,In_857);
nor U1592 (N_1592,In_1172,In_1142);
or U1593 (N_1593,In_506,In_1480);
or U1594 (N_1594,In_744,In_1028);
nand U1595 (N_1595,In_1134,In_1257);
nand U1596 (N_1596,In_554,In_236);
xor U1597 (N_1597,In_1144,In_1130);
nor U1598 (N_1598,In_1241,In_1207);
nand U1599 (N_1599,In_88,In_1229);
and U1600 (N_1600,In_616,In_433);
xnor U1601 (N_1601,In_37,In_823);
nand U1602 (N_1602,In_4,In_1411);
xnor U1603 (N_1603,In_1379,In_309);
nand U1604 (N_1604,In_337,In_576);
nand U1605 (N_1605,In_919,In_646);
xor U1606 (N_1606,In_46,In_1109);
and U1607 (N_1607,In_1225,In_1412);
nand U1608 (N_1608,In_586,In_821);
xnor U1609 (N_1609,In_614,In_710);
xnor U1610 (N_1610,In_797,In_1009);
or U1611 (N_1611,In_874,In_607);
nor U1612 (N_1612,In_111,In_882);
xor U1613 (N_1613,In_1048,In_861);
nor U1614 (N_1614,In_930,In_1262);
nor U1615 (N_1615,In_1037,In_47);
xnor U1616 (N_1616,In_707,In_981);
and U1617 (N_1617,In_1471,In_807);
and U1618 (N_1618,In_1447,In_721);
nand U1619 (N_1619,In_235,In_1193);
xor U1620 (N_1620,In_1007,In_1179);
nand U1621 (N_1621,In_313,In_1267);
nor U1622 (N_1622,In_80,In_54);
nand U1623 (N_1623,In_1065,In_703);
or U1624 (N_1624,In_270,In_929);
nand U1625 (N_1625,In_1288,In_315);
or U1626 (N_1626,In_249,In_827);
xnor U1627 (N_1627,In_119,In_24);
xor U1628 (N_1628,In_87,In_760);
nand U1629 (N_1629,In_955,In_1485);
xnor U1630 (N_1630,In_1168,In_225);
and U1631 (N_1631,In_72,In_50);
nand U1632 (N_1632,In_461,In_604);
or U1633 (N_1633,In_1398,In_542);
nor U1634 (N_1634,In_1477,In_816);
and U1635 (N_1635,In_914,In_1389);
or U1636 (N_1636,In_1211,In_573);
and U1637 (N_1637,In_739,In_482);
xor U1638 (N_1638,In_314,In_410);
and U1639 (N_1639,In_824,In_1440);
nand U1640 (N_1640,In_55,In_599);
or U1641 (N_1641,In_870,In_1326);
xor U1642 (N_1642,In_1285,In_829);
or U1643 (N_1643,In_370,In_185);
xnor U1644 (N_1644,In_842,In_676);
or U1645 (N_1645,In_634,In_250);
nand U1646 (N_1646,In_150,In_328);
or U1647 (N_1647,In_241,In_624);
and U1648 (N_1648,In_499,In_665);
or U1649 (N_1649,In_825,In_422);
and U1650 (N_1650,In_1291,In_1134);
nor U1651 (N_1651,In_379,In_281);
nor U1652 (N_1652,In_863,In_458);
nand U1653 (N_1653,In_179,In_1386);
nand U1654 (N_1654,In_1133,In_9);
or U1655 (N_1655,In_261,In_161);
or U1656 (N_1656,In_23,In_777);
and U1657 (N_1657,In_392,In_1126);
xor U1658 (N_1658,In_938,In_718);
or U1659 (N_1659,In_192,In_1158);
nand U1660 (N_1660,In_1179,In_715);
xnor U1661 (N_1661,In_1365,In_335);
and U1662 (N_1662,In_921,In_1424);
and U1663 (N_1663,In_488,In_39);
or U1664 (N_1664,In_186,In_448);
nand U1665 (N_1665,In_391,In_668);
nand U1666 (N_1666,In_311,In_359);
nand U1667 (N_1667,In_624,In_1320);
or U1668 (N_1668,In_162,In_258);
or U1669 (N_1669,In_779,In_1409);
nor U1670 (N_1670,In_607,In_482);
nor U1671 (N_1671,In_822,In_1018);
nand U1672 (N_1672,In_937,In_1423);
or U1673 (N_1673,In_1062,In_6);
nor U1674 (N_1674,In_1282,In_431);
xnor U1675 (N_1675,In_1173,In_541);
or U1676 (N_1676,In_1101,In_634);
or U1677 (N_1677,In_103,In_1497);
and U1678 (N_1678,In_1147,In_1275);
and U1679 (N_1679,In_278,In_1046);
nand U1680 (N_1680,In_679,In_1298);
nor U1681 (N_1681,In_31,In_22);
or U1682 (N_1682,In_631,In_103);
nand U1683 (N_1683,In_1081,In_791);
xor U1684 (N_1684,In_801,In_1112);
xnor U1685 (N_1685,In_202,In_1043);
and U1686 (N_1686,In_181,In_354);
and U1687 (N_1687,In_293,In_443);
or U1688 (N_1688,In_1104,In_1390);
nor U1689 (N_1689,In_704,In_1398);
and U1690 (N_1690,In_393,In_491);
or U1691 (N_1691,In_564,In_361);
and U1692 (N_1692,In_964,In_579);
or U1693 (N_1693,In_1112,In_868);
nor U1694 (N_1694,In_131,In_1497);
and U1695 (N_1695,In_1419,In_431);
xnor U1696 (N_1696,In_329,In_655);
and U1697 (N_1697,In_918,In_259);
or U1698 (N_1698,In_267,In_667);
or U1699 (N_1699,In_1049,In_544);
xnor U1700 (N_1700,In_553,In_1452);
nand U1701 (N_1701,In_1390,In_1066);
nor U1702 (N_1702,In_439,In_666);
nor U1703 (N_1703,In_177,In_1290);
nor U1704 (N_1704,In_1004,In_561);
nand U1705 (N_1705,In_377,In_1397);
nor U1706 (N_1706,In_1152,In_1221);
or U1707 (N_1707,In_1428,In_125);
nand U1708 (N_1708,In_1291,In_300);
and U1709 (N_1709,In_147,In_364);
or U1710 (N_1710,In_995,In_1403);
xor U1711 (N_1711,In_1429,In_1324);
nand U1712 (N_1712,In_1409,In_362);
nor U1713 (N_1713,In_387,In_808);
nor U1714 (N_1714,In_621,In_559);
xor U1715 (N_1715,In_860,In_443);
nor U1716 (N_1716,In_1442,In_769);
nand U1717 (N_1717,In_199,In_1119);
nor U1718 (N_1718,In_658,In_849);
xnor U1719 (N_1719,In_1388,In_415);
and U1720 (N_1720,In_948,In_545);
nor U1721 (N_1721,In_638,In_204);
nor U1722 (N_1722,In_133,In_544);
or U1723 (N_1723,In_1434,In_1079);
nand U1724 (N_1724,In_177,In_133);
or U1725 (N_1725,In_1078,In_392);
nand U1726 (N_1726,In_1091,In_479);
and U1727 (N_1727,In_241,In_687);
nor U1728 (N_1728,In_1047,In_470);
or U1729 (N_1729,In_1006,In_238);
and U1730 (N_1730,In_481,In_1408);
nand U1731 (N_1731,In_64,In_513);
and U1732 (N_1732,In_1206,In_750);
xnor U1733 (N_1733,In_1198,In_1476);
nor U1734 (N_1734,In_44,In_13);
nand U1735 (N_1735,In_1136,In_850);
xor U1736 (N_1736,In_878,In_854);
or U1737 (N_1737,In_250,In_1161);
or U1738 (N_1738,In_90,In_48);
nor U1739 (N_1739,In_861,In_162);
or U1740 (N_1740,In_1036,In_579);
nand U1741 (N_1741,In_22,In_397);
or U1742 (N_1742,In_900,In_946);
or U1743 (N_1743,In_155,In_367);
nor U1744 (N_1744,In_598,In_1056);
xor U1745 (N_1745,In_721,In_1057);
and U1746 (N_1746,In_552,In_1199);
xnor U1747 (N_1747,In_239,In_311);
or U1748 (N_1748,In_641,In_1299);
and U1749 (N_1749,In_1209,In_1256);
nor U1750 (N_1750,In_153,In_1175);
nor U1751 (N_1751,In_788,In_731);
nand U1752 (N_1752,In_705,In_251);
and U1753 (N_1753,In_478,In_607);
xor U1754 (N_1754,In_202,In_167);
or U1755 (N_1755,In_1185,In_300);
and U1756 (N_1756,In_1305,In_1006);
nor U1757 (N_1757,In_108,In_1058);
nand U1758 (N_1758,In_19,In_914);
or U1759 (N_1759,In_715,In_1103);
or U1760 (N_1760,In_774,In_369);
and U1761 (N_1761,In_280,In_213);
and U1762 (N_1762,In_6,In_669);
or U1763 (N_1763,In_632,In_779);
or U1764 (N_1764,In_332,In_1328);
nand U1765 (N_1765,In_1165,In_971);
nand U1766 (N_1766,In_1353,In_1209);
or U1767 (N_1767,In_1119,In_168);
nor U1768 (N_1768,In_750,In_706);
or U1769 (N_1769,In_241,In_485);
nor U1770 (N_1770,In_106,In_227);
xnor U1771 (N_1771,In_422,In_778);
or U1772 (N_1772,In_327,In_281);
nand U1773 (N_1773,In_440,In_40);
or U1774 (N_1774,In_1225,In_1045);
xor U1775 (N_1775,In_587,In_1457);
nor U1776 (N_1776,In_822,In_1107);
xnor U1777 (N_1777,In_48,In_25);
xor U1778 (N_1778,In_1056,In_688);
and U1779 (N_1779,In_325,In_1309);
nor U1780 (N_1780,In_1122,In_193);
and U1781 (N_1781,In_533,In_1207);
xnor U1782 (N_1782,In_773,In_462);
nor U1783 (N_1783,In_160,In_591);
nor U1784 (N_1784,In_408,In_1463);
nor U1785 (N_1785,In_939,In_956);
and U1786 (N_1786,In_5,In_128);
and U1787 (N_1787,In_773,In_472);
nand U1788 (N_1788,In_186,In_160);
nor U1789 (N_1789,In_961,In_1488);
xor U1790 (N_1790,In_624,In_138);
nand U1791 (N_1791,In_569,In_957);
nor U1792 (N_1792,In_51,In_1130);
or U1793 (N_1793,In_1239,In_888);
nand U1794 (N_1794,In_119,In_1351);
and U1795 (N_1795,In_1180,In_25);
nand U1796 (N_1796,In_1120,In_915);
and U1797 (N_1797,In_860,In_576);
and U1798 (N_1798,In_88,In_1172);
nand U1799 (N_1799,In_99,In_759);
and U1800 (N_1800,In_1059,In_469);
xnor U1801 (N_1801,In_452,In_1313);
or U1802 (N_1802,In_1398,In_281);
and U1803 (N_1803,In_616,In_1283);
xnor U1804 (N_1804,In_305,In_1172);
or U1805 (N_1805,In_518,In_1142);
nor U1806 (N_1806,In_690,In_875);
nand U1807 (N_1807,In_1282,In_1253);
nor U1808 (N_1808,In_393,In_516);
and U1809 (N_1809,In_1088,In_502);
nor U1810 (N_1810,In_335,In_727);
or U1811 (N_1811,In_1427,In_1385);
nand U1812 (N_1812,In_1142,In_260);
xnor U1813 (N_1813,In_408,In_1079);
nor U1814 (N_1814,In_969,In_603);
nand U1815 (N_1815,In_569,In_283);
nor U1816 (N_1816,In_1200,In_347);
or U1817 (N_1817,In_560,In_111);
or U1818 (N_1818,In_268,In_854);
xnor U1819 (N_1819,In_672,In_550);
nand U1820 (N_1820,In_407,In_216);
or U1821 (N_1821,In_382,In_1052);
nor U1822 (N_1822,In_162,In_1006);
or U1823 (N_1823,In_414,In_1172);
xnor U1824 (N_1824,In_66,In_1415);
nand U1825 (N_1825,In_1304,In_385);
nand U1826 (N_1826,In_1355,In_458);
and U1827 (N_1827,In_1136,In_1085);
nand U1828 (N_1828,In_940,In_898);
or U1829 (N_1829,In_886,In_1421);
or U1830 (N_1830,In_685,In_656);
and U1831 (N_1831,In_83,In_892);
nand U1832 (N_1832,In_1181,In_1298);
nor U1833 (N_1833,In_162,In_1444);
or U1834 (N_1834,In_60,In_655);
nor U1835 (N_1835,In_154,In_588);
and U1836 (N_1836,In_1403,In_580);
nand U1837 (N_1837,In_668,In_739);
and U1838 (N_1838,In_1363,In_590);
nor U1839 (N_1839,In_1324,In_630);
xnor U1840 (N_1840,In_1032,In_1358);
nor U1841 (N_1841,In_805,In_898);
and U1842 (N_1842,In_462,In_570);
and U1843 (N_1843,In_161,In_500);
or U1844 (N_1844,In_534,In_922);
or U1845 (N_1845,In_1190,In_239);
nor U1846 (N_1846,In_580,In_437);
or U1847 (N_1847,In_1444,In_656);
nand U1848 (N_1848,In_570,In_224);
nor U1849 (N_1849,In_890,In_954);
xor U1850 (N_1850,In_941,In_724);
nand U1851 (N_1851,In_1165,In_489);
or U1852 (N_1852,In_390,In_711);
xor U1853 (N_1853,In_417,In_1291);
or U1854 (N_1854,In_1409,In_705);
xor U1855 (N_1855,In_857,In_688);
nand U1856 (N_1856,In_324,In_476);
nand U1857 (N_1857,In_853,In_1179);
nand U1858 (N_1858,In_119,In_580);
nand U1859 (N_1859,In_1458,In_711);
and U1860 (N_1860,In_1112,In_288);
nor U1861 (N_1861,In_772,In_1323);
or U1862 (N_1862,In_1032,In_466);
nand U1863 (N_1863,In_241,In_559);
or U1864 (N_1864,In_516,In_766);
and U1865 (N_1865,In_1369,In_31);
xnor U1866 (N_1866,In_132,In_175);
nor U1867 (N_1867,In_839,In_929);
and U1868 (N_1868,In_991,In_103);
or U1869 (N_1869,In_710,In_1084);
or U1870 (N_1870,In_589,In_1267);
or U1871 (N_1871,In_1312,In_1276);
xnor U1872 (N_1872,In_591,In_167);
nand U1873 (N_1873,In_1047,In_1254);
or U1874 (N_1874,In_604,In_1142);
or U1875 (N_1875,In_1094,In_1062);
or U1876 (N_1876,In_49,In_1223);
or U1877 (N_1877,In_440,In_1224);
or U1878 (N_1878,In_31,In_1164);
nand U1879 (N_1879,In_695,In_935);
and U1880 (N_1880,In_514,In_552);
or U1881 (N_1881,In_184,In_216);
and U1882 (N_1882,In_931,In_751);
nand U1883 (N_1883,In_1139,In_1183);
xor U1884 (N_1884,In_419,In_1135);
nand U1885 (N_1885,In_1470,In_792);
nand U1886 (N_1886,In_490,In_658);
and U1887 (N_1887,In_720,In_1394);
nand U1888 (N_1888,In_1474,In_278);
nor U1889 (N_1889,In_665,In_813);
nand U1890 (N_1890,In_500,In_960);
and U1891 (N_1891,In_1441,In_369);
nor U1892 (N_1892,In_765,In_911);
or U1893 (N_1893,In_342,In_896);
and U1894 (N_1894,In_889,In_242);
or U1895 (N_1895,In_911,In_610);
nand U1896 (N_1896,In_642,In_650);
or U1897 (N_1897,In_268,In_1318);
xnor U1898 (N_1898,In_301,In_1494);
or U1899 (N_1899,In_478,In_241);
and U1900 (N_1900,In_554,In_447);
xnor U1901 (N_1901,In_596,In_1067);
nor U1902 (N_1902,In_1353,In_416);
nand U1903 (N_1903,In_1253,In_386);
nand U1904 (N_1904,In_1181,In_1280);
and U1905 (N_1905,In_1471,In_421);
and U1906 (N_1906,In_1026,In_1404);
nor U1907 (N_1907,In_354,In_1075);
nand U1908 (N_1908,In_656,In_1199);
nor U1909 (N_1909,In_782,In_1033);
nand U1910 (N_1910,In_406,In_21);
xor U1911 (N_1911,In_131,In_483);
nand U1912 (N_1912,In_249,In_822);
and U1913 (N_1913,In_1164,In_300);
and U1914 (N_1914,In_166,In_338);
nand U1915 (N_1915,In_62,In_605);
nor U1916 (N_1916,In_528,In_105);
nor U1917 (N_1917,In_19,In_169);
and U1918 (N_1918,In_353,In_1220);
nand U1919 (N_1919,In_1263,In_822);
or U1920 (N_1920,In_1111,In_867);
xnor U1921 (N_1921,In_1073,In_96);
and U1922 (N_1922,In_448,In_284);
nand U1923 (N_1923,In_29,In_828);
nor U1924 (N_1924,In_548,In_940);
nor U1925 (N_1925,In_985,In_26);
nor U1926 (N_1926,In_454,In_1472);
and U1927 (N_1927,In_260,In_840);
nand U1928 (N_1928,In_647,In_1422);
nor U1929 (N_1929,In_1464,In_317);
and U1930 (N_1930,In_583,In_1464);
and U1931 (N_1931,In_1258,In_385);
and U1932 (N_1932,In_1446,In_1114);
or U1933 (N_1933,In_215,In_1255);
nand U1934 (N_1934,In_205,In_1368);
and U1935 (N_1935,In_1187,In_1286);
or U1936 (N_1936,In_1347,In_1387);
or U1937 (N_1937,In_399,In_1362);
or U1938 (N_1938,In_1141,In_578);
and U1939 (N_1939,In_911,In_1131);
xnor U1940 (N_1940,In_809,In_1394);
nor U1941 (N_1941,In_1224,In_835);
nand U1942 (N_1942,In_1380,In_1463);
xnor U1943 (N_1943,In_224,In_743);
and U1944 (N_1944,In_917,In_977);
and U1945 (N_1945,In_114,In_1087);
nand U1946 (N_1946,In_959,In_1328);
xor U1947 (N_1947,In_485,In_1452);
xnor U1948 (N_1948,In_52,In_610);
and U1949 (N_1949,In_580,In_899);
or U1950 (N_1950,In_1067,In_1480);
nor U1951 (N_1951,In_298,In_300);
and U1952 (N_1952,In_1476,In_1353);
nand U1953 (N_1953,In_776,In_255);
nor U1954 (N_1954,In_1107,In_1262);
nand U1955 (N_1955,In_707,In_910);
or U1956 (N_1956,In_1114,In_1334);
xnor U1957 (N_1957,In_684,In_436);
xnor U1958 (N_1958,In_220,In_665);
xnor U1959 (N_1959,In_779,In_119);
or U1960 (N_1960,In_531,In_745);
nand U1961 (N_1961,In_196,In_881);
or U1962 (N_1962,In_222,In_618);
nand U1963 (N_1963,In_433,In_428);
nand U1964 (N_1964,In_1261,In_1310);
nor U1965 (N_1965,In_602,In_573);
nor U1966 (N_1966,In_648,In_1447);
nor U1967 (N_1967,In_874,In_905);
or U1968 (N_1968,In_351,In_449);
and U1969 (N_1969,In_730,In_1474);
nand U1970 (N_1970,In_1301,In_789);
nor U1971 (N_1971,In_407,In_1375);
and U1972 (N_1972,In_284,In_1119);
and U1973 (N_1973,In_959,In_681);
nor U1974 (N_1974,In_836,In_21);
xnor U1975 (N_1975,In_1173,In_824);
nor U1976 (N_1976,In_1396,In_801);
nand U1977 (N_1977,In_484,In_1483);
nor U1978 (N_1978,In_170,In_751);
xor U1979 (N_1979,In_535,In_16);
nand U1980 (N_1980,In_751,In_1429);
nor U1981 (N_1981,In_85,In_966);
nor U1982 (N_1982,In_347,In_1354);
and U1983 (N_1983,In_1352,In_917);
or U1984 (N_1984,In_1131,In_1129);
and U1985 (N_1985,In_312,In_417);
nand U1986 (N_1986,In_714,In_547);
xor U1987 (N_1987,In_3,In_505);
and U1988 (N_1988,In_109,In_1092);
nand U1989 (N_1989,In_983,In_1454);
xnor U1990 (N_1990,In_940,In_82);
nand U1991 (N_1991,In_720,In_1441);
xnor U1992 (N_1992,In_1174,In_676);
nor U1993 (N_1993,In_398,In_617);
nand U1994 (N_1994,In_1226,In_1413);
and U1995 (N_1995,In_1070,In_450);
nand U1996 (N_1996,In_203,In_471);
xor U1997 (N_1997,In_293,In_1269);
xor U1998 (N_1998,In_1418,In_490);
xnor U1999 (N_1999,In_1002,In_939);
xnor U2000 (N_2000,In_319,In_1199);
and U2001 (N_2001,In_208,In_235);
nor U2002 (N_2002,In_34,In_1436);
or U2003 (N_2003,In_630,In_1106);
or U2004 (N_2004,In_272,In_1192);
or U2005 (N_2005,In_688,In_1407);
or U2006 (N_2006,In_406,In_1406);
xor U2007 (N_2007,In_1307,In_777);
or U2008 (N_2008,In_1375,In_576);
or U2009 (N_2009,In_278,In_61);
xnor U2010 (N_2010,In_81,In_555);
xor U2011 (N_2011,In_286,In_914);
nor U2012 (N_2012,In_999,In_1499);
or U2013 (N_2013,In_391,In_845);
or U2014 (N_2014,In_1131,In_90);
xor U2015 (N_2015,In_189,In_1136);
nand U2016 (N_2016,In_141,In_888);
or U2017 (N_2017,In_73,In_672);
nor U2018 (N_2018,In_1327,In_1313);
or U2019 (N_2019,In_925,In_395);
nand U2020 (N_2020,In_1315,In_1047);
nand U2021 (N_2021,In_1380,In_715);
nor U2022 (N_2022,In_1062,In_1137);
nand U2023 (N_2023,In_1329,In_235);
and U2024 (N_2024,In_400,In_847);
and U2025 (N_2025,In_1114,In_503);
and U2026 (N_2026,In_1091,In_283);
nor U2027 (N_2027,In_508,In_820);
xor U2028 (N_2028,In_79,In_40);
nor U2029 (N_2029,In_83,In_1202);
nor U2030 (N_2030,In_651,In_259);
nand U2031 (N_2031,In_294,In_472);
xnor U2032 (N_2032,In_115,In_417);
nand U2033 (N_2033,In_1385,In_1047);
and U2034 (N_2034,In_697,In_446);
xnor U2035 (N_2035,In_198,In_536);
xor U2036 (N_2036,In_742,In_1374);
xnor U2037 (N_2037,In_841,In_421);
nor U2038 (N_2038,In_762,In_33);
nor U2039 (N_2039,In_972,In_590);
xnor U2040 (N_2040,In_1211,In_1419);
xor U2041 (N_2041,In_761,In_1237);
nand U2042 (N_2042,In_554,In_138);
xnor U2043 (N_2043,In_873,In_480);
or U2044 (N_2044,In_1134,In_174);
or U2045 (N_2045,In_249,In_160);
or U2046 (N_2046,In_1230,In_860);
xnor U2047 (N_2047,In_714,In_334);
or U2048 (N_2048,In_493,In_447);
nor U2049 (N_2049,In_405,In_1283);
and U2050 (N_2050,In_530,In_519);
nor U2051 (N_2051,In_127,In_999);
or U2052 (N_2052,In_270,In_581);
nor U2053 (N_2053,In_780,In_980);
or U2054 (N_2054,In_1478,In_1484);
nand U2055 (N_2055,In_178,In_29);
nor U2056 (N_2056,In_970,In_1151);
and U2057 (N_2057,In_883,In_72);
xnor U2058 (N_2058,In_184,In_1044);
nand U2059 (N_2059,In_215,In_305);
nor U2060 (N_2060,In_174,In_1041);
nor U2061 (N_2061,In_550,In_1346);
nand U2062 (N_2062,In_880,In_824);
and U2063 (N_2063,In_150,In_867);
xnor U2064 (N_2064,In_258,In_1380);
nor U2065 (N_2065,In_1137,In_44);
xor U2066 (N_2066,In_149,In_138);
and U2067 (N_2067,In_1005,In_245);
and U2068 (N_2068,In_732,In_1077);
xnor U2069 (N_2069,In_213,In_44);
or U2070 (N_2070,In_582,In_574);
nand U2071 (N_2071,In_874,In_230);
nor U2072 (N_2072,In_974,In_706);
nor U2073 (N_2073,In_686,In_611);
or U2074 (N_2074,In_1306,In_930);
and U2075 (N_2075,In_281,In_666);
and U2076 (N_2076,In_925,In_872);
and U2077 (N_2077,In_1208,In_1434);
or U2078 (N_2078,In_323,In_1004);
nand U2079 (N_2079,In_689,In_1331);
nand U2080 (N_2080,In_1372,In_1295);
or U2081 (N_2081,In_755,In_1331);
xnor U2082 (N_2082,In_475,In_83);
or U2083 (N_2083,In_322,In_1121);
nor U2084 (N_2084,In_140,In_367);
nor U2085 (N_2085,In_1265,In_636);
xnor U2086 (N_2086,In_105,In_1282);
and U2087 (N_2087,In_873,In_987);
or U2088 (N_2088,In_417,In_586);
or U2089 (N_2089,In_953,In_957);
nor U2090 (N_2090,In_396,In_45);
xnor U2091 (N_2091,In_134,In_641);
nand U2092 (N_2092,In_240,In_711);
xor U2093 (N_2093,In_1470,In_536);
nand U2094 (N_2094,In_1225,In_615);
or U2095 (N_2095,In_709,In_1048);
xnor U2096 (N_2096,In_940,In_728);
and U2097 (N_2097,In_1213,In_106);
or U2098 (N_2098,In_285,In_198);
nor U2099 (N_2099,In_213,In_881);
nand U2100 (N_2100,In_1418,In_733);
and U2101 (N_2101,In_1111,In_754);
and U2102 (N_2102,In_173,In_1130);
nor U2103 (N_2103,In_758,In_1028);
nor U2104 (N_2104,In_455,In_1456);
and U2105 (N_2105,In_798,In_579);
xor U2106 (N_2106,In_1430,In_276);
nand U2107 (N_2107,In_0,In_1390);
nor U2108 (N_2108,In_476,In_827);
nor U2109 (N_2109,In_779,In_404);
nor U2110 (N_2110,In_1359,In_526);
nor U2111 (N_2111,In_49,In_1030);
nand U2112 (N_2112,In_1287,In_950);
nor U2113 (N_2113,In_550,In_1111);
and U2114 (N_2114,In_211,In_413);
or U2115 (N_2115,In_996,In_1087);
or U2116 (N_2116,In_424,In_55);
nor U2117 (N_2117,In_180,In_956);
or U2118 (N_2118,In_716,In_845);
and U2119 (N_2119,In_447,In_1288);
xnor U2120 (N_2120,In_1125,In_994);
nor U2121 (N_2121,In_276,In_343);
and U2122 (N_2122,In_1034,In_1013);
xor U2123 (N_2123,In_109,In_1452);
or U2124 (N_2124,In_880,In_555);
nor U2125 (N_2125,In_1442,In_716);
xor U2126 (N_2126,In_664,In_1216);
nor U2127 (N_2127,In_1046,In_1024);
nand U2128 (N_2128,In_422,In_668);
nor U2129 (N_2129,In_642,In_140);
nand U2130 (N_2130,In_1489,In_886);
and U2131 (N_2131,In_548,In_1056);
nor U2132 (N_2132,In_955,In_1281);
nand U2133 (N_2133,In_1182,In_278);
nor U2134 (N_2134,In_475,In_147);
nor U2135 (N_2135,In_45,In_1237);
xor U2136 (N_2136,In_581,In_1043);
nor U2137 (N_2137,In_990,In_878);
nand U2138 (N_2138,In_136,In_707);
and U2139 (N_2139,In_290,In_1087);
and U2140 (N_2140,In_1461,In_1081);
or U2141 (N_2141,In_290,In_65);
nor U2142 (N_2142,In_750,In_954);
nand U2143 (N_2143,In_1445,In_121);
or U2144 (N_2144,In_1018,In_630);
or U2145 (N_2145,In_974,In_555);
nor U2146 (N_2146,In_181,In_1031);
nor U2147 (N_2147,In_1011,In_153);
nand U2148 (N_2148,In_255,In_256);
xor U2149 (N_2149,In_1139,In_1338);
nor U2150 (N_2150,In_993,In_1250);
and U2151 (N_2151,In_1213,In_384);
nor U2152 (N_2152,In_45,In_73);
nor U2153 (N_2153,In_339,In_578);
nand U2154 (N_2154,In_1337,In_490);
xor U2155 (N_2155,In_1409,In_1294);
xnor U2156 (N_2156,In_1162,In_299);
nand U2157 (N_2157,In_13,In_91);
nand U2158 (N_2158,In_1076,In_505);
nor U2159 (N_2159,In_476,In_70);
xnor U2160 (N_2160,In_602,In_108);
or U2161 (N_2161,In_1133,In_18);
and U2162 (N_2162,In_827,In_373);
nand U2163 (N_2163,In_912,In_144);
and U2164 (N_2164,In_352,In_1439);
or U2165 (N_2165,In_1235,In_411);
or U2166 (N_2166,In_297,In_89);
or U2167 (N_2167,In_1330,In_458);
nor U2168 (N_2168,In_864,In_940);
and U2169 (N_2169,In_1089,In_649);
and U2170 (N_2170,In_1193,In_360);
nor U2171 (N_2171,In_125,In_1225);
nor U2172 (N_2172,In_1151,In_245);
or U2173 (N_2173,In_354,In_899);
or U2174 (N_2174,In_382,In_949);
nand U2175 (N_2175,In_115,In_191);
nor U2176 (N_2176,In_828,In_163);
and U2177 (N_2177,In_1327,In_685);
xor U2178 (N_2178,In_314,In_283);
and U2179 (N_2179,In_14,In_102);
nor U2180 (N_2180,In_1296,In_711);
xnor U2181 (N_2181,In_16,In_176);
and U2182 (N_2182,In_1336,In_733);
nand U2183 (N_2183,In_178,In_798);
nand U2184 (N_2184,In_912,In_1294);
xor U2185 (N_2185,In_324,In_1396);
or U2186 (N_2186,In_194,In_326);
xor U2187 (N_2187,In_807,In_430);
xnor U2188 (N_2188,In_53,In_1027);
nand U2189 (N_2189,In_471,In_1086);
nor U2190 (N_2190,In_615,In_521);
nand U2191 (N_2191,In_767,In_1491);
nand U2192 (N_2192,In_280,In_811);
nand U2193 (N_2193,In_714,In_789);
or U2194 (N_2194,In_1059,In_832);
or U2195 (N_2195,In_1101,In_571);
and U2196 (N_2196,In_1428,In_1295);
and U2197 (N_2197,In_1306,In_778);
xnor U2198 (N_2198,In_264,In_1418);
nand U2199 (N_2199,In_117,In_969);
and U2200 (N_2200,In_594,In_1461);
and U2201 (N_2201,In_1189,In_1138);
xor U2202 (N_2202,In_1395,In_163);
xor U2203 (N_2203,In_886,In_992);
nor U2204 (N_2204,In_548,In_841);
xor U2205 (N_2205,In_415,In_882);
nand U2206 (N_2206,In_46,In_1213);
nor U2207 (N_2207,In_930,In_683);
or U2208 (N_2208,In_343,In_623);
nand U2209 (N_2209,In_791,In_78);
nand U2210 (N_2210,In_155,In_638);
nand U2211 (N_2211,In_1092,In_883);
nand U2212 (N_2212,In_739,In_145);
nor U2213 (N_2213,In_1352,In_725);
nor U2214 (N_2214,In_491,In_205);
nand U2215 (N_2215,In_866,In_576);
or U2216 (N_2216,In_97,In_393);
nand U2217 (N_2217,In_941,In_586);
nand U2218 (N_2218,In_1179,In_32);
or U2219 (N_2219,In_1274,In_269);
nor U2220 (N_2220,In_990,In_980);
nor U2221 (N_2221,In_864,In_491);
or U2222 (N_2222,In_202,In_1116);
and U2223 (N_2223,In_1318,In_643);
and U2224 (N_2224,In_690,In_185);
nor U2225 (N_2225,In_876,In_525);
or U2226 (N_2226,In_889,In_679);
nand U2227 (N_2227,In_1377,In_320);
or U2228 (N_2228,In_1334,In_933);
xnor U2229 (N_2229,In_100,In_626);
and U2230 (N_2230,In_1294,In_785);
and U2231 (N_2231,In_894,In_973);
nor U2232 (N_2232,In_1071,In_900);
nand U2233 (N_2233,In_405,In_785);
or U2234 (N_2234,In_1115,In_1068);
nor U2235 (N_2235,In_951,In_1306);
or U2236 (N_2236,In_1265,In_497);
and U2237 (N_2237,In_1005,In_87);
or U2238 (N_2238,In_373,In_969);
nand U2239 (N_2239,In_677,In_280);
xor U2240 (N_2240,In_667,In_464);
and U2241 (N_2241,In_803,In_682);
xor U2242 (N_2242,In_550,In_1378);
and U2243 (N_2243,In_59,In_859);
nor U2244 (N_2244,In_1154,In_1043);
or U2245 (N_2245,In_756,In_1450);
or U2246 (N_2246,In_1277,In_489);
nand U2247 (N_2247,In_498,In_1493);
and U2248 (N_2248,In_658,In_1139);
xnor U2249 (N_2249,In_748,In_1393);
or U2250 (N_2250,In_624,In_773);
nor U2251 (N_2251,In_942,In_246);
or U2252 (N_2252,In_1454,In_1180);
nand U2253 (N_2253,In_212,In_1103);
nor U2254 (N_2254,In_692,In_955);
or U2255 (N_2255,In_89,In_62);
nor U2256 (N_2256,In_774,In_98);
and U2257 (N_2257,In_538,In_552);
nand U2258 (N_2258,In_415,In_712);
and U2259 (N_2259,In_1368,In_849);
nand U2260 (N_2260,In_301,In_717);
nand U2261 (N_2261,In_1143,In_348);
nor U2262 (N_2262,In_756,In_490);
xnor U2263 (N_2263,In_506,In_298);
nor U2264 (N_2264,In_828,In_410);
nor U2265 (N_2265,In_1172,In_207);
xnor U2266 (N_2266,In_124,In_1321);
or U2267 (N_2267,In_1299,In_218);
nand U2268 (N_2268,In_671,In_255);
xor U2269 (N_2269,In_1073,In_205);
nor U2270 (N_2270,In_939,In_535);
or U2271 (N_2271,In_1089,In_771);
or U2272 (N_2272,In_26,In_658);
nand U2273 (N_2273,In_1161,In_494);
or U2274 (N_2274,In_1302,In_646);
nand U2275 (N_2275,In_1006,In_92);
nand U2276 (N_2276,In_1143,In_1150);
nor U2277 (N_2277,In_1437,In_809);
nand U2278 (N_2278,In_459,In_1039);
or U2279 (N_2279,In_1097,In_592);
nor U2280 (N_2280,In_506,In_621);
nor U2281 (N_2281,In_947,In_708);
nand U2282 (N_2282,In_943,In_1498);
nand U2283 (N_2283,In_1211,In_989);
nand U2284 (N_2284,In_1469,In_1115);
nand U2285 (N_2285,In_1466,In_251);
xnor U2286 (N_2286,In_468,In_70);
and U2287 (N_2287,In_761,In_1072);
nand U2288 (N_2288,In_1126,In_991);
and U2289 (N_2289,In_1222,In_59);
and U2290 (N_2290,In_752,In_101);
or U2291 (N_2291,In_86,In_616);
and U2292 (N_2292,In_1335,In_663);
nand U2293 (N_2293,In_759,In_9);
nor U2294 (N_2294,In_518,In_502);
nor U2295 (N_2295,In_970,In_9);
or U2296 (N_2296,In_1049,In_570);
or U2297 (N_2297,In_95,In_791);
or U2298 (N_2298,In_1267,In_1469);
nor U2299 (N_2299,In_601,In_245);
nand U2300 (N_2300,In_203,In_1121);
xor U2301 (N_2301,In_368,In_248);
nor U2302 (N_2302,In_1028,In_75);
nand U2303 (N_2303,In_917,In_683);
xor U2304 (N_2304,In_1279,In_373);
or U2305 (N_2305,In_1246,In_158);
nand U2306 (N_2306,In_228,In_1492);
or U2307 (N_2307,In_1104,In_941);
nand U2308 (N_2308,In_546,In_101);
or U2309 (N_2309,In_261,In_1058);
and U2310 (N_2310,In_1455,In_520);
nor U2311 (N_2311,In_584,In_1191);
nand U2312 (N_2312,In_687,In_1410);
and U2313 (N_2313,In_16,In_1283);
xnor U2314 (N_2314,In_1453,In_1438);
nand U2315 (N_2315,In_850,In_1289);
and U2316 (N_2316,In_106,In_1118);
or U2317 (N_2317,In_230,In_575);
and U2318 (N_2318,In_789,In_760);
or U2319 (N_2319,In_185,In_1365);
and U2320 (N_2320,In_137,In_524);
nor U2321 (N_2321,In_405,In_838);
and U2322 (N_2322,In_1473,In_1334);
and U2323 (N_2323,In_597,In_420);
xnor U2324 (N_2324,In_790,In_710);
nand U2325 (N_2325,In_958,In_28);
and U2326 (N_2326,In_202,In_1090);
nor U2327 (N_2327,In_990,In_443);
xnor U2328 (N_2328,In_252,In_1094);
nand U2329 (N_2329,In_307,In_1462);
xnor U2330 (N_2330,In_1055,In_479);
nand U2331 (N_2331,In_878,In_455);
nand U2332 (N_2332,In_1039,In_428);
nor U2333 (N_2333,In_422,In_101);
xor U2334 (N_2334,In_393,In_1446);
xnor U2335 (N_2335,In_665,In_900);
and U2336 (N_2336,In_401,In_283);
nand U2337 (N_2337,In_391,In_1195);
or U2338 (N_2338,In_1410,In_463);
or U2339 (N_2339,In_194,In_766);
xor U2340 (N_2340,In_1294,In_1491);
or U2341 (N_2341,In_184,In_148);
nand U2342 (N_2342,In_1293,In_1105);
nor U2343 (N_2343,In_929,In_176);
and U2344 (N_2344,In_741,In_85);
xor U2345 (N_2345,In_852,In_649);
xor U2346 (N_2346,In_563,In_190);
nand U2347 (N_2347,In_983,In_223);
nand U2348 (N_2348,In_625,In_654);
nor U2349 (N_2349,In_735,In_19);
xnor U2350 (N_2350,In_358,In_708);
xnor U2351 (N_2351,In_1407,In_1270);
and U2352 (N_2352,In_824,In_127);
nand U2353 (N_2353,In_1028,In_535);
or U2354 (N_2354,In_572,In_740);
nand U2355 (N_2355,In_123,In_544);
nor U2356 (N_2356,In_1351,In_83);
or U2357 (N_2357,In_1178,In_1010);
nand U2358 (N_2358,In_386,In_1021);
xnor U2359 (N_2359,In_73,In_695);
nand U2360 (N_2360,In_123,In_1406);
nand U2361 (N_2361,In_569,In_936);
nor U2362 (N_2362,In_766,In_1367);
and U2363 (N_2363,In_683,In_573);
nand U2364 (N_2364,In_1077,In_762);
xnor U2365 (N_2365,In_477,In_1285);
nand U2366 (N_2366,In_296,In_35);
and U2367 (N_2367,In_262,In_66);
xor U2368 (N_2368,In_1038,In_1224);
and U2369 (N_2369,In_51,In_797);
or U2370 (N_2370,In_885,In_22);
xor U2371 (N_2371,In_988,In_753);
nor U2372 (N_2372,In_859,In_1398);
or U2373 (N_2373,In_953,In_369);
nor U2374 (N_2374,In_816,In_1385);
and U2375 (N_2375,In_67,In_160);
or U2376 (N_2376,In_1144,In_952);
xor U2377 (N_2377,In_588,In_756);
xnor U2378 (N_2378,In_138,In_1329);
and U2379 (N_2379,In_1357,In_1353);
and U2380 (N_2380,In_1337,In_536);
and U2381 (N_2381,In_663,In_1486);
nand U2382 (N_2382,In_483,In_846);
and U2383 (N_2383,In_868,In_584);
xnor U2384 (N_2384,In_1274,In_766);
and U2385 (N_2385,In_1331,In_655);
nand U2386 (N_2386,In_691,In_1286);
nor U2387 (N_2387,In_1234,In_1243);
xor U2388 (N_2388,In_1494,In_233);
and U2389 (N_2389,In_1465,In_340);
nand U2390 (N_2390,In_934,In_1239);
or U2391 (N_2391,In_1480,In_1488);
nand U2392 (N_2392,In_749,In_1449);
or U2393 (N_2393,In_48,In_782);
nand U2394 (N_2394,In_213,In_63);
or U2395 (N_2395,In_330,In_929);
nor U2396 (N_2396,In_639,In_366);
or U2397 (N_2397,In_474,In_1075);
nand U2398 (N_2398,In_1308,In_220);
xnor U2399 (N_2399,In_211,In_844);
nor U2400 (N_2400,In_553,In_576);
nor U2401 (N_2401,In_739,In_228);
nor U2402 (N_2402,In_609,In_1251);
nand U2403 (N_2403,In_97,In_106);
xor U2404 (N_2404,In_950,In_1383);
xnor U2405 (N_2405,In_1020,In_1385);
nand U2406 (N_2406,In_1488,In_827);
xnor U2407 (N_2407,In_1208,In_106);
xnor U2408 (N_2408,In_1292,In_1381);
nand U2409 (N_2409,In_1262,In_832);
xor U2410 (N_2410,In_1357,In_1041);
nor U2411 (N_2411,In_1213,In_617);
nand U2412 (N_2412,In_621,In_1375);
and U2413 (N_2413,In_1025,In_562);
and U2414 (N_2414,In_424,In_1066);
xor U2415 (N_2415,In_1343,In_786);
or U2416 (N_2416,In_862,In_733);
nor U2417 (N_2417,In_954,In_179);
nor U2418 (N_2418,In_154,In_555);
nand U2419 (N_2419,In_1490,In_748);
and U2420 (N_2420,In_167,In_532);
and U2421 (N_2421,In_496,In_444);
nor U2422 (N_2422,In_205,In_1079);
nor U2423 (N_2423,In_520,In_1305);
nor U2424 (N_2424,In_1318,In_695);
nand U2425 (N_2425,In_357,In_993);
nand U2426 (N_2426,In_1357,In_1124);
or U2427 (N_2427,In_552,In_143);
nor U2428 (N_2428,In_344,In_1109);
nor U2429 (N_2429,In_112,In_665);
or U2430 (N_2430,In_1216,In_1143);
nand U2431 (N_2431,In_649,In_1325);
nand U2432 (N_2432,In_949,In_1007);
xor U2433 (N_2433,In_813,In_666);
and U2434 (N_2434,In_704,In_1457);
nor U2435 (N_2435,In_492,In_1027);
xnor U2436 (N_2436,In_586,In_1380);
nand U2437 (N_2437,In_608,In_710);
and U2438 (N_2438,In_155,In_1109);
and U2439 (N_2439,In_373,In_37);
xor U2440 (N_2440,In_687,In_158);
xnor U2441 (N_2441,In_648,In_407);
nor U2442 (N_2442,In_398,In_335);
nand U2443 (N_2443,In_586,In_1130);
xor U2444 (N_2444,In_632,In_117);
and U2445 (N_2445,In_916,In_1230);
nand U2446 (N_2446,In_1254,In_1006);
xnor U2447 (N_2447,In_842,In_931);
xnor U2448 (N_2448,In_1365,In_584);
nand U2449 (N_2449,In_364,In_191);
or U2450 (N_2450,In_93,In_921);
or U2451 (N_2451,In_1437,In_903);
and U2452 (N_2452,In_179,In_628);
or U2453 (N_2453,In_484,In_1256);
and U2454 (N_2454,In_1321,In_1365);
and U2455 (N_2455,In_1374,In_324);
nand U2456 (N_2456,In_1106,In_1430);
and U2457 (N_2457,In_155,In_788);
nand U2458 (N_2458,In_381,In_1292);
or U2459 (N_2459,In_623,In_383);
and U2460 (N_2460,In_346,In_294);
nor U2461 (N_2461,In_331,In_695);
nor U2462 (N_2462,In_821,In_499);
nor U2463 (N_2463,In_15,In_1110);
and U2464 (N_2464,In_757,In_807);
or U2465 (N_2465,In_850,In_1444);
or U2466 (N_2466,In_1177,In_918);
and U2467 (N_2467,In_1295,In_78);
and U2468 (N_2468,In_739,In_131);
xor U2469 (N_2469,In_133,In_566);
nor U2470 (N_2470,In_1462,In_1221);
and U2471 (N_2471,In_440,In_1126);
nand U2472 (N_2472,In_372,In_775);
or U2473 (N_2473,In_1094,In_1281);
or U2474 (N_2474,In_509,In_570);
or U2475 (N_2475,In_1119,In_876);
or U2476 (N_2476,In_1044,In_452);
and U2477 (N_2477,In_139,In_80);
xor U2478 (N_2478,In_99,In_815);
or U2479 (N_2479,In_98,In_70);
and U2480 (N_2480,In_292,In_1217);
or U2481 (N_2481,In_267,In_1236);
or U2482 (N_2482,In_1092,In_654);
or U2483 (N_2483,In_394,In_1459);
nand U2484 (N_2484,In_1405,In_935);
xnor U2485 (N_2485,In_1405,In_501);
and U2486 (N_2486,In_1042,In_1067);
and U2487 (N_2487,In_993,In_1481);
and U2488 (N_2488,In_939,In_643);
nand U2489 (N_2489,In_970,In_413);
or U2490 (N_2490,In_647,In_710);
nor U2491 (N_2491,In_1056,In_118);
and U2492 (N_2492,In_677,In_772);
xnor U2493 (N_2493,In_827,In_1110);
nand U2494 (N_2494,In_812,In_26);
nor U2495 (N_2495,In_1007,In_352);
nor U2496 (N_2496,In_1291,In_1195);
nand U2497 (N_2497,In_948,In_287);
nor U2498 (N_2498,In_1383,In_569);
nand U2499 (N_2499,In_603,In_318);
nor U2500 (N_2500,In_1109,In_1480);
nand U2501 (N_2501,In_1017,In_173);
and U2502 (N_2502,In_1174,In_183);
and U2503 (N_2503,In_1068,In_936);
xor U2504 (N_2504,In_204,In_395);
nand U2505 (N_2505,In_755,In_919);
xor U2506 (N_2506,In_226,In_1300);
or U2507 (N_2507,In_784,In_748);
nor U2508 (N_2508,In_205,In_56);
nor U2509 (N_2509,In_634,In_135);
or U2510 (N_2510,In_322,In_3);
xnor U2511 (N_2511,In_409,In_399);
or U2512 (N_2512,In_1232,In_134);
and U2513 (N_2513,In_964,In_214);
or U2514 (N_2514,In_1128,In_371);
or U2515 (N_2515,In_581,In_252);
xnor U2516 (N_2516,In_1349,In_1321);
or U2517 (N_2517,In_708,In_1283);
xnor U2518 (N_2518,In_1452,In_777);
nor U2519 (N_2519,In_353,In_430);
and U2520 (N_2520,In_451,In_416);
nor U2521 (N_2521,In_849,In_861);
or U2522 (N_2522,In_280,In_1057);
nand U2523 (N_2523,In_756,In_549);
nor U2524 (N_2524,In_2,In_1251);
or U2525 (N_2525,In_776,In_100);
and U2526 (N_2526,In_404,In_1144);
and U2527 (N_2527,In_797,In_453);
nand U2528 (N_2528,In_1494,In_557);
xnor U2529 (N_2529,In_526,In_1035);
or U2530 (N_2530,In_1451,In_793);
and U2531 (N_2531,In_521,In_1336);
nand U2532 (N_2532,In_195,In_4);
nor U2533 (N_2533,In_465,In_810);
and U2534 (N_2534,In_127,In_535);
nand U2535 (N_2535,In_1084,In_1470);
nor U2536 (N_2536,In_601,In_502);
and U2537 (N_2537,In_927,In_80);
xor U2538 (N_2538,In_743,In_565);
nor U2539 (N_2539,In_634,In_1158);
or U2540 (N_2540,In_7,In_966);
xnor U2541 (N_2541,In_257,In_823);
xnor U2542 (N_2542,In_380,In_1367);
nand U2543 (N_2543,In_617,In_1080);
xor U2544 (N_2544,In_1374,In_102);
nor U2545 (N_2545,In_1450,In_3);
and U2546 (N_2546,In_887,In_1044);
nand U2547 (N_2547,In_1464,In_156);
xnor U2548 (N_2548,In_1035,In_517);
xnor U2549 (N_2549,In_1389,In_776);
xnor U2550 (N_2550,In_523,In_1197);
nand U2551 (N_2551,In_613,In_234);
nand U2552 (N_2552,In_759,In_364);
and U2553 (N_2553,In_37,In_1435);
and U2554 (N_2554,In_828,In_1375);
nand U2555 (N_2555,In_391,In_1251);
and U2556 (N_2556,In_594,In_428);
or U2557 (N_2557,In_1359,In_959);
or U2558 (N_2558,In_625,In_1474);
nor U2559 (N_2559,In_1415,In_1412);
nor U2560 (N_2560,In_138,In_7);
or U2561 (N_2561,In_106,In_1128);
or U2562 (N_2562,In_803,In_1035);
nor U2563 (N_2563,In_1292,In_392);
xor U2564 (N_2564,In_872,In_401);
nor U2565 (N_2565,In_460,In_659);
nor U2566 (N_2566,In_1024,In_761);
nor U2567 (N_2567,In_961,In_10);
or U2568 (N_2568,In_1136,In_705);
nor U2569 (N_2569,In_538,In_171);
xor U2570 (N_2570,In_1213,In_1352);
xor U2571 (N_2571,In_1102,In_820);
or U2572 (N_2572,In_909,In_405);
or U2573 (N_2573,In_978,In_207);
or U2574 (N_2574,In_1045,In_1169);
xor U2575 (N_2575,In_732,In_1044);
nand U2576 (N_2576,In_414,In_98);
nand U2577 (N_2577,In_46,In_927);
and U2578 (N_2578,In_1430,In_1208);
nor U2579 (N_2579,In_1114,In_216);
and U2580 (N_2580,In_1293,In_583);
or U2581 (N_2581,In_1356,In_530);
or U2582 (N_2582,In_831,In_421);
xor U2583 (N_2583,In_359,In_132);
or U2584 (N_2584,In_922,In_981);
or U2585 (N_2585,In_608,In_796);
xnor U2586 (N_2586,In_402,In_679);
xnor U2587 (N_2587,In_1054,In_555);
xnor U2588 (N_2588,In_619,In_812);
and U2589 (N_2589,In_258,In_882);
xnor U2590 (N_2590,In_1476,In_1266);
or U2591 (N_2591,In_597,In_1187);
and U2592 (N_2592,In_794,In_1048);
nor U2593 (N_2593,In_33,In_252);
nor U2594 (N_2594,In_591,In_710);
nor U2595 (N_2595,In_1196,In_112);
nor U2596 (N_2596,In_925,In_412);
xnor U2597 (N_2597,In_856,In_810);
or U2598 (N_2598,In_341,In_655);
xnor U2599 (N_2599,In_1218,In_1270);
and U2600 (N_2600,In_1341,In_688);
xnor U2601 (N_2601,In_476,In_1102);
nor U2602 (N_2602,In_1456,In_367);
and U2603 (N_2603,In_987,In_721);
and U2604 (N_2604,In_976,In_629);
xor U2605 (N_2605,In_169,In_184);
xnor U2606 (N_2606,In_1335,In_938);
or U2607 (N_2607,In_1330,In_1424);
or U2608 (N_2608,In_694,In_582);
or U2609 (N_2609,In_504,In_525);
xor U2610 (N_2610,In_190,In_936);
nand U2611 (N_2611,In_1191,In_27);
and U2612 (N_2612,In_371,In_701);
nor U2613 (N_2613,In_937,In_1216);
xor U2614 (N_2614,In_61,In_959);
xnor U2615 (N_2615,In_1493,In_505);
nor U2616 (N_2616,In_1098,In_998);
xnor U2617 (N_2617,In_622,In_567);
or U2618 (N_2618,In_674,In_291);
and U2619 (N_2619,In_127,In_1415);
nor U2620 (N_2620,In_1163,In_1434);
and U2621 (N_2621,In_1183,In_899);
xnor U2622 (N_2622,In_442,In_984);
nor U2623 (N_2623,In_289,In_733);
or U2624 (N_2624,In_791,In_691);
or U2625 (N_2625,In_327,In_257);
and U2626 (N_2626,In_54,In_195);
xnor U2627 (N_2627,In_439,In_1273);
nor U2628 (N_2628,In_482,In_1358);
nand U2629 (N_2629,In_263,In_279);
or U2630 (N_2630,In_1043,In_621);
nor U2631 (N_2631,In_1144,In_831);
nand U2632 (N_2632,In_436,In_239);
or U2633 (N_2633,In_934,In_1415);
nor U2634 (N_2634,In_838,In_1092);
and U2635 (N_2635,In_743,In_321);
or U2636 (N_2636,In_244,In_357);
xnor U2637 (N_2637,In_303,In_499);
and U2638 (N_2638,In_1470,In_159);
xor U2639 (N_2639,In_1210,In_1086);
nor U2640 (N_2640,In_1265,In_686);
or U2641 (N_2641,In_1091,In_731);
nand U2642 (N_2642,In_574,In_1082);
nand U2643 (N_2643,In_1351,In_1070);
xnor U2644 (N_2644,In_360,In_341);
and U2645 (N_2645,In_1140,In_702);
or U2646 (N_2646,In_1130,In_688);
and U2647 (N_2647,In_561,In_877);
or U2648 (N_2648,In_1335,In_1355);
xor U2649 (N_2649,In_81,In_1206);
xor U2650 (N_2650,In_1026,In_44);
nand U2651 (N_2651,In_922,In_233);
or U2652 (N_2652,In_893,In_679);
nor U2653 (N_2653,In_928,In_193);
xnor U2654 (N_2654,In_1311,In_96);
and U2655 (N_2655,In_1476,In_1433);
nor U2656 (N_2656,In_721,In_601);
nor U2657 (N_2657,In_279,In_206);
nand U2658 (N_2658,In_1203,In_569);
nor U2659 (N_2659,In_1216,In_206);
or U2660 (N_2660,In_1451,In_998);
xor U2661 (N_2661,In_1231,In_653);
nor U2662 (N_2662,In_668,In_1154);
nand U2663 (N_2663,In_335,In_190);
xnor U2664 (N_2664,In_1358,In_1253);
nand U2665 (N_2665,In_10,In_1332);
xor U2666 (N_2666,In_1299,In_252);
and U2667 (N_2667,In_490,In_1006);
or U2668 (N_2668,In_619,In_1219);
or U2669 (N_2669,In_261,In_568);
and U2670 (N_2670,In_280,In_392);
nor U2671 (N_2671,In_741,In_765);
nor U2672 (N_2672,In_1055,In_1377);
and U2673 (N_2673,In_1444,In_1497);
and U2674 (N_2674,In_785,In_827);
xnor U2675 (N_2675,In_1498,In_1384);
and U2676 (N_2676,In_1023,In_175);
or U2677 (N_2677,In_1420,In_258);
nor U2678 (N_2678,In_475,In_1067);
or U2679 (N_2679,In_11,In_91);
or U2680 (N_2680,In_114,In_908);
nand U2681 (N_2681,In_1004,In_413);
xor U2682 (N_2682,In_73,In_946);
or U2683 (N_2683,In_1136,In_1098);
nor U2684 (N_2684,In_1271,In_734);
nor U2685 (N_2685,In_615,In_440);
xor U2686 (N_2686,In_516,In_1172);
xnor U2687 (N_2687,In_259,In_1377);
or U2688 (N_2688,In_1298,In_879);
nor U2689 (N_2689,In_1348,In_333);
nand U2690 (N_2690,In_19,In_214);
and U2691 (N_2691,In_246,In_1071);
xor U2692 (N_2692,In_592,In_1067);
or U2693 (N_2693,In_1269,In_1125);
nand U2694 (N_2694,In_144,In_875);
nand U2695 (N_2695,In_1298,In_1383);
xor U2696 (N_2696,In_809,In_1035);
xor U2697 (N_2697,In_421,In_1262);
nand U2698 (N_2698,In_623,In_1426);
xnor U2699 (N_2699,In_1023,In_1091);
or U2700 (N_2700,In_215,In_314);
xor U2701 (N_2701,In_1152,In_810);
xnor U2702 (N_2702,In_362,In_36);
nor U2703 (N_2703,In_571,In_1142);
xor U2704 (N_2704,In_931,In_730);
nand U2705 (N_2705,In_937,In_1118);
and U2706 (N_2706,In_252,In_886);
xor U2707 (N_2707,In_1287,In_394);
xnor U2708 (N_2708,In_545,In_472);
or U2709 (N_2709,In_959,In_113);
or U2710 (N_2710,In_714,In_1308);
or U2711 (N_2711,In_822,In_133);
and U2712 (N_2712,In_1366,In_512);
or U2713 (N_2713,In_326,In_950);
nor U2714 (N_2714,In_1418,In_1238);
nor U2715 (N_2715,In_1397,In_763);
xor U2716 (N_2716,In_1405,In_863);
and U2717 (N_2717,In_1103,In_478);
or U2718 (N_2718,In_954,In_542);
nand U2719 (N_2719,In_487,In_939);
nand U2720 (N_2720,In_1339,In_368);
xor U2721 (N_2721,In_193,In_525);
nor U2722 (N_2722,In_199,In_515);
nor U2723 (N_2723,In_943,In_613);
nor U2724 (N_2724,In_1447,In_825);
and U2725 (N_2725,In_112,In_680);
and U2726 (N_2726,In_567,In_1037);
xor U2727 (N_2727,In_1338,In_339);
and U2728 (N_2728,In_378,In_1074);
nor U2729 (N_2729,In_494,In_1083);
or U2730 (N_2730,In_1328,In_700);
nand U2731 (N_2731,In_1342,In_858);
nor U2732 (N_2732,In_1115,In_129);
and U2733 (N_2733,In_177,In_484);
nand U2734 (N_2734,In_1414,In_721);
nand U2735 (N_2735,In_174,In_817);
nand U2736 (N_2736,In_288,In_1347);
and U2737 (N_2737,In_799,In_654);
xnor U2738 (N_2738,In_925,In_437);
nor U2739 (N_2739,In_1141,In_949);
xnor U2740 (N_2740,In_47,In_837);
xor U2741 (N_2741,In_333,In_1375);
or U2742 (N_2742,In_915,In_629);
nor U2743 (N_2743,In_377,In_504);
and U2744 (N_2744,In_314,In_190);
and U2745 (N_2745,In_467,In_236);
xor U2746 (N_2746,In_1444,In_150);
or U2747 (N_2747,In_744,In_651);
xor U2748 (N_2748,In_560,In_584);
and U2749 (N_2749,In_1183,In_451);
nor U2750 (N_2750,In_622,In_519);
nand U2751 (N_2751,In_970,In_1057);
xnor U2752 (N_2752,In_478,In_1208);
nor U2753 (N_2753,In_1080,In_43);
and U2754 (N_2754,In_615,In_685);
nor U2755 (N_2755,In_1325,In_645);
and U2756 (N_2756,In_573,In_1010);
nand U2757 (N_2757,In_1159,In_364);
and U2758 (N_2758,In_192,In_289);
nor U2759 (N_2759,In_238,In_1382);
nand U2760 (N_2760,In_1102,In_171);
and U2761 (N_2761,In_777,In_799);
and U2762 (N_2762,In_779,In_1373);
or U2763 (N_2763,In_268,In_1380);
nand U2764 (N_2764,In_943,In_1462);
nand U2765 (N_2765,In_1400,In_933);
or U2766 (N_2766,In_473,In_1249);
nor U2767 (N_2767,In_137,In_46);
nand U2768 (N_2768,In_544,In_783);
nand U2769 (N_2769,In_742,In_888);
and U2770 (N_2770,In_1200,In_736);
nand U2771 (N_2771,In_612,In_1445);
and U2772 (N_2772,In_211,In_170);
and U2773 (N_2773,In_406,In_896);
nor U2774 (N_2774,In_785,In_1128);
nor U2775 (N_2775,In_985,In_407);
nand U2776 (N_2776,In_1480,In_67);
or U2777 (N_2777,In_1437,In_1051);
or U2778 (N_2778,In_1338,In_1357);
nor U2779 (N_2779,In_248,In_94);
nor U2780 (N_2780,In_501,In_410);
nor U2781 (N_2781,In_15,In_1226);
nor U2782 (N_2782,In_692,In_457);
or U2783 (N_2783,In_953,In_884);
nand U2784 (N_2784,In_344,In_937);
and U2785 (N_2785,In_1123,In_1178);
nor U2786 (N_2786,In_53,In_1276);
or U2787 (N_2787,In_1108,In_539);
xnor U2788 (N_2788,In_360,In_1106);
or U2789 (N_2789,In_937,In_1167);
or U2790 (N_2790,In_1144,In_283);
and U2791 (N_2791,In_542,In_614);
or U2792 (N_2792,In_1343,In_1226);
and U2793 (N_2793,In_1343,In_282);
nor U2794 (N_2794,In_378,In_833);
nand U2795 (N_2795,In_895,In_863);
xnor U2796 (N_2796,In_899,In_1128);
nor U2797 (N_2797,In_1155,In_667);
nor U2798 (N_2798,In_366,In_785);
nor U2799 (N_2799,In_945,In_481);
xnor U2800 (N_2800,In_1317,In_738);
xor U2801 (N_2801,In_154,In_155);
or U2802 (N_2802,In_1002,In_294);
nand U2803 (N_2803,In_405,In_487);
nor U2804 (N_2804,In_349,In_565);
and U2805 (N_2805,In_1297,In_351);
and U2806 (N_2806,In_748,In_1264);
and U2807 (N_2807,In_584,In_1338);
nor U2808 (N_2808,In_994,In_1228);
nand U2809 (N_2809,In_850,In_1432);
and U2810 (N_2810,In_1076,In_1261);
nand U2811 (N_2811,In_139,In_632);
or U2812 (N_2812,In_1439,In_821);
or U2813 (N_2813,In_534,In_1009);
xor U2814 (N_2814,In_438,In_72);
xnor U2815 (N_2815,In_1241,In_373);
xnor U2816 (N_2816,In_76,In_1318);
xnor U2817 (N_2817,In_930,In_180);
xnor U2818 (N_2818,In_334,In_608);
xnor U2819 (N_2819,In_835,In_1434);
and U2820 (N_2820,In_148,In_1012);
or U2821 (N_2821,In_130,In_1295);
and U2822 (N_2822,In_1392,In_416);
xnor U2823 (N_2823,In_572,In_379);
nor U2824 (N_2824,In_49,In_1258);
xnor U2825 (N_2825,In_69,In_87);
nor U2826 (N_2826,In_311,In_541);
nand U2827 (N_2827,In_27,In_1346);
and U2828 (N_2828,In_573,In_982);
or U2829 (N_2829,In_471,In_785);
xor U2830 (N_2830,In_615,In_911);
nand U2831 (N_2831,In_1238,In_1111);
nor U2832 (N_2832,In_966,In_447);
nor U2833 (N_2833,In_135,In_265);
xor U2834 (N_2834,In_764,In_1143);
or U2835 (N_2835,In_250,In_410);
nor U2836 (N_2836,In_463,In_434);
or U2837 (N_2837,In_1339,In_871);
and U2838 (N_2838,In_1284,In_608);
nor U2839 (N_2839,In_1376,In_1415);
xnor U2840 (N_2840,In_1032,In_3);
or U2841 (N_2841,In_1477,In_591);
xor U2842 (N_2842,In_1245,In_1325);
nor U2843 (N_2843,In_700,In_957);
or U2844 (N_2844,In_656,In_326);
and U2845 (N_2845,In_343,In_1180);
xnor U2846 (N_2846,In_485,In_80);
or U2847 (N_2847,In_263,In_373);
nor U2848 (N_2848,In_1431,In_468);
and U2849 (N_2849,In_1408,In_354);
xnor U2850 (N_2850,In_195,In_305);
xnor U2851 (N_2851,In_1471,In_748);
xnor U2852 (N_2852,In_343,In_1385);
or U2853 (N_2853,In_920,In_933);
nand U2854 (N_2854,In_1445,In_113);
or U2855 (N_2855,In_793,In_533);
nand U2856 (N_2856,In_1411,In_17);
or U2857 (N_2857,In_1427,In_92);
or U2858 (N_2858,In_1392,In_1322);
or U2859 (N_2859,In_410,In_194);
nor U2860 (N_2860,In_559,In_460);
nor U2861 (N_2861,In_79,In_48);
nand U2862 (N_2862,In_1224,In_1153);
nand U2863 (N_2863,In_812,In_362);
and U2864 (N_2864,In_1115,In_816);
and U2865 (N_2865,In_1120,In_1376);
or U2866 (N_2866,In_1409,In_782);
and U2867 (N_2867,In_633,In_916);
xor U2868 (N_2868,In_1223,In_132);
nor U2869 (N_2869,In_1044,In_1411);
and U2870 (N_2870,In_212,In_534);
and U2871 (N_2871,In_1268,In_1291);
xnor U2872 (N_2872,In_492,In_721);
and U2873 (N_2873,In_906,In_205);
nor U2874 (N_2874,In_568,In_1242);
xor U2875 (N_2875,In_736,In_654);
nor U2876 (N_2876,In_542,In_446);
xnor U2877 (N_2877,In_383,In_1479);
xnor U2878 (N_2878,In_1210,In_623);
xnor U2879 (N_2879,In_1331,In_143);
or U2880 (N_2880,In_379,In_832);
and U2881 (N_2881,In_1247,In_520);
nor U2882 (N_2882,In_1112,In_300);
nor U2883 (N_2883,In_260,In_182);
or U2884 (N_2884,In_235,In_190);
or U2885 (N_2885,In_1371,In_857);
and U2886 (N_2886,In_401,In_94);
or U2887 (N_2887,In_322,In_1110);
or U2888 (N_2888,In_1218,In_414);
or U2889 (N_2889,In_68,In_44);
nor U2890 (N_2890,In_200,In_1205);
nand U2891 (N_2891,In_1283,In_833);
nor U2892 (N_2892,In_1407,In_1400);
nor U2893 (N_2893,In_124,In_873);
or U2894 (N_2894,In_932,In_671);
nor U2895 (N_2895,In_206,In_692);
nand U2896 (N_2896,In_798,In_1298);
nor U2897 (N_2897,In_1271,In_313);
xnor U2898 (N_2898,In_467,In_898);
or U2899 (N_2899,In_569,In_1067);
or U2900 (N_2900,In_972,In_509);
nor U2901 (N_2901,In_115,In_613);
and U2902 (N_2902,In_1146,In_1461);
or U2903 (N_2903,In_147,In_119);
and U2904 (N_2904,In_448,In_1071);
xnor U2905 (N_2905,In_1161,In_455);
and U2906 (N_2906,In_1223,In_1138);
or U2907 (N_2907,In_1436,In_1447);
xor U2908 (N_2908,In_395,In_462);
nor U2909 (N_2909,In_754,In_1176);
and U2910 (N_2910,In_60,In_184);
and U2911 (N_2911,In_1411,In_107);
or U2912 (N_2912,In_628,In_197);
and U2913 (N_2913,In_546,In_1381);
and U2914 (N_2914,In_978,In_980);
nand U2915 (N_2915,In_69,In_520);
xnor U2916 (N_2916,In_1366,In_131);
nor U2917 (N_2917,In_663,In_195);
nor U2918 (N_2918,In_566,In_175);
or U2919 (N_2919,In_217,In_840);
xnor U2920 (N_2920,In_319,In_422);
nor U2921 (N_2921,In_504,In_973);
and U2922 (N_2922,In_1061,In_995);
nor U2923 (N_2923,In_950,In_1411);
and U2924 (N_2924,In_666,In_809);
nand U2925 (N_2925,In_1274,In_1215);
nand U2926 (N_2926,In_913,In_1148);
and U2927 (N_2927,In_1327,In_1105);
nor U2928 (N_2928,In_1169,In_678);
nor U2929 (N_2929,In_1278,In_1057);
xor U2930 (N_2930,In_388,In_586);
and U2931 (N_2931,In_958,In_61);
nand U2932 (N_2932,In_798,In_59);
and U2933 (N_2933,In_196,In_511);
or U2934 (N_2934,In_709,In_614);
nand U2935 (N_2935,In_674,In_829);
and U2936 (N_2936,In_319,In_99);
and U2937 (N_2937,In_771,In_598);
and U2938 (N_2938,In_23,In_1086);
nor U2939 (N_2939,In_431,In_1257);
and U2940 (N_2940,In_1130,In_1217);
nor U2941 (N_2941,In_115,In_1035);
or U2942 (N_2942,In_676,In_764);
xnor U2943 (N_2943,In_1082,In_638);
xnor U2944 (N_2944,In_951,In_519);
or U2945 (N_2945,In_681,In_406);
xor U2946 (N_2946,In_613,In_326);
xor U2947 (N_2947,In_711,In_441);
or U2948 (N_2948,In_530,In_1146);
or U2949 (N_2949,In_513,In_113);
and U2950 (N_2950,In_1275,In_315);
or U2951 (N_2951,In_1405,In_101);
xnor U2952 (N_2952,In_1353,In_1094);
xnor U2953 (N_2953,In_211,In_137);
nand U2954 (N_2954,In_201,In_484);
and U2955 (N_2955,In_706,In_872);
xnor U2956 (N_2956,In_627,In_1278);
and U2957 (N_2957,In_1100,In_544);
nor U2958 (N_2958,In_1261,In_214);
xor U2959 (N_2959,In_1436,In_1187);
nand U2960 (N_2960,In_1297,In_169);
nor U2961 (N_2961,In_866,In_415);
or U2962 (N_2962,In_457,In_378);
xnor U2963 (N_2963,In_1290,In_321);
or U2964 (N_2964,In_529,In_1467);
nor U2965 (N_2965,In_941,In_803);
nor U2966 (N_2966,In_1049,In_28);
nand U2967 (N_2967,In_1203,In_1247);
or U2968 (N_2968,In_338,In_573);
and U2969 (N_2969,In_1346,In_108);
xor U2970 (N_2970,In_1331,In_796);
and U2971 (N_2971,In_465,In_1462);
and U2972 (N_2972,In_87,In_1361);
or U2973 (N_2973,In_494,In_386);
nor U2974 (N_2974,In_164,In_965);
nand U2975 (N_2975,In_672,In_215);
or U2976 (N_2976,In_74,In_679);
and U2977 (N_2977,In_193,In_699);
nand U2978 (N_2978,In_1043,In_390);
nand U2979 (N_2979,In_924,In_686);
nor U2980 (N_2980,In_451,In_546);
xnor U2981 (N_2981,In_136,In_959);
xnor U2982 (N_2982,In_499,In_124);
xor U2983 (N_2983,In_257,In_408);
and U2984 (N_2984,In_1363,In_791);
and U2985 (N_2985,In_1201,In_863);
nand U2986 (N_2986,In_1497,In_222);
nand U2987 (N_2987,In_699,In_732);
nor U2988 (N_2988,In_77,In_1144);
and U2989 (N_2989,In_245,In_752);
or U2990 (N_2990,In_946,In_336);
xnor U2991 (N_2991,In_1344,In_1249);
xnor U2992 (N_2992,In_631,In_969);
xnor U2993 (N_2993,In_197,In_393);
and U2994 (N_2994,In_678,In_201);
xor U2995 (N_2995,In_492,In_760);
or U2996 (N_2996,In_943,In_294);
xor U2997 (N_2997,In_1377,In_431);
and U2998 (N_2998,In_772,In_441);
or U2999 (N_2999,In_842,In_1306);
or U3000 (N_3000,N_107,N_2388);
nand U3001 (N_3001,N_1560,N_1702);
and U3002 (N_3002,N_2766,N_2896);
and U3003 (N_3003,N_1191,N_1917);
or U3004 (N_3004,N_766,N_2994);
or U3005 (N_3005,N_1641,N_81);
nor U3006 (N_3006,N_205,N_968);
and U3007 (N_3007,N_1382,N_2007);
or U3008 (N_3008,N_2708,N_488);
xnor U3009 (N_3009,N_2082,N_2436);
nor U3010 (N_3010,N_1777,N_178);
nor U3011 (N_3011,N_1350,N_2386);
xor U3012 (N_3012,N_1930,N_1646);
and U3013 (N_3013,N_1345,N_2130);
nor U3014 (N_3014,N_1750,N_1054);
nor U3015 (N_3015,N_2963,N_2264);
nand U3016 (N_3016,N_1062,N_275);
nor U3017 (N_3017,N_1261,N_670);
xnor U3018 (N_3018,N_2794,N_1996);
and U3019 (N_3019,N_191,N_2441);
xnor U3020 (N_3020,N_2735,N_1706);
or U3021 (N_3021,N_2623,N_285);
nand U3022 (N_3022,N_2062,N_2661);
or U3023 (N_3023,N_1774,N_1419);
nand U3024 (N_3024,N_491,N_610);
and U3025 (N_3025,N_1763,N_2779);
and U3026 (N_3026,N_2087,N_1584);
or U3027 (N_3027,N_459,N_522);
nor U3028 (N_3028,N_588,N_2822);
xor U3029 (N_3029,N_224,N_2685);
xnor U3030 (N_3030,N_1070,N_739);
and U3031 (N_3031,N_1950,N_370);
nor U3032 (N_3032,N_1301,N_152);
xor U3033 (N_3033,N_1211,N_302);
nor U3034 (N_3034,N_953,N_2450);
nand U3035 (N_3035,N_2621,N_111);
nor U3036 (N_3036,N_2048,N_2391);
nor U3037 (N_3037,N_2194,N_2959);
nand U3038 (N_3038,N_2868,N_1632);
or U3039 (N_3039,N_1764,N_1119);
nor U3040 (N_3040,N_166,N_1146);
or U3041 (N_3041,N_2298,N_1431);
xnor U3042 (N_3042,N_733,N_2714);
nand U3043 (N_3043,N_142,N_554);
or U3044 (N_3044,N_2697,N_2080);
or U3045 (N_3045,N_497,N_305);
nor U3046 (N_3046,N_2049,N_2282);
xor U3047 (N_3047,N_2244,N_2395);
nor U3048 (N_3048,N_852,N_1615);
and U3049 (N_3049,N_403,N_1708);
nor U3050 (N_3050,N_223,N_25);
nand U3051 (N_3051,N_2478,N_2227);
nor U3052 (N_3052,N_635,N_2625);
nor U3053 (N_3053,N_2104,N_425);
and U3054 (N_3054,N_1694,N_1246);
xor U3055 (N_3055,N_263,N_1056);
nand U3056 (N_3056,N_432,N_1843);
or U3057 (N_3057,N_2144,N_2635);
xor U3058 (N_3058,N_1459,N_225);
or U3059 (N_3059,N_331,N_335);
or U3060 (N_3060,N_2040,N_2549);
xor U3061 (N_3061,N_1289,N_2502);
xnor U3062 (N_3062,N_723,N_2129);
nor U3063 (N_3063,N_1883,N_2153);
xor U3064 (N_3064,N_311,N_385);
nand U3065 (N_3065,N_2469,N_580);
nand U3066 (N_3066,N_64,N_1300);
nand U3067 (N_3067,N_313,N_82);
or U3068 (N_3068,N_2182,N_1287);
nor U3069 (N_3069,N_1791,N_552);
xnor U3070 (N_3070,N_2446,N_1753);
nand U3071 (N_3071,N_1463,N_2921);
nand U3072 (N_3072,N_1011,N_898);
xnor U3073 (N_3073,N_2791,N_2204);
xor U3074 (N_3074,N_1554,N_1666);
nand U3075 (N_3075,N_653,N_1609);
nor U3076 (N_3076,N_2232,N_833);
or U3077 (N_3077,N_2060,N_2727);
nand U3078 (N_3078,N_493,N_637);
nor U3079 (N_3079,N_79,N_1675);
nand U3080 (N_3080,N_1597,N_787);
nand U3081 (N_3081,N_603,N_557);
xnor U3082 (N_3082,N_2366,N_394);
or U3083 (N_3083,N_1735,N_924);
or U3084 (N_3084,N_238,N_2190);
nor U3085 (N_3085,N_1716,N_2657);
or U3086 (N_3086,N_1681,N_1712);
nor U3087 (N_3087,N_727,N_1826);
nand U3088 (N_3088,N_375,N_2793);
nor U3089 (N_3089,N_2590,N_1687);
and U3090 (N_3090,N_874,N_1749);
nand U3091 (N_3091,N_805,N_424);
nor U3092 (N_3092,N_276,N_2234);
and U3093 (N_3093,N_1730,N_500);
xor U3094 (N_3094,N_1332,N_803);
nor U3095 (N_3095,N_1538,N_1649);
nand U3096 (N_3096,N_2103,N_1668);
and U3097 (N_3097,N_2715,N_2169);
and U3098 (N_3098,N_807,N_190);
nor U3099 (N_3099,N_1890,N_1860);
xnor U3100 (N_3100,N_1150,N_2583);
nor U3101 (N_3101,N_95,N_2967);
nor U3102 (N_3102,N_1206,N_1804);
nor U3103 (N_3103,N_2856,N_2663);
nand U3104 (N_3104,N_1500,N_1734);
nand U3105 (N_3105,N_2954,N_2081);
nand U3106 (N_3106,N_2909,N_369);
xnor U3107 (N_3107,N_886,N_1907);
or U3108 (N_3108,N_2420,N_33);
and U3109 (N_3109,N_2317,N_1628);
nand U3110 (N_3110,N_686,N_2164);
and U3111 (N_3111,N_353,N_1693);
xor U3112 (N_3112,N_1293,N_2730);
nor U3113 (N_3113,N_2464,N_980);
xnor U3114 (N_3114,N_986,N_1648);
or U3115 (N_3115,N_1717,N_157);
nand U3116 (N_3116,N_2107,N_464);
xnor U3117 (N_3117,N_1812,N_136);
xor U3118 (N_3118,N_88,N_1178);
nor U3119 (N_3119,N_2574,N_1933);
and U3120 (N_3120,N_2326,N_2415);
nand U3121 (N_3121,N_330,N_673);
nand U3122 (N_3122,N_1509,N_2167);
nand U3123 (N_3123,N_729,N_761);
nand U3124 (N_3124,N_1444,N_2154);
nor U3125 (N_3125,N_1400,N_2515);
xor U3126 (N_3126,N_565,N_211);
nand U3127 (N_3127,N_2068,N_1082);
nand U3128 (N_3128,N_719,N_2545);
nand U3129 (N_3129,N_2218,N_606);
xor U3130 (N_3130,N_2397,N_1691);
and U3131 (N_3131,N_625,N_2680);
and U3132 (N_3132,N_608,N_520);
and U3133 (N_3133,N_1469,N_1193);
xnor U3134 (N_3134,N_154,N_2548);
and U3135 (N_3135,N_2764,N_546);
or U3136 (N_3136,N_273,N_1553);
nand U3137 (N_3137,N_14,N_1532);
nor U3138 (N_3138,N_869,N_1661);
xnor U3139 (N_3139,N_2944,N_586);
nand U3140 (N_3140,N_1778,N_204);
nor U3141 (N_3141,N_1346,N_2600);
or U3142 (N_3142,N_2166,N_881);
nor U3143 (N_3143,N_2102,N_1829);
and U3144 (N_3144,N_2782,N_519);
xor U3145 (N_3145,N_663,N_1428);
xnor U3146 (N_3146,N_2393,N_2656);
and U3147 (N_3147,N_1481,N_1026);
nor U3148 (N_3148,N_1058,N_75);
and U3149 (N_3149,N_133,N_195);
xnor U3150 (N_3150,N_1231,N_1226);
and U3151 (N_3151,N_530,N_471);
or U3152 (N_3152,N_1028,N_2615);
and U3153 (N_3153,N_1363,N_2830);
or U3154 (N_3154,N_1336,N_438);
or U3155 (N_3155,N_2936,N_993);
and U3156 (N_3156,N_2212,N_1517);
nand U3157 (N_3157,N_2297,N_2271);
or U3158 (N_3158,N_202,N_443);
xnor U3159 (N_3159,N_1063,N_2767);
and U3160 (N_3160,N_1898,N_507);
nor U3161 (N_3161,N_36,N_850);
nand U3162 (N_3162,N_2845,N_2920);
or U3163 (N_3163,N_1789,N_2706);
nor U3164 (N_3164,N_710,N_1700);
nand U3165 (N_3165,N_243,N_357);
or U3166 (N_3166,N_925,N_1832);
nand U3167 (N_3167,N_220,N_802);
xor U3168 (N_3168,N_640,N_2185);
nand U3169 (N_3169,N_1470,N_2718);
nand U3170 (N_3170,N_288,N_1551);
xnor U3171 (N_3171,N_102,N_1227);
nor U3172 (N_3172,N_2105,N_1850);
xor U3173 (N_3173,N_96,N_2756);
nand U3174 (N_3174,N_2044,N_1217);
xnor U3175 (N_3175,N_1592,N_728);
and U3176 (N_3176,N_1258,N_1698);
xnor U3177 (N_3177,N_560,N_1642);
nor U3178 (N_3178,N_2527,N_829);
and U3179 (N_3179,N_1266,N_2965);
or U3180 (N_3180,N_696,N_1415);
nand U3181 (N_3181,N_1928,N_1674);
and U3182 (N_3182,N_215,N_2310);
or U3183 (N_3183,N_1130,N_1160);
nand U3184 (N_3184,N_2681,N_1203);
and U3185 (N_3185,N_1034,N_899);
nor U3186 (N_3186,N_2260,N_1680);
nand U3187 (N_3187,N_2351,N_1233);
nand U3188 (N_3188,N_617,N_917);
xor U3189 (N_3189,N_1934,N_1887);
or U3190 (N_3190,N_2400,N_2698);
xor U3191 (N_3191,N_892,N_253);
or U3192 (N_3192,N_592,N_1079);
nor U3193 (N_3193,N_322,N_2783);
xor U3194 (N_3194,N_319,N_1873);
nand U3195 (N_3195,N_421,N_1904);
or U3196 (N_3196,N_992,N_244);
nor U3197 (N_3197,N_1100,N_404);
or U3198 (N_3198,N_938,N_2544);
nor U3199 (N_3199,N_2795,N_2307);
or U3200 (N_3200,N_1645,N_361);
nor U3201 (N_3201,N_159,N_1484);
or U3202 (N_3202,N_2359,N_181);
or U3203 (N_3203,N_2461,N_314);
xnor U3204 (N_3204,N_1068,N_631);
nor U3205 (N_3205,N_1557,N_1651);
xor U3206 (N_3206,N_689,N_2753);
and U3207 (N_3207,N_78,N_2966);
xnor U3208 (N_3208,N_613,N_1920);
nor U3209 (N_3209,N_1433,N_1085);
and U3210 (N_3210,N_2134,N_2242);
and U3211 (N_3211,N_1663,N_336);
or U3212 (N_3212,N_1072,N_1434);
nor U3213 (N_3213,N_1073,N_2976);
and U3214 (N_3214,N_1783,N_66);
nand U3215 (N_3215,N_2928,N_1099);
xnor U3216 (N_3216,N_571,N_619);
or U3217 (N_3217,N_1071,N_650);
and U3218 (N_3218,N_68,N_1868);
nand U3219 (N_3219,N_490,N_2065);
nand U3220 (N_3220,N_564,N_423);
xor U3221 (N_3221,N_1869,N_1991);
nor U3222 (N_3222,N_71,N_446);
or U3223 (N_3223,N_356,N_2488);
xor U3224 (N_3224,N_2693,N_2286);
or U3225 (N_3225,N_648,N_1733);
xor U3226 (N_3226,N_307,N_2025);
nor U3227 (N_3227,N_405,N_2611);
nand U3228 (N_3228,N_1775,N_2061);
or U3229 (N_3229,N_641,N_1480);
and U3230 (N_3230,N_2946,N_168);
and U3231 (N_3231,N_1000,N_2970);
nand U3232 (N_3232,N_2018,N_1477);
nor U3233 (N_3233,N_1205,N_376);
nor U3234 (N_3234,N_1264,N_651);
and U3235 (N_3235,N_827,N_1851);
or U3236 (N_3236,N_1214,N_652);
or U3237 (N_3237,N_2943,N_1170);
or U3238 (N_3238,N_1813,N_2823);
nor U3239 (N_3239,N_1183,N_2803);
xor U3240 (N_3240,N_753,N_2224);
nand U3241 (N_3241,N_902,N_1420);
nor U3242 (N_3242,N_2832,N_2014);
xor U3243 (N_3243,N_1485,N_2734);
xor U3244 (N_3244,N_2883,N_1252);
nand U3245 (N_3245,N_2669,N_2792);
xor U3246 (N_3246,N_2809,N_2159);
nand U3247 (N_3247,N_2305,N_861);
nand U3248 (N_3248,N_1269,N_2724);
and U3249 (N_3249,N_1357,N_1726);
nor U3250 (N_3250,N_1508,N_1089);
or U3251 (N_3251,N_374,N_2926);
or U3252 (N_3252,N_1547,N_1952);
nor U3253 (N_3253,N_1937,N_2489);
or U3254 (N_3254,N_1187,N_2449);
nor U3255 (N_3255,N_2263,N_2231);
and U3256 (N_3256,N_1616,N_1552);
nand U3257 (N_3257,N_834,N_2591);
and U3258 (N_3258,N_2438,N_1326);
nor U3259 (N_3259,N_2220,N_523);
nand U3260 (N_3260,N_1656,N_513);
nand U3261 (N_3261,N_2587,N_939);
nand U3262 (N_3262,N_1916,N_2160);
and U3263 (N_3263,N_1044,N_2655);
nor U3264 (N_3264,N_627,N_2406);
xor U3265 (N_3265,N_2041,N_1882);
xnor U3266 (N_3266,N_2240,N_2373);
xor U3267 (N_3267,N_2662,N_108);
nor U3268 (N_3268,N_2408,N_2844);
nand U3269 (N_3269,N_1334,N_2606);
xnor U3270 (N_3270,N_2914,N_105);
nand U3271 (N_3271,N_2002,N_442);
xor U3272 (N_3272,N_1565,N_352);
and U3273 (N_3273,N_515,N_873);
nand U3274 (N_3274,N_903,N_1247);
nand U3275 (N_3275,N_2091,N_2020);
xor U3276 (N_3276,N_1241,N_1834);
nand U3277 (N_3277,N_1751,N_1257);
and U3278 (N_3278,N_1384,N_866);
and U3279 (N_3279,N_846,N_1229);
nor U3280 (N_3280,N_2175,N_2618);
nand U3281 (N_3281,N_2195,N_2075);
or U3282 (N_3282,N_505,N_1412);
nand U3283 (N_3283,N_1474,N_1047);
xnor U3284 (N_3284,N_1958,N_1291);
nor U3285 (N_3285,N_851,N_2992);
nand U3286 (N_3286,N_98,N_2911);
xor U3287 (N_3287,N_45,N_414);
or U3288 (N_3288,N_2180,N_137);
nor U3289 (N_3289,N_1926,N_1002);
nand U3290 (N_3290,N_2362,N_662);
nor U3291 (N_3291,N_2751,N_2287);
nand U3292 (N_3292,N_1243,N_452);
or U3293 (N_3293,N_2624,N_844);
and U3294 (N_3294,N_1960,N_1600);
xnor U3295 (N_3295,N_2897,N_841);
and U3296 (N_3296,N_2146,N_2165);
or U3297 (N_3297,N_1133,N_1055);
or U3298 (N_3298,N_1817,N_2906);
and U3299 (N_3299,N_822,N_741);
nand U3300 (N_3300,N_758,N_2427);
and U3301 (N_3301,N_2045,N_1006);
nor U3302 (N_3302,N_2499,N_717);
xnor U3303 (N_3303,N_130,N_309);
nand U3304 (N_3304,N_266,N_919);
nor U3305 (N_3305,N_1719,N_1152);
nand U3306 (N_3306,N_1936,N_975);
nor U3307 (N_3307,N_1493,N_2721);
and U3308 (N_3308,N_2026,N_1237);
nor U3309 (N_3309,N_1440,N_1727);
nor U3310 (N_3310,N_1259,N_735);
nor U3311 (N_3311,N_745,N_2719);
or U3312 (N_3312,N_1115,N_561);
or U3313 (N_3313,N_1541,N_1081);
and U3314 (N_3314,N_2426,N_2016);
or U3315 (N_3315,N_2859,N_173);
nand U3316 (N_3316,N_2733,N_2202);
or U3317 (N_3317,N_2673,N_1114);
nor U3318 (N_3318,N_1242,N_1841);
nand U3319 (N_3319,N_2999,N_1889);
nor U3320 (N_3320,N_1871,N_660);
nor U3321 (N_3321,N_1808,N_76);
nor U3322 (N_3322,N_2984,N_1931);
nor U3323 (N_3323,N_770,N_407);
xor U3324 (N_3324,N_2831,N_790);
xor U3325 (N_3325,N_1947,N_528);
nand U3326 (N_3326,N_611,N_2369);
and U3327 (N_3327,N_2017,N_1109);
xor U3328 (N_3328,N_1207,N_2122);
xnor U3329 (N_3329,N_575,N_2875);
or U3330 (N_3330,N_1184,N_1894);
xor U3331 (N_3331,N_2565,N_2505);
nand U3332 (N_3332,N_887,N_2757);
and U3333 (N_3333,N_2895,N_103);
nor U3334 (N_3334,N_1980,N_77);
or U3335 (N_3335,N_2935,N_1340);
xnor U3336 (N_3336,N_2410,N_2463);
or U3337 (N_3337,N_2742,N_2035);
and U3338 (N_3338,N_2932,N_1491);
and U3339 (N_3339,N_1131,N_579);
nor U3340 (N_3340,N_2686,N_93);
and U3341 (N_3341,N_888,N_2414);
xor U3342 (N_3342,N_2986,N_2381);
nor U3343 (N_3343,N_1588,N_2781);
nand U3344 (N_3344,N_1280,N_487);
and U3345 (N_3345,N_1250,N_462);
and U3346 (N_3346,N_2891,N_1769);
nor U3347 (N_3347,N_1310,N_772);
or U3348 (N_3348,N_657,N_2024);
nand U3349 (N_3349,N_988,N_2128);
or U3350 (N_3350,N_2700,N_1720);
nor U3351 (N_3351,N_2550,N_448);
and U3352 (N_3352,N_249,N_1323);
nor U3353 (N_3353,N_1424,N_985);
nand U3354 (N_3354,N_1041,N_1782);
and U3355 (N_3355,N_1807,N_2535);
or U3356 (N_3356,N_1244,N_1507);
or U3357 (N_3357,N_502,N_984);
or U3358 (N_3358,N_412,N_1288);
and U3359 (N_3359,N_2849,N_2953);
nor U3360 (N_3360,N_726,N_2323);
xor U3361 (N_3361,N_6,N_2829);
nand U3362 (N_3362,N_1267,N_135);
xor U3363 (N_3363,N_1624,N_478);
xnor U3364 (N_3364,N_1910,N_1189);
or U3365 (N_3365,N_2632,N_1969);
or U3366 (N_3366,N_1144,N_114);
xnor U3367 (N_3367,N_1134,N_1274);
nand U3368 (N_3368,N_1155,N_1248);
or U3369 (N_3369,N_675,N_649);
and U3370 (N_3370,N_282,N_1);
nand U3371 (N_3371,N_2701,N_2892);
xor U3372 (N_3372,N_2133,N_1398);
nor U3373 (N_3373,N_2452,N_2855);
nand U3374 (N_3374,N_1251,N_1505);
nand U3375 (N_3375,N_1810,N_1486);
and U3376 (N_3376,N_2008,N_2413);
nor U3377 (N_3377,N_540,N_476);
or U3378 (N_3378,N_1621,N_2726);
or U3379 (N_3379,N_2346,N_171);
nand U3380 (N_3380,N_2846,N_2274);
and U3381 (N_3381,N_1408,N_16);
or U3382 (N_3382,N_935,N_2585);
nand U3383 (N_3383,N_1643,N_1526);
xnor U3384 (N_3384,N_1136,N_239);
xor U3385 (N_3385,N_1620,N_158);
and U3386 (N_3386,N_2786,N_473);
xnor U3387 (N_3387,N_666,N_308);
and U3388 (N_3388,N_2775,N_566);
xnor U3389 (N_3389,N_961,N_2930);
nand U3390 (N_3390,N_708,N_1515);
nand U3391 (N_3391,N_2631,N_2399);
and U3392 (N_3392,N_2857,N_2329);
nand U3393 (N_3393,N_2266,N_2760);
xor U3394 (N_3394,N_2815,N_1306);
xor U3395 (N_3395,N_929,N_1862);
nand U3396 (N_3396,N_569,N_1221);
xor U3397 (N_3397,N_2155,N_1043);
and U3398 (N_3398,N_2094,N_2233);
xor U3399 (N_3399,N_1617,N_1447);
nand U3400 (N_3400,N_2496,N_2084);
xor U3401 (N_3401,N_918,N_2302);
nor U3402 (N_3402,N_2058,N_2258);
xnor U3403 (N_3403,N_1723,N_2711);
nand U3404 (N_3404,N_2501,N_954);
and U3405 (N_3405,N_2684,N_1017);
or U3406 (N_3406,N_2610,N_541);
nand U3407 (N_3407,N_2731,N_1356);
xor U3408 (N_3408,N_52,N_2525);
nor U3409 (N_3409,N_2428,N_2006);
and U3410 (N_3410,N_2720,N_58);
nand U3411 (N_3411,N_2113,N_1536);
nor U3412 (N_3412,N_2125,N_1224);
nand U3413 (N_3413,N_1732,N_1478);
and U3414 (N_3414,N_609,N_2116);
xor U3415 (N_3415,N_843,N_1741);
nand U3416 (N_3416,N_325,N_2604);
nor U3417 (N_3417,N_773,N_2230);
nand U3418 (N_3418,N_2772,N_1878);
nor U3419 (N_3419,N_691,N_1570);
and U3420 (N_3420,N_1204,N_684);
and U3421 (N_3421,N_2495,N_879);
or U3422 (N_3422,N_1040,N_2931);
and U3423 (N_3423,N_437,N_1467);
nor U3424 (N_3424,N_781,N_1697);
and U3425 (N_3425,N_1956,N_2658);
xnor U3426 (N_3426,N_2380,N_470);
nor U3427 (N_3427,N_864,N_1057);
xnor U3428 (N_3428,N_1093,N_1742);
and U3429 (N_3429,N_607,N_2046);
and U3430 (N_3430,N_199,N_1030);
nand U3431 (N_3431,N_2197,N_1436);
or U3432 (N_3432,N_2272,N_50);
or U3433 (N_3433,N_2101,N_237);
and U3434 (N_3434,N_667,N_1128);
and U3435 (N_3435,N_408,N_2352);
xor U3436 (N_3436,N_1149,N_1003);
nand U3437 (N_3437,N_1086,N_2279);
nor U3438 (N_3438,N_1831,N_2597);
and U3439 (N_3439,N_489,N_2561);
or U3440 (N_3440,N_164,N_2392);
or U3441 (N_3441,N_655,N_2995);
or U3442 (N_3442,N_2177,N_1853);
nand U3443 (N_3443,N_326,N_836);
nor U3444 (N_3444,N_1035,N_2411);
xor U3445 (N_3445,N_1285,N_186);
nor U3446 (N_3446,N_1122,N_1074);
and U3447 (N_3447,N_1858,N_1501);
xnor U3448 (N_3448,N_2667,N_894);
xor U3449 (N_3449,N_2531,N_2801);
and U3450 (N_3450,N_1094,N_390);
and U3451 (N_3451,N_2213,N_989);
xnor U3452 (N_3452,N_121,N_2385);
xor U3453 (N_3453,N_299,N_38);
xnor U3454 (N_3454,N_257,N_616);
or U3455 (N_3455,N_669,N_2072);
or U3456 (N_3456,N_2148,N_333);
xor U3457 (N_3457,N_2509,N_2957);
nor U3458 (N_3458,N_2481,N_2334);
nand U3459 (N_3459,N_1245,N_1613);
or U3460 (N_3460,N_2763,N_1176);
nand U3461 (N_3461,N_44,N_2870);
nand U3462 (N_3462,N_392,N_647);
xor U3463 (N_3463,N_659,N_1967);
xnor U3464 (N_3464,N_1512,N_2762);
nand U3465 (N_3465,N_1390,N_1069);
xnor U3466 (N_3466,N_2372,N_1090);
nor U3467 (N_3467,N_1612,N_1962);
nand U3468 (N_3468,N_596,N_454);
or U3469 (N_3469,N_884,N_1548);
and U3470 (N_3470,N_116,N_2314);
or U3471 (N_3471,N_1163,N_1239);
or U3472 (N_3472,N_2540,N_144);
nand U3473 (N_3473,N_747,N_567);
nand U3474 (N_3474,N_1985,N_2908);
nor U3475 (N_3475,N_2512,N_1429);
nand U3476 (N_3476,N_399,N_2412);
and U3477 (N_3477,N_2884,N_1562);
xnor U3478 (N_3478,N_2788,N_2135);
or U3479 (N_3479,N_973,N_1833);
and U3480 (N_3480,N_2066,N_923);
nor U3481 (N_3481,N_1328,N_122);
nor U3482 (N_3482,N_1514,N_24);
xor U3483 (N_3483,N_1254,N_2969);
and U3484 (N_3484,N_1608,N_581);
xnor U3485 (N_3485,N_909,N_345);
xor U3486 (N_3486,N_2047,N_1837);
xor U3487 (N_3487,N_2704,N_42);
nor U3488 (N_3488,N_624,N_937);
nor U3489 (N_3489,N_548,N_1208);
or U3490 (N_3490,N_2207,N_1836);
nor U3491 (N_3491,N_538,N_1430);
nand U3492 (N_3492,N_143,N_1886);
xor U3493 (N_3493,N_172,N_831);
xnor U3494 (N_3494,N_636,N_54);
and U3495 (N_3495,N_1315,N_683);
or U3496 (N_3496,N_1915,N_2192);
nand U3497 (N_3497,N_896,N_1001);
nand U3498 (N_3498,N_2250,N_1728);
xor U3499 (N_3499,N_1510,N_1249);
nor U3500 (N_3500,N_2813,N_509);
nand U3501 (N_3501,N_1036,N_1308);
and U3502 (N_3502,N_1238,N_1335);
xor U3503 (N_3503,N_1135,N_977);
nand U3504 (N_3504,N_2929,N_1758);
or U3505 (N_3505,N_828,N_915);
or U3506 (N_3506,N_1321,N_1032);
or U3507 (N_3507,N_1260,N_2745);
xor U3508 (N_3508,N_486,N_304);
and U3509 (N_3509,N_101,N_2665);
nand U3510 (N_3510,N_676,N_1604);
nor U3511 (N_3511,N_1295,N_100);
nand U3512 (N_3512,N_177,N_2402);
nor U3513 (N_3513,N_2443,N_832);
xor U3514 (N_3514,N_2176,N_2467);
xor U3515 (N_3515,N_1979,N_913);
nor U3516 (N_3516,N_1639,N_731);
nor U3517 (N_3517,N_300,N_1669);
or U3518 (N_3518,N_722,N_284);
and U3519 (N_3519,N_1696,N_1685);
nand U3520 (N_3520,N_2879,N_495);
and U3521 (N_3521,N_2522,N_2653);
nor U3522 (N_3522,N_928,N_387);
or U3523 (N_3523,N_1992,N_1194);
or U3524 (N_3524,N_2578,N_1296);
xnor U3525 (N_3525,N_1881,N_1633);
nand U3526 (N_3526,N_1722,N_583);
and U3527 (N_3527,N_26,N_1626);
or U3528 (N_3528,N_2073,N_643);
xnor U3529 (N_3529,N_1162,N_472);
xor U3530 (N_3530,N_1531,N_457);
xnor U3531 (N_3531,N_1954,N_2120);
and U3532 (N_3532,N_665,N_2249);
or U3533 (N_3533,N_2405,N_931);
xor U3534 (N_3534,N_890,N_499);
nand U3535 (N_3535,N_574,N_524);
and U3536 (N_3536,N_576,N_946);
nor U3537 (N_3537,N_1603,N_534);
nor U3538 (N_3538,N_2695,N_1282);
nor U3539 (N_3539,N_2437,N_2077);
nand U3540 (N_3540,N_1797,N_274);
and U3541 (N_3541,N_1983,N_328);
nand U3542 (N_3542,N_431,N_123);
xor U3543 (N_3543,N_5,N_794);
and U3544 (N_3544,N_1012,N_1004);
nand U3545 (N_3545,N_2818,N_1273);
nand U3546 (N_3546,N_2215,N_1066);
xnor U3547 (N_3547,N_1550,N_1815);
or U3548 (N_3548,N_342,N_740);
nand U3549 (N_3549,N_184,N_1294);
nand U3550 (N_3550,N_1145,N_2200);
or U3551 (N_3551,N_1401,N_1380);
nand U3552 (N_3552,N_703,N_2376);
nor U3553 (N_3553,N_2296,N_465);
or U3554 (N_3554,N_1676,N_1840);
nor U3555 (N_3555,N_222,N_2354);
or U3556 (N_3556,N_1213,N_533);
xor U3557 (N_3557,N_767,N_0);
xor U3558 (N_3558,N_2293,N_2542);
nand U3559 (N_3559,N_549,N_1938);
and U3560 (N_3560,N_746,N_2338);
nand U3561 (N_3561,N_1766,N_1405);
xnor U3562 (N_3562,N_1761,N_878);
nand U3563 (N_3563,N_1468,N_131);
or U3564 (N_3564,N_53,N_1818);
xnor U3565 (N_3565,N_1499,N_1579);
xnor U3566 (N_3566,N_628,N_900);
and U3567 (N_3567,N_2814,N_1416);
or U3568 (N_3568,N_39,N_558);
xnor U3569 (N_3569,N_511,N_2841);
and U3570 (N_3570,N_814,N_2033);
nand U3571 (N_3571,N_1046,N_2517);
or U3572 (N_3572,N_2268,N_1684);
xnor U3573 (N_3573,N_504,N_1594);
nor U3574 (N_3574,N_2728,N_2993);
xnor U3575 (N_3575,N_2511,N_388);
nand U3576 (N_3576,N_287,N_1729);
or U3577 (N_3577,N_1835,N_1494);
nand U3578 (N_3578,N_820,N_2012);
and U3579 (N_3579,N_73,N_780);
or U3580 (N_3580,N_2915,N_1361);
nor U3581 (N_3581,N_1568,N_1098);
xor U3582 (N_3582,N_15,N_1080);
xor U3583 (N_3583,N_1895,N_344);
nor U3584 (N_3584,N_1688,N_2447);
nand U3585 (N_3585,N_1638,N_296);
and U3586 (N_3586,N_455,N_1619);
nand U3587 (N_3587,N_1116,N_2960);
or U3588 (N_3588,N_1359,N_1051);
or U3589 (N_3589,N_2171,N_2407);
nand U3590 (N_3590,N_1234,N_1496);
nand U3591 (N_3591,N_2643,N_1175);
and U3592 (N_3592,N_1460,N_2722);
xnor U3593 (N_3593,N_1718,N_216);
nor U3594 (N_3594,N_2005,N_30);
and U3595 (N_3595,N_1138,N_2032);
xor U3596 (N_3596,N_1352,N_1795);
nand U3597 (N_3597,N_170,N_1759);
and U3598 (N_3598,N_1112,N_970);
and U3599 (N_3599,N_1622,N_2445);
and U3600 (N_3600,N_2785,N_2123);
nor U3601 (N_3601,N_2161,N_867);
and U3602 (N_3602,N_2255,N_1378);
nand U3603 (N_3603,N_933,N_2790);
nand U3604 (N_3604,N_227,N_1385);
nor U3605 (N_3605,N_1892,N_364);
nand U3606 (N_3606,N_2773,N_1577);
xnor U3607 (N_3607,N_2628,N_2530);
nand U3608 (N_3608,N_1545,N_1441);
nor U3609 (N_3609,N_2339,N_229);
nand U3610 (N_3610,N_230,N_2894);
nand U3611 (N_3611,N_1998,N_2483);
and U3612 (N_3612,N_2537,N_1374);
nor U3613 (N_3613,N_2682,N_1566);
nor U3614 (N_3614,N_2217,N_1773);
or U3615 (N_3615,N_749,N_1988);
or U3616 (N_3616,N_51,N_2333);
or U3617 (N_3617,N_769,N_1278);
or U3618 (N_3618,N_1559,N_629);
or U3619 (N_3619,N_734,N_163);
and U3620 (N_3620,N_461,N_2648);
or U3621 (N_3621,N_1386,N_234);
or U3622 (N_3622,N_1327,N_269);
and U3623 (N_3623,N_70,N_1110);
nor U3624 (N_3624,N_2453,N_2852);
or U3625 (N_3625,N_132,N_2214);
or U3626 (N_3626,N_826,N_1271);
or U3627 (N_3627,N_279,N_2952);
or U3628 (N_3628,N_1644,N_795);
and U3629 (N_3629,N_531,N_605);
xor U3630 (N_3630,N_1629,N_176);
and U3631 (N_3631,N_2184,N_1589);
and U3632 (N_3632,N_681,N_8);
nand U3633 (N_3633,N_2038,N_1455);
nand U3634 (N_3634,N_1316,N_2457);
xnor U3635 (N_3635,N_1502,N_2647);
nand U3636 (N_3636,N_2988,N_572);
or U3637 (N_3637,N_198,N_1276);
and U3638 (N_3638,N_1856,N_1779);
xor U3639 (N_3639,N_1746,N_768);
nand U3640 (N_3640,N_1870,N_1425);
or U3641 (N_3641,N_2039,N_2559);
nand U3642 (N_3642,N_139,N_2472);
nand U3643 (N_3643,N_1053,N_1520);
nor U3644 (N_3644,N_219,N_1324);
and U3645 (N_3645,N_1452,N_240);
and U3646 (N_3646,N_1802,N_21);
nor U3647 (N_3647,N_1885,N_2828);
and U3648 (N_3648,N_2358,N_804);
and U3649 (N_3649,N_340,N_2886);
xnor U3650 (N_3650,N_594,N_926);
nand U3651 (N_3651,N_2280,N_2893);
or U3652 (N_3652,N_1593,N_1513);
and U3653 (N_3653,N_1479,N_1827);
xor U3654 (N_3654,N_798,N_167);
and U3655 (N_3655,N_1918,N_1872);
nand U3656 (N_3656,N_503,N_277);
nor U3657 (N_3657,N_2115,N_477);
or U3658 (N_3658,N_2599,N_1528);
nand U3659 (N_3659,N_2473,N_2973);
or U3660 (N_3660,N_927,N_2158);
nor U3661 (N_3661,N_397,N_1305);
xnor U3662 (N_3662,N_1329,N_2810);
or U3663 (N_3663,N_351,N_395);
xor U3664 (N_3664,N_687,N_2363);
nand U3665 (N_3665,N_1921,N_1605);
or U3666 (N_3666,N_1671,N_658);
nand U3667 (N_3667,N_1951,N_2816);
or U3668 (N_3668,N_738,N_301);
nor U3669 (N_3669,N_2827,N_2528);
nor U3670 (N_3670,N_2676,N_2833);
nand U3671 (N_3671,N_539,N_705);
nand U3672 (N_3672,N_1366,N_1943);
xor U3673 (N_3673,N_2096,N_763);
xnor U3674 (N_3674,N_1065,N_942);
nor U3675 (N_3675,N_595,N_907);
nand U3676 (N_3676,N_2678,N_318);
nor U3677 (N_3677,N_430,N_2170);
and U3678 (N_3678,N_1490,N_2289);
and U3679 (N_3679,N_1544,N_2620);
nand U3680 (N_3680,N_2580,N_2117);
nor U3681 (N_3681,N_2341,N_1307);
nor U3682 (N_3682,N_401,N_2031);
or U3683 (N_3683,N_1014,N_1816);
or U3684 (N_3684,N_776,N_1309);
or U3685 (N_3685,N_1623,N_1743);
or U3686 (N_3686,N_1796,N_456);
nand U3687 (N_3687,N_1167,N_2099);
or U3688 (N_3688,N_1443,N_479);
xor U3689 (N_3689,N_1768,N_323);
nand U3690 (N_3690,N_2651,N_730);
xor U3691 (N_3691,N_1748,N_1731);
and U3692 (N_3692,N_2208,N_626);
nand U3693 (N_3693,N_22,N_74);
nand U3694 (N_3694,N_943,N_2371);
or U3695 (N_3695,N_427,N_2683);
and U3696 (N_3696,N_1427,N_601);
xnor U3697 (N_3697,N_2252,N_634);
or U3698 (N_3698,N_2143,N_2311);
nand U3699 (N_3699,N_904,N_2554);
and U3700 (N_3700,N_1558,N_800);
and U3701 (N_3701,N_771,N_2181);
nand U3702 (N_3702,N_882,N_2746);
nor U3703 (N_3703,N_2645,N_1546);
and U3704 (N_3704,N_1140,N_1824);
nand U3705 (N_3705,N_1839,N_2253);
xnor U3706 (N_3706,N_1192,N_2616);
nor U3707 (N_3707,N_600,N_976);
xor U3708 (N_3708,N_501,N_1798);
nor U3709 (N_3709,N_2301,N_1981);
and U3710 (N_3710,N_1337,N_1198);
or U3711 (N_3711,N_86,N_2265);
or U3712 (N_3712,N_348,N_2927);
nand U3713 (N_3713,N_2941,N_2251);
nor U3714 (N_3714,N_748,N_2613);
nand U3715 (N_3715,N_671,N_543);
nand U3716 (N_3716,N_1989,N_1290);
nor U3717 (N_3717,N_28,N_2900);
or U3718 (N_3718,N_2098,N_2558);
nand U3719 (N_3719,N_622,N_265);
nand U3720 (N_3720,N_1575,N_1201);
nor U3721 (N_3721,N_213,N_2741);
xor U3722 (N_3722,N_521,N_124);
xor U3723 (N_3723,N_295,N_258);
nand U3724 (N_3724,N_2675,N_1874);
nor U3725 (N_3725,N_2462,N_2749);
and U3726 (N_3726,N_2800,N_1801);
and U3727 (N_3727,N_2423,N_1670);
nand U3728 (N_3728,N_1143,N_2974);
nand U3729 (N_3729,N_83,N_91);
nor U3730 (N_3730,N_2627,N_996);
nor U3731 (N_3731,N_2327,N_145);
or U3732 (N_3732,N_2254,N_2140);
and U3733 (N_3733,N_2563,N_272);
xnor U3734 (N_3734,N_441,N_1387);
or U3735 (N_3735,N_612,N_2288);
or U3736 (N_3736,N_161,N_732);
or U3737 (N_3737,N_1903,N_1286);
nor U3738 (N_3738,N_2384,N_2536);
nand U3739 (N_3739,N_1262,N_1805);
nor U3740 (N_3740,N_685,N_363);
or U3741 (N_3741,N_1556,N_1535);
or U3742 (N_3742,N_1171,N_532);
xor U3743 (N_3743,N_1987,N_2743);
xor U3744 (N_3744,N_2882,N_2836);
or U3745 (N_3745,N_2431,N_2433);
xnor U3746 (N_3746,N_2516,N_2109);
nor U3747 (N_3747,N_1472,N_2036);
xnor U3748 (N_3748,N_2664,N_2270);
and U3749 (N_3749,N_1599,N_402);
nand U3750 (N_3750,N_2560,N_2557);
nor U3751 (N_3751,N_542,N_1602);
xor U3752 (N_3752,N_955,N_1475);
or U3753 (N_3753,N_964,N_2796);
xnor U3754 (N_3754,N_2229,N_1375);
nor U3755 (N_3755,N_1075,N_621);
and U3756 (N_3756,N_2567,N_1393);
nand U3757 (N_3757,N_585,N_2913);
and U3758 (N_3758,N_396,N_233);
or U3759 (N_3759,N_2510,N_11);
xor U3760 (N_3760,N_1202,N_1970);
or U3761 (N_3761,N_932,N_371);
xnor U3762 (N_3762,N_1667,N_2064);
and U3763 (N_3763,N_1901,N_614);
nor U3764 (N_3764,N_987,N_189);
xnor U3765 (N_3765,N_1929,N_1518);
nand U3766 (N_3766,N_2834,N_1739);
nand U3767 (N_3767,N_2152,N_792);
and U3768 (N_3768,N_2063,N_1029);
or U3769 (N_3769,N_2573,N_842);
and U3770 (N_3770,N_2330,N_434);
xnor U3771 (N_3771,N_1106,N_2881);
xor U3772 (N_3772,N_2622,N_1800);
or U3773 (N_3773,N_1580,N_1540);
or U3774 (N_3774,N_2837,N_848);
or U3775 (N_3775,N_2114,N_2124);
nor U3776 (N_3776,N_2028,N_962);
nor U3777 (N_3777,N_1705,N_1690);
nand U3778 (N_3778,N_232,N_2880);
or U3779 (N_3779,N_2533,N_880);
xor U3780 (N_3780,N_1713,N_2674);
and U3781 (N_3781,N_1021,N_1409);
or U3782 (N_3782,N_1516,N_1913);
xnor U3783 (N_3783,N_1880,N_2848);
nand U3784 (N_3784,N_2865,N_4);
xor U3785 (N_3785,N_1737,N_1174);
nand U3786 (N_3786,N_1113,N_591);
nor U3787 (N_3787,N_760,N_1281);
or U3788 (N_3788,N_496,N_1064);
nand U3789 (N_3789,N_1423,N_2021);
xor U3790 (N_3790,N_354,N_949);
and U3791 (N_3791,N_2577,N_40);
nand U3792 (N_3792,N_2688,N_944);
nand U3793 (N_3793,N_94,N_2299);
and U3794 (N_3794,N_245,N_1222);
xnor U3795 (N_3795,N_895,N_207);
nor U3796 (N_3796,N_981,N_120);
nor U3797 (N_3797,N_960,N_1451);
or U3798 (N_3798,N_1971,N_872);
and U3799 (N_3799,N_775,N_1059);
nand U3800 (N_3800,N_1924,N_1120);
and U3801 (N_3801,N_2752,N_1781);
and U3802 (N_3802,N_1844,N_1453);
nor U3803 (N_3803,N_2454,N_338);
xor U3804 (N_3804,N_2409,N_1857);
nor U3805 (N_3805,N_1673,N_2485);
nand U3806 (N_3806,N_1524,N_2566);
nor U3807 (N_3807,N_786,N_206);
and U3808 (N_3808,N_1905,N_1591);
and U3809 (N_3809,N_547,N_2357);
xor U3810 (N_3810,N_654,N_2295);
xnor U3811 (N_3811,N_778,N_2404);
or U3812 (N_3812,N_1127,N_2284);
or U3813 (N_3813,N_2235,N_1330);
or U3814 (N_3814,N_41,N_1784);
nor U3815 (N_3815,N_1407,N_1223);
and U3816 (N_3816,N_12,N_1317);
or U3817 (N_3817,N_1973,N_439);
and U3818 (N_3818,N_85,N_2555);
and U3819 (N_3819,N_1492,N_1787);
nor U3820 (N_3820,N_1159,N_2347);
nor U3821 (N_3821,N_1097,N_2901);
nand U3822 (N_3822,N_347,N_2626);
or U3823 (N_3823,N_1182,N_934);
xor U3824 (N_3824,N_690,N_2336);
or U3825 (N_3825,N_458,N_2210);
or U3826 (N_3826,N_856,N_1631);
xor U3827 (N_3827,N_908,N_563);
or U3828 (N_3828,N_774,N_791);
xnor U3829 (N_3829,N_2487,N_1349);
and U3830 (N_3830,N_2466,N_995);
nand U3831 (N_3831,N_1105,N_1255);
or U3832 (N_3832,N_194,N_1319);
nor U3833 (N_3833,N_1372,N_1754);
nor U3834 (N_3834,N_2564,N_1446);
and U3835 (N_3835,N_2086,N_860);
or U3836 (N_3836,N_2602,N_1095);
xor U3837 (N_3837,N_1102,N_1462);
or U3838 (N_3838,N_10,N_2572);
nor U3839 (N_3839,N_306,N_854);
nand U3840 (N_3840,N_2945,N_2850);
and U3841 (N_3841,N_2292,N_97);
and U3842 (N_3842,N_2471,N_1331);
xnor U3843 (N_3843,N_1581,N_2383);
or U3844 (N_3844,N_2639,N_1027);
xor U3845 (N_3845,N_782,N_1650);
xor U3846 (N_3846,N_1955,N_320);
xor U3847 (N_3847,N_197,N_2905);
nor U3848 (N_3848,N_1355,N_155);
or U3849 (N_3849,N_2571,N_1964);
xor U3850 (N_3850,N_796,N_615);
and U3851 (N_3851,N_1195,N_1935);
xnor U3852 (N_3852,N_1974,N_2594);
or U3853 (N_3853,N_260,N_1945);
and U3854 (N_3854,N_324,N_2425);
nand U3855 (N_3855,N_1725,N_553);
and U3856 (N_3856,N_2817,N_1465);
or U3857 (N_3857,N_2888,N_688);
or U3858 (N_3858,N_1031,N_289);
nand U3859 (N_3859,N_1413,N_1314);
xnor U3860 (N_3860,N_1009,N_963);
nor U3861 (N_3861,N_855,N_2029);
xnor U3862 (N_3862,N_2237,N_1590);
xor U3863 (N_3863,N_208,N_956);
and U3864 (N_3864,N_2193,N_808);
or U3865 (N_3865,N_2350,N_2853);
and U3866 (N_3866,N_713,N_1172);
xnor U3867 (N_3867,N_383,N_35);
or U3868 (N_3868,N_411,N_1569);
and U3869 (N_3869,N_332,N_2907);
xnor U3870 (N_3870,N_2997,N_815);
xor U3871 (N_3871,N_2644,N_317);
or U3872 (N_3872,N_1025,N_2916);
or U3873 (N_3873,N_469,N_1096);
and U3874 (N_3874,N_292,N_1067);
xor U3875 (N_3875,N_293,N_49);
or U3876 (N_3876,N_2556,N_89);
xnor U3877 (N_3877,N_920,N_84);
and U3878 (N_3878,N_1506,N_556);
and U3879 (N_3879,N_1965,N_623);
xnor U3880 (N_3880,N_725,N_2898);
nand U3881 (N_3881,N_2309,N_67);
nor U3882 (N_3882,N_2150,N_2429);
nand U3883 (N_3883,N_2864,N_1912);
xor U3884 (N_3884,N_2878,N_2090);
nand U3885 (N_3885,N_259,N_1563);
nor U3886 (N_3886,N_2598,N_334);
nor U3887 (N_3887,N_2919,N_959);
nand U3888 (N_3888,N_2172,N_2239);
nand U3889 (N_3889,N_1888,N_2977);
or U3890 (N_3890,N_2699,N_1533);
xnor U3891 (N_3891,N_380,N_1091);
and U3892 (N_3892,N_147,N_218);
or U3893 (N_3893,N_1362,N_2980);
nor U3894 (N_3894,N_349,N_1397);
and U3895 (N_3895,N_1740,N_140);
or U3896 (N_3896,N_2947,N_2470);
xor U3897 (N_3897,N_2324,N_1236);
xor U3898 (N_3898,N_468,N_2416);
or U3899 (N_3899,N_2825,N_1946);
nand U3900 (N_3900,N_845,N_1896);
nor U3901 (N_3901,N_664,N_174);
xnor U3902 (N_3902,N_2617,N_1148);
and U3903 (N_3903,N_2092,N_2276);
or U3904 (N_3904,N_367,N_2111);
nand U3905 (N_3905,N_578,N_418);
and U3906 (N_3906,N_2964,N_1396);
and U3907 (N_3907,N_1785,N_386);
or U3908 (N_3908,N_2744,N_2398);
nor U3909 (N_3909,N_2304,N_597);
nand U3910 (N_3910,N_2607,N_508);
nand U3911 (N_3911,N_1298,N_1019);
or U3912 (N_3912,N_1793,N_889);
nand U3913 (N_3913,N_2067,N_2401);
or U3914 (N_3914,N_1318,N_2187);
nor U3915 (N_3915,N_2052,N_2211);
or U3916 (N_3916,N_1199,N_1820);
or U3917 (N_3917,N_645,N_2377);
and U3918 (N_3918,N_1371,N_1838);
nor U3919 (N_3919,N_599,N_180);
or U3920 (N_3920,N_1292,N_2396);
and U3921 (N_3921,N_823,N_268);
xor U3922 (N_3922,N_1402,N_715);
xnor U3923 (N_3923,N_1606,N_971);
or U3924 (N_3924,N_1571,N_1092);
or U3925 (N_3925,N_2183,N_2189);
nand U3926 (N_3926,N_825,N_1849);
nor U3927 (N_3927,N_697,N_870);
xnor U3928 (N_3928,N_372,N_1709);
nor U3929 (N_3929,N_2010,N_1151);
nor U3930 (N_3930,N_1634,N_2987);
and U3931 (N_3931,N_2011,N_426);
and U3932 (N_3932,N_281,N_755);
or U3933 (N_3933,N_1333,N_2821);
xor U3934 (N_3934,N_1190,N_527);
nor U3935 (N_3935,N_2281,N_34);
or U3936 (N_3936,N_1383,N_1487);
nand U3937 (N_3937,N_1365,N_298);
nand U3938 (N_3938,N_9,N_1978);
xor U3939 (N_3939,N_589,N_1765);
xor U3940 (N_3940,N_551,N_2858);
or U3941 (N_3941,N_1304,N_2677);
xor U3942 (N_3942,N_2465,N_577);
and U3943 (N_3943,N_1421,N_602);
xnor U3944 (N_3944,N_2370,N_1503);
xnor U3945 (N_3945,N_362,N_2238);
and U3946 (N_3946,N_682,N_1197);
nor U3947 (N_3947,N_72,N_1561);
xnor U3948 (N_3948,N_2285,N_1389);
xor U3949 (N_3949,N_2949,N_1230);
xor U3950 (N_3950,N_1235,N_2950);
and U3951 (N_3951,N_736,N_2508);
or U3952 (N_3952,N_329,N_2275);
nand U3953 (N_3953,N_2328,N_969);
and U3954 (N_3954,N_1297,N_799);
nor U3955 (N_3955,N_1049,N_695);
nand U3956 (N_3956,N_2322,N_1662);
nand U3957 (N_3957,N_1449,N_2493);
or U3958 (N_3958,N_117,N_242);
nand U3959 (N_3959,N_555,N_1961);
or U3960 (N_3960,N_2780,N_2784);
nor U3961 (N_3961,N_2996,N_2876);
nor U3962 (N_3962,N_2191,N_2991);
nand U3963 (N_3963,N_1376,N_2009);
nor U3964 (N_3964,N_2345,N_1156);
or U3965 (N_3965,N_1897,N_2003);
or U3966 (N_3966,N_1977,N_2051);
or U3967 (N_3967,N_2201,N_2660);
nor U3968 (N_3968,N_1438,N_1392);
nor U3969 (N_3969,N_2126,N_2422);
and U3970 (N_3970,N_17,N_2608);
or U3971 (N_3971,N_698,N_598);
or U3972 (N_3972,N_1525,N_482);
xnor U3973 (N_3973,N_1821,N_1863);
xor U3974 (N_3974,N_1185,N_632);
and U3975 (N_3975,N_1636,N_2321);
or U3976 (N_3976,N_700,N_2799);
xor U3977 (N_3977,N_43,N_947);
nor U3978 (N_3978,N_1129,N_435);
and U3979 (N_3979,N_63,N_2492);
and U3980 (N_3980,N_2948,N_1360);
nor U3981 (N_3981,N_1891,N_966);
nor U3982 (N_3982,N_2589,N_2340);
and U3983 (N_3983,N_2332,N_2241);
and U3984 (N_3984,N_90,N_246);
or U3985 (N_3985,N_1168,N_1179);
and U3986 (N_3986,N_817,N_201);
or U3987 (N_3987,N_2089,N_756);
and U3988 (N_3988,N_1414,N_2468);
nor U3989 (N_3989,N_377,N_656);
nand U3990 (N_3990,N_1699,N_517);
nand U3991 (N_3991,N_1790,N_2712);
xnor U3992 (N_3992,N_2811,N_2961);
xor U3993 (N_3993,N_1437,N_1865);
xor U3994 (N_3994,N_1303,N_2513);
and U3995 (N_3995,N_20,N_858);
xor U3996 (N_3996,N_1164,N_2552);
and U3997 (N_3997,N_1714,N_29);
nand U3998 (N_3998,N_1659,N_2534);
xor U3999 (N_3999,N_2053,N_1005);
or U4000 (N_4000,N_2981,N_2903);
nor U4001 (N_4001,N_1710,N_1220);
or U4002 (N_4002,N_2937,N_1141);
and U4003 (N_4003,N_1814,N_2459);
and U4004 (N_4004,N_1107,N_283);
nor U4005 (N_4005,N_2642,N_179);
nand U4006 (N_4006,N_278,N_1050);
nor U4007 (N_4007,N_2112,N_1111);
nor U4008 (N_4008,N_2917,N_1448);
and U4009 (N_4009,N_2514,N_2054);
and U4010 (N_4010,N_1039,N_1018);
and U4011 (N_4011,N_1158,N_1445);
xor U4012 (N_4012,N_2173,N_2417);
and U4013 (N_4013,N_366,N_1549);
or U4014 (N_4014,N_1876,N_1664);
nor U4015 (N_4015,N_1275,N_2851);
xnor U4016 (N_4016,N_250,N_1995);
nand U4017 (N_4017,N_2568,N_1033);
nand U4018 (N_4018,N_1045,N_141);
xnor U4019 (N_4019,N_2494,N_677);
xor U4020 (N_4020,N_247,N_252);
nand U4021 (N_4021,N_1919,N_2245);
and U4022 (N_4022,N_1103,N_1543);
nand U4023 (N_4023,N_2364,N_1825);
xor U4024 (N_4024,N_1630,N_2529);
and U4025 (N_4025,N_264,N_2283);
xor U4026 (N_4026,N_2524,N_409);
and U4027 (N_4027,N_847,N_1153);
xnor U4028 (N_4028,N_514,N_1010);
and U4029 (N_4029,N_1618,N_2174);
and U4030 (N_4030,N_2581,N_2355);
nand U4031 (N_4031,N_2000,N_2592);
xnor U4032 (N_4032,N_231,N_1755);
and U4033 (N_4033,N_1344,N_862);
or U4034 (N_4034,N_2670,N_2768);
and U4035 (N_4035,N_2294,N_1422);
and U4036 (N_4036,N_704,N_1406);
and U4037 (N_4037,N_1845,N_1351);
or U4038 (N_4038,N_752,N_422);
or U4039 (N_4039,N_1625,N_957);
or U4040 (N_4040,N_1994,N_853);
nor U4041 (N_4041,N_1439,N_1020);
or U4042 (N_4042,N_1403,N_2939);
nor U4043 (N_4043,N_2778,N_1277);
or U4044 (N_4044,N_1482,N_1391);
xnor U4045 (N_4045,N_2659,N_2486);
nand U4046 (N_4046,N_2820,N_2455);
nor U4047 (N_4047,N_1132,N_720);
xor U4048 (N_4048,N_1442,N_2506);
nor U4049 (N_4049,N_419,N_453);
nand U4050 (N_4050,N_2206,N_1165);
or U4051 (N_4051,N_1939,N_1689);
nand U4052 (N_4052,N_1982,N_1993);
nand U4053 (N_4053,N_358,N_2277);
nand U4054 (N_4054,N_463,N_1125);
xor U4055 (N_4055,N_2804,N_702);
nor U4056 (N_4056,N_1037,N_1283);
or U4057 (N_4057,N_1511,N_1108);
nor U4058 (N_4058,N_1752,N_1555);
and U4059 (N_4059,N_2802,N_1302);
and U4060 (N_4060,N_911,N_1341);
or U4061 (N_4061,N_2955,N_1139);
nand U4062 (N_4062,N_2634,N_1997);
xor U4063 (N_4063,N_2854,N_1944);
or U4064 (N_4064,N_2899,N_1660);
nor U4065 (N_4065,N_87,N_118);
or U4066 (N_4066,N_379,N_570);
and U4067 (N_4067,N_550,N_2303);
and U4068 (N_4068,N_1677,N_1861);
nand U4069 (N_4069,N_1692,N_840);
nand U4070 (N_4070,N_2078,N_1537);
or U4071 (N_4071,N_2526,N_346);
and U4072 (N_4072,N_261,N_1695);
and U4073 (N_4073,N_2188,N_2389);
nand U4074 (N_4074,N_2641,N_573);
or U4075 (N_4075,N_119,N_2923);
or U4076 (N_4076,N_1940,N_813);
xor U4077 (N_4077,N_398,N_484);
and U4078 (N_4078,N_256,N_584);
nor U4079 (N_4079,N_1461,N_327);
or U4080 (N_4080,N_1738,N_151);
xor U4081 (N_4081,N_2710,N_2343);
or U4082 (N_4082,N_498,N_1232);
and U4083 (N_4083,N_1780,N_2490);
nor U4084 (N_4084,N_812,N_1121);
nor U4085 (N_4085,N_835,N_1585);
and U4086 (N_4086,N_945,N_1358);
xnor U4087 (N_4087,N_126,N_2070);
nand U4088 (N_4088,N_1925,N_2758);
xor U4089 (N_4089,N_188,N_129);
nor U4090 (N_4090,N_784,N_2100);
nand U4091 (N_4091,N_545,N_1893);
xnor U4092 (N_4092,N_2807,N_1426);
nor U4093 (N_4093,N_474,N_2924);
nor U4094 (N_4094,N_1867,N_1984);
nor U4095 (N_4095,N_2149,N_2553);
nor U4096 (N_4096,N_2867,N_2546);
xor U4097 (N_4097,N_59,N_948);
or U4098 (N_4098,N_1976,N_2839);
nor U4099 (N_4099,N_1875,N_381);
or U4100 (N_4100,N_1786,N_1313);
and U4101 (N_4101,N_3,N_661);
xnor U4102 (N_4102,N_2716,N_400);
xnor U4103 (N_4103,N_2547,N_2765);
and U4104 (N_4104,N_1497,N_2375);
nor U4105 (N_4105,N_2451,N_1744);
xnor U4106 (N_4106,N_2866,N_901);
and U4107 (N_4107,N_2612,N_940);
xor U4108 (N_4108,N_23,N_2729);
xnor U4109 (N_4109,N_420,N_494);
or U4110 (N_4110,N_2649,N_2717);
nor U4111 (N_4111,N_2419,N_2889);
nor U4112 (N_4112,N_2209,N_1200);
nor U4113 (N_4113,N_2228,N_1212);
nand U4114 (N_4114,N_1268,N_1084);
xor U4115 (N_4115,N_2956,N_2042);
or U4116 (N_4116,N_2131,N_818);
and U4117 (N_4117,N_2394,N_1180);
or U4118 (N_4118,N_321,N_196);
nand U4119 (N_4119,N_2030,N_1325);
or U4120 (N_4120,N_885,N_1788);
xnor U4121 (N_4121,N_2316,N_912);
or U4122 (N_4122,N_1147,N_2055);
and U4123 (N_4123,N_1756,N_2057);
nand U4124 (N_4124,N_1567,N_2588);
nor U4125 (N_4125,N_2918,N_2374);
or U4126 (N_4126,N_254,N_2748);
xnor U4127 (N_4127,N_1124,N_193);
nor U4128 (N_4128,N_952,N_368);
nor U4129 (N_4129,N_2259,N_1450);
xnor U4130 (N_4130,N_226,N_1367);
nor U4131 (N_4131,N_1118,N_125);
nor U4132 (N_4132,N_1013,N_1923);
xnor U4133 (N_4133,N_2975,N_587);
nand U4134 (N_4134,N_2925,N_2562);
nor U4135 (N_4135,N_819,N_48);
nor U4136 (N_4136,N_2739,N_1745);
and U4137 (N_4137,N_809,N_2862);
xor U4138 (N_4138,N_214,N_789);
nor U4139 (N_4139,N_537,N_1637);
xor U4140 (N_4140,N_1061,N_2761);
nor U4141 (N_4141,N_2982,N_1902);
xnor U4142 (N_4142,N_406,N_2805);
nand U4143 (N_4143,N_2269,N_2435);
and U4144 (N_4144,N_350,N_2353);
nor U4145 (N_4145,N_1583,N_1949);
xor U4146 (N_4146,N_2887,N_267);
and U4147 (N_4147,N_2186,N_2247);
nor U4148 (N_4148,N_2291,N_182);
and U4149 (N_4149,N_762,N_1169);
nand U4150 (N_4150,N_2835,N_2737);
xor U4151 (N_4151,N_693,N_990);
xor U4152 (N_4152,N_757,N_2787);
nor U4153 (N_4153,N_863,N_2979);
or U4154 (N_4154,N_1504,N_109);
and U4155 (N_4155,N_871,N_2872);
or U4156 (N_4156,N_701,N_1772);
nand U4157 (N_4157,N_1256,N_2873);
or U4158 (N_4158,N_1473,N_2933);
and U4159 (N_4159,N_2942,N_113);
xnor U4160 (N_4160,N_1052,N_1711);
or U4161 (N_4161,N_436,N_2300);
and U4162 (N_4162,N_410,N_200);
nand U4163 (N_4163,N_1529,N_982);
nor U4164 (N_4164,N_2582,N_2262);
and U4165 (N_4165,N_972,N_1823);
nor U4166 (N_4166,N_2874,N_2236);
and U4167 (N_4167,N_1582,N_2226);
or U4168 (N_4168,N_2013,N_1522);
xnor U4169 (N_4169,N_56,N_2922);
and U4170 (N_4170,N_389,N_2747);
or U4171 (N_4171,N_203,N_1299);
and U4172 (N_4172,N_2119,N_1986);
or U4173 (N_4173,N_2037,N_1864);
and U4174 (N_4174,N_2088,N_1975);
xor U4175 (N_4175,N_1142,N_1672);
and U4176 (N_4176,N_2145,N_2541);
nor U4177 (N_4177,N_2798,N_2379);
nor U4178 (N_4178,N_2633,N_1707);
nor U4179 (N_4179,N_2056,N_2069);
nand U4180 (N_4180,N_1942,N_967);
xor U4181 (N_4181,N_2985,N_2754);
and U4182 (N_4182,N_210,N_997);
or U4183 (N_4183,N_2071,N_2938);
or U4184 (N_4184,N_1899,N_492);
and U4185 (N_4185,N_1530,N_1173);
nor U4186 (N_4186,N_2951,N_428);
or U4187 (N_4187,N_620,N_2521);
or U4188 (N_4188,N_1854,N_291);
xnor U4189 (N_4189,N_2707,N_2842);
nor U4190 (N_4190,N_2614,N_830);
nand U4191 (N_4191,N_1922,N_286);
or U4192 (N_4192,N_801,N_875);
xnor U4193 (N_4193,N_2430,N_839);
xor U4194 (N_4194,N_134,N_384);
or U4195 (N_4195,N_2543,N_1263);
and U4196 (N_4196,N_2696,N_2059);
or U4197 (N_4197,N_2313,N_788);
or U4198 (N_4198,N_2771,N_290);
nand U4199 (N_4199,N_2221,N_922);
nand U4200 (N_4200,N_1799,N_450);
and U4201 (N_4201,N_1154,N_859);
and U4202 (N_4202,N_2019,N_1411);
xnor U4203 (N_4203,N_816,N_868);
and U4204 (N_4204,N_2689,N_310);
nand U4205 (N_4205,N_1762,N_639);
or U4206 (N_4206,N_721,N_2442);
xor U4207 (N_4207,N_883,N_2702);
or U4208 (N_4208,N_241,N_1767);
xnor U4209 (N_4209,N_62,N_1008);
or U4210 (N_4210,N_1653,N_106);
or U4211 (N_4211,N_562,N_2603);
or U4212 (N_4212,N_1595,N_1999);
or U4213 (N_4213,N_2789,N_2349);
nor U4214 (N_4214,N_582,N_2538);
nor U4215 (N_4215,N_460,N_824);
or U4216 (N_4216,N_2335,N_2424);
nand U4217 (N_4217,N_2679,N_1614);
and U4218 (N_4218,N_914,N_1640);
xnor U4219 (N_4219,N_951,N_1859);
or U4220 (N_4220,N_217,N_2520);
nand U4221 (N_4221,N_1279,N_153);
nand U4222 (N_4222,N_672,N_297);
nor U4223 (N_4223,N_37,N_1968);
nand U4224 (N_4224,N_974,N_1104);
nor U4225 (N_4225,N_2484,N_1417);
xor U4226 (N_4226,N_1015,N_674);
and U4227 (N_4227,N_1948,N_2640);
nand U4228 (N_4228,N_724,N_646);
and U4229 (N_4229,N_2121,N_679);
or U4230 (N_4230,N_169,N_998);
and U4231 (N_4231,N_2093,N_2703);
nand U4232 (N_4232,N_192,N_339);
and U4233 (N_4233,N_2694,N_2320);
xnor U4234 (N_4234,N_2503,N_2477);
and U4235 (N_4235,N_2050,N_1489);
and U4236 (N_4236,N_1914,N_2);
xnor U4237 (N_4237,N_714,N_235);
or U4238 (N_4238,N_270,N_27);
nor U4239 (N_4239,N_2034,N_2797);
or U4240 (N_4240,N_2826,N_1715);
nor U4241 (N_4241,N_2636,N_512);
xor U4242 (N_4242,N_1678,N_429);
nor U4243 (N_4243,N_737,N_2076);
nor U4244 (N_4244,N_921,N_2456);
and U4245 (N_4245,N_2890,N_1038);
nor U4246 (N_4246,N_1181,N_1209);
or U4247 (N_4247,N_1339,N_1265);
and U4248 (N_4248,N_764,N_57);
or U4249 (N_4249,N_444,N_1369);
xor U4250 (N_4250,N_1601,N_1471);
and U4251 (N_4251,N_1016,N_110);
and U4252 (N_4252,N_2127,N_2958);
nand U4253 (N_4253,N_2027,N_1410);
nand U4254 (N_4254,N_337,N_506);
nand U4255 (N_4255,N_451,N_2518);
nor U4256 (N_4256,N_1353,N_1483);
and U4257 (N_4257,N_2222,N_2079);
or U4258 (N_4258,N_837,N_906);
or U4259 (N_4259,N_1312,N_2256);
xnor U4260 (N_4260,N_2732,N_2043);
nor U4261 (N_4261,N_481,N_2750);
xnor U4262 (N_4262,N_1186,N_2740);
xor U4263 (N_4263,N_1776,N_718);
nor U4264 (N_4264,N_2519,N_1395);
xor U4265 (N_4265,N_80,N_2593);
and U4266 (N_4266,N_7,N_2713);
or U4267 (N_4267,N_535,N_2248);
nand U4268 (N_4268,N_262,N_2983);
xor U4269 (N_4269,N_1704,N_2178);
xor U4270 (N_4270,N_92,N_127);
xor U4271 (N_4271,N_2637,N_355);
xor U4272 (N_4272,N_475,N_55);
nor U4273 (N_4273,N_1900,N_699);
xor U4274 (N_4274,N_1166,N_2532);
and U4275 (N_4275,N_2142,N_236);
or U4276 (N_4276,N_2022,N_271);
or U4277 (N_4277,N_2575,N_1679);
and U4278 (N_4278,N_2198,N_910);
and U4279 (N_4279,N_1655,N_2306);
xnor U4280 (N_4280,N_897,N_2147);
nor U4281 (N_4281,N_115,N_1219);
xnor U4282 (N_4282,N_2595,N_2576);
nand U4283 (N_4283,N_1218,N_393);
xor U4284 (N_4284,N_1240,N_2871);
nor U4285 (N_4285,N_2497,N_209);
and U4286 (N_4286,N_1909,N_413);
or U4287 (N_4287,N_638,N_2968);
nor U4288 (N_4288,N_2971,N_2219);
nor U4289 (N_4289,N_1573,N_2273);
nand U4290 (N_4290,N_2877,N_1966);
or U4291 (N_4291,N_2308,N_248);
or U4292 (N_4292,N_750,N_2806);
or U4293 (N_4293,N_2203,N_2458);
nor U4294 (N_4294,N_1830,N_930);
and U4295 (N_4295,N_1023,N_2319);
nand U4296 (N_4296,N_1157,N_2843);
or U4297 (N_4297,N_979,N_2474);
or U4298 (N_4298,N_2539,N_2106);
nor U4299 (N_4299,N_2110,N_865);
or U4300 (N_4300,N_1454,N_2759);
nand U4301 (N_4301,N_315,N_1990);
xor U4302 (N_4302,N_1388,N_2770);
nand U4303 (N_4303,N_1347,N_2095);
or U4304 (N_4304,N_1972,N_2015);
or U4305 (N_4305,N_1161,N_1488);
nand U4306 (N_4306,N_1932,N_99);
xnor U4307 (N_4307,N_1364,N_1809);
nand U4308 (N_4308,N_936,N_2725);
nand U4309 (N_4309,N_433,N_162);
xnor U4310 (N_4310,N_1757,N_2136);
and U4311 (N_4311,N_1760,N_744);
or U4312 (N_4312,N_2479,N_1587);
and U4313 (N_4313,N_1022,N_2083);
nand U4314 (N_4314,N_1848,N_1665);
or U4315 (N_4315,N_1647,N_1792);
xor U4316 (N_4316,N_1320,N_1348);
nor U4317 (N_4317,N_228,N_694);
nand U4318 (N_4318,N_751,N_2723);
nor U4319 (N_4319,N_359,N_1457);
or U4320 (N_4320,N_112,N_678);
xnor U4321 (N_4321,N_2196,N_1343);
and U4322 (N_4322,N_2223,N_146);
nand U4323 (N_4323,N_2434,N_2998);
xnor U4324 (N_4324,N_2097,N_2569);
nand U4325 (N_4325,N_46,N_2378);
or U4326 (N_4326,N_559,N_1354);
nor U4327 (N_4327,N_466,N_2138);
or U4328 (N_4328,N_1078,N_104);
nand U4329 (N_4329,N_1338,N_1311);
nand U4330 (N_4330,N_360,N_2824);
and U4331 (N_4331,N_2691,N_1399);
or U4332 (N_4332,N_13,N_1048);
and U4333 (N_4333,N_1610,N_1137);
nand U4334 (N_4334,N_175,N_483);
xor U4335 (N_4335,N_2978,N_1572);
nor U4336 (N_4336,N_1088,N_2243);
nand U4337 (N_4337,N_2630,N_994);
or U4338 (N_4338,N_2605,N_978);
or U4339 (N_4339,N_849,N_544);
and U4340 (N_4340,N_2387,N_2551);
xor U4341 (N_4341,N_1953,N_1771);
xor U4342 (N_4342,N_1087,N_1196);
xnor U4343 (N_4343,N_312,N_1683);
and U4344 (N_4344,N_1060,N_2840);
xnor U4345 (N_4345,N_891,N_2331);
or U4346 (N_4346,N_467,N_2074);
nand U4347 (N_4347,N_983,N_2666);
and U4348 (N_4348,N_415,N_1879);
and U4349 (N_4349,N_485,N_2132);
and U4350 (N_4350,N_2500,N_2934);
nor U4351 (N_4351,N_1578,N_2444);
nor U4352 (N_4352,N_1216,N_2972);
nor U4353 (N_4353,N_2596,N_1042);
and U4354 (N_4354,N_373,N_378);
or U4355 (N_4355,N_1542,N_2507);
nand U4356 (N_4356,N_716,N_1024);
nand U4357 (N_4357,N_742,N_445);
xnor U4358 (N_4358,N_1607,N_630);
xor U4359 (N_4359,N_905,N_2368);
or U4360 (N_4360,N_2861,N_916);
or U4361 (N_4361,N_1404,N_2205);
or U4362 (N_4362,N_516,N_518);
or U4363 (N_4363,N_2403,N_1270);
or U4364 (N_4364,N_2863,N_642);
and U4365 (N_4365,N_2579,N_61);
xnor U4366 (N_4366,N_1927,N_1701);
xor U4367 (N_4367,N_1822,N_1534);
and U4368 (N_4368,N_1586,N_1177);
nor U4369 (N_4369,N_680,N_1852);
xnor U4370 (N_4370,N_1117,N_1519);
xor U4371 (N_4371,N_2990,N_2344);
nand U4372 (N_4372,N_2163,N_2738);
nand U4373 (N_4373,N_2261,N_2382);
nor U4374 (N_4374,N_2672,N_2475);
or U4375 (N_4375,N_1476,N_876);
and U4376 (N_4376,N_1521,N_1657);
and U4377 (N_4377,N_965,N_1884);
or U4378 (N_4378,N_2523,N_759);
nand U4379 (N_4379,N_536,N_1076);
xnor U4380 (N_4380,N_2312,N_590);
xnor U4381 (N_4381,N_2418,N_2199);
or U4382 (N_4382,N_529,N_316);
nand U4383 (N_4383,N_480,N_2001);
nand U4384 (N_4384,N_2085,N_2460);
xnor U4385 (N_4385,N_1272,N_1574);
or U4386 (N_4386,N_2278,N_838);
and U4387 (N_4387,N_1225,N_2904);
nand U4388 (N_4388,N_1747,N_150);
nor U4389 (N_4389,N_1498,N_2432);
xor U4390 (N_4390,N_2023,N_2912);
and U4391 (N_4391,N_754,N_857);
or U4392 (N_4392,N_2325,N_19);
nor U4393 (N_4393,N_212,N_2910);
or U4394 (N_4394,N_138,N_1908);
nor U4395 (N_4395,N_294,N_1373);
xor U4396 (N_4396,N_1523,N_2584);
nand U4397 (N_4397,N_711,N_47);
nand U4398 (N_4398,N_417,N_1458);
nand U4399 (N_4399,N_1811,N_1126);
or U4400 (N_4400,N_709,N_1284);
xor U4401 (N_4401,N_1539,N_633);
xor U4402 (N_4402,N_593,N_1564);
nand U4403 (N_4403,N_251,N_2156);
nor U4404 (N_4404,N_1855,N_185);
nand U4405 (N_4405,N_941,N_1736);
nand U4406 (N_4406,N_604,N_2692);
nor U4407 (N_4407,N_2812,N_1652);
nand U4408 (N_4408,N_2847,N_821);
nand U4409 (N_4409,N_526,N_779);
xnor U4410 (N_4410,N_303,N_1370);
and U4411 (N_4411,N_2690,N_806);
and U4412 (N_4412,N_1210,N_2141);
or U4413 (N_4413,N_2777,N_2646);
nor U4414 (N_4414,N_797,N_165);
xnor U4415 (N_4415,N_1911,N_2838);
or U4416 (N_4416,N_2668,N_2162);
xor U4417 (N_4417,N_2769,N_32);
or U4418 (N_4418,N_1627,N_1598);
or U4419 (N_4419,N_2337,N_1847);
nand U4420 (N_4420,N_1123,N_1957);
and U4421 (N_4421,N_2808,N_1846);
xnor U4422 (N_4422,N_2290,N_1464);
and U4423 (N_4423,N_440,N_1466);
nor U4424 (N_4424,N_1435,N_2439);
xor U4425 (N_4425,N_2629,N_1635);
nand U4426 (N_4426,N_2650,N_1215);
or U4427 (N_4427,N_2504,N_2004);
and U4428 (N_4428,N_2962,N_183);
nand U4429 (N_4429,N_1188,N_2705);
xor U4430 (N_4430,N_2774,N_2885);
nor U4431 (N_4431,N_31,N_2671);
nand U4432 (N_4432,N_1866,N_1527);
or U4433 (N_4433,N_1654,N_2586);
nand U4434 (N_4434,N_2367,N_2498);
nand U4435 (N_4435,N_692,N_2267);
or U4436 (N_4436,N_2476,N_743);
and U4437 (N_4437,N_783,N_2246);
xnor U4438 (N_4438,N_1842,N_1077);
nor U4439 (N_4439,N_1794,N_2356);
or U4440 (N_4440,N_447,N_1703);
nor U4441 (N_4441,N_2480,N_1394);
or U4442 (N_4442,N_2638,N_2654);
or U4443 (N_4443,N_1253,N_1007);
nor U4444 (N_4444,N_668,N_2361);
nor U4445 (N_4445,N_2860,N_1806);
nand U4446 (N_4446,N_2940,N_449);
and U4447 (N_4447,N_877,N_1906);
or U4448 (N_4448,N_149,N_2365);
xor U4449 (N_4449,N_1596,N_2216);
nor U4450 (N_4450,N_1228,N_1083);
nand U4451 (N_4451,N_1682,N_2179);
or U4452 (N_4452,N_2448,N_765);
xnor U4453 (N_4453,N_1963,N_1959);
or U4454 (N_4454,N_2570,N_1770);
or U4455 (N_4455,N_644,N_69);
and U4456 (N_4456,N_893,N_2902);
and U4457 (N_4457,N_525,N_958);
nand U4458 (N_4458,N_2225,N_416);
and U4459 (N_4459,N_712,N_810);
nor U4460 (N_4460,N_1819,N_707);
or U4461 (N_4461,N_1322,N_1342);
and U4462 (N_4462,N_1377,N_2108);
nor U4463 (N_4463,N_65,N_999);
nor U4464 (N_4464,N_18,N_2869);
and U4465 (N_4465,N_2360,N_2755);
or U4466 (N_4466,N_221,N_341);
nor U4467 (N_4467,N_2137,N_2440);
or U4468 (N_4468,N_60,N_793);
nand U4469 (N_4469,N_1368,N_2609);
nor U4470 (N_4470,N_1432,N_343);
xnor U4471 (N_4471,N_148,N_2342);
nand U4472 (N_4472,N_1877,N_1658);
and U4473 (N_4473,N_2652,N_2989);
nand U4474 (N_4474,N_2390,N_2491);
nor U4475 (N_4475,N_2687,N_510);
or U4476 (N_4476,N_2318,N_2482);
xnor U4477 (N_4477,N_1456,N_2619);
nor U4478 (N_4478,N_365,N_2776);
xnor U4479 (N_4479,N_1724,N_2315);
nand U4480 (N_4480,N_1803,N_2601);
xnor U4481 (N_4481,N_777,N_2157);
nor U4482 (N_4482,N_2168,N_1101);
nor U4483 (N_4483,N_950,N_785);
and U4484 (N_4484,N_811,N_2819);
or U4485 (N_4485,N_280,N_2257);
xor U4486 (N_4486,N_160,N_1418);
xnor U4487 (N_4487,N_2421,N_991);
xnor U4488 (N_4488,N_128,N_1721);
xnor U4489 (N_4489,N_706,N_1576);
xnor U4490 (N_4490,N_255,N_1381);
nor U4491 (N_4491,N_2118,N_1828);
nand U4492 (N_4492,N_2139,N_2151);
nand U4493 (N_4493,N_391,N_568);
nor U4494 (N_4494,N_1611,N_382);
nand U4495 (N_4495,N_1686,N_2348);
nor U4496 (N_4496,N_1941,N_1379);
xor U4497 (N_4497,N_1495,N_156);
nand U4498 (N_4498,N_618,N_2709);
nor U4499 (N_4499,N_187,N_2736);
nand U4500 (N_4500,N_1512,N_510);
nand U4501 (N_4501,N_1838,N_388);
nor U4502 (N_4502,N_483,N_2295);
or U4503 (N_4503,N_559,N_2168);
nor U4504 (N_4504,N_2756,N_671);
xor U4505 (N_4505,N_2495,N_1461);
and U4506 (N_4506,N_2597,N_2412);
nor U4507 (N_4507,N_347,N_1078);
nand U4508 (N_4508,N_1881,N_588);
and U4509 (N_4509,N_264,N_827);
xor U4510 (N_4510,N_2732,N_1960);
nand U4511 (N_4511,N_1569,N_2706);
and U4512 (N_4512,N_1344,N_2579);
and U4513 (N_4513,N_471,N_1121);
xor U4514 (N_4514,N_1207,N_2882);
nand U4515 (N_4515,N_637,N_1085);
nand U4516 (N_4516,N_1766,N_1467);
nor U4517 (N_4517,N_1425,N_849);
xor U4518 (N_4518,N_404,N_94);
nor U4519 (N_4519,N_1941,N_167);
and U4520 (N_4520,N_2900,N_2992);
nand U4521 (N_4521,N_744,N_2790);
or U4522 (N_4522,N_1371,N_488);
xnor U4523 (N_4523,N_1698,N_424);
xnor U4524 (N_4524,N_878,N_1891);
xnor U4525 (N_4525,N_1313,N_649);
or U4526 (N_4526,N_273,N_103);
and U4527 (N_4527,N_1086,N_1368);
nor U4528 (N_4528,N_173,N_1233);
xnor U4529 (N_4529,N_2771,N_2127);
or U4530 (N_4530,N_2795,N_205);
nor U4531 (N_4531,N_2103,N_446);
nor U4532 (N_4532,N_2590,N_2438);
nor U4533 (N_4533,N_676,N_1937);
xnor U4534 (N_4534,N_2392,N_2767);
or U4535 (N_4535,N_680,N_2069);
or U4536 (N_4536,N_0,N_2973);
or U4537 (N_4537,N_1748,N_1970);
nand U4538 (N_4538,N_1032,N_947);
and U4539 (N_4539,N_1920,N_407);
and U4540 (N_4540,N_1523,N_2250);
xnor U4541 (N_4541,N_1190,N_187);
and U4542 (N_4542,N_2752,N_1971);
nor U4543 (N_4543,N_2177,N_1574);
nor U4544 (N_4544,N_207,N_2912);
and U4545 (N_4545,N_1792,N_1600);
nand U4546 (N_4546,N_1161,N_1817);
xnor U4547 (N_4547,N_2257,N_643);
nor U4548 (N_4548,N_401,N_2363);
nand U4549 (N_4549,N_632,N_2822);
xor U4550 (N_4550,N_2064,N_1558);
nor U4551 (N_4551,N_2435,N_604);
and U4552 (N_4552,N_2893,N_201);
nor U4553 (N_4553,N_1729,N_1784);
nor U4554 (N_4554,N_2136,N_682);
or U4555 (N_4555,N_887,N_1030);
and U4556 (N_4556,N_1881,N_1561);
and U4557 (N_4557,N_341,N_2488);
nor U4558 (N_4558,N_1426,N_587);
or U4559 (N_4559,N_2530,N_2314);
and U4560 (N_4560,N_1704,N_2153);
and U4561 (N_4561,N_929,N_2534);
and U4562 (N_4562,N_656,N_708);
xor U4563 (N_4563,N_2201,N_1845);
xnor U4564 (N_4564,N_1462,N_1625);
and U4565 (N_4565,N_103,N_2298);
and U4566 (N_4566,N_2289,N_1400);
xnor U4567 (N_4567,N_44,N_2473);
nand U4568 (N_4568,N_2250,N_421);
nor U4569 (N_4569,N_434,N_1831);
and U4570 (N_4570,N_417,N_1774);
or U4571 (N_4571,N_2448,N_2644);
or U4572 (N_4572,N_76,N_1963);
or U4573 (N_4573,N_2477,N_299);
and U4574 (N_4574,N_328,N_2409);
xnor U4575 (N_4575,N_1655,N_1338);
nand U4576 (N_4576,N_2043,N_2472);
nor U4577 (N_4577,N_399,N_230);
nand U4578 (N_4578,N_2438,N_2758);
xnor U4579 (N_4579,N_2305,N_1916);
nor U4580 (N_4580,N_2978,N_2532);
or U4581 (N_4581,N_2612,N_1445);
and U4582 (N_4582,N_2111,N_432);
or U4583 (N_4583,N_1195,N_1088);
or U4584 (N_4584,N_277,N_1951);
xor U4585 (N_4585,N_2140,N_803);
nor U4586 (N_4586,N_2479,N_1454);
nor U4587 (N_4587,N_363,N_1679);
or U4588 (N_4588,N_2119,N_71);
or U4589 (N_4589,N_941,N_1169);
nand U4590 (N_4590,N_147,N_1400);
nor U4591 (N_4591,N_2901,N_596);
xor U4592 (N_4592,N_791,N_225);
nand U4593 (N_4593,N_179,N_2325);
and U4594 (N_4594,N_1548,N_2157);
and U4595 (N_4595,N_300,N_1941);
xnor U4596 (N_4596,N_1166,N_234);
nand U4597 (N_4597,N_2296,N_1369);
nand U4598 (N_4598,N_2119,N_2186);
xnor U4599 (N_4599,N_488,N_2916);
or U4600 (N_4600,N_701,N_2600);
and U4601 (N_4601,N_1492,N_2006);
nor U4602 (N_4602,N_882,N_391);
xnor U4603 (N_4603,N_807,N_559);
xnor U4604 (N_4604,N_1980,N_440);
nand U4605 (N_4605,N_713,N_2388);
and U4606 (N_4606,N_885,N_2264);
and U4607 (N_4607,N_1583,N_1908);
nand U4608 (N_4608,N_336,N_2371);
nand U4609 (N_4609,N_2564,N_1074);
and U4610 (N_4610,N_1960,N_1285);
or U4611 (N_4611,N_317,N_952);
or U4612 (N_4612,N_430,N_1983);
nand U4613 (N_4613,N_1130,N_738);
xnor U4614 (N_4614,N_2343,N_2531);
nand U4615 (N_4615,N_696,N_552);
xor U4616 (N_4616,N_877,N_153);
and U4617 (N_4617,N_2988,N_982);
xor U4618 (N_4618,N_1546,N_1691);
xnor U4619 (N_4619,N_1278,N_2518);
xor U4620 (N_4620,N_2912,N_2134);
xnor U4621 (N_4621,N_1436,N_305);
xnor U4622 (N_4622,N_1881,N_591);
nand U4623 (N_4623,N_1943,N_1854);
nor U4624 (N_4624,N_853,N_719);
and U4625 (N_4625,N_103,N_169);
or U4626 (N_4626,N_624,N_2460);
nor U4627 (N_4627,N_258,N_1720);
or U4628 (N_4628,N_766,N_338);
nand U4629 (N_4629,N_2027,N_1927);
nor U4630 (N_4630,N_369,N_2303);
and U4631 (N_4631,N_2515,N_2389);
nand U4632 (N_4632,N_2197,N_1113);
nand U4633 (N_4633,N_1405,N_651);
nor U4634 (N_4634,N_2221,N_1923);
nor U4635 (N_4635,N_84,N_2748);
xnor U4636 (N_4636,N_252,N_1126);
and U4637 (N_4637,N_258,N_2103);
or U4638 (N_4638,N_31,N_1002);
nand U4639 (N_4639,N_2732,N_156);
nand U4640 (N_4640,N_1545,N_677);
xor U4641 (N_4641,N_2497,N_1481);
nand U4642 (N_4642,N_2355,N_796);
nand U4643 (N_4643,N_1201,N_646);
nand U4644 (N_4644,N_336,N_2889);
nor U4645 (N_4645,N_2813,N_966);
nand U4646 (N_4646,N_2371,N_2127);
nor U4647 (N_4647,N_1052,N_1892);
or U4648 (N_4648,N_2985,N_308);
and U4649 (N_4649,N_2280,N_1744);
nor U4650 (N_4650,N_2008,N_1436);
nand U4651 (N_4651,N_2091,N_116);
or U4652 (N_4652,N_2717,N_715);
or U4653 (N_4653,N_2804,N_1334);
nand U4654 (N_4654,N_1402,N_1592);
or U4655 (N_4655,N_2532,N_131);
and U4656 (N_4656,N_1495,N_222);
nor U4657 (N_4657,N_2462,N_552);
nor U4658 (N_4658,N_2349,N_1277);
xnor U4659 (N_4659,N_432,N_1730);
or U4660 (N_4660,N_1174,N_1201);
nor U4661 (N_4661,N_2898,N_2839);
and U4662 (N_4662,N_1720,N_1895);
and U4663 (N_4663,N_632,N_2051);
nand U4664 (N_4664,N_2881,N_697);
or U4665 (N_4665,N_2498,N_2826);
nand U4666 (N_4666,N_1988,N_146);
xnor U4667 (N_4667,N_114,N_2080);
xnor U4668 (N_4668,N_1918,N_1189);
or U4669 (N_4669,N_2970,N_2120);
nand U4670 (N_4670,N_2332,N_2109);
nor U4671 (N_4671,N_367,N_153);
and U4672 (N_4672,N_1816,N_1737);
nand U4673 (N_4673,N_334,N_1478);
xnor U4674 (N_4674,N_718,N_1822);
nor U4675 (N_4675,N_1619,N_881);
and U4676 (N_4676,N_639,N_1309);
nand U4677 (N_4677,N_859,N_1834);
or U4678 (N_4678,N_1576,N_168);
and U4679 (N_4679,N_2421,N_1340);
nor U4680 (N_4680,N_2415,N_2362);
or U4681 (N_4681,N_2222,N_1634);
xor U4682 (N_4682,N_2521,N_1077);
or U4683 (N_4683,N_2895,N_169);
nor U4684 (N_4684,N_574,N_1798);
xnor U4685 (N_4685,N_2366,N_756);
xor U4686 (N_4686,N_318,N_343);
nor U4687 (N_4687,N_1130,N_1689);
nor U4688 (N_4688,N_110,N_2786);
or U4689 (N_4689,N_2881,N_20);
xnor U4690 (N_4690,N_2158,N_2502);
nor U4691 (N_4691,N_1584,N_1411);
xnor U4692 (N_4692,N_2221,N_594);
xor U4693 (N_4693,N_983,N_1902);
xor U4694 (N_4694,N_897,N_2281);
and U4695 (N_4695,N_2435,N_2905);
nand U4696 (N_4696,N_2560,N_2344);
or U4697 (N_4697,N_1564,N_1855);
or U4698 (N_4698,N_1720,N_1732);
nor U4699 (N_4699,N_2340,N_1439);
and U4700 (N_4700,N_2144,N_2071);
or U4701 (N_4701,N_1780,N_6);
xor U4702 (N_4702,N_31,N_40);
nor U4703 (N_4703,N_906,N_743);
nor U4704 (N_4704,N_823,N_1898);
nand U4705 (N_4705,N_1034,N_235);
nor U4706 (N_4706,N_1697,N_952);
xnor U4707 (N_4707,N_1204,N_410);
nand U4708 (N_4708,N_1177,N_1679);
xnor U4709 (N_4709,N_1297,N_296);
or U4710 (N_4710,N_275,N_574);
or U4711 (N_4711,N_2027,N_1159);
or U4712 (N_4712,N_2947,N_1644);
nor U4713 (N_4713,N_695,N_1940);
or U4714 (N_4714,N_1393,N_534);
and U4715 (N_4715,N_1566,N_1529);
or U4716 (N_4716,N_2345,N_2395);
nand U4717 (N_4717,N_641,N_569);
and U4718 (N_4718,N_2586,N_1827);
and U4719 (N_4719,N_2669,N_830);
or U4720 (N_4720,N_2812,N_1384);
nor U4721 (N_4721,N_2024,N_190);
nor U4722 (N_4722,N_786,N_2525);
or U4723 (N_4723,N_586,N_2140);
and U4724 (N_4724,N_1192,N_252);
and U4725 (N_4725,N_2598,N_2249);
nor U4726 (N_4726,N_2672,N_374);
nor U4727 (N_4727,N_2511,N_2309);
nand U4728 (N_4728,N_213,N_750);
nand U4729 (N_4729,N_539,N_1328);
xor U4730 (N_4730,N_2808,N_1106);
nand U4731 (N_4731,N_1320,N_2170);
and U4732 (N_4732,N_1399,N_1756);
nor U4733 (N_4733,N_761,N_2354);
and U4734 (N_4734,N_2113,N_541);
nand U4735 (N_4735,N_1541,N_573);
nor U4736 (N_4736,N_2280,N_1379);
and U4737 (N_4737,N_1151,N_2617);
xnor U4738 (N_4738,N_2625,N_2833);
nand U4739 (N_4739,N_167,N_1522);
nor U4740 (N_4740,N_920,N_1624);
and U4741 (N_4741,N_2354,N_1264);
xnor U4742 (N_4742,N_358,N_2796);
nand U4743 (N_4743,N_2716,N_963);
and U4744 (N_4744,N_945,N_1773);
nor U4745 (N_4745,N_686,N_1135);
xnor U4746 (N_4746,N_642,N_1195);
and U4747 (N_4747,N_523,N_2587);
nor U4748 (N_4748,N_2395,N_2071);
and U4749 (N_4749,N_1065,N_2797);
nand U4750 (N_4750,N_2201,N_377);
nand U4751 (N_4751,N_766,N_848);
nand U4752 (N_4752,N_1573,N_2689);
or U4753 (N_4753,N_2900,N_2200);
nor U4754 (N_4754,N_639,N_762);
xor U4755 (N_4755,N_1193,N_2907);
nor U4756 (N_4756,N_2034,N_1962);
nand U4757 (N_4757,N_2910,N_724);
and U4758 (N_4758,N_1614,N_404);
nor U4759 (N_4759,N_1176,N_2994);
and U4760 (N_4760,N_1092,N_104);
nand U4761 (N_4761,N_2924,N_504);
xor U4762 (N_4762,N_431,N_2303);
and U4763 (N_4763,N_2111,N_148);
nand U4764 (N_4764,N_2653,N_2226);
nor U4765 (N_4765,N_352,N_2690);
nand U4766 (N_4766,N_1808,N_2991);
or U4767 (N_4767,N_368,N_1403);
xnor U4768 (N_4768,N_1509,N_2);
nor U4769 (N_4769,N_1798,N_623);
xnor U4770 (N_4770,N_1404,N_471);
and U4771 (N_4771,N_1595,N_197);
and U4772 (N_4772,N_2421,N_2012);
nand U4773 (N_4773,N_1787,N_2208);
xnor U4774 (N_4774,N_1721,N_606);
xnor U4775 (N_4775,N_1118,N_1085);
nand U4776 (N_4776,N_1641,N_2885);
nand U4777 (N_4777,N_2141,N_510);
xor U4778 (N_4778,N_782,N_259);
and U4779 (N_4779,N_1369,N_2848);
and U4780 (N_4780,N_2377,N_1874);
or U4781 (N_4781,N_2037,N_2872);
or U4782 (N_4782,N_2136,N_329);
and U4783 (N_4783,N_1031,N_1956);
nor U4784 (N_4784,N_2673,N_565);
and U4785 (N_4785,N_498,N_1108);
and U4786 (N_4786,N_2491,N_1978);
and U4787 (N_4787,N_1351,N_1254);
xnor U4788 (N_4788,N_569,N_1626);
and U4789 (N_4789,N_286,N_1802);
xor U4790 (N_4790,N_2629,N_728);
and U4791 (N_4791,N_999,N_2325);
nand U4792 (N_4792,N_2098,N_1777);
and U4793 (N_4793,N_423,N_1121);
or U4794 (N_4794,N_709,N_66);
or U4795 (N_4795,N_813,N_1478);
xnor U4796 (N_4796,N_2667,N_2523);
nor U4797 (N_4797,N_969,N_227);
nor U4798 (N_4798,N_2473,N_2058);
nand U4799 (N_4799,N_257,N_1976);
nor U4800 (N_4800,N_1701,N_1508);
nand U4801 (N_4801,N_9,N_1873);
nor U4802 (N_4802,N_957,N_1768);
or U4803 (N_4803,N_2367,N_465);
nand U4804 (N_4804,N_1317,N_1473);
or U4805 (N_4805,N_294,N_30);
or U4806 (N_4806,N_572,N_800);
nor U4807 (N_4807,N_1828,N_2431);
nor U4808 (N_4808,N_562,N_2656);
nand U4809 (N_4809,N_1652,N_604);
nor U4810 (N_4810,N_1868,N_1913);
xor U4811 (N_4811,N_134,N_1478);
nand U4812 (N_4812,N_2745,N_1473);
nor U4813 (N_4813,N_387,N_837);
nor U4814 (N_4814,N_2811,N_293);
nand U4815 (N_4815,N_2912,N_2132);
nor U4816 (N_4816,N_2526,N_450);
xnor U4817 (N_4817,N_2340,N_988);
xnor U4818 (N_4818,N_1068,N_2595);
xnor U4819 (N_4819,N_299,N_2005);
and U4820 (N_4820,N_194,N_922);
and U4821 (N_4821,N_1767,N_1981);
or U4822 (N_4822,N_20,N_710);
nand U4823 (N_4823,N_829,N_109);
and U4824 (N_4824,N_2037,N_2691);
or U4825 (N_4825,N_914,N_2331);
nor U4826 (N_4826,N_2603,N_2169);
nand U4827 (N_4827,N_363,N_2377);
nor U4828 (N_4828,N_745,N_170);
nand U4829 (N_4829,N_2109,N_890);
or U4830 (N_4830,N_1438,N_2561);
xnor U4831 (N_4831,N_522,N_1963);
nand U4832 (N_4832,N_1480,N_289);
and U4833 (N_4833,N_1734,N_616);
nor U4834 (N_4834,N_2744,N_10);
or U4835 (N_4835,N_1672,N_2382);
and U4836 (N_4836,N_1604,N_478);
nor U4837 (N_4837,N_885,N_635);
or U4838 (N_4838,N_1804,N_2769);
xnor U4839 (N_4839,N_260,N_2483);
and U4840 (N_4840,N_1063,N_307);
nor U4841 (N_4841,N_2581,N_187);
or U4842 (N_4842,N_1460,N_487);
nand U4843 (N_4843,N_2557,N_2858);
or U4844 (N_4844,N_1661,N_1344);
nand U4845 (N_4845,N_1361,N_771);
nor U4846 (N_4846,N_2282,N_1598);
or U4847 (N_4847,N_2697,N_253);
and U4848 (N_4848,N_1750,N_1175);
nand U4849 (N_4849,N_2601,N_175);
nand U4850 (N_4850,N_2173,N_2775);
xor U4851 (N_4851,N_1100,N_712);
or U4852 (N_4852,N_2005,N_224);
nor U4853 (N_4853,N_2518,N_1046);
nand U4854 (N_4854,N_1824,N_2638);
nand U4855 (N_4855,N_636,N_1138);
and U4856 (N_4856,N_1095,N_1728);
nand U4857 (N_4857,N_2919,N_729);
nand U4858 (N_4858,N_1401,N_2570);
or U4859 (N_4859,N_2568,N_1182);
nor U4860 (N_4860,N_1435,N_2352);
nor U4861 (N_4861,N_1805,N_631);
nand U4862 (N_4862,N_863,N_689);
nor U4863 (N_4863,N_991,N_2703);
and U4864 (N_4864,N_1809,N_1664);
nand U4865 (N_4865,N_504,N_136);
or U4866 (N_4866,N_250,N_2936);
and U4867 (N_4867,N_1847,N_742);
nor U4868 (N_4868,N_2650,N_2114);
nor U4869 (N_4869,N_1977,N_2108);
or U4870 (N_4870,N_936,N_320);
nand U4871 (N_4871,N_1575,N_1118);
xnor U4872 (N_4872,N_1130,N_1073);
xor U4873 (N_4873,N_2476,N_143);
nor U4874 (N_4874,N_1570,N_757);
or U4875 (N_4875,N_2741,N_1210);
nor U4876 (N_4876,N_2676,N_2586);
nand U4877 (N_4877,N_1606,N_1541);
nand U4878 (N_4878,N_2659,N_1676);
nor U4879 (N_4879,N_1175,N_1453);
nor U4880 (N_4880,N_2100,N_375);
or U4881 (N_4881,N_2817,N_558);
and U4882 (N_4882,N_347,N_424);
nand U4883 (N_4883,N_2371,N_2668);
nand U4884 (N_4884,N_263,N_1287);
nand U4885 (N_4885,N_2435,N_2341);
nor U4886 (N_4886,N_2932,N_2064);
nand U4887 (N_4887,N_419,N_2867);
xor U4888 (N_4888,N_476,N_138);
xor U4889 (N_4889,N_1443,N_226);
or U4890 (N_4890,N_1598,N_432);
xnor U4891 (N_4891,N_2001,N_2902);
nand U4892 (N_4892,N_364,N_2833);
nor U4893 (N_4893,N_1965,N_2298);
nand U4894 (N_4894,N_733,N_1933);
xor U4895 (N_4895,N_1126,N_2186);
and U4896 (N_4896,N_1822,N_2892);
nand U4897 (N_4897,N_2386,N_2336);
and U4898 (N_4898,N_1436,N_2578);
nand U4899 (N_4899,N_2123,N_1616);
nand U4900 (N_4900,N_2104,N_2949);
nor U4901 (N_4901,N_692,N_84);
nor U4902 (N_4902,N_145,N_823);
or U4903 (N_4903,N_91,N_2698);
xor U4904 (N_4904,N_2610,N_441);
and U4905 (N_4905,N_2841,N_1599);
or U4906 (N_4906,N_2153,N_1518);
nor U4907 (N_4907,N_2502,N_1498);
and U4908 (N_4908,N_1044,N_1852);
nand U4909 (N_4909,N_817,N_1354);
nand U4910 (N_4910,N_146,N_1927);
nor U4911 (N_4911,N_2103,N_297);
xnor U4912 (N_4912,N_1499,N_127);
or U4913 (N_4913,N_767,N_868);
nand U4914 (N_4914,N_2289,N_191);
nor U4915 (N_4915,N_663,N_1271);
nand U4916 (N_4916,N_2916,N_2209);
xnor U4917 (N_4917,N_120,N_2519);
nand U4918 (N_4918,N_2159,N_1112);
nor U4919 (N_4919,N_2106,N_108);
and U4920 (N_4920,N_1201,N_1079);
xor U4921 (N_4921,N_363,N_946);
nand U4922 (N_4922,N_251,N_1402);
and U4923 (N_4923,N_1654,N_1796);
or U4924 (N_4924,N_2148,N_1594);
nand U4925 (N_4925,N_346,N_2781);
or U4926 (N_4926,N_87,N_1410);
and U4927 (N_4927,N_1543,N_1089);
nor U4928 (N_4928,N_1127,N_2592);
nand U4929 (N_4929,N_2322,N_1833);
xnor U4930 (N_4930,N_2732,N_1560);
or U4931 (N_4931,N_2053,N_1405);
and U4932 (N_4932,N_1414,N_2822);
nand U4933 (N_4933,N_2011,N_1701);
xnor U4934 (N_4934,N_1629,N_2845);
nand U4935 (N_4935,N_0,N_1408);
nand U4936 (N_4936,N_897,N_2303);
and U4937 (N_4937,N_347,N_1021);
or U4938 (N_4938,N_2270,N_1169);
nand U4939 (N_4939,N_1210,N_775);
or U4940 (N_4940,N_1118,N_2699);
xnor U4941 (N_4941,N_2827,N_224);
or U4942 (N_4942,N_1903,N_2448);
nor U4943 (N_4943,N_2028,N_285);
nor U4944 (N_4944,N_719,N_2770);
or U4945 (N_4945,N_610,N_1448);
xnor U4946 (N_4946,N_1459,N_942);
nor U4947 (N_4947,N_2489,N_170);
nor U4948 (N_4948,N_2476,N_2621);
nor U4949 (N_4949,N_1616,N_533);
and U4950 (N_4950,N_1473,N_2423);
and U4951 (N_4951,N_607,N_220);
xor U4952 (N_4952,N_575,N_921);
nand U4953 (N_4953,N_447,N_249);
and U4954 (N_4954,N_2003,N_398);
xor U4955 (N_4955,N_2127,N_2725);
and U4956 (N_4956,N_2668,N_1707);
nand U4957 (N_4957,N_1904,N_1748);
xnor U4958 (N_4958,N_197,N_2511);
or U4959 (N_4959,N_2746,N_2306);
nor U4960 (N_4960,N_2108,N_707);
nand U4961 (N_4961,N_1983,N_2933);
nand U4962 (N_4962,N_2936,N_2970);
nor U4963 (N_4963,N_135,N_2665);
xor U4964 (N_4964,N_2773,N_2559);
nor U4965 (N_4965,N_2865,N_1899);
xor U4966 (N_4966,N_1276,N_2621);
and U4967 (N_4967,N_446,N_2204);
nor U4968 (N_4968,N_2860,N_2124);
nor U4969 (N_4969,N_42,N_2525);
nor U4970 (N_4970,N_775,N_2737);
nor U4971 (N_4971,N_2355,N_1368);
xnor U4972 (N_4972,N_2268,N_1813);
xnor U4973 (N_4973,N_226,N_803);
or U4974 (N_4974,N_1726,N_2144);
or U4975 (N_4975,N_2730,N_251);
xnor U4976 (N_4976,N_1303,N_439);
and U4977 (N_4977,N_1563,N_1346);
nor U4978 (N_4978,N_136,N_774);
xor U4979 (N_4979,N_2670,N_882);
nand U4980 (N_4980,N_431,N_1254);
or U4981 (N_4981,N_2910,N_46);
or U4982 (N_4982,N_2816,N_414);
nor U4983 (N_4983,N_110,N_2825);
and U4984 (N_4984,N_358,N_593);
or U4985 (N_4985,N_166,N_2618);
or U4986 (N_4986,N_1381,N_2154);
or U4987 (N_4987,N_1061,N_2175);
or U4988 (N_4988,N_2594,N_1160);
nor U4989 (N_4989,N_543,N_1188);
nand U4990 (N_4990,N_2404,N_2445);
or U4991 (N_4991,N_2982,N_2939);
nand U4992 (N_4992,N_2746,N_1832);
and U4993 (N_4993,N_1200,N_1051);
or U4994 (N_4994,N_2789,N_1853);
and U4995 (N_4995,N_1513,N_188);
nor U4996 (N_4996,N_258,N_2438);
xnor U4997 (N_4997,N_2381,N_3);
nand U4998 (N_4998,N_2838,N_1473);
or U4999 (N_4999,N_430,N_2850);
xor U5000 (N_5000,N_471,N_932);
xor U5001 (N_5001,N_136,N_1513);
nand U5002 (N_5002,N_1840,N_1479);
or U5003 (N_5003,N_2345,N_838);
or U5004 (N_5004,N_2694,N_2148);
or U5005 (N_5005,N_1355,N_97);
or U5006 (N_5006,N_1664,N_1739);
nand U5007 (N_5007,N_2601,N_1434);
nand U5008 (N_5008,N_49,N_1821);
and U5009 (N_5009,N_1822,N_2172);
or U5010 (N_5010,N_1487,N_932);
nand U5011 (N_5011,N_1496,N_973);
nor U5012 (N_5012,N_1582,N_2202);
nand U5013 (N_5013,N_2421,N_1253);
nor U5014 (N_5014,N_433,N_1550);
and U5015 (N_5015,N_41,N_399);
xor U5016 (N_5016,N_1168,N_652);
nor U5017 (N_5017,N_140,N_1573);
nor U5018 (N_5018,N_607,N_2148);
or U5019 (N_5019,N_2158,N_762);
nor U5020 (N_5020,N_1274,N_2885);
and U5021 (N_5021,N_361,N_1144);
or U5022 (N_5022,N_2405,N_607);
xnor U5023 (N_5023,N_2654,N_1624);
or U5024 (N_5024,N_240,N_1025);
xnor U5025 (N_5025,N_867,N_2987);
nor U5026 (N_5026,N_1536,N_1961);
nor U5027 (N_5027,N_51,N_1861);
xnor U5028 (N_5028,N_329,N_1174);
and U5029 (N_5029,N_1738,N_1797);
and U5030 (N_5030,N_715,N_1541);
nor U5031 (N_5031,N_1665,N_251);
and U5032 (N_5032,N_1879,N_1222);
or U5033 (N_5033,N_423,N_1886);
nor U5034 (N_5034,N_2423,N_1503);
or U5035 (N_5035,N_2051,N_2645);
xor U5036 (N_5036,N_728,N_610);
nand U5037 (N_5037,N_1113,N_2762);
nand U5038 (N_5038,N_1916,N_1054);
nor U5039 (N_5039,N_902,N_2212);
nor U5040 (N_5040,N_442,N_739);
and U5041 (N_5041,N_1764,N_1878);
and U5042 (N_5042,N_1799,N_669);
nand U5043 (N_5043,N_2305,N_251);
nand U5044 (N_5044,N_2598,N_1195);
nand U5045 (N_5045,N_575,N_2182);
and U5046 (N_5046,N_1813,N_2170);
nor U5047 (N_5047,N_73,N_1303);
nor U5048 (N_5048,N_1666,N_2316);
or U5049 (N_5049,N_1510,N_2182);
nor U5050 (N_5050,N_1593,N_1586);
or U5051 (N_5051,N_1751,N_2789);
nor U5052 (N_5052,N_1037,N_445);
xor U5053 (N_5053,N_2430,N_2935);
nor U5054 (N_5054,N_686,N_455);
xor U5055 (N_5055,N_1907,N_87);
nor U5056 (N_5056,N_227,N_2999);
or U5057 (N_5057,N_1959,N_1540);
nand U5058 (N_5058,N_391,N_892);
and U5059 (N_5059,N_1069,N_716);
and U5060 (N_5060,N_2927,N_1408);
or U5061 (N_5061,N_290,N_404);
xnor U5062 (N_5062,N_671,N_333);
xor U5063 (N_5063,N_2202,N_2252);
and U5064 (N_5064,N_1950,N_755);
nand U5065 (N_5065,N_2349,N_1865);
and U5066 (N_5066,N_367,N_2806);
and U5067 (N_5067,N_2602,N_2066);
and U5068 (N_5068,N_2420,N_2074);
nand U5069 (N_5069,N_2624,N_133);
or U5070 (N_5070,N_952,N_845);
xnor U5071 (N_5071,N_879,N_2220);
or U5072 (N_5072,N_1465,N_933);
and U5073 (N_5073,N_730,N_2062);
xor U5074 (N_5074,N_2837,N_1805);
and U5075 (N_5075,N_2945,N_2894);
nor U5076 (N_5076,N_1714,N_1193);
nor U5077 (N_5077,N_1347,N_1464);
or U5078 (N_5078,N_2576,N_1125);
nand U5079 (N_5079,N_623,N_792);
nand U5080 (N_5080,N_811,N_976);
xor U5081 (N_5081,N_1718,N_2170);
nor U5082 (N_5082,N_2140,N_2517);
and U5083 (N_5083,N_926,N_2572);
and U5084 (N_5084,N_1578,N_1947);
nor U5085 (N_5085,N_1701,N_2418);
xor U5086 (N_5086,N_2952,N_2723);
xor U5087 (N_5087,N_932,N_560);
nand U5088 (N_5088,N_2490,N_1550);
or U5089 (N_5089,N_285,N_2218);
nand U5090 (N_5090,N_904,N_273);
or U5091 (N_5091,N_1034,N_1005);
xnor U5092 (N_5092,N_1013,N_2590);
xor U5093 (N_5093,N_2564,N_453);
nand U5094 (N_5094,N_1169,N_1736);
nor U5095 (N_5095,N_1075,N_2161);
nor U5096 (N_5096,N_1217,N_751);
nor U5097 (N_5097,N_1536,N_487);
nor U5098 (N_5098,N_2247,N_1859);
xor U5099 (N_5099,N_1720,N_2514);
and U5100 (N_5100,N_1873,N_2056);
nor U5101 (N_5101,N_1932,N_1254);
xor U5102 (N_5102,N_1179,N_1952);
and U5103 (N_5103,N_1256,N_1818);
and U5104 (N_5104,N_383,N_1766);
nor U5105 (N_5105,N_948,N_1776);
xor U5106 (N_5106,N_2050,N_801);
or U5107 (N_5107,N_1841,N_1093);
or U5108 (N_5108,N_2762,N_2350);
or U5109 (N_5109,N_339,N_1612);
nor U5110 (N_5110,N_391,N_1040);
xor U5111 (N_5111,N_28,N_2333);
or U5112 (N_5112,N_1910,N_65);
and U5113 (N_5113,N_1174,N_2045);
xnor U5114 (N_5114,N_1001,N_712);
or U5115 (N_5115,N_629,N_248);
nand U5116 (N_5116,N_567,N_2606);
nand U5117 (N_5117,N_68,N_2529);
nand U5118 (N_5118,N_2248,N_1159);
and U5119 (N_5119,N_2297,N_491);
nand U5120 (N_5120,N_1121,N_1315);
xor U5121 (N_5121,N_2323,N_1677);
and U5122 (N_5122,N_2305,N_940);
nand U5123 (N_5123,N_2576,N_311);
xnor U5124 (N_5124,N_2481,N_1489);
nor U5125 (N_5125,N_1662,N_2360);
and U5126 (N_5126,N_858,N_1008);
nor U5127 (N_5127,N_1745,N_1138);
nand U5128 (N_5128,N_2766,N_1782);
or U5129 (N_5129,N_628,N_2819);
or U5130 (N_5130,N_1760,N_1667);
xor U5131 (N_5131,N_2967,N_2406);
xnor U5132 (N_5132,N_2320,N_2875);
nand U5133 (N_5133,N_1740,N_262);
xor U5134 (N_5134,N_1477,N_670);
nor U5135 (N_5135,N_524,N_1768);
nor U5136 (N_5136,N_1880,N_2685);
nor U5137 (N_5137,N_2258,N_2151);
xor U5138 (N_5138,N_174,N_584);
or U5139 (N_5139,N_670,N_919);
nand U5140 (N_5140,N_461,N_2447);
xnor U5141 (N_5141,N_2983,N_148);
nor U5142 (N_5142,N_308,N_790);
or U5143 (N_5143,N_2778,N_556);
nor U5144 (N_5144,N_2180,N_277);
and U5145 (N_5145,N_1063,N_694);
xnor U5146 (N_5146,N_2702,N_1720);
or U5147 (N_5147,N_1050,N_2252);
nor U5148 (N_5148,N_112,N_2413);
and U5149 (N_5149,N_1030,N_1880);
or U5150 (N_5150,N_487,N_945);
and U5151 (N_5151,N_450,N_154);
xor U5152 (N_5152,N_2059,N_564);
xnor U5153 (N_5153,N_2293,N_2274);
xnor U5154 (N_5154,N_1386,N_1034);
xnor U5155 (N_5155,N_1531,N_1673);
nand U5156 (N_5156,N_2001,N_1576);
or U5157 (N_5157,N_606,N_1277);
and U5158 (N_5158,N_2453,N_47);
or U5159 (N_5159,N_2140,N_2440);
nor U5160 (N_5160,N_266,N_78);
or U5161 (N_5161,N_785,N_2048);
nand U5162 (N_5162,N_2554,N_2096);
and U5163 (N_5163,N_625,N_973);
xnor U5164 (N_5164,N_907,N_1107);
or U5165 (N_5165,N_2549,N_932);
or U5166 (N_5166,N_2643,N_19);
or U5167 (N_5167,N_2847,N_1257);
or U5168 (N_5168,N_492,N_754);
nor U5169 (N_5169,N_1359,N_797);
nor U5170 (N_5170,N_2016,N_292);
and U5171 (N_5171,N_2707,N_2557);
nand U5172 (N_5172,N_2458,N_278);
or U5173 (N_5173,N_302,N_2366);
xnor U5174 (N_5174,N_2703,N_1866);
and U5175 (N_5175,N_2480,N_2302);
xnor U5176 (N_5176,N_2757,N_717);
xor U5177 (N_5177,N_530,N_460);
or U5178 (N_5178,N_155,N_2196);
nor U5179 (N_5179,N_2343,N_1548);
xor U5180 (N_5180,N_441,N_268);
xor U5181 (N_5181,N_2271,N_2694);
and U5182 (N_5182,N_1461,N_351);
xnor U5183 (N_5183,N_2513,N_2991);
nand U5184 (N_5184,N_1374,N_325);
nand U5185 (N_5185,N_1442,N_2647);
nor U5186 (N_5186,N_263,N_1216);
nand U5187 (N_5187,N_2479,N_1110);
nor U5188 (N_5188,N_2381,N_773);
nand U5189 (N_5189,N_1021,N_2925);
or U5190 (N_5190,N_2695,N_2791);
xnor U5191 (N_5191,N_2160,N_2826);
or U5192 (N_5192,N_1663,N_1068);
and U5193 (N_5193,N_1429,N_2086);
xnor U5194 (N_5194,N_330,N_2264);
or U5195 (N_5195,N_2713,N_2721);
nand U5196 (N_5196,N_1604,N_1421);
nand U5197 (N_5197,N_2887,N_664);
nor U5198 (N_5198,N_655,N_1894);
or U5199 (N_5199,N_2602,N_1929);
and U5200 (N_5200,N_152,N_862);
nand U5201 (N_5201,N_987,N_1777);
or U5202 (N_5202,N_2841,N_1533);
or U5203 (N_5203,N_1858,N_2266);
xor U5204 (N_5204,N_2701,N_1833);
or U5205 (N_5205,N_797,N_551);
or U5206 (N_5206,N_1159,N_999);
nand U5207 (N_5207,N_15,N_926);
xor U5208 (N_5208,N_2168,N_2403);
xor U5209 (N_5209,N_1461,N_366);
and U5210 (N_5210,N_1781,N_1757);
and U5211 (N_5211,N_2230,N_2406);
xor U5212 (N_5212,N_1835,N_2173);
and U5213 (N_5213,N_1695,N_992);
nand U5214 (N_5214,N_1571,N_1486);
or U5215 (N_5215,N_1435,N_76);
nand U5216 (N_5216,N_1500,N_609);
nand U5217 (N_5217,N_1802,N_2604);
nor U5218 (N_5218,N_82,N_1303);
and U5219 (N_5219,N_2256,N_1132);
nand U5220 (N_5220,N_758,N_236);
xnor U5221 (N_5221,N_1956,N_1815);
nor U5222 (N_5222,N_1083,N_1275);
nor U5223 (N_5223,N_1409,N_2931);
nand U5224 (N_5224,N_2726,N_2734);
or U5225 (N_5225,N_2906,N_433);
nor U5226 (N_5226,N_2424,N_1656);
nand U5227 (N_5227,N_2232,N_512);
and U5228 (N_5228,N_1008,N_2457);
xnor U5229 (N_5229,N_2250,N_2641);
or U5230 (N_5230,N_2928,N_2273);
nand U5231 (N_5231,N_1444,N_2109);
xnor U5232 (N_5232,N_179,N_2833);
and U5233 (N_5233,N_851,N_1457);
xnor U5234 (N_5234,N_17,N_1623);
nor U5235 (N_5235,N_793,N_1065);
xnor U5236 (N_5236,N_2685,N_1032);
and U5237 (N_5237,N_1805,N_1884);
nor U5238 (N_5238,N_2816,N_2524);
or U5239 (N_5239,N_2517,N_190);
nor U5240 (N_5240,N_2859,N_459);
xnor U5241 (N_5241,N_426,N_71);
nor U5242 (N_5242,N_839,N_1876);
nand U5243 (N_5243,N_884,N_2217);
nand U5244 (N_5244,N_2460,N_2);
and U5245 (N_5245,N_2394,N_746);
or U5246 (N_5246,N_606,N_106);
or U5247 (N_5247,N_2098,N_1727);
and U5248 (N_5248,N_2389,N_2922);
nor U5249 (N_5249,N_1094,N_1519);
nor U5250 (N_5250,N_284,N_2594);
xnor U5251 (N_5251,N_200,N_2759);
nand U5252 (N_5252,N_624,N_16);
nand U5253 (N_5253,N_2551,N_359);
nand U5254 (N_5254,N_415,N_2976);
nor U5255 (N_5255,N_1911,N_2831);
and U5256 (N_5256,N_2280,N_2385);
nand U5257 (N_5257,N_205,N_1241);
xnor U5258 (N_5258,N_1740,N_2163);
nand U5259 (N_5259,N_2781,N_1103);
nand U5260 (N_5260,N_2272,N_689);
nand U5261 (N_5261,N_2492,N_2536);
and U5262 (N_5262,N_2505,N_2070);
xnor U5263 (N_5263,N_2932,N_2232);
nand U5264 (N_5264,N_2994,N_993);
or U5265 (N_5265,N_1719,N_1144);
xor U5266 (N_5266,N_512,N_2294);
and U5267 (N_5267,N_2486,N_1069);
xnor U5268 (N_5268,N_570,N_2554);
nor U5269 (N_5269,N_1298,N_2127);
xnor U5270 (N_5270,N_1897,N_1868);
nor U5271 (N_5271,N_556,N_2988);
or U5272 (N_5272,N_803,N_517);
xnor U5273 (N_5273,N_2371,N_2434);
and U5274 (N_5274,N_1612,N_2728);
or U5275 (N_5275,N_2403,N_2218);
nor U5276 (N_5276,N_2896,N_1783);
and U5277 (N_5277,N_1582,N_402);
nand U5278 (N_5278,N_1222,N_1272);
nand U5279 (N_5279,N_216,N_950);
and U5280 (N_5280,N_2657,N_2983);
or U5281 (N_5281,N_2349,N_596);
nor U5282 (N_5282,N_518,N_370);
xnor U5283 (N_5283,N_1917,N_2395);
and U5284 (N_5284,N_518,N_1107);
xnor U5285 (N_5285,N_759,N_2698);
or U5286 (N_5286,N_1952,N_1802);
nand U5287 (N_5287,N_2111,N_1552);
or U5288 (N_5288,N_1189,N_2244);
xnor U5289 (N_5289,N_1261,N_996);
nor U5290 (N_5290,N_2246,N_540);
or U5291 (N_5291,N_2627,N_2748);
nand U5292 (N_5292,N_2220,N_51);
or U5293 (N_5293,N_2515,N_1039);
or U5294 (N_5294,N_437,N_1455);
nor U5295 (N_5295,N_1844,N_2439);
xor U5296 (N_5296,N_1693,N_2505);
and U5297 (N_5297,N_1192,N_2606);
and U5298 (N_5298,N_1047,N_484);
nor U5299 (N_5299,N_486,N_869);
nor U5300 (N_5300,N_2368,N_810);
nand U5301 (N_5301,N_253,N_600);
xor U5302 (N_5302,N_395,N_1847);
nor U5303 (N_5303,N_2251,N_1003);
xor U5304 (N_5304,N_7,N_2980);
and U5305 (N_5305,N_2258,N_2664);
nand U5306 (N_5306,N_2942,N_413);
xnor U5307 (N_5307,N_1378,N_2931);
and U5308 (N_5308,N_2747,N_61);
nand U5309 (N_5309,N_1390,N_1904);
and U5310 (N_5310,N_672,N_1037);
or U5311 (N_5311,N_1445,N_1988);
and U5312 (N_5312,N_1917,N_2756);
nor U5313 (N_5313,N_1948,N_261);
and U5314 (N_5314,N_184,N_2166);
nor U5315 (N_5315,N_1826,N_2949);
nand U5316 (N_5316,N_65,N_1083);
nor U5317 (N_5317,N_600,N_2507);
and U5318 (N_5318,N_423,N_2067);
nor U5319 (N_5319,N_1947,N_562);
nor U5320 (N_5320,N_2305,N_528);
nand U5321 (N_5321,N_1205,N_977);
and U5322 (N_5322,N_1315,N_2940);
xnor U5323 (N_5323,N_2509,N_1270);
or U5324 (N_5324,N_880,N_2390);
nand U5325 (N_5325,N_1029,N_1856);
nor U5326 (N_5326,N_2753,N_2801);
xnor U5327 (N_5327,N_1387,N_2087);
xor U5328 (N_5328,N_1047,N_1400);
or U5329 (N_5329,N_1435,N_2236);
nor U5330 (N_5330,N_2464,N_2168);
nor U5331 (N_5331,N_1221,N_2572);
or U5332 (N_5332,N_1438,N_2592);
nand U5333 (N_5333,N_1115,N_2687);
and U5334 (N_5334,N_894,N_2420);
xor U5335 (N_5335,N_1019,N_1983);
xnor U5336 (N_5336,N_1581,N_2049);
or U5337 (N_5337,N_2378,N_1233);
or U5338 (N_5338,N_1531,N_1890);
or U5339 (N_5339,N_1775,N_2294);
xor U5340 (N_5340,N_779,N_1146);
xnor U5341 (N_5341,N_1300,N_172);
or U5342 (N_5342,N_2417,N_868);
nor U5343 (N_5343,N_203,N_2970);
nor U5344 (N_5344,N_1851,N_2415);
nor U5345 (N_5345,N_1383,N_2492);
or U5346 (N_5346,N_2087,N_68);
nor U5347 (N_5347,N_507,N_1694);
xor U5348 (N_5348,N_2757,N_410);
and U5349 (N_5349,N_2437,N_1724);
or U5350 (N_5350,N_2276,N_1858);
xnor U5351 (N_5351,N_749,N_598);
and U5352 (N_5352,N_1521,N_977);
nor U5353 (N_5353,N_1208,N_262);
xnor U5354 (N_5354,N_438,N_748);
nor U5355 (N_5355,N_2446,N_2419);
nand U5356 (N_5356,N_2080,N_1142);
nor U5357 (N_5357,N_2866,N_1195);
and U5358 (N_5358,N_2735,N_587);
nor U5359 (N_5359,N_908,N_699);
or U5360 (N_5360,N_1387,N_2287);
nor U5361 (N_5361,N_1449,N_913);
or U5362 (N_5362,N_2022,N_1576);
and U5363 (N_5363,N_2720,N_829);
and U5364 (N_5364,N_2156,N_878);
or U5365 (N_5365,N_1481,N_1797);
or U5366 (N_5366,N_748,N_566);
xnor U5367 (N_5367,N_1933,N_540);
or U5368 (N_5368,N_456,N_1897);
nand U5369 (N_5369,N_14,N_2269);
nand U5370 (N_5370,N_2597,N_2404);
xor U5371 (N_5371,N_2615,N_1196);
xnor U5372 (N_5372,N_1390,N_6);
nand U5373 (N_5373,N_611,N_1845);
nor U5374 (N_5374,N_469,N_161);
or U5375 (N_5375,N_483,N_120);
nor U5376 (N_5376,N_1811,N_1476);
or U5377 (N_5377,N_2004,N_2688);
nand U5378 (N_5378,N_352,N_1629);
nor U5379 (N_5379,N_1866,N_611);
nand U5380 (N_5380,N_97,N_2224);
nand U5381 (N_5381,N_1011,N_697);
and U5382 (N_5382,N_1386,N_1553);
nand U5383 (N_5383,N_1346,N_1991);
xor U5384 (N_5384,N_2512,N_2397);
nand U5385 (N_5385,N_2993,N_2509);
nor U5386 (N_5386,N_717,N_2039);
and U5387 (N_5387,N_812,N_2339);
xnor U5388 (N_5388,N_2796,N_676);
nand U5389 (N_5389,N_699,N_2936);
nand U5390 (N_5390,N_1898,N_1971);
xor U5391 (N_5391,N_1271,N_445);
and U5392 (N_5392,N_1972,N_2292);
nor U5393 (N_5393,N_1490,N_2917);
xor U5394 (N_5394,N_1519,N_729);
and U5395 (N_5395,N_528,N_1693);
nand U5396 (N_5396,N_1398,N_1808);
or U5397 (N_5397,N_425,N_2535);
or U5398 (N_5398,N_1736,N_2151);
and U5399 (N_5399,N_2960,N_1572);
or U5400 (N_5400,N_2982,N_2376);
nand U5401 (N_5401,N_917,N_1418);
and U5402 (N_5402,N_534,N_136);
nand U5403 (N_5403,N_919,N_1064);
and U5404 (N_5404,N_2754,N_1707);
xnor U5405 (N_5405,N_2951,N_2723);
nor U5406 (N_5406,N_1116,N_1589);
xnor U5407 (N_5407,N_2592,N_761);
nand U5408 (N_5408,N_1517,N_1929);
nor U5409 (N_5409,N_2578,N_2831);
nor U5410 (N_5410,N_2038,N_540);
or U5411 (N_5411,N_2364,N_84);
or U5412 (N_5412,N_2932,N_2664);
nor U5413 (N_5413,N_413,N_837);
nor U5414 (N_5414,N_2413,N_530);
xor U5415 (N_5415,N_638,N_1051);
nor U5416 (N_5416,N_137,N_2859);
nand U5417 (N_5417,N_2759,N_1027);
xor U5418 (N_5418,N_2140,N_2461);
nor U5419 (N_5419,N_2403,N_785);
xnor U5420 (N_5420,N_2181,N_2664);
or U5421 (N_5421,N_1711,N_479);
nand U5422 (N_5422,N_2927,N_291);
xor U5423 (N_5423,N_880,N_70);
xor U5424 (N_5424,N_174,N_1280);
or U5425 (N_5425,N_2459,N_2701);
nor U5426 (N_5426,N_1849,N_2114);
nand U5427 (N_5427,N_1519,N_2669);
nor U5428 (N_5428,N_712,N_1598);
and U5429 (N_5429,N_2631,N_746);
nand U5430 (N_5430,N_635,N_860);
and U5431 (N_5431,N_1402,N_824);
xor U5432 (N_5432,N_1291,N_625);
nor U5433 (N_5433,N_510,N_1011);
nand U5434 (N_5434,N_987,N_1273);
and U5435 (N_5435,N_2438,N_289);
nand U5436 (N_5436,N_134,N_2646);
nand U5437 (N_5437,N_424,N_2569);
xor U5438 (N_5438,N_852,N_1283);
and U5439 (N_5439,N_1071,N_453);
and U5440 (N_5440,N_2622,N_68);
nor U5441 (N_5441,N_2185,N_2528);
nor U5442 (N_5442,N_184,N_380);
or U5443 (N_5443,N_2283,N_794);
and U5444 (N_5444,N_2270,N_1702);
xor U5445 (N_5445,N_1256,N_2882);
nor U5446 (N_5446,N_1805,N_1453);
nor U5447 (N_5447,N_1439,N_1467);
or U5448 (N_5448,N_2055,N_460);
nand U5449 (N_5449,N_264,N_2593);
and U5450 (N_5450,N_1154,N_870);
nor U5451 (N_5451,N_1771,N_1708);
xnor U5452 (N_5452,N_168,N_224);
nand U5453 (N_5453,N_229,N_53);
xnor U5454 (N_5454,N_2414,N_1383);
nand U5455 (N_5455,N_707,N_2326);
xor U5456 (N_5456,N_562,N_2563);
nor U5457 (N_5457,N_2039,N_1615);
xor U5458 (N_5458,N_1788,N_184);
or U5459 (N_5459,N_2902,N_1377);
nand U5460 (N_5460,N_2298,N_1731);
nor U5461 (N_5461,N_695,N_322);
and U5462 (N_5462,N_2470,N_211);
nand U5463 (N_5463,N_920,N_2703);
or U5464 (N_5464,N_1943,N_2912);
xor U5465 (N_5465,N_261,N_818);
nor U5466 (N_5466,N_1686,N_1546);
nor U5467 (N_5467,N_1924,N_2531);
and U5468 (N_5468,N_2229,N_1081);
and U5469 (N_5469,N_1404,N_1591);
and U5470 (N_5470,N_1706,N_365);
or U5471 (N_5471,N_1121,N_1477);
and U5472 (N_5472,N_183,N_334);
and U5473 (N_5473,N_242,N_1682);
or U5474 (N_5474,N_678,N_2986);
xor U5475 (N_5475,N_846,N_442);
xnor U5476 (N_5476,N_2794,N_2070);
xnor U5477 (N_5477,N_2039,N_1120);
xor U5478 (N_5478,N_2568,N_629);
xnor U5479 (N_5479,N_1247,N_869);
nand U5480 (N_5480,N_2482,N_2170);
nand U5481 (N_5481,N_1151,N_2569);
xor U5482 (N_5482,N_2788,N_209);
nor U5483 (N_5483,N_2189,N_2327);
or U5484 (N_5484,N_2951,N_2032);
and U5485 (N_5485,N_908,N_2735);
nand U5486 (N_5486,N_2770,N_2985);
xnor U5487 (N_5487,N_983,N_2970);
or U5488 (N_5488,N_1714,N_1464);
and U5489 (N_5489,N_2694,N_840);
nand U5490 (N_5490,N_903,N_1363);
nor U5491 (N_5491,N_1235,N_2527);
nand U5492 (N_5492,N_2937,N_720);
nor U5493 (N_5493,N_1455,N_1253);
xnor U5494 (N_5494,N_1832,N_1965);
nand U5495 (N_5495,N_541,N_207);
and U5496 (N_5496,N_928,N_1152);
xnor U5497 (N_5497,N_357,N_1439);
or U5498 (N_5498,N_1005,N_2228);
and U5499 (N_5499,N_2697,N_2046);
xor U5500 (N_5500,N_2709,N_1532);
xnor U5501 (N_5501,N_101,N_1895);
and U5502 (N_5502,N_1425,N_329);
nand U5503 (N_5503,N_1338,N_1933);
nor U5504 (N_5504,N_2602,N_1778);
and U5505 (N_5505,N_471,N_2054);
or U5506 (N_5506,N_2616,N_887);
or U5507 (N_5507,N_123,N_2947);
and U5508 (N_5508,N_470,N_15);
nor U5509 (N_5509,N_1218,N_652);
and U5510 (N_5510,N_2258,N_782);
xnor U5511 (N_5511,N_2680,N_710);
nand U5512 (N_5512,N_1322,N_1410);
nor U5513 (N_5513,N_802,N_2013);
nor U5514 (N_5514,N_858,N_1729);
or U5515 (N_5515,N_2169,N_1211);
nor U5516 (N_5516,N_541,N_2881);
nor U5517 (N_5517,N_1727,N_1519);
xor U5518 (N_5518,N_2783,N_785);
or U5519 (N_5519,N_2016,N_2303);
nor U5520 (N_5520,N_2635,N_2082);
and U5521 (N_5521,N_265,N_143);
nor U5522 (N_5522,N_2917,N_1797);
or U5523 (N_5523,N_745,N_1023);
and U5524 (N_5524,N_856,N_2960);
nor U5525 (N_5525,N_46,N_673);
or U5526 (N_5526,N_1329,N_1350);
nand U5527 (N_5527,N_21,N_827);
or U5528 (N_5528,N_2818,N_1241);
nand U5529 (N_5529,N_2544,N_2464);
and U5530 (N_5530,N_1874,N_282);
or U5531 (N_5531,N_823,N_2299);
nand U5532 (N_5532,N_2032,N_165);
and U5533 (N_5533,N_2392,N_2836);
nor U5534 (N_5534,N_806,N_1418);
or U5535 (N_5535,N_2691,N_1131);
nand U5536 (N_5536,N_2347,N_1415);
or U5537 (N_5537,N_81,N_859);
nand U5538 (N_5538,N_409,N_904);
xnor U5539 (N_5539,N_1921,N_857);
nand U5540 (N_5540,N_4,N_1542);
nor U5541 (N_5541,N_1008,N_317);
nor U5542 (N_5542,N_381,N_148);
nor U5543 (N_5543,N_717,N_1776);
xnor U5544 (N_5544,N_1060,N_2951);
or U5545 (N_5545,N_2979,N_2239);
and U5546 (N_5546,N_1250,N_711);
nor U5547 (N_5547,N_2444,N_1694);
nand U5548 (N_5548,N_1332,N_2448);
or U5549 (N_5549,N_812,N_883);
or U5550 (N_5550,N_888,N_2457);
or U5551 (N_5551,N_1773,N_1914);
nor U5552 (N_5552,N_479,N_875);
and U5553 (N_5553,N_978,N_123);
nor U5554 (N_5554,N_2017,N_2515);
nor U5555 (N_5555,N_507,N_966);
or U5556 (N_5556,N_2509,N_418);
nand U5557 (N_5557,N_2907,N_2931);
or U5558 (N_5558,N_2377,N_1264);
xnor U5559 (N_5559,N_462,N_2318);
or U5560 (N_5560,N_2264,N_1878);
nand U5561 (N_5561,N_365,N_486);
nor U5562 (N_5562,N_2783,N_2127);
nor U5563 (N_5563,N_1035,N_1319);
nand U5564 (N_5564,N_1566,N_2962);
nor U5565 (N_5565,N_2923,N_749);
or U5566 (N_5566,N_2536,N_2791);
xor U5567 (N_5567,N_1166,N_1778);
and U5568 (N_5568,N_2242,N_224);
xnor U5569 (N_5569,N_1491,N_2087);
and U5570 (N_5570,N_333,N_2647);
and U5571 (N_5571,N_527,N_714);
xor U5572 (N_5572,N_653,N_1713);
nand U5573 (N_5573,N_2923,N_2174);
xnor U5574 (N_5574,N_1607,N_42);
or U5575 (N_5575,N_1321,N_1354);
xnor U5576 (N_5576,N_590,N_2067);
nand U5577 (N_5577,N_10,N_2895);
xor U5578 (N_5578,N_1381,N_2113);
nor U5579 (N_5579,N_1383,N_295);
nor U5580 (N_5580,N_2832,N_1512);
nor U5581 (N_5581,N_602,N_210);
xor U5582 (N_5582,N_1164,N_2311);
xor U5583 (N_5583,N_2692,N_132);
and U5584 (N_5584,N_2037,N_2956);
nand U5585 (N_5585,N_2227,N_2266);
nand U5586 (N_5586,N_1513,N_2783);
nand U5587 (N_5587,N_970,N_1879);
nor U5588 (N_5588,N_872,N_152);
xnor U5589 (N_5589,N_705,N_2145);
xor U5590 (N_5590,N_519,N_2182);
nor U5591 (N_5591,N_810,N_2682);
nor U5592 (N_5592,N_1713,N_2240);
nand U5593 (N_5593,N_1281,N_1693);
and U5594 (N_5594,N_1794,N_1221);
nor U5595 (N_5595,N_1036,N_1882);
nand U5596 (N_5596,N_2334,N_989);
nor U5597 (N_5597,N_1077,N_630);
nor U5598 (N_5598,N_1504,N_1168);
xnor U5599 (N_5599,N_1031,N_2356);
or U5600 (N_5600,N_10,N_1938);
or U5601 (N_5601,N_1561,N_2175);
nand U5602 (N_5602,N_2819,N_841);
and U5603 (N_5603,N_932,N_1472);
and U5604 (N_5604,N_2499,N_2380);
nand U5605 (N_5605,N_933,N_2280);
or U5606 (N_5606,N_1482,N_987);
or U5607 (N_5607,N_1510,N_2261);
or U5608 (N_5608,N_1655,N_2340);
nand U5609 (N_5609,N_1441,N_1973);
xnor U5610 (N_5610,N_2803,N_2561);
and U5611 (N_5611,N_1682,N_2275);
and U5612 (N_5612,N_1057,N_1133);
nand U5613 (N_5613,N_1827,N_335);
and U5614 (N_5614,N_1967,N_1327);
nor U5615 (N_5615,N_2164,N_642);
and U5616 (N_5616,N_934,N_609);
nor U5617 (N_5617,N_2466,N_136);
and U5618 (N_5618,N_2002,N_1072);
xor U5619 (N_5619,N_897,N_1600);
xor U5620 (N_5620,N_2471,N_28);
nor U5621 (N_5621,N_833,N_649);
and U5622 (N_5622,N_1341,N_17);
xnor U5623 (N_5623,N_1577,N_2099);
xor U5624 (N_5624,N_235,N_1282);
nand U5625 (N_5625,N_1462,N_292);
nand U5626 (N_5626,N_2052,N_660);
or U5627 (N_5627,N_41,N_1753);
xor U5628 (N_5628,N_1550,N_345);
nor U5629 (N_5629,N_760,N_113);
nand U5630 (N_5630,N_1927,N_956);
nor U5631 (N_5631,N_447,N_2737);
or U5632 (N_5632,N_2514,N_2309);
and U5633 (N_5633,N_1612,N_864);
and U5634 (N_5634,N_2678,N_499);
xor U5635 (N_5635,N_2879,N_1942);
or U5636 (N_5636,N_2591,N_1816);
xnor U5637 (N_5637,N_1307,N_1653);
and U5638 (N_5638,N_1650,N_340);
nor U5639 (N_5639,N_925,N_2149);
xor U5640 (N_5640,N_2238,N_1355);
nand U5641 (N_5641,N_761,N_2781);
or U5642 (N_5642,N_429,N_2988);
or U5643 (N_5643,N_89,N_875);
nand U5644 (N_5644,N_1319,N_2143);
and U5645 (N_5645,N_1484,N_1257);
nand U5646 (N_5646,N_213,N_498);
and U5647 (N_5647,N_1064,N_506);
nor U5648 (N_5648,N_816,N_2807);
or U5649 (N_5649,N_1655,N_1634);
and U5650 (N_5650,N_1571,N_1610);
nand U5651 (N_5651,N_2924,N_698);
nand U5652 (N_5652,N_2132,N_2597);
or U5653 (N_5653,N_2950,N_1156);
or U5654 (N_5654,N_2637,N_2108);
and U5655 (N_5655,N_330,N_1309);
or U5656 (N_5656,N_2171,N_1520);
and U5657 (N_5657,N_132,N_945);
nand U5658 (N_5658,N_2948,N_2783);
xnor U5659 (N_5659,N_2542,N_1088);
or U5660 (N_5660,N_2203,N_2465);
and U5661 (N_5661,N_2057,N_516);
xor U5662 (N_5662,N_2059,N_1039);
and U5663 (N_5663,N_1806,N_694);
and U5664 (N_5664,N_286,N_2133);
or U5665 (N_5665,N_567,N_616);
nor U5666 (N_5666,N_2547,N_472);
nand U5667 (N_5667,N_2758,N_1918);
xor U5668 (N_5668,N_2401,N_894);
and U5669 (N_5669,N_707,N_113);
nor U5670 (N_5670,N_2052,N_2764);
nand U5671 (N_5671,N_1648,N_1055);
or U5672 (N_5672,N_1783,N_2086);
and U5673 (N_5673,N_1787,N_2437);
and U5674 (N_5674,N_1795,N_1740);
nor U5675 (N_5675,N_1435,N_1274);
xor U5676 (N_5676,N_173,N_1614);
or U5677 (N_5677,N_503,N_2358);
nor U5678 (N_5678,N_1919,N_2224);
and U5679 (N_5679,N_734,N_1128);
or U5680 (N_5680,N_682,N_2056);
nand U5681 (N_5681,N_2541,N_438);
xor U5682 (N_5682,N_513,N_2883);
or U5683 (N_5683,N_708,N_728);
nor U5684 (N_5684,N_2629,N_976);
or U5685 (N_5685,N_2500,N_281);
xnor U5686 (N_5686,N_2882,N_1900);
nor U5687 (N_5687,N_244,N_2264);
and U5688 (N_5688,N_1980,N_594);
nand U5689 (N_5689,N_2375,N_2052);
xor U5690 (N_5690,N_55,N_1620);
nand U5691 (N_5691,N_836,N_2361);
nand U5692 (N_5692,N_246,N_1216);
xor U5693 (N_5693,N_1724,N_1205);
or U5694 (N_5694,N_254,N_1503);
nor U5695 (N_5695,N_1585,N_1270);
nand U5696 (N_5696,N_1594,N_556);
nand U5697 (N_5697,N_2947,N_2400);
nor U5698 (N_5698,N_119,N_748);
xor U5699 (N_5699,N_2824,N_1950);
and U5700 (N_5700,N_177,N_452);
xnor U5701 (N_5701,N_843,N_2480);
nand U5702 (N_5702,N_174,N_566);
xnor U5703 (N_5703,N_1371,N_2252);
nand U5704 (N_5704,N_800,N_2111);
nor U5705 (N_5705,N_266,N_1278);
and U5706 (N_5706,N_1850,N_2779);
or U5707 (N_5707,N_3,N_2137);
xnor U5708 (N_5708,N_758,N_1897);
nor U5709 (N_5709,N_992,N_2700);
nand U5710 (N_5710,N_1096,N_1590);
nand U5711 (N_5711,N_664,N_1544);
nand U5712 (N_5712,N_2146,N_1605);
or U5713 (N_5713,N_967,N_999);
and U5714 (N_5714,N_2679,N_812);
and U5715 (N_5715,N_1276,N_2512);
nand U5716 (N_5716,N_730,N_1065);
xor U5717 (N_5717,N_43,N_1120);
and U5718 (N_5718,N_1009,N_1809);
xnor U5719 (N_5719,N_2022,N_41);
or U5720 (N_5720,N_1748,N_2561);
or U5721 (N_5721,N_607,N_1380);
and U5722 (N_5722,N_1681,N_446);
nand U5723 (N_5723,N_2206,N_1404);
or U5724 (N_5724,N_2148,N_6);
xor U5725 (N_5725,N_1465,N_2995);
or U5726 (N_5726,N_1213,N_2944);
or U5727 (N_5727,N_1440,N_2510);
nand U5728 (N_5728,N_361,N_2457);
and U5729 (N_5729,N_1861,N_1388);
and U5730 (N_5730,N_23,N_2677);
or U5731 (N_5731,N_815,N_1424);
nand U5732 (N_5732,N_1024,N_2474);
nor U5733 (N_5733,N_2455,N_2655);
or U5734 (N_5734,N_1542,N_1915);
nor U5735 (N_5735,N_291,N_1648);
nor U5736 (N_5736,N_1282,N_1089);
nor U5737 (N_5737,N_264,N_2022);
xor U5738 (N_5738,N_1261,N_1081);
and U5739 (N_5739,N_1925,N_445);
and U5740 (N_5740,N_1205,N_2317);
or U5741 (N_5741,N_2806,N_186);
nand U5742 (N_5742,N_1633,N_2846);
nor U5743 (N_5743,N_1398,N_348);
xor U5744 (N_5744,N_2771,N_2294);
and U5745 (N_5745,N_1386,N_1162);
xnor U5746 (N_5746,N_2364,N_256);
and U5747 (N_5747,N_1932,N_1231);
nand U5748 (N_5748,N_1377,N_166);
or U5749 (N_5749,N_357,N_1014);
nand U5750 (N_5750,N_1249,N_2877);
nor U5751 (N_5751,N_554,N_359);
xnor U5752 (N_5752,N_2748,N_271);
nand U5753 (N_5753,N_1047,N_2383);
nand U5754 (N_5754,N_1024,N_309);
xor U5755 (N_5755,N_753,N_2222);
nand U5756 (N_5756,N_420,N_365);
and U5757 (N_5757,N_2844,N_2044);
nor U5758 (N_5758,N_904,N_2701);
nor U5759 (N_5759,N_1625,N_1472);
nor U5760 (N_5760,N_1552,N_765);
nor U5761 (N_5761,N_1506,N_2818);
and U5762 (N_5762,N_2529,N_1905);
and U5763 (N_5763,N_537,N_1096);
or U5764 (N_5764,N_1423,N_1254);
xor U5765 (N_5765,N_1859,N_1692);
and U5766 (N_5766,N_1985,N_913);
nand U5767 (N_5767,N_2741,N_768);
and U5768 (N_5768,N_513,N_765);
nand U5769 (N_5769,N_1383,N_1089);
xor U5770 (N_5770,N_552,N_66);
or U5771 (N_5771,N_2133,N_432);
nand U5772 (N_5772,N_2027,N_2178);
and U5773 (N_5773,N_1875,N_264);
or U5774 (N_5774,N_2006,N_242);
or U5775 (N_5775,N_1942,N_620);
or U5776 (N_5776,N_934,N_2303);
xnor U5777 (N_5777,N_783,N_1175);
or U5778 (N_5778,N_2780,N_156);
or U5779 (N_5779,N_408,N_58);
and U5780 (N_5780,N_1227,N_225);
and U5781 (N_5781,N_500,N_2071);
nand U5782 (N_5782,N_1977,N_2500);
nand U5783 (N_5783,N_2547,N_1348);
xor U5784 (N_5784,N_924,N_3);
and U5785 (N_5785,N_1587,N_659);
and U5786 (N_5786,N_2740,N_204);
and U5787 (N_5787,N_1050,N_1719);
nand U5788 (N_5788,N_269,N_2820);
nor U5789 (N_5789,N_1285,N_2383);
or U5790 (N_5790,N_2281,N_438);
xor U5791 (N_5791,N_1810,N_2347);
or U5792 (N_5792,N_1543,N_2089);
or U5793 (N_5793,N_925,N_2716);
nand U5794 (N_5794,N_506,N_297);
nor U5795 (N_5795,N_2325,N_2267);
xor U5796 (N_5796,N_1828,N_2973);
and U5797 (N_5797,N_246,N_504);
xnor U5798 (N_5798,N_2942,N_332);
xor U5799 (N_5799,N_1231,N_1776);
xor U5800 (N_5800,N_635,N_423);
or U5801 (N_5801,N_2424,N_1940);
or U5802 (N_5802,N_2857,N_2635);
xor U5803 (N_5803,N_572,N_1762);
and U5804 (N_5804,N_2280,N_1442);
xnor U5805 (N_5805,N_2256,N_2616);
xnor U5806 (N_5806,N_341,N_1018);
or U5807 (N_5807,N_1789,N_419);
nor U5808 (N_5808,N_730,N_635);
and U5809 (N_5809,N_1920,N_2869);
nor U5810 (N_5810,N_948,N_1609);
and U5811 (N_5811,N_1696,N_40);
nand U5812 (N_5812,N_2588,N_2035);
or U5813 (N_5813,N_708,N_1711);
and U5814 (N_5814,N_2921,N_2365);
xnor U5815 (N_5815,N_550,N_1855);
nand U5816 (N_5816,N_2624,N_1114);
nand U5817 (N_5817,N_2609,N_2797);
nand U5818 (N_5818,N_2611,N_381);
xor U5819 (N_5819,N_1154,N_2055);
nand U5820 (N_5820,N_2784,N_2980);
nor U5821 (N_5821,N_164,N_1782);
xnor U5822 (N_5822,N_716,N_1113);
and U5823 (N_5823,N_1541,N_1762);
and U5824 (N_5824,N_2159,N_1019);
and U5825 (N_5825,N_1360,N_199);
xor U5826 (N_5826,N_2145,N_422);
or U5827 (N_5827,N_370,N_2926);
or U5828 (N_5828,N_2827,N_706);
or U5829 (N_5829,N_623,N_1875);
and U5830 (N_5830,N_2563,N_428);
nand U5831 (N_5831,N_2411,N_922);
xor U5832 (N_5832,N_901,N_111);
xor U5833 (N_5833,N_1171,N_2521);
xor U5834 (N_5834,N_2131,N_1969);
or U5835 (N_5835,N_817,N_2533);
nand U5836 (N_5836,N_907,N_673);
and U5837 (N_5837,N_232,N_1267);
nor U5838 (N_5838,N_2406,N_1359);
xnor U5839 (N_5839,N_2574,N_715);
nand U5840 (N_5840,N_2416,N_2525);
nor U5841 (N_5841,N_761,N_336);
or U5842 (N_5842,N_890,N_767);
or U5843 (N_5843,N_1378,N_658);
nor U5844 (N_5844,N_441,N_1433);
nand U5845 (N_5845,N_2851,N_659);
and U5846 (N_5846,N_1116,N_2638);
nand U5847 (N_5847,N_1278,N_726);
or U5848 (N_5848,N_2619,N_2167);
and U5849 (N_5849,N_742,N_1202);
xnor U5850 (N_5850,N_225,N_1410);
nand U5851 (N_5851,N_521,N_1638);
and U5852 (N_5852,N_2116,N_715);
nor U5853 (N_5853,N_993,N_1263);
and U5854 (N_5854,N_688,N_2670);
and U5855 (N_5855,N_2223,N_1339);
and U5856 (N_5856,N_1645,N_2501);
xnor U5857 (N_5857,N_1547,N_724);
and U5858 (N_5858,N_986,N_2537);
xor U5859 (N_5859,N_1396,N_502);
and U5860 (N_5860,N_2820,N_267);
and U5861 (N_5861,N_2584,N_2066);
and U5862 (N_5862,N_1527,N_670);
or U5863 (N_5863,N_1544,N_1816);
xnor U5864 (N_5864,N_2016,N_1797);
xor U5865 (N_5865,N_329,N_2);
nor U5866 (N_5866,N_2540,N_656);
or U5867 (N_5867,N_698,N_2458);
and U5868 (N_5868,N_1134,N_1443);
xnor U5869 (N_5869,N_1200,N_2464);
or U5870 (N_5870,N_1178,N_1036);
nand U5871 (N_5871,N_1859,N_2119);
xnor U5872 (N_5872,N_2043,N_1054);
nor U5873 (N_5873,N_2958,N_636);
and U5874 (N_5874,N_357,N_1765);
and U5875 (N_5875,N_1284,N_1875);
nor U5876 (N_5876,N_485,N_194);
xor U5877 (N_5877,N_2510,N_2469);
nand U5878 (N_5878,N_749,N_1572);
xnor U5879 (N_5879,N_1831,N_2256);
xnor U5880 (N_5880,N_2469,N_2268);
nand U5881 (N_5881,N_1118,N_2973);
xor U5882 (N_5882,N_1660,N_543);
xnor U5883 (N_5883,N_1006,N_306);
xor U5884 (N_5884,N_214,N_701);
and U5885 (N_5885,N_32,N_1157);
or U5886 (N_5886,N_1851,N_1750);
and U5887 (N_5887,N_2961,N_2604);
nand U5888 (N_5888,N_1946,N_2999);
xor U5889 (N_5889,N_470,N_572);
xor U5890 (N_5890,N_1532,N_948);
nand U5891 (N_5891,N_582,N_2976);
nor U5892 (N_5892,N_1163,N_304);
and U5893 (N_5893,N_1154,N_1267);
and U5894 (N_5894,N_2315,N_724);
xor U5895 (N_5895,N_1974,N_2551);
xnor U5896 (N_5896,N_1038,N_285);
nor U5897 (N_5897,N_1273,N_1051);
nand U5898 (N_5898,N_397,N_2338);
and U5899 (N_5899,N_2297,N_1474);
xnor U5900 (N_5900,N_1109,N_656);
xor U5901 (N_5901,N_2970,N_2573);
nor U5902 (N_5902,N_2436,N_1875);
nor U5903 (N_5903,N_2626,N_579);
nand U5904 (N_5904,N_253,N_801);
nand U5905 (N_5905,N_1666,N_2881);
nand U5906 (N_5906,N_2584,N_1285);
and U5907 (N_5907,N_2066,N_2087);
and U5908 (N_5908,N_2947,N_1022);
nand U5909 (N_5909,N_505,N_2250);
xor U5910 (N_5910,N_1276,N_111);
nand U5911 (N_5911,N_805,N_1634);
xnor U5912 (N_5912,N_161,N_450);
nor U5913 (N_5913,N_2919,N_2859);
nand U5914 (N_5914,N_1266,N_1508);
and U5915 (N_5915,N_1206,N_1572);
and U5916 (N_5916,N_734,N_1180);
and U5917 (N_5917,N_2943,N_61);
nand U5918 (N_5918,N_2815,N_2898);
or U5919 (N_5919,N_2267,N_1748);
nand U5920 (N_5920,N_2345,N_2063);
xor U5921 (N_5921,N_2822,N_2211);
or U5922 (N_5922,N_1553,N_225);
and U5923 (N_5923,N_628,N_1042);
and U5924 (N_5924,N_975,N_2997);
nor U5925 (N_5925,N_2195,N_362);
xnor U5926 (N_5926,N_1979,N_2839);
or U5927 (N_5927,N_805,N_2982);
or U5928 (N_5928,N_2816,N_1264);
nand U5929 (N_5929,N_2640,N_1196);
or U5930 (N_5930,N_960,N_103);
or U5931 (N_5931,N_30,N_1410);
nand U5932 (N_5932,N_481,N_2894);
and U5933 (N_5933,N_505,N_2105);
nand U5934 (N_5934,N_1719,N_839);
or U5935 (N_5935,N_874,N_803);
nor U5936 (N_5936,N_2799,N_28);
xor U5937 (N_5937,N_1387,N_1767);
and U5938 (N_5938,N_1950,N_354);
nor U5939 (N_5939,N_2244,N_1431);
nand U5940 (N_5940,N_1039,N_737);
or U5941 (N_5941,N_2660,N_585);
or U5942 (N_5942,N_1391,N_2486);
xor U5943 (N_5943,N_1342,N_2236);
and U5944 (N_5944,N_2423,N_47);
nor U5945 (N_5945,N_695,N_1098);
or U5946 (N_5946,N_715,N_1942);
nor U5947 (N_5947,N_1235,N_1997);
nor U5948 (N_5948,N_1791,N_1804);
nand U5949 (N_5949,N_1152,N_943);
xnor U5950 (N_5950,N_1177,N_2078);
nand U5951 (N_5951,N_2177,N_2975);
or U5952 (N_5952,N_763,N_1752);
or U5953 (N_5953,N_2482,N_1040);
or U5954 (N_5954,N_416,N_2741);
nor U5955 (N_5955,N_555,N_1112);
nor U5956 (N_5956,N_1615,N_2318);
or U5957 (N_5957,N_1565,N_1814);
nand U5958 (N_5958,N_841,N_1603);
or U5959 (N_5959,N_1,N_288);
and U5960 (N_5960,N_382,N_787);
nand U5961 (N_5961,N_1993,N_1059);
and U5962 (N_5962,N_2731,N_2473);
or U5963 (N_5963,N_1157,N_2591);
or U5964 (N_5964,N_634,N_2474);
nor U5965 (N_5965,N_2574,N_2188);
xnor U5966 (N_5966,N_2482,N_493);
nand U5967 (N_5967,N_1365,N_823);
nor U5968 (N_5968,N_2222,N_2585);
xnor U5969 (N_5969,N_1812,N_2280);
xor U5970 (N_5970,N_216,N_979);
nor U5971 (N_5971,N_56,N_2263);
nand U5972 (N_5972,N_2404,N_989);
nand U5973 (N_5973,N_367,N_130);
nor U5974 (N_5974,N_605,N_3);
and U5975 (N_5975,N_2688,N_2259);
nand U5976 (N_5976,N_123,N_829);
nand U5977 (N_5977,N_167,N_2102);
nor U5978 (N_5978,N_1022,N_1671);
or U5979 (N_5979,N_2492,N_559);
nand U5980 (N_5980,N_1154,N_2277);
or U5981 (N_5981,N_2816,N_1634);
or U5982 (N_5982,N_1446,N_425);
and U5983 (N_5983,N_1005,N_744);
xnor U5984 (N_5984,N_588,N_104);
nand U5985 (N_5985,N_248,N_1154);
nand U5986 (N_5986,N_308,N_1464);
nor U5987 (N_5987,N_425,N_1860);
xor U5988 (N_5988,N_2583,N_734);
xor U5989 (N_5989,N_26,N_2549);
xor U5990 (N_5990,N_1176,N_1471);
nand U5991 (N_5991,N_1624,N_562);
or U5992 (N_5992,N_2172,N_993);
nand U5993 (N_5993,N_385,N_103);
and U5994 (N_5994,N_175,N_2244);
nor U5995 (N_5995,N_416,N_1359);
xnor U5996 (N_5996,N_501,N_2450);
nand U5997 (N_5997,N_1948,N_733);
xor U5998 (N_5998,N_2663,N_190);
or U5999 (N_5999,N_681,N_1625);
or U6000 (N_6000,N_5525,N_5388);
nand U6001 (N_6001,N_5673,N_4303);
nor U6002 (N_6002,N_5489,N_3616);
and U6003 (N_6003,N_5804,N_5888);
or U6004 (N_6004,N_4444,N_4557);
nand U6005 (N_6005,N_3056,N_5212);
and U6006 (N_6006,N_4091,N_5091);
nor U6007 (N_6007,N_5275,N_4970);
or U6008 (N_6008,N_4057,N_4314);
and U6009 (N_6009,N_3910,N_4025);
and U6010 (N_6010,N_4428,N_3707);
xor U6011 (N_6011,N_4002,N_5995);
nor U6012 (N_6012,N_4814,N_4561);
nand U6013 (N_6013,N_5485,N_4518);
and U6014 (N_6014,N_5934,N_3730);
nor U6015 (N_6015,N_3259,N_3870);
or U6016 (N_6016,N_5653,N_5740);
nand U6017 (N_6017,N_4865,N_3545);
nor U6018 (N_6018,N_4842,N_5831);
nor U6019 (N_6019,N_4938,N_4829);
xnor U6020 (N_6020,N_5389,N_5067);
or U6021 (N_6021,N_5768,N_3580);
or U6022 (N_6022,N_5955,N_3725);
xor U6023 (N_6023,N_5199,N_4045);
and U6024 (N_6024,N_5614,N_5724);
and U6025 (N_6025,N_4902,N_4704);
nor U6026 (N_6026,N_3272,N_5780);
and U6027 (N_6027,N_4188,N_4388);
or U6028 (N_6028,N_5984,N_3785);
nor U6029 (N_6029,N_3524,N_4223);
nand U6030 (N_6030,N_3138,N_4221);
or U6031 (N_6031,N_4526,N_3869);
nand U6032 (N_6032,N_5432,N_3495);
xor U6033 (N_6033,N_4151,N_4701);
or U6034 (N_6034,N_4610,N_5259);
nor U6035 (N_6035,N_3302,N_3890);
xor U6036 (N_6036,N_3742,N_5428);
or U6037 (N_6037,N_4978,N_4370);
and U6038 (N_6038,N_4772,N_5070);
xor U6039 (N_6039,N_4852,N_4476);
and U6040 (N_6040,N_5945,N_5017);
nand U6041 (N_6041,N_4949,N_5741);
nand U6042 (N_6042,N_5878,N_3084);
and U6043 (N_6043,N_5403,N_5548);
or U6044 (N_6044,N_5564,N_5876);
and U6045 (N_6045,N_5985,N_5441);
or U6046 (N_6046,N_5932,N_4964);
nor U6047 (N_6047,N_4300,N_4523);
xor U6048 (N_6048,N_4257,N_5265);
nand U6049 (N_6049,N_4510,N_4318);
and U6050 (N_6050,N_4966,N_4089);
or U6051 (N_6051,N_4888,N_4307);
and U6052 (N_6052,N_3195,N_3666);
or U6053 (N_6053,N_3090,N_5881);
or U6054 (N_6054,N_3876,N_4098);
or U6055 (N_6055,N_3823,N_3796);
or U6056 (N_6056,N_4622,N_5197);
or U6057 (N_6057,N_5574,N_4912);
xnor U6058 (N_6058,N_5851,N_5782);
or U6059 (N_6059,N_3954,N_5603);
xor U6060 (N_6060,N_3689,N_5762);
xor U6061 (N_6061,N_3368,N_3743);
nand U6062 (N_6062,N_3546,N_5620);
xor U6063 (N_6063,N_4359,N_4077);
nand U6064 (N_6064,N_3511,N_4786);
nand U6065 (N_6065,N_5993,N_4178);
or U6066 (N_6066,N_3288,N_4943);
nor U6067 (N_6067,N_4216,N_3875);
xnor U6068 (N_6068,N_4122,N_3203);
and U6069 (N_6069,N_4236,N_3585);
or U6070 (N_6070,N_4560,N_3759);
and U6071 (N_6071,N_4874,N_4352);
or U6072 (N_6072,N_3283,N_4791);
xnor U6073 (N_6073,N_3590,N_4075);
nor U6074 (N_6074,N_3162,N_4164);
and U6075 (N_6075,N_4000,N_4773);
and U6076 (N_6076,N_4714,N_4958);
nand U6077 (N_6077,N_5186,N_4722);
nor U6078 (N_6078,N_5447,N_3924);
or U6079 (N_6079,N_5010,N_5412);
and U6080 (N_6080,N_3083,N_3281);
and U6081 (N_6081,N_5665,N_4816);
or U6082 (N_6082,N_5555,N_5503);
nand U6083 (N_6083,N_3547,N_5511);
nand U6084 (N_6084,N_5474,N_3502);
or U6085 (N_6085,N_5990,N_5766);
or U6086 (N_6086,N_5090,N_3168);
nor U6087 (N_6087,N_3454,N_4652);
nor U6088 (N_6088,N_5732,N_5788);
nor U6089 (N_6089,N_5068,N_5772);
nand U6090 (N_6090,N_3335,N_3817);
nand U6091 (N_6091,N_3134,N_4372);
xor U6092 (N_6092,N_4778,N_5889);
nand U6093 (N_6093,N_5746,N_4932);
nand U6094 (N_6094,N_4528,N_3466);
xnor U6095 (N_6095,N_4607,N_5882);
or U6096 (N_6096,N_5280,N_3717);
nand U6097 (N_6097,N_3223,N_4042);
or U6098 (N_6098,N_3777,N_3933);
and U6099 (N_6099,N_5373,N_3212);
and U6100 (N_6100,N_5506,N_4500);
and U6101 (N_6101,N_5334,N_3993);
and U6102 (N_6102,N_5736,N_4290);
xor U6103 (N_6103,N_3934,N_3755);
or U6104 (N_6104,N_3520,N_4915);
xor U6105 (N_6105,N_3818,N_5970);
or U6106 (N_6106,N_3367,N_3053);
and U6107 (N_6107,N_4577,N_5825);
nor U6108 (N_6108,N_4394,N_3529);
xor U6109 (N_6109,N_4491,N_4564);
and U6110 (N_6110,N_4276,N_3155);
or U6111 (N_6111,N_3481,N_5187);
xnor U6112 (N_6112,N_4161,N_3437);
or U6113 (N_6113,N_3709,N_5534);
nor U6114 (N_6114,N_5348,N_5697);
or U6115 (N_6115,N_5361,N_4945);
or U6116 (N_6116,N_4447,N_3381);
nand U6117 (N_6117,N_3112,N_4203);
xor U6118 (N_6118,N_5180,N_5501);
and U6119 (N_6119,N_5700,N_5211);
nor U6120 (N_6120,N_3323,N_4123);
xor U6121 (N_6121,N_3810,N_5947);
or U6122 (N_6122,N_5537,N_3800);
nand U6123 (N_6123,N_4777,N_4142);
xnor U6124 (N_6124,N_3308,N_5434);
and U6125 (N_6125,N_5834,N_5602);
xnor U6126 (N_6126,N_5758,N_5685);
or U6127 (N_6127,N_4097,N_4039);
and U6128 (N_6128,N_3807,N_3263);
or U6129 (N_6129,N_3643,N_3158);
nand U6130 (N_6130,N_5647,N_5591);
nor U6131 (N_6131,N_3157,N_3034);
xor U6132 (N_6132,N_3932,N_5482);
nand U6133 (N_6133,N_4726,N_3496);
and U6134 (N_6134,N_3067,N_5917);
or U6135 (N_6135,N_5638,N_3718);
and U6136 (N_6136,N_5101,N_4190);
nor U6137 (N_6137,N_5797,N_3955);
xnor U6138 (N_6138,N_5705,N_5290);
nand U6139 (N_6139,N_3864,N_5808);
nor U6140 (N_6140,N_3037,N_5026);
xnor U6141 (N_6141,N_5805,N_4730);
nor U6142 (N_6142,N_5706,N_3284);
or U6143 (N_6143,N_4118,N_4272);
or U6144 (N_6144,N_4116,N_4141);
nor U6145 (N_6145,N_4803,N_4304);
and U6146 (N_6146,N_3901,N_4661);
or U6147 (N_6147,N_5337,N_4796);
nand U6148 (N_6148,N_3975,N_4611);
or U6149 (N_6149,N_3136,N_4343);
nor U6150 (N_6150,N_3413,N_5580);
nor U6151 (N_6151,N_3277,N_4189);
nand U6152 (N_6152,N_3710,N_4544);
xor U6153 (N_6153,N_5451,N_3541);
nor U6154 (N_6154,N_4595,N_3645);
nand U6155 (N_6155,N_4844,N_4267);
nand U6156 (N_6156,N_5387,N_4815);
or U6157 (N_6157,N_5627,N_4270);
and U6158 (N_6158,N_4515,N_5530);
xor U6159 (N_6159,N_5579,N_4612);
or U6160 (N_6160,N_3235,N_5321);
nor U6161 (N_6161,N_4843,N_3172);
nor U6162 (N_6162,N_4132,N_4674);
nand U6163 (N_6163,N_5146,N_5927);
and U6164 (N_6164,N_4056,N_3861);
xor U6165 (N_6165,N_5483,N_5452);
xnor U6166 (N_6166,N_3724,N_4527);
and U6167 (N_6167,N_3105,N_5427);
or U6168 (N_6168,N_5058,N_4997);
nor U6169 (N_6169,N_5196,N_4185);
nand U6170 (N_6170,N_3074,N_5000);
and U6171 (N_6171,N_3720,N_4402);
nand U6172 (N_6172,N_4727,N_3018);
nand U6173 (N_6173,N_3706,N_3399);
or U6174 (N_6174,N_3300,N_5301);
xnor U6175 (N_6175,N_5975,N_5004);
nor U6176 (N_6176,N_4382,N_3179);
nor U6177 (N_6177,N_4933,N_5251);
or U6178 (N_6178,N_5898,N_5274);
xor U6179 (N_6179,N_4846,N_5689);
and U6180 (N_6180,N_5130,N_4639);
xnor U6181 (N_6181,N_3280,N_4348);
nor U6182 (N_6182,N_5380,N_4043);
nor U6183 (N_6183,N_3160,N_3116);
and U6184 (N_6184,N_3394,N_4569);
xor U6185 (N_6185,N_5332,N_3668);
and U6186 (N_6186,N_4451,N_5553);
xor U6187 (N_6187,N_3363,N_3349);
nor U6188 (N_6188,N_5462,N_5966);
xnor U6189 (N_6189,N_3998,N_5405);
nand U6190 (N_6190,N_3415,N_5264);
or U6191 (N_6191,N_5271,N_5129);
nand U6192 (N_6192,N_5919,N_4017);
and U6193 (N_6193,N_5473,N_3544);
nor U6194 (N_6194,N_5976,N_3703);
xnor U6195 (N_6195,N_5436,N_4710);
xnor U6196 (N_6196,N_4209,N_5406);
nor U6197 (N_6197,N_3698,N_5909);
or U6198 (N_6198,N_5939,N_4277);
or U6199 (N_6199,N_4385,N_4358);
and U6200 (N_6200,N_3749,N_3611);
and U6201 (N_6201,N_3214,N_4899);
xnor U6202 (N_6202,N_3863,N_3741);
or U6203 (N_6203,N_4512,N_4897);
xnor U6204 (N_6204,N_4921,N_5841);
nand U6205 (N_6205,N_4060,N_4242);
nor U6206 (N_6206,N_3566,N_4884);
nand U6207 (N_6207,N_4636,N_3103);
and U6208 (N_6208,N_5637,N_3151);
and U6209 (N_6209,N_3485,N_4241);
nand U6210 (N_6210,N_3120,N_4825);
nand U6211 (N_6211,N_3561,N_3336);
and U6212 (N_6212,N_4081,N_5254);
xnor U6213 (N_6213,N_5079,N_4963);
or U6214 (N_6214,N_5830,N_3574);
xor U6215 (N_6215,N_5366,N_5495);
or U6216 (N_6216,N_4826,N_5941);
or U6217 (N_6217,N_4302,N_4919);
xnor U6218 (N_6218,N_4881,N_4731);
and U6219 (N_6219,N_4634,N_3608);
xor U6220 (N_6220,N_4836,N_4227);
nor U6221 (N_6221,N_4166,N_3442);
nor U6222 (N_6222,N_5069,N_5832);
or U6223 (N_6223,N_3327,N_3145);
xor U6224 (N_6224,N_4054,N_4996);
and U6225 (N_6225,N_4766,N_5690);
or U6226 (N_6226,N_5549,N_3745);
and U6227 (N_6227,N_3441,N_4479);
nand U6228 (N_6228,N_4432,N_3497);
nand U6229 (N_6229,N_3445,N_3313);
or U6230 (N_6230,N_5873,N_4985);
nand U6231 (N_6231,N_3530,N_3218);
xor U6232 (N_6232,N_3129,N_4441);
nand U6233 (N_6233,N_5370,N_5105);
and U6234 (N_6234,N_5583,N_5551);
and U6235 (N_6235,N_5817,N_3588);
and U6236 (N_6236,N_4086,N_3695);
or U6237 (N_6237,N_4935,N_3683);
xor U6238 (N_6238,N_5519,N_3965);
xor U6239 (N_6239,N_5184,N_4617);
xor U6240 (N_6240,N_3356,N_3141);
or U6241 (N_6241,N_3477,N_3029);
nand U6242 (N_6242,N_4923,N_5250);
nor U6243 (N_6243,N_4589,N_3872);
and U6244 (N_6244,N_4708,N_4376);
and U6245 (N_6245,N_5520,N_3728);
nor U6246 (N_6246,N_3686,N_4279);
nand U6247 (N_6247,N_5731,N_4551);
nor U6248 (N_6248,N_5677,N_4538);
nand U6249 (N_6249,N_5468,N_5409);
nand U6250 (N_6250,N_5982,N_3781);
nor U6251 (N_6251,N_4632,N_5465);
and U6252 (N_6252,N_4941,N_5936);
or U6253 (N_6253,N_4619,N_3811);
and U6254 (N_6254,N_4357,N_4981);
nor U6255 (N_6255,N_3512,N_3312);
and U6256 (N_6256,N_5131,N_5860);
and U6257 (N_6257,N_4156,N_4378);
and U6258 (N_6258,N_5981,N_5987);
or U6259 (N_6259,N_3365,N_5112);
nand U6260 (N_6260,N_3884,N_3310);
xnor U6261 (N_6261,N_4239,N_5718);
nor U6262 (N_6262,N_4130,N_5542);
xor U6263 (N_6263,N_3265,N_5439);
xnor U6264 (N_6264,N_4524,N_3767);
nor U6265 (N_6265,N_3221,N_3828);
or U6266 (N_6266,N_5656,N_4102);
nor U6267 (N_6267,N_4988,N_4109);
xor U6268 (N_6268,N_3422,N_4396);
nand U6269 (N_6269,N_3137,N_5011);
xor U6270 (N_6270,N_5419,N_3022);
nand U6271 (N_6271,N_5381,N_5815);
nor U6272 (N_6272,N_3531,N_4680);
nor U6273 (N_6273,N_4289,N_3476);
or U6274 (N_6274,N_3079,N_4615);
nor U6275 (N_6275,N_3516,N_3017);
nand U6276 (N_6276,N_3681,N_5566);
xor U6277 (N_6277,N_5526,N_3460);
nand U6278 (N_6278,N_5569,N_5233);
nand U6279 (N_6279,N_3052,N_3009);
or U6280 (N_6280,N_5471,N_5613);
and U6281 (N_6281,N_4858,N_5231);
and U6282 (N_6282,N_3921,N_4474);
nor U6283 (N_6283,N_5765,N_3847);
nand U6284 (N_6284,N_3325,N_4651);
nor U6285 (N_6285,N_5365,N_4608);
nand U6286 (N_6286,N_5127,N_4404);
nand U6287 (N_6287,N_4115,N_5488);
or U6288 (N_6288,N_5426,N_3661);
or U6289 (N_6289,N_3233,N_4516);
xor U6290 (N_6290,N_5385,N_4292);
and U6291 (N_6291,N_3478,N_4658);
xor U6292 (N_6292,N_5002,N_4295);
or U6293 (N_6293,N_3679,N_3920);
and U6294 (N_6294,N_5901,N_5260);
or U6295 (N_6295,N_3963,N_5824);
xnor U6296 (N_6296,N_3417,N_5783);
nand U6297 (N_6297,N_4495,N_3007);
nor U6298 (N_6298,N_4138,N_4575);
nand U6299 (N_6299,N_5034,N_4698);
or U6300 (N_6300,N_3628,N_4763);
nand U6301 (N_6301,N_5124,N_3500);
nor U6302 (N_6302,N_5375,N_3459);
or U6303 (N_6303,N_5437,N_4268);
xor U6304 (N_6304,N_4266,N_4519);
nand U6305 (N_6305,N_5601,N_5498);
xor U6306 (N_6306,N_5449,N_3040);
nor U6307 (N_6307,N_3788,N_3046);
or U6308 (N_6308,N_3935,N_3789);
and U6309 (N_6309,N_4793,N_5796);
or U6310 (N_6310,N_3328,N_5794);
nand U6311 (N_6311,N_3114,N_5065);
or U6312 (N_6312,N_4992,N_3946);
and U6313 (N_6313,N_3860,N_4746);
and U6314 (N_6314,N_3945,N_4546);
and U6315 (N_6315,N_3069,N_5650);
or U6316 (N_6316,N_3187,N_4646);
nand U6317 (N_6317,N_4271,N_3489);
nor U6318 (N_6318,N_5237,N_3694);
or U6319 (N_6319,N_4940,N_4226);
and U6320 (N_6320,N_5351,N_4321);
nand U6321 (N_6321,N_4602,N_5561);
nor U6322 (N_6322,N_4720,N_4979);
nand U6323 (N_6323,N_3771,N_3806);
nand U6324 (N_6324,N_5216,N_5054);
and U6325 (N_6325,N_3450,N_4275);
or U6326 (N_6326,N_4715,N_4711);
and U6327 (N_6327,N_4063,N_4194);
nor U6328 (N_6328,N_5390,N_4851);
or U6329 (N_6329,N_3982,N_3347);
or U6330 (N_6330,N_4336,N_3224);
xnor U6331 (N_6331,N_5720,N_5223);
xnor U6332 (N_6332,N_5175,N_4489);
and U6333 (N_6333,N_4106,N_3840);
xnor U6334 (N_6334,N_4211,N_4001);
and U6335 (N_6335,N_4162,N_5745);
and U6336 (N_6336,N_3101,N_5019);
nand U6337 (N_6337,N_5914,N_3229);
nor U6338 (N_6338,N_4670,N_4145);
nor U6339 (N_6339,N_4008,N_5377);
or U6340 (N_6340,N_3086,N_4215);
xor U6341 (N_6341,N_3438,N_5368);
xor U6342 (N_6342,N_5203,N_4663);
xnor U6343 (N_6343,N_4584,N_5022);
nor U6344 (N_6344,N_3358,N_4010);
and U6345 (N_6345,N_3464,N_5560);
or U6346 (N_6346,N_4628,N_3410);
and U6347 (N_6347,N_4513,N_4464);
xor U6348 (N_6348,N_5973,N_4984);
and U6349 (N_6349,N_5836,N_4395);
or U6350 (N_6350,N_5826,N_5494);
or U6351 (N_6351,N_5543,N_4709);
xor U6352 (N_6352,N_4414,N_5342);
or U6353 (N_6353,N_4568,N_3401);
xnor U6354 (N_6354,N_4386,N_5969);
nand U6355 (N_6355,N_3050,N_3264);
nand U6356 (N_6356,N_4049,N_4532);
nor U6357 (N_6357,N_3360,N_3593);
and U6358 (N_6358,N_3534,N_3239);
and U6359 (N_6359,N_3513,N_3904);
and U6360 (N_6360,N_3238,N_5930);
xnor U6361 (N_6361,N_3715,N_4136);
and U6362 (N_6362,N_4790,N_4427);
xor U6363 (N_6363,N_5194,N_3342);
or U6364 (N_6364,N_5717,N_3487);
xnor U6365 (N_6365,N_5658,N_3652);
nor U6366 (N_6366,N_5801,N_4547);
nand U6367 (N_6367,N_4693,N_5557);
nor U6368 (N_6368,N_3631,N_3411);
nor U6369 (N_6369,N_5722,N_5554);
nor U6370 (N_6370,N_4436,N_4186);
or U6371 (N_6371,N_5989,N_3304);
or U6372 (N_6372,N_4251,N_4671);
or U6373 (N_6373,N_3483,N_4768);
nor U6374 (N_6374,N_5209,N_3968);
nand U6375 (N_6375,N_5958,N_5476);
and U6376 (N_6376,N_4411,N_5983);
or U6377 (N_6377,N_4809,N_4878);
or U6378 (N_6378,N_5350,N_3020);
nor U6379 (N_6379,N_3311,N_5335);
or U6380 (N_6380,N_3783,N_3254);
nand U6381 (N_6381,N_3468,N_4204);
xnor U6382 (N_6382,N_5719,N_4662);
nand U6383 (N_6383,N_3688,N_4019);
and U6384 (N_6384,N_3038,N_4805);
nor U6385 (N_6385,N_5311,N_5053);
xor U6386 (N_6386,N_4509,N_4015);
xor U6387 (N_6387,N_3372,N_4853);
nand U6388 (N_6388,N_3929,N_4975);
nor U6389 (N_6389,N_4305,N_5528);
and U6390 (N_6390,N_3440,N_4762);
nor U6391 (N_6391,N_5208,N_3196);
or U6392 (N_6392,N_3232,N_3307);
or U6393 (N_6393,N_3913,N_4688);
nand U6394 (N_6394,N_3927,N_5813);
xor U6395 (N_6395,N_5967,N_3309);
xnor U6396 (N_6396,N_4410,N_5659);
xnor U6397 (N_6397,N_3882,N_5800);
or U6398 (N_6398,N_4250,N_4535);
or U6399 (N_6399,N_5964,N_3491);
nor U6400 (N_6400,N_3230,N_3554);
xnor U6401 (N_6401,N_5082,N_4496);
xnor U6402 (N_6402,N_3331,N_4167);
nand U6403 (N_6403,N_3149,N_3226);
or U6404 (N_6404,N_5305,N_5059);
or U6405 (N_6405,N_4265,N_3937);
nand U6406 (N_6406,N_3031,N_5571);
nand U6407 (N_6407,N_3607,N_4700);
and U6408 (N_6408,N_3292,N_4244);
nand U6409 (N_6409,N_5657,N_4240);
nand U6410 (N_6410,N_3990,N_4176);
or U6411 (N_6411,N_4459,N_5663);
and U6412 (N_6412,N_4064,N_4398);
nand U6413 (N_6413,N_4213,N_5077);
and U6414 (N_6414,N_3987,N_3190);
or U6415 (N_6415,N_5630,N_4012);
xor U6416 (N_6416,N_5809,N_4706);
xnor U6417 (N_6417,N_4920,N_4055);
xor U6418 (N_6418,N_3687,N_4332);
nor U6419 (N_6419,N_4287,N_5852);
xnor U6420 (N_6420,N_4906,N_4264);
or U6421 (N_6421,N_5573,N_5297);
xnor U6422 (N_6422,N_4732,N_3775);
and U6423 (N_6423,N_3154,N_4383);
nor U6424 (N_6424,N_5870,N_5003);
nor U6425 (N_6425,N_3470,N_3075);
nor U6426 (N_6426,N_3064,N_4859);
nand U6427 (N_6427,N_4177,N_5725);
nand U6428 (N_6428,N_3750,N_3274);
nand U6429 (N_6429,N_5159,N_4999);
nand U6430 (N_6430,N_5032,N_3797);
or U6431 (N_6431,N_3886,N_4249);
nand U6432 (N_6432,N_3769,N_4795);
or U6433 (N_6433,N_4890,N_4534);
and U6434 (N_6434,N_4096,N_4417);
nand U6435 (N_6435,N_4296,N_4455);
xor U6436 (N_6436,N_4928,N_4195);
and U6437 (N_6437,N_3727,N_5675);
nand U6438 (N_6438,N_5522,N_3174);
nand U6439 (N_6439,N_5959,N_5430);
xnor U6440 (N_6440,N_4092,N_3278);
nand U6441 (N_6441,N_4672,N_5227);
nor U6442 (N_6442,N_5621,N_3831);
xor U6443 (N_6443,N_5323,N_3205);
nand U6444 (N_6444,N_5532,N_4744);
or U6445 (N_6445,N_3739,N_3418);
nand U6446 (N_6446,N_3733,N_5752);
or U6447 (N_6447,N_4253,N_5048);
xnor U6448 (N_6448,N_4368,N_3200);
nand U6449 (N_6449,N_4013,N_4574);
and U6450 (N_6450,N_5942,N_3508);
nand U6451 (N_6451,N_3598,N_4152);
or U6452 (N_6452,N_5152,N_4004);
xor U6453 (N_6453,N_5183,N_3093);
or U6454 (N_6454,N_3255,N_5153);
and U6455 (N_6455,N_3337,N_3883);
or U6456 (N_6456,N_5714,N_4445);
or U6457 (N_6457,N_3473,N_3412);
xnor U6458 (N_6458,N_5221,N_4369);
or U6459 (N_6459,N_4736,N_3964);
and U6460 (N_6460,N_3858,N_5651);
nor U6461 (N_6461,N_5905,N_5908);
or U6462 (N_6462,N_5325,N_3291);
nand U6463 (N_6463,N_4419,N_4586);
xor U6464 (N_6464,N_5167,N_4643);
and U6465 (N_6465,N_4477,N_3603);
nand U6466 (N_6466,N_3856,N_3655);
or U6467 (N_6467,N_5492,N_4182);
nand U6468 (N_6468,N_4614,N_4552);
xor U6469 (N_6469,N_4649,N_5938);
xnor U6470 (N_6470,N_3953,N_4678);
nand U6471 (N_6471,N_4283,N_4620);
nor U6472 (N_6472,N_4655,N_3294);
and U6473 (N_6473,N_4280,N_5455);
or U6474 (N_6474,N_5458,N_3943);
nor U6475 (N_6475,N_5885,N_3549);
xor U6476 (N_6476,N_4642,N_5163);
xnor U6477 (N_6477,N_4175,N_3197);
xor U6478 (N_6478,N_5352,N_3532);
xor U6479 (N_6479,N_4488,N_3322);
nand U6480 (N_6480,N_5541,N_4924);
xnor U6481 (N_6481,N_4522,N_3731);
or U6482 (N_6482,N_5143,N_4724);
nor U6483 (N_6483,N_5100,N_3537);
or U6484 (N_6484,N_5702,N_4345);
nor U6485 (N_6485,N_4007,N_4601);
nor U6486 (N_6486,N_3439,N_4752);
and U6487 (N_6487,N_5968,N_4199);
and U6488 (N_6488,N_3618,N_3726);
nand U6489 (N_6489,N_4898,N_5978);
nand U6490 (N_6490,N_3428,N_4059);
nand U6491 (N_6491,N_3177,N_3117);
and U6492 (N_6492,N_3124,N_4549);
nor U6493 (N_6493,N_5998,N_5247);
nand U6494 (N_6494,N_4960,N_4016);
or U6495 (N_6495,N_4862,N_3714);
nor U6496 (N_6496,N_4517,N_5679);
nand U6497 (N_6497,N_4033,N_5716);
or U6498 (N_6498,N_4324,N_5915);
or U6499 (N_6499,N_4037,N_4695);
and U6500 (N_6500,N_3515,N_5150);
xor U6501 (N_6501,N_4764,N_4035);
nor U6502 (N_6502,N_5811,N_3748);
or U6503 (N_6503,N_5097,N_3094);
nor U6504 (N_6504,N_5001,N_5040);
xor U6505 (N_6505,N_5461,N_5469);
nor U6506 (N_6506,N_4624,N_4430);
or U6507 (N_6507,N_5454,N_4469);
xnor U6508 (N_6508,N_5819,N_3676);
or U6509 (N_6509,N_3822,N_5868);
and U6510 (N_6510,N_3630,N_5193);
xnor U6511 (N_6511,N_4355,N_4487);
and U6512 (N_6512,N_5661,N_4962);
nor U6513 (N_6513,N_3005,N_5165);
or U6514 (N_6514,N_4687,N_5974);
xor U6515 (N_6515,N_4212,N_4857);
and U6516 (N_6516,N_3579,N_5980);
nor U6517 (N_6517,N_3868,N_3245);
nor U6518 (N_6518,N_3370,N_3306);
and U6519 (N_6519,N_4463,N_3297);
or U6520 (N_6520,N_4514,N_5098);
nor U6521 (N_6521,N_4458,N_4679);
and U6522 (N_6522,N_3721,N_5246);
xor U6523 (N_6523,N_4375,N_3885);
xnor U6524 (N_6524,N_5397,N_4117);
and U6525 (N_6525,N_3150,N_4645);
or U6526 (N_6526,N_3564,N_3183);
or U6527 (N_6527,N_4003,N_5750);
nor U6528 (N_6528,N_3405,N_5562);
nand U6529 (N_6529,N_3165,N_4067);
nor U6530 (N_6530,N_3402,N_5570);
or U6531 (N_6531,N_3251,N_4446);
xnor U6532 (N_6532,N_3452,N_3036);
nor U6533 (N_6533,N_4471,N_5916);
or U6534 (N_6534,N_5148,N_3219);
or U6535 (N_6535,N_5273,N_4539);
xnor U6536 (N_6536,N_3557,N_3670);
or U6537 (N_6537,N_3950,N_4238);
and U6538 (N_6538,N_3374,N_5926);
nor U6539 (N_6539,N_4756,N_5546);
or U6540 (N_6540,N_4505,N_3045);
or U6541 (N_6541,N_5345,N_4408);
xor U6542 (N_6542,N_4580,N_3471);
xnor U6543 (N_6543,N_5844,N_5676);
or U6544 (N_6544,N_3791,N_4237);
or U6545 (N_6545,N_3248,N_5126);
nor U6546 (N_6546,N_3048,N_5464);
xor U6547 (N_6547,N_5715,N_5249);
and U6548 (N_6548,N_3166,N_4637);
or U6549 (N_6549,N_4088,N_4641);
nand U6550 (N_6550,N_3184,N_4429);
xor U6551 (N_6551,N_5491,N_3770);
or U6552 (N_6552,N_4090,N_4282);
nand U6553 (N_6553,N_5684,N_5453);
or U6554 (N_6554,N_4099,N_3560);
nor U6555 (N_6555,N_4206,N_3217);
xnor U6556 (N_6556,N_4163,N_5877);
or U6557 (N_6557,N_5539,N_4987);
and U6558 (N_6558,N_3572,N_5833);
nand U6559 (N_6559,N_5948,N_5935);
xnor U6560 (N_6560,N_4165,N_3296);
nand U6561 (N_6561,N_5372,N_3510);
nor U6562 (N_6562,N_4644,N_3974);
xor U6563 (N_6563,N_4074,N_5244);
and U6564 (N_6564,N_5156,N_5303);
nor U6565 (N_6565,N_3133,N_3474);
nor U6566 (N_6566,N_3766,N_5642);
xor U6567 (N_6567,N_5652,N_4755);
nor U6568 (N_6568,N_5006,N_5042);
or U6569 (N_6569,N_5701,N_3448);
nor U6570 (N_6570,N_3614,N_5671);
xor U6571 (N_6571,N_5754,N_4837);
or U6572 (N_6572,N_5828,N_4931);
or U6573 (N_6573,N_4880,N_5735);
nor U6574 (N_6574,N_3109,N_3866);
and U6575 (N_6575,N_5139,N_3078);
xnor U6576 (N_6576,N_4692,N_5241);
nor U6577 (N_6577,N_4113,N_4944);
nor U6578 (N_6578,N_3629,N_5504);
nor U6579 (N_6579,N_3436,N_3527);
nand U6580 (N_6580,N_4588,N_3625);
or U6581 (N_6581,N_3106,N_5738);
or U6582 (N_6582,N_4686,N_3260);
and U6583 (N_6583,N_4330,N_5703);
xnor U6584 (N_6584,N_4076,N_4320);
xor U6585 (N_6585,N_5837,N_4848);
and U6586 (N_6586,N_4694,N_3210);
and U6587 (N_6587,N_4579,N_3916);
xor U6588 (N_6588,N_3125,N_5587);
nand U6589 (N_6589,N_5151,N_4625);
nor U6590 (N_6590,N_5119,N_3073);
nand U6591 (N_6591,N_5288,N_4407);
or U6592 (N_6592,N_4058,N_5394);
or U6593 (N_6593,N_4301,N_3361);
or U6594 (N_6594,N_4835,N_3049);
nor U6595 (N_6595,N_5178,N_5088);
or U6596 (N_6596,N_4864,N_4571);
nor U6597 (N_6597,N_5189,N_5463);
xnor U6598 (N_6598,N_4111,N_4900);
and U6599 (N_6599,N_4405,N_5857);
and U6600 (N_6600,N_3862,N_5787);
xor U6601 (N_6601,N_4952,N_4503);
and U6602 (N_6602,N_3877,N_5295);
and U6603 (N_6603,N_3812,N_5814);
nor U6604 (N_6604,N_3406,N_4834);
nand U6605 (N_6605,N_5071,N_3793);
and U6606 (N_6606,N_5517,N_5018);
and U6607 (N_6607,N_4110,N_5440);
or U6608 (N_6608,N_4465,N_5681);
or U6609 (N_6609,N_3584,N_5438);
and U6610 (N_6610,N_3568,N_5318);
xnor U6611 (N_6611,N_4681,N_4737);
xor U6612 (N_6612,N_4585,N_3303);
nor U6613 (N_6613,N_4124,N_3228);
nand U6614 (N_6614,N_3784,N_4220);
and U6615 (N_6615,N_5523,N_4139);
nand U6616 (N_6616,N_5362,N_3169);
or U6617 (N_6617,N_4424,N_5820);
nor U6618 (N_6618,N_3305,N_3553);
xnor U6619 (N_6619,N_4434,N_4506);
or U6620 (N_6620,N_5266,N_5029);
and U6621 (N_6621,N_5739,N_4903);
and U6622 (N_6622,N_4550,N_3012);
or U6623 (N_6623,N_4160,N_3054);
nor U6624 (N_6624,N_3708,N_3222);
nand U6625 (N_6625,N_5737,N_5417);
nor U6626 (N_6626,N_4093,N_3175);
or U6627 (N_6627,N_4146,N_5309);
nor U6628 (N_6628,N_3243,N_3737);
xor U6629 (N_6629,N_4684,N_4719);
and U6630 (N_6630,N_5236,N_4072);
xor U6631 (N_6631,N_3981,N_5484);
nand U6632 (N_6632,N_4869,N_3888);
or U6633 (N_6633,N_3493,N_5294);
nor U6634 (N_6634,N_4929,N_5626);
nor U6635 (N_6635,N_4667,N_4377);
and U6636 (N_6636,N_5478,N_4761);
or U6637 (N_6637,N_5316,N_4169);
or U6638 (N_6638,N_3507,N_4930);
nor U6639 (N_6639,N_5624,N_4020);
nor U6640 (N_6640,N_4274,N_3633);
and U6641 (N_6641,N_4543,N_5645);
and U6642 (N_6642,N_4245,N_5308);
nor U6643 (N_6643,N_3925,N_3484);
xnor U6644 (N_6644,N_4827,N_3700);
nor U6645 (N_6645,N_5393,N_5662);
nand U6646 (N_6646,N_3632,N_3390);
xor U6647 (N_6647,N_5374,N_4050);
nand U6648 (N_6648,N_4802,N_4840);
nand U6649 (N_6649,N_5166,N_4380);
or U6650 (N_6650,N_3189,N_5664);
or U6651 (N_6651,N_4740,N_4769);
nor U6652 (N_6652,N_4590,N_4626);
xnor U6653 (N_6653,N_3562,N_3619);
xor U6654 (N_6654,N_3426,N_3835);
or U6655 (N_6655,N_5014,N_5141);
nor U6656 (N_6656,N_5578,N_4507);
and U6657 (N_6657,N_5314,N_4078);
and U6658 (N_6658,N_4953,N_3573);
and U6659 (N_6659,N_5344,N_3702);
nand U6660 (N_6660,N_4183,N_5655);
or U6661 (N_6661,N_3634,N_4340);
nor U6662 (N_6662,N_3364,N_4501);
and U6663 (N_6663,N_5043,N_5565);
and U6664 (N_6664,N_3772,N_4593);
nor U6665 (N_6665,N_4627,N_4754);
xor U6666 (N_6666,N_3680,N_5891);
and U6667 (N_6667,N_4027,N_4051);
and U6668 (N_6668,N_5516,N_5396);
and U6669 (N_6669,N_3991,N_5606);
nor U6670 (N_6670,N_3723,N_5232);
nand U6671 (N_6671,N_4748,N_5358);
and U6672 (N_6672,N_3786,N_5899);
and U6673 (N_6673,N_4219,N_3782);
nor U6674 (N_6674,N_3732,N_4936);
and U6675 (N_6675,N_4563,N_4046);
or U6676 (N_6676,N_5267,N_3080);
or U6677 (N_6677,N_5890,N_4937);
and U6678 (N_6678,N_5508,N_4170);
or U6679 (N_6679,N_3995,N_3578);
and U6680 (N_6680,N_4134,N_4107);
nand U6681 (N_6681,N_5329,N_3764);
nand U6682 (N_6682,N_5729,N_5683);
xnor U6683 (N_6683,N_5252,N_3826);
nand U6684 (N_6684,N_5424,N_3622);
nand U6685 (N_6685,N_5225,N_3701);
xor U6686 (N_6686,N_5604,N_4397);
nand U6687 (N_6687,N_3693,N_3768);
nor U6688 (N_6688,N_5005,N_3602);
nor U6689 (N_6689,N_5333,N_4202);
xnor U6690 (N_6690,N_3960,N_4466);
nor U6691 (N_6691,N_5568,N_4572);
xnor U6692 (N_6692,N_5979,N_5111);
xor U6693 (N_6693,N_5445,N_4052);
nand U6694 (N_6694,N_5477,N_3346);
nand U6695 (N_6695,N_5790,N_5270);
xnor U6696 (N_6696,N_4365,N_3126);
and U6697 (N_6697,N_4418,N_3514);
and U6698 (N_6698,N_5922,N_5084);
and U6699 (N_6699,N_5545,N_4664);
xnor U6700 (N_6700,N_3601,N_3609);
or U6701 (N_6701,N_4082,N_3366);
nor U6702 (N_6702,N_3637,N_3032);
or U6703 (N_6703,N_5008,N_5763);
or U6704 (N_6704,N_3377,N_3359);
xnor U6705 (N_6705,N_4891,N_5289);
and U6706 (N_6706,N_5081,N_3928);
and U6707 (N_6707,N_5402,N_3908);
or U6708 (N_6708,N_5060,N_3833);
nor U6709 (N_6709,N_4860,N_3085);
xor U6710 (N_6710,N_5219,N_4750);
nand U6711 (N_6711,N_5558,N_4387);
nand U6712 (N_6712,N_5535,N_3463);
xor U6713 (N_6713,N_4886,N_4657);
and U6714 (N_6714,N_5928,N_4233);
and U6715 (N_6715,N_5640,N_3906);
nor U6716 (N_6716,N_4873,N_4968);
nand U6717 (N_6717,N_5253,N_3298);
xor U6718 (N_6718,N_4603,N_5929);
nor U6719 (N_6719,N_5698,N_4196);
nor U6720 (N_6720,N_4235,N_5442);
and U6721 (N_6721,N_4149,N_4894);
and U6722 (N_6722,N_5678,N_4855);
nor U6723 (N_6723,N_3857,N_4567);
and U6724 (N_6724,N_4606,N_4457);
nand U6725 (N_6725,N_5191,N_4482);
nand U6726 (N_6726,N_4946,N_4635);
and U6727 (N_6727,N_4497,N_3753);
xnor U6728 (N_6728,N_5369,N_5410);
or U6729 (N_6729,N_3236,N_5041);
and U6730 (N_6730,N_3178,N_4871);
or U6731 (N_6731,N_4473,N_3345);
and U6732 (N_6732,N_5164,N_4200);
xnor U6733 (N_6733,N_4977,N_5020);
and U6734 (N_6734,N_5622,N_3270);
and U6735 (N_6735,N_4733,N_4775);
and U6736 (N_6736,N_5238,N_4131);
xor U6737 (N_6737,N_3369,N_4225);
and U6738 (N_6738,N_3249,N_5505);
nand U6739 (N_6739,N_4461,N_4159);
and U6740 (N_6740,N_3446,N_3859);
or U6741 (N_6741,N_5798,N_5224);
xor U6742 (N_6742,N_4062,N_3589);
nor U6743 (N_6743,N_5075,N_3123);
xnor U6744 (N_6744,N_5343,N_3429);
nand U6745 (N_6745,N_5171,N_3986);
or U6746 (N_6746,N_4760,N_5281);
and U6747 (N_6747,N_5835,N_5472);
or U6748 (N_6748,N_3824,N_4011);
and U6749 (N_6749,N_3841,N_5298);
nor U6750 (N_6750,N_5147,N_5431);
nor U6751 (N_6751,N_3814,N_4023);
nor U6752 (N_6752,N_3639,N_4438);
or U6753 (N_6753,N_4148,N_4665);
nor U6754 (N_6754,N_5292,N_4363);
and U6755 (N_6755,N_4782,N_3836);
nor U6756 (N_6756,N_3834,N_4470);
or U6757 (N_6757,N_4591,N_5268);
or U6758 (N_6758,N_5756,N_5608);
or U6759 (N_6759,N_5330,N_3023);
and U6760 (N_6760,N_3128,N_3762);
nand U6761 (N_6761,N_5415,N_3059);
or U6762 (N_6762,N_4120,N_4353);
nand U6763 (N_6763,N_3518,N_3188);
and U6764 (N_6764,N_4576,N_4697);
xor U6765 (N_6765,N_4485,N_5354);
nor U6766 (N_6766,N_5154,N_3139);
and U6767 (N_6767,N_5030,N_3482);
and U6768 (N_6768,N_3674,N_4556);
nand U6769 (N_6769,N_3207,N_3690);
xnor U6770 (N_6770,N_4030,N_5986);
and U6771 (N_6771,N_5248,N_3605);
nor U6772 (N_6772,N_3389,N_5086);
nand U6773 (N_6773,N_3492,N_4403);
or U6774 (N_6774,N_4817,N_4808);
xor U6775 (N_6775,N_3504,N_3420);
nand U6776 (N_6776,N_4210,N_4454);
nand U6777 (N_6777,N_3842,N_4319);
xor U6778 (N_6778,N_3976,N_5202);
nor U6779 (N_6779,N_5304,N_3131);
nor U6780 (N_6780,N_4707,N_3761);
nand U6781 (N_6781,N_4094,N_4222);
and U6782 (N_6782,N_5028,N_5616);
and U6783 (N_6783,N_3543,N_5696);
xor U6784 (N_6784,N_5625,N_4431);
nand U6785 (N_6785,N_5629,N_5781);
and U6786 (N_6786,N_4258,N_3352);
and U6787 (N_6787,N_5121,N_4914);
nand U6788 (N_6788,N_5514,N_4327);
nand U6789 (N_6789,N_5952,N_5550);
xor U6790 (N_6790,N_3997,N_4558);
or U6791 (N_6791,N_5263,N_3211);
nor U6792 (N_6792,N_5687,N_5822);
nor U6793 (N_6793,N_4562,N_5423);
nand U6794 (N_6794,N_3181,N_3242);
xnor U6795 (N_6795,N_5138,N_3167);
nor U6796 (N_6796,N_5307,N_5161);
or U6797 (N_6797,N_4047,N_3849);
xnor U6798 (N_6798,N_5222,N_4119);
nand U6799 (N_6799,N_3719,N_4892);
or U6800 (N_6800,N_4976,N_3923);
nor U6801 (N_6801,N_4922,N_5823);
nor U6802 (N_6802,N_4942,N_5272);
xor U6803 (N_6803,N_3837,N_5185);
nand U6804 (N_6804,N_4776,N_4934);
xor U6805 (N_6805,N_5092,N_5599);
nand U6806 (N_6806,N_3646,N_3096);
nor U6807 (N_6807,N_4133,N_4423);
nand U6808 (N_6808,N_3902,N_4508);
nand U6809 (N_6809,N_5810,N_4638);
xor U6810 (N_6810,N_3486,N_5816);
and U6811 (N_6811,N_4950,N_3135);
or U6812 (N_6812,N_5062,N_4771);
nor U6813 (N_6813,N_5855,N_3315);
and U6814 (N_6814,N_5904,N_4781);
xor U6815 (N_6815,N_4916,N_4957);
or U6816 (N_6816,N_3751,N_3988);
nand U6817 (N_6817,N_5422,N_3747);
nand U6818 (N_6818,N_4845,N_3192);
xnor U6819 (N_6819,N_4876,N_3408);
nand U6820 (N_6820,N_4416,N_5845);
xnor U6821 (N_6821,N_5609,N_4847);
nor U6822 (N_6822,N_3343,N_4794);
xnor U6823 (N_6823,N_5880,N_4765);
or U6824 (N_6824,N_4566,N_4481);
and U6825 (N_6825,N_4721,N_3237);
xnor U6826 (N_6826,N_3378,N_3874);
or U6827 (N_6827,N_4918,N_4286);
nor U6828 (N_6828,N_4308,N_4259);
nor U6829 (N_6829,N_4316,N_4153);
nor U6830 (N_6830,N_4101,N_4536);
and U6831 (N_6831,N_4725,N_3651);
nand U6832 (N_6832,N_3846,N_4983);
or U6833 (N_6833,N_5544,N_5965);
xnor U6834 (N_6834,N_4361,N_4367);
and U6835 (N_6835,N_4450,N_3790);
nor U6836 (N_6836,N_3432,N_4833);
or U6837 (N_6837,N_3978,N_5122);
and U6838 (N_6838,N_4334,N_3971);
nor U6839 (N_6839,N_5951,N_5322);
or U6840 (N_6840,N_3261,N_4310);
nor U6841 (N_6841,N_3348,N_3461);
and U6842 (N_6842,N_5413,N_5095);
nand U6843 (N_6843,N_3650,N_4656);
and U6844 (N_6844,N_5181,N_4565);
nand U6845 (N_6845,N_5997,N_4974);
nand U6846 (N_6846,N_4504,N_3744);
or U6847 (N_6847,N_4070,N_4618);
nor U6848 (N_6848,N_4647,N_4356);
xor U6849 (N_6849,N_4028,N_5786);
nor U6850 (N_6850,N_5045,N_3350);
nor U6851 (N_6851,N_3555,N_5961);
nand U6852 (N_6852,N_3384,N_3623);
and U6853 (N_6853,N_3250,N_4337);
or U6854 (N_6854,N_3640,N_3984);
nor U6855 (N_6855,N_5906,N_3108);
or U6856 (N_6856,N_3006,N_4349);
and U6857 (N_6857,N_3076,N_5871);
and U6858 (N_6858,N_3380,N_5864);
or U6859 (N_6859,N_5639,N_3110);
or U6860 (N_6860,N_5400,N_3506);
nor U6861 (N_6861,N_3253,N_4247);
xor U6862 (N_6862,N_3567,N_4374);
xnor U6863 (N_6863,N_5764,N_3878);
nand U6864 (N_6864,N_5727,N_3774);
and U6865 (N_6865,N_5326,N_3209);
and U6866 (N_6866,N_5012,N_4391);
nand U6867 (N_6867,N_4798,N_3077);
nor U6868 (N_6868,N_4596,N_3973);
nand U6869 (N_6869,N_5869,N_4197);
xor U6870 (N_6870,N_4676,N_3010);
or U6871 (N_6871,N_5336,N_4068);
and U6872 (N_6872,N_3992,N_5479);
nor U6873 (N_6873,N_5747,N_5999);
or U6874 (N_6874,N_4797,N_5214);
xor U6875 (N_6875,N_4812,N_5283);
nor U6876 (N_6876,N_3521,N_4044);
and U6877 (N_6877,N_4467,N_4592);
nand U6878 (N_6878,N_3552,N_5734);
and U6879 (N_6879,N_4648,N_4168);
xnor U6880 (N_6880,N_3026,N_3341);
nand U6881 (N_6881,N_5672,N_3142);
xnor U6882 (N_6882,N_4741,N_3082);
or U6883 (N_6883,N_3400,N_4616);
nand U6884 (N_6884,N_5015,N_4993);
nand U6885 (N_6885,N_5950,N_5009);
nand U6886 (N_6886,N_3853,N_3333);
nand U6887 (N_6887,N_3540,N_5691);
nor U6888 (N_6888,N_4022,N_4738);
nor U6889 (N_6889,N_3582,N_5711);
and U6890 (N_6890,N_3182,N_4947);
or U6891 (N_6891,N_4799,N_4955);
xnor U6892 (N_6892,N_5900,N_4273);
xor U6893 (N_6893,N_3821,N_5407);
and U6894 (N_6894,N_3832,N_4312);
and U6895 (N_6895,N_3268,N_5893);
nand U6896 (N_6896,N_5179,N_4412);
nand U6897 (N_6897,N_4998,N_4850);
xnor U6898 (N_6898,N_5324,N_5039);
nand U6899 (N_6899,N_5584,N_3740);
nor U6900 (N_6900,N_4415,N_3240);
or U6901 (N_6901,N_5839,N_5670);
and U6902 (N_6902,N_3386,N_3019);
xnor U6903 (N_6903,N_4217,N_5142);
nand U6904 (N_6904,N_3419,N_3025);
nand U6905 (N_6905,N_4379,N_3063);
nand U6906 (N_6906,N_3805,N_3592);
xnor U6907 (N_6907,N_3947,N_3095);
and U6908 (N_6908,N_4278,N_4254);
nand U6909 (N_6909,N_4529,N_3803);
nand U6910 (N_6910,N_3430,N_5894);
nand U6911 (N_6911,N_3542,N_5085);
xnor U6912 (N_6912,N_3930,N_5667);
xor U6913 (N_6913,N_5109,N_3966);
nor U6914 (N_6914,N_4231,N_5450);
xor U6915 (N_6915,N_3569,N_4806);
nor U6916 (N_6916,N_4323,N_5721);
nor U6917 (N_6917,N_5116,N_3194);
nand U6918 (N_6918,N_5963,N_3244);
and U6919 (N_6919,N_4913,N_3423);
or U6920 (N_6920,N_3467,N_5818);
and U6921 (N_6921,N_5497,N_4347);
xnor U6922 (N_6922,N_3897,N_3659);
nand U6923 (N_6923,N_3776,N_3705);
nor U6924 (N_6924,N_3845,N_3610);
or U6925 (N_6925,N_5025,N_4269);
nand U6926 (N_6926,N_3898,N_3558);
xnor U6927 (N_6927,N_3014,N_4187);
nor U6928 (N_6928,N_3848,N_5577);
and U6929 (N_6929,N_3736,N_5592);
xnor U6930 (N_6930,N_4785,N_5007);
xor U6931 (N_6931,N_5708,N_5046);
and U6932 (N_6932,N_3393,N_3392);
nand U6933 (N_6933,N_4910,N_5200);
or U6934 (N_6934,N_3922,N_3027);
or U6935 (N_6935,N_4026,N_5931);
nand U6936 (N_6936,N_5031,N_3403);
nand U6937 (N_6937,N_4677,N_4291);
and U6938 (N_6938,N_4982,N_5132);
nand U6939 (N_6939,N_4735,N_3066);
xnor U6940 (N_6940,N_3061,N_3959);
nor U6941 (N_6941,N_5421,N_5956);
nor U6942 (N_6942,N_4229,N_5524);
nor U6943 (N_6943,N_4439,N_5674);
nand U6944 (N_6944,N_5226,N_5617);
and U6945 (N_6945,N_3216,N_5760);
xor U6946 (N_6946,N_5827,N_5013);
and U6947 (N_6947,N_5774,N_4066);
nand U6948 (N_6948,N_4689,N_5285);
xnor U6949 (N_6949,N_3338,N_4144);
xnor U6950 (N_6950,N_3669,N_5744);
and U6951 (N_6951,N_4425,N_4548);
xor U6952 (N_6952,N_4889,N_4486);
or U6953 (N_6953,N_5104,N_3696);
nand U6954 (N_6954,N_5628,N_3479);
nand U6955 (N_6955,N_4832,N_3115);
nor U6956 (N_6956,N_5957,N_4181);
nor U6957 (N_6957,N_5669,N_5331);
nor U6958 (N_6958,N_3647,N_4137);
nor U6959 (N_6959,N_4956,N_5055);
xor U6960 (N_6960,N_4014,N_3273);
and U6961 (N_6961,N_5257,N_5512);
nor U6962 (N_6962,N_5913,N_3662);
nor U6963 (N_6963,N_3193,N_5654);
and U6964 (N_6964,N_3282,N_4192);
and U6965 (N_6965,N_5777,N_4545);
nor U6966 (N_6966,N_4198,N_5128);
xnor U6967 (N_6967,N_4413,N_5946);
or U6968 (N_6968,N_5486,N_4813);
nor U6969 (N_6969,N_5038,N_5133);
or U6970 (N_6970,N_5074,N_5502);
xnor U6971 (N_6971,N_4838,N_5812);
and U6972 (N_6972,N_5228,N_4967);
nor U6973 (N_6973,N_4409,N_4703);
and U6974 (N_6974,N_5971,N_3829);
nor U6975 (N_6975,N_4135,N_5598);
nand U6976 (N_6976,N_5588,N_3620);
xnor U6977 (N_6977,N_4071,N_5648);
nand U6978 (N_6978,N_5357,N_4284);
and U6979 (N_6979,N_3234,N_5773);
xor U6980 (N_6980,N_3156,N_5027);
xor U6981 (N_6981,N_3967,N_3451);
nand U6982 (N_6982,N_4006,N_3996);
nor U6983 (N_6983,N_4885,N_3208);
or U6984 (N_6984,N_5115,N_3021);
nor U6985 (N_6985,N_3713,N_3779);
or U6986 (N_6986,N_3301,N_3186);
nor U6987 (N_6987,N_3815,N_5123);
or U6988 (N_6988,N_4329,N_5610);
and U6989 (N_6989,N_3926,N_5401);
xnor U6990 (N_6990,N_5467,N_5044);
nand U6991 (N_6991,N_5459,N_5278);
xor U6992 (N_6992,N_3433,N_5572);
xnor U6993 (N_6993,N_3001,N_3658);
nor U6994 (N_6994,N_4085,N_5632);
or U6995 (N_6995,N_5328,N_3642);
or U6996 (N_6996,N_3595,N_4511);
and U6997 (N_6997,N_3752,N_4774);
nand U6998 (N_6998,N_5078,N_3635);
nor U6999 (N_6999,N_5218,N_5680);
or U7000 (N_7000,N_5751,N_3317);
xor U7001 (N_7001,N_4494,N_4630);
xor U7002 (N_7002,N_4699,N_5594);
nand U7003 (N_7003,N_3844,N_3551);
and U7004 (N_7004,N_3641,N_5207);
nand U7005 (N_7005,N_4650,N_4866);
nor U7006 (N_7006,N_5849,N_3427);
nand U7007 (N_7007,N_5924,N_5921);
or U7008 (N_7008,N_3213,N_3176);
or U7009 (N_7009,N_3202,N_3985);
or U7010 (N_7010,N_4597,N_4224);
nor U7011 (N_7011,N_4112,N_3613);
nand U7012 (N_7012,N_5158,N_5113);
and U7013 (N_7013,N_5170,N_3068);
nand U7014 (N_7014,N_5856,N_4256);
nand U7015 (N_7015,N_4533,N_4281);
and U7016 (N_7016,N_4554,N_3127);
nand U7017 (N_7017,N_4633,N_3615);
xor U7018 (N_7018,N_5761,N_5466);
and U7019 (N_7019,N_5954,N_3684);
or U7020 (N_7020,N_4819,N_4605);
nor U7021 (N_7021,N_5619,N_5269);
nand U7022 (N_7022,N_4021,N_4818);
nand U7023 (N_7023,N_3648,N_5277);
xnor U7024 (N_7024,N_4986,N_5341);
nand U7025 (N_7025,N_5590,N_3891);
or U7026 (N_7026,N_5120,N_4053);
xnor U7027 (N_7027,N_4965,N_3977);
nor U7028 (N_7028,N_5339,N_4104);
or U7029 (N_7029,N_4406,N_4745);
xor U7030 (N_7030,N_5360,N_3539);
nor U7031 (N_7031,N_5160,N_5563);
or U7032 (N_7032,N_5414,N_3102);
xor U7033 (N_7033,N_5346,N_3107);
nor U7034 (N_7034,N_3324,N_4582);
or U7035 (N_7035,N_5195,N_3957);
and U7036 (N_7036,N_5803,N_5533);
xnor U7037 (N_7037,N_4173,N_5853);
or U7038 (N_7038,N_3013,N_3354);
and U7039 (N_7039,N_5210,N_3999);
and U7040 (N_7040,N_5859,N_3008);
xor U7041 (N_7041,N_4939,N_3256);
nand U7042 (N_7042,N_4883,N_3058);
or U7043 (N_7043,N_5865,N_5135);
or U7044 (N_7044,N_3871,N_5897);
xnor U7045 (N_7045,N_4442,N_3326);
xnor U7046 (N_7046,N_5446,N_4691);
xor U7047 (N_7047,N_3057,N_5728);
xnor U7048 (N_7048,N_5310,N_4462);
and U7049 (N_7049,N_4553,N_5649);
or U7050 (N_7050,N_5087,N_5944);
and U7051 (N_7051,N_5408,N_3663);
nand U7052 (N_7052,N_4743,N_4333);
and U7053 (N_7053,N_3673,N_3915);
or U7054 (N_7054,N_4666,N_3376);
xor U7055 (N_7055,N_5605,N_5507);
and U7056 (N_7056,N_5866,N_5024);
nor U7057 (N_7057,N_5215,N_5861);
or U7058 (N_7058,N_4555,N_5755);
or U7059 (N_7059,N_3397,N_4629);
xnor U7060 (N_7060,N_4087,N_5887);
nand U7061 (N_7061,N_3919,N_5872);
or U7062 (N_7062,N_3002,N_5595);
and U7063 (N_7063,N_5327,N_5064);
or U7064 (N_7064,N_3039,N_3526);
and U7065 (N_7065,N_3498,N_3765);
xnor U7066 (N_7066,N_4559,N_3952);
xor U7067 (N_7067,N_4948,N_3033);
or U7068 (N_7068,N_5157,N_3314);
and U7069 (N_7069,N_5612,N_5096);
nand U7070 (N_7070,N_4877,N_5618);
nand U7071 (N_7071,N_3729,N_5258);
nand U7072 (N_7072,N_5395,N_4653);
xor U7073 (N_7073,N_3030,N_4810);
xnor U7074 (N_7074,N_4154,N_3672);
and U7075 (N_7075,N_3792,N_4351);
or U7076 (N_7076,N_4261,N_5172);
nand U7077 (N_7077,N_4032,N_3780);
nand U7078 (N_7078,N_5235,N_4335);
and U7079 (N_7079,N_4371,N_5371);
nand U7080 (N_7080,N_4824,N_5460);
and U7081 (N_7081,N_5907,N_4784);
and U7082 (N_7082,N_3143,N_5842);
nor U7083 (N_7083,N_3586,N_5444);
xor U7084 (N_7084,N_4804,N_5838);
xor U7085 (N_7085,N_4540,N_3855);
and U7086 (N_7086,N_3269,N_4456);
and U7087 (N_7087,N_5693,N_5347);
or U7088 (N_7088,N_4103,N_4364);
nor U7089 (N_7089,N_3227,N_4440);
xnor U7090 (N_7090,N_5429,N_5636);
or U7091 (N_7091,N_5585,N_3035);
or U7092 (N_7092,N_5996,N_4905);
xor U7093 (N_7093,N_3969,N_5050);
and U7094 (N_7094,N_5874,N_4800);
or U7095 (N_7095,N_3299,N_4158);
and U7096 (N_7096,N_3970,N_5559);
xnor U7097 (N_7097,N_3691,N_4705);
nand U7098 (N_7098,N_4443,N_5083);
xor U7099 (N_7099,N_5080,N_5879);
nor U7100 (N_7100,N_3914,N_4293);
or U7101 (N_7101,N_4520,N_3434);
nand U7102 (N_7102,N_5242,N_4437);
or U7103 (N_7103,N_4180,N_4484);
nor U7104 (N_7104,N_4980,N_4392);
xnor U7105 (N_7105,N_3435,N_4384);
nand U7106 (N_7106,N_3712,N_5793);
or U7107 (N_7107,N_5312,N_4285);
or U7108 (N_7108,N_3424,N_4660);
xor U7109 (N_7109,N_4255,N_3576);
xor U7110 (N_7110,N_3678,N_4326);
nand U7111 (N_7111,N_3949,N_3357);
nand U7112 (N_7112,N_5282,N_3907);
and U7113 (N_7113,N_3675,N_3656);
and U7114 (N_7114,N_4341,N_3711);
and U7115 (N_7115,N_4325,N_5213);
nor U7116 (N_7116,N_5749,N_5510);
or U7117 (N_7117,N_4901,N_4475);
and U7118 (N_7118,N_5713,N_4959);
xor U7119 (N_7119,N_5806,N_4468);
xnor U7120 (N_7120,N_3447,N_4822);
nor U7121 (N_7121,N_5748,N_4243);
nand U7122 (N_7122,N_3340,N_4034);
or U7123 (N_7123,N_3899,N_4907);
nand U7124 (N_7124,N_4668,N_4121);
xnor U7125 (N_7125,N_3119,N_4525);
nand U7126 (N_7126,N_4718,N_5992);
xnor U7127 (N_7127,N_5245,N_5937);
and U7128 (N_7128,N_4828,N_3591);
nand U7129 (N_7129,N_5399,N_5356);
nand U7130 (N_7130,N_5575,N_4420);
or U7131 (N_7131,N_5391,N_5182);
or U7132 (N_7132,N_5633,N_3850);
or U7133 (N_7133,N_4252,N_5262);
nand U7134 (N_7134,N_4362,N_5902);
or U7135 (N_7135,N_3071,N_3657);
xnor U7136 (N_7136,N_5276,N_5136);
or U7137 (N_7137,N_5313,N_4483);
nand U7138 (N_7138,N_3820,N_4421);
nand U7139 (N_7139,N_4009,N_5296);
nor U7140 (N_7140,N_3425,N_4712);
xnor U7141 (N_7141,N_5552,N_5896);
or U7142 (N_7142,N_5623,N_4911);
and U7143 (N_7143,N_4954,N_3519);
nand U7144 (N_7144,N_3556,N_4126);
and U7145 (N_7145,N_4344,N_3091);
and U7146 (N_7146,N_3626,N_3881);
nor U7147 (N_7147,N_5846,N_3121);
xor U7148 (N_7148,N_5500,N_5168);
xnor U7149 (N_7149,N_3956,N_4232);
xnor U7150 (N_7150,N_3958,N_3146);
nand U7151 (N_7151,N_5229,N_3773);
and U7152 (N_7152,N_4702,N_5692);
nor U7153 (N_7153,N_5789,N_5315);
and U7154 (N_7154,N_5063,N_4991);
and U7155 (N_7155,N_5771,N_3917);
or U7156 (N_7156,N_5349,N_4073);
nand U7157 (N_7157,N_3624,N_3147);
or U7158 (N_7158,N_3980,N_4581);
or U7159 (N_7159,N_5201,N_3931);
nand U7160 (N_7160,N_3042,N_4313);
or U7161 (N_7161,N_5712,N_4788);
or U7162 (N_7162,N_4306,N_5688);
xnor U7163 (N_7163,N_3469,N_3287);
xnor U7164 (N_7164,N_5317,N_4767);
xor U7165 (N_7165,N_3617,N_5840);
nor U7166 (N_7166,N_3388,N_5117);
xnor U7167 (N_7167,N_3535,N_5404);
or U7168 (N_7168,N_3132,N_3293);
nand U7169 (N_7169,N_5600,N_5607);
and U7170 (N_7170,N_4174,N_3170);
nor U7171 (N_7171,N_4927,N_3353);
nor U7172 (N_7172,N_4125,N_5037);
nor U7173 (N_7173,N_4201,N_3113);
or U7174 (N_7174,N_5496,N_4179);
xnor U7175 (N_7175,N_5293,N_3677);
and U7176 (N_7176,N_5821,N_5261);
and U7177 (N_7177,N_3332,N_5547);
and U7178 (N_7178,N_5862,N_3290);
xnor U7179 (N_7179,N_4973,N_3565);
nand U7180 (N_7180,N_5521,N_4100);
nand U7181 (N_7181,N_5940,N_3088);
nand U7182 (N_7182,N_5240,N_5829);
and U7183 (N_7183,N_4230,N_3880);
nand U7184 (N_7184,N_4690,N_3295);
or U7185 (N_7185,N_5903,N_3517);
and U7186 (N_7186,N_3734,N_5847);
and U7187 (N_7187,N_3289,N_3494);
or U7188 (N_7188,N_4604,N_5205);
and U7189 (N_7189,N_3994,N_5695);
nand U7190 (N_7190,N_5433,N_4789);
xor U7191 (N_7191,N_3756,N_4095);
nor U7192 (N_7192,N_3062,N_3409);
nand U7193 (N_7193,N_5359,N_3746);
or U7194 (N_7194,N_3813,N_5110);
and U7195 (N_7195,N_5378,N_4031);
nand U7196 (N_7196,N_3697,N_5475);
and U7197 (N_7197,N_3989,N_3979);
or U7198 (N_7198,N_3852,N_5418);
and U7199 (N_7199,N_3895,N_4830);
or U7200 (N_7200,N_5994,N_4114);
and U7201 (N_7201,N_5686,N_4801);
nor U7202 (N_7202,N_5398,N_4989);
nand U7203 (N_7203,N_5884,N_5682);
xnor U7204 (N_7204,N_5527,N_5125);
nand U7205 (N_7205,N_3942,N_4821);
xor U7206 (N_7206,N_5094,N_3004);
or U7207 (N_7207,N_4854,N_3396);
nand U7208 (N_7208,N_3787,N_3538);
nand U7209 (N_7209,N_5875,N_4716);
nor U7210 (N_7210,N_5753,N_4029);
or U7211 (N_7211,N_5481,N_5291);
or U7212 (N_7212,N_4309,N_3587);
xor U7213 (N_7213,N_3667,N_5641);
nand U7214 (N_7214,N_3936,N_4621);
nand U7215 (N_7215,N_4193,N_4298);
or U7216 (N_7216,N_3509,N_5243);
and U7217 (N_7217,N_5093,N_5456);
or U7218 (N_7218,N_3488,N_3649);
or U7219 (N_7219,N_4542,N_4311);
and U7220 (N_7220,N_5972,N_5962);
nor U7221 (N_7221,N_5300,N_3951);
xnor U7222 (N_7222,N_3559,N_3819);
nor U7223 (N_7223,N_5644,N_4631);
xor U7224 (N_7224,N_5383,N_5118);
xor U7225 (N_7225,N_4040,N_3778);
xor U7226 (N_7226,N_5302,N_5379);
nor U7227 (N_7227,N_4917,N_4787);
and U7228 (N_7228,N_5376,N_5364);
or U7229 (N_7229,N_3653,N_3528);
nand U7230 (N_7230,N_3398,N_3636);
or U7231 (N_7231,N_4951,N_5480);
or U7232 (N_7232,N_5382,N_4172);
nor U7233 (N_7233,N_3252,N_4904);
nand U7234 (N_7234,N_3665,N_5102);
or U7235 (N_7235,N_3757,N_4990);
nand U7236 (N_7236,N_4895,N_4770);
xor U7237 (N_7237,N_5704,N_3246);
nand U7238 (N_7238,N_3794,N_3612);
nand U7239 (N_7239,N_5807,N_3330);
and U7240 (N_7240,N_3896,N_4317);
nor U7241 (N_7241,N_3802,N_4129);
nor U7242 (N_7242,N_4995,N_3431);
nor U7243 (N_7243,N_3838,N_3889);
nand U7244 (N_7244,N_3140,N_4381);
or U7245 (N_7245,N_4140,N_4521);
and U7246 (N_7246,N_4246,N_4831);
and U7247 (N_7247,N_5509,N_3804);
xor U7248 (N_7248,N_4080,N_4729);
or U7249 (N_7249,N_5854,N_3900);
nand U7250 (N_7250,N_5056,N_4105);
nor U7251 (N_7251,N_3458,N_4502);
or U7252 (N_7252,N_5960,N_3051);
nor U7253 (N_7253,N_5016,N_5792);
or U7254 (N_7254,N_5918,N_5490);
xor U7255 (N_7255,N_3462,N_3407);
or U7256 (N_7256,N_5912,N_4342);
and U7257 (N_7257,N_3621,N_4909);
nor U7258 (N_7258,N_3941,N_4882);
or U7259 (N_7259,N_5204,N_4328);
and U7260 (N_7260,N_3873,N_4717);
and U7261 (N_7261,N_5769,N_3404);
or U7262 (N_7262,N_5411,N_3180);
nand U7263 (N_7263,N_3911,N_3499);
or U7264 (N_7264,N_5047,N_5089);
or U7265 (N_7265,N_5035,N_4872);
nand U7266 (N_7266,N_4587,N_5234);
or U7267 (N_7267,N_4373,N_3801);
xnor U7268 (N_7268,N_3948,N_5953);
nor U7269 (N_7269,N_3015,N_3339);
and U7270 (N_7270,N_3201,N_5743);
xor U7271 (N_7271,N_4478,N_3972);
nor U7272 (N_7272,N_5858,N_3596);
and U7273 (N_7273,N_3597,N_5895);
and U7274 (N_7274,N_3571,N_4758);
nor U7275 (N_7275,N_3939,N_4260);
and U7276 (N_7276,N_3060,N_4460);
xnor U7277 (N_7277,N_4143,N_3455);
nor U7278 (N_7278,N_5925,N_5883);
xnor U7279 (N_7279,N_3258,N_4393);
nor U7280 (N_7280,N_4811,N_4297);
and U7281 (N_7281,N_4839,N_3600);
xor U7282 (N_7282,N_3961,N_4299);
nand U7283 (N_7283,N_3275,N_4972);
nor U7284 (N_7284,N_4041,N_4926);
xor U7285 (N_7285,N_5597,N_3443);
or U7286 (N_7286,N_5173,N_3809);
and U7287 (N_7287,N_4354,N_3604);
or U7288 (N_7288,N_4753,N_4262);
nand U7289 (N_7289,N_3654,N_3475);
nand U7290 (N_7290,N_3286,N_3047);
nor U7291 (N_7291,N_3163,N_5886);
or U7292 (N_7292,N_3865,N_3267);
nor U7293 (N_7293,N_5757,N_3144);
xnor U7294 (N_7294,N_5615,N_5425);
nand U7295 (N_7295,N_3089,N_4366);
and U7296 (N_7296,N_5140,N_5169);
and U7297 (N_7297,N_3825,N_5778);
xnor U7298 (N_7298,N_3905,N_3355);
xnor U7299 (N_7299,N_5911,N_5923);
and U7300 (N_7300,N_3044,N_5386);
nor U7301 (N_7301,N_4315,N_4613);
xor U7302 (N_7302,N_3316,N_4191);
and U7303 (N_7303,N_3148,N_3016);
nand U7304 (N_7304,N_4248,N_5707);
or U7305 (N_7305,N_3198,N_3944);
nand U7306 (N_7306,N_3318,N_4331);
nor U7307 (N_7307,N_3758,N_4208);
xor U7308 (N_7308,N_5538,N_4389);
or U7309 (N_7309,N_5114,N_5255);
nor U7310 (N_7310,N_4339,N_4609);
nor U7311 (N_7311,N_4868,N_5850);
nand U7312 (N_7312,N_5582,N_5531);
nor U7313 (N_7313,N_4841,N_3692);
nor U7314 (N_7314,N_3072,N_3271);
nand U7315 (N_7315,N_5867,N_5392);
nor U7316 (N_7316,N_4541,N_5646);
nand U7317 (N_7317,N_4448,N_3453);
and U7318 (N_7318,N_4493,N_4875);
and U7319 (N_7319,N_3449,N_4018);
nand U7320 (N_7320,N_5384,N_3329);
xor U7321 (N_7321,N_3414,N_4452);
or U7322 (N_7322,N_4780,N_4867);
or U7323 (N_7323,N_4654,N_4472);
and U7324 (N_7324,N_3122,N_5949);
nor U7325 (N_7325,N_3799,N_3570);
nand U7326 (N_7326,N_5634,N_3893);
nand U7327 (N_7327,N_5367,N_3241);
nor U7328 (N_7328,N_3065,N_5198);
xor U7329 (N_7329,N_3231,N_5843);
nand U7330 (N_7330,N_3391,N_3382);
nand U7331 (N_7331,N_4723,N_3795);
or U7332 (N_7332,N_3456,N_4322);
and U7333 (N_7333,N_3000,N_4499);
or U7334 (N_7334,N_4792,N_3843);
and U7335 (N_7335,N_5220,N_5694);
xnor U7336 (N_7336,N_3225,N_4682);
or U7337 (N_7337,N_3319,N_4024);
xor U7338 (N_7338,N_4570,N_3164);
xnor U7339 (N_7339,N_4583,N_5355);
or U7340 (N_7340,N_5699,N_3320);
nand U7341 (N_7341,N_4128,N_5660);
xnor U7342 (N_7342,N_5076,N_4623);
or U7343 (N_7343,N_4600,N_5286);
nand U7344 (N_7344,N_4856,N_5776);
nand U7345 (N_7345,N_3581,N_3099);
nand U7346 (N_7346,N_3490,N_5287);
and U7347 (N_7347,N_3043,N_3351);
and U7348 (N_7348,N_5099,N_4065);
nand U7349 (N_7349,N_5144,N_3152);
nand U7350 (N_7350,N_5596,N_3940);
and U7351 (N_7351,N_3918,N_5785);
xor U7352 (N_7352,N_3983,N_5206);
and U7353 (N_7353,N_4537,N_5239);
and U7354 (N_7354,N_5784,N_4360);
or U7355 (N_7355,N_3276,N_5767);
or U7356 (N_7356,N_3266,N_3501);
or U7357 (N_7357,N_4757,N_4683);
nor U7358 (N_7358,N_5108,N_3416);
and U7359 (N_7359,N_4157,N_5567);
nand U7360 (N_7360,N_3321,N_5188);
nand U7361 (N_7361,N_3130,N_5363);
xnor U7362 (N_7362,N_3041,N_4594);
or U7363 (N_7363,N_3457,N_4578);
and U7364 (N_7364,N_5457,N_5176);
nand U7365 (N_7365,N_5611,N_4908);
nor U7366 (N_7366,N_3204,N_5493);
and U7367 (N_7367,N_4228,N_4739);
and U7368 (N_7368,N_4433,N_3536);
xor U7369 (N_7369,N_3472,N_3575);
or U7370 (N_7370,N_5863,N_3839);
xnor U7371 (N_7371,N_4893,N_4346);
xor U7372 (N_7372,N_4759,N_4498);
and U7373 (N_7373,N_5443,N_4969);
nand U7374 (N_7374,N_3738,N_4971);
and U7375 (N_7375,N_3606,N_3671);
or U7376 (N_7376,N_3362,N_5635);
xnor U7377 (N_7377,N_4005,N_4925);
or U7378 (N_7378,N_4728,N_5709);
and U7379 (N_7379,N_4490,N_4530);
nor U7380 (N_7380,N_4887,N_4288);
xor U7381 (N_7381,N_5051,N_4108);
and U7382 (N_7382,N_3199,N_4422);
or U7383 (N_7383,N_5581,N_5435);
xnor U7384 (N_7384,N_5106,N_5733);
or U7385 (N_7385,N_5487,N_5155);
and U7386 (N_7386,N_4449,N_3279);
xnor U7387 (N_7387,N_4294,N_4673);
nand U7388 (N_7388,N_4127,N_5107);
xnor U7389 (N_7389,N_5795,N_4599);
nor U7390 (N_7390,N_5066,N_3024);
and U7391 (N_7391,N_5177,N_5149);
and U7392 (N_7392,N_5174,N_5589);
nand U7393 (N_7393,N_3257,N_3379);
or U7394 (N_7394,N_5991,N_3664);
and U7395 (N_7395,N_4084,N_5284);
and U7396 (N_7396,N_3722,N_3682);
nand U7397 (N_7397,N_3215,N_5556);
nand U7398 (N_7398,N_4401,N_3159);
and U7399 (N_7399,N_3480,N_5033);
nand U7400 (N_7400,N_3563,N_4961);
xor U7401 (N_7401,N_4861,N_5892);
xnor U7402 (N_7402,N_3583,N_3104);
nor U7403 (N_7403,N_4492,N_4870);
or U7404 (N_7404,N_5353,N_3685);
or U7405 (N_7405,N_5137,N_3522);
nor U7406 (N_7406,N_4036,N_3153);
nand U7407 (N_7407,N_3523,N_5230);
xor U7408 (N_7408,N_3118,N_4659);
or U7409 (N_7409,N_4171,N_4823);
and U7410 (N_7410,N_4573,N_5518);
or U7411 (N_7411,N_5779,N_3011);
nor U7412 (N_7412,N_5217,N_5848);
and U7413 (N_7413,N_5726,N_5023);
nand U7414 (N_7414,N_4263,N_3070);
or U7415 (N_7415,N_4994,N_3421);
and U7416 (N_7416,N_5448,N_3879);
and U7417 (N_7417,N_3505,N_4749);
and U7418 (N_7418,N_4083,N_5145);
nor U7419 (N_7419,N_4150,N_4184);
or U7420 (N_7420,N_5910,N_4435);
and U7421 (N_7421,N_4048,N_5052);
nand U7422 (N_7422,N_3854,N_4734);
nand U7423 (N_7423,N_4685,N_4751);
and U7424 (N_7424,N_3003,N_3912);
nand U7425 (N_7425,N_5943,N_4338);
nand U7426 (N_7426,N_5791,N_5540);
or U7427 (N_7427,N_4207,N_5072);
xor U7428 (N_7428,N_4675,N_3830);
nor U7429 (N_7429,N_3098,N_3334);
nor U7430 (N_7430,N_4234,N_5103);
nand U7431 (N_7431,N_4713,N_3081);
and U7432 (N_7432,N_5513,N_4038);
or U7433 (N_7433,N_3887,N_3760);
nand U7434 (N_7434,N_5775,N_3894);
and U7435 (N_7435,N_3185,N_3962);
nand U7436 (N_7436,N_4453,N_3247);
nand U7437 (N_7437,N_5049,N_5306);
nand U7438 (N_7438,N_4696,N_3525);
xor U7439 (N_7439,N_3533,N_4069);
nand U7440 (N_7440,N_3161,N_3699);
xor U7441 (N_7441,N_4779,N_4218);
nor U7442 (N_7442,N_5742,N_3191);
and U7443 (N_7443,N_3385,N_3798);
nor U7444 (N_7444,N_3503,N_4205);
nand U7445 (N_7445,N_5529,N_5643);
or U7446 (N_7446,N_4598,N_3550);
nor U7447 (N_7447,N_3028,N_3387);
and U7448 (N_7448,N_3465,N_5499);
nor U7449 (N_7449,N_5710,N_4879);
and U7450 (N_7450,N_4390,N_3644);
nand U7451 (N_7451,N_5416,N_4820);
xnor U7452 (N_7452,N_3716,N_3704);
nor U7453 (N_7453,N_5470,N_5666);
nand U7454 (N_7454,N_5668,N_5162);
nor U7455 (N_7455,N_4863,N_3171);
nand U7456 (N_7456,N_5586,N_5515);
xor U7457 (N_7457,N_4742,N_3638);
nor U7458 (N_7458,N_5802,N_4480);
and U7459 (N_7459,N_5061,N_4896);
or U7460 (N_7460,N_4061,N_5420);
xor U7461 (N_7461,N_5920,N_5631);
and U7462 (N_7462,N_5977,N_3097);
and U7463 (N_7463,N_3444,N_5319);
nor U7464 (N_7464,N_4807,N_5340);
nand U7465 (N_7465,N_5021,N_5320);
nand U7466 (N_7466,N_5192,N_4849);
or U7467 (N_7467,N_3763,N_5073);
xnor U7468 (N_7468,N_5933,N_4426);
and U7469 (N_7469,N_3548,N_5759);
nand U7470 (N_7470,N_5338,N_5593);
or U7471 (N_7471,N_4783,N_3577);
or U7472 (N_7472,N_3220,N_3344);
or U7473 (N_7473,N_4747,N_3395);
nor U7474 (N_7474,N_4155,N_5723);
nand U7475 (N_7475,N_5730,N_4669);
xnor U7476 (N_7476,N_3087,N_4214);
nor U7477 (N_7477,N_3373,N_3173);
or U7478 (N_7478,N_4399,N_3754);
xnor U7479 (N_7479,N_3262,N_5057);
or U7480 (N_7480,N_5799,N_3100);
or U7481 (N_7481,N_4350,N_3735);
nand U7482 (N_7482,N_5256,N_4640);
nand U7483 (N_7483,N_3938,N_3599);
nor U7484 (N_7484,N_3851,N_3371);
and U7485 (N_7485,N_3816,N_3111);
and U7486 (N_7486,N_3903,N_3627);
and U7487 (N_7487,N_3808,N_4531);
and U7488 (N_7488,N_3285,N_5134);
and U7489 (N_7489,N_3867,N_4147);
nand U7490 (N_7490,N_3892,N_3375);
nand U7491 (N_7491,N_3206,N_3660);
xor U7492 (N_7492,N_5299,N_5279);
or U7493 (N_7493,N_5036,N_4079);
and U7494 (N_7494,N_3055,N_3909);
and U7495 (N_7495,N_3827,N_5576);
or U7496 (N_7496,N_3092,N_3594);
xor U7497 (N_7497,N_4400,N_5770);
nor U7498 (N_7498,N_3383,N_5988);
and U7499 (N_7499,N_5536,N_5190);
or U7500 (N_7500,N_3477,N_4855);
or U7501 (N_7501,N_5900,N_4969);
nor U7502 (N_7502,N_4652,N_3743);
xor U7503 (N_7503,N_3800,N_3106);
xnor U7504 (N_7504,N_3331,N_3303);
or U7505 (N_7505,N_5853,N_3239);
nor U7506 (N_7506,N_4774,N_3173);
nand U7507 (N_7507,N_3059,N_3140);
or U7508 (N_7508,N_3232,N_5881);
nand U7509 (N_7509,N_4309,N_5798);
xor U7510 (N_7510,N_4815,N_5777);
nand U7511 (N_7511,N_5401,N_4633);
nor U7512 (N_7512,N_5295,N_3700);
nand U7513 (N_7513,N_4831,N_3096);
and U7514 (N_7514,N_5549,N_3263);
nor U7515 (N_7515,N_3882,N_5889);
nor U7516 (N_7516,N_5312,N_4514);
or U7517 (N_7517,N_3443,N_4685);
xnor U7518 (N_7518,N_5596,N_3626);
xnor U7519 (N_7519,N_3507,N_5635);
xor U7520 (N_7520,N_3759,N_5304);
nor U7521 (N_7521,N_4751,N_4820);
nand U7522 (N_7522,N_3802,N_4542);
nand U7523 (N_7523,N_4839,N_4620);
or U7524 (N_7524,N_4074,N_4429);
xor U7525 (N_7525,N_3113,N_4403);
xor U7526 (N_7526,N_4115,N_3851);
and U7527 (N_7527,N_4573,N_4675);
nand U7528 (N_7528,N_4296,N_5328);
xnor U7529 (N_7529,N_4870,N_4230);
nand U7530 (N_7530,N_5646,N_4455);
nor U7531 (N_7531,N_3268,N_3470);
nand U7532 (N_7532,N_4838,N_3257);
or U7533 (N_7533,N_5425,N_5271);
xor U7534 (N_7534,N_5714,N_5645);
nor U7535 (N_7535,N_4678,N_3075);
or U7536 (N_7536,N_3994,N_5321);
nand U7537 (N_7537,N_5620,N_3674);
xor U7538 (N_7538,N_5093,N_4515);
nor U7539 (N_7539,N_3617,N_3071);
xor U7540 (N_7540,N_4119,N_3040);
xor U7541 (N_7541,N_5252,N_4907);
nand U7542 (N_7542,N_4546,N_5054);
and U7543 (N_7543,N_4113,N_3649);
or U7544 (N_7544,N_5257,N_3328);
and U7545 (N_7545,N_3786,N_4464);
xnor U7546 (N_7546,N_3614,N_3911);
nand U7547 (N_7547,N_3306,N_3403);
or U7548 (N_7548,N_4197,N_3948);
nor U7549 (N_7549,N_3962,N_4550);
xnor U7550 (N_7550,N_5982,N_3364);
nand U7551 (N_7551,N_5306,N_3684);
nand U7552 (N_7552,N_3485,N_5874);
xor U7553 (N_7553,N_5294,N_4292);
or U7554 (N_7554,N_5097,N_4768);
nor U7555 (N_7555,N_5408,N_4231);
nor U7556 (N_7556,N_5616,N_3943);
nand U7557 (N_7557,N_3626,N_3504);
nor U7558 (N_7558,N_5738,N_4831);
nand U7559 (N_7559,N_5481,N_4996);
nor U7560 (N_7560,N_3726,N_5807);
or U7561 (N_7561,N_3437,N_5094);
nand U7562 (N_7562,N_5318,N_3897);
and U7563 (N_7563,N_4485,N_3573);
or U7564 (N_7564,N_5892,N_5202);
xnor U7565 (N_7565,N_3142,N_3284);
nand U7566 (N_7566,N_3957,N_3186);
nand U7567 (N_7567,N_4567,N_4500);
xnor U7568 (N_7568,N_4945,N_5369);
and U7569 (N_7569,N_5019,N_3813);
xor U7570 (N_7570,N_3408,N_3461);
and U7571 (N_7571,N_3753,N_5110);
or U7572 (N_7572,N_4572,N_4018);
and U7573 (N_7573,N_3749,N_3005);
and U7574 (N_7574,N_4928,N_5363);
xnor U7575 (N_7575,N_4965,N_4142);
nand U7576 (N_7576,N_4673,N_3608);
and U7577 (N_7577,N_3030,N_4717);
nand U7578 (N_7578,N_3070,N_5552);
and U7579 (N_7579,N_5480,N_4319);
xor U7580 (N_7580,N_4903,N_4646);
xor U7581 (N_7581,N_4628,N_3987);
xnor U7582 (N_7582,N_3841,N_4829);
or U7583 (N_7583,N_4109,N_5345);
nand U7584 (N_7584,N_3503,N_3397);
nand U7585 (N_7585,N_3726,N_3420);
xor U7586 (N_7586,N_4199,N_3290);
and U7587 (N_7587,N_4317,N_3159);
and U7588 (N_7588,N_5125,N_3773);
or U7589 (N_7589,N_4148,N_4802);
and U7590 (N_7590,N_3233,N_4369);
or U7591 (N_7591,N_5894,N_5122);
and U7592 (N_7592,N_3550,N_4871);
xnor U7593 (N_7593,N_4943,N_3674);
nand U7594 (N_7594,N_5457,N_4624);
and U7595 (N_7595,N_5312,N_5995);
and U7596 (N_7596,N_5784,N_5391);
or U7597 (N_7597,N_4443,N_5116);
or U7598 (N_7598,N_5065,N_5002);
and U7599 (N_7599,N_3728,N_4303);
xnor U7600 (N_7600,N_4741,N_5293);
xnor U7601 (N_7601,N_3440,N_4373);
xor U7602 (N_7602,N_4228,N_5035);
or U7603 (N_7603,N_3778,N_4431);
and U7604 (N_7604,N_4884,N_5972);
or U7605 (N_7605,N_5264,N_3834);
nand U7606 (N_7606,N_3853,N_5865);
or U7607 (N_7607,N_4732,N_3980);
and U7608 (N_7608,N_4180,N_5342);
and U7609 (N_7609,N_5303,N_5166);
or U7610 (N_7610,N_3016,N_5590);
and U7611 (N_7611,N_4216,N_4699);
xnor U7612 (N_7612,N_5993,N_3537);
xor U7613 (N_7613,N_3695,N_4615);
xor U7614 (N_7614,N_3929,N_3607);
or U7615 (N_7615,N_3641,N_4039);
nor U7616 (N_7616,N_3038,N_4319);
and U7617 (N_7617,N_3589,N_5553);
or U7618 (N_7618,N_5741,N_5963);
and U7619 (N_7619,N_4672,N_3521);
nand U7620 (N_7620,N_5861,N_3062);
and U7621 (N_7621,N_5472,N_4211);
nand U7622 (N_7622,N_4685,N_3428);
nor U7623 (N_7623,N_4283,N_4230);
xor U7624 (N_7624,N_5037,N_3631);
and U7625 (N_7625,N_5449,N_5204);
nand U7626 (N_7626,N_5408,N_5230);
xnor U7627 (N_7627,N_5125,N_5070);
nand U7628 (N_7628,N_4582,N_3169);
or U7629 (N_7629,N_3478,N_5719);
nor U7630 (N_7630,N_4765,N_4865);
xnor U7631 (N_7631,N_3994,N_3569);
and U7632 (N_7632,N_3481,N_3135);
nor U7633 (N_7633,N_4223,N_3892);
nand U7634 (N_7634,N_4049,N_5818);
and U7635 (N_7635,N_3747,N_3300);
or U7636 (N_7636,N_5164,N_5085);
nor U7637 (N_7637,N_4277,N_4137);
nand U7638 (N_7638,N_5562,N_4586);
and U7639 (N_7639,N_5909,N_5914);
or U7640 (N_7640,N_3147,N_3103);
nor U7641 (N_7641,N_5588,N_5114);
and U7642 (N_7642,N_5627,N_3326);
or U7643 (N_7643,N_5541,N_3578);
nand U7644 (N_7644,N_4347,N_3827);
or U7645 (N_7645,N_5898,N_4051);
or U7646 (N_7646,N_3551,N_5460);
and U7647 (N_7647,N_4467,N_3337);
xnor U7648 (N_7648,N_4881,N_4310);
and U7649 (N_7649,N_5658,N_5970);
xnor U7650 (N_7650,N_4316,N_5974);
or U7651 (N_7651,N_4304,N_5486);
nand U7652 (N_7652,N_5932,N_3411);
nand U7653 (N_7653,N_5016,N_5166);
or U7654 (N_7654,N_5941,N_5972);
and U7655 (N_7655,N_3187,N_5153);
nor U7656 (N_7656,N_3536,N_3595);
and U7657 (N_7657,N_4383,N_4818);
and U7658 (N_7658,N_5881,N_3690);
and U7659 (N_7659,N_4122,N_5966);
nand U7660 (N_7660,N_5730,N_4179);
xor U7661 (N_7661,N_3691,N_5678);
nor U7662 (N_7662,N_5359,N_4226);
xor U7663 (N_7663,N_3176,N_3068);
or U7664 (N_7664,N_5117,N_5758);
nor U7665 (N_7665,N_3314,N_4545);
or U7666 (N_7666,N_5876,N_3900);
xnor U7667 (N_7667,N_5252,N_4360);
nand U7668 (N_7668,N_5681,N_4624);
or U7669 (N_7669,N_4791,N_3878);
xor U7670 (N_7670,N_3500,N_5278);
nand U7671 (N_7671,N_5599,N_5108);
xnor U7672 (N_7672,N_4620,N_3730);
or U7673 (N_7673,N_4137,N_3972);
xor U7674 (N_7674,N_3698,N_4124);
nand U7675 (N_7675,N_4799,N_5048);
nand U7676 (N_7676,N_5369,N_3669);
and U7677 (N_7677,N_5461,N_4309);
xor U7678 (N_7678,N_5346,N_4469);
nor U7679 (N_7679,N_5160,N_4855);
and U7680 (N_7680,N_3788,N_3452);
nor U7681 (N_7681,N_4283,N_5828);
and U7682 (N_7682,N_4594,N_5994);
xor U7683 (N_7683,N_5086,N_3970);
nor U7684 (N_7684,N_5176,N_5325);
xnor U7685 (N_7685,N_3884,N_5571);
or U7686 (N_7686,N_5205,N_3469);
nor U7687 (N_7687,N_5440,N_3332);
and U7688 (N_7688,N_5617,N_3623);
xnor U7689 (N_7689,N_5042,N_5150);
and U7690 (N_7690,N_4171,N_5832);
xor U7691 (N_7691,N_3321,N_5578);
and U7692 (N_7692,N_4450,N_4529);
or U7693 (N_7693,N_3523,N_5229);
nor U7694 (N_7694,N_5340,N_4192);
nand U7695 (N_7695,N_4283,N_3381);
xnor U7696 (N_7696,N_3653,N_4305);
nand U7697 (N_7697,N_4632,N_5946);
and U7698 (N_7698,N_5050,N_5364);
nand U7699 (N_7699,N_4984,N_3873);
nand U7700 (N_7700,N_4719,N_4418);
xor U7701 (N_7701,N_4562,N_5918);
or U7702 (N_7702,N_5014,N_5989);
or U7703 (N_7703,N_5089,N_4957);
or U7704 (N_7704,N_3698,N_3731);
nor U7705 (N_7705,N_4068,N_5377);
or U7706 (N_7706,N_4652,N_4935);
xnor U7707 (N_7707,N_3767,N_5593);
nor U7708 (N_7708,N_4273,N_3120);
nor U7709 (N_7709,N_3087,N_4982);
nand U7710 (N_7710,N_3891,N_5538);
or U7711 (N_7711,N_5885,N_3150);
nor U7712 (N_7712,N_4294,N_5518);
and U7713 (N_7713,N_3324,N_4358);
or U7714 (N_7714,N_4570,N_4566);
nand U7715 (N_7715,N_4145,N_4163);
or U7716 (N_7716,N_5799,N_4181);
xnor U7717 (N_7717,N_4814,N_5498);
or U7718 (N_7718,N_4075,N_3402);
and U7719 (N_7719,N_4245,N_4467);
nor U7720 (N_7720,N_4903,N_3026);
nor U7721 (N_7721,N_3353,N_4078);
nand U7722 (N_7722,N_4969,N_4638);
or U7723 (N_7723,N_3091,N_4526);
and U7724 (N_7724,N_5911,N_3474);
xnor U7725 (N_7725,N_5597,N_4053);
or U7726 (N_7726,N_4505,N_5347);
or U7727 (N_7727,N_5386,N_5816);
nor U7728 (N_7728,N_5774,N_5299);
or U7729 (N_7729,N_5399,N_3782);
nor U7730 (N_7730,N_3130,N_4817);
nor U7731 (N_7731,N_3457,N_4128);
nor U7732 (N_7732,N_4027,N_5987);
nor U7733 (N_7733,N_3548,N_5725);
xor U7734 (N_7734,N_3814,N_5189);
xnor U7735 (N_7735,N_5149,N_4070);
and U7736 (N_7736,N_4857,N_5766);
nor U7737 (N_7737,N_4957,N_4289);
or U7738 (N_7738,N_4613,N_3739);
nand U7739 (N_7739,N_3430,N_5845);
xor U7740 (N_7740,N_3770,N_5319);
or U7741 (N_7741,N_5329,N_5613);
nor U7742 (N_7742,N_5254,N_4004);
nand U7743 (N_7743,N_4602,N_3360);
xnor U7744 (N_7744,N_3437,N_3471);
or U7745 (N_7745,N_4996,N_3402);
xor U7746 (N_7746,N_3410,N_3307);
and U7747 (N_7747,N_4217,N_5046);
xnor U7748 (N_7748,N_3019,N_5077);
and U7749 (N_7749,N_3299,N_5275);
or U7750 (N_7750,N_3200,N_3862);
xnor U7751 (N_7751,N_4551,N_3734);
nand U7752 (N_7752,N_4680,N_4582);
nor U7753 (N_7753,N_5428,N_3001);
nand U7754 (N_7754,N_5218,N_3423);
nand U7755 (N_7755,N_4203,N_5158);
xnor U7756 (N_7756,N_5951,N_3537);
and U7757 (N_7757,N_4873,N_4916);
xor U7758 (N_7758,N_3794,N_5621);
xnor U7759 (N_7759,N_5581,N_4677);
nand U7760 (N_7760,N_4733,N_3862);
or U7761 (N_7761,N_4650,N_4976);
or U7762 (N_7762,N_3985,N_5443);
xor U7763 (N_7763,N_3287,N_4596);
xnor U7764 (N_7764,N_4512,N_3651);
nor U7765 (N_7765,N_4661,N_3404);
xnor U7766 (N_7766,N_3409,N_3534);
xnor U7767 (N_7767,N_5806,N_4255);
nand U7768 (N_7768,N_4405,N_4100);
nor U7769 (N_7769,N_5255,N_3740);
nor U7770 (N_7770,N_3658,N_5382);
and U7771 (N_7771,N_3438,N_3904);
or U7772 (N_7772,N_5693,N_5678);
or U7773 (N_7773,N_5686,N_3288);
or U7774 (N_7774,N_3727,N_4569);
xor U7775 (N_7775,N_5000,N_3871);
or U7776 (N_7776,N_4981,N_5818);
or U7777 (N_7777,N_5259,N_3264);
and U7778 (N_7778,N_3237,N_5401);
xor U7779 (N_7779,N_4607,N_4902);
xnor U7780 (N_7780,N_4991,N_3820);
nor U7781 (N_7781,N_4709,N_5568);
and U7782 (N_7782,N_4614,N_5894);
and U7783 (N_7783,N_3501,N_5347);
and U7784 (N_7784,N_4281,N_4048);
nor U7785 (N_7785,N_5957,N_5396);
xnor U7786 (N_7786,N_3096,N_5996);
nor U7787 (N_7787,N_3238,N_3222);
nor U7788 (N_7788,N_3824,N_5010);
or U7789 (N_7789,N_3899,N_5070);
nor U7790 (N_7790,N_3950,N_5854);
or U7791 (N_7791,N_5581,N_5550);
or U7792 (N_7792,N_4053,N_3265);
or U7793 (N_7793,N_5995,N_3374);
and U7794 (N_7794,N_3914,N_3302);
nor U7795 (N_7795,N_3545,N_5500);
nor U7796 (N_7796,N_5422,N_3451);
or U7797 (N_7797,N_4740,N_4462);
or U7798 (N_7798,N_3087,N_5855);
or U7799 (N_7799,N_3426,N_5172);
nor U7800 (N_7800,N_4679,N_4782);
xnor U7801 (N_7801,N_4911,N_5553);
or U7802 (N_7802,N_3113,N_4434);
nand U7803 (N_7803,N_5987,N_5106);
nand U7804 (N_7804,N_5145,N_3528);
nor U7805 (N_7805,N_5217,N_4756);
xor U7806 (N_7806,N_3507,N_5117);
xor U7807 (N_7807,N_5572,N_4918);
and U7808 (N_7808,N_5676,N_4201);
nand U7809 (N_7809,N_3348,N_4517);
nand U7810 (N_7810,N_3253,N_3262);
xnor U7811 (N_7811,N_5701,N_5790);
xor U7812 (N_7812,N_3040,N_4013);
xnor U7813 (N_7813,N_3798,N_5816);
xnor U7814 (N_7814,N_5259,N_4142);
and U7815 (N_7815,N_5310,N_4625);
nor U7816 (N_7816,N_4377,N_5941);
nor U7817 (N_7817,N_5062,N_3555);
nand U7818 (N_7818,N_5836,N_5298);
nor U7819 (N_7819,N_5976,N_4759);
and U7820 (N_7820,N_3884,N_3888);
nor U7821 (N_7821,N_3270,N_3721);
or U7822 (N_7822,N_5644,N_3112);
nand U7823 (N_7823,N_4488,N_4603);
or U7824 (N_7824,N_3758,N_3914);
and U7825 (N_7825,N_4934,N_3589);
xor U7826 (N_7826,N_4559,N_4530);
xnor U7827 (N_7827,N_5977,N_4273);
nor U7828 (N_7828,N_5080,N_4334);
and U7829 (N_7829,N_5368,N_3520);
nor U7830 (N_7830,N_5379,N_3068);
nor U7831 (N_7831,N_5159,N_5706);
or U7832 (N_7832,N_4187,N_3622);
xnor U7833 (N_7833,N_3725,N_4430);
xnor U7834 (N_7834,N_5217,N_4559);
nor U7835 (N_7835,N_5557,N_4082);
nand U7836 (N_7836,N_4408,N_5682);
nor U7837 (N_7837,N_5463,N_3566);
and U7838 (N_7838,N_3162,N_5609);
or U7839 (N_7839,N_5243,N_5080);
nand U7840 (N_7840,N_4783,N_5791);
or U7841 (N_7841,N_5567,N_4619);
nand U7842 (N_7842,N_3727,N_4462);
nor U7843 (N_7843,N_5376,N_3532);
nand U7844 (N_7844,N_4011,N_3805);
nand U7845 (N_7845,N_3927,N_5834);
nor U7846 (N_7846,N_4181,N_4468);
nand U7847 (N_7847,N_3466,N_4405);
or U7848 (N_7848,N_4965,N_5617);
and U7849 (N_7849,N_4590,N_5948);
nand U7850 (N_7850,N_3023,N_3970);
and U7851 (N_7851,N_4793,N_3441);
xor U7852 (N_7852,N_3993,N_4773);
nand U7853 (N_7853,N_4154,N_3215);
xor U7854 (N_7854,N_3594,N_3515);
and U7855 (N_7855,N_5845,N_5574);
nand U7856 (N_7856,N_4748,N_4635);
nor U7857 (N_7857,N_5042,N_4537);
and U7858 (N_7858,N_3100,N_3003);
nand U7859 (N_7859,N_4118,N_5554);
nand U7860 (N_7860,N_4142,N_3712);
nor U7861 (N_7861,N_5019,N_4780);
or U7862 (N_7862,N_4084,N_5628);
nor U7863 (N_7863,N_5016,N_4709);
nor U7864 (N_7864,N_3489,N_5455);
nand U7865 (N_7865,N_4822,N_5224);
and U7866 (N_7866,N_3313,N_4208);
nor U7867 (N_7867,N_4207,N_4656);
or U7868 (N_7868,N_4111,N_5129);
and U7869 (N_7869,N_5594,N_4219);
or U7870 (N_7870,N_3577,N_5297);
nand U7871 (N_7871,N_3923,N_5139);
and U7872 (N_7872,N_3870,N_4096);
or U7873 (N_7873,N_5609,N_5713);
or U7874 (N_7874,N_3751,N_4936);
nand U7875 (N_7875,N_3202,N_3929);
and U7876 (N_7876,N_4804,N_4096);
and U7877 (N_7877,N_4980,N_3552);
or U7878 (N_7878,N_5185,N_4746);
nor U7879 (N_7879,N_5717,N_4464);
and U7880 (N_7880,N_4096,N_4150);
nor U7881 (N_7881,N_5562,N_3760);
or U7882 (N_7882,N_4823,N_5605);
or U7883 (N_7883,N_3526,N_4532);
and U7884 (N_7884,N_5370,N_5462);
or U7885 (N_7885,N_3703,N_3362);
and U7886 (N_7886,N_4857,N_5239);
xnor U7887 (N_7887,N_4999,N_4451);
xnor U7888 (N_7888,N_5338,N_5963);
nand U7889 (N_7889,N_3905,N_4079);
nor U7890 (N_7890,N_5308,N_4591);
xnor U7891 (N_7891,N_3772,N_3352);
xnor U7892 (N_7892,N_3465,N_3525);
and U7893 (N_7893,N_4648,N_4664);
and U7894 (N_7894,N_4028,N_4725);
xnor U7895 (N_7895,N_3603,N_3872);
xor U7896 (N_7896,N_4803,N_3719);
xor U7897 (N_7897,N_4591,N_5581);
nor U7898 (N_7898,N_4071,N_5062);
and U7899 (N_7899,N_3983,N_5878);
xor U7900 (N_7900,N_3317,N_5128);
and U7901 (N_7901,N_4193,N_3685);
nand U7902 (N_7902,N_3793,N_5206);
and U7903 (N_7903,N_5047,N_4344);
nand U7904 (N_7904,N_4554,N_3935);
xnor U7905 (N_7905,N_4720,N_3503);
xnor U7906 (N_7906,N_5413,N_4832);
or U7907 (N_7907,N_5563,N_5140);
nor U7908 (N_7908,N_4941,N_5614);
xnor U7909 (N_7909,N_5593,N_5312);
and U7910 (N_7910,N_5831,N_5851);
nor U7911 (N_7911,N_4416,N_5789);
or U7912 (N_7912,N_4646,N_3246);
and U7913 (N_7913,N_3562,N_5284);
and U7914 (N_7914,N_4217,N_4040);
and U7915 (N_7915,N_3444,N_5231);
xnor U7916 (N_7916,N_3897,N_5897);
nand U7917 (N_7917,N_3057,N_5706);
xor U7918 (N_7918,N_5376,N_3413);
nor U7919 (N_7919,N_5467,N_5313);
and U7920 (N_7920,N_4214,N_4175);
nor U7921 (N_7921,N_5159,N_3923);
xnor U7922 (N_7922,N_5213,N_4324);
or U7923 (N_7923,N_4212,N_3060);
or U7924 (N_7924,N_5927,N_5206);
nor U7925 (N_7925,N_4652,N_3614);
or U7926 (N_7926,N_5775,N_3423);
or U7927 (N_7927,N_4271,N_3910);
nand U7928 (N_7928,N_4179,N_5391);
and U7929 (N_7929,N_4998,N_3212);
nand U7930 (N_7930,N_3283,N_3265);
and U7931 (N_7931,N_3015,N_4117);
nand U7932 (N_7932,N_4079,N_5265);
xnor U7933 (N_7933,N_5385,N_3207);
xnor U7934 (N_7934,N_5674,N_3020);
nand U7935 (N_7935,N_5010,N_4129);
nand U7936 (N_7936,N_3039,N_5543);
xnor U7937 (N_7937,N_5822,N_4953);
and U7938 (N_7938,N_4284,N_5025);
xnor U7939 (N_7939,N_4843,N_3067);
nor U7940 (N_7940,N_4769,N_5302);
and U7941 (N_7941,N_3593,N_4488);
or U7942 (N_7942,N_4494,N_5242);
or U7943 (N_7943,N_4604,N_3310);
nand U7944 (N_7944,N_4215,N_5082);
and U7945 (N_7945,N_4043,N_3505);
and U7946 (N_7946,N_4033,N_4755);
or U7947 (N_7947,N_5185,N_5680);
nor U7948 (N_7948,N_3813,N_5281);
and U7949 (N_7949,N_3330,N_3562);
and U7950 (N_7950,N_3288,N_4007);
or U7951 (N_7951,N_4033,N_3333);
nand U7952 (N_7952,N_4505,N_5628);
and U7953 (N_7953,N_5636,N_4515);
and U7954 (N_7954,N_5819,N_5705);
or U7955 (N_7955,N_4895,N_3279);
or U7956 (N_7956,N_4606,N_3271);
nor U7957 (N_7957,N_5405,N_3336);
xor U7958 (N_7958,N_3631,N_4548);
xnor U7959 (N_7959,N_3825,N_3083);
nand U7960 (N_7960,N_3658,N_3534);
and U7961 (N_7961,N_4794,N_5319);
xnor U7962 (N_7962,N_5122,N_3166);
and U7963 (N_7963,N_4373,N_5011);
nor U7964 (N_7964,N_3007,N_4615);
nand U7965 (N_7965,N_3454,N_3122);
nand U7966 (N_7966,N_4808,N_4656);
or U7967 (N_7967,N_5475,N_3676);
and U7968 (N_7968,N_4600,N_4981);
xnor U7969 (N_7969,N_5610,N_5883);
and U7970 (N_7970,N_5840,N_5023);
nor U7971 (N_7971,N_5744,N_3812);
and U7972 (N_7972,N_4329,N_5002);
nand U7973 (N_7973,N_5059,N_3964);
and U7974 (N_7974,N_5282,N_3097);
or U7975 (N_7975,N_5940,N_3352);
xnor U7976 (N_7976,N_5630,N_4915);
or U7977 (N_7977,N_4046,N_3411);
xor U7978 (N_7978,N_3614,N_5927);
nand U7979 (N_7979,N_5528,N_5831);
and U7980 (N_7980,N_4689,N_5245);
nor U7981 (N_7981,N_3878,N_5057);
and U7982 (N_7982,N_3876,N_3108);
xor U7983 (N_7983,N_4733,N_3042);
or U7984 (N_7984,N_4376,N_4950);
nor U7985 (N_7985,N_5751,N_4760);
nand U7986 (N_7986,N_4193,N_4009);
nand U7987 (N_7987,N_5511,N_3743);
and U7988 (N_7988,N_4052,N_3924);
or U7989 (N_7989,N_5694,N_5793);
and U7990 (N_7990,N_5875,N_4009);
nand U7991 (N_7991,N_3126,N_3268);
or U7992 (N_7992,N_4742,N_3648);
and U7993 (N_7993,N_4872,N_5638);
nor U7994 (N_7994,N_3239,N_4015);
xnor U7995 (N_7995,N_3822,N_3901);
nor U7996 (N_7996,N_4861,N_4001);
nor U7997 (N_7997,N_5547,N_5832);
xor U7998 (N_7998,N_5715,N_3826);
or U7999 (N_7999,N_5439,N_3085);
nor U8000 (N_8000,N_5568,N_4407);
nor U8001 (N_8001,N_4708,N_3756);
or U8002 (N_8002,N_3480,N_4809);
and U8003 (N_8003,N_3879,N_4508);
and U8004 (N_8004,N_5688,N_5990);
nor U8005 (N_8005,N_4721,N_4909);
and U8006 (N_8006,N_3514,N_3226);
nand U8007 (N_8007,N_5180,N_3042);
and U8008 (N_8008,N_4218,N_3053);
nor U8009 (N_8009,N_5659,N_5351);
xnor U8010 (N_8010,N_5005,N_4229);
and U8011 (N_8011,N_4338,N_5676);
and U8012 (N_8012,N_3139,N_5114);
xnor U8013 (N_8013,N_4783,N_3573);
or U8014 (N_8014,N_5837,N_3235);
or U8015 (N_8015,N_5926,N_5095);
or U8016 (N_8016,N_3302,N_4786);
xor U8017 (N_8017,N_4531,N_5789);
xnor U8018 (N_8018,N_4312,N_5631);
and U8019 (N_8019,N_5352,N_5563);
or U8020 (N_8020,N_3456,N_4735);
nor U8021 (N_8021,N_3144,N_3440);
nor U8022 (N_8022,N_4558,N_5578);
or U8023 (N_8023,N_5866,N_5765);
xnor U8024 (N_8024,N_4911,N_4043);
xnor U8025 (N_8025,N_3036,N_4527);
or U8026 (N_8026,N_4548,N_4127);
and U8027 (N_8027,N_5273,N_5784);
nand U8028 (N_8028,N_3794,N_3252);
and U8029 (N_8029,N_4580,N_4914);
nor U8030 (N_8030,N_3029,N_5716);
and U8031 (N_8031,N_4233,N_5806);
xnor U8032 (N_8032,N_5151,N_3723);
or U8033 (N_8033,N_5859,N_3427);
or U8034 (N_8034,N_3446,N_3063);
nand U8035 (N_8035,N_4288,N_4900);
nor U8036 (N_8036,N_4437,N_3851);
or U8037 (N_8037,N_4074,N_5137);
and U8038 (N_8038,N_4354,N_3978);
or U8039 (N_8039,N_4602,N_4658);
nand U8040 (N_8040,N_5854,N_5883);
or U8041 (N_8041,N_4149,N_3076);
nor U8042 (N_8042,N_3720,N_3070);
or U8043 (N_8043,N_5521,N_5821);
nor U8044 (N_8044,N_5896,N_4628);
or U8045 (N_8045,N_4848,N_4283);
nor U8046 (N_8046,N_4362,N_3017);
xor U8047 (N_8047,N_5511,N_5555);
and U8048 (N_8048,N_5122,N_4447);
xor U8049 (N_8049,N_4353,N_4392);
or U8050 (N_8050,N_4439,N_3322);
or U8051 (N_8051,N_5583,N_3787);
nand U8052 (N_8052,N_3292,N_5848);
or U8053 (N_8053,N_4250,N_5099);
nand U8054 (N_8054,N_3743,N_4163);
nor U8055 (N_8055,N_5514,N_5701);
and U8056 (N_8056,N_5084,N_4327);
or U8057 (N_8057,N_5830,N_3005);
or U8058 (N_8058,N_5257,N_5967);
nand U8059 (N_8059,N_4806,N_3783);
or U8060 (N_8060,N_4875,N_5557);
nand U8061 (N_8061,N_4955,N_5765);
or U8062 (N_8062,N_4472,N_4881);
nor U8063 (N_8063,N_5376,N_3816);
or U8064 (N_8064,N_5833,N_5146);
xnor U8065 (N_8065,N_5535,N_4183);
and U8066 (N_8066,N_3422,N_3000);
and U8067 (N_8067,N_3457,N_4471);
nand U8068 (N_8068,N_5838,N_4053);
xor U8069 (N_8069,N_4048,N_3428);
or U8070 (N_8070,N_4370,N_3392);
or U8071 (N_8071,N_3128,N_3793);
or U8072 (N_8072,N_3991,N_3027);
xor U8073 (N_8073,N_3112,N_4769);
xnor U8074 (N_8074,N_5996,N_4234);
nand U8075 (N_8075,N_4320,N_5546);
and U8076 (N_8076,N_3823,N_4244);
nand U8077 (N_8077,N_5899,N_4214);
nand U8078 (N_8078,N_5177,N_3987);
and U8079 (N_8079,N_3368,N_5739);
and U8080 (N_8080,N_4470,N_4016);
nor U8081 (N_8081,N_4023,N_3210);
nand U8082 (N_8082,N_4871,N_3498);
and U8083 (N_8083,N_3730,N_3133);
or U8084 (N_8084,N_5545,N_3100);
or U8085 (N_8085,N_3016,N_5585);
nor U8086 (N_8086,N_5067,N_3351);
nand U8087 (N_8087,N_3581,N_4605);
nor U8088 (N_8088,N_5331,N_3174);
or U8089 (N_8089,N_3963,N_3711);
xor U8090 (N_8090,N_4773,N_3314);
or U8091 (N_8091,N_4966,N_3277);
xor U8092 (N_8092,N_3222,N_4814);
or U8093 (N_8093,N_4176,N_4423);
and U8094 (N_8094,N_3804,N_4466);
and U8095 (N_8095,N_4027,N_4881);
and U8096 (N_8096,N_4558,N_4148);
and U8097 (N_8097,N_4125,N_5333);
and U8098 (N_8098,N_5169,N_3118);
and U8099 (N_8099,N_5799,N_5433);
nor U8100 (N_8100,N_5276,N_3621);
or U8101 (N_8101,N_3403,N_3817);
xor U8102 (N_8102,N_4803,N_5560);
xnor U8103 (N_8103,N_4366,N_5044);
xor U8104 (N_8104,N_3537,N_3701);
nand U8105 (N_8105,N_5646,N_3045);
xor U8106 (N_8106,N_4849,N_4287);
or U8107 (N_8107,N_3996,N_4895);
or U8108 (N_8108,N_3421,N_3243);
nand U8109 (N_8109,N_5361,N_5509);
and U8110 (N_8110,N_4479,N_4023);
nor U8111 (N_8111,N_4831,N_5466);
and U8112 (N_8112,N_4637,N_3448);
nor U8113 (N_8113,N_4662,N_4230);
and U8114 (N_8114,N_5537,N_5148);
nand U8115 (N_8115,N_4826,N_3599);
nand U8116 (N_8116,N_3362,N_4476);
nor U8117 (N_8117,N_3924,N_5328);
nor U8118 (N_8118,N_5006,N_4884);
and U8119 (N_8119,N_3667,N_5216);
nand U8120 (N_8120,N_3352,N_3221);
and U8121 (N_8121,N_3540,N_4031);
nor U8122 (N_8122,N_3832,N_3665);
nand U8123 (N_8123,N_5257,N_5175);
xor U8124 (N_8124,N_5195,N_4101);
or U8125 (N_8125,N_3179,N_4471);
and U8126 (N_8126,N_5472,N_4735);
nand U8127 (N_8127,N_4190,N_4353);
or U8128 (N_8128,N_5132,N_4143);
nor U8129 (N_8129,N_5672,N_4055);
and U8130 (N_8130,N_4499,N_3402);
and U8131 (N_8131,N_5633,N_4855);
nand U8132 (N_8132,N_5666,N_5993);
nand U8133 (N_8133,N_3616,N_4789);
nand U8134 (N_8134,N_5270,N_4913);
xor U8135 (N_8135,N_4336,N_5498);
and U8136 (N_8136,N_5346,N_3459);
or U8137 (N_8137,N_3287,N_3121);
nor U8138 (N_8138,N_5784,N_5020);
nand U8139 (N_8139,N_3189,N_5909);
or U8140 (N_8140,N_4950,N_4537);
xor U8141 (N_8141,N_4820,N_4634);
nor U8142 (N_8142,N_3103,N_4910);
or U8143 (N_8143,N_5504,N_4713);
and U8144 (N_8144,N_3353,N_4215);
nor U8145 (N_8145,N_3098,N_5092);
nor U8146 (N_8146,N_3685,N_4240);
or U8147 (N_8147,N_3604,N_4065);
and U8148 (N_8148,N_5954,N_3966);
xnor U8149 (N_8149,N_3864,N_5674);
or U8150 (N_8150,N_3437,N_4503);
xnor U8151 (N_8151,N_3016,N_5000);
and U8152 (N_8152,N_5240,N_3669);
and U8153 (N_8153,N_5029,N_3563);
xnor U8154 (N_8154,N_4789,N_5852);
and U8155 (N_8155,N_3679,N_3708);
or U8156 (N_8156,N_5959,N_5140);
nand U8157 (N_8157,N_4154,N_3199);
nand U8158 (N_8158,N_3800,N_4783);
nand U8159 (N_8159,N_3193,N_5038);
or U8160 (N_8160,N_5555,N_5785);
or U8161 (N_8161,N_5131,N_5228);
xor U8162 (N_8162,N_5209,N_3909);
or U8163 (N_8163,N_4778,N_5491);
nand U8164 (N_8164,N_4560,N_3383);
or U8165 (N_8165,N_3776,N_3352);
nand U8166 (N_8166,N_3694,N_3671);
xnor U8167 (N_8167,N_3243,N_5805);
nor U8168 (N_8168,N_5955,N_3227);
or U8169 (N_8169,N_3392,N_5370);
xnor U8170 (N_8170,N_4144,N_5538);
nand U8171 (N_8171,N_3073,N_4460);
nor U8172 (N_8172,N_5799,N_5497);
nand U8173 (N_8173,N_4665,N_4950);
and U8174 (N_8174,N_5562,N_4416);
nor U8175 (N_8175,N_4537,N_3158);
xor U8176 (N_8176,N_4342,N_4633);
xor U8177 (N_8177,N_5346,N_5848);
nand U8178 (N_8178,N_3376,N_5421);
and U8179 (N_8179,N_5213,N_4357);
and U8180 (N_8180,N_5690,N_5356);
or U8181 (N_8181,N_5488,N_5037);
xnor U8182 (N_8182,N_4008,N_4128);
nor U8183 (N_8183,N_4032,N_3234);
xnor U8184 (N_8184,N_5858,N_3361);
xor U8185 (N_8185,N_4971,N_5191);
nand U8186 (N_8186,N_5080,N_3560);
nand U8187 (N_8187,N_5900,N_4645);
or U8188 (N_8188,N_3287,N_5503);
xor U8189 (N_8189,N_5375,N_5285);
and U8190 (N_8190,N_5205,N_5169);
nor U8191 (N_8191,N_4994,N_5475);
and U8192 (N_8192,N_4767,N_4262);
and U8193 (N_8193,N_4816,N_3494);
or U8194 (N_8194,N_5213,N_3077);
nand U8195 (N_8195,N_5091,N_4881);
or U8196 (N_8196,N_5841,N_4881);
nor U8197 (N_8197,N_5687,N_3209);
xor U8198 (N_8198,N_5889,N_5960);
nor U8199 (N_8199,N_5380,N_5408);
xnor U8200 (N_8200,N_5854,N_3476);
or U8201 (N_8201,N_5182,N_4362);
nand U8202 (N_8202,N_5453,N_5056);
xnor U8203 (N_8203,N_5147,N_3838);
xnor U8204 (N_8204,N_3174,N_5850);
nor U8205 (N_8205,N_3567,N_3510);
and U8206 (N_8206,N_5034,N_3325);
and U8207 (N_8207,N_4467,N_5995);
nand U8208 (N_8208,N_5474,N_5532);
xor U8209 (N_8209,N_4756,N_4367);
xor U8210 (N_8210,N_3528,N_3654);
xor U8211 (N_8211,N_3438,N_5489);
or U8212 (N_8212,N_5117,N_4307);
xor U8213 (N_8213,N_3202,N_5414);
and U8214 (N_8214,N_3656,N_3635);
nor U8215 (N_8215,N_5209,N_4233);
and U8216 (N_8216,N_3338,N_5114);
nor U8217 (N_8217,N_3828,N_4160);
or U8218 (N_8218,N_4256,N_5527);
xnor U8219 (N_8219,N_3694,N_3836);
nor U8220 (N_8220,N_3355,N_5332);
or U8221 (N_8221,N_5772,N_5759);
xnor U8222 (N_8222,N_5860,N_5349);
or U8223 (N_8223,N_3751,N_3178);
nand U8224 (N_8224,N_5997,N_3526);
nand U8225 (N_8225,N_3341,N_3754);
nor U8226 (N_8226,N_5622,N_3973);
nand U8227 (N_8227,N_4811,N_5478);
nand U8228 (N_8228,N_3305,N_4204);
or U8229 (N_8229,N_5610,N_3828);
and U8230 (N_8230,N_3996,N_5695);
nor U8231 (N_8231,N_3718,N_3738);
nor U8232 (N_8232,N_4875,N_5990);
xor U8233 (N_8233,N_3608,N_4484);
nand U8234 (N_8234,N_4047,N_5901);
nor U8235 (N_8235,N_5990,N_3337);
and U8236 (N_8236,N_5818,N_3699);
xor U8237 (N_8237,N_4730,N_4573);
and U8238 (N_8238,N_5855,N_4925);
xnor U8239 (N_8239,N_5780,N_3376);
and U8240 (N_8240,N_5612,N_5087);
nor U8241 (N_8241,N_4357,N_4609);
or U8242 (N_8242,N_3308,N_4507);
nand U8243 (N_8243,N_4662,N_3507);
xor U8244 (N_8244,N_5010,N_5194);
xnor U8245 (N_8245,N_5763,N_4720);
or U8246 (N_8246,N_4269,N_5793);
or U8247 (N_8247,N_4748,N_4031);
nand U8248 (N_8248,N_5593,N_4791);
or U8249 (N_8249,N_4478,N_4254);
nand U8250 (N_8250,N_3541,N_4692);
nand U8251 (N_8251,N_3962,N_4081);
and U8252 (N_8252,N_3895,N_3534);
and U8253 (N_8253,N_5114,N_4007);
xnor U8254 (N_8254,N_3172,N_3814);
nand U8255 (N_8255,N_4455,N_5020);
or U8256 (N_8256,N_4565,N_5550);
or U8257 (N_8257,N_5429,N_5495);
nor U8258 (N_8258,N_4802,N_4304);
or U8259 (N_8259,N_3882,N_4073);
nand U8260 (N_8260,N_3073,N_3636);
xnor U8261 (N_8261,N_3469,N_5891);
xor U8262 (N_8262,N_3798,N_4176);
or U8263 (N_8263,N_4540,N_3781);
nand U8264 (N_8264,N_3609,N_3031);
xnor U8265 (N_8265,N_3773,N_3467);
or U8266 (N_8266,N_3546,N_3211);
nor U8267 (N_8267,N_3047,N_4083);
nor U8268 (N_8268,N_3743,N_3390);
nand U8269 (N_8269,N_5050,N_4109);
and U8270 (N_8270,N_5023,N_5709);
xor U8271 (N_8271,N_4740,N_5382);
nand U8272 (N_8272,N_3720,N_4485);
nor U8273 (N_8273,N_4357,N_4439);
and U8274 (N_8274,N_3760,N_4787);
or U8275 (N_8275,N_4891,N_5639);
and U8276 (N_8276,N_5296,N_3092);
or U8277 (N_8277,N_5356,N_5782);
xnor U8278 (N_8278,N_3152,N_5442);
nor U8279 (N_8279,N_4166,N_4833);
nand U8280 (N_8280,N_3563,N_3701);
xor U8281 (N_8281,N_5458,N_5988);
nand U8282 (N_8282,N_4704,N_3914);
or U8283 (N_8283,N_3855,N_3829);
xor U8284 (N_8284,N_4851,N_5972);
xor U8285 (N_8285,N_4541,N_5828);
nor U8286 (N_8286,N_4187,N_4907);
nor U8287 (N_8287,N_4146,N_4516);
nand U8288 (N_8288,N_5290,N_3849);
xor U8289 (N_8289,N_3852,N_4116);
or U8290 (N_8290,N_3382,N_3021);
nand U8291 (N_8291,N_5969,N_3883);
xnor U8292 (N_8292,N_3666,N_4597);
nor U8293 (N_8293,N_5034,N_5324);
xnor U8294 (N_8294,N_3533,N_5241);
nor U8295 (N_8295,N_5145,N_4112);
and U8296 (N_8296,N_5615,N_3668);
nor U8297 (N_8297,N_3856,N_5610);
nor U8298 (N_8298,N_5363,N_3936);
and U8299 (N_8299,N_3487,N_3288);
or U8300 (N_8300,N_4834,N_3930);
xnor U8301 (N_8301,N_3409,N_5620);
xor U8302 (N_8302,N_3520,N_3528);
xnor U8303 (N_8303,N_3040,N_4107);
nand U8304 (N_8304,N_4092,N_4264);
xor U8305 (N_8305,N_4151,N_3609);
xnor U8306 (N_8306,N_3728,N_3005);
xor U8307 (N_8307,N_3466,N_3245);
and U8308 (N_8308,N_3433,N_3428);
xor U8309 (N_8309,N_3593,N_4253);
nor U8310 (N_8310,N_3761,N_4796);
nor U8311 (N_8311,N_5221,N_5587);
xnor U8312 (N_8312,N_5473,N_3529);
xor U8313 (N_8313,N_5185,N_3427);
nand U8314 (N_8314,N_5832,N_3764);
and U8315 (N_8315,N_5668,N_4561);
xnor U8316 (N_8316,N_3701,N_4903);
and U8317 (N_8317,N_3191,N_4288);
nand U8318 (N_8318,N_5489,N_3283);
and U8319 (N_8319,N_5419,N_5188);
xor U8320 (N_8320,N_5819,N_3194);
nor U8321 (N_8321,N_4722,N_4943);
or U8322 (N_8322,N_3728,N_5670);
nand U8323 (N_8323,N_5930,N_5471);
and U8324 (N_8324,N_3432,N_5685);
xnor U8325 (N_8325,N_3976,N_4682);
nor U8326 (N_8326,N_5554,N_5056);
xor U8327 (N_8327,N_3127,N_5932);
or U8328 (N_8328,N_4616,N_4975);
and U8329 (N_8329,N_5121,N_4814);
and U8330 (N_8330,N_5083,N_3042);
xor U8331 (N_8331,N_5789,N_3041);
and U8332 (N_8332,N_4973,N_4966);
xor U8333 (N_8333,N_5309,N_5765);
and U8334 (N_8334,N_5319,N_4989);
and U8335 (N_8335,N_5375,N_4335);
or U8336 (N_8336,N_4704,N_3381);
nor U8337 (N_8337,N_5880,N_5366);
and U8338 (N_8338,N_5369,N_5576);
xor U8339 (N_8339,N_5708,N_3965);
nor U8340 (N_8340,N_3497,N_3235);
nand U8341 (N_8341,N_4576,N_3077);
nor U8342 (N_8342,N_3885,N_5451);
nor U8343 (N_8343,N_5646,N_3905);
nand U8344 (N_8344,N_5625,N_5800);
nor U8345 (N_8345,N_4346,N_4201);
nand U8346 (N_8346,N_3410,N_4834);
and U8347 (N_8347,N_4011,N_4438);
or U8348 (N_8348,N_3795,N_5595);
xnor U8349 (N_8349,N_4689,N_4232);
and U8350 (N_8350,N_5476,N_4915);
nand U8351 (N_8351,N_5220,N_5438);
or U8352 (N_8352,N_5994,N_4798);
and U8353 (N_8353,N_4351,N_5029);
and U8354 (N_8354,N_5827,N_5007);
xnor U8355 (N_8355,N_5332,N_5673);
and U8356 (N_8356,N_5220,N_4548);
nor U8357 (N_8357,N_4752,N_5758);
and U8358 (N_8358,N_3174,N_3889);
or U8359 (N_8359,N_5607,N_4058);
and U8360 (N_8360,N_3188,N_5800);
and U8361 (N_8361,N_5990,N_3944);
xnor U8362 (N_8362,N_4296,N_5524);
nand U8363 (N_8363,N_4520,N_4423);
nand U8364 (N_8364,N_5785,N_5769);
xor U8365 (N_8365,N_4051,N_3203);
or U8366 (N_8366,N_4611,N_5486);
nor U8367 (N_8367,N_5314,N_3459);
nor U8368 (N_8368,N_3981,N_5142);
and U8369 (N_8369,N_3411,N_4768);
and U8370 (N_8370,N_3345,N_3729);
nand U8371 (N_8371,N_4002,N_3649);
nand U8372 (N_8372,N_5255,N_5414);
xor U8373 (N_8373,N_4020,N_5978);
or U8374 (N_8374,N_4061,N_3543);
and U8375 (N_8375,N_4494,N_3323);
and U8376 (N_8376,N_5764,N_3741);
nor U8377 (N_8377,N_4998,N_5929);
and U8378 (N_8378,N_4635,N_4220);
xor U8379 (N_8379,N_4056,N_4407);
nor U8380 (N_8380,N_3937,N_5032);
nand U8381 (N_8381,N_4180,N_4697);
or U8382 (N_8382,N_5786,N_5482);
and U8383 (N_8383,N_3779,N_5232);
nor U8384 (N_8384,N_4962,N_4531);
nand U8385 (N_8385,N_5477,N_3483);
and U8386 (N_8386,N_5819,N_3518);
xor U8387 (N_8387,N_5612,N_5259);
xnor U8388 (N_8388,N_3582,N_4162);
nand U8389 (N_8389,N_3778,N_5799);
or U8390 (N_8390,N_5194,N_3220);
xnor U8391 (N_8391,N_5206,N_3192);
nand U8392 (N_8392,N_5464,N_4753);
nor U8393 (N_8393,N_5944,N_3079);
or U8394 (N_8394,N_3744,N_4965);
or U8395 (N_8395,N_3639,N_5837);
nor U8396 (N_8396,N_5952,N_4222);
xor U8397 (N_8397,N_4662,N_4774);
nand U8398 (N_8398,N_4796,N_4870);
or U8399 (N_8399,N_5124,N_5959);
xor U8400 (N_8400,N_3068,N_4905);
xnor U8401 (N_8401,N_3635,N_4149);
nor U8402 (N_8402,N_4769,N_3470);
xnor U8403 (N_8403,N_3338,N_4889);
nand U8404 (N_8404,N_5885,N_4500);
or U8405 (N_8405,N_3391,N_4059);
nor U8406 (N_8406,N_3273,N_4980);
nor U8407 (N_8407,N_3534,N_5241);
or U8408 (N_8408,N_4680,N_5672);
or U8409 (N_8409,N_3600,N_5198);
xnor U8410 (N_8410,N_5317,N_4145);
and U8411 (N_8411,N_4456,N_3243);
xor U8412 (N_8412,N_3327,N_5383);
nand U8413 (N_8413,N_3553,N_3470);
and U8414 (N_8414,N_3063,N_5647);
nand U8415 (N_8415,N_4850,N_5908);
and U8416 (N_8416,N_4440,N_4456);
nand U8417 (N_8417,N_3693,N_3388);
nor U8418 (N_8418,N_5140,N_3211);
or U8419 (N_8419,N_5682,N_3771);
and U8420 (N_8420,N_4669,N_3543);
nand U8421 (N_8421,N_3093,N_4097);
nor U8422 (N_8422,N_4201,N_5226);
nand U8423 (N_8423,N_4785,N_5184);
nand U8424 (N_8424,N_4046,N_4486);
nand U8425 (N_8425,N_3072,N_5600);
nand U8426 (N_8426,N_3002,N_5157);
nor U8427 (N_8427,N_4563,N_4213);
nand U8428 (N_8428,N_5576,N_3595);
nand U8429 (N_8429,N_3748,N_4540);
nand U8430 (N_8430,N_5144,N_4979);
or U8431 (N_8431,N_3075,N_3590);
and U8432 (N_8432,N_4712,N_3032);
and U8433 (N_8433,N_3472,N_5597);
nor U8434 (N_8434,N_3027,N_3481);
xnor U8435 (N_8435,N_4563,N_3736);
nand U8436 (N_8436,N_4304,N_5453);
and U8437 (N_8437,N_3071,N_4901);
and U8438 (N_8438,N_4699,N_5176);
or U8439 (N_8439,N_4577,N_4297);
nor U8440 (N_8440,N_4366,N_3698);
nand U8441 (N_8441,N_4324,N_3784);
and U8442 (N_8442,N_3408,N_4734);
or U8443 (N_8443,N_3905,N_5911);
and U8444 (N_8444,N_4307,N_4442);
nand U8445 (N_8445,N_5915,N_3742);
nand U8446 (N_8446,N_4954,N_4765);
and U8447 (N_8447,N_4473,N_4184);
xnor U8448 (N_8448,N_5902,N_4104);
nor U8449 (N_8449,N_5141,N_4612);
or U8450 (N_8450,N_5847,N_3990);
nand U8451 (N_8451,N_5561,N_4375);
or U8452 (N_8452,N_3675,N_4647);
or U8453 (N_8453,N_5085,N_5371);
and U8454 (N_8454,N_4590,N_4224);
and U8455 (N_8455,N_4836,N_5253);
xnor U8456 (N_8456,N_4999,N_5571);
nand U8457 (N_8457,N_3013,N_4999);
and U8458 (N_8458,N_5265,N_5029);
or U8459 (N_8459,N_4648,N_5484);
or U8460 (N_8460,N_5075,N_5439);
xnor U8461 (N_8461,N_3789,N_4535);
nand U8462 (N_8462,N_4803,N_4026);
and U8463 (N_8463,N_5366,N_4989);
and U8464 (N_8464,N_5773,N_5569);
and U8465 (N_8465,N_5904,N_3468);
nand U8466 (N_8466,N_5191,N_5443);
xor U8467 (N_8467,N_5128,N_4884);
nand U8468 (N_8468,N_4858,N_5523);
and U8469 (N_8469,N_3648,N_4239);
nand U8470 (N_8470,N_3119,N_5552);
nor U8471 (N_8471,N_5489,N_3589);
nand U8472 (N_8472,N_3294,N_5080);
xor U8473 (N_8473,N_4468,N_3288);
or U8474 (N_8474,N_5774,N_3192);
and U8475 (N_8475,N_3081,N_3995);
nand U8476 (N_8476,N_5861,N_4645);
nand U8477 (N_8477,N_3580,N_4953);
or U8478 (N_8478,N_5125,N_3928);
and U8479 (N_8479,N_3555,N_3578);
nor U8480 (N_8480,N_3872,N_4359);
and U8481 (N_8481,N_5765,N_3678);
nor U8482 (N_8482,N_5176,N_5842);
or U8483 (N_8483,N_4224,N_4499);
and U8484 (N_8484,N_4564,N_5678);
xor U8485 (N_8485,N_4245,N_3655);
nor U8486 (N_8486,N_4413,N_5582);
or U8487 (N_8487,N_5825,N_4212);
or U8488 (N_8488,N_4095,N_4242);
nor U8489 (N_8489,N_4558,N_5925);
or U8490 (N_8490,N_3391,N_3642);
nor U8491 (N_8491,N_5356,N_3050);
nor U8492 (N_8492,N_5860,N_4961);
nor U8493 (N_8493,N_4956,N_3974);
or U8494 (N_8494,N_4089,N_3539);
xnor U8495 (N_8495,N_5795,N_5355);
nand U8496 (N_8496,N_4727,N_5209);
nand U8497 (N_8497,N_3504,N_3578);
xor U8498 (N_8498,N_5558,N_3934);
or U8499 (N_8499,N_5097,N_4242);
or U8500 (N_8500,N_5545,N_4194);
nand U8501 (N_8501,N_5368,N_4001);
and U8502 (N_8502,N_5583,N_4898);
and U8503 (N_8503,N_5933,N_5323);
nand U8504 (N_8504,N_5009,N_3732);
nand U8505 (N_8505,N_4562,N_5178);
nor U8506 (N_8506,N_5859,N_5867);
nand U8507 (N_8507,N_3565,N_3137);
nand U8508 (N_8508,N_4214,N_3547);
and U8509 (N_8509,N_3101,N_3928);
nand U8510 (N_8510,N_4185,N_5180);
nor U8511 (N_8511,N_5524,N_5185);
or U8512 (N_8512,N_5562,N_3708);
xnor U8513 (N_8513,N_4432,N_5638);
xnor U8514 (N_8514,N_3275,N_5080);
or U8515 (N_8515,N_4574,N_5376);
xor U8516 (N_8516,N_3817,N_5153);
nand U8517 (N_8517,N_4716,N_4972);
xor U8518 (N_8518,N_5666,N_3965);
and U8519 (N_8519,N_4979,N_3611);
nor U8520 (N_8520,N_5535,N_5150);
and U8521 (N_8521,N_4994,N_3694);
or U8522 (N_8522,N_3399,N_4228);
and U8523 (N_8523,N_4462,N_4120);
and U8524 (N_8524,N_4221,N_4774);
nand U8525 (N_8525,N_3404,N_4613);
or U8526 (N_8526,N_5827,N_4431);
xnor U8527 (N_8527,N_3847,N_3267);
and U8528 (N_8528,N_5919,N_5984);
or U8529 (N_8529,N_5722,N_3145);
xor U8530 (N_8530,N_5770,N_3497);
or U8531 (N_8531,N_3448,N_5422);
xor U8532 (N_8532,N_3821,N_5751);
nor U8533 (N_8533,N_5471,N_3727);
or U8534 (N_8534,N_5505,N_4351);
or U8535 (N_8535,N_5684,N_4055);
nor U8536 (N_8536,N_3666,N_4996);
nand U8537 (N_8537,N_4391,N_4578);
or U8538 (N_8538,N_4082,N_5087);
or U8539 (N_8539,N_3802,N_4477);
and U8540 (N_8540,N_5686,N_5768);
and U8541 (N_8541,N_4495,N_3253);
nand U8542 (N_8542,N_3023,N_4777);
nor U8543 (N_8543,N_5100,N_4545);
nand U8544 (N_8544,N_5358,N_3282);
and U8545 (N_8545,N_4901,N_5934);
nor U8546 (N_8546,N_3724,N_4865);
nor U8547 (N_8547,N_3401,N_5430);
or U8548 (N_8548,N_3679,N_4926);
xor U8549 (N_8549,N_5746,N_3479);
xnor U8550 (N_8550,N_3439,N_5050);
or U8551 (N_8551,N_5394,N_3009);
and U8552 (N_8552,N_5981,N_3313);
nand U8553 (N_8553,N_4603,N_5956);
or U8554 (N_8554,N_3102,N_3505);
or U8555 (N_8555,N_4396,N_4507);
nand U8556 (N_8556,N_5163,N_4436);
or U8557 (N_8557,N_3082,N_3079);
and U8558 (N_8558,N_3352,N_4444);
or U8559 (N_8559,N_5160,N_5430);
or U8560 (N_8560,N_4609,N_4912);
nor U8561 (N_8561,N_3116,N_4543);
xnor U8562 (N_8562,N_3389,N_4504);
and U8563 (N_8563,N_4768,N_3315);
nor U8564 (N_8564,N_3005,N_4466);
and U8565 (N_8565,N_4007,N_5144);
nor U8566 (N_8566,N_4755,N_3060);
xor U8567 (N_8567,N_5489,N_3945);
and U8568 (N_8568,N_4457,N_4785);
nor U8569 (N_8569,N_3299,N_3053);
and U8570 (N_8570,N_4731,N_3080);
or U8571 (N_8571,N_5320,N_4555);
nand U8572 (N_8572,N_4123,N_3175);
xnor U8573 (N_8573,N_3332,N_4371);
xor U8574 (N_8574,N_5304,N_3801);
nor U8575 (N_8575,N_5467,N_4884);
nand U8576 (N_8576,N_4726,N_4328);
and U8577 (N_8577,N_4877,N_3924);
or U8578 (N_8578,N_3160,N_5489);
nand U8579 (N_8579,N_4309,N_3939);
nand U8580 (N_8580,N_4983,N_3013);
nor U8581 (N_8581,N_4117,N_3876);
xor U8582 (N_8582,N_4981,N_3942);
nand U8583 (N_8583,N_3814,N_3213);
nand U8584 (N_8584,N_4868,N_4572);
nor U8585 (N_8585,N_4637,N_3936);
nor U8586 (N_8586,N_5746,N_5321);
or U8587 (N_8587,N_3844,N_3233);
nor U8588 (N_8588,N_4279,N_3925);
or U8589 (N_8589,N_4656,N_5819);
or U8590 (N_8590,N_3365,N_3888);
and U8591 (N_8591,N_5330,N_5886);
and U8592 (N_8592,N_3488,N_4273);
xor U8593 (N_8593,N_5396,N_5662);
nor U8594 (N_8594,N_3472,N_4494);
nor U8595 (N_8595,N_4062,N_3238);
xor U8596 (N_8596,N_3143,N_4352);
nand U8597 (N_8597,N_4252,N_3636);
xnor U8598 (N_8598,N_5363,N_3608);
and U8599 (N_8599,N_5731,N_4945);
and U8600 (N_8600,N_4508,N_5532);
xor U8601 (N_8601,N_5594,N_5542);
or U8602 (N_8602,N_4965,N_5951);
or U8603 (N_8603,N_5077,N_3308);
nand U8604 (N_8604,N_3900,N_5623);
or U8605 (N_8605,N_5278,N_5762);
xnor U8606 (N_8606,N_5078,N_4070);
nand U8607 (N_8607,N_3718,N_4333);
nand U8608 (N_8608,N_5249,N_3970);
nand U8609 (N_8609,N_4323,N_3862);
and U8610 (N_8610,N_3703,N_5310);
and U8611 (N_8611,N_3729,N_3538);
nand U8612 (N_8612,N_4261,N_5104);
xor U8613 (N_8613,N_5029,N_4936);
xnor U8614 (N_8614,N_5343,N_5228);
xnor U8615 (N_8615,N_3568,N_5380);
xnor U8616 (N_8616,N_5486,N_3833);
nor U8617 (N_8617,N_5810,N_5513);
xnor U8618 (N_8618,N_5723,N_4047);
and U8619 (N_8619,N_3837,N_4536);
and U8620 (N_8620,N_3839,N_5566);
or U8621 (N_8621,N_5189,N_4391);
nor U8622 (N_8622,N_4537,N_5085);
nand U8623 (N_8623,N_5925,N_3282);
and U8624 (N_8624,N_5768,N_5985);
nor U8625 (N_8625,N_3870,N_5890);
or U8626 (N_8626,N_4151,N_3720);
or U8627 (N_8627,N_3543,N_3219);
nor U8628 (N_8628,N_5848,N_3546);
and U8629 (N_8629,N_4339,N_5809);
nor U8630 (N_8630,N_3484,N_5920);
and U8631 (N_8631,N_4149,N_4713);
xor U8632 (N_8632,N_5008,N_3947);
or U8633 (N_8633,N_3298,N_4662);
or U8634 (N_8634,N_3918,N_4868);
nand U8635 (N_8635,N_4101,N_3449);
xnor U8636 (N_8636,N_4189,N_5697);
xor U8637 (N_8637,N_5978,N_4000);
and U8638 (N_8638,N_5661,N_5939);
and U8639 (N_8639,N_5269,N_3496);
nor U8640 (N_8640,N_5900,N_3947);
nor U8641 (N_8641,N_5756,N_4963);
or U8642 (N_8642,N_4672,N_5651);
nor U8643 (N_8643,N_5226,N_5791);
and U8644 (N_8644,N_3584,N_4154);
nor U8645 (N_8645,N_4297,N_5771);
xnor U8646 (N_8646,N_3833,N_5147);
and U8647 (N_8647,N_5135,N_5192);
xnor U8648 (N_8648,N_4860,N_5007);
or U8649 (N_8649,N_5753,N_5630);
nand U8650 (N_8650,N_5007,N_3553);
nor U8651 (N_8651,N_5880,N_4797);
and U8652 (N_8652,N_3498,N_4657);
and U8653 (N_8653,N_5741,N_4786);
or U8654 (N_8654,N_3294,N_4287);
nor U8655 (N_8655,N_4830,N_4334);
xnor U8656 (N_8656,N_3955,N_5309);
xor U8657 (N_8657,N_5354,N_4402);
or U8658 (N_8658,N_3121,N_3820);
nor U8659 (N_8659,N_4050,N_4164);
and U8660 (N_8660,N_4692,N_5770);
xor U8661 (N_8661,N_3657,N_4791);
xnor U8662 (N_8662,N_4896,N_3177);
nor U8663 (N_8663,N_5310,N_5786);
xnor U8664 (N_8664,N_3932,N_3477);
nor U8665 (N_8665,N_4635,N_5096);
or U8666 (N_8666,N_4489,N_4929);
or U8667 (N_8667,N_4383,N_3753);
or U8668 (N_8668,N_5360,N_5372);
nand U8669 (N_8669,N_3064,N_5694);
nand U8670 (N_8670,N_4268,N_5077);
nand U8671 (N_8671,N_3399,N_4051);
and U8672 (N_8672,N_5182,N_4749);
and U8673 (N_8673,N_4009,N_4760);
nand U8674 (N_8674,N_5046,N_4716);
nand U8675 (N_8675,N_4697,N_5115);
or U8676 (N_8676,N_5777,N_3707);
nor U8677 (N_8677,N_3746,N_4008);
xnor U8678 (N_8678,N_4208,N_3730);
xor U8679 (N_8679,N_4721,N_3717);
or U8680 (N_8680,N_5360,N_5089);
and U8681 (N_8681,N_5381,N_5598);
or U8682 (N_8682,N_3084,N_5140);
and U8683 (N_8683,N_3546,N_5105);
xnor U8684 (N_8684,N_5800,N_3860);
or U8685 (N_8685,N_4718,N_3705);
or U8686 (N_8686,N_4720,N_4311);
or U8687 (N_8687,N_3592,N_4856);
xor U8688 (N_8688,N_4680,N_4452);
nand U8689 (N_8689,N_4106,N_3990);
nand U8690 (N_8690,N_3264,N_4783);
and U8691 (N_8691,N_3433,N_5183);
nand U8692 (N_8692,N_5569,N_4305);
and U8693 (N_8693,N_3814,N_5277);
nand U8694 (N_8694,N_3958,N_3550);
or U8695 (N_8695,N_4826,N_3821);
nand U8696 (N_8696,N_3698,N_3619);
nor U8697 (N_8697,N_4559,N_4892);
nand U8698 (N_8698,N_4111,N_3587);
and U8699 (N_8699,N_3130,N_5518);
nor U8700 (N_8700,N_3494,N_4367);
xnor U8701 (N_8701,N_4623,N_3803);
and U8702 (N_8702,N_3685,N_3086);
or U8703 (N_8703,N_3148,N_4379);
and U8704 (N_8704,N_5131,N_4516);
or U8705 (N_8705,N_5637,N_5896);
or U8706 (N_8706,N_4647,N_5467);
and U8707 (N_8707,N_5627,N_3172);
nor U8708 (N_8708,N_5675,N_5648);
nand U8709 (N_8709,N_5501,N_3952);
or U8710 (N_8710,N_5113,N_4196);
and U8711 (N_8711,N_5697,N_3992);
or U8712 (N_8712,N_5193,N_5470);
nand U8713 (N_8713,N_4536,N_5704);
or U8714 (N_8714,N_5743,N_4178);
and U8715 (N_8715,N_4413,N_5509);
xnor U8716 (N_8716,N_5002,N_3073);
xnor U8717 (N_8717,N_5029,N_3094);
xnor U8718 (N_8718,N_4063,N_4973);
nor U8719 (N_8719,N_3087,N_3449);
and U8720 (N_8720,N_4337,N_3838);
xor U8721 (N_8721,N_4661,N_3169);
or U8722 (N_8722,N_3687,N_3362);
or U8723 (N_8723,N_5235,N_3693);
or U8724 (N_8724,N_5803,N_5928);
or U8725 (N_8725,N_4607,N_5201);
nor U8726 (N_8726,N_5537,N_4644);
nor U8727 (N_8727,N_4408,N_5454);
nand U8728 (N_8728,N_3648,N_5979);
or U8729 (N_8729,N_3876,N_5089);
and U8730 (N_8730,N_3978,N_5910);
or U8731 (N_8731,N_4494,N_5314);
and U8732 (N_8732,N_5975,N_4209);
nand U8733 (N_8733,N_4466,N_4556);
or U8734 (N_8734,N_5999,N_3181);
xor U8735 (N_8735,N_3191,N_5217);
xor U8736 (N_8736,N_3035,N_4946);
xnor U8737 (N_8737,N_4454,N_4840);
nor U8738 (N_8738,N_3627,N_3467);
nor U8739 (N_8739,N_5520,N_4301);
or U8740 (N_8740,N_5412,N_5331);
nor U8741 (N_8741,N_4418,N_5822);
nor U8742 (N_8742,N_3467,N_4921);
nor U8743 (N_8743,N_4396,N_3363);
or U8744 (N_8744,N_3857,N_5291);
nand U8745 (N_8745,N_3921,N_4557);
nor U8746 (N_8746,N_5251,N_4813);
nor U8747 (N_8747,N_4459,N_5148);
nor U8748 (N_8748,N_4493,N_3069);
nor U8749 (N_8749,N_5256,N_3471);
or U8750 (N_8750,N_5688,N_5453);
nand U8751 (N_8751,N_4473,N_5073);
or U8752 (N_8752,N_5209,N_5157);
and U8753 (N_8753,N_3969,N_4195);
nand U8754 (N_8754,N_3740,N_5294);
nand U8755 (N_8755,N_3206,N_3968);
nand U8756 (N_8756,N_4798,N_5405);
xnor U8757 (N_8757,N_3294,N_5948);
nand U8758 (N_8758,N_3965,N_5487);
or U8759 (N_8759,N_3799,N_4051);
nor U8760 (N_8760,N_4459,N_5081);
xor U8761 (N_8761,N_3668,N_4627);
and U8762 (N_8762,N_3726,N_4812);
and U8763 (N_8763,N_4608,N_4200);
or U8764 (N_8764,N_3023,N_5203);
nand U8765 (N_8765,N_3161,N_4652);
and U8766 (N_8766,N_3835,N_5857);
xor U8767 (N_8767,N_3770,N_3925);
nor U8768 (N_8768,N_5873,N_4966);
and U8769 (N_8769,N_4768,N_3088);
nand U8770 (N_8770,N_3982,N_3719);
nand U8771 (N_8771,N_5358,N_5857);
and U8772 (N_8772,N_3793,N_4751);
nand U8773 (N_8773,N_3001,N_5413);
xor U8774 (N_8774,N_3598,N_5995);
and U8775 (N_8775,N_3377,N_5508);
nand U8776 (N_8776,N_5974,N_3895);
and U8777 (N_8777,N_4360,N_4069);
xor U8778 (N_8778,N_5003,N_4820);
and U8779 (N_8779,N_3299,N_4230);
and U8780 (N_8780,N_3674,N_5177);
xor U8781 (N_8781,N_4582,N_5811);
or U8782 (N_8782,N_5515,N_5935);
or U8783 (N_8783,N_4008,N_4553);
or U8784 (N_8784,N_5842,N_3473);
nor U8785 (N_8785,N_4487,N_3434);
nor U8786 (N_8786,N_3564,N_4063);
or U8787 (N_8787,N_3788,N_3224);
and U8788 (N_8788,N_3162,N_4207);
and U8789 (N_8789,N_5859,N_5620);
nand U8790 (N_8790,N_5357,N_4076);
nand U8791 (N_8791,N_5840,N_3405);
or U8792 (N_8792,N_4066,N_3360);
and U8793 (N_8793,N_4969,N_4141);
xor U8794 (N_8794,N_3213,N_5346);
xor U8795 (N_8795,N_3972,N_5389);
nor U8796 (N_8796,N_5078,N_3927);
and U8797 (N_8797,N_4493,N_3124);
xor U8798 (N_8798,N_4351,N_4664);
and U8799 (N_8799,N_3733,N_3347);
nand U8800 (N_8800,N_5507,N_3670);
or U8801 (N_8801,N_4413,N_5889);
xnor U8802 (N_8802,N_5736,N_5471);
or U8803 (N_8803,N_5312,N_5128);
and U8804 (N_8804,N_3816,N_4808);
and U8805 (N_8805,N_4864,N_5158);
xor U8806 (N_8806,N_3099,N_4540);
or U8807 (N_8807,N_5318,N_3736);
xor U8808 (N_8808,N_5307,N_3095);
xnor U8809 (N_8809,N_5809,N_3925);
nand U8810 (N_8810,N_5372,N_4062);
or U8811 (N_8811,N_5449,N_4073);
and U8812 (N_8812,N_5517,N_3674);
and U8813 (N_8813,N_3994,N_5879);
nor U8814 (N_8814,N_3522,N_5356);
or U8815 (N_8815,N_3063,N_3463);
or U8816 (N_8816,N_3850,N_5864);
nor U8817 (N_8817,N_5835,N_5230);
and U8818 (N_8818,N_4316,N_5305);
and U8819 (N_8819,N_3876,N_5494);
and U8820 (N_8820,N_5622,N_4688);
and U8821 (N_8821,N_4544,N_3061);
or U8822 (N_8822,N_3131,N_4331);
and U8823 (N_8823,N_5312,N_5119);
and U8824 (N_8824,N_5020,N_3443);
nor U8825 (N_8825,N_3500,N_4567);
and U8826 (N_8826,N_4808,N_3644);
or U8827 (N_8827,N_3378,N_3926);
nor U8828 (N_8828,N_3181,N_3402);
nor U8829 (N_8829,N_3941,N_4897);
or U8830 (N_8830,N_4927,N_5085);
xnor U8831 (N_8831,N_3202,N_3907);
or U8832 (N_8832,N_4392,N_4563);
xor U8833 (N_8833,N_5541,N_5548);
or U8834 (N_8834,N_3937,N_4478);
or U8835 (N_8835,N_3505,N_4918);
nor U8836 (N_8836,N_4913,N_5946);
xnor U8837 (N_8837,N_5897,N_4639);
or U8838 (N_8838,N_5182,N_3467);
and U8839 (N_8839,N_5622,N_5623);
xor U8840 (N_8840,N_3977,N_5975);
or U8841 (N_8841,N_4132,N_3131);
nor U8842 (N_8842,N_3694,N_5422);
nor U8843 (N_8843,N_3877,N_3916);
xor U8844 (N_8844,N_4465,N_5736);
or U8845 (N_8845,N_4485,N_3101);
and U8846 (N_8846,N_4294,N_5483);
xor U8847 (N_8847,N_4169,N_4068);
or U8848 (N_8848,N_4800,N_3170);
xnor U8849 (N_8849,N_5831,N_5468);
nor U8850 (N_8850,N_4704,N_3772);
and U8851 (N_8851,N_3474,N_3428);
xnor U8852 (N_8852,N_4964,N_4426);
and U8853 (N_8853,N_4509,N_3032);
xor U8854 (N_8854,N_3002,N_4647);
and U8855 (N_8855,N_4874,N_3817);
and U8856 (N_8856,N_4971,N_5551);
or U8857 (N_8857,N_5931,N_3971);
xnor U8858 (N_8858,N_5236,N_5420);
xor U8859 (N_8859,N_5897,N_5901);
xor U8860 (N_8860,N_5284,N_5760);
nand U8861 (N_8861,N_3050,N_5450);
or U8862 (N_8862,N_4827,N_3394);
nor U8863 (N_8863,N_4187,N_4850);
and U8864 (N_8864,N_5966,N_3801);
nor U8865 (N_8865,N_4154,N_5268);
nor U8866 (N_8866,N_3090,N_5116);
and U8867 (N_8867,N_5055,N_4517);
nor U8868 (N_8868,N_5153,N_4329);
nor U8869 (N_8869,N_3264,N_3869);
and U8870 (N_8870,N_5651,N_3888);
or U8871 (N_8871,N_3992,N_3956);
nand U8872 (N_8872,N_4191,N_5382);
nand U8873 (N_8873,N_3166,N_4960);
nand U8874 (N_8874,N_3201,N_3215);
or U8875 (N_8875,N_4725,N_5825);
and U8876 (N_8876,N_5836,N_4388);
xnor U8877 (N_8877,N_5191,N_3384);
nand U8878 (N_8878,N_3968,N_4398);
nand U8879 (N_8879,N_3199,N_5772);
nand U8880 (N_8880,N_3471,N_4544);
or U8881 (N_8881,N_5202,N_4919);
and U8882 (N_8882,N_5288,N_4790);
nand U8883 (N_8883,N_4142,N_3265);
and U8884 (N_8884,N_5323,N_5557);
nor U8885 (N_8885,N_5260,N_3084);
and U8886 (N_8886,N_5742,N_4957);
xor U8887 (N_8887,N_4744,N_3634);
nor U8888 (N_8888,N_3573,N_3470);
xnor U8889 (N_8889,N_5071,N_3462);
or U8890 (N_8890,N_4089,N_5799);
xor U8891 (N_8891,N_5437,N_5113);
xor U8892 (N_8892,N_3942,N_4252);
nor U8893 (N_8893,N_4083,N_4372);
or U8894 (N_8894,N_4537,N_4123);
xnor U8895 (N_8895,N_4668,N_3290);
nand U8896 (N_8896,N_5630,N_5893);
and U8897 (N_8897,N_3000,N_5134);
nor U8898 (N_8898,N_3549,N_4982);
nand U8899 (N_8899,N_3256,N_3142);
nor U8900 (N_8900,N_3862,N_4234);
nand U8901 (N_8901,N_5935,N_3668);
xor U8902 (N_8902,N_3990,N_3177);
and U8903 (N_8903,N_3002,N_3567);
nand U8904 (N_8904,N_4910,N_4817);
nand U8905 (N_8905,N_4257,N_5529);
and U8906 (N_8906,N_5250,N_5382);
nor U8907 (N_8907,N_5234,N_5917);
or U8908 (N_8908,N_3060,N_3326);
or U8909 (N_8909,N_5264,N_3610);
or U8910 (N_8910,N_5522,N_3008);
xor U8911 (N_8911,N_4941,N_3635);
nand U8912 (N_8912,N_3510,N_5910);
nor U8913 (N_8913,N_3384,N_5895);
xnor U8914 (N_8914,N_3032,N_3264);
and U8915 (N_8915,N_4014,N_4328);
nand U8916 (N_8916,N_4748,N_5548);
or U8917 (N_8917,N_3689,N_3925);
nand U8918 (N_8918,N_4820,N_5273);
or U8919 (N_8919,N_3074,N_3425);
or U8920 (N_8920,N_3278,N_4133);
nand U8921 (N_8921,N_5355,N_3463);
xor U8922 (N_8922,N_3799,N_3812);
nand U8923 (N_8923,N_4129,N_3759);
nand U8924 (N_8924,N_3061,N_4205);
nor U8925 (N_8925,N_3574,N_5552);
nor U8926 (N_8926,N_3006,N_4465);
and U8927 (N_8927,N_5052,N_5862);
nand U8928 (N_8928,N_3454,N_4035);
or U8929 (N_8929,N_5917,N_3609);
and U8930 (N_8930,N_5303,N_5835);
nor U8931 (N_8931,N_4760,N_3328);
nor U8932 (N_8932,N_4957,N_4119);
and U8933 (N_8933,N_5288,N_5215);
or U8934 (N_8934,N_3350,N_5370);
or U8935 (N_8935,N_3440,N_4844);
or U8936 (N_8936,N_4421,N_4481);
or U8937 (N_8937,N_4126,N_3116);
and U8938 (N_8938,N_5136,N_3152);
nand U8939 (N_8939,N_5270,N_3097);
nand U8940 (N_8940,N_5346,N_5750);
or U8941 (N_8941,N_4157,N_5759);
nand U8942 (N_8942,N_4814,N_3845);
nand U8943 (N_8943,N_3773,N_3100);
nor U8944 (N_8944,N_4143,N_5195);
nor U8945 (N_8945,N_5621,N_3510);
nor U8946 (N_8946,N_3816,N_4912);
nand U8947 (N_8947,N_4482,N_3936);
and U8948 (N_8948,N_3424,N_4328);
or U8949 (N_8949,N_3997,N_3870);
xor U8950 (N_8950,N_5028,N_4675);
and U8951 (N_8951,N_5661,N_5760);
xor U8952 (N_8952,N_3777,N_5473);
and U8953 (N_8953,N_4267,N_4450);
or U8954 (N_8954,N_5644,N_3165);
xor U8955 (N_8955,N_4633,N_3015);
xnor U8956 (N_8956,N_5353,N_3566);
nor U8957 (N_8957,N_3465,N_4485);
nor U8958 (N_8958,N_3224,N_5482);
or U8959 (N_8959,N_3880,N_4545);
nand U8960 (N_8960,N_4682,N_3119);
nor U8961 (N_8961,N_3020,N_4068);
nor U8962 (N_8962,N_3907,N_5067);
or U8963 (N_8963,N_4305,N_4427);
or U8964 (N_8964,N_5678,N_4946);
and U8965 (N_8965,N_5018,N_3350);
nor U8966 (N_8966,N_4004,N_4034);
nor U8967 (N_8967,N_4513,N_5554);
nor U8968 (N_8968,N_5773,N_3065);
or U8969 (N_8969,N_4753,N_5913);
nand U8970 (N_8970,N_4667,N_3472);
nor U8971 (N_8971,N_4562,N_4111);
xnor U8972 (N_8972,N_4763,N_5943);
xnor U8973 (N_8973,N_5935,N_3834);
nor U8974 (N_8974,N_3392,N_3492);
and U8975 (N_8975,N_3789,N_5480);
or U8976 (N_8976,N_3149,N_5005);
or U8977 (N_8977,N_4230,N_4987);
and U8978 (N_8978,N_3242,N_4373);
nor U8979 (N_8979,N_5953,N_5206);
or U8980 (N_8980,N_4871,N_3796);
and U8981 (N_8981,N_4219,N_5969);
nand U8982 (N_8982,N_5626,N_5814);
xor U8983 (N_8983,N_4352,N_3635);
xor U8984 (N_8984,N_5514,N_5688);
or U8985 (N_8985,N_4459,N_5116);
nand U8986 (N_8986,N_5252,N_5120);
nand U8987 (N_8987,N_5807,N_5707);
xor U8988 (N_8988,N_3087,N_5599);
nor U8989 (N_8989,N_5802,N_5834);
nand U8990 (N_8990,N_5373,N_4868);
nor U8991 (N_8991,N_4353,N_3343);
nor U8992 (N_8992,N_3207,N_3259);
nand U8993 (N_8993,N_5928,N_5793);
nand U8994 (N_8994,N_4797,N_5887);
xnor U8995 (N_8995,N_4984,N_3404);
and U8996 (N_8996,N_4223,N_4739);
nor U8997 (N_8997,N_4645,N_4733);
nor U8998 (N_8998,N_3374,N_5975);
nor U8999 (N_8999,N_3171,N_3147);
or U9000 (N_9000,N_8659,N_8543);
xnor U9001 (N_9001,N_6555,N_6533);
and U9002 (N_9002,N_7515,N_7288);
nand U9003 (N_9003,N_6327,N_8434);
and U9004 (N_9004,N_7652,N_7095);
xor U9005 (N_9005,N_8680,N_8250);
nand U9006 (N_9006,N_8896,N_7446);
nor U9007 (N_9007,N_7384,N_7956);
nand U9008 (N_9008,N_7035,N_8197);
nand U9009 (N_9009,N_7858,N_8656);
nand U9010 (N_9010,N_6652,N_6791);
nor U9011 (N_9011,N_6385,N_7782);
nor U9012 (N_9012,N_7818,N_6066);
nand U9013 (N_9013,N_8001,N_7200);
xnor U9014 (N_9014,N_8232,N_8162);
nand U9015 (N_9015,N_7995,N_8331);
nor U9016 (N_9016,N_7826,N_7933);
nand U9017 (N_9017,N_7112,N_7969);
nand U9018 (N_9018,N_6232,N_7841);
or U9019 (N_9019,N_6844,N_8525);
and U9020 (N_9020,N_7081,N_7978);
nand U9021 (N_9021,N_7239,N_6128);
or U9022 (N_9022,N_8509,N_8992);
or U9023 (N_9023,N_8120,N_7934);
nor U9024 (N_9024,N_6629,N_8606);
xor U9025 (N_9025,N_7186,N_7698);
nor U9026 (N_9026,N_7071,N_7359);
or U9027 (N_9027,N_8990,N_8645);
nand U9028 (N_9028,N_7373,N_8712);
or U9029 (N_9029,N_7151,N_8164);
or U9030 (N_9030,N_7092,N_7983);
and U9031 (N_9031,N_6820,N_7816);
nor U9032 (N_9032,N_7353,N_7753);
or U9033 (N_9033,N_6985,N_6019);
and U9034 (N_9034,N_8215,N_7465);
xnor U9035 (N_9035,N_8345,N_8475);
and U9036 (N_9036,N_7810,N_6548);
xor U9037 (N_9037,N_6477,N_6658);
or U9038 (N_9038,N_7883,N_6503);
xnor U9039 (N_9039,N_7972,N_6220);
nand U9040 (N_9040,N_6416,N_8826);
xnor U9041 (N_9041,N_8796,N_6235);
xnor U9042 (N_9042,N_8751,N_6002);
nand U9043 (N_9043,N_6297,N_7851);
or U9044 (N_9044,N_8426,N_7792);
nor U9045 (N_9045,N_7120,N_8445);
nand U9046 (N_9046,N_7477,N_8088);
or U9047 (N_9047,N_8378,N_7119);
and U9048 (N_9048,N_7561,N_6344);
xor U9049 (N_9049,N_7820,N_6885);
and U9050 (N_9050,N_7715,N_8711);
nor U9051 (N_9051,N_8844,N_6901);
and U9052 (N_9052,N_8581,N_7617);
xor U9053 (N_9053,N_8756,N_8316);
and U9054 (N_9054,N_8291,N_7107);
or U9055 (N_9055,N_8562,N_6606);
and U9056 (N_9056,N_6971,N_8192);
nand U9057 (N_9057,N_7322,N_8810);
or U9058 (N_9058,N_6902,N_7909);
xnor U9059 (N_9059,N_6014,N_7419);
nand U9060 (N_9060,N_7575,N_8731);
and U9061 (N_9061,N_7130,N_8633);
xnor U9062 (N_9062,N_7868,N_6701);
xor U9063 (N_9063,N_6252,N_6254);
nand U9064 (N_9064,N_6990,N_7136);
or U9065 (N_9065,N_6412,N_8256);
nand U9066 (N_9066,N_7847,N_8596);
xnor U9067 (N_9067,N_8179,N_6445);
xor U9068 (N_9068,N_7448,N_7478);
and U9069 (N_9069,N_7884,N_8949);
xnor U9070 (N_9070,N_6177,N_8743);
nor U9071 (N_9071,N_7835,N_7098);
and U9072 (N_9072,N_7572,N_6660);
nor U9073 (N_9073,N_7040,N_6143);
or U9074 (N_9074,N_7512,N_7655);
and U9075 (N_9075,N_8785,N_7552);
and U9076 (N_9076,N_7226,N_8255);
nand U9077 (N_9077,N_7270,N_6741);
and U9078 (N_9078,N_7844,N_8501);
xnor U9079 (N_9079,N_8056,N_7400);
nand U9080 (N_9080,N_6358,N_8038);
and U9081 (N_9081,N_6012,N_8940);
or U9082 (N_9082,N_6432,N_7704);
xnor U9083 (N_9083,N_6541,N_8683);
xnor U9084 (N_9084,N_6546,N_6871);
or U9085 (N_9085,N_7410,N_8403);
or U9086 (N_9086,N_6435,N_8512);
and U9087 (N_9087,N_8853,N_8758);
xor U9088 (N_9088,N_8350,N_6936);
nor U9089 (N_9089,N_6053,N_8715);
xor U9090 (N_9090,N_7308,N_7965);
nor U9091 (N_9091,N_8762,N_8640);
or U9092 (N_9092,N_7295,N_8690);
and U9093 (N_9093,N_8004,N_6245);
and U9094 (N_9094,N_8200,N_6389);
nor U9095 (N_9095,N_8086,N_6894);
and U9096 (N_9096,N_7436,N_6137);
nand U9097 (N_9097,N_7372,N_7897);
or U9098 (N_9098,N_7754,N_8040);
nand U9099 (N_9099,N_6896,N_8817);
xnor U9100 (N_9100,N_8809,N_8486);
xor U9101 (N_9101,N_8182,N_8076);
nor U9102 (N_9102,N_7018,N_7605);
or U9103 (N_9103,N_7251,N_6746);
nor U9104 (N_9104,N_8789,N_8852);
xor U9105 (N_9105,N_8891,N_6476);
nor U9106 (N_9106,N_8318,N_7705);
xor U9107 (N_9107,N_6035,N_7767);
xnor U9108 (N_9108,N_7519,N_6005);
nor U9109 (N_9109,N_6628,N_6459);
nor U9110 (N_9110,N_7929,N_8140);
nand U9111 (N_9111,N_6838,N_8689);
and U9112 (N_9112,N_7452,N_7959);
or U9113 (N_9113,N_6011,N_7985);
and U9114 (N_9114,N_7639,N_6227);
xor U9115 (N_9115,N_6281,N_8152);
nor U9116 (N_9116,N_8334,N_8110);
nand U9117 (N_9117,N_8439,N_7079);
xnor U9118 (N_9118,N_6188,N_6931);
nor U9119 (N_9119,N_6591,N_6353);
xnor U9120 (N_9120,N_8611,N_6041);
xor U9121 (N_9121,N_6133,N_8832);
nor U9122 (N_9122,N_7356,N_7195);
nor U9123 (N_9123,N_6860,N_6168);
xnor U9124 (N_9124,N_6830,N_8221);
or U9125 (N_9125,N_6626,N_8700);
nand U9126 (N_9126,N_7537,N_7779);
xor U9127 (N_9127,N_8150,N_8929);
xor U9128 (N_9128,N_7730,N_7689);
nand U9129 (N_9129,N_8580,N_6185);
nand U9130 (N_9130,N_7197,N_8091);
or U9131 (N_9131,N_7520,N_7756);
nand U9132 (N_9132,N_6560,N_7574);
nand U9133 (N_9133,N_6106,N_7840);
and U9134 (N_9134,N_7357,N_8511);
or U9135 (N_9135,N_6020,N_8871);
nand U9136 (N_9136,N_6715,N_8154);
and U9137 (N_9137,N_8095,N_7582);
nand U9138 (N_9138,N_6178,N_8505);
or U9139 (N_9139,N_8764,N_7522);
and U9140 (N_9140,N_7598,N_7640);
or U9141 (N_9141,N_8269,N_8630);
xor U9142 (N_9142,N_7694,N_7194);
nand U9143 (N_9143,N_7049,N_8414);
or U9144 (N_9144,N_7966,N_7862);
nor U9145 (N_9145,N_6260,N_7333);
and U9146 (N_9146,N_8499,N_6393);
xor U9147 (N_9147,N_8588,N_6813);
nand U9148 (N_9148,N_6515,N_6157);
nor U9149 (N_9149,N_6236,N_8917);
nor U9150 (N_9150,N_7674,N_8208);
nor U9151 (N_9151,N_7736,N_8904);
nor U9152 (N_9152,N_8365,N_8695);
or U9153 (N_9153,N_6898,N_7707);
nor U9154 (N_9154,N_8377,N_6025);
xor U9155 (N_9155,N_6161,N_6600);
or U9156 (N_9156,N_8558,N_8209);
and U9157 (N_9157,N_6602,N_7800);
nand U9158 (N_9158,N_7409,N_8792);
and U9159 (N_9159,N_7039,N_7155);
nor U9160 (N_9160,N_8777,N_8135);
nand U9161 (N_9161,N_7977,N_8216);
or U9162 (N_9162,N_8233,N_7695);
xnor U9163 (N_9163,N_8382,N_7102);
nor U9164 (N_9164,N_8530,N_6132);
nor U9165 (N_9165,N_6292,N_7882);
xor U9166 (N_9166,N_8077,N_6149);
nand U9167 (N_9167,N_7463,N_8213);
nor U9168 (N_9168,N_7693,N_8615);
nor U9169 (N_9169,N_8390,N_8666);
nand U9170 (N_9170,N_7660,N_8142);
and U9171 (N_9171,N_8470,N_7544);
and U9172 (N_9172,N_7922,N_6247);
nand U9173 (N_9173,N_6109,N_7115);
nand U9174 (N_9174,N_8790,N_7848);
nor U9175 (N_9175,N_7108,N_7449);
xor U9176 (N_9176,N_6290,N_8986);
nor U9177 (N_9177,N_7662,N_6273);
xor U9178 (N_9178,N_8778,N_7341);
xor U9179 (N_9179,N_8648,N_7626);
nand U9180 (N_9180,N_7257,N_7044);
nor U9181 (N_9181,N_6582,N_7623);
xnor U9182 (N_9182,N_6145,N_7555);
and U9183 (N_9183,N_8863,N_6234);
nor U9184 (N_9184,N_8719,N_8031);
xnor U9185 (N_9185,N_8921,N_8612);
nor U9186 (N_9186,N_7292,N_8014);
and U9187 (N_9187,N_7163,N_8768);
or U9188 (N_9188,N_6499,N_7427);
nand U9189 (N_9189,N_7228,N_8673);
nor U9190 (N_9190,N_6342,N_6140);
and U9191 (N_9191,N_8103,N_8181);
and U9192 (N_9192,N_6552,N_6265);
nand U9193 (N_9193,N_8663,N_6315);
xor U9194 (N_9194,N_7828,N_8676);
nand U9195 (N_9195,N_7627,N_6309);
nand U9196 (N_9196,N_6904,N_8429);
xnor U9197 (N_9197,N_6138,N_6561);
nor U9198 (N_9198,N_7369,N_6704);
or U9199 (N_9199,N_6259,N_8157);
and U9200 (N_9200,N_6664,N_8902);
nand U9201 (N_9201,N_6593,N_8447);
xor U9202 (N_9202,N_8653,N_6105);
or U9203 (N_9203,N_6864,N_7113);
xnor U9204 (N_9204,N_6821,N_7303);
and U9205 (N_9205,N_6368,N_6598);
or U9206 (N_9206,N_6070,N_6840);
or U9207 (N_9207,N_7732,N_6121);
or U9208 (N_9208,N_8293,N_8259);
xor U9209 (N_9209,N_8498,N_6886);
or U9210 (N_9210,N_8988,N_8727);
nand U9211 (N_9211,N_6967,N_8463);
or U9212 (N_9212,N_6521,N_8123);
nor U9213 (N_9213,N_7618,N_6073);
nor U9214 (N_9214,N_6566,N_7731);
and U9215 (N_9215,N_6766,N_6078);
nor U9216 (N_9216,N_6743,N_7164);
nand U9217 (N_9217,N_7880,N_6513);
or U9218 (N_9218,N_6524,N_7533);
or U9219 (N_9219,N_6150,N_7233);
or U9220 (N_9220,N_6246,N_7720);
nor U9221 (N_9221,N_8951,N_8258);
or U9222 (N_9222,N_7172,N_7406);
or U9223 (N_9223,N_6243,N_6468);
xnor U9224 (N_9224,N_8053,N_7344);
or U9225 (N_9225,N_6376,N_8189);
and U9226 (N_9226,N_8803,N_8257);
or U9227 (N_9227,N_8959,N_6869);
nand U9228 (N_9228,N_7700,N_7518);
or U9229 (N_9229,N_6549,N_7930);
nand U9230 (N_9230,N_8857,N_6190);
xor U9231 (N_9231,N_8322,N_6090);
and U9232 (N_9232,N_6721,N_6302);
and U9233 (N_9233,N_8254,N_8178);
or U9234 (N_9234,N_8129,N_8707);
nand U9235 (N_9235,N_6239,N_7149);
or U9236 (N_9236,N_8834,N_6303);
nor U9237 (N_9237,N_6547,N_7718);
xnor U9238 (N_9238,N_8818,N_6287);
nor U9239 (N_9239,N_7162,N_8093);
xor U9240 (N_9240,N_6843,N_6230);
or U9241 (N_9241,N_6540,N_8313);
nand U9242 (N_9242,N_7907,N_8087);
xnor U9243 (N_9243,N_7622,N_6672);
nand U9244 (N_9244,N_8609,N_8728);
nand U9245 (N_9245,N_7370,N_8554);
or U9246 (N_9246,N_7747,N_8537);
or U9247 (N_9247,N_8206,N_6941);
nand U9248 (N_9248,N_7009,N_6427);
nor U9249 (N_9249,N_8880,N_6648);
and U9250 (N_9250,N_6553,N_6777);
nor U9251 (N_9251,N_7528,N_7248);
or U9252 (N_9252,N_6848,N_8854);
and U9253 (N_9253,N_7974,N_6845);
or U9254 (N_9254,N_7986,N_6768);
nand U9255 (N_9255,N_7952,N_6313);
xnor U9256 (N_9256,N_7403,N_8211);
xnor U9257 (N_9257,N_8416,N_7258);
nor U9258 (N_9258,N_7794,N_8991);
and U9259 (N_9259,N_6293,N_6331);
xnor U9260 (N_9260,N_7814,N_6055);
xnor U9261 (N_9261,N_6630,N_8819);
and U9262 (N_9262,N_8829,N_6951);
or U9263 (N_9263,N_7212,N_6980);
xnor U9264 (N_9264,N_6594,N_7831);
nand U9265 (N_9265,N_7843,N_7566);
and U9266 (N_9266,N_7179,N_8926);
or U9267 (N_9267,N_8718,N_8165);
or U9268 (N_9268,N_8999,N_8346);
nor U9269 (N_9269,N_7760,N_8235);
xor U9270 (N_9270,N_8627,N_7424);
nand U9271 (N_9271,N_6021,N_8954);
nand U9272 (N_9272,N_6029,N_8526);
nand U9273 (N_9273,N_8850,N_7713);
or U9274 (N_9274,N_8772,N_8133);
and U9275 (N_9275,N_7834,N_6206);
nand U9276 (N_9276,N_6905,N_6584);
nor U9277 (N_9277,N_7371,N_7000);
or U9278 (N_9278,N_8924,N_7545);
and U9279 (N_9279,N_6643,N_7289);
xnor U9280 (N_9280,N_8000,N_6175);
and U9281 (N_9281,N_7709,N_8565);
nor U9282 (N_9282,N_6530,N_6436);
xnor U9283 (N_9283,N_8280,N_8945);
nor U9284 (N_9284,N_7964,N_6891);
nor U9285 (N_9285,N_8708,N_6329);
or U9286 (N_9286,N_8557,N_7171);
or U9287 (N_9287,N_7062,N_8376);
nand U9288 (N_9288,N_8669,N_7672);
xnor U9289 (N_9289,N_6983,N_7159);
nor U9290 (N_9290,N_6054,N_6559);
nor U9291 (N_9291,N_8117,N_6879);
xnor U9292 (N_9292,N_6018,N_8412);
and U9293 (N_9293,N_7529,N_7932);
or U9294 (N_9294,N_6097,N_7808);
xnor U9295 (N_9295,N_6127,N_7799);
or U9296 (N_9296,N_7766,N_6386);
xnor U9297 (N_9297,N_7309,N_7323);
nand U9298 (N_9298,N_8387,N_8464);
nand U9299 (N_9299,N_8224,N_8138);
or U9300 (N_9300,N_7253,N_7650);
nor U9301 (N_9301,N_8618,N_6264);
nor U9302 (N_9302,N_8248,N_7474);
nor U9303 (N_9303,N_8396,N_8413);
nand U9304 (N_9304,N_6597,N_6650);
or U9305 (N_9305,N_7690,N_8273);
nand U9306 (N_9306,N_7022,N_7464);
nor U9307 (N_9307,N_6839,N_8935);
nor U9308 (N_9308,N_7990,N_6214);
or U9309 (N_9309,N_8845,N_6982);
nor U9310 (N_9310,N_6948,N_7712);
and U9311 (N_9311,N_6224,N_8374);
or U9312 (N_9312,N_6362,N_8214);
and U9313 (N_9313,N_6976,N_8620);
nor U9314 (N_9314,N_7085,N_8134);
nor U9315 (N_9315,N_8828,N_7404);
nor U9316 (N_9316,N_7502,N_7152);
nand U9317 (N_9317,N_8568,N_6280);
nand U9318 (N_9318,N_6815,N_6670);
xnor U9319 (N_9319,N_6732,N_7319);
nand U9320 (N_9320,N_6348,N_6796);
and U9321 (N_9321,N_8239,N_7935);
and U9322 (N_9322,N_7468,N_7348);
and U9323 (N_9323,N_6666,N_7230);
or U9324 (N_9324,N_6216,N_7422);
and U9325 (N_9325,N_6801,N_7578);
or U9326 (N_9326,N_7174,N_7511);
or U9327 (N_9327,N_7823,N_7679);
nand U9328 (N_9328,N_6663,N_8641);
nor U9329 (N_9329,N_6174,N_7265);
and U9330 (N_9330,N_6166,N_7277);
nor U9331 (N_9331,N_6656,N_7648);
or U9332 (N_9332,N_8220,N_8393);
nand U9333 (N_9333,N_8160,N_6441);
and U9334 (N_9334,N_8617,N_6863);
and U9335 (N_9335,N_8518,N_8685);
and U9336 (N_9336,N_7856,N_7165);
and U9337 (N_9337,N_7614,N_8981);
and U9338 (N_9338,N_7073,N_7889);
or U9339 (N_9339,N_8514,N_8781);
xor U9340 (N_9340,N_8922,N_8102);
nand U9341 (N_9341,N_8602,N_6738);
nand U9342 (N_9342,N_8825,N_8422);
or U9343 (N_9343,N_6938,N_6159);
and U9344 (N_9344,N_6209,N_7931);
and U9345 (N_9345,N_7314,N_7781);
nand U9346 (N_9346,N_7750,N_6364);
nor U9347 (N_9347,N_8864,N_7514);
nor U9348 (N_9348,N_7176,N_6424);
or U9349 (N_9349,N_8025,N_7505);
and U9350 (N_9350,N_7047,N_7992);
or U9351 (N_9351,N_7066,N_8372);
and U9352 (N_9352,N_8655,N_8879);
and U9353 (N_9353,N_7524,N_8311);
xor U9354 (N_9354,N_8462,N_7287);
xor U9355 (N_9355,N_6409,N_8983);
nor U9356 (N_9356,N_7493,N_7306);
or U9357 (N_9357,N_6024,N_7530);
and U9358 (N_9358,N_6330,N_8952);
nand U9359 (N_9359,N_6739,N_6271);
nand U9360 (N_9360,N_8381,N_8106);
and U9361 (N_9361,N_6696,N_6420);
nand U9362 (N_9362,N_6085,N_6500);
or U9363 (N_9363,N_6764,N_8912);
xnor U9364 (N_9364,N_7989,N_7236);
or U9365 (N_9365,N_7571,N_7435);
or U9366 (N_9366,N_7878,N_7282);
nor U9367 (N_9367,N_7778,N_6927);
and U9368 (N_9368,N_6022,N_8099);
nor U9369 (N_9369,N_8353,N_8684);
xnor U9370 (N_9370,N_8191,N_7378);
nand U9371 (N_9371,N_8698,N_7645);
nor U9372 (N_9372,N_6398,N_8636);
nand U9373 (N_9373,N_6867,N_7874);
nand U9374 (N_9374,N_6295,N_7157);
xor U9375 (N_9375,N_6966,N_6550);
xnor U9376 (N_9376,N_7338,N_6542);
nor U9377 (N_9377,N_6651,N_7998);
or U9378 (N_9378,N_8720,N_8262);
or U9379 (N_9379,N_7094,N_6760);
nand U9380 (N_9380,N_8104,N_7898);
nand U9381 (N_9381,N_8306,N_8210);
nand U9382 (N_9382,N_8996,N_7527);
nor U9383 (N_9383,N_8029,N_8428);
or U9384 (N_9384,N_6251,N_7927);
nor U9385 (N_9385,N_8533,N_7203);
or U9386 (N_9386,N_6917,N_8808);
or U9387 (N_9387,N_8173,N_7007);
and U9388 (N_9388,N_8515,N_8765);
xnor U9389 (N_9389,N_7680,N_6478);
nand U9390 (N_9390,N_6167,N_6103);
xor U9391 (N_9391,N_7812,N_7122);
nand U9392 (N_9392,N_6633,N_8253);
or U9393 (N_9393,N_6852,N_8234);
nor U9394 (N_9394,N_6835,N_6609);
or U9395 (N_9395,N_8049,N_6599);
nand U9396 (N_9396,N_7688,N_7421);
nand U9397 (N_9397,N_6915,N_7489);
xnor U9398 (N_9398,N_8180,N_8228);
and U9399 (N_9399,N_6356,N_8096);
xor U9400 (N_9400,N_8094,N_8885);
or U9401 (N_9401,N_8174,N_6687);
and U9402 (N_9402,N_7084,N_8510);
nand U9403 (N_9403,N_7012,N_6590);
and U9404 (N_9404,N_7391,N_7202);
nand U9405 (N_9405,N_8843,N_6993);
xnor U9406 (N_9406,N_8691,N_7173);
xor U9407 (N_9407,N_7137,N_7414);
nor U9408 (N_9408,N_7426,N_7788);
nand U9409 (N_9409,N_6678,N_8392);
or U9410 (N_9410,N_7397,N_6102);
and U9411 (N_9411,N_8692,N_7548);
and U9412 (N_9412,N_7456,N_8265);
nor U9413 (N_9413,N_8171,N_6802);
and U9414 (N_9414,N_7268,N_6562);
and U9415 (N_9415,N_8406,N_8156);
xnor U9416 (N_9416,N_6792,N_8035);
and U9417 (N_9417,N_7472,N_8783);
or U9418 (N_9418,N_7616,N_6793);
and U9419 (N_9419,N_6182,N_6854);
or U9420 (N_9420,N_8534,N_6505);
and U9421 (N_9421,N_6893,N_6786);
and U9422 (N_9422,N_7111,N_7991);
and U9423 (N_9423,N_8763,N_6907);
nand U9424 (N_9424,N_7169,N_6810);
nor U9425 (N_9425,N_8915,N_8199);
and U9426 (N_9426,N_7342,N_6525);
or U9427 (N_9427,N_6622,N_7182);
nand U9428 (N_9428,N_6977,N_6383);
and U9429 (N_9429,N_6442,N_6874);
xnor U9430 (N_9430,N_6984,N_7774);
and U9431 (N_9431,N_8497,N_7661);
nand U9432 (N_9432,N_8185,N_6415);
and U9433 (N_9433,N_6113,N_6842);
or U9434 (N_9434,N_6229,N_6072);
and U9435 (N_9435,N_8846,N_8137);
and U9436 (N_9436,N_7875,N_7250);
nand U9437 (N_9437,N_6595,N_8517);
nand U9438 (N_9438,N_8305,N_7015);
and U9439 (N_9439,N_7402,N_8744);
and U9440 (N_9440,N_8941,N_6636);
nor U9441 (N_9441,N_8139,N_6935);
and U9442 (N_9442,N_7070,N_7559);
or U9443 (N_9443,N_8882,N_8908);
nor U9444 (N_9444,N_8993,N_8423);
xor U9445 (N_9445,N_6900,N_8621);
nor U9446 (N_9446,N_6605,N_7219);
nor U9447 (N_9447,N_8046,N_7337);
nand U9448 (N_9448,N_6814,N_7361);
or U9449 (N_9449,N_6646,N_6564);
and U9450 (N_9450,N_6272,N_7328);
nand U9451 (N_9451,N_7735,N_8592);
or U9452 (N_9452,N_6501,N_7543);
nand U9453 (N_9453,N_6308,N_7600);
xor U9454 (N_9454,N_7673,N_8070);
nand U9455 (N_9455,N_7266,N_7153);
nand U9456 (N_9456,N_8321,N_7532);
nor U9457 (N_9457,N_6059,N_7646);
xnor U9458 (N_9458,N_8674,N_6472);
or U9459 (N_9459,N_6180,N_6667);
nor U9460 (N_9460,N_8761,N_7829);
xnor U9461 (N_9461,N_6205,N_6887);
xnor U9462 (N_9462,N_8100,N_7293);
nor U9463 (N_9463,N_6092,N_8585);
nand U9464 (N_9464,N_6527,N_6833);
nor U9465 (N_9465,N_8726,N_8082);
or U9466 (N_9466,N_8176,N_8433);
xor U9467 (N_9467,N_8485,N_7852);
and U9468 (N_9468,N_6139,N_6173);
xor U9469 (N_9469,N_7891,N_6061);
xnor U9470 (N_9470,N_7975,N_8714);
or U9471 (N_9471,N_6702,N_8401);
or U9472 (N_9472,N_6467,N_6352);
or U9473 (N_9473,N_8292,N_8937);
and U9474 (N_9474,N_7860,N_6675);
and U9475 (N_9475,N_6705,N_6288);
xnor U9476 (N_9476,N_7089,N_8974);
xnor U9477 (N_9477,N_6575,N_8605);
nand U9478 (N_9478,N_7658,N_6765);
nor U9479 (N_9479,N_8755,N_8041);
nand U9480 (N_9480,N_6405,N_8753);
nand U9481 (N_9481,N_8802,N_7383);
or U9482 (N_9482,N_7432,N_8007);
or U9483 (N_9483,N_8686,N_6475);
nand U9484 (N_9484,N_6576,N_7540);
or U9485 (N_9485,N_6627,N_8170);
and U9486 (N_9486,N_8649,N_6339);
nand U9487 (N_9487,N_6510,N_7670);
xor U9488 (N_9488,N_8252,N_7984);
xor U9489 (N_9489,N_7041,N_7940);
nor U9490 (N_9490,N_6752,N_6099);
or U9491 (N_9491,N_6526,N_7077);
or U9492 (N_9492,N_6381,N_8347);
xor U9493 (N_9493,N_7597,N_6811);
and U9494 (N_9494,N_8024,N_8298);
nor U9495 (N_9495,N_8892,N_6987);
nor U9496 (N_9496,N_7025,N_7096);
xor U9497 (N_9497,N_7791,N_6380);
or U9498 (N_9498,N_7768,N_6470);
xor U9499 (N_9499,N_8861,N_7387);
nor U9500 (N_9500,N_7280,N_6062);
nor U9501 (N_9501,N_6425,N_8840);
nor U9502 (N_9502,N_6222,N_8793);
or U9503 (N_9503,N_7607,N_7486);
nand U9504 (N_9504,N_6058,N_8923);
nand U9505 (N_9505,N_8600,N_7584);
and U9506 (N_9506,N_8811,N_7595);
nor U9507 (N_9507,N_8011,N_8194);
nand U9508 (N_9508,N_6289,N_8107);
and U9509 (N_9509,N_7722,N_7769);
or U9510 (N_9510,N_6337,N_6728);
nor U9511 (N_9511,N_6581,N_6294);
nor U9512 (N_9512,N_8938,N_8874);
and U9513 (N_9513,N_8646,N_6603);
nand U9514 (N_9514,N_8159,N_8061);
and U9515 (N_9515,N_8184,N_8905);
xnor U9516 (N_9516,N_7926,N_7216);
nand U9517 (N_9517,N_6535,N_7612);
xnor U9518 (N_9518,N_8071,N_7615);
nor U9519 (N_9519,N_6240,N_7238);
xor U9520 (N_9520,N_6892,N_8402);
and U9521 (N_9521,N_6518,N_7492);
nor U9522 (N_9522,N_6890,N_8052);
or U9523 (N_9523,N_8386,N_6074);
xnor U9524 (N_9524,N_6350,N_6828);
or U9525 (N_9525,N_6640,N_8798);
nor U9526 (N_9526,N_6975,N_6808);
nand U9527 (N_9527,N_8677,N_6758);
or U9528 (N_9528,N_8866,N_7232);
and U9529 (N_9529,N_8607,N_6889);
xor U9530 (N_9530,N_8431,N_6158);
nor U9531 (N_9531,N_7755,N_7517);
and U9532 (N_9532,N_8639,N_6611);
and U9533 (N_9533,N_7951,N_7339);
nand U9534 (N_9534,N_6955,N_7031);
or U9535 (N_9535,N_6233,N_8335);
or U9536 (N_9536,N_7676,N_7547);
xor U9537 (N_9537,N_7916,N_6403);
and U9538 (N_9538,N_6578,N_6165);
nor U9539 (N_9539,N_6779,N_6558);
nand U9540 (N_9540,N_7939,N_6722);
nor U9541 (N_9541,N_7064,N_6100);
xnor U9542 (N_9542,N_8187,N_7034);
nand U9543 (N_9543,N_7054,N_8651);
or U9544 (N_9544,N_8327,N_7981);
nand U9545 (N_9545,N_6668,N_8218);
or U9546 (N_9546,N_6397,N_7326);
and U9547 (N_9547,N_8397,N_7013);
or U9548 (N_9548,N_8504,N_8021);
xor U9549 (N_9549,N_7494,N_8008);
nor U9550 (N_9550,N_6676,N_8821);
and U9551 (N_9551,N_6079,N_6032);
and U9552 (N_9552,N_8590,N_8155);
nor U9553 (N_9553,N_6387,N_8804);
or U9554 (N_9554,N_8824,N_6355);
and U9555 (N_9555,N_8297,N_6241);
or U9556 (N_9556,N_7350,N_8979);
or U9557 (N_9557,N_6207,N_8242);
and U9558 (N_9558,N_8198,N_7033);
xnor U9559 (N_9559,N_8446,N_7088);
or U9560 (N_9560,N_7921,N_6677);
nand U9561 (N_9561,N_6536,N_7330);
xnor U9562 (N_9562,N_6278,N_7043);
and U9563 (N_9563,N_6763,N_7531);
and U9564 (N_9564,N_6703,N_8204);
or U9565 (N_9565,N_6154,N_7010);
and U9566 (N_9566,N_7501,N_8420);
or U9567 (N_9567,N_6610,N_8287);
or U9568 (N_9568,N_6734,N_6419);
xor U9569 (N_9569,N_8309,N_6218);
or U9570 (N_9570,N_7300,N_6873);
nor U9571 (N_9571,N_6125,N_7599);
nand U9572 (N_9572,N_7729,N_7104);
or U9573 (N_9573,N_6969,N_6195);
nor U9574 (N_9574,N_8274,N_8652);
xnor U9575 (N_9575,N_7118,N_6706);
and U9576 (N_9576,N_6081,N_8290);
nor U9577 (N_9577,N_7428,N_7893);
or U9578 (N_9578,N_6316,N_6949);
and U9579 (N_9579,N_8328,N_8400);
or U9580 (N_9580,N_6261,N_6699);
nand U9581 (N_9581,N_7302,N_8805);
and U9582 (N_9582,N_8489,N_8304);
or U9583 (N_9583,N_6880,N_8482);
xnor U9584 (N_9584,N_6096,N_6794);
nor U9585 (N_9585,N_8784,N_8125);
and U9586 (N_9586,N_7017,N_6928);
nand U9587 (N_9587,N_6338,N_7667);
or U9588 (N_9588,N_7681,N_7377);
or U9589 (N_9589,N_6131,N_6333);
or U9590 (N_9590,N_6800,N_7177);
and U9591 (N_9591,N_6870,N_8492);
and U9592 (N_9592,N_6798,N_8593);
or U9593 (N_9593,N_8472,N_6554);
nor U9594 (N_9594,N_8670,N_6517);
or U9595 (N_9595,N_7240,N_8303);
xnor U9596 (N_9596,N_6645,N_7272);
and U9597 (N_9597,N_8126,N_6714);
nor U9598 (N_9598,N_8479,N_6034);
nand U9599 (N_9599,N_6319,N_7905);
or U9600 (N_9600,N_6816,N_8085);
nand U9601 (N_9601,N_8343,N_6080);
nor U9602 (N_9602,N_7587,N_8555);
nand U9603 (N_9603,N_7692,N_6181);
xnor U9604 (N_9604,N_8260,N_6506);
and U9605 (N_9605,N_8203,N_6944);
or U9606 (N_9606,N_8359,N_8454);
nor U9607 (N_9607,N_6068,N_7471);
and U9608 (N_9608,N_8773,N_6989);
xnor U9609 (N_9609,N_7147,N_7601);
nor U9610 (N_9610,N_7093,N_6831);
or U9611 (N_9611,N_8918,N_8424);
or U9612 (N_9612,N_8528,N_6580);
nand U9613 (N_9613,N_6000,N_7273);
or U9614 (N_9614,N_6172,N_7221);
or U9615 (N_9615,N_6992,N_8058);
nor U9616 (N_9616,N_7804,N_7467);
nor U9617 (N_9617,N_7822,N_6489);
nor U9618 (N_9618,N_6819,N_6471);
nor U9619 (N_9619,N_6876,N_7873);
or U9620 (N_9620,N_8870,N_7687);
nand U9621 (N_9621,N_6396,N_6123);
and U9622 (N_9622,N_6680,N_8500);
xnor U9623 (N_9623,N_6248,N_7154);
nand U9624 (N_9624,N_8760,N_6392);
xnor U9625 (N_9625,N_7839,N_7635);
and U9626 (N_9626,N_7294,N_6946);
nor U9627 (N_9627,N_6514,N_7853);
nor U9628 (N_9628,N_6846,N_6269);
xnor U9629 (N_9629,N_7741,N_8083);
or U9630 (N_9630,N_7483,N_7946);
and U9631 (N_9631,N_7589,N_6130);
and U9632 (N_9632,N_6784,N_6903);
xor U9633 (N_9633,N_6556,N_8286);
nor U9634 (N_9634,N_7764,N_8028);
nand U9635 (N_9635,N_6428,N_8391);
and U9636 (N_9636,N_7305,N_6507);
or U9637 (N_9637,N_7894,N_6749);
xnor U9638 (N_9638,N_7550,N_6301);
nand U9639 (N_9639,N_6466,N_6266);
and U9640 (N_9640,N_7244,N_8266);
or U9641 (N_9641,N_6144,N_6653);
or U9642 (N_9642,N_8831,N_6458);
or U9643 (N_9643,N_6634,N_8409);
nand U9644 (N_9644,N_6963,N_8966);
nand U9645 (N_9645,N_8080,N_8681);
nor U9646 (N_9646,N_6211,N_7696);
xor U9647 (N_9647,N_6401,N_8586);
or U9648 (N_9648,N_8319,N_8595);
or U9649 (N_9649,N_8101,N_8738);
or U9650 (N_9650,N_6730,N_6731);
or U9651 (N_9651,N_6225,N_7863);
or U9652 (N_9652,N_7444,N_6249);
or U9653 (N_9653,N_6994,N_8502);
nand U9654 (N_9654,N_8893,N_6030);
nand U9655 (N_9655,N_8249,N_7610);
nor U9656 (N_9656,N_8907,N_8750);
and U9657 (N_9657,N_7837,N_8830);
nor U9658 (N_9658,N_8894,N_6809);
or U9659 (N_9659,N_7993,N_7521);
nor U9660 (N_9660,N_7534,N_6868);
xnor U9661 (N_9661,N_6720,N_6539);
xnor U9662 (N_9662,N_7360,N_8748);
nor U9663 (N_9663,N_7411,N_8594);
or U9664 (N_9664,N_7324,N_7955);
or U9665 (N_9665,N_8022,N_8559);
or U9666 (N_9666,N_6780,N_7748);
and U9667 (N_9667,N_8055,N_6444);
xnor U9668 (N_9668,N_7242,N_6298);
xor U9669 (N_9669,N_6529,N_7442);
xnor U9670 (N_9670,N_7274,N_6347);
and U9671 (N_9671,N_7220,N_8953);
nor U9672 (N_9672,N_8856,N_6142);
xor U9673 (N_9673,N_8398,N_8355);
nand U9674 (N_9674,N_8556,N_8635);
and U9675 (N_9675,N_6110,N_6711);
xor U9676 (N_9676,N_8629,N_8749);
nor U9677 (N_9677,N_8136,N_8236);
nor U9678 (N_9678,N_6557,N_6343);
or U9679 (N_9679,N_7859,N_7011);
or U9680 (N_9680,N_8268,N_7376);
xor U9681 (N_9681,N_6422,N_7208);
and U9682 (N_9682,N_6455,N_7105);
nand U9683 (N_9683,N_8587,N_7286);
nand U9684 (N_9684,N_8267,N_6827);
nand U9685 (N_9685,N_8065,N_7229);
nand U9686 (N_9686,N_8148,N_6713);
nand U9687 (N_9687,N_8342,N_6391);
and U9688 (N_9688,N_8442,N_6351);
and U9689 (N_9689,N_6279,N_6511);
nand U9690 (N_9690,N_8956,N_6400);
nand U9691 (N_9691,N_6908,N_6770);
nor U9692 (N_9692,N_7255,N_7401);
nand U9693 (N_9693,N_8141,N_6803);
and U9694 (N_9694,N_6997,N_8067);
nor U9695 (N_9695,N_8769,N_7457);
nand U9696 (N_9696,N_8705,N_6408);
xor U9697 (N_9697,N_8440,N_8075);
xor U9698 (N_9698,N_8862,N_7283);
and U9699 (N_9699,N_8963,N_8575);
or U9700 (N_9700,N_8576,N_6063);
xnor U9701 (N_9701,N_8147,N_6767);
nand U9702 (N_9702,N_8042,N_8539);
or U9703 (N_9703,N_7004,N_6379);
nor U9704 (N_9704,N_8578,N_7198);
nand U9705 (N_9705,N_8661,N_7503);
and U9706 (N_9706,N_8295,N_8296);
nand U9707 (N_9707,N_7131,N_6747);
nor U9708 (N_9708,N_7473,N_8109);
nand U9709 (N_9709,N_8112,N_8090);
nand U9710 (N_9710,N_6939,N_7313);
xor U9711 (N_9711,N_7669,N_6748);
xor U9712 (N_9712,N_8368,N_8132);
and U9713 (N_9713,N_8550,N_6543);
nor U9714 (N_9714,N_7262,N_7842);
and U9715 (N_9715,N_6060,N_6050);
and U9716 (N_9716,N_8207,N_6932);
nor U9717 (N_9717,N_6832,N_8480);
and U9718 (N_9718,N_6978,N_7708);
or U9719 (N_9719,N_7797,N_7063);
and U9720 (N_9720,N_8452,N_7145);
or U9721 (N_9721,N_7028,N_8244);
xnor U9722 (N_9722,N_8251,N_7659);
nor U9723 (N_9723,N_8418,N_7415);
xnor U9724 (N_9724,N_7609,N_7817);
xor U9725 (N_9725,N_6884,N_8842);
nand U9726 (N_9726,N_6250,N_7144);
nand U9727 (N_9727,N_8521,N_6162);
nand U9728 (N_9728,N_6134,N_8363);
nor U9729 (N_9729,N_8212,N_6775);
nor U9730 (N_9730,N_8895,N_6862);
xnor U9731 (N_9731,N_8704,N_8713);
or U9732 (N_9732,N_7777,N_6270);
nand U9733 (N_9733,N_7807,N_8186);
or U9734 (N_9734,N_7437,N_8143);
nand U9735 (N_9735,N_7237,N_7761);
nor U9736 (N_9736,N_8920,N_8358);
nand U9737 (N_9737,N_6001,N_7407);
or U9738 (N_9738,N_8989,N_6474);
nor U9739 (N_9739,N_6023,N_6523);
or U9740 (N_9740,N_7970,N_8544);
xnor U9741 (N_9741,N_7475,N_7606);
nor U9742 (N_9742,N_7796,N_7895);
nand U9743 (N_9743,N_6563,N_6681);
nor U9744 (N_9744,N_6617,N_6095);
and U9745 (N_9745,N_8503,N_8084);
or U9746 (N_9746,N_6457,N_7187);
xor U9747 (N_9747,N_8223,N_6875);
nor U9748 (N_9748,N_6919,N_7317);
nor U9749 (N_9749,N_6601,N_7743);
or U9750 (N_9750,N_8867,N_6788);
or U9751 (N_9751,N_6712,N_6755);
nor U9752 (N_9752,N_8980,N_6335);
and U9753 (N_9753,N_7918,N_8724);
and U9754 (N_9754,N_8299,N_6464);
or U9755 (N_9755,N_8399,N_8059);
nand U9756 (N_9756,N_7947,N_8166);
xor U9757 (N_9757,N_7281,N_8942);
xnor U9758 (N_9758,N_8740,N_7310);
and U9759 (N_9759,N_7312,N_6359);
nor U9760 (N_9760,N_7352,N_6141);
nor U9761 (N_9761,N_7919,N_6545);
nor U9762 (N_9762,N_6200,N_7484);
and U9763 (N_9763,N_8634,N_8227);
nor U9764 (N_9764,N_8583,N_8407);
nor U9765 (N_9765,N_7438,N_6346);
or U9766 (N_9766,N_7380,N_7008);
and U9767 (N_9767,N_8508,N_8626);
and U9768 (N_9768,N_7048,N_8373);
nand U9769 (N_9769,N_6736,N_8167);
and U9770 (N_9770,N_8456,N_7385);
and U9771 (N_9771,N_6953,N_6772);
nor U9772 (N_9772,N_8277,N_7497);
xor U9773 (N_9773,N_6307,N_6374);
nor U9774 (N_9774,N_6371,N_6744);
xor U9775 (N_9775,N_6589,N_8637);
or U9776 (N_9776,N_6754,N_7830);
nand U9777 (N_9777,N_8610,N_8717);
xor U9778 (N_9778,N_7447,N_7381);
or U9779 (N_9779,N_7936,N_8477);
or U9780 (N_9780,N_7836,N_8944);
nand U9781 (N_9781,N_6156,N_8441);
xor U9782 (N_9782,N_6108,N_6778);
nor U9783 (N_9783,N_8351,N_7362);
nor U9784 (N_9784,N_7653,N_7052);
and U9785 (N_9785,N_7591,N_6761);
nand U9786 (N_9786,N_6957,N_6429);
nor U9787 (N_9787,N_7999,N_6454);
nor U9788 (N_9788,N_8457,N_6069);
xor U9789 (N_9789,N_8348,N_7542);
or U9790 (N_9790,N_8308,N_7346);
and U9791 (N_9791,N_8163,N_8873);
or U9792 (N_9792,N_6013,N_8427);
xor U9793 (N_9793,N_7190,N_6437);
or U9794 (N_9794,N_7116,N_7558);
xnor U9795 (N_9795,N_6929,N_7210);
xor U9796 (N_9796,N_6238,N_8177);
nor U9797 (N_9797,N_6357,N_6574);
or U9798 (N_9798,N_7068,N_8496);
and U9799 (N_9799,N_6382,N_7243);
nor U9800 (N_9800,N_8002,N_6502);
or U9801 (N_9801,N_7042,N_7055);
nand U9802 (N_9802,N_7666,N_6945);
nand U9803 (N_9803,N_8385,N_6671);
and U9804 (N_9804,N_7714,N_8622);
nor U9805 (N_9805,N_7958,N_6729);
nand U9806 (N_9806,N_7567,N_8560);
and U9807 (N_9807,N_8903,N_8230);
nand U9808 (N_9808,N_7643,N_6116);
nor U9809 (N_9809,N_7334,N_7269);
xnor U9810 (N_9810,N_6285,N_7861);
and U9811 (N_9811,N_7634,N_8946);
nand U9812 (N_9812,N_6858,N_6310);
nand U9813 (N_9813,N_8950,N_7368);
nor U9814 (N_9814,N_7183,N_8081);
nand U9815 (N_9815,N_8675,N_7006);
or U9816 (N_9816,N_6257,N_7740);
nor U9817 (N_9817,N_6853,N_7291);
nor U9818 (N_9818,N_6733,N_7461);
or U9819 (N_9819,N_6850,N_8694);
nor U9820 (N_9820,N_8884,N_6583);
nand U9821 (N_9821,N_8483,N_8601);
nand U9822 (N_9822,N_7513,N_6282);
nand U9823 (N_9823,N_8394,N_6164);
nand U9824 (N_9824,N_7611,N_7374);
nor U9825 (N_9825,N_8632,N_6926);
nand U9826 (N_9826,N_7390,N_7733);
xnor U9827 (N_9827,N_7196,N_7101);
nand U9828 (N_9828,N_7087,N_7016);
and U9829 (N_9829,N_6488,N_6544);
or U9830 (N_9830,N_8364,N_8383);
and U9831 (N_9831,N_6958,N_7045);
nand U9832 (N_9832,N_7060,N_8127);
or U9833 (N_9833,N_7420,N_7942);
xnor U9834 (N_9834,N_8806,N_8812);
or U9835 (N_9835,N_6112,N_7920);
nor U9836 (N_9836,N_8549,N_7389);
and U9837 (N_9837,N_8919,N_8018);
nor U9838 (N_9838,N_7900,N_7785);
xnor U9839 (N_9839,N_8312,N_6790);
nor U9840 (N_9840,N_8060,N_6686);
nand U9841 (N_9841,N_6710,N_6504);
nor U9842 (N_9842,N_8909,N_7784);
nand U9843 (N_9843,N_8188,N_8775);
nor U9844 (N_9844,N_8231,N_8948);
xor U9845 (N_9845,N_7425,N_6179);
or U9846 (N_9846,N_8118,N_7780);
xnor U9847 (N_9847,N_6450,N_6328);
or U9848 (N_9848,N_7546,N_6118);
and U9849 (N_9849,N_8716,N_7592);
and U9850 (N_9850,N_8776,N_6228);
nand U9851 (N_9851,N_8947,N_8701);
nor U9852 (N_9852,N_8116,N_7752);
nor U9853 (N_9853,N_7913,N_6217);
nand U9854 (N_9854,N_6537,N_8430);
and U9855 (N_9855,N_8967,N_7762);
or U9856 (N_9856,N_8371,N_7539);
or U9857 (N_9857,N_6184,N_7139);
nand U9858 (N_9858,N_8168,N_7364);
and U9859 (N_9859,N_8044,N_8013);
xor U9860 (N_9860,N_8589,N_8465);
nor U9861 (N_9861,N_7161,N_8072);
or U9862 (N_9862,N_6136,N_6135);
or U9863 (N_9863,N_7140,N_8339);
and U9864 (N_9864,N_8964,N_6751);
xor U9865 (N_9865,N_7507,N_7855);
xnor U9866 (N_9866,N_8933,N_7886);
xor U9867 (N_9867,N_8461,N_8410);
xor U9868 (N_9868,N_6056,N_8598);
nand U9869 (N_9869,N_6120,N_7719);
or U9870 (N_9870,N_8384,N_6119);
or U9871 (N_9871,N_8914,N_7734);
xnor U9872 (N_9872,N_8190,N_8016);
nor U9873 (N_9873,N_6592,N_8994);
or U9874 (N_9874,N_7331,N_6049);
and U9875 (N_9875,N_6981,N_7725);
or U9876 (N_9876,N_7469,N_8771);
or U9877 (N_9877,N_6805,N_8816);
xor U9878 (N_9878,N_8302,N_8356);
nand U9879 (N_9879,N_7580,N_7980);
nand U9880 (N_9880,N_6849,N_7412);
nand U9881 (N_9881,N_7392,N_6147);
nor U9882 (N_9882,N_7019,N_6213);
and U9883 (N_9883,N_7490,N_7329);
or U9884 (N_9884,N_7738,N_6988);
nand U9885 (N_9885,N_8516,N_8723);
nor U9886 (N_9886,N_6433,N_6460);
nor U9887 (N_9887,N_6750,N_7211);
nor U9888 (N_9888,N_6531,N_8978);
or U9889 (N_9889,N_7872,N_8471);
xor U9890 (N_9890,N_7395,N_7343);
nand U9891 (N_9891,N_7885,N_8579);
and U9892 (N_9892,N_7254,N_6226);
or U9893 (N_9893,N_7466,N_8613);
or U9894 (N_9894,N_8913,N_8419);
or U9895 (N_9895,N_7256,N_8710);
nand U9896 (N_9896,N_6189,N_7789);
or U9897 (N_9897,N_6950,N_7647);
nand U9898 (N_9898,N_6692,N_7845);
nand U9899 (N_9899,N_8647,N_7249);
nand U9900 (N_9900,N_7866,N_8567);
nand U9901 (N_9901,N_6043,N_8366);
nand U9902 (N_9902,N_8955,N_6776);
nor U9903 (N_9903,N_7218,N_6823);
nand U9904 (N_9904,N_6332,N_8453);
or U9905 (N_9905,N_7298,N_6995);
nor U9906 (N_9906,N_6924,N_7217);
nor U9907 (N_9907,N_6986,N_6153);
nor U9908 (N_9908,N_6596,N_6952);
nor U9909 (N_9909,N_6759,N_6661);
nand U9910 (N_9910,N_7168,N_8752);
and U9911 (N_9911,N_7551,N_7059);
and U9912 (N_9912,N_6960,N_7776);
xnor U9913 (N_9913,N_8005,N_7443);
nor U9914 (N_9914,N_7345,N_6719);
or U9915 (N_9915,N_8217,N_6469);
xnor U9916 (N_9916,N_8573,N_7354);
nand U9917 (N_9917,N_6799,N_8326);
and U9918 (N_9918,N_6045,N_7798);
or U9919 (N_9919,N_7504,N_7604);
and U9920 (N_9920,N_7908,N_6007);
or U9921 (N_9921,N_6735,N_6641);
and U9922 (N_9922,N_6451,N_7386);
and U9923 (N_9923,N_7394,N_7053);
and U9924 (N_9924,N_8887,N_7206);
xnor U9925 (N_9925,N_8800,N_7644);
and U9926 (N_9926,N_7535,N_7441);
nand U9927 (N_9927,N_7937,N_6942);
xor U9928 (N_9928,N_6426,N_7677);
or U9929 (N_9929,N_7460,N_8523);
or U9930 (N_9930,N_6148,N_7963);
or U9931 (N_9931,N_8284,N_6812);
xor U9932 (N_9932,N_8973,N_8272);
and U9933 (N_9933,N_8438,N_6317);
nor U9934 (N_9934,N_8522,N_7026);
nand U9935 (N_9935,N_8340,N_8310);
nand U9936 (N_9936,N_8301,N_8417);
xnor U9937 (N_9937,N_8144,N_6117);
nor U9938 (N_9938,N_6498,N_6388);
and U9939 (N_9939,N_7664,N_8625);
xnor U9940 (N_9940,N_6847,N_7278);
and U9941 (N_9941,N_6771,N_6782);
xnor U9942 (N_9942,N_6882,N_7691);
nand U9943 (N_9943,N_6659,N_8644);
nor U9944 (N_9944,N_6492,N_6635);
xor U9945 (N_9945,N_7620,N_6888);
nor U9946 (N_9946,N_8767,N_6569);
and U9947 (N_9947,N_8995,N_8360);
nor U9948 (N_9948,N_6618,N_6300);
or U9949 (N_9949,N_7222,N_8459);
and U9950 (N_9950,N_6620,N_8687);
nor U9951 (N_9951,N_8039,N_7223);
xor U9952 (N_9952,N_7925,N_6742);
nor U9953 (N_9953,N_8927,N_8774);
xnor U9954 (N_9954,N_7510,N_6322);
nor U9955 (N_9955,N_7123,N_8786);
nor U9956 (N_9956,N_6349,N_7214);
nor U9957 (N_9957,N_8664,N_6447);
and U9958 (N_9958,N_6258,N_7192);
xnor U9959 (N_9959,N_6155,N_6625);
nand U9960 (N_9960,N_8965,N_7065);
nand U9961 (N_9961,N_7765,N_6146);
or U9962 (N_9962,N_8451,N_6336);
or U9963 (N_9963,N_7150,N_7737);
nand U9964 (N_9964,N_8657,N_7577);
nand U9965 (N_9965,N_7057,N_6726);
nand U9966 (N_9966,N_6774,N_7316);
xor U9967 (N_9967,N_7114,N_8513);
and U9968 (N_9968,N_7325,N_6276);
nor U9969 (N_9969,N_7910,N_8823);
nor U9970 (N_9970,N_6740,N_6413);
and U9971 (N_9971,N_6920,N_8119);
or U9972 (N_9972,N_6482,N_6657);
nor U9973 (N_9973,N_7124,N_8063);
or U9974 (N_9974,N_6623,N_8851);
nor U9975 (N_9975,N_7072,N_7225);
xnor U9976 (N_9976,N_8108,N_7129);
or U9977 (N_9977,N_6959,N_8890);
xnor U9978 (N_9978,N_8928,N_7462);
or U9979 (N_9979,N_8089,N_6395);
nand U9980 (N_9980,N_8531,N_6621);
nor U9981 (N_9981,N_7642,N_8283);
nand U9982 (N_9982,N_7949,N_8435);
xnor U9983 (N_9983,N_8314,N_7902);
nor U9984 (N_9984,N_8519,N_6970);
xor U9985 (N_9985,N_6616,N_7702);
xnor U9986 (N_9986,N_7987,N_8421);
nor U9987 (N_9987,N_6198,N_8124);
nor U9988 (N_9988,N_6277,N_7516);
or U9989 (N_9989,N_7175,N_8276);
nand U9990 (N_9990,N_6785,N_7685);
nand U9991 (N_9991,N_6201,N_8939);
or U9992 (N_9992,N_8865,N_7241);
nor U9993 (N_9993,N_8017,N_7275);
or U9994 (N_9994,N_6866,N_8969);
nor U9995 (N_9995,N_6027,N_7869);
or U9996 (N_9996,N_8671,N_8281);
nor U9997 (N_9997,N_6783,N_8012);
or U9998 (N_9998,N_6456,N_8279);
xor U9999 (N_9999,N_6923,N_6861);
or U10000 (N_10000,N_6717,N_6323);
and U10001 (N_10001,N_6916,N_6439);
nand U10002 (N_10002,N_7581,N_6363);
and U10003 (N_10003,N_7074,N_7181);
xor U10004 (N_10004,N_8219,N_8264);
xnor U10005 (N_10005,N_8997,N_7665);
nor U10006 (N_10006,N_7480,N_8658);
and U10007 (N_10007,N_6231,N_7260);
nand U10008 (N_10008,N_8113,N_7440);
or U10009 (N_10009,N_8561,N_6587);
and U10010 (N_10010,N_6275,N_8899);
xor U10011 (N_10011,N_6694,N_7619);
or U10012 (N_10012,N_6320,N_6191);
or U10013 (N_10013,N_6567,N_7967);
nand U10014 (N_10014,N_6091,N_6631);
and U10015 (N_10015,N_8702,N_8357);
xor U10016 (N_10016,N_7117,N_8970);
or U10017 (N_10017,N_7099,N_7957);
nor U10018 (N_10018,N_6199,N_6372);
xnor U10019 (N_10019,N_8729,N_6716);
or U10020 (N_10020,N_8263,N_8332);
or U10021 (N_10021,N_7654,N_7683);
nand U10022 (N_10022,N_7121,N_7790);
and U10023 (N_10023,N_7100,N_8437);
xor U10024 (N_10024,N_7960,N_7746);
nor U10025 (N_10025,N_6283,N_6568);
or U10026 (N_10026,N_8288,N_6015);
xnor U10027 (N_10027,N_6423,N_7982);
nand U10028 (N_10028,N_6709,N_6934);
nor U10029 (N_10029,N_6083,N_8225);
nor U10030 (N_10030,N_7924,N_8547);
and U10031 (N_10031,N_8571,N_6341);
and U10032 (N_10032,N_6911,N_7899);
and U10033 (N_10033,N_7832,N_8468);
xor U10034 (N_10034,N_8033,N_6943);
nand U10035 (N_10035,N_8491,N_7568);
nand U10036 (N_10036,N_6044,N_8958);
nand U10037 (N_10037,N_6274,N_8195);
and U10038 (N_10038,N_8553,N_6493);
xnor U10039 (N_10039,N_6490,N_7803);
nand U10040 (N_10040,N_7570,N_8527);
xnor U10041 (N_10041,N_7727,N_8934);
or U10042 (N_10042,N_8984,N_7973);
and U10043 (N_10043,N_8006,N_8051);
nand U10044 (N_10044,N_7349,N_8754);
nand U10045 (N_10045,N_6613,N_7160);
or U10046 (N_10046,N_6077,N_6585);
xnor U10047 (N_10047,N_7367,N_6797);
or U10048 (N_10048,N_8183,N_7434);
nor U10049 (N_10049,N_6052,N_6769);
nor U10050 (N_10050,N_8352,N_8529);
xnor U10051 (N_10051,N_8706,N_8642);
and U10052 (N_10052,N_7706,N_8476);
or U10053 (N_10053,N_7056,N_7697);
or U10054 (N_10054,N_8307,N_7491);
xnor U10055 (N_10055,N_6961,N_7311);
nor U10056 (N_10056,N_8535,N_6972);
xnor U10057 (N_10057,N_8010,N_7682);
xor U10058 (N_10058,N_7815,N_8484);
xnor U10059 (N_10059,N_8977,N_8742);
xor U10060 (N_10060,N_7245,N_8408);
nor U10061 (N_10061,N_6452,N_8285);
nand U10062 (N_10062,N_7744,N_6010);
or U10063 (N_10063,N_7488,N_7824);
and U10064 (N_10064,N_6296,N_8604);
nand U10065 (N_10065,N_7917,N_8432);
nor U10066 (N_10066,N_7775,N_7433);
xnor U10067 (N_10067,N_6673,N_6818);
and U10068 (N_10068,N_6375,N_7030);
or U10069 (N_10069,N_6004,N_7649);
nor U10070 (N_10070,N_8859,N_7146);
nand U10071 (N_10071,N_6065,N_6360);
or U10072 (N_10072,N_8034,N_6519);
xor U10073 (N_10073,N_8697,N_8925);
xnor U10074 (N_10074,N_6446,N_7110);
nand U10075 (N_10075,N_7613,N_7624);
nor U10076 (N_10076,N_6718,N_7506);
nor U10077 (N_10077,N_7067,N_6968);
nand U10078 (N_10078,N_8813,N_6851);
nor U10079 (N_10079,N_7772,N_7742);
or U10080 (N_10080,N_7479,N_7948);
nand U10081 (N_10081,N_6407,N_6991);
nor U10082 (N_10082,N_6017,N_6522);
and U10083 (N_10083,N_7996,N_7125);
nand U10084 (N_10084,N_6064,N_7603);
xnor U10085 (N_10085,N_7499,N_8975);
nor U10086 (N_10086,N_7971,N_7485);
nor U10087 (N_10087,N_8961,N_8875);
xnor U10088 (N_10088,N_6051,N_7002);
xnor U10089 (N_10089,N_6737,N_8336);
nand U10090 (N_10090,N_6009,N_6434);
xnor U10091 (N_10091,N_8161,N_7413);
nor U10092 (N_10092,N_6122,N_6508);
and U10093 (N_10093,N_8570,N_6370);
or U10094 (N_10094,N_7355,N_8878);
xnor U10095 (N_10095,N_7470,N_7086);
xnor U10096 (N_10096,N_8976,N_6075);
xor U10097 (N_10097,N_7994,N_8043);
and U10098 (N_10098,N_6579,N_7724);
xnor U10099 (N_10099,N_7979,N_6913);
or U10100 (N_10100,N_7633,N_6773);
xor U10101 (N_10101,N_6841,N_8900);
or U10102 (N_10102,N_7296,N_8545);
nor U10103 (N_10103,N_8815,N_7711);
xnor U10104 (N_10104,N_6689,N_8624);
and U10105 (N_10105,N_8591,N_6438);
or U10106 (N_10106,N_6203,N_7363);
and U10107 (N_10107,N_6373,N_8759);
and U10108 (N_10108,N_6124,N_6026);
or U10109 (N_10109,N_7668,N_6979);
nand U10110 (N_10110,N_6354,N_7630);
nor U10111 (N_10111,N_6325,N_6003);
or U10112 (N_10112,N_7912,N_7297);
nor U10113 (N_10113,N_6286,N_8146);
and U10114 (N_10114,N_7850,N_8079);
nand U10115 (N_10115,N_6006,N_6695);
and U10116 (N_10116,N_8665,N_8361);
nor U10117 (N_10117,N_8467,N_7763);
or U10118 (N_10118,N_6909,N_7656);
xor U10119 (N_10119,N_8872,N_7911);
or U10120 (N_10120,N_6082,N_6321);
or U10121 (N_10121,N_7109,N_8582);
nand U10122 (N_10122,N_6912,N_8725);
nand U10123 (N_10123,N_8069,N_8506);
nand U10124 (N_10124,N_8631,N_7867);
nand U10125 (N_10125,N_7536,N_6700);
nor U10126 (N_10126,N_8354,N_7787);
xor U10127 (N_10127,N_8145,N_8009);
nor U10128 (N_10128,N_8494,N_6256);
or U10129 (N_10129,N_8478,N_7227);
xnor U10130 (N_10130,N_7944,N_8822);
or U10131 (N_10131,N_6366,N_7451);
nand U10132 (N_10132,N_7082,N_8469);
nand U10133 (N_10133,N_7651,N_7809);
and U10134 (N_10134,N_6367,N_8699);
and U10135 (N_10135,N_7864,N_7135);
or U10136 (N_10136,N_8448,N_8741);
nor U10137 (N_10137,N_7588,N_8078);
nor U10138 (N_10138,N_8757,N_7128);
xnor U10139 (N_10139,N_7327,N_7090);
and U10140 (N_10140,N_6806,N_8569);
nand U10141 (N_10141,N_8278,N_8149);
and U10142 (N_10142,N_6872,N_6463);
nor U10143 (N_10143,N_8032,N_6479);
or U10144 (N_10144,N_7029,N_8444);
xor U10145 (N_10145,N_7906,N_8241);
and U10146 (N_10146,N_7318,N_7051);
and U10147 (N_10147,N_7158,N_8289);
or U10148 (N_10148,N_8650,N_7199);
nor U10149 (N_10149,N_7141,N_6268);
and U10150 (N_10150,N_7498,N_7284);
nand U10151 (N_10151,N_7408,N_7418);
nand U10152 (N_10152,N_7271,N_8936);
and U10153 (N_10153,N_6877,N_6449);
and U10154 (N_10154,N_6837,N_6324);
or U10155 (N_10155,N_6312,N_6443);
xnor U10156 (N_10156,N_7583,N_7950);
xnor U10157 (N_10157,N_8709,N_6473);
and U10158 (N_10158,N_6962,N_6067);
or U10159 (N_10159,N_7180,N_6314);
and U10160 (N_10160,N_8662,N_7388);
xnor U10161 (N_10161,N_7264,N_6918);
xor U10162 (N_10162,N_8971,N_6679);
and U10163 (N_10163,N_6033,N_7838);
or U10164 (N_10164,N_7020,N_8175);
or U10165 (N_10165,N_8794,N_6817);
xnor U10166 (N_10166,N_6572,N_8787);
nand U10167 (N_10167,N_8599,N_6163);
or U10168 (N_10168,N_6365,N_6088);
xor U10169 (N_10169,N_8050,N_8425);
nand U10170 (N_10170,N_7560,N_8733);
nand U10171 (N_10171,N_6973,N_6637);
xnor U10172 (N_10172,N_6588,N_7209);
nand U10173 (N_10173,N_6608,N_8238);
xnor U10174 (N_10174,N_8998,N_7749);
nor U10175 (N_10175,N_7632,N_8507);
xnor U10176 (N_10176,N_8551,N_6822);
and U10177 (N_10177,N_8449,N_7285);
nand U10178 (N_10178,N_7675,N_7854);
or U10179 (N_10179,N_7304,N_7621);
nand U10180 (N_10180,N_8722,N_7579);
or U10181 (N_10181,N_7430,N_6724);
nand U10182 (N_10182,N_7213,N_7833);
nand U10183 (N_10183,N_8487,N_7701);
xnor U10184 (N_10184,N_7594,N_6878);
nor U10185 (N_10185,N_8721,N_8889);
nand U10186 (N_10186,N_7078,N_7953);
nor U10187 (N_10187,N_7416,N_8577);
nor U10188 (N_10188,N_8202,N_6789);
nand U10189 (N_10189,N_7585,N_8030);
and U10190 (N_10190,N_7745,N_8130);
nor U10191 (N_10191,N_6565,N_8901);
and U10192 (N_10192,N_6291,N_6036);
and U10193 (N_10193,N_7728,N_6448);
nand U10194 (N_10194,N_7625,N_7142);
or U10195 (N_10195,N_6683,N_6855);
or U10196 (N_10196,N_8960,N_7458);
nand U10197 (N_10197,N_7061,N_8628);
and U10198 (N_10198,N_7525,N_7382);
and U10199 (N_10199,N_8972,N_7751);
and U10200 (N_10200,N_6196,N_7340);
xnor U10201 (N_10201,N_6170,N_6462);
or U10202 (N_10202,N_6076,N_8532);
or U10203 (N_10203,N_6390,N_7375);
or U10204 (N_10204,N_6340,N_7954);
xor U10205 (N_10205,N_8158,N_8574);
xor U10206 (N_10206,N_7132,N_6334);
nand U10207 (N_10207,N_8395,N_8968);
nor U10208 (N_10208,N_7526,N_8538);
and U10209 (N_10209,N_8836,N_8985);
nand U10210 (N_10210,N_7508,N_7231);
nand U10211 (N_10211,N_7641,N_7596);
xor U10212 (N_10212,N_6418,N_7178);
or U10213 (N_10213,N_7819,N_7523);
nand U10214 (N_10214,N_8795,N_6647);
nor U10215 (N_10215,N_7896,N_6115);
xor U10216 (N_10216,N_7487,N_8982);
and U10217 (N_10217,N_6804,N_7496);
and U10218 (N_10218,N_6410,N_8660);
or U10219 (N_10219,N_7663,N_6008);
nand U10220 (N_10220,N_7076,N_6881);
nor U10221 (N_10221,N_7246,N_8682);
and U10222 (N_10222,N_8466,N_8362);
nor U10223 (N_10223,N_6399,N_8693);
and U10224 (N_10224,N_8869,N_7657);
or U10225 (N_10225,N_6193,N_8703);
xor U10226 (N_10226,N_6836,N_8062);
and U10227 (N_10227,N_6906,N_6965);
and U10228 (N_10228,N_7968,N_7106);
xnor U10229 (N_10229,N_7771,N_6825);
nand U10230 (N_10230,N_6834,N_7716);
and U10231 (N_10231,N_6192,N_6219);
xnor U10232 (N_10232,N_7001,N_6632);
or U10233 (N_10233,N_7565,N_7608);
nor U10234 (N_10234,N_7877,N_7439);
nand U10235 (N_10235,N_6930,N_8092);
or U10236 (N_10236,N_6384,N_8495);
nor U10237 (N_10237,N_7299,N_6649);
xnor U10238 (N_10238,N_7938,N_6996);
xnor U10239 (N_10239,N_7075,N_7204);
nand U10240 (N_10240,N_8074,N_7050);
nand U10241 (N_10241,N_7166,N_8455);
and U10242 (N_10242,N_7134,N_6570);
nand U10243 (N_10243,N_6512,N_8696);
or U10244 (N_10244,N_7207,N_6897);
xnor U10245 (N_10245,N_8667,N_7686);
nand U10246 (N_10246,N_8247,N_8524);
or U10247 (N_10247,N_8105,N_6674);
nor U10248 (N_10248,N_6655,N_6402);
or U10249 (N_10249,N_6954,N_8098);
nand U10250 (N_10250,N_6028,N_7976);
xnor U10251 (N_10251,N_8566,N_8458);
nand U10252 (N_10252,N_6378,N_6727);
nand U10253 (N_10253,N_7091,N_7557);
nand U10254 (N_10254,N_7802,N_7569);
nand U10255 (N_10255,N_8858,N_7538);
and U10256 (N_10256,N_6638,N_8801);
or U10257 (N_10257,N_8490,N_7083);
or U10258 (N_10258,N_7710,N_8436);
or U10259 (N_10259,N_7038,N_8678);
or U10260 (N_10260,N_7636,N_8294);
nand U10261 (N_10261,N_7793,N_8745);
nand U10262 (N_10262,N_6311,N_8460);
or U10263 (N_10263,N_6654,N_8246);
and U10264 (N_10264,N_8003,N_6883);
nand U10265 (N_10265,N_6665,N_6781);
nor U10266 (N_10266,N_7901,N_8608);
nand U10267 (N_10267,N_7553,N_8172);
xnor U10268 (N_10268,N_6707,N_8205);
or U10269 (N_10269,N_8324,N_6087);
nor U10270 (N_10270,N_6484,N_7252);
or U10271 (N_10271,N_7366,N_8564);
xnor U10272 (N_10272,N_7857,N_6481);
xor U10273 (N_10273,N_8542,N_8196);
and U10274 (N_10274,N_7865,N_6639);
nor U10275 (N_10275,N_6642,N_8597);
or U10276 (N_10276,N_7887,N_8380);
or U10277 (N_10277,N_8746,N_7307);
nand U10278 (N_10278,N_7997,N_6480);
nand U10279 (N_10279,N_7148,N_6244);
nand U10280 (N_10280,N_6495,N_8488);
nor U10281 (N_10281,N_6345,N_8910);
and U10282 (N_10282,N_7431,N_8835);
nor U10283 (N_10283,N_7806,N_7138);
and U10284 (N_10284,N_7904,N_8073);
nand U10285 (N_10285,N_8883,N_6084);
nand U10286 (N_10286,N_6284,N_8779);
nor U10287 (N_10287,N_7482,N_8245);
xor U10288 (N_10288,N_6829,N_6038);
and U10289 (N_10289,N_6040,N_6202);
and U10290 (N_10290,N_7915,N_7396);
nor U10291 (N_10291,N_6745,N_8066);
or U10292 (N_10292,N_8548,N_6197);
and U10293 (N_10293,N_6183,N_8849);
or U10294 (N_10294,N_6369,N_7193);
nand U10295 (N_10295,N_7703,N_8855);
nor U10296 (N_10296,N_6223,N_7573);
xor U10297 (N_10297,N_7335,N_6921);
xnor U10298 (N_10298,N_8019,N_8367);
nor U10299 (N_10299,N_8338,N_6318);
nor U10300 (N_10300,N_8886,N_8275);
nor U10301 (N_10301,N_6486,N_8877);
or U10302 (N_10302,N_7923,N_7450);
xor U10303 (N_10303,N_6037,N_8770);
xnor U10304 (N_10304,N_7347,N_6612);
or U10305 (N_10305,N_6204,N_8057);
nor U10306 (N_10306,N_8111,N_8300);
and U10307 (N_10307,N_7726,N_7783);
and U10308 (N_10308,N_6586,N_7563);
nor U10309 (N_10309,N_6494,N_7593);
and U10310 (N_10310,N_6111,N_8814);
or U10311 (N_10311,N_7881,N_7871);
xor U10312 (N_10312,N_8654,N_7336);
and U10313 (N_10313,N_7758,N_7638);
nand U10314 (N_10314,N_8541,N_7455);
nor U10315 (N_10315,N_8325,N_8026);
or U10316 (N_10316,N_6509,N_7127);
nand U10317 (N_10317,N_8020,N_8572);
and U10318 (N_10318,N_7903,N_7321);
or U10319 (N_10319,N_7170,N_8638);
or U10320 (N_10320,N_7205,N_8037);
nor U10321 (N_10321,N_7167,N_6614);
and U10322 (N_10322,N_7549,N_7184);
nor U10323 (N_10323,N_6690,N_8837);
or U10324 (N_10324,N_8799,N_6684);
xnor U10325 (N_10325,N_8474,N_7014);
or U10326 (N_10326,N_8603,N_6644);
or U10327 (N_10327,N_7069,N_6406);
or U10328 (N_10328,N_7825,N_7201);
nor U10329 (N_10329,N_6757,N_7032);
xnor U10330 (N_10330,N_6306,N_6974);
or U10331 (N_10331,N_7365,N_6534);
xnor U10332 (N_10332,N_7024,N_8201);
xor U10333 (N_10333,N_6305,N_7631);
nor U10334 (N_10334,N_6169,N_8036);
xnor U10335 (N_10335,N_7185,N_6394);
nand U10336 (N_10336,N_7126,N_6160);
or U10337 (N_10337,N_8349,N_7247);
xor U10338 (N_10338,N_7037,N_8114);
nand U10339 (N_10339,N_6485,N_7279);
and U10340 (N_10340,N_6262,N_8643);
nor U10341 (N_10341,N_8222,N_7721);
xor U10342 (N_10342,N_8688,N_8054);
xnor U10343 (N_10343,N_6604,N_8552);
or U10344 (N_10344,N_7541,N_7454);
nand U10345 (N_10345,N_7263,N_6114);
xnor U10346 (N_10346,N_8838,N_6361);
nand U10347 (N_10347,N_8122,N_8847);
or U10348 (N_10348,N_8584,N_7576);
nand U10349 (N_10349,N_6046,N_7870);
or U10350 (N_10350,N_7892,N_8736);
and U10351 (N_10351,N_7379,N_7556);
nand U10352 (N_10352,N_6693,N_6857);
nand U10353 (N_10353,N_8732,N_6151);
xor U10354 (N_10354,N_6212,N_6532);
xor U10355 (N_10355,N_8619,N_6299);
nand U10356 (N_10356,N_6215,N_7801);
or U10357 (N_10357,N_7509,N_6685);
and U10358 (N_10358,N_6430,N_6326);
nand U10359 (N_10359,N_6865,N_6304);
and U10360 (N_10360,N_8315,N_6624);
nor U10361 (N_10361,N_7757,N_6465);
nor U10362 (N_10362,N_7805,N_6933);
xnor U10363 (N_10363,N_6461,N_6756);
or U10364 (N_10364,N_7215,N_7554);
nand U10365 (N_10365,N_7021,N_8881);
nor U10366 (N_10366,N_7602,N_6047);
or U10367 (N_10367,N_8737,N_8115);
nor U10368 (N_10368,N_7023,N_7476);
xor U10369 (N_10369,N_8443,N_8261);
or U10370 (N_10370,N_7445,N_6697);
or U10371 (N_10371,N_8064,N_6089);
nand U10372 (N_10372,N_6682,N_8323);
nor U10373 (N_10373,N_8045,N_8906);
or U10374 (N_10374,N_7723,N_8027);
or U10375 (N_10375,N_8766,N_6242);
nand U10376 (N_10376,N_8987,N_7259);
or U10377 (N_10377,N_6708,N_7453);
nor U10378 (N_10378,N_6071,N_7261);
or U10379 (N_10379,N_7103,N_7301);
or U10380 (N_10380,N_8860,N_8048);
nor U10381 (N_10381,N_7058,N_7962);
and U10382 (N_10382,N_7717,N_8520);
and U10383 (N_10383,N_8317,N_8930);
or U10384 (N_10384,N_7890,N_6528);
xor U10385 (N_10385,N_8369,N_6762);
nand U10386 (N_10386,N_8848,N_7481);
nor U10387 (N_10387,N_7027,N_8672);
or U10388 (N_10388,N_7562,N_7945);
xor U10389 (N_10389,N_7500,N_7813);
or U10390 (N_10390,N_8375,N_7678);
nor U10391 (N_10391,N_8668,N_6237);
nand U10392 (N_10392,N_6826,N_6048);
nand U10393 (N_10393,N_6691,N_8807);
or U10394 (N_10394,N_7398,N_7879);
xnor U10395 (N_10395,N_7003,N_8897);
xor U10396 (N_10396,N_7224,N_7188);
nand U10397 (N_10397,N_8388,N_7590);
nor U10398 (N_10398,N_6571,N_7080);
and U10399 (N_10399,N_6107,N_8888);
nand U10400 (N_10400,N_7143,N_6093);
xnor U10401 (N_10401,N_8237,N_8820);
xnor U10402 (N_10402,N_7914,N_8679);
or U10403 (N_10403,N_6039,N_8614);
or U10404 (N_10404,N_8957,N_7811);
and U10405 (N_10405,N_8169,N_6187);
or U10406 (N_10406,N_8876,N_7586);
nand U10407 (N_10407,N_8411,N_7097);
xnor U10408 (N_10408,N_8450,N_6453);
nand U10409 (N_10409,N_8563,N_6807);
or U10410 (N_10410,N_8916,N_8415);
xnor U10411 (N_10411,N_7628,N_8962);
nor U10412 (N_10412,N_6496,N_6947);
nand U10413 (N_10413,N_7699,N_7637);
nand U10414 (N_10414,N_6956,N_8023);
nand U10415 (N_10415,N_8151,N_6129);
or U10416 (N_10416,N_8229,N_6483);
and U10417 (N_10417,N_6824,N_8780);
nand U10418 (N_10418,N_6208,N_7393);
or U10419 (N_10419,N_7770,N_6031);
nor U10420 (N_10420,N_8734,N_8747);
nor U10421 (N_10421,N_8868,N_6615);
xnor U10422 (N_10422,N_8341,N_8782);
xor U10423 (N_10423,N_7036,N_6098);
nand U10424 (N_10424,N_7133,N_8370);
nand U10425 (N_10425,N_7234,N_8730);
or U10426 (N_10426,N_6086,N_6573);
nor U10427 (N_10427,N_7267,N_6520);
or U10428 (N_10428,N_6914,N_8333);
and U10429 (N_10429,N_7888,N_8337);
nand U10430 (N_10430,N_7961,N_7046);
nor U10431 (N_10431,N_6856,N_6538);
nor U10432 (N_10432,N_8841,N_6662);
and U10433 (N_10433,N_8735,N_6491);
and U10434 (N_10434,N_6688,N_7417);
and U10435 (N_10435,N_6186,N_8931);
or U10436 (N_10436,N_8270,N_7849);
xor U10437 (N_10437,N_8911,N_7235);
xor U10438 (N_10438,N_6267,N_6221);
nor U10439 (N_10439,N_7943,N_8226);
nand U10440 (N_10440,N_6152,N_8193);
or U10441 (N_10441,N_8097,N_8827);
or U10442 (N_10442,N_8344,N_8943);
nand U10443 (N_10443,N_7786,N_6126);
nand U10444 (N_10444,N_6940,N_8833);
or U10445 (N_10445,N_8047,N_7941);
or U10446 (N_10446,N_8739,N_7671);
nor U10447 (N_10447,N_7399,N_6998);
or U10448 (N_10448,N_7156,N_7988);
nand U10449 (N_10449,N_6999,N_8320);
or U10450 (N_10450,N_8493,N_6795);
xor U10451 (N_10451,N_8153,N_8131);
and U10452 (N_10452,N_6497,N_7928);
xnor U10453 (N_10453,N_6042,N_8898);
xor U10454 (N_10454,N_6171,N_6255);
xnor U10455 (N_10455,N_7827,N_7739);
or U10456 (N_10456,N_8546,N_8616);
nor U10457 (N_10457,N_6101,N_8330);
and U10458 (N_10458,N_8015,N_8405);
nor U10459 (N_10459,N_6417,N_8329);
nor U10460 (N_10460,N_6925,N_8379);
nor U10461 (N_10461,N_6104,N_8243);
nor U10462 (N_10462,N_7005,N_6194);
or U10463 (N_10463,N_6487,N_6753);
nand U10464 (N_10464,N_7459,N_6263);
or U10465 (N_10465,N_8932,N_8788);
nand U10466 (N_10466,N_8481,N_6922);
nor U10467 (N_10467,N_8791,N_7191);
or U10468 (N_10468,N_6016,N_6411);
or U10469 (N_10469,N_7332,N_7358);
xnor U10470 (N_10470,N_7315,N_7290);
and U10471 (N_10471,N_8473,N_6404);
xor U10472 (N_10472,N_7276,N_7423);
nand U10473 (N_10473,N_8068,N_6210);
nor U10474 (N_10474,N_7495,N_8389);
xnor U10475 (N_10475,N_6094,N_6377);
and U10476 (N_10476,N_6577,N_6698);
nor U10477 (N_10477,N_6910,N_7629);
nor U10478 (N_10478,N_7795,N_7821);
or U10479 (N_10479,N_6253,N_6669);
or U10480 (N_10480,N_8271,N_6899);
nor U10481 (N_10481,N_7189,N_6431);
nand U10482 (N_10482,N_6964,N_7846);
nor U10483 (N_10483,N_6787,N_8623);
nand U10484 (N_10484,N_6414,N_8128);
xnor U10485 (N_10485,N_7684,N_7773);
xor U10486 (N_10486,N_7320,N_6725);
and U10487 (N_10487,N_6421,N_7351);
xor U10488 (N_10488,N_6895,N_6619);
nand U10489 (N_10489,N_7429,N_7405);
nor U10490 (N_10490,N_6057,N_6937);
and U10491 (N_10491,N_8540,N_8839);
or U10492 (N_10492,N_6176,N_6723);
nor U10493 (N_10493,N_6607,N_6551);
or U10494 (N_10494,N_8797,N_8240);
nand U10495 (N_10495,N_6440,N_8282);
nand U10496 (N_10496,N_8404,N_7876);
or U10497 (N_10497,N_7564,N_6516);
or U10498 (N_10498,N_8536,N_6859);
or U10499 (N_10499,N_8121,N_7759);
nor U10500 (N_10500,N_7314,N_8495);
and U10501 (N_10501,N_7121,N_8347);
nor U10502 (N_10502,N_6969,N_8395);
nor U10503 (N_10503,N_7020,N_6963);
nand U10504 (N_10504,N_8809,N_7248);
nand U10505 (N_10505,N_7100,N_8648);
and U10506 (N_10506,N_6738,N_7477);
and U10507 (N_10507,N_6107,N_8240);
xnor U10508 (N_10508,N_8336,N_8540);
or U10509 (N_10509,N_6048,N_7658);
xor U10510 (N_10510,N_7509,N_6599);
xnor U10511 (N_10511,N_8149,N_7102);
or U10512 (N_10512,N_6809,N_7655);
and U10513 (N_10513,N_6247,N_7697);
and U10514 (N_10514,N_7200,N_6644);
nor U10515 (N_10515,N_6973,N_8040);
xor U10516 (N_10516,N_8287,N_8977);
xnor U10517 (N_10517,N_8989,N_7206);
nor U10518 (N_10518,N_8443,N_7294);
or U10519 (N_10519,N_7276,N_6117);
and U10520 (N_10520,N_6346,N_8520);
and U10521 (N_10521,N_7216,N_7297);
and U10522 (N_10522,N_7709,N_8444);
and U10523 (N_10523,N_7969,N_6470);
nand U10524 (N_10524,N_8450,N_7277);
xor U10525 (N_10525,N_6856,N_6008);
nor U10526 (N_10526,N_8303,N_8601);
nand U10527 (N_10527,N_8339,N_8056);
and U10528 (N_10528,N_7079,N_6466);
nand U10529 (N_10529,N_6411,N_7413);
nand U10530 (N_10530,N_6513,N_7634);
xnor U10531 (N_10531,N_6893,N_8105);
nor U10532 (N_10532,N_8761,N_6413);
and U10533 (N_10533,N_7293,N_8542);
nand U10534 (N_10534,N_7011,N_6980);
nand U10535 (N_10535,N_7801,N_8761);
xnor U10536 (N_10536,N_7292,N_8911);
xor U10537 (N_10537,N_6247,N_6126);
nand U10538 (N_10538,N_6220,N_7673);
nor U10539 (N_10539,N_6570,N_6002);
nand U10540 (N_10540,N_6731,N_7998);
or U10541 (N_10541,N_7397,N_7774);
and U10542 (N_10542,N_7226,N_6856);
or U10543 (N_10543,N_7211,N_8294);
and U10544 (N_10544,N_7105,N_6402);
nand U10545 (N_10545,N_7175,N_8098);
xnor U10546 (N_10546,N_7010,N_6334);
nand U10547 (N_10547,N_7516,N_8938);
or U10548 (N_10548,N_7457,N_8893);
nand U10549 (N_10549,N_8541,N_7024);
or U10550 (N_10550,N_6569,N_6476);
xnor U10551 (N_10551,N_7437,N_6363);
xor U10552 (N_10552,N_6391,N_7061);
xnor U10553 (N_10553,N_8365,N_8147);
nor U10554 (N_10554,N_8727,N_6482);
xnor U10555 (N_10555,N_8327,N_6625);
nand U10556 (N_10556,N_6560,N_7205);
xnor U10557 (N_10557,N_6044,N_8478);
xnor U10558 (N_10558,N_7743,N_7053);
nor U10559 (N_10559,N_8097,N_6963);
xnor U10560 (N_10560,N_7046,N_8202);
and U10561 (N_10561,N_6632,N_6261);
and U10562 (N_10562,N_6687,N_6260);
or U10563 (N_10563,N_7117,N_6270);
nand U10564 (N_10564,N_7320,N_8876);
and U10565 (N_10565,N_7740,N_6513);
nand U10566 (N_10566,N_6071,N_8516);
xor U10567 (N_10567,N_6699,N_6014);
and U10568 (N_10568,N_7389,N_6983);
nor U10569 (N_10569,N_6548,N_6960);
nand U10570 (N_10570,N_8835,N_7386);
or U10571 (N_10571,N_8769,N_7780);
nand U10572 (N_10572,N_6612,N_7289);
nor U10573 (N_10573,N_8552,N_8302);
xor U10574 (N_10574,N_7278,N_8664);
or U10575 (N_10575,N_8792,N_6785);
xor U10576 (N_10576,N_7377,N_6079);
nor U10577 (N_10577,N_8875,N_7501);
and U10578 (N_10578,N_6695,N_6503);
nand U10579 (N_10579,N_8865,N_7487);
or U10580 (N_10580,N_7075,N_7196);
nand U10581 (N_10581,N_8346,N_6416);
nor U10582 (N_10582,N_8285,N_7253);
and U10583 (N_10583,N_8954,N_6530);
xnor U10584 (N_10584,N_8393,N_7049);
and U10585 (N_10585,N_7519,N_7473);
and U10586 (N_10586,N_6229,N_6605);
or U10587 (N_10587,N_6548,N_7020);
or U10588 (N_10588,N_7495,N_6458);
and U10589 (N_10589,N_8810,N_7282);
nand U10590 (N_10590,N_8284,N_8088);
nor U10591 (N_10591,N_6453,N_7072);
nor U10592 (N_10592,N_8775,N_6504);
nand U10593 (N_10593,N_7505,N_8577);
xnor U10594 (N_10594,N_7976,N_8586);
and U10595 (N_10595,N_6693,N_6848);
nand U10596 (N_10596,N_6166,N_6532);
nand U10597 (N_10597,N_7308,N_8489);
nor U10598 (N_10598,N_8559,N_8069);
nor U10599 (N_10599,N_8841,N_8252);
or U10600 (N_10600,N_8689,N_8633);
and U10601 (N_10601,N_8915,N_8571);
nand U10602 (N_10602,N_7282,N_6543);
nand U10603 (N_10603,N_7436,N_6021);
nor U10604 (N_10604,N_8960,N_6696);
xnor U10605 (N_10605,N_8774,N_8269);
xor U10606 (N_10606,N_7105,N_8364);
and U10607 (N_10607,N_8855,N_6696);
and U10608 (N_10608,N_6918,N_8914);
nand U10609 (N_10609,N_6167,N_7355);
xor U10610 (N_10610,N_6880,N_6539);
or U10611 (N_10611,N_7882,N_8187);
nand U10612 (N_10612,N_6732,N_8238);
or U10613 (N_10613,N_7617,N_8239);
nor U10614 (N_10614,N_6035,N_6627);
nand U10615 (N_10615,N_6395,N_7489);
and U10616 (N_10616,N_7563,N_8776);
or U10617 (N_10617,N_7939,N_8537);
xnor U10618 (N_10618,N_7585,N_7142);
or U10619 (N_10619,N_6827,N_6649);
and U10620 (N_10620,N_7902,N_8450);
and U10621 (N_10621,N_8626,N_7317);
xnor U10622 (N_10622,N_8474,N_6998);
or U10623 (N_10623,N_7305,N_8749);
nor U10624 (N_10624,N_7133,N_8792);
or U10625 (N_10625,N_6374,N_6350);
or U10626 (N_10626,N_8298,N_8678);
nand U10627 (N_10627,N_8398,N_7944);
xor U10628 (N_10628,N_7523,N_6230);
nor U10629 (N_10629,N_6726,N_7147);
nand U10630 (N_10630,N_6792,N_6747);
xor U10631 (N_10631,N_7086,N_6850);
or U10632 (N_10632,N_8977,N_6584);
xor U10633 (N_10633,N_6144,N_7525);
nor U10634 (N_10634,N_8026,N_7247);
or U10635 (N_10635,N_8735,N_7961);
nor U10636 (N_10636,N_7700,N_6045);
xnor U10637 (N_10637,N_6953,N_6679);
nor U10638 (N_10638,N_8117,N_7550);
nand U10639 (N_10639,N_7948,N_8632);
xnor U10640 (N_10640,N_8978,N_6153);
nor U10641 (N_10641,N_7633,N_8798);
xnor U10642 (N_10642,N_8109,N_6752);
nand U10643 (N_10643,N_7098,N_7941);
xnor U10644 (N_10644,N_8838,N_8680);
and U10645 (N_10645,N_7553,N_7921);
nor U10646 (N_10646,N_6590,N_6940);
and U10647 (N_10647,N_6221,N_6260);
or U10648 (N_10648,N_7641,N_8709);
nor U10649 (N_10649,N_6346,N_8435);
and U10650 (N_10650,N_6695,N_7751);
xor U10651 (N_10651,N_7031,N_8466);
and U10652 (N_10652,N_6660,N_8917);
xor U10653 (N_10653,N_7554,N_8480);
nor U10654 (N_10654,N_6412,N_7620);
nor U10655 (N_10655,N_8674,N_7147);
and U10656 (N_10656,N_8624,N_6305);
nor U10657 (N_10657,N_7575,N_8308);
nor U10658 (N_10658,N_6166,N_6561);
nor U10659 (N_10659,N_8616,N_8014);
nand U10660 (N_10660,N_6970,N_7708);
xnor U10661 (N_10661,N_8340,N_6597);
nand U10662 (N_10662,N_8470,N_8321);
and U10663 (N_10663,N_8213,N_7415);
nand U10664 (N_10664,N_8457,N_7541);
nand U10665 (N_10665,N_8485,N_7787);
xor U10666 (N_10666,N_7518,N_7052);
nand U10667 (N_10667,N_7853,N_7321);
or U10668 (N_10668,N_8681,N_7374);
nor U10669 (N_10669,N_8914,N_7288);
or U10670 (N_10670,N_6094,N_6105);
or U10671 (N_10671,N_6852,N_7761);
and U10672 (N_10672,N_6538,N_7586);
nand U10673 (N_10673,N_8854,N_7334);
and U10674 (N_10674,N_7407,N_6576);
nor U10675 (N_10675,N_8664,N_8160);
and U10676 (N_10676,N_8160,N_7100);
nand U10677 (N_10677,N_8707,N_8157);
or U10678 (N_10678,N_6408,N_8564);
or U10679 (N_10679,N_7659,N_8346);
and U10680 (N_10680,N_8089,N_7644);
and U10681 (N_10681,N_7552,N_8170);
xnor U10682 (N_10682,N_8685,N_7566);
nand U10683 (N_10683,N_8807,N_6022);
nand U10684 (N_10684,N_6099,N_8675);
and U10685 (N_10685,N_6938,N_8473);
nor U10686 (N_10686,N_6247,N_8902);
nor U10687 (N_10687,N_6210,N_7836);
xor U10688 (N_10688,N_8785,N_6584);
xor U10689 (N_10689,N_6758,N_8379);
nor U10690 (N_10690,N_6948,N_8994);
nor U10691 (N_10691,N_6213,N_8399);
nand U10692 (N_10692,N_8239,N_7965);
xnor U10693 (N_10693,N_7221,N_7662);
or U10694 (N_10694,N_6990,N_8850);
xnor U10695 (N_10695,N_7458,N_8080);
and U10696 (N_10696,N_8711,N_7615);
nor U10697 (N_10697,N_6776,N_6642);
nor U10698 (N_10698,N_7752,N_8230);
nand U10699 (N_10699,N_8430,N_8398);
nand U10700 (N_10700,N_7635,N_6270);
nand U10701 (N_10701,N_8984,N_8215);
nor U10702 (N_10702,N_8116,N_7325);
nor U10703 (N_10703,N_8244,N_8464);
xnor U10704 (N_10704,N_7140,N_8900);
and U10705 (N_10705,N_8081,N_8849);
nor U10706 (N_10706,N_8434,N_6089);
xor U10707 (N_10707,N_7373,N_8218);
xnor U10708 (N_10708,N_6912,N_6567);
and U10709 (N_10709,N_6183,N_6802);
nor U10710 (N_10710,N_8842,N_6896);
and U10711 (N_10711,N_8530,N_6186);
or U10712 (N_10712,N_7636,N_8283);
xnor U10713 (N_10713,N_8618,N_8346);
or U10714 (N_10714,N_6876,N_6431);
nand U10715 (N_10715,N_8311,N_8191);
nor U10716 (N_10716,N_7364,N_8425);
nand U10717 (N_10717,N_7869,N_8506);
nor U10718 (N_10718,N_6526,N_6372);
nor U10719 (N_10719,N_6904,N_7195);
or U10720 (N_10720,N_6838,N_7442);
nor U10721 (N_10721,N_8914,N_7414);
xor U10722 (N_10722,N_7329,N_7273);
nor U10723 (N_10723,N_6750,N_8039);
and U10724 (N_10724,N_8200,N_8188);
xnor U10725 (N_10725,N_6952,N_7219);
and U10726 (N_10726,N_6192,N_7439);
nand U10727 (N_10727,N_6637,N_8144);
nand U10728 (N_10728,N_7355,N_6905);
or U10729 (N_10729,N_8173,N_7562);
nand U10730 (N_10730,N_7091,N_8092);
nor U10731 (N_10731,N_8982,N_7742);
and U10732 (N_10732,N_7857,N_7582);
nand U10733 (N_10733,N_7737,N_6960);
nor U10734 (N_10734,N_7093,N_6482);
or U10735 (N_10735,N_6631,N_6889);
xor U10736 (N_10736,N_8486,N_8982);
or U10737 (N_10737,N_8531,N_6566);
nand U10738 (N_10738,N_6469,N_7500);
xor U10739 (N_10739,N_8148,N_6936);
nand U10740 (N_10740,N_8052,N_7073);
nor U10741 (N_10741,N_6607,N_7058);
nor U10742 (N_10742,N_7681,N_7515);
xor U10743 (N_10743,N_8459,N_7522);
nand U10744 (N_10744,N_7499,N_6283);
nand U10745 (N_10745,N_7407,N_7326);
nor U10746 (N_10746,N_7987,N_7890);
nor U10747 (N_10747,N_8733,N_8210);
nand U10748 (N_10748,N_6725,N_8314);
and U10749 (N_10749,N_7764,N_7567);
nor U10750 (N_10750,N_8181,N_7619);
or U10751 (N_10751,N_7932,N_6721);
or U10752 (N_10752,N_7967,N_6915);
nand U10753 (N_10753,N_7349,N_6102);
or U10754 (N_10754,N_6637,N_7588);
or U10755 (N_10755,N_6470,N_7191);
and U10756 (N_10756,N_8712,N_8372);
nand U10757 (N_10757,N_8446,N_7781);
or U10758 (N_10758,N_7671,N_8203);
or U10759 (N_10759,N_7357,N_6672);
xor U10760 (N_10760,N_6396,N_7200);
nand U10761 (N_10761,N_8362,N_8722);
or U10762 (N_10762,N_6292,N_8073);
or U10763 (N_10763,N_8270,N_8104);
nand U10764 (N_10764,N_7661,N_8121);
nor U10765 (N_10765,N_8465,N_7981);
or U10766 (N_10766,N_7172,N_6253);
nand U10767 (N_10767,N_6392,N_7306);
or U10768 (N_10768,N_8140,N_8742);
or U10769 (N_10769,N_8627,N_6610);
or U10770 (N_10770,N_7738,N_8819);
xnor U10771 (N_10771,N_6314,N_7431);
xnor U10772 (N_10772,N_8082,N_8004);
and U10773 (N_10773,N_8632,N_7339);
nand U10774 (N_10774,N_8236,N_8349);
nor U10775 (N_10775,N_6709,N_6047);
or U10776 (N_10776,N_8448,N_7912);
or U10777 (N_10777,N_7821,N_7258);
nor U10778 (N_10778,N_6951,N_8919);
nor U10779 (N_10779,N_7883,N_7044);
or U10780 (N_10780,N_8300,N_6489);
and U10781 (N_10781,N_7277,N_7087);
xor U10782 (N_10782,N_8124,N_8560);
and U10783 (N_10783,N_6395,N_7661);
and U10784 (N_10784,N_8207,N_7329);
or U10785 (N_10785,N_7074,N_7305);
nand U10786 (N_10786,N_7540,N_8480);
nor U10787 (N_10787,N_8703,N_6826);
xor U10788 (N_10788,N_7254,N_8679);
nor U10789 (N_10789,N_8575,N_6590);
xnor U10790 (N_10790,N_8998,N_8494);
and U10791 (N_10791,N_6592,N_6694);
xnor U10792 (N_10792,N_6086,N_7455);
or U10793 (N_10793,N_6009,N_6371);
or U10794 (N_10794,N_8229,N_7118);
nor U10795 (N_10795,N_8320,N_7418);
nor U10796 (N_10796,N_7961,N_6024);
xnor U10797 (N_10797,N_6507,N_6257);
and U10798 (N_10798,N_6241,N_8078);
nor U10799 (N_10799,N_6836,N_7248);
and U10800 (N_10800,N_8061,N_8480);
and U10801 (N_10801,N_6727,N_7987);
nand U10802 (N_10802,N_8283,N_6655);
and U10803 (N_10803,N_6983,N_6599);
xor U10804 (N_10804,N_8862,N_7705);
or U10805 (N_10805,N_7970,N_6206);
nor U10806 (N_10806,N_6009,N_8602);
or U10807 (N_10807,N_6244,N_6438);
or U10808 (N_10808,N_6975,N_7308);
and U10809 (N_10809,N_6390,N_8516);
and U10810 (N_10810,N_6251,N_8286);
nor U10811 (N_10811,N_6078,N_6545);
and U10812 (N_10812,N_6764,N_6468);
nor U10813 (N_10813,N_8438,N_6171);
or U10814 (N_10814,N_6113,N_8267);
nand U10815 (N_10815,N_8756,N_8058);
nand U10816 (N_10816,N_8087,N_7744);
xnor U10817 (N_10817,N_7720,N_7920);
nand U10818 (N_10818,N_8876,N_7120);
xnor U10819 (N_10819,N_8906,N_6554);
and U10820 (N_10820,N_8432,N_7049);
nand U10821 (N_10821,N_8072,N_8212);
and U10822 (N_10822,N_7854,N_7596);
and U10823 (N_10823,N_7011,N_8686);
nor U10824 (N_10824,N_8191,N_7690);
and U10825 (N_10825,N_8754,N_7533);
and U10826 (N_10826,N_8008,N_7919);
or U10827 (N_10827,N_8304,N_8510);
nand U10828 (N_10828,N_8818,N_8848);
or U10829 (N_10829,N_8511,N_7912);
nor U10830 (N_10830,N_7232,N_6505);
nand U10831 (N_10831,N_6629,N_7254);
and U10832 (N_10832,N_7907,N_6434);
nand U10833 (N_10833,N_8824,N_7461);
nand U10834 (N_10834,N_6528,N_7807);
or U10835 (N_10835,N_8825,N_7084);
nand U10836 (N_10836,N_7959,N_7667);
or U10837 (N_10837,N_7352,N_6124);
nor U10838 (N_10838,N_8636,N_6080);
nand U10839 (N_10839,N_7383,N_6821);
nor U10840 (N_10840,N_7781,N_7582);
and U10841 (N_10841,N_8082,N_7393);
nor U10842 (N_10842,N_7855,N_7942);
or U10843 (N_10843,N_8844,N_7273);
or U10844 (N_10844,N_6269,N_8594);
xor U10845 (N_10845,N_8953,N_8777);
or U10846 (N_10846,N_6085,N_8754);
and U10847 (N_10847,N_6978,N_8551);
nand U10848 (N_10848,N_7490,N_7094);
or U10849 (N_10849,N_8620,N_7859);
nor U10850 (N_10850,N_7994,N_8549);
nand U10851 (N_10851,N_8411,N_7719);
and U10852 (N_10852,N_6112,N_8785);
nor U10853 (N_10853,N_7965,N_6959);
nor U10854 (N_10854,N_7252,N_7274);
and U10855 (N_10855,N_6526,N_6384);
xor U10856 (N_10856,N_7580,N_7402);
nor U10857 (N_10857,N_8042,N_6389);
or U10858 (N_10858,N_8255,N_8044);
xor U10859 (N_10859,N_6172,N_6822);
and U10860 (N_10860,N_8923,N_6195);
and U10861 (N_10861,N_8793,N_6251);
xor U10862 (N_10862,N_7047,N_8994);
nor U10863 (N_10863,N_7592,N_8539);
xnor U10864 (N_10864,N_6639,N_8794);
nor U10865 (N_10865,N_6822,N_8048);
or U10866 (N_10866,N_8217,N_8254);
nand U10867 (N_10867,N_7009,N_7981);
xnor U10868 (N_10868,N_7422,N_7207);
xnor U10869 (N_10869,N_6710,N_6656);
nand U10870 (N_10870,N_8634,N_6915);
nor U10871 (N_10871,N_7817,N_8640);
nor U10872 (N_10872,N_6033,N_8124);
xnor U10873 (N_10873,N_7136,N_7407);
xnor U10874 (N_10874,N_6839,N_7964);
nand U10875 (N_10875,N_8501,N_6918);
nor U10876 (N_10876,N_6966,N_6339);
or U10877 (N_10877,N_7455,N_7317);
or U10878 (N_10878,N_8169,N_6547);
xor U10879 (N_10879,N_6497,N_6219);
and U10880 (N_10880,N_7396,N_6721);
or U10881 (N_10881,N_8541,N_8605);
nand U10882 (N_10882,N_6973,N_7569);
nand U10883 (N_10883,N_7384,N_6266);
and U10884 (N_10884,N_7824,N_6651);
and U10885 (N_10885,N_7383,N_7514);
and U10886 (N_10886,N_6739,N_7723);
nand U10887 (N_10887,N_8080,N_7555);
xor U10888 (N_10888,N_7844,N_7105);
nand U10889 (N_10889,N_7173,N_8220);
nand U10890 (N_10890,N_7190,N_7222);
and U10891 (N_10891,N_6912,N_7135);
or U10892 (N_10892,N_7832,N_8846);
xor U10893 (N_10893,N_7003,N_8265);
nand U10894 (N_10894,N_6268,N_6181);
nand U10895 (N_10895,N_8537,N_7582);
nor U10896 (N_10896,N_8465,N_7911);
xnor U10897 (N_10897,N_8694,N_6203);
nor U10898 (N_10898,N_8439,N_7930);
or U10899 (N_10899,N_6044,N_8139);
nand U10900 (N_10900,N_6540,N_6979);
or U10901 (N_10901,N_7611,N_6133);
xor U10902 (N_10902,N_6255,N_6130);
and U10903 (N_10903,N_6101,N_7660);
or U10904 (N_10904,N_6974,N_6454);
nand U10905 (N_10905,N_6591,N_8243);
xor U10906 (N_10906,N_7063,N_7650);
nand U10907 (N_10907,N_7380,N_7953);
and U10908 (N_10908,N_7021,N_8831);
or U10909 (N_10909,N_7326,N_6337);
xnor U10910 (N_10910,N_8265,N_6369);
or U10911 (N_10911,N_7678,N_7393);
and U10912 (N_10912,N_8938,N_8324);
and U10913 (N_10913,N_7363,N_7141);
and U10914 (N_10914,N_7163,N_8373);
or U10915 (N_10915,N_6064,N_7911);
nor U10916 (N_10916,N_6236,N_7972);
and U10917 (N_10917,N_6254,N_8198);
xor U10918 (N_10918,N_6064,N_6932);
and U10919 (N_10919,N_7994,N_6924);
or U10920 (N_10920,N_7262,N_6153);
or U10921 (N_10921,N_8067,N_7472);
nand U10922 (N_10922,N_7259,N_8390);
nor U10923 (N_10923,N_7213,N_8815);
and U10924 (N_10924,N_6119,N_6434);
or U10925 (N_10925,N_8282,N_8081);
nor U10926 (N_10926,N_7741,N_8251);
nor U10927 (N_10927,N_7000,N_6606);
or U10928 (N_10928,N_8241,N_7858);
or U10929 (N_10929,N_8477,N_8324);
nand U10930 (N_10930,N_8725,N_7204);
xnor U10931 (N_10931,N_7280,N_7367);
xnor U10932 (N_10932,N_7507,N_7888);
nand U10933 (N_10933,N_6607,N_7875);
nor U10934 (N_10934,N_8216,N_7667);
xor U10935 (N_10935,N_8081,N_6204);
nor U10936 (N_10936,N_8958,N_7770);
nor U10937 (N_10937,N_7367,N_8454);
nor U10938 (N_10938,N_8910,N_7203);
and U10939 (N_10939,N_6816,N_8683);
or U10940 (N_10940,N_8166,N_7422);
xnor U10941 (N_10941,N_8696,N_8068);
nor U10942 (N_10942,N_8231,N_7022);
or U10943 (N_10943,N_7340,N_7302);
nand U10944 (N_10944,N_6843,N_8054);
nor U10945 (N_10945,N_7823,N_8459);
nand U10946 (N_10946,N_7787,N_7019);
nand U10947 (N_10947,N_6296,N_7380);
xnor U10948 (N_10948,N_7666,N_6130);
nor U10949 (N_10949,N_6671,N_8339);
or U10950 (N_10950,N_7800,N_8168);
and U10951 (N_10951,N_7941,N_7318);
xnor U10952 (N_10952,N_6083,N_6318);
and U10953 (N_10953,N_6418,N_7526);
xor U10954 (N_10954,N_6102,N_6765);
nor U10955 (N_10955,N_7354,N_6875);
xnor U10956 (N_10956,N_8467,N_6285);
and U10957 (N_10957,N_8816,N_6309);
and U10958 (N_10958,N_7582,N_7695);
and U10959 (N_10959,N_8018,N_7521);
nand U10960 (N_10960,N_6443,N_8408);
or U10961 (N_10961,N_6626,N_6670);
or U10962 (N_10962,N_8827,N_8215);
and U10963 (N_10963,N_7489,N_8378);
nor U10964 (N_10964,N_8946,N_6981);
and U10965 (N_10965,N_7536,N_8441);
nor U10966 (N_10966,N_7372,N_7459);
nand U10967 (N_10967,N_6859,N_7116);
and U10968 (N_10968,N_7741,N_7739);
and U10969 (N_10969,N_8818,N_6364);
nor U10970 (N_10970,N_7480,N_7834);
xnor U10971 (N_10971,N_8052,N_8679);
nor U10972 (N_10972,N_7074,N_7478);
nor U10973 (N_10973,N_6364,N_6806);
nand U10974 (N_10974,N_6740,N_8524);
and U10975 (N_10975,N_6737,N_6237);
nor U10976 (N_10976,N_7801,N_7471);
nand U10977 (N_10977,N_6539,N_6435);
nand U10978 (N_10978,N_8688,N_7685);
or U10979 (N_10979,N_6940,N_7409);
nor U10980 (N_10980,N_8368,N_8871);
nor U10981 (N_10981,N_8226,N_8286);
nand U10982 (N_10982,N_6716,N_8090);
xnor U10983 (N_10983,N_7728,N_7298);
xnor U10984 (N_10984,N_8698,N_6566);
or U10985 (N_10985,N_8111,N_7157);
and U10986 (N_10986,N_7776,N_8248);
nor U10987 (N_10987,N_8515,N_7274);
nor U10988 (N_10988,N_7330,N_6057);
nor U10989 (N_10989,N_7103,N_6025);
nand U10990 (N_10990,N_8739,N_7261);
nor U10991 (N_10991,N_8941,N_6802);
nor U10992 (N_10992,N_8291,N_8205);
or U10993 (N_10993,N_7104,N_8136);
or U10994 (N_10994,N_6717,N_6964);
and U10995 (N_10995,N_7428,N_6161);
or U10996 (N_10996,N_7588,N_6031);
and U10997 (N_10997,N_6457,N_6948);
xor U10998 (N_10998,N_7535,N_7558);
nor U10999 (N_10999,N_7750,N_8866);
nor U11000 (N_11000,N_7700,N_6981);
xnor U11001 (N_11001,N_8082,N_8431);
xnor U11002 (N_11002,N_8964,N_7113);
xnor U11003 (N_11003,N_6415,N_7900);
and U11004 (N_11004,N_7926,N_8453);
nor U11005 (N_11005,N_6981,N_6581);
nor U11006 (N_11006,N_6504,N_7098);
or U11007 (N_11007,N_6689,N_7484);
xor U11008 (N_11008,N_6337,N_7134);
nand U11009 (N_11009,N_8444,N_8325);
xor U11010 (N_11010,N_8997,N_6268);
and U11011 (N_11011,N_7206,N_6226);
nor U11012 (N_11012,N_6003,N_8377);
nand U11013 (N_11013,N_8065,N_8199);
and U11014 (N_11014,N_6413,N_7641);
and U11015 (N_11015,N_7851,N_6625);
or U11016 (N_11016,N_7344,N_8198);
xnor U11017 (N_11017,N_7846,N_6119);
xor U11018 (N_11018,N_7322,N_8420);
xnor U11019 (N_11019,N_6522,N_6964);
and U11020 (N_11020,N_6274,N_6275);
xor U11021 (N_11021,N_8055,N_6185);
and U11022 (N_11022,N_8084,N_7140);
nand U11023 (N_11023,N_6192,N_8743);
and U11024 (N_11024,N_8017,N_8159);
nor U11025 (N_11025,N_6884,N_7641);
nand U11026 (N_11026,N_8149,N_8106);
xnor U11027 (N_11027,N_6074,N_8756);
and U11028 (N_11028,N_8254,N_7986);
nand U11029 (N_11029,N_7940,N_8067);
xor U11030 (N_11030,N_6817,N_7056);
xnor U11031 (N_11031,N_6889,N_8504);
or U11032 (N_11032,N_8746,N_8468);
nor U11033 (N_11033,N_6840,N_7575);
nor U11034 (N_11034,N_6986,N_6904);
or U11035 (N_11035,N_6831,N_7484);
nand U11036 (N_11036,N_6930,N_8588);
nor U11037 (N_11037,N_7474,N_6408);
or U11038 (N_11038,N_7288,N_7172);
and U11039 (N_11039,N_6575,N_6263);
and U11040 (N_11040,N_7810,N_7582);
nor U11041 (N_11041,N_6256,N_7328);
nor U11042 (N_11042,N_7571,N_7676);
xnor U11043 (N_11043,N_7416,N_8352);
and U11044 (N_11044,N_7772,N_7962);
nand U11045 (N_11045,N_7728,N_6818);
xor U11046 (N_11046,N_8450,N_7322);
xnor U11047 (N_11047,N_7725,N_6831);
and U11048 (N_11048,N_6136,N_8512);
nor U11049 (N_11049,N_6947,N_7813);
and U11050 (N_11050,N_6943,N_7999);
nand U11051 (N_11051,N_8366,N_7343);
or U11052 (N_11052,N_6512,N_7154);
and U11053 (N_11053,N_8735,N_8009);
nand U11054 (N_11054,N_7269,N_7532);
nand U11055 (N_11055,N_7835,N_8253);
xor U11056 (N_11056,N_7401,N_6423);
or U11057 (N_11057,N_8445,N_7920);
nand U11058 (N_11058,N_6255,N_6960);
nor U11059 (N_11059,N_8236,N_8820);
xor U11060 (N_11060,N_6536,N_7947);
nand U11061 (N_11061,N_7471,N_8107);
xor U11062 (N_11062,N_8080,N_8903);
xor U11063 (N_11063,N_8144,N_7140);
or U11064 (N_11064,N_6120,N_6654);
nor U11065 (N_11065,N_7828,N_7813);
and U11066 (N_11066,N_7008,N_6681);
and U11067 (N_11067,N_6036,N_6570);
nand U11068 (N_11068,N_8857,N_7164);
nand U11069 (N_11069,N_8633,N_8026);
and U11070 (N_11070,N_6315,N_7957);
or U11071 (N_11071,N_7757,N_7304);
nand U11072 (N_11072,N_8266,N_7163);
nor U11073 (N_11073,N_7035,N_6245);
xnor U11074 (N_11074,N_8544,N_7982);
nand U11075 (N_11075,N_8695,N_6256);
xor U11076 (N_11076,N_8482,N_7299);
or U11077 (N_11077,N_6576,N_8922);
xnor U11078 (N_11078,N_8148,N_7566);
or U11079 (N_11079,N_7694,N_7539);
or U11080 (N_11080,N_8034,N_6395);
nor U11081 (N_11081,N_8942,N_6259);
xnor U11082 (N_11082,N_6564,N_7587);
and U11083 (N_11083,N_6095,N_7190);
nand U11084 (N_11084,N_8379,N_8480);
or U11085 (N_11085,N_6199,N_8461);
and U11086 (N_11086,N_8739,N_6741);
or U11087 (N_11087,N_6510,N_6492);
xnor U11088 (N_11088,N_7631,N_8654);
and U11089 (N_11089,N_8756,N_6014);
nor U11090 (N_11090,N_6758,N_8453);
nand U11091 (N_11091,N_7082,N_8174);
and U11092 (N_11092,N_7137,N_7647);
or U11093 (N_11093,N_8550,N_7178);
and U11094 (N_11094,N_8664,N_6758);
and U11095 (N_11095,N_6446,N_7518);
nor U11096 (N_11096,N_6431,N_8606);
nand U11097 (N_11097,N_8381,N_7052);
nand U11098 (N_11098,N_7439,N_7876);
and U11099 (N_11099,N_7491,N_6528);
nand U11100 (N_11100,N_7881,N_7788);
xnor U11101 (N_11101,N_6948,N_6016);
xnor U11102 (N_11102,N_6871,N_6955);
xnor U11103 (N_11103,N_7395,N_6191);
and U11104 (N_11104,N_6959,N_7494);
or U11105 (N_11105,N_7285,N_6010);
or U11106 (N_11106,N_8059,N_7718);
or U11107 (N_11107,N_8267,N_6037);
xnor U11108 (N_11108,N_7230,N_7566);
nor U11109 (N_11109,N_7302,N_8130);
nor U11110 (N_11110,N_7064,N_7971);
nand U11111 (N_11111,N_6350,N_8319);
or U11112 (N_11112,N_7301,N_6177);
or U11113 (N_11113,N_8606,N_8170);
and U11114 (N_11114,N_6314,N_7448);
xnor U11115 (N_11115,N_6812,N_6070);
xor U11116 (N_11116,N_7819,N_7741);
or U11117 (N_11117,N_7358,N_7036);
nor U11118 (N_11118,N_6282,N_8228);
and U11119 (N_11119,N_8415,N_8269);
or U11120 (N_11120,N_7368,N_8900);
nor U11121 (N_11121,N_7550,N_6316);
xor U11122 (N_11122,N_6819,N_7226);
or U11123 (N_11123,N_8891,N_7680);
xor U11124 (N_11124,N_8633,N_6555);
or U11125 (N_11125,N_7276,N_6499);
nor U11126 (N_11126,N_6703,N_7009);
nand U11127 (N_11127,N_7233,N_8903);
xnor U11128 (N_11128,N_8135,N_6392);
nand U11129 (N_11129,N_6982,N_8417);
xor U11130 (N_11130,N_8124,N_8534);
and U11131 (N_11131,N_8766,N_6379);
or U11132 (N_11132,N_6883,N_7982);
nand U11133 (N_11133,N_7909,N_7309);
xor U11134 (N_11134,N_6151,N_8764);
nor U11135 (N_11135,N_6243,N_6542);
xor U11136 (N_11136,N_8669,N_8366);
or U11137 (N_11137,N_6942,N_7668);
nor U11138 (N_11138,N_7257,N_6371);
and U11139 (N_11139,N_6016,N_7667);
xnor U11140 (N_11140,N_8339,N_6856);
and U11141 (N_11141,N_8749,N_7495);
or U11142 (N_11142,N_6137,N_8618);
nor U11143 (N_11143,N_8748,N_8373);
and U11144 (N_11144,N_7734,N_8042);
nand U11145 (N_11145,N_7780,N_6238);
nor U11146 (N_11146,N_6453,N_6581);
nor U11147 (N_11147,N_6679,N_7197);
nand U11148 (N_11148,N_6246,N_6298);
nand U11149 (N_11149,N_7764,N_7231);
or U11150 (N_11150,N_6112,N_6638);
and U11151 (N_11151,N_7406,N_6194);
and U11152 (N_11152,N_7244,N_6192);
and U11153 (N_11153,N_6134,N_6648);
xor U11154 (N_11154,N_6186,N_6921);
nand U11155 (N_11155,N_6155,N_7828);
nand U11156 (N_11156,N_7654,N_6669);
or U11157 (N_11157,N_7534,N_7177);
nand U11158 (N_11158,N_6915,N_6174);
or U11159 (N_11159,N_8953,N_8197);
and U11160 (N_11160,N_6744,N_6476);
and U11161 (N_11161,N_8177,N_6480);
xor U11162 (N_11162,N_7378,N_6985);
nor U11163 (N_11163,N_6497,N_6851);
nand U11164 (N_11164,N_6691,N_7538);
and U11165 (N_11165,N_8492,N_8135);
nand U11166 (N_11166,N_7826,N_7486);
and U11167 (N_11167,N_6703,N_8178);
or U11168 (N_11168,N_6356,N_7792);
xnor U11169 (N_11169,N_8338,N_8321);
or U11170 (N_11170,N_7431,N_8976);
nand U11171 (N_11171,N_7300,N_6177);
and U11172 (N_11172,N_6295,N_6636);
and U11173 (N_11173,N_8145,N_6814);
xor U11174 (N_11174,N_7776,N_6160);
xnor U11175 (N_11175,N_7515,N_8801);
nor U11176 (N_11176,N_7486,N_6733);
nand U11177 (N_11177,N_7680,N_6900);
nor U11178 (N_11178,N_7478,N_6596);
nor U11179 (N_11179,N_7663,N_8412);
nor U11180 (N_11180,N_8282,N_6014);
and U11181 (N_11181,N_6812,N_7886);
or U11182 (N_11182,N_8436,N_6424);
nand U11183 (N_11183,N_7295,N_7870);
xor U11184 (N_11184,N_6254,N_7529);
xnor U11185 (N_11185,N_6231,N_8700);
or U11186 (N_11186,N_8311,N_8871);
nand U11187 (N_11187,N_7202,N_6961);
nand U11188 (N_11188,N_7766,N_7453);
xnor U11189 (N_11189,N_7002,N_6927);
and U11190 (N_11190,N_8005,N_6861);
or U11191 (N_11191,N_8414,N_7305);
nand U11192 (N_11192,N_7054,N_8556);
or U11193 (N_11193,N_8989,N_6191);
and U11194 (N_11194,N_6105,N_7363);
or U11195 (N_11195,N_7387,N_7242);
and U11196 (N_11196,N_7974,N_8754);
and U11197 (N_11197,N_6336,N_7111);
xor U11198 (N_11198,N_8125,N_8841);
nand U11199 (N_11199,N_7663,N_8049);
nand U11200 (N_11200,N_8226,N_7595);
nand U11201 (N_11201,N_6050,N_7572);
or U11202 (N_11202,N_6401,N_6244);
or U11203 (N_11203,N_6398,N_7975);
and U11204 (N_11204,N_6968,N_7349);
xnor U11205 (N_11205,N_8526,N_8708);
nand U11206 (N_11206,N_6488,N_8899);
and U11207 (N_11207,N_8299,N_8607);
nand U11208 (N_11208,N_6820,N_7063);
nor U11209 (N_11209,N_8094,N_7056);
nor U11210 (N_11210,N_6550,N_8690);
and U11211 (N_11211,N_8470,N_7961);
nand U11212 (N_11212,N_6601,N_8472);
nor U11213 (N_11213,N_7057,N_6718);
or U11214 (N_11214,N_8783,N_7786);
or U11215 (N_11215,N_6600,N_7023);
xor U11216 (N_11216,N_6853,N_8794);
or U11217 (N_11217,N_6392,N_6800);
and U11218 (N_11218,N_8607,N_6080);
or U11219 (N_11219,N_7453,N_7783);
or U11220 (N_11220,N_8556,N_7794);
or U11221 (N_11221,N_6784,N_8846);
nand U11222 (N_11222,N_8071,N_6732);
xor U11223 (N_11223,N_8546,N_6555);
or U11224 (N_11224,N_6636,N_6082);
and U11225 (N_11225,N_6140,N_7493);
nor U11226 (N_11226,N_8292,N_8408);
and U11227 (N_11227,N_6782,N_8248);
or U11228 (N_11228,N_8800,N_8105);
nor U11229 (N_11229,N_7796,N_7968);
nor U11230 (N_11230,N_7450,N_8453);
xnor U11231 (N_11231,N_8505,N_7791);
nor U11232 (N_11232,N_6117,N_6489);
or U11233 (N_11233,N_6956,N_7796);
and U11234 (N_11234,N_6888,N_8261);
xor U11235 (N_11235,N_8118,N_8856);
nor U11236 (N_11236,N_7786,N_7422);
nor U11237 (N_11237,N_7160,N_7689);
nor U11238 (N_11238,N_8399,N_6424);
xor U11239 (N_11239,N_8241,N_6036);
nand U11240 (N_11240,N_7842,N_8132);
xnor U11241 (N_11241,N_6780,N_6118);
nand U11242 (N_11242,N_6059,N_8309);
or U11243 (N_11243,N_6770,N_6048);
and U11244 (N_11244,N_6808,N_6508);
or U11245 (N_11245,N_7691,N_6090);
nand U11246 (N_11246,N_8900,N_7740);
nor U11247 (N_11247,N_6734,N_7564);
xnor U11248 (N_11248,N_6680,N_8856);
or U11249 (N_11249,N_8114,N_7684);
or U11250 (N_11250,N_8847,N_6212);
nand U11251 (N_11251,N_7216,N_7753);
and U11252 (N_11252,N_6147,N_8856);
nor U11253 (N_11253,N_7665,N_8085);
and U11254 (N_11254,N_8273,N_7928);
nand U11255 (N_11255,N_8159,N_7461);
xor U11256 (N_11256,N_8853,N_6755);
or U11257 (N_11257,N_7736,N_7438);
xnor U11258 (N_11258,N_8944,N_6957);
and U11259 (N_11259,N_6010,N_8721);
or U11260 (N_11260,N_7832,N_6217);
xnor U11261 (N_11261,N_6215,N_7654);
xnor U11262 (N_11262,N_8292,N_6895);
or U11263 (N_11263,N_6018,N_6320);
nand U11264 (N_11264,N_8197,N_6307);
or U11265 (N_11265,N_8008,N_7373);
or U11266 (N_11266,N_6023,N_7078);
and U11267 (N_11267,N_7662,N_7233);
nand U11268 (N_11268,N_8237,N_8244);
nand U11269 (N_11269,N_8529,N_6463);
and U11270 (N_11270,N_7270,N_6383);
nor U11271 (N_11271,N_6248,N_7532);
nor U11272 (N_11272,N_7025,N_6208);
xnor U11273 (N_11273,N_7529,N_8749);
or U11274 (N_11274,N_8927,N_6028);
nand U11275 (N_11275,N_7654,N_8247);
nand U11276 (N_11276,N_8220,N_8192);
and U11277 (N_11277,N_6005,N_8232);
xnor U11278 (N_11278,N_8960,N_6770);
nand U11279 (N_11279,N_7056,N_6591);
and U11280 (N_11280,N_6953,N_6187);
or U11281 (N_11281,N_7349,N_8040);
or U11282 (N_11282,N_6183,N_8324);
or U11283 (N_11283,N_8511,N_6363);
xnor U11284 (N_11284,N_8456,N_6794);
nor U11285 (N_11285,N_6762,N_6588);
nor U11286 (N_11286,N_7195,N_8647);
or U11287 (N_11287,N_8967,N_7794);
nand U11288 (N_11288,N_7368,N_6229);
or U11289 (N_11289,N_7820,N_8594);
xnor U11290 (N_11290,N_6670,N_6620);
xnor U11291 (N_11291,N_8506,N_7677);
xor U11292 (N_11292,N_8181,N_6697);
or U11293 (N_11293,N_7736,N_6694);
nand U11294 (N_11294,N_7113,N_7645);
nor U11295 (N_11295,N_6908,N_8109);
or U11296 (N_11296,N_6390,N_7762);
xnor U11297 (N_11297,N_6993,N_6329);
and U11298 (N_11298,N_7719,N_8897);
or U11299 (N_11299,N_7917,N_8263);
xnor U11300 (N_11300,N_7891,N_7807);
nor U11301 (N_11301,N_6010,N_6181);
nor U11302 (N_11302,N_8087,N_6780);
nor U11303 (N_11303,N_8384,N_8365);
nand U11304 (N_11304,N_8360,N_8524);
and U11305 (N_11305,N_7501,N_8617);
nand U11306 (N_11306,N_6861,N_6492);
nor U11307 (N_11307,N_6317,N_7968);
nand U11308 (N_11308,N_6043,N_6290);
or U11309 (N_11309,N_8897,N_6830);
and U11310 (N_11310,N_7195,N_7827);
nand U11311 (N_11311,N_8735,N_8234);
or U11312 (N_11312,N_8080,N_6281);
xor U11313 (N_11313,N_7358,N_6580);
and U11314 (N_11314,N_7763,N_8603);
or U11315 (N_11315,N_8232,N_6814);
or U11316 (N_11316,N_7688,N_8971);
and U11317 (N_11317,N_8786,N_8159);
xor U11318 (N_11318,N_7164,N_6314);
nand U11319 (N_11319,N_8366,N_8512);
nand U11320 (N_11320,N_8657,N_7871);
nor U11321 (N_11321,N_7602,N_6889);
or U11322 (N_11322,N_7517,N_6008);
nor U11323 (N_11323,N_6082,N_7122);
xor U11324 (N_11324,N_6220,N_6694);
nand U11325 (N_11325,N_7976,N_7843);
nor U11326 (N_11326,N_8121,N_7146);
nand U11327 (N_11327,N_7078,N_7734);
nor U11328 (N_11328,N_8418,N_6703);
and U11329 (N_11329,N_7298,N_7980);
nand U11330 (N_11330,N_6710,N_8216);
or U11331 (N_11331,N_8653,N_6023);
xor U11332 (N_11332,N_6000,N_8595);
nand U11333 (N_11333,N_7005,N_6182);
nand U11334 (N_11334,N_6798,N_7791);
or U11335 (N_11335,N_7639,N_7588);
or U11336 (N_11336,N_8593,N_7448);
or U11337 (N_11337,N_7861,N_8236);
and U11338 (N_11338,N_7045,N_8505);
or U11339 (N_11339,N_8518,N_7598);
and U11340 (N_11340,N_8009,N_6040);
xnor U11341 (N_11341,N_8393,N_7178);
nor U11342 (N_11342,N_7227,N_7487);
and U11343 (N_11343,N_8123,N_8365);
nor U11344 (N_11344,N_8698,N_7838);
or U11345 (N_11345,N_8839,N_6739);
or U11346 (N_11346,N_6738,N_6511);
nand U11347 (N_11347,N_6746,N_8035);
nand U11348 (N_11348,N_7065,N_6272);
nand U11349 (N_11349,N_7471,N_6447);
and U11350 (N_11350,N_6301,N_7764);
nand U11351 (N_11351,N_6557,N_8354);
xnor U11352 (N_11352,N_7999,N_6229);
xnor U11353 (N_11353,N_8431,N_6413);
or U11354 (N_11354,N_7295,N_8453);
and U11355 (N_11355,N_6975,N_7656);
or U11356 (N_11356,N_7194,N_6595);
and U11357 (N_11357,N_6681,N_7096);
and U11358 (N_11358,N_7296,N_8880);
nand U11359 (N_11359,N_6108,N_7959);
nor U11360 (N_11360,N_7342,N_7981);
nor U11361 (N_11361,N_7259,N_6078);
nor U11362 (N_11362,N_6240,N_8505);
xnor U11363 (N_11363,N_8195,N_6373);
and U11364 (N_11364,N_8591,N_7167);
and U11365 (N_11365,N_8447,N_7188);
xor U11366 (N_11366,N_8710,N_7889);
nand U11367 (N_11367,N_6531,N_8609);
nor U11368 (N_11368,N_6568,N_6828);
xnor U11369 (N_11369,N_8697,N_7717);
and U11370 (N_11370,N_6015,N_7787);
or U11371 (N_11371,N_8743,N_7187);
nor U11372 (N_11372,N_8611,N_6207);
or U11373 (N_11373,N_7633,N_8035);
xor U11374 (N_11374,N_6991,N_7633);
or U11375 (N_11375,N_6937,N_6383);
xnor U11376 (N_11376,N_6561,N_8646);
and U11377 (N_11377,N_8238,N_6156);
nand U11378 (N_11378,N_8934,N_7053);
nand U11379 (N_11379,N_8247,N_8103);
and U11380 (N_11380,N_7879,N_6545);
and U11381 (N_11381,N_8009,N_6893);
and U11382 (N_11382,N_6788,N_6643);
nand U11383 (N_11383,N_6398,N_7601);
nand U11384 (N_11384,N_8727,N_7288);
xnor U11385 (N_11385,N_8525,N_6912);
or U11386 (N_11386,N_6024,N_6780);
xor U11387 (N_11387,N_7385,N_6517);
nor U11388 (N_11388,N_8205,N_8790);
nand U11389 (N_11389,N_8183,N_6400);
nand U11390 (N_11390,N_6845,N_8712);
nand U11391 (N_11391,N_6436,N_8623);
xor U11392 (N_11392,N_8240,N_7385);
nand U11393 (N_11393,N_8218,N_7184);
xor U11394 (N_11394,N_7520,N_7336);
and U11395 (N_11395,N_8403,N_6131);
nand U11396 (N_11396,N_6190,N_6462);
and U11397 (N_11397,N_6697,N_7581);
nor U11398 (N_11398,N_7252,N_6364);
xnor U11399 (N_11399,N_7810,N_8059);
or U11400 (N_11400,N_6804,N_7868);
and U11401 (N_11401,N_6151,N_6357);
nor U11402 (N_11402,N_6066,N_6958);
nor U11403 (N_11403,N_6111,N_6582);
or U11404 (N_11404,N_6310,N_6331);
xnor U11405 (N_11405,N_7529,N_8845);
or U11406 (N_11406,N_8084,N_7854);
nand U11407 (N_11407,N_8680,N_6273);
and U11408 (N_11408,N_6843,N_7871);
nor U11409 (N_11409,N_6424,N_7493);
xor U11410 (N_11410,N_7745,N_8408);
nand U11411 (N_11411,N_6978,N_7265);
and U11412 (N_11412,N_8758,N_6748);
nor U11413 (N_11413,N_7687,N_6060);
or U11414 (N_11414,N_6324,N_7729);
xor U11415 (N_11415,N_8564,N_6330);
nor U11416 (N_11416,N_7344,N_8892);
nand U11417 (N_11417,N_6689,N_8124);
and U11418 (N_11418,N_6442,N_6923);
or U11419 (N_11419,N_8967,N_7524);
xnor U11420 (N_11420,N_6140,N_8198);
or U11421 (N_11421,N_7882,N_7725);
nand U11422 (N_11422,N_7298,N_7519);
or U11423 (N_11423,N_7274,N_7352);
nand U11424 (N_11424,N_7621,N_7313);
nand U11425 (N_11425,N_7393,N_6963);
or U11426 (N_11426,N_8235,N_7070);
xnor U11427 (N_11427,N_6306,N_6489);
nor U11428 (N_11428,N_7179,N_6527);
and U11429 (N_11429,N_8167,N_8386);
nor U11430 (N_11430,N_7262,N_8393);
xor U11431 (N_11431,N_6958,N_6987);
and U11432 (N_11432,N_6582,N_8761);
nor U11433 (N_11433,N_6645,N_8731);
and U11434 (N_11434,N_7411,N_6743);
and U11435 (N_11435,N_7387,N_7634);
nand U11436 (N_11436,N_8966,N_8429);
xor U11437 (N_11437,N_8767,N_8061);
nand U11438 (N_11438,N_8092,N_6376);
or U11439 (N_11439,N_8252,N_7455);
or U11440 (N_11440,N_8180,N_6381);
or U11441 (N_11441,N_6627,N_6222);
nor U11442 (N_11442,N_6336,N_8839);
nor U11443 (N_11443,N_8143,N_6953);
nand U11444 (N_11444,N_6047,N_7975);
nor U11445 (N_11445,N_6779,N_6407);
and U11446 (N_11446,N_8851,N_7595);
nor U11447 (N_11447,N_6277,N_6663);
or U11448 (N_11448,N_7969,N_7941);
and U11449 (N_11449,N_7109,N_6458);
or U11450 (N_11450,N_7336,N_6169);
and U11451 (N_11451,N_7647,N_6976);
or U11452 (N_11452,N_7835,N_7787);
xor U11453 (N_11453,N_7398,N_6041);
nand U11454 (N_11454,N_8847,N_7618);
xor U11455 (N_11455,N_6653,N_6305);
nand U11456 (N_11456,N_6211,N_6962);
or U11457 (N_11457,N_7519,N_6482);
xnor U11458 (N_11458,N_7530,N_7042);
or U11459 (N_11459,N_7319,N_6074);
nand U11460 (N_11460,N_6498,N_8132);
and U11461 (N_11461,N_8460,N_8879);
nor U11462 (N_11462,N_8483,N_6122);
nor U11463 (N_11463,N_7815,N_8460);
nand U11464 (N_11464,N_6315,N_8969);
xor U11465 (N_11465,N_6927,N_8201);
or U11466 (N_11466,N_6382,N_7555);
xor U11467 (N_11467,N_6840,N_8042);
or U11468 (N_11468,N_6175,N_7158);
or U11469 (N_11469,N_7509,N_7994);
or U11470 (N_11470,N_6612,N_7215);
nor U11471 (N_11471,N_7498,N_7775);
nor U11472 (N_11472,N_7948,N_8781);
or U11473 (N_11473,N_6279,N_6934);
or U11474 (N_11474,N_8435,N_8468);
or U11475 (N_11475,N_6117,N_7798);
xor U11476 (N_11476,N_8968,N_7062);
nand U11477 (N_11477,N_7419,N_8913);
xnor U11478 (N_11478,N_7854,N_8545);
nor U11479 (N_11479,N_8786,N_6665);
xor U11480 (N_11480,N_6222,N_8834);
xnor U11481 (N_11481,N_6904,N_8820);
and U11482 (N_11482,N_6407,N_7432);
nand U11483 (N_11483,N_8612,N_6019);
nor U11484 (N_11484,N_7107,N_6498);
or U11485 (N_11485,N_6152,N_6912);
nand U11486 (N_11486,N_8107,N_6342);
nand U11487 (N_11487,N_7124,N_6118);
xnor U11488 (N_11488,N_7278,N_6573);
nor U11489 (N_11489,N_6428,N_6412);
and U11490 (N_11490,N_6242,N_7522);
xor U11491 (N_11491,N_7279,N_6281);
xor U11492 (N_11492,N_8083,N_6766);
nand U11493 (N_11493,N_7102,N_6193);
xnor U11494 (N_11494,N_8490,N_7916);
nand U11495 (N_11495,N_7764,N_7592);
and U11496 (N_11496,N_6112,N_8450);
nor U11497 (N_11497,N_6859,N_8544);
nor U11498 (N_11498,N_7253,N_6344);
nor U11499 (N_11499,N_7873,N_6248);
nand U11500 (N_11500,N_8776,N_8631);
xnor U11501 (N_11501,N_8012,N_6843);
nand U11502 (N_11502,N_8043,N_8514);
nor U11503 (N_11503,N_6860,N_7699);
xnor U11504 (N_11504,N_7046,N_6753);
nor U11505 (N_11505,N_8851,N_7491);
nand U11506 (N_11506,N_7597,N_6849);
or U11507 (N_11507,N_7532,N_8208);
xor U11508 (N_11508,N_6220,N_8683);
and U11509 (N_11509,N_8290,N_7640);
nor U11510 (N_11510,N_7566,N_6236);
or U11511 (N_11511,N_8786,N_7321);
and U11512 (N_11512,N_8070,N_8268);
nand U11513 (N_11513,N_7310,N_6566);
nand U11514 (N_11514,N_8909,N_7874);
or U11515 (N_11515,N_6827,N_8285);
or U11516 (N_11516,N_7949,N_6129);
or U11517 (N_11517,N_6318,N_6919);
xnor U11518 (N_11518,N_8705,N_7975);
xor U11519 (N_11519,N_6564,N_7064);
nor U11520 (N_11520,N_8869,N_8560);
or U11521 (N_11521,N_7754,N_6773);
or U11522 (N_11522,N_7210,N_8102);
and U11523 (N_11523,N_7381,N_8932);
nand U11524 (N_11524,N_8126,N_8251);
nor U11525 (N_11525,N_6198,N_8113);
xor U11526 (N_11526,N_8103,N_8292);
xor U11527 (N_11527,N_6935,N_8134);
nor U11528 (N_11528,N_8669,N_6620);
and U11529 (N_11529,N_8163,N_8795);
and U11530 (N_11530,N_6516,N_7569);
and U11531 (N_11531,N_6035,N_7782);
and U11532 (N_11532,N_7922,N_7264);
nor U11533 (N_11533,N_8060,N_8845);
nand U11534 (N_11534,N_8580,N_8050);
nand U11535 (N_11535,N_7169,N_8241);
nand U11536 (N_11536,N_8631,N_8572);
nor U11537 (N_11537,N_7186,N_7788);
nor U11538 (N_11538,N_6770,N_7300);
and U11539 (N_11539,N_7940,N_6392);
or U11540 (N_11540,N_7335,N_8506);
or U11541 (N_11541,N_6919,N_7383);
xnor U11542 (N_11542,N_7888,N_8480);
nor U11543 (N_11543,N_7047,N_6431);
and U11544 (N_11544,N_8566,N_7043);
nand U11545 (N_11545,N_6028,N_8922);
and U11546 (N_11546,N_8459,N_8010);
xnor U11547 (N_11547,N_6351,N_7730);
xnor U11548 (N_11548,N_7024,N_8111);
nor U11549 (N_11549,N_8046,N_7091);
nor U11550 (N_11550,N_8820,N_6931);
nand U11551 (N_11551,N_7987,N_7216);
nor U11552 (N_11552,N_8386,N_6398);
and U11553 (N_11553,N_8490,N_6779);
and U11554 (N_11554,N_6577,N_6167);
and U11555 (N_11555,N_8288,N_8846);
or U11556 (N_11556,N_8783,N_6745);
xor U11557 (N_11557,N_7267,N_6374);
nand U11558 (N_11558,N_8355,N_8098);
nor U11559 (N_11559,N_8845,N_7293);
xnor U11560 (N_11560,N_6000,N_8150);
or U11561 (N_11561,N_6262,N_7547);
and U11562 (N_11562,N_8597,N_8952);
and U11563 (N_11563,N_6489,N_8196);
xnor U11564 (N_11564,N_6715,N_7129);
nor U11565 (N_11565,N_6031,N_8497);
and U11566 (N_11566,N_8046,N_8392);
or U11567 (N_11567,N_6151,N_8863);
and U11568 (N_11568,N_8273,N_8212);
or U11569 (N_11569,N_6972,N_7694);
nor U11570 (N_11570,N_6281,N_7539);
or U11571 (N_11571,N_8249,N_7370);
nor U11572 (N_11572,N_6219,N_7428);
or U11573 (N_11573,N_7869,N_7242);
or U11574 (N_11574,N_6330,N_8629);
or U11575 (N_11575,N_6761,N_6832);
or U11576 (N_11576,N_6117,N_6035);
and U11577 (N_11577,N_6980,N_8761);
nand U11578 (N_11578,N_7618,N_6112);
xnor U11579 (N_11579,N_6521,N_7701);
and U11580 (N_11580,N_6246,N_6169);
nand U11581 (N_11581,N_7544,N_6004);
nor U11582 (N_11582,N_8908,N_6133);
xor U11583 (N_11583,N_6798,N_6203);
or U11584 (N_11584,N_7096,N_6030);
xor U11585 (N_11585,N_6829,N_8724);
or U11586 (N_11586,N_6328,N_7093);
nand U11587 (N_11587,N_8077,N_7639);
or U11588 (N_11588,N_8160,N_6553);
nand U11589 (N_11589,N_6726,N_7289);
nand U11590 (N_11590,N_7762,N_6125);
or U11591 (N_11591,N_8627,N_7380);
or U11592 (N_11592,N_6790,N_8428);
nor U11593 (N_11593,N_6504,N_7677);
and U11594 (N_11594,N_6397,N_7579);
or U11595 (N_11595,N_6722,N_8073);
or U11596 (N_11596,N_8170,N_8916);
xnor U11597 (N_11597,N_7597,N_8511);
xor U11598 (N_11598,N_8226,N_7723);
xor U11599 (N_11599,N_6382,N_8593);
xnor U11600 (N_11600,N_8064,N_6563);
nor U11601 (N_11601,N_8511,N_7862);
or U11602 (N_11602,N_7880,N_7501);
xor U11603 (N_11603,N_6691,N_6476);
and U11604 (N_11604,N_7334,N_7011);
xor U11605 (N_11605,N_6565,N_6313);
nor U11606 (N_11606,N_8308,N_7292);
xnor U11607 (N_11607,N_7964,N_8029);
or U11608 (N_11608,N_6933,N_8616);
xnor U11609 (N_11609,N_8500,N_7594);
xnor U11610 (N_11610,N_7059,N_8869);
nand U11611 (N_11611,N_8002,N_6668);
or U11612 (N_11612,N_8339,N_8455);
or U11613 (N_11613,N_6672,N_6264);
nor U11614 (N_11614,N_6640,N_8742);
and U11615 (N_11615,N_6637,N_6326);
or U11616 (N_11616,N_7199,N_6608);
or U11617 (N_11617,N_8280,N_8051);
nand U11618 (N_11618,N_7143,N_7255);
and U11619 (N_11619,N_7023,N_8946);
nand U11620 (N_11620,N_6733,N_6253);
or U11621 (N_11621,N_8546,N_8432);
and U11622 (N_11622,N_6270,N_6398);
nor U11623 (N_11623,N_6786,N_7196);
and U11624 (N_11624,N_7403,N_6155);
nand U11625 (N_11625,N_6276,N_8441);
xor U11626 (N_11626,N_6018,N_6459);
nor U11627 (N_11627,N_6582,N_8714);
and U11628 (N_11628,N_8754,N_8013);
nor U11629 (N_11629,N_8980,N_7262);
and U11630 (N_11630,N_7854,N_6382);
nand U11631 (N_11631,N_6205,N_6575);
or U11632 (N_11632,N_6209,N_7804);
xor U11633 (N_11633,N_6870,N_8636);
xor U11634 (N_11634,N_8608,N_6416);
or U11635 (N_11635,N_6691,N_7967);
nor U11636 (N_11636,N_8803,N_7729);
nand U11637 (N_11637,N_6066,N_7514);
xor U11638 (N_11638,N_7566,N_8813);
xor U11639 (N_11639,N_6512,N_7047);
or U11640 (N_11640,N_8093,N_6073);
or U11641 (N_11641,N_8805,N_8560);
nand U11642 (N_11642,N_8359,N_8805);
xnor U11643 (N_11643,N_7364,N_8235);
nor U11644 (N_11644,N_6159,N_7070);
or U11645 (N_11645,N_6425,N_7263);
nor U11646 (N_11646,N_8636,N_7906);
xor U11647 (N_11647,N_7407,N_8855);
nor U11648 (N_11648,N_6708,N_7849);
nand U11649 (N_11649,N_7622,N_8900);
nand U11650 (N_11650,N_7378,N_7794);
nand U11651 (N_11651,N_7286,N_7974);
and U11652 (N_11652,N_6890,N_7666);
xnor U11653 (N_11653,N_8068,N_7449);
xor U11654 (N_11654,N_6839,N_6188);
or U11655 (N_11655,N_8035,N_7990);
and U11656 (N_11656,N_6349,N_8858);
and U11657 (N_11657,N_6386,N_8132);
nor U11658 (N_11658,N_8157,N_7385);
or U11659 (N_11659,N_6852,N_7573);
nor U11660 (N_11660,N_7412,N_8726);
and U11661 (N_11661,N_6885,N_6336);
nand U11662 (N_11662,N_6105,N_6712);
nand U11663 (N_11663,N_8578,N_8777);
xnor U11664 (N_11664,N_7138,N_7530);
nor U11665 (N_11665,N_8019,N_7665);
or U11666 (N_11666,N_7058,N_6112);
xor U11667 (N_11667,N_8213,N_6938);
xnor U11668 (N_11668,N_6034,N_7104);
and U11669 (N_11669,N_6648,N_8765);
nor U11670 (N_11670,N_7803,N_7397);
and U11671 (N_11671,N_8075,N_6410);
nand U11672 (N_11672,N_6670,N_7854);
nor U11673 (N_11673,N_6796,N_8808);
or U11674 (N_11674,N_7413,N_7769);
or U11675 (N_11675,N_8809,N_6340);
or U11676 (N_11676,N_7717,N_7223);
nor U11677 (N_11677,N_7865,N_6096);
nor U11678 (N_11678,N_8689,N_8934);
and U11679 (N_11679,N_6676,N_6126);
or U11680 (N_11680,N_7462,N_6719);
xor U11681 (N_11681,N_7865,N_7753);
xor U11682 (N_11682,N_6145,N_7048);
nor U11683 (N_11683,N_8730,N_8647);
or U11684 (N_11684,N_7138,N_7158);
nand U11685 (N_11685,N_8183,N_8547);
or U11686 (N_11686,N_6228,N_8154);
nand U11687 (N_11687,N_7086,N_6347);
nand U11688 (N_11688,N_7720,N_8762);
xor U11689 (N_11689,N_6373,N_7008);
nor U11690 (N_11690,N_6769,N_8832);
or U11691 (N_11691,N_8278,N_7163);
and U11692 (N_11692,N_8030,N_7768);
nand U11693 (N_11693,N_7708,N_6112);
or U11694 (N_11694,N_6822,N_7562);
nand U11695 (N_11695,N_8641,N_6869);
nand U11696 (N_11696,N_8943,N_6775);
xor U11697 (N_11697,N_8555,N_6101);
or U11698 (N_11698,N_8590,N_7176);
nor U11699 (N_11699,N_8597,N_7085);
xor U11700 (N_11700,N_6086,N_6306);
xnor U11701 (N_11701,N_8316,N_7379);
nand U11702 (N_11702,N_8984,N_8315);
or U11703 (N_11703,N_8527,N_8918);
or U11704 (N_11704,N_8759,N_8995);
nor U11705 (N_11705,N_6668,N_8861);
or U11706 (N_11706,N_6250,N_7885);
nor U11707 (N_11707,N_7243,N_7545);
nand U11708 (N_11708,N_6838,N_7985);
or U11709 (N_11709,N_7105,N_7912);
nor U11710 (N_11710,N_6909,N_6428);
nor U11711 (N_11711,N_7719,N_6817);
nor U11712 (N_11712,N_6691,N_8030);
nand U11713 (N_11713,N_6169,N_6154);
or U11714 (N_11714,N_6968,N_7705);
nand U11715 (N_11715,N_8431,N_8049);
or U11716 (N_11716,N_7021,N_7394);
nand U11717 (N_11717,N_7828,N_7695);
and U11718 (N_11718,N_8533,N_8271);
and U11719 (N_11719,N_6421,N_7590);
or U11720 (N_11720,N_8693,N_8122);
and U11721 (N_11721,N_8276,N_8431);
nand U11722 (N_11722,N_6555,N_6974);
nand U11723 (N_11723,N_8741,N_8657);
and U11724 (N_11724,N_8621,N_8370);
nor U11725 (N_11725,N_6877,N_6190);
xor U11726 (N_11726,N_7627,N_6068);
xor U11727 (N_11727,N_8281,N_8869);
nand U11728 (N_11728,N_8394,N_8527);
xor U11729 (N_11729,N_8766,N_8293);
nor U11730 (N_11730,N_8858,N_7597);
nand U11731 (N_11731,N_7147,N_7471);
nor U11732 (N_11732,N_8417,N_6564);
or U11733 (N_11733,N_7487,N_6277);
or U11734 (N_11734,N_6344,N_7852);
nand U11735 (N_11735,N_7901,N_7177);
and U11736 (N_11736,N_8088,N_7182);
nand U11737 (N_11737,N_7871,N_7666);
xor U11738 (N_11738,N_6682,N_6072);
and U11739 (N_11739,N_8530,N_7071);
or U11740 (N_11740,N_6517,N_6145);
and U11741 (N_11741,N_6107,N_8686);
or U11742 (N_11742,N_7373,N_6340);
and U11743 (N_11743,N_7509,N_7548);
nor U11744 (N_11744,N_7401,N_6040);
and U11745 (N_11745,N_7270,N_6224);
and U11746 (N_11746,N_8446,N_7216);
xnor U11747 (N_11747,N_6532,N_6983);
nor U11748 (N_11748,N_8055,N_7270);
nor U11749 (N_11749,N_7208,N_7261);
xor U11750 (N_11750,N_8939,N_6252);
nor U11751 (N_11751,N_7109,N_6009);
xnor U11752 (N_11752,N_7991,N_6331);
or U11753 (N_11753,N_8028,N_7385);
nand U11754 (N_11754,N_7051,N_8372);
or U11755 (N_11755,N_7033,N_6862);
or U11756 (N_11756,N_6373,N_7733);
nand U11757 (N_11757,N_7459,N_7001);
or U11758 (N_11758,N_6485,N_6254);
or U11759 (N_11759,N_7892,N_7364);
nand U11760 (N_11760,N_6353,N_7109);
nor U11761 (N_11761,N_8995,N_7225);
nand U11762 (N_11762,N_7474,N_7603);
or U11763 (N_11763,N_8192,N_8201);
nor U11764 (N_11764,N_7667,N_7552);
nor U11765 (N_11765,N_6531,N_7555);
and U11766 (N_11766,N_8350,N_6632);
nand U11767 (N_11767,N_8777,N_7492);
or U11768 (N_11768,N_7994,N_7897);
xor U11769 (N_11769,N_6427,N_8834);
xnor U11770 (N_11770,N_7776,N_6945);
and U11771 (N_11771,N_8912,N_7236);
or U11772 (N_11772,N_7448,N_6050);
or U11773 (N_11773,N_7681,N_7318);
and U11774 (N_11774,N_8252,N_8151);
nor U11775 (N_11775,N_6698,N_8154);
xnor U11776 (N_11776,N_6129,N_6452);
nand U11777 (N_11777,N_8729,N_7736);
xor U11778 (N_11778,N_7674,N_6997);
or U11779 (N_11779,N_8525,N_8967);
nor U11780 (N_11780,N_7471,N_7086);
xnor U11781 (N_11781,N_7261,N_7907);
nand U11782 (N_11782,N_6589,N_6903);
or U11783 (N_11783,N_8329,N_6906);
and U11784 (N_11784,N_8386,N_8958);
nor U11785 (N_11785,N_6190,N_7175);
nand U11786 (N_11786,N_7142,N_6277);
and U11787 (N_11787,N_8148,N_7354);
and U11788 (N_11788,N_7268,N_7831);
xnor U11789 (N_11789,N_8756,N_6716);
xnor U11790 (N_11790,N_7695,N_7760);
xnor U11791 (N_11791,N_8470,N_7013);
and U11792 (N_11792,N_6108,N_8213);
xor U11793 (N_11793,N_7614,N_6260);
xnor U11794 (N_11794,N_8582,N_6298);
and U11795 (N_11795,N_6639,N_6955);
nand U11796 (N_11796,N_6567,N_6106);
and U11797 (N_11797,N_6181,N_7394);
or U11798 (N_11798,N_7936,N_7601);
or U11799 (N_11799,N_6195,N_6208);
nand U11800 (N_11800,N_6051,N_7900);
or U11801 (N_11801,N_6712,N_7405);
and U11802 (N_11802,N_6289,N_8214);
xnor U11803 (N_11803,N_7280,N_6912);
or U11804 (N_11804,N_7477,N_8759);
and U11805 (N_11805,N_6573,N_8683);
and U11806 (N_11806,N_8754,N_6701);
nand U11807 (N_11807,N_6961,N_8811);
nor U11808 (N_11808,N_6340,N_6156);
nor U11809 (N_11809,N_8025,N_7865);
nand U11810 (N_11810,N_6475,N_7294);
nor U11811 (N_11811,N_6379,N_7718);
and U11812 (N_11812,N_6105,N_6154);
xor U11813 (N_11813,N_7679,N_6254);
nor U11814 (N_11814,N_6848,N_7267);
and U11815 (N_11815,N_8802,N_8518);
nand U11816 (N_11816,N_6681,N_6887);
or U11817 (N_11817,N_7471,N_6260);
nor U11818 (N_11818,N_8593,N_6205);
or U11819 (N_11819,N_8858,N_7584);
or U11820 (N_11820,N_8524,N_8799);
or U11821 (N_11821,N_7230,N_7236);
xor U11822 (N_11822,N_6998,N_6414);
xor U11823 (N_11823,N_8511,N_6119);
xnor U11824 (N_11824,N_6830,N_7073);
xnor U11825 (N_11825,N_6390,N_7793);
and U11826 (N_11826,N_8747,N_8704);
nand U11827 (N_11827,N_7053,N_6866);
and U11828 (N_11828,N_8283,N_7524);
or U11829 (N_11829,N_7970,N_7728);
xnor U11830 (N_11830,N_8184,N_7761);
and U11831 (N_11831,N_6829,N_6131);
nor U11832 (N_11832,N_7815,N_7866);
xor U11833 (N_11833,N_7557,N_8152);
and U11834 (N_11834,N_6568,N_7086);
nand U11835 (N_11835,N_7688,N_7584);
nor U11836 (N_11836,N_8185,N_6734);
nor U11837 (N_11837,N_7917,N_8631);
or U11838 (N_11838,N_8984,N_6830);
nor U11839 (N_11839,N_7402,N_6387);
or U11840 (N_11840,N_7534,N_7712);
xor U11841 (N_11841,N_7721,N_6225);
xor U11842 (N_11842,N_7526,N_7829);
xnor U11843 (N_11843,N_8302,N_7220);
nand U11844 (N_11844,N_7680,N_7913);
or U11845 (N_11845,N_6799,N_8919);
nor U11846 (N_11846,N_6106,N_6673);
xor U11847 (N_11847,N_8108,N_7293);
nor U11848 (N_11848,N_6637,N_7182);
or U11849 (N_11849,N_7183,N_8496);
nand U11850 (N_11850,N_7795,N_6384);
xor U11851 (N_11851,N_6488,N_8736);
or U11852 (N_11852,N_8529,N_6453);
xnor U11853 (N_11853,N_6917,N_8110);
nand U11854 (N_11854,N_7849,N_7916);
xnor U11855 (N_11855,N_8759,N_8682);
xor U11856 (N_11856,N_8985,N_6269);
and U11857 (N_11857,N_6486,N_7295);
nor U11858 (N_11858,N_8351,N_6282);
and U11859 (N_11859,N_7731,N_7992);
or U11860 (N_11860,N_7631,N_7454);
and U11861 (N_11861,N_6975,N_8862);
nor U11862 (N_11862,N_8576,N_6262);
nor U11863 (N_11863,N_7284,N_7615);
or U11864 (N_11864,N_6514,N_6584);
nand U11865 (N_11865,N_6134,N_6752);
or U11866 (N_11866,N_8265,N_7763);
and U11867 (N_11867,N_8480,N_6883);
or U11868 (N_11868,N_6540,N_6773);
nor U11869 (N_11869,N_7039,N_8557);
nand U11870 (N_11870,N_7083,N_6600);
and U11871 (N_11871,N_6258,N_8638);
nand U11872 (N_11872,N_6505,N_8239);
and U11873 (N_11873,N_8846,N_8331);
or U11874 (N_11874,N_6291,N_7663);
xor U11875 (N_11875,N_7199,N_6523);
and U11876 (N_11876,N_7119,N_6957);
and U11877 (N_11877,N_6394,N_7142);
xnor U11878 (N_11878,N_6810,N_8402);
nor U11879 (N_11879,N_7327,N_6137);
nor U11880 (N_11880,N_6226,N_7932);
or U11881 (N_11881,N_8596,N_8677);
nor U11882 (N_11882,N_8384,N_8910);
nand U11883 (N_11883,N_6976,N_7244);
and U11884 (N_11884,N_6962,N_6755);
and U11885 (N_11885,N_8682,N_8860);
nand U11886 (N_11886,N_7091,N_6711);
or U11887 (N_11887,N_8069,N_7105);
nor U11888 (N_11888,N_7677,N_6577);
or U11889 (N_11889,N_8383,N_7480);
or U11890 (N_11890,N_6241,N_8872);
nor U11891 (N_11891,N_8678,N_6191);
xor U11892 (N_11892,N_7787,N_7417);
nor U11893 (N_11893,N_8072,N_6525);
and U11894 (N_11894,N_6792,N_7060);
nand U11895 (N_11895,N_8253,N_7396);
nor U11896 (N_11896,N_8817,N_7551);
or U11897 (N_11897,N_8096,N_7946);
and U11898 (N_11898,N_7272,N_6482);
nor U11899 (N_11899,N_6010,N_6073);
and U11900 (N_11900,N_6276,N_6432);
xor U11901 (N_11901,N_6619,N_8089);
xnor U11902 (N_11902,N_8363,N_8491);
nor U11903 (N_11903,N_6695,N_7675);
and U11904 (N_11904,N_8407,N_7041);
xnor U11905 (N_11905,N_8429,N_6636);
nand U11906 (N_11906,N_6483,N_8232);
or U11907 (N_11907,N_7559,N_8204);
xnor U11908 (N_11908,N_6388,N_6247);
xor U11909 (N_11909,N_8017,N_7331);
nand U11910 (N_11910,N_8855,N_6796);
or U11911 (N_11911,N_7965,N_8574);
or U11912 (N_11912,N_6902,N_7585);
xnor U11913 (N_11913,N_6280,N_6268);
nand U11914 (N_11914,N_8535,N_7955);
and U11915 (N_11915,N_7414,N_6950);
or U11916 (N_11916,N_7411,N_8558);
nand U11917 (N_11917,N_7840,N_7411);
nand U11918 (N_11918,N_8716,N_8217);
or U11919 (N_11919,N_8038,N_7612);
xnor U11920 (N_11920,N_8349,N_7885);
nand U11921 (N_11921,N_6517,N_8244);
xor U11922 (N_11922,N_6552,N_6325);
nor U11923 (N_11923,N_8051,N_6733);
nor U11924 (N_11924,N_7451,N_8797);
xnor U11925 (N_11925,N_6482,N_7415);
xor U11926 (N_11926,N_8248,N_6310);
nor U11927 (N_11927,N_8479,N_7303);
nand U11928 (N_11928,N_6767,N_7118);
xnor U11929 (N_11929,N_8382,N_7297);
xnor U11930 (N_11930,N_7495,N_6620);
or U11931 (N_11931,N_7330,N_8626);
nand U11932 (N_11932,N_7113,N_6534);
nand U11933 (N_11933,N_8658,N_8617);
xor U11934 (N_11934,N_6739,N_7189);
nor U11935 (N_11935,N_7187,N_8201);
xnor U11936 (N_11936,N_6617,N_6682);
or U11937 (N_11937,N_6897,N_6314);
or U11938 (N_11938,N_8559,N_6197);
nor U11939 (N_11939,N_7711,N_8669);
and U11940 (N_11940,N_7621,N_6906);
or U11941 (N_11941,N_8679,N_6877);
xnor U11942 (N_11942,N_8830,N_8274);
and U11943 (N_11943,N_6804,N_8596);
nand U11944 (N_11944,N_8609,N_7046);
nand U11945 (N_11945,N_7684,N_8193);
nor U11946 (N_11946,N_8787,N_7324);
xnor U11947 (N_11947,N_7410,N_8002);
nand U11948 (N_11948,N_8878,N_7804);
nor U11949 (N_11949,N_7984,N_7762);
nand U11950 (N_11950,N_8172,N_8713);
and U11951 (N_11951,N_6744,N_6664);
and U11952 (N_11952,N_7699,N_7007);
nor U11953 (N_11953,N_8379,N_7898);
xor U11954 (N_11954,N_6542,N_6281);
xnor U11955 (N_11955,N_8461,N_8192);
xor U11956 (N_11956,N_7096,N_7780);
nor U11957 (N_11957,N_7402,N_7576);
nor U11958 (N_11958,N_6592,N_6915);
nor U11959 (N_11959,N_6023,N_8595);
or U11960 (N_11960,N_6330,N_7705);
nand U11961 (N_11961,N_6198,N_8780);
and U11962 (N_11962,N_8910,N_6227);
xnor U11963 (N_11963,N_7694,N_6796);
xor U11964 (N_11964,N_8984,N_6896);
and U11965 (N_11965,N_6716,N_6155);
or U11966 (N_11966,N_6179,N_8605);
nand U11967 (N_11967,N_8879,N_7344);
nor U11968 (N_11968,N_6673,N_6360);
xor U11969 (N_11969,N_6057,N_8214);
and U11970 (N_11970,N_6201,N_6242);
nor U11971 (N_11971,N_8261,N_6777);
and U11972 (N_11972,N_8694,N_8845);
nand U11973 (N_11973,N_8850,N_7937);
and U11974 (N_11974,N_6068,N_8185);
xor U11975 (N_11975,N_7594,N_7518);
and U11976 (N_11976,N_7390,N_8982);
or U11977 (N_11977,N_7190,N_6703);
or U11978 (N_11978,N_7604,N_8718);
nand U11979 (N_11979,N_7983,N_8188);
nand U11980 (N_11980,N_6355,N_8127);
nor U11981 (N_11981,N_6150,N_7616);
nand U11982 (N_11982,N_7645,N_8010);
nor U11983 (N_11983,N_7565,N_6601);
or U11984 (N_11984,N_6090,N_8321);
or U11985 (N_11985,N_6181,N_7545);
xor U11986 (N_11986,N_7261,N_7536);
xnor U11987 (N_11987,N_7686,N_7654);
or U11988 (N_11988,N_8297,N_7459);
xor U11989 (N_11989,N_7050,N_8552);
nand U11990 (N_11990,N_7919,N_7219);
xnor U11991 (N_11991,N_6705,N_7836);
nand U11992 (N_11992,N_7809,N_7307);
or U11993 (N_11993,N_7967,N_7247);
nand U11994 (N_11994,N_8273,N_6823);
nand U11995 (N_11995,N_6745,N_7355);
nand U11996 (N_11996,N_6972,N_8028);
nor U11997 (N_11997,N_6032,N_7863);
nor U11998 (N_11998,N_6543,N_7044);
nor U11999 (N_11999,N_8818,N_7706);
and U12000 (N_12000,N_9539,N_9924);
nor U12001 (N_12001,N_9068,N_11663);
or U12002 (N_12002,N_9935,N_11604);
or U12003 (N_12003,N_9323,N_11708);
xor U12004 (N_12004,N_9882,N_9511);
and U12005 (N_12005,N_10002,N_11119);
or U12006 (N_12006,N_10332,N_9582);
xnor U12007 (N_12007,N_9691,N_11463);
or U12008 (N_12008,N_9457,N_10765);
nand U12009 (N_12009,N_11169,N_11652);
or U12010 (N_12010,N_10891,N_9571);
nor U12011 (N_12011,N_11156,N_10851);
and U12012 (N_12012,N_11061,N_9167);
xnor U12013 (N_12013,N_10262,N_11151);
nand U12014 (N_12014,N_9586,N_10515);
nand U12015 (N_12015,N_10907,N_11741);
or U12016 (N_12016,N_11395,N_9273);
xnor U12017 (N_12017,N_10822,N_11396);
nand U12018 (N_12018,N_11357,N_11097);
xor U12019 (N_12019,N_9812,N_9821);
or U12020 (N_12020,N_11812,N_10229);
nor U12021 (N_12021,N_11908,N_9763);
or U12022 (N_12022,N_10609,N_9578);
xor U12023 (N_12023,N_10673,N_10812);
and U12024 (N_12024,N_11497,N_9561);
or U12025 (N_12025,N_9491,N_9253);
nand U12026 (N_12026,N_11719,N_9341);
or U12027 (N_12027,N_11041,N_10846);
nand U12028 (N_12028,N_10892,N_9408);
nor U12029 (N_12029,N_10434,N_11465);
nor U12030 (N_12030,N_11054,N_9676);
nor U12031 (N_12031,N_9029,N_9121);
and U12032 (N_12032,N_11832,N_10992);
or U12033 (N_12033,N_10204,N_11434);
or U12034 (N_12034,N_11849,N_9061);
or U12035 (N_12035,N_10773,N_11569);
nor U12036 (N_12036,N_9100,N_11455);
or U12037 (N_12037,N_11593,N_10076);
nand U12038 (N_12038,N_9410,N_9805);
nand U12039 (N_12039,N_9002,N_9831);
nand U12040 (N_12040,N_9069,N_11913);
nand U12041 (N_12041,N_9976,N_9795);
nand U12042 (N_12042,N_9439,N_9466);
or U12043 (N_12043,N_10792,N_10875);
and U12044 (N_12044,N_11304,N_10728);
xnor U12045 (N_12045,N_10420,N_9462);
nor U12046 (N_12046,N_11992,N_11748);
nor U12047 (N_12047,N_9200,N_9858);
and U12048 (N_12048,N_9208,N_11608);
or U12049 (N_12049,N_9105,N_10122);
xor U12050 (N_12050,N_11583,N_9572);
and U12051 (N_12051,N_11784,N_10209);
or U12052 (N_12052,N_9475,N_9468);
nor U12053 (N_12053,N_11934,N_11603);
and U12054 (N_12054,N_9728,N_11090);
and U12055 (N_12055,N_9168,N_10772);
nor U12056 (N_12056,N_10705,N_11763);
and U12057 (N_12057,N_9897,N_9957);
and U12058 (N_12058,N_9127,N_10624);
or U12059 (N_12059,N_11888,N_10326);
nor U12060 (N_12060,N_11870,N_10422);
xor U12061 (N_12061,N_11247,N_10459);
and U12062 (N_12062,N_10201,N_10651);
or U12063 (N_12063,N_10713,N_9126);
nor U12064 (N_12064,N_10330,N_9404);
xor U12065 (N_12065,N_11843,N_10981);
and U12066 (N_12066,N_9875,N_11922);
and U12067 (N_12067,N_11354,N_11044);
or U12068 (N_12068,N_10180,N_9204);
nor U12069 (N_12069,N_10775,N_10176);
nor U12070 (N_12070,N_11880,N_11523);
xnor U12071 (N_12071,N_9237,N_9946);
nor U12072 (N_12072,N_9284,N_9715);
xor U12073 (N_12073,N_10887,N_9723);
nand U12074 (N_12074,N_11493,N_11915);
nand U12075 (N_12075,N_11785,N_9714);
and U12076 (N_12076,N_11985,N_11745);
nand U12077 (N_12077,N_9624,N_9879);
or U12078 (N_12078,N_9137,N_10516);
and U12079 (N_12079,N_11052,N_9358);
nand U12080 (N_12080,N_10505,N_9318);
nand U12081 (N_12081,N_11294,N_11494);
xor U12082 (N_12082,N_9067,N_9617);
xnor U12083 (N_12083,N_9667,N_9832);
nand U12084 (N_12084,N_9095,N_10782);
xor U12085 (N_12085,N_11997,N_9652);
nor U12086 (N_12086,N_11162,N_10649);
xor U12087 (N_12087,N_10636,N_9816);
nor U12088 (N_12088,N_11794,N_11651);
and U12089 (N_12089,N_9635,N_11215);
and U12090 (N_12090,N_11557,N_10831);
and U12091 (N_12091,N_9809,N_9163);
nor U12092 (N_12092,N_11083,N_10294);
and U12093 (N_12093,N_11877,N_10921);
nand U12094 (N_12094,N_11799,N_9209);
and U12095 (N_12095,N_11034,N_10223);
xor U12096 (N_12096,N_10743,N_11895);
nor U12097 (N_12097,N_10170,N_10716);
nand U12098 (N_12098,N_9923,N_9140);
or U12099 (N_12099,N_9604,N_11264);
or U12100 (N_12100,N_9931,N_9449);
or U12101 (N_12101,N_9428,N_9490);
nor U12102 (N_12102,N_10724,N_9071);
and U12103 (N_12103,N_9009,N_11805);
nand U12104 (N_12104,N_11925,N_9302);
or U12105 (N_12105,N_11277,N_9735);
and U12106 (N_12106,N_11687,N_11062);
xor U12107 (N_12107,N_9709,N_10087);
nand U12108 (N_12108,N_9696,N_10449);
nand U12109 (N_12109,N_9919,N_9264);
nand U12110 (N_12110,N_9603,N_11136);
nor U12111 (N_12111,N_11372,N_10579);
nand U12112 (N_12112,N_11195,N_10581);
nand U12113 (N_12113,N_9899,N_10856);
and U12114 (N_12114,N_9514,N_10497);
and U12115 (N_12115,N_9164,N_11007);
or U12116 (N_12116,N_10469,N_10686);
xor U12117 (N_12117,N_11017,N_11636);
nor U12118 (N_12118,N_9834,N_10642);
nor U12119 (N_12119,N_9672,N_9568);
nand U12120 (N_12120,N_10273,N_11358);
nor U12121 (N_12121,N_11756,N_11871);
xor U12122 (N_12122,N_9848,N_9089);
and U12123 (N_12123,N_9355,N_9653);
and U12124 (N_12124,N_10553,N_11689);
nor U12125 (N_12125,N_10460,N_11365);
and U12126 (N_12126,N_10308,N_9978);
xor U12127 (N_12127,N_9927,N_11001);
and U12128 (N_12128,N_9049,N_11541);
and U12129 (N_12129,N_11677,N_10654);
xnor U12130 (N_12130,N_9835,N_9540);
nor U12131 (N_12131,N_10928,N_10898);
or U12132 (N_12132,N_10361,N_9786);
and U12133 (N_12133,N_10166,N_9869);
and U12134 (N_12134,N_11182,N_9116);
nand U12135 (N_12135,N_9373,N_10997);
and U12136 (N_12136,N_10770,N_9296);
nand U12137 (N_12137,N_10450,N_11456);
and U12138 (N_12138,N_10755,N_11158);
or U12139 (N_12139,N_10196,N_10036);
or U12140 (N_12140,N_11907,N_10511);
nand U12141 (N_12141,N_11701,N_9390);
or U12142 (N_12142,N_11927,N_10025);
nor U12143 (N_12143,N_10000,N_10185);
and U12144 (N_12144,N_10888,N_9352);
nor U12145 (N_12145,N_9308,N_10070);
nand U12146 (N_12146,N_9291,N_9001);
or U12147 (N_12147,N_10710,N_9228);
and U12148 (N_12148,N_11046,N_9732);
or U12149 (N_12149,N_9937,N_9782);
nand U12150 (N_12150,N_11959,N_11290);
and U12151 (N_12151,N_11937,N_11644);
xor U12152 (N_12152,N_10969,N_11574);
and U12153 (N_12153,N_11248,N_10530);
xnor U12154 (N_12154,N_11953,N_9815);
or U12155 (N_12155,N_10671,N_10726);
xor U12156 (N_12156,N_9194,N_10408);
nand U12157 (N_12157,N_9954,N_10576);
nor U12158 (N_12158,N_10554,N_10913);
nor U12159 (N_12159,N_9960,N_10005);
nor U12160 (N_12160,N_9144,N_11690);
and U12161 (N_12161,N_10104,N_10022);
nand U12162 (N_12162,N_9893,N_10599);
or U12163 (N_12163,N_10869,N_11814);
nor U12164 (N_12164,N_11637,N_11060);
nand U12165 (N_12165,N_10144,N_9533);
nor U12166 (N_12166,N_9781,N_10098);
nor U12167 (N_12167,N_11536,N_9399);
or U12168 (N_12168,N_9365,N_10396);
and U12169 (N_12169,N_10964,N_11906);
and U12170 (N_12170,N_10682,N_10717);
or U12171 (N_12171,N_9531,N_11274);
xor U12172 (N_12172,N_9925,N_10764);
xor U12173 (N_12173,N_10946,N_10054);
or U12174 (N_12174,N_11964,N_10954);
nor U12175 (N_12175,N_9701,N_11946);
xnor U12176 (N_12176,N_11955,N_10539);
xor U12177 (N_12177,N_9799,N_11995);
nor U12178 (N_12178,N_9698,N_9006);
xnor U12179 (N_12179,N_10238,N_10043);
or U12180 (N_12180,N_11691,N_10967);
xor U12181 (N_12181,N_11682,N_10035);
and U12182 (N_12182,N_10307,N_10081);
nor U12183 (N_12183,N_9827,N_9917);
and U12184 (N_12184,N_9138,N_11932);
or U12185 (N_12185,N_10323,N_11257);
nand U12186 (N_12186,N_9377,N_11234);
nand U12187 (N_12187,N_9972,N_9523);
and U12188 (N_12188,N_11478,N_11028);
and U12189 (N_12189,N_9471,N_11129);
xor U12190 (N_12190,N_11101,N_10565);
or U12191 (N_12191,N_10694,N_10252);
or U12192 (N_12192,N_11170,N_11683);
or U12193 (N_12193,N_11951,N_11591);
and U12194 (N_12194,N_11567,N_11408);
or U12195 (N_12195,N_9883,N_9712);
or U12196 (N_12196,N_9780,N_11853);
nor U12197 (N_12197,N_11271,N_10142);
and U12198 (N_12198,N_9150,N_9565);
nor U12199 (N_12199,N_11822,N_9814);
nor U12200 (N_12200,N_10476,N_11808);
and U12201 (N_12201,N_11551,N_10503);
or U12202 (N_12202,N_11440,N_11505);
or U12203 (N_12203,N_9015,N_10113);
and U12204 (N_12204,N_11080,N_9430);
nor U12205 (N_12205,N_11473,N_9460);
nor U12206 (N_12206,N_10135,N_11602);
nor U12207 (N_12207,N_9785,N_11232);
and U12208 (N_12208,N_9620,N_9804);
nand U12209 (N_12209,N_10795,N_10498);
and U12210 (N_12210,N_11199,N_10653);
or U12211 (N_12211,N_10894,N_10067);
xnor U12212 (N_12212,N_10443,N_10518);
nor U12213 (N_12213,N_9711,N_11680);
xnor U12214 (N_12214,N_10612,N_11426);
nand U12215 (N_12215,N_10998,N_9246);
nor U12216 (N_12216,N_11219,N_10883);
or U12217 (N_12217,N_11511,N_9211);
and U12218 (N_12218,N_11786,N_10814);
and U12219 (N_12219,N_11163,N_9479);
xor U12220 (N_12220,N_10030,N_10573);
nor U12221 (N_12221,N_10102,N_10933);
and U12222 (N_12222,N_9555,N_10520);
or U12223 (N_12223,N_9614,N_10232);
or U12224 (N_12224,N_10521,N_11464);
xnor U12225 (N_12225,N_9195,N_10438);
xnor U12226 (N_12226,N_10622,N_9829);
nor U12227 (N_12227,N_11367,N_9192);
nand U12228 (N_12228,N_9287,N_11297);
and U12229 (N_12229,N_11949,N_9379);
or U12230 (N_12230,N_10629,N_9091);
nand U12231 (N_12231,N_9496,N_10645);
nor U12232 (N_12232,N_9492,N_11578);
and U12233 (N_12233,N_11999,N_9156);
xnor U12234 (N_12234,N_10344,N_9594);
or U12235 (N_12235,N_11622,N_10314);
xor U12236 (N_12236,N_11935,N_11560);
nor U12237 (N_12237,N_9376,N_11758);
nor U12238 (N_12238,N_11890,N_9864);
xnor U12239 (N_12239,N_10300,N_9359);
nand U12240 (N_12240,N_10251,N_10152);
and U12241 (N_12241,N_11150,N_9332);
xnor U12242 (N_12242,N_9054,N_10631);
nor U12243 (N_12243,N_9940,N_9744);
and U12244 (N_12244,N_9996,N_9463);
nand U12245 (N_12245,N_9928,N_11834);
xnor U12246 (N_12246,N_11283,N_9650);
xor U12247 (N_12247,N_11082,N_9991);
and U12248 (N_12248,N_9967,N_10820);
nand U12249 (N_12249,N_10555,N_9538);
or U12250 (N_12250,N_9175,N_11127);
nor U12251 (N_12251,N_9421,N_9870);
xnor U12252 (N_12252,N_11811,N_9980);
or U12253 (N_12253,N_10362,N_10392);
xnor U12254 (N_12254,N_10889,N_11522);
or U12255 (N_12255,N_10721,N_9682);
or U12256 (N_12256,N_9304,N_11516);
or U12257 (N_12257,N_11809,N_10077);
nand U12258 (N_12258,N_11334,N_10661);
nor U12259 (N_12259,N_10341,N_11423);
xnor U12260 (N_12260,N_10777,N_10970);
xor U12261 (N_12261,N_9292,N_10588);
nor U12262 (N_12262,N_11614,N_10130);
or U12263 (N_12263,N_11787,N_11045);
xnor U12264 (N_12264,N_11032,N_11432);
xor U12265 (N_12265,N_10213,N_11980);
or U12266 (N_12266,N_9685,N_10684);
and U12267 (N_12267,N_9939,N_11236);
nor U12268 (N_12268,N_10269,N_11280);
or U12269 (N_12269,N_9139,N_10372);
and U12270 (N_12270,N_11855,N_11111);
xnor U12271 (N_12271,N_11209,N_11078);
xor U12272 (N_12272,N_10802,N_9549);
nor U12273 (N_12273,N_10377,N_11149);
nand U12274 (N_12274,N_9753,N_10864);
nand U12275 (N_12275,N_11308,N_9766);
nand U12276 (N_12276,N_11715,N_9317);
xor U12277 (N_12277,N_10853,N_10837);
nand U12278 (N_12278,N_10725,N_9933);
and U12279 (N_12279,N_10492,N_9674);
or U12280 (N_12280,N_11771,N_11442);
nand U12281 (N_12281,N_10955,N_10348);
nor U12282 (N_12282,N_11030,N_10698);
and U12283 (N_12283,N_11342,N_11769);
and U12284 (N_12284,N_10474,N_10940);
or U12285 (N_12285,N_9312,N_10138);
nor U12286 (N_12286,N_10123,N_9043);
xor U12287 (N_12287,N_9014,N_10762);
nor U12288 (N_12288,N_9385,N_10606);
nor U12289 (N_12289,N_11901,N_11008);
and U12290 (N_12290,N_11712,N_11295);
nor U12291 (N_12291,N_9193,N_9784);
nor U12292 (N_12292,N_9160,N_11393);
and U12293 (N_12293,N_11036,N_11508);
nand U12294 (N_12294,N_11923,N_10711);
xnor U12295 (N_12295,N_11495,N_10256);
xor U12296 (N_12296,N_10932,N_10013);
and U12297 (N_12297,N_9665,N_9575);
or U12298 (N_12298,N_10595,N_11875);
nand U12299 (N_12299,N_9099,N_10215);
nand U12300 (N_12300,N_9597,N_10454);
or U12301 (N_12301,N_11065,N_9666);
or U12302 (N_12302,N_9506,N_11392);
or U12303 (N_12303,N_9039,N_11400);
and U12304 (N_12304,N_9670,N_9495);
xor U12305 (N_12305,N_10212,N_11472);
or U12306 (N_12306,N_11053,N_11340);
nand U12307 (N_12307,N_11592,N_10452);
nand U12308 (N_12308,N_9649,N_10137);
xnor U12309 (N_12309,N_10024,N_10089);
or U12310 (N_12310,N_11343,N_11255);
nand U12311 (N_12311,N_11040,N_11279);
nand U12312 (N_12312,N_11641,N_9181);
nor U12313 (N_12313,N_11931,N_10331);
and U12314 (N_12314,N_10739,N_9431);
or U12315 (N_12315,N_10304,N_10991);
nor U12316 (N_12316,N_9016,N_10284);
nor U12317 (N_12317,N_11211,N_11619);
nor U12318 (N_12318,N_9473,N_11015);
nor U12319 (N_12319,N_11282,N_10867);
nor U12320 (N_12320,N_9148,N_10982);
nand U12321 (N_12321,N_10761,N_9543);
xor U12322 (N_12322,N_10766,N_10780);
nor U12323 (N_12323,N_11327,N_11135);
and U12324 (N_12324,N_10283,N_10403);
nor U12325 (N_12325,N_11941,N_9427);
or U12326 (N_12326,N_10914,N_10345);
xor U12327 (N_12327,N_10097,N_9726);
nor U12328 (N_12328,N_11410,N_10064);
and U12329 (N_12329,N_11540,N_10821);
and U12330 (N_12330,N_10689,N_9664);
nor U12331 (N_12331,N_10281,N_9601);
and U12332 (N_12332,N_9129,N_11231);
or U12333 (N_12333,N_9087,N_11596);
nand U12334 (N_12334,N_10563,N_10436);
nor U12335 (N_12335,N_10297,N_11402);
or U12336 (N_12336,N_10816,N_10712);
nand U12337 (N_12337,N_11218,N_10900);
and U12338 (N_12338,N_10676,N_11315);
or U12339 (N_12339,N_11095,N_11382);
and U12340 (N_12340,N_9310,N_10927);
nor U12341 (N_12341,N_9411,N_9743);
nor U12342 (N_12342,N_11164,N_9529);
or U12343 (N_12343,N_11978,N_10590);
nor U12344 (N_12344,N_11984,N_10321);
xnor U12345 (N_12345,N_11605,N_10745);
and U12346 (N_12346,N_9968,N_9884);
nor U12347 (N_12347,N_10715,N_10029);
and U12348 (N_12348,N_10248,N_10222);
nor U12349 (N_12349,N_11178,N_10159);
or U12350 (N_12350,N_9364,N_10552);
or U12351 (N_12351,N_10390,N_9407);
xnor U12352 (N_12352,N_9372,N_11798);
xor U12353 (N_12353,N_9335,N_10803);
and U12354 (N_12354,N_9557,N_10243);
and U12355 (N_12355,N_10401,N_11138);
nand U12356 (N_12356,N_9438,N_9964);
xor U12357 (N_12357,N_9777,N_10560);
xor U12358 (N_12358,N_10990,N_9521);
nor U12359 (N_12359,N_9545,N_9589);
or U12360 (N_12360,N_11801,N_9461);
and U12361 (N_12361,N_11079,N_11933);
and U12362 (N_12362,N_9904,N_9337);
and U12363 (N_12363,N_9792,N_11161);
nand U12364 (N_12364,N_11502,N_11291);
and U12365 (N_12365,N_11662,N_10410);
xor U12366 (N_12366,N_9227,N_11134);
or U12367 (N_12367,N_9342,N_10621);
and U12368 (N_12368,N_10291,N_9500);
or U12369 (N_12369,N_9678,N_9267);
and U12370 (N_12370,N_9697,N_10187);
or U12371 (N_12371,N_11289,N_11697);
nand U12372 (N_12372,N_10136,N_11005);
nand U12373 (N_12373,N_11731,N_10627);
or U12374 (N_12374,N_10605,N_9590);
or U12375 (N_12375,N_9891,N_11568);
and U12376 (N_12376,N_9269,N_9853);
or U12377 (N_12377,N_10120,N_9081);
and U12378 (N_12378,N_11986,N_10971);
xnor U12379 (N_12379,N_9789,N_9961);
and U12380 (N_12380,N_9737,N_11318);
nand U12381 (N_12381,N_9623,N_9695);
and U12382 (N_12382,N_9602,N_10619);
or U12383 (N_12383,N_9559,N_11020);
xor U12384 (N_12384,N_9052,N_10417);
nor U12385 (N_12385,N_9608,N_10194);
xor U12386 (N_12386,N_10574,N_10440);
or U12387 (N_12387,N_10873,N_11789);
xnor U12388 (N_12388,N_11293,N_11706);
nand U12389 (N_12389,N_9080,N_10161);
and U12390 (N_12390,N_10095,N_11117);
xor U12391 (N_12391,N_9902,N_11887);
xor U12392 (N_12392,N_10100,N_9019);
nor U12393 (N_12393,N_9648,N_11130);
or U12394 (N_12394,N_10117,N_10221);
and U12395 (N_12395,N_9563,N_11673);
and U12396 (N_12396,N_9909,N_9405);
and U12397 (N_12397,N_11921,N_9450);
and U12398 (N_12398,N_11518,N_9658);
nand U12399 (N_12399,N_11886,N_9679);
xnor U12400 (N_12400,N_10744,N_11561);
or U12401 (N_12401,N_11728,N_9881);
nor U12402 (N_12402,N_11369,N_11881);
xor U12403 (N_12403,N_9618,N_10513);
or U12404 (N_12404,N_10550,N_9485);
and U12405 (N_12405,N_10668,N_11326);
or U12406 (N_12406,N_9713,N_10363);
nand U12407 (N_12407,N_11698,N_10220);
nor U12408 (N_12408,N_10360,N_9199);
and U12409 (N_12409,N_10861,N_10068);
nor U12410 (N_12410,N_11833,N_10727);
nand U12411 (N_12411,N_10917,N_10828);
nor U12412 (N_12412,N_11470,N_10429);
and U12413 (N_12413,N_11051,N_10637);
or U12414 (N_12414,N_10165,N_10972);
and U12415 (N_12415,N_11048,N_10655);
nand U12416 (N_12416,N_9392,N_9244);
nand U12417 (N_12417,N_11813,N_11792);
nand U12418 (N_12418,N_9381,N_11404);
xnor U12419 (N_12419,N_9088,N_11196);
or U12420 (N_12420,N_10532,N_9520);
nor U12421 (N_12421,N_11383,N_9519);
nand U12422 (N_12422,N_11348,N_9186);
xor U12423 (N_12423,N_10542,N_11147);
and U12424 (N_12424,N_10254,N_11725);
and U12425 (N_12425,N_11821,N_10486);
nand U12426 (N_12426,N_11067,N_10327);
or U12427 (N_12427,N_10587,N_11524);
nand U12428 (N_12428,N_11742,N_10028);
or U12429 (N_12429,N_9020,N_9914);
nor U12430 (N_12430,N_9515,N_11322);
nand U12431 (N_12431,N_9110,N_10523);
nand U12432 (N_12432,N_11534,N_9971);
xor U12433 (N_12433,N_9348,N_9239);
nor U12434 (N_12434,N_10356,N_9857);
xor U12435 (N_12435,N_10490,N_10038);
or U12436 (N_12436,N_10324,N_9477);
nor U12437 (N_12437,N_10050,N_9028);
nand U12438 (N_12438,N_10027,N_10278);
nor U12439 (N_12439,N_9993,N_10722);
and U12440 (N_12440,N_10545,N_10247);
and U12441 (N_12441,N_10551,N_10033);
nand U12442 (N_12442,N_9012,N_9588);
nand U12443 (N_12443,N_11220,N_9558);
or U12444 (N_12444,N_11462,N_10826);
nor U12445 (N_12445,N_11757,N_9045);
xnor U12446 (N_12446,N_9295,N_11916);
or U12447 (N_12447,N_10522,N_9532);
nand U12448 (N_12448,N_11626,N_11320);
xor U12449 (N_12449,N_10966,N_9083);
nand U12450 (N_12450,N_11613,N_9943);
xor U12451 (N_12451,N_10746,N_10617);
nand U12452 (N_12452,N_9741,N_11056);
or U12453 (N_12453,N_10870,N_10845);
or U12454 (N_12454,N_11982,N_10150);
or U12455 (N_12455,N_9103,N_11852);
and U12456 (N_12456,N_9580,N_9478);
xnor U12457 (N_12457,N_10325,N_9177);
or U12458 (N_12458,N_11033,N_9973);
nand U12459 (N_12459,N_11185,N_10148);
and U12460 (N_12460,N_10956,N_9433);
nand U12461 (N_12461,N_11844,N_10813);
nor U12462 (N_12462,N_9414,N_10594);
and U12463 (N_12463,N_10863,N_10525);
or U12464 (N_12464,N_10384,N_10738);
nor U12465 (N_12465,N_10567,N_9871);
and U12466 (N_12466,N_11276,N_11430);
xnor U12467 (N_12467,N_9950,N_9347);
nor U12468 (N_12468,N_9115,N_9900);
xnor U12469 (N_12469,N_10806,N_10754);
nor U12470 (N_12470,N_9579,N_9426);
nand U12471 (N_12471,N_10596,N_10623);
nand U12472 (N_12472,N_11292,N_10797);
nand U12473 (N_12473,N_10707,N_10255);
and U12474 (N_12474,N_11038,N_11635);
or U12475 (N_12475,N_9331,N_9632);
or U12476 (N_12476,N_11858,N_9742);
or U12477 (N_12477,N_9013,N_9030);
or U12478 (N_12478,N_10391,N_11063);
xor U12479 (N_12479,N_10480,N_11058);
nor U12480 (N_12480,N_11965,N_9704);
nand U12481 (N_12481,N_10389,N_11165);
or U12482 (N_12482,N_10266,N_11137);
or U12483 (N_12483,N_9918,N_11928);
or U12484 (N_12484,N_10174,N_10317);
nor U12485 (N_12485,N_11003,N_9487);
nand U12486 (N_12486,N_10640,N_10471);
or U12487 (N_12487,N_11422,N_10882);
or U12488 (N_12488,N_10834,N_10865);
nor U12489 (N_12489,N_10948,N_9338);
nor U12490 (N_12490,N_9775,N_10646);
and U12491 (N_12491,N_10696,N_11957);
xor U12492 (N_12492,N_11301,N_11443);
or U12493 (N_12493,N_11089,N_10302);
xnor U12494 (N_12494,N_10519,N_10611);
nand U12495 (N_12495,N_10145,N_11990);
or U12496 (N_12496,N_10398,N_9659);
nor U12497 (N_12497,N_11310,N_11123);
nand U12498 (N_12498,N_9154,N_11267);
xor U12499 (N_12499,N_10210,N_10091);
or U12500 (N_12500,N_9486,N_9862);
nand U12501 (N_12501,N_11510,N_9056);
and U12502 (N_12502,N_10757,N_10312);
or U12503 (N_12503,N_10249,N_11107);
nor U12504 (N_12504,N_11363,N_11306);
or U12505 (N_12505,N_11103,N_11245);
or U12506 (N_12506,N_9866,N_11856);
xnor U12507 (N_12507,N_11407,N_11893);
nand U12508 (N_12508,N_9265,N_10078);
nand U12509 (N_12509,N_9339,N_11011);
nand U12510 (N_12510,N_11329,N_11338);
and U12511 (N_12511,N_9576,N_10040);
or U12512 (N_12512,N_11242,N_11528);
nor U12513 (N_12513,N_10128,N_10285);
nor U12514 (N_12514,N_11938,N_9262);
xor U12515 (N_12515,N_9550,N_10364);
xnor U12516 (N_12516,N_10227,N_10546);
or U12517 (N_12517,N_10929,N_9412);
or U12518 (N_12518,N_11006,N_10318);
xnor U12519 (N_12519,N_9818,N_10557);
and U12520 (N_12520,N_9333,N_11643);
nand U12521 (N_12521,N_11212,N_11412);
xnor U12522 (N_12522,N_10908,N_11839);
nor U12523 (N_12523,N_11042,N_9293);
xor U12524 (N_12524,N_9010,N_11804);
xor U12525 (N_12525,N_9898,N_9513);
and U12526 (N_12526,N_10809,N_9938);
xor U12527 (N_12527,N_10421,N_10547);
nand U12528 (N_12528,N_11155,N_11189);
nand U12529 (N_12529,N_9573,N_11016);
nand U12530 (N_12530,N_11634,N_10852);
or U12531 (N_12531,N_10009,N_9482);
and U12532 (N_12532,N_9041,N_9082);
or U12533 (N_12533,N_10616,N_9794);
xor U12534 (N_12534,N_9320,N_11835);
or U12535 (N_12535,N_10985,N_9707);
and U12536 (N_12536,N_9261,N_9391);
nor U12537 (N_12537,N_11695,N_9703);
or U12538 (N_12538,N_10042,N_9770);
or U12539 (N_12539,N_10878,N_10234);
xnor U12540 (N_12540,N_10072,N_10177);
nor U12541 (N_12541,N_10311,N_11268);
nand U12542 (N_12542,N_9249,N_11590);
nor U12543 (N_12543,N_11521,N_10121);
or U12544 (N_12544,N_11724,N_9941);
or U12545 (N_12545,N_9075,N_11971);
and U12546 (N_12546,N_10974,N_9113);
nand U12547 (N_12547,N_11620,N_10231);
and U12548 (N_12548,N_11251,N_9669);
nand U12549 (N_12549,N_9509,N_9188);
and U12550 (N_12550,N_9525,N_9970);
and U12551 (N_12551,N_11059,N_11678);
xor U12552 (N_12552,N_9616,N_10272);
or U12553 (N_12553,N_10110,N_11694);
or U12554 (N_12554,N_11896,N_11380);
nand U12555 (N_12555,N_9361,N_9158);
and U12556 (N_12556,N_11606,N_10347);
or U12557 (N_12557,N_11377,N_10504);
nor U12558 (N_12558,N_10019,N_10049);
nand U12559 (N_12559,N_10527,N_9501);
nand U12560 (N_12560,N_11353,N_10274);
or U12561 (N_12561,N_10265,N_11874);
xor U12562 (N_12562,N_9722,N_9546);
nand U12563 (N_12563,N_9926,N_10178);
nor U12564 (N_12564,N_9417,N_11816);
nor U12565 (N_12565,N_11122,N_10535);
xnor U12566 (N_12566,N_9951,N_10899);
nand U12567 (N_12567,N_9047,N_9360);
nor U12568 (N_12568,N_11675,N_10483);
and U12569 (N_12569,N_11836,N_10192);
nand U12570 (N_12570,N_10926,N_11829);
and U12571 (N_12571,N_10186,N_9910);
and U12572 (N_12572,N_9402,N_11445);
and U12573 (N_12573,N_9849,N_10189);
xor U12574 (N_12574,N_9677,N_9432);
xnor U12575 (N_12575,N_9595,N_11716);
xor U12576 (N_12576,N_11846,N_10499);
xnor U12577 (N_12577,N_9610,N_10920);
and U12578 (N_12578,N_11599,N_9178);
and U12579 (N_12579,N_10703,N_9123);
or U12580 (N_12580,N_9638,N_9544);
and U12581 (N_12581,N_10670,N_10510);
and U12582 (N_12582,N_11081,N_11898);
or U12583 (N_12583,N_11945,N_10413);
nor U12584 (N_12584,N_10298,N_11665);
or U12585 (N_12585,N_10729,N_11570);
or U12586 (N_12586,N_11409,N_11070);
xor U12587 (N_12587,N_11441,N_11197);
nor U12588 (N_12588,N_11142,N_9908);
xor U12589 (N_12589,N_10630,N_10001);
nand U12590 (N_12590,N_10781,N_10464);
nor U12591 (N_12591,N_11554,N_10800);
xnor U12592 (N_12592,N_9101,N_10409);
and U12593 (N_12593,N_11710,N_9774);
nor U12594 (N_12594,N_10839,N_11566);
nor U12595 (N_12595,N_9894,N_10507);
nand U12596 (N_12596,N_9066,N_9464);
or U12597 (N_12597,N_9063,N_10798);
xnor U12598 (N_12598,N_9569,N_9643);
nand U12599 (N_12599,N_9005,N_9574);
xor U12600 (N_12600,N_10890,N_9257);
nand U12601 (N_12601,N_10672,N_11981);
or U12602 (N_12602,N_11623,N_11143);
nand U12603 (N_12603,N_9097,N_9472);
nand U12604 (N_12604,N_10129,N_9740);
or U12605 (N_12605,N_9222,N_9989);
or U12606 (N_12606,N_11559,N_9528);
xnor U12607 (N_12607,N_9983,N_9146);
xor U12608 (N_12608,N_10406,N_11956);
nor U12609 (N_12609,N_9671,N_9238);
and U12610 (N_12610,N_11777,N_10692);
xnor U12611 (N_12611,N_11944,N_9745);
xnor U12612 (N_12612,N_11370,N_11974);
and U12613 (N_12613,N_9141,N_11580);
xor U12614 (N_12614,N_10500,N_10872);
xor U12615 (N_12615,N_10667,N_10157);
or U12616 (N_12616,N_9499,N_9240);
and U12617 (N_12617,N_11727,N_11309);
or U12618 (N_12618,N_11002,N_10437);
nand U12619 (N_12619,N_11692,N_10771);
and U12620 (N_12620,N_10182,N_10315);
nor U12621 (N_12621,N_10886,N_10763);
or U12622 (N_12622,N_9425,N_11076);
or U12623 (N_12623,N_10381,N_11657);
xor U12624 (N_12624,N_10179,N_10736);
nor U12625 (N_12625,N_11043,N_10310);
nand U12626 (N_12626,N_9833,N_11202);
nor U12627 (N_12627,N_11538,N_11625);
and U12628 (N_12628,N_11543,N_10163);
and U12629 (N_12629,N_11740,N_10140);
xnor U12630 (N_12630,N_10368,N_10016);
and U12631 (N_12631,N_9306,N_9929);
or U12632 (N_12632,N_10414,N_9459);
or U12633 (N_12633,N_10748,N_11581);
or U12634 (N_12634,N_9564,N_10099);
nor U12635 (N_12635,N_9437,N_11050);
nor U12636 (N_12636,N_11514,N_10463);
and U12637 (N_12637,N_11391,N_10885);
or U12638 (N_12638,N_9203,N_9328);
and U12639 (N_12639,N_10062,N_11782);
or U12640 (N_12640,N_11387,N_11278);
nand U12641 (N_12641,N_9998,N_11351);
or U12642 (N_12642,N_11860,N_11361);
and U12643 (N_12643,N_10647,N_9729);
xnor U12644 (N_12644,N_10086,N_11824);
xnor U12645 (N_12645,N_10680,N_11037);
xnor U12646 (N_12646,N_9975,N_11598);
xor U12647 (N_12647,N_11720,N_10394);
and U12648 (N_12648,N_9184,N_9944);
or U12649 (N_12649,N_9008,N_11869);
nand U12650 (N_12650,N_10206,N_11879);
or U12651 (N_12651,N_9286,N_9032);
nor U12652 (N_12652,N_9662,N_9647);
nor U12653 (N_12653,N_11810,N_9422);
xor U12654 (N_12654,N_9684,N_11761);
nor U12655 (N_12655,N_9959,N_10734);
and U12656 (N_12656,N_10959,N_10774);
nor U12657 (N_12657,N_10351,N_9687);
nor U12658 (N_12658,N_9783,N_9124);
nand U12659 (N_12659,N_9813,N_9739);
nand U12660 (N_12660,N_10134,N_10370);
and U12661 (N_12661,N_9541,N_11437);
nor U12662 (N_12662,N_10583,N_10173);
nor U12663 (N_12663,N_10032,N_11713);
or U12664 (N_12664,N_11153,N_9584);
or U12665 (N_12665,N_9183,N_11256);
or U12666 (N_12666,N_10369,N_10011);
and U12667 (N_12667,N_10191,N_9185);
and U12668 (N_12668,N_10842,N_9230);
and U12669 (N_12669,N_9560,N_10825);
xnor U12670 (N_12670,N_10904,N_10108);
and U12671 (N_12671,N_9905,N_11624);
nand U12672 (N_12672,N_9474,N_11968);
nand U12673 (N_12673,N_9162,N_11615);
nand U12674 (N_12674,N_10493,N_9629);
nand U12675 (N_12675,N_9370,N_10171);
or U12676 (N_12676,N_11390,N_10776);
and U12677 (N_12677,N_10276,N_10584);
and U12678 (N_12678,N_11772,N_10664);
nor U12679 (N_12679,N_11723,N_9583);
and U12680 (N_12680,N_11684,N_9934);
xnor U12681 (N_12681,N_10962,N_11258);
nor U12682 (N_12682,N_9277,N_9443);
nor U12683 (N_12683,N_10020,N_10769);
xor U12684 (N_12684,N_11520,N_11610);
nand U12685 (N_12685,N_10441,N_11120);
xor U12686 (N_12686,N_11996,N_11128);
nor U12687 (N_12687,N_10211,N_10709);
or U12688 (N_12688,N_11399,N_11611);
nand U12689 (N_12689,N_11373,N_10730);
and U12690 (N_12690,N_10063,N_10943);
nor U12691 (N_12691,N_11205,N_10586);
and U12692 (N_12692,N_9673,N_9429);
nor U12693 (N_12693,N_9057,N_11460);
xor U12694 (N_12694,N_9930,N_10945);
or U12695 (N_12695,N_11729,N_10228);
and U12696 (N_12696,N_10484,N_10259);
nand U12697 (N_12697,N_11783,N_11198);
xnor U12698 (N_12698,N_9811,N_9787);
xor U12699 (N_12699,N_9681,N_11347);
nor U12700 (N_12700,N_9187,N_10984);
nor U12701 (N_12701,N_9702,N_9748);
or U12702 (N_12702,N_11201,N_10541);
nor U12703 (N_12703,N_11225,N_9889);
nor U12704 (N_12704,N_11104,N_9936);
xor U12705 (N_12705,N_11630,N_9548);
nor U12706 (N_12706,N_9343,N_11337);
xnor U12707 (N_12707,N_10526,N_11722);
or U12708 (N_12708,N_10111,N_11023);
nor U12709 (N_12709,N_10548,N_10577);
nor U12710 (N_12710,N_11966,N_11154);
or U12711 (N_12711,N_10397,N_11884);
nor U12712 (N_12712,N_10112,N_9969);
nor U12713 (N_12713,N_11797,N_10808);
and U12714 (N_12714,N_11850,N_10768);
xor U12715 (N_12715,N_10149,N_11031);
or U12716 (N_12716,N_11401,N_9994);
nand U12717 (N_12717,N_11364,N_9260);
and U12718 (N_12718,N_10090,N_11830);
or U12719 (N_12719,N_9334,N_11587);
nor U12720 (N_12720,N_10756,N_11867);
or U12721 (N_12721,N_9756,N_9288);
nand U12722 (N_12722,N_10733,N_11190);
nand U12723 (N_12723,N_10660,N_10988);
nor U12724 (N_12724,N_11436,N_11669);
xor U12725 (N_12725,N_11435,N_10415);
xor U12726 (N_12726,N_10309,N_11431);
xor U12727 (N_12727,N_11250,N_9798);
xor U12728 (N_12728,N_10371,N_11993);
or U12729 (N_12729,N_10004,N_10912);
and U12730 (N_12730,N_11702,N_9050);
nor U12731 (N_12731,N_11467,N_11717);
xnor U12732 (N_12732,N_10740,N_11262);
or U12733 (N_12733,N_10708,N_11558);
or U12734 (N_12734,N_10055,N_11273);
xnor U12735 (N_12735,N_10752,N_9362);
xnor U12736 (N_12736,N_11768,N_11108);
nand U12737 (N_12737,N_9822,N_10352);
and U12738 (N_12738,N_11948,N_10339);
nor U12739 (N_12739,N_11807,N_10382);
and U12740 (N_12740,N_11654,N_11405);
nand U12741 (N_12741,N_11181,N_11718);
or U12742 (N_12742,N_10482,N_9688);
nor U12743 (N_12743,N_9026,N_11228);
or U12744 (N_12744,N_10402,N_9446);
nor U12745 (N_12745,N_11321,N_11961);
nand U12746 (N_12746,N_9680,N_11014);
and U12747 (N_12747,N_10634,N_11806);
and U12748 (N_12748,N_10608,N_11429);
xor U12749 (N_12749,N_10975,N_10644);
or U12750 (N_12750,N_11263,N_10939);
and U12751 (N_12751,N_10026,N_10107);
xnor U12752 (N_12752,N_9340,N_9076);
and U12753 (N_12753,N_9987,N_11166);
or U12754 (N_12754,N_9587,N_10874);
nand U12755 (N_12755,N_11324,N_11296);
or U12756 (N_12756,N_9502,N_9458);
nand U12757 (N_12757,N_10688,N_11350);
and U12758 (N_12758,N_11679,N_10796);
nor U12759 (N_12759,N_11878,N_10387);
or U12760 (N_12760,N_11897,N_10060);
and U12761 (N_12761,N_9455,N_11498);
or U12762 (N_12762,N_11449,N_11144);
and U12763 (N_12763,N_10349,N_9136);
or U12764 (N_12764,N_11577,N_10791);
or U12765 (N_12765,N_11447,N_11244);
nand U12766 (N_12766,N_9773,N_10329);
nand U12767 (N_12767,N_10479,N_11899);
nand U12768 (N_12768,N_10947,N_9494);
and U12769 (N_12769,N_10467,N_10428);
nand U12770 (N_12770,N_11330,N_11109);
and U12771 (N_12771,N_11093,N_11656);
or U12772 (N_12772,N_10855,N_11229);
nor U12773 (N_12773,N_10282,N_10558);
nand U12774 (N_12774,N_9508,N_11504);
xor U12775 (N_12775,N_9394,N_9336);
nor U12776 (N_12776,N_11827,N_11627);
nand U12777 (N_12777,N_9734,N_10217);
xor U12778 (N_12778,N_9442,N_11239);
xnor U12779 (N_12779,N_10656,N_9218);
nor U12780 (N_12780,N_11892,N_9058);
or U12781 (N_12781,N_11859,N_11779);
xor U12782 (N_12782,N_11658,N_11238);
nand U12783 (N_12783,N_11909,N_11802);
xor U12784 (N_12784,N_9383,N_11428);
or U12785 (N_12785,N_9516,N_10133);
nor U12786 (N_12786,N_10977,N_9593);
nor U12787 (N_12787,N_9527,N_10799);
or U12788 (N_12788,N_11967,N_9298);
nand U12789 (N_12789,N_11452,N_10731);
nor U12790 (N_12790,N_11600,N_11439);
nand U12791 (N_12791,N_9626,N_11735);
xnor U12792 (N_12792,N_11173,N_10700);
xor U12793 (N_12793,N_9198,N_9803);
xnor U12794 (N_12794,N_10041,N_9214);
nor U12795 (N_12795,N_10299,N_10979);
nor U12796 (N_12796,N_10674,N_9247);
or U12797 (N_12797,N_11187,N_10818);
nand U12798 (N_12798,N_9229,N_11734);
nand U12799 (N_12799,N_9503,N_9363);
nor U12800 (N_12800,N_9512,N_10202);
nor U12801 (N_12801,N_11796,N_10448);
or U12802 (N_12802,N_10881,N_10169);
or U12803 (N_12803,N_9591,N_10264);
xor U12804 (N_12804,N_11457,N_10662);
and U12805 (N_12805,N_11113,N_9488);
nand U12806 (N_12806,N_10021,N_9000);
and U12807 (N_12807,N_9467,N_10815);
xnor U12808 (N_12808,N_9725,N_11087);
nor U12809 (N_12809,N_10677,N_11857);
xor U12810 (N_12810,N_10181,N_11612);
nor U12811 (N_12811,N_9077,N_10827);
nor U12812 (N_12812,N_9846,N_9566);
xnor U12813 (N_12813,N_10333,N_9134);
and U12814 (N_12814,N_9906,N_10509);
nand U12815 (N_12815,N_10079,N_11529);
and U12816 (N_12816,N_10749,N_11126);
and U12817 (N_12817,N_11545,N_11905);
or U12818 (N_12818,N_9915,N_10279);
nand U12819 (N_12819,N_10580,N_11260);
or U12820 (N_12820,N_10880,N_9155);
nand U12821 (N_12821,N_10334,N_11359);
xor U12822 (N_12822,N_10790,N_9705);
nor U12823 (N_12823,N_10237,N_11952);
nor U12824 (N_12824,N_9171,N_10200);
and U12825 (N_12825,N_9090,N_10195);
or U12826 (N_12826,N_10506,N_10286);
xnor U12827 (N_12827,N_10293,N_9451);
or U12828 (N_12828,N_9315,N_11681);
and U12829 (N_12829,N_10502,N_11595);
nor U12830 (N_12830,N_9801,N_10337);
or U12831 (N_12831,N_11601,N_10268);
nor U12832 (N_12832,N_10995,N_9530);
and U12833 (N_12833,N_9986,N_10528);
and U12834 (N_12834,N_9654,N_10575);
nor U12835 (N_12835,N_11838,N_11483);
nor U12836 (N_12836,N_9605,N_10597);
or U12837 (N_12837,N_9021,N_10069);
nor U12838 (N_12838,N_11597,N_11222);
xnor U12839 (N_12839,N_11989,N_11018);
nor U12840 (N_12840,N_9406,N_11642);
xor U12841 (N_12841,N_11069,N_9307);
or U12842 (N_12842,N_11146,N_10783);
nor U12843 (N_12843,N_9400,N_10296);
nor U12844 (N_12844,N_9854,N_9639);
or U12845 (N_12845,N_9368,N_10767);
nand U12846 (N_12846,N_10399,N_10524);
nand U12847 (N_12847,N_9828,N_10061);
or U12848 (N_12848,N_9498,N_11286);
xor U12849 (N_12849,N_10987,N_9031);
nand U12850 (N_12850,N_9250,N_10017);
nand U12851 (N_12851,N_11672,N_10562);
xor U12852 (N_12852,N_11249,N_9327);
and U12853 (N_12853,N_11458,N_11817);
nor U12854 (N_12854,N_10162,N_11609);
and U12855 (N_12855,N_9111,N_10934);
xnor U12856 (N_12856,N_9505,N_11714);
nor U12857 (N_12857,N_11628,N_9350);
or U12858 (N_12858,N_10681,N_9793);
nor U12859 (N_12859,N_10909,N_9294);
nor U12860 (N_12860,N_11533,N_9949);
xor U12861 (N_12861,N_11385,N_10570);
nor U12862 (N_12862,N_10848,N_9434);
nand U12863 (N_12863,N_10963,N_10529);
nor U12864 (N_12864,N_11451,N_10335);
nand U12865 (N_12865,N_11584,N_9668);
xnor U12866 (N_12866,N_10338,N_10699);
xor U12867 (N_12867,N_11227,N_10442);
and U12868 (N_12868,N_9048,N_9064);
nor U12869 (N_12869,N_10517,N_9992);
xor U12870 (N_12870,N_10942,N_9631);
or U12871 (N_12871,N_10993,N_9859);
nand U12872 (N_12872,N_9965,N_9301);
nor U12873 (N_12873,N_11466,N_11096);
xor U12874 (N_12874,N_11366,N_11730);
xor U12875 (N_12875,N_9011,N_10214);
or U12876 (N_12876,N_10051,N_10271);
nand U12877 (N_12877,N_10355,N_9830);
xnor U12878 (N_12878,N_11841,N_9752);
or U12879 (N_12879,N_10008,N_10568);
nand U12880 (N_12880,N_10877,N_11765);
xor U12881 (N_12881,N_10641,N_11650);
nand U12882 (N_12882,N_9627,N_11275);
and U12883 (N_12883,N_9197,N_11918);
and U12884 (N_12884,N_9863,N_10849);
nand U12885 (N_12885,N_11411,N_9117);
nand U12886 (N_12886,N_9118,N_9634);
or U12887 (N_12887,N_10706,N_11589);
nor U12888 (N_12888,N_9152,N_11639);
and U12889 (N_12889,N_11920,N_11755);
nor U12890 (N_12890,N_9771,N_11421);
nor U12891 (N_12891,N_10447,N_10127);
nor U12892 (N_12892,N_9398,N_11700);
nand U12893 (N_12893,N_11696,N_11848);
and U12894 (N_12894,N_9216,N_10614);
or U12895 (N_12895,N_9447,N_10859);
or U12896 (N_12896,N_10960,N_9232);
xnor U12897 (N_12897,N_10896,N_11762);
nor U12898 (N_12898,N_11496,N_9885);
nor U12899 (N_12899,N_10538,N_9716);
nand U12900 (N_12900,N_9445,N_9481);
or U12901 (N_12901,N_11988,N_10693);
nand U12902 (N_12902,N_9252,N_11688);
nor U12903 (N_12903,N_9196,N_9754);
xor U12904 (N_12904,N_9476,N_9609);
nor U12905 (N_12905,N_9259,N_10319);
nand U12906 (N_12906,N_11480,N_10288);
xnor U12907 (N_12907,N_10431,N_11515);
nand U12908 (N_12908,N_11842,N_10059);
and U12909 (N_12909,N_10559,N_9607);
nor U12910 (N_12910,N_9084,N_10175);
nor U12911 (N_12911,N_10986,N_9628);
nand U12912 (N_12912,N_11091,N_11929);
xor U12913 (N_12913,N_10253,N_11171);
and U12914 (N_12914,N_11298,N_11394);
or U12915 (N_12915,N_9622,N_9074);
xor U12916 (N_12916,N_9235,N_9003);
xnor U12917 (N_12917,N_9281,N_11573);
nor U12918 (N_12918,N_11024,N_9108);
or U12919 (N_12919,N_10589,N_10961);
and U12920 (N_12920,N_9769,N_9988);
and U12921 (N_12921,N_11152,N_11379);
or U12922 (N_12922,N_10472,N_9630);
and U12923 (N_12923,N_10139,N_9309);
or U12924 (N_12924,N_11919,N_10126);
or U12925 (N_12925,N_10468,N_9321);
nand U12926 (N_12926,N_11552,N_11660);
nor U12927 (N_12927,N_10052,N_11141);
or U12928 (N_12928,N_11174,N_11025);
and U12929 (N_12929,N_11618,N_10056);
or U12930 (N_12930,N_10953,N_9098);
or U12931 (N_12931,N_9022,N_9985);
nand U12932 (N_12932,N_11471,N_11075);
nor U12933 (N_12933,N_10957,N_9637);
nor U12934 (N_12934,N_11346,N_10488);
nand U12935 (N_12935,N_9241,N_11709);
xor U12936 (N_12936,N_9389,N_9371);
nand U12937 (N_12937,N_10923,N_9393);
xnor U12938 (N_12938,N_9955,N_9646);
and U12939 (N_12939,N_11851,N_9718);
nand U12940 (N_12940,N_9810,N_11542);
xor U12941 (N_12941,N_10066,N_9382);
and U12942 (N_12942,N_11179,N_10188);
or U12943 (N_12943,N_11184,N_10830);
nor U12944 (N_12944,N_9750,N_9553);
nand U12945 (N_12945,N_11406,N_9132);
xor U12946 (N_12946,N_9416,N_11240);
or U12947 (N_12947,N_9867,N_9824);
nand U12948 (N_12948,N_11425,N_10810);
nor U12949 (N_12949,N_9730,N_9397);
or U12950 (N_12950,N_10114,N_10944);
or U12951 (N_12951,N_11132,N_11446);
xor U12952 (N_12952,N_10824,N_11509);
xnor U12953 (N_12953,N_10679,N_10835);
nand U12954 (N_12954,N_10328,N_9844);
and U12955 (N_12955,N_10225,N_9717);
nand U12956 (N_12956,N_9305,N_9522);
and U12957 (N_12957,N_11072,N_9314);
nand U12958 (N_12958,N_10080,N_10501);
and U12959 (N_12959,N_10305,N_9825);
and U12960 (N_12960,N_9690,N_9356);
and U12961 (N_12961,N_11433,N_11019);
nor U12962 (N_12962,N_11328,N_11667);
nand U12963 (N_12963,N_11563,N_10613);
nor U12964 (N_12964,N_10340,N_9112);
nor U12965 (N_12965,N_9044,N_9297);
and U12966 (N_12966,N_10902,N_9093);
or U12967 (N_12967,N_9166,N_10582);
and U12968 (N_12968,N_10531,N_11764);
nor U12969 (N_12969,N_10336,N_9719);
nand U12970 (N_12970,N_11943,N_11736);
and U12971 (N_12971,N_9282,N_10359);
and U12972 (N_12972,N_10514,N_11607);
nand U12973 (N_12973,N_9409,N_10543);
xor U12974 (N_12974,N_11066,N_10427);
nand U12975 (N_12975,N_9480,N_9552);
nand U12976 (N_12976,N_11417,N_9151);
nor U12977 (N_12977,N_11356,N_10105);
or U12978 (N_12978,N_11491,N_10607);
and U12979 (N_12979,N_11503,N_11549);
and U12980 (N_12980,N_11790,N_11629);
xor U12981 (N_12981,N_9855,N_10458);
or U12982 (N_12982,N_9841,N_9319);
and U12983 (N_12983,N_9645,N_10585);
nor U12984 (N_12984,N_9655,N_11397);
nor U12985 (N_12985,N_11616,N_9329);
nor U12986 (N_12986,N_10556,N_11344);
and U12987 (N_12987,N_11287,N_11319);
xnor U12988 (N_12988,N_9720,N_11148);
xor U12989 (N_12989,N_11500,N_9143);
nor U12990 (N_12990,N_11230,N_10491);
and U12991 (N_12991,N_9621,N_11192);
nand U12992 (N_12992,N_10860,N_9663);
and U12993 (N_12993,N_11270,N_10275);
nand U12994 (N_12994,N_9161,N_11254);
or U12995 (N_12995,N_9191,N_9266);
nand U12996 (N_12996,N_11281,N_11646);
or U12997 (N_12997,N_10380,N_9790);
nor U12998 (N_12998,N_9109,N_10322);
nand U12999 (N_12999,N_10190,N_11770);
nor U13000 (N_13000,N_10461,N_10633);
or U13001 (N_13001,N_11550,N_9598);
and U13002 (N_13002,N_9357,N_11300);
and U13003 (N_13003,N_10895,N_10924);
xor U13004 (N_13004,N_9731,N_10751);
and U13005 (N_13005,N_11854,N_11311);
nand U13006 (N_13006,N_11272,N_9207);
xor U13007 (N_13007,N_10003,N_11026);
nor U13008 (N_13008,N_10006,N_9311);
nand U13009 (N_13009,N_11035,N_11074);
and U13010 (N_13010,N_11902,N_9912);
and U13011 (N_13011,N_10386,N_11579);
nand U13012 (N_13012,N_10534,N_10495);
xor U13013 (N_13013,N_10065,N_10132);
xnor U13014 (N_13014,N_9963,N_9640);
nor U13015 (N_13015,N_9493,N_9226);
xor U13016 (N_13016,N_11333,N_11049);
or U13017 (N_13017,N_11004,N_10456);
or U13018 (N_13018,N_9223,N_9060);
and U13019 (N_13019,N_11954,N_9577);
or U13020 (N_13020,N_11204,N_11339);
or U13021 (N_13021,N_10905,N_11876);
xnor U13022 (N_13022,N_11207,N_10841);
and U13023 (N_13023,N_9233,N_10395);
or U13024 (N_13024,N_10233,N_10156);
nand U13025 (N_13025,N_11305,N_10216);
nand U13026 (N_13026,N_10598,N_11862);
xnor U13027 (N_13027,N_11711,N_10719);
nand U13028 (N_13028,N_10496,N_11991);
xor U13029 (N_13029,N_11335,N_9757);
and U13030 (N_13030,N_9435,N_11261);
xor U13031 (N_13031,N_10965,N_9845);
and U13032 (N_13032,N_10257,N_11490);
and U13033 (N_13033,N_10578,N_10950);
nand U13034 (N_13034,N_10626,N_9219);
nand U13035 (N_13035,N_11513,N_11863);
xnor U13036 (N_13036,N_10023,N_9396);
nand U13037 (N_13037,N_10789,N_11299);
or U13038 (N_13038,N_11998,N_10477);
nand U13039 (N_13039,N_11180,N_10643);
nand U13040 (N_13040,N_9388,N_9202);
and U13041 (N_13041,N_10373,N_9887);
nor U13042 (N_13042,N_11766,N_11415);
and U13043 (N_13043,N_10457,N_10375);
or U13044 (N_13044,N_11564,N_10058);
or U13045 (N_13045,N_9135,N_11732);
and U13046 (N_13046,N_11253,N_10445);
nor U13047 (N_13047,N_10172,N_11537);
and U13048 (N_13048,N_10084,N_11284);
nand U13049 (N_13049,N_11685,N_11721);
and U13050 (N_13050,N_9007,N_11468);
or U13051 (N_13051,N_10044,N_9689);
nor U13052 (N_13052,N_10466,N_9683);
nand U13053 (N_13053,N_10075,N_11633);
or U13054 (N_13054,N_10018,N_10941);
xnor U13055 (N_13055,N_11726,N_9779);
xor U13056 (N_13056,N_10455,N_10154);
xor U13057 (N_13057,N_10242,N_9644);
nor U13058 (N_13058,N_10037,N_10197);
xnor U13059 (N_13059,N_9504,N_10376);
nor U13060 (N_13060,N_9860,N_9212);
xnor U13061 (N_13061,N_11200,N_11704);
xor U13062 (N_13062,N_9221,N_10936);
and U13063 (N_13063,N_9708,N_10444);
and U13064 (N_13064,N_9611,N_9153);
nor U13065 (N_13065,N_9038,N_10378);
nor U13066 (N_13066,N_9641,N_9256);
nor U13067 (N_13067,N_10836,N_11963);
nand U13068 (N_13068,N_11477,N_11168);
nand U13069 (N_13069,N_11631,N_9159);
nand U13070 (N_13070,N_9035,N_11818);
xnor U13071 (N_13071,N_9133,N_9271);
and U13072 (N_13072,N_10915,N_10854);
nand U13073 (N_13073,N_11420,N_10735);
nor U13074 (N_13074,N_11360,N_9243);
and U13075 (N_13075,N_10096,N_10785);
nand U13076 (N_13076,N_11947,N_9448);
xnor U13077 (N_13077,N_11760,N_9190);
xor U13078 (N_13078,N_10635,N_10405);
and U13079 (N_13079,N_11418,N_9042);
xor U13080 (N_13080,N_9114,N_9033);
nor U13081 (N_13081,N_10657,N_9554);
or U13082 (N_13082,N_11223,N_10198);
nand U13083 (N_13083,N_11213,N_11313);
and U13084 (N_13084,N_9242,N_11773);
nand U13085 (N_13085,N_11131,N_11094);
xor U13086 (N_13086,N_10868,N_9415);
or U13087 (N_13087,N_9724,N_11413);
or U13088 (N_13088,N_10404,N_10316);
xnor U13089 (N_13089,N_9510,N_9201);
and U13090 (N_13090,N_11556,N_11475);
and U13091 (N_13091,N_9839,N_10153);
and U13092 (N_13092,N_9079,N_11571);
and U13093 (N_13093,N_11525,N_10666);
xor U13094 (N_13094,N_10685,N_9440);
nor U13095 (N_13095,N_10357,N_9551);
xnor U13096 (N_13096,N_9325,N_10610);
nand U13097 (N_13097,N_10919,N_10779);
or U13098 (N_13098,N_11177,N_9600);
nor U13099 (N_13099,N_11352,N_9299);
xor U13100 (N_13100,N_11670,N_11100);
or U13101 (N_13101,N_9788,N_11167);
or U13102 (N_13102,N_11224,N_9534);
xnor U13103 (N_13103,N_9979,N_10817);
and U13104 (N_13104,N_11655,N_9086);
or U13105 (N_13105,N_11621,N_9210);
nor U13106 (N_13106,N_10289,N_11252);
or U13107 (N_13107,N_10620,N_11507);
nor U13108 (N_13108,N_9517,N_11586);
nand U13109 (N_13109,N_10164,N_11973);
or U13110 (N_13110,N_11499,N_9263);
nand U13111 (N_13111,N_10697,N_10866);
nor U13112 (N_13112,N_11926,N_9353);
and U13113 (N_13113,N_11039,N_11139);
and U13114 (N_13114,N_11265,N_9051);
nor U13115 (N_13115,N_9220,N_11776);
nor U13116 (N_13116,N_9764,N_11555);
or U13117 (N_13117,N_10240,N_9436);
nand U13118 (N_13118,N_11962,N_9547);
nor U13119 (N_13119,N_11693,N_9874);
xor U13120 (N_13120,N_11791,N_10784);
nor U13121 (N_13121,N_10549,N_10601);
nor U13122 (N_13122,N_11193,N_9182);
xor U13123 (N_13123,N_11488,N_9349);
xnor U13124 (N_13124,N_9004,N_11013);
xor U13125 (N_13125,N_10147,N_11826);
or U13126 (N_13126,N_10628,N_11640);
and U13127 (N_13127,N_11389,N_11172);
xor U13128 (N_13128,N_11266,N_10536);
nor U13129 (N_13129,N_10983,N_10512);
xor U13130 (N_13130,N_9861,N_10683);
or U13131 (N_13131,N_10031,N_9254);
or U13132 (N_13132,N_10301,N_11572);
and U13133 (N_13133,N_10374,N_10400);
nand U13134 (N_13134,N_10561,N_10416);
nor U13135 (N_13135,N_10385,N_9791);
xor U13136 (N_13136,N_11750,N_11975);
nand U13137 (N_13137,N_11133,N_11064);
nand U13138 (N_13138,N_9778,N_9895);
or U13139 (N_13139,N_10879,N_11482);
nor U13140 (N_13140,N_11501,N_11865);
nand U13141 (N_13141,N_9213,N_9386);
and U13142 (N_13142,N_10012,N_9489);
and U13143 (N_13143,N_9102,N_11746);
nand U13144 (N_13144,N_9149,N_10435);
nor U13145 (N_13145,N_10805,N_9441);
nand U13146 (N_13146,N_10592,N_11414);
nor U13147 (N_13147,N_11664,N_11939);
xor U13148 (N_13148,N_10303,N_11535);
and U13149 (N_13149,N_9258,N_11914);
and U13150 (N_13150,N_9686,N_11183);
or U13151 (N_13151,N_9418,N_10082);
xor U13152 (N_13152,N_10823,N_11705);
nand U13153 (N_13153,N_9746,N_11781);
and U13154 (N_13154,N_9145,N_10342);
nor U13155 (N_13155,N_11124,N_9956);
xnor U13156 (N_13156,N_11699,N_9419);
xnor U13157 (N_13157,N_11479,N_11485);
nand U13158 (N_13158,N_9694,N_10958);
and U13159 (N_13159,N_9366,N_11114);
or U13160 (N_13160,N_11073,N_10678);
nor U13161 (N_13161,N_9535,N_10829);
and U13162 (N_13162,N_11638,N_9172);
and U13163 (N_13163,N_10167,N_10663);
or U13164 (N_13164,N_10893,N_10632);
or U13165 (N_13165,N_11226,N_11994);
and U13166 (N_13166,N_10794,N_10615);
and U13167 (N_13167,N_9710,N_10267);
xor U13168 (N_13168,N_9749,N_9037);
xnor U13169 (N_13169,N_11419,N_9040);
nand U13170 (N_13170,N_11831,N_10533);
or U13171 (N_13171,N_11071,N_9865);
nor U13172 (N_13172,N_9843,N_10704);
and U13173 (N_13173,N_9800,N_10124);
xnor U13174 (N_13174,N_10968,N_11979);
xor U13175 (N_13175,N_11077,N_11121);
and U13176 (N_13176,N_10618,N_10014);
nor U13177 (N_13177,N_9316,N_10687);
nor U13178 (N_13178,N_11288,N_9330);
nand U13179 (N_13179,N_10489,N_11316);
nand U13180 (N_13180,N_11317,N_11738);
or U13181 (N_13181,N_9581,N_9981);
nand U13182 (N_13182,N_9542,N_11649);
or U13183 (N_13183,N_9886,N_11246);
and U13184 (N_13184,N_10843,N_11924);
and U13185 (N_13185,N_10473,N_10871);
xor U13186 (N_13186,N_9901,N_11487);
or U13187 (N_13187,N_10910,N_11332);
nand U13188 (N_13188,N_11868,N_10151);
or U13189 (N_13189,N_11186,N_9275);
nand U13190 (N_13190,N_9344,N_10481);
xor U13191 (N_13191,N_10419,N_9078);
nor U13192 (N_13192,N_10280,N_11527);
nor U13193 (N_13193,N_9890,N_10115);
nor U13194 (N_13194,N_10850,N_10354);
nand U13195 (N_13195,N_9802,N_9189);
and U13196 (N_13196,N_9470,N_10951);
or U13197 (N_13197,N_10203,N_9072);
or U13198 (N_13198,N_10109,N_11323);
or U13199 (N_13199,N_10423,N_11666);
nor U13200 (N_13200,N_10786,N_9692);
or U13201 (N_13201,N_9612,N_10665);
xnor U13202 (N_13202,N_9808,N_9420);
nor U13203 (N_13203,N_11575,N_11803);
and U13204 (N_13204,N_10141,N_10160);
nor U13205 (N_13205,N_9636,N_11303);
nor U13206 (N_13206,N_11588,N_11010);
nand U13207 (N_13207,N_10897,N_9507);
nand U13208 (N_13208,N_11206,N_11526);
xnor U13209 (N_13209,N_11531,N_10116);
nand U13210 (N_13210,N_9721,N_10659);
nand U13211 (N_13211,N_9444,N_9034);
or U13212 (N_13212,N_9911,N_11825);
or U13213 (N_13213,N_11331,N_9537);
or U13214 (N_13214,N_10652,N_11086);
xnor U13215 (N_13215,N_10732,N_9606);
xor U13216 (N_13216,N_11241,N_9872);
or U13217 (N_13217,N_10258,N_10088);
and U13218 (N_13218,N_9065,N_9765);
xnor U13219 (N_13219,N_9847,N_11532);
nand U13220 (N_13220,N_9179,N_11900);
and U13221 (N_13221,N_9916,N_9806);
and U13222 (N_13222,N_11341,N_9401);
or U13223 (N_13223,N_9836,N_11936);
xnor U13224 (N_13224,N_11085,N_9326);
nand U13225 (N_13225,N_9807,N_11217);
nor U13226 (N_13226,N_9120,N_11029);
nand U13227 (N_13227,N_9036,N_9374);
nor U13228 (N_13228,N_10648,N_9130);
nand U13229 (N_13229,N_9107,N_11362);
nand U13230 (N_13230,N_10313,N_9285);
and U13231 (N_13231,N_10007,N_10393);
nor U13232 (N_13232,N_9351,N_9567);
nand U13233 (N_13233,N_9272,N_10650);
xor U13234 (N_13234,N_11594,N_10010);
nor U13235 (N_13235,N_9300,N_10388);
nand U13236 (N_13236,N_11828,N_11582);
nand U13237 (N_13237,N_9727,N_10235);
nor U13238 (N_13238,N_11047,N_10446);
and U13239 (N_13239,N_9877,N_11454);
or U13240 (N_13240,N_11739,N_10639);
and U13241 (N_13241,N_10801,N_10658);
xor U13242 (N_13242,N_9215,N_9999);
nand U13243 (N_13243,N_10989,N_10270);
nand U13244 (N_13244,N_10085,N_10718);
or U13245 (N_13245,N_11506,N_9027);
or U13246 (N_13246,N_9642,N_11903);
nor U13247 (N_13247,N_10350,N_11098);
nor U13248 (N_13248,N_10306,N_10353);
nor U13249 (N_13249,N_10487,N_11530);
and U13250 (N_13250,N_11243,N_10508);
xor U13251 (N_13251,N_10168,N_9657);
nand U13252 (N_13252,N_10092,N_11375);
nand U13253 (N_13253,N_10101,N_10226);
xor U13254 (N_13254,N_11022,N_11099);
xor U13255 (N_13255,N_9106,N_9142);
nand U13256 (N_13256,N_9046,N_9903);
and U13257 (N_13257,N_10199,N_10219);
nand U13258 (N_13258,N_11565,N_11743);
nand U13259 (N_13259,N_9888,N_11388);
nor U13260 (N_13260,N_9424,N_10451);
nand U13261 (N_13261,N_9454,N_10465);
xor U13262 (N_13262,N_11940,N_9369);
or U13263 (N_13263,N_11368,N_11885);
or U13264 (N_13264,N_9997,N_9205);
nor U13265 (N_13265,N_9820,N_10224);
and U13266 (N_13266,N_11950,N_9367);
nand U13267 (N_13267,N_10544,N_11845);
nand U13268 (N_13268,N_11661,N_9767);
nand U13269 (N_13269,N_11910,N_9751);
nor U13270 (N_13270,N_11092,N_10365);
or U13271 (N_13271,N_11911,N_9947);
and U13272 (N_13272,N_9585,N_10844);
or U13273 (N_13273,N_11647,N_10938);
xnor U13274 (N_13274,N_10295,N_9982);
or U13275 (N_13275,N_10758,N_11381);
nor U13276 (N_13276,N_10426,N_9225);
xnor U13277 (N_13277,N_9456,N_11977);
or U13278 (N_13278,N_10236,N_11112);
or U13279 (N_13279,N_9660,N_10430);
or U13280 (N_13280,N_10741,N_9290);
nand U13281 (N_13281,N_9059,N_11744);
nor U13282 (N_13282,N_11378,N_9147);
nand U13283 (N_13283,N_9384,N_11188);
nor U13284 (N_13284,N_9920,N_10246);
nand U13285 (N_13285,N_11176,N_11175);
xor U13286 (N_13286,N_10930,N_11882);
and U13287 (N_13287,N_10478,N_9289);
xnor U13288 (N_13288,N_11969,N_9823);
and U13289 (N_13289,N_11349,N_10675);
nand U13290 (N_13290,N_9856,N_11987);
xor U13291 (N_13291,N_10935,N_11216);
nand U13292 (N_13292,N_10566,N_9736);
xor U13293 (N_13293,N_10158,N_10847);
or U13294 (N_13294,N_10669,N_10906);
and U13295 (N_13295,N_9119,N_10925);
or U13296 (N_13296,N_10261,N_9974);
and U13297 (N_13297,N_9217,N_11068);
or U13298 (N_13298,N_10747,N_10759);
xor U13299 (N_13299,N_11285,N_11872);
nand U13300 (N_13300,N_10106,N_11733);
and U13301 (N_13301,N_9518,N_10857);
or U13302 (N_13302,N_10737,N_10690);
xor U13303 (N_13303,N_10876,N_9483);
nor U13304 (N_13304,N_10701,N_11676);
and U13305 (N_13305,N_10918,N_11084);
nand U13306 (N_13306,N_11000,N_10540);
and U13307 (N_13307,N_9656,N_9942);
or U13308 (N_13308,N_10804,N_10980);
and U13309 (N_13309,N_11562,N_9768);
xor U13310 (N_13310,N_10155,N_11972);
xor U13311 (N_13311,N_10379,N_11312);
and U13312 (N_13312,N_9613,N_9125);
and U13313 (N_13313,N_11088,N_9596);
nor U13314 (N_13314,N_9234,N_11233);
or U13315 (N_13315,N_9880,N_11840);
nor U13316 (N_13316,N_10537,N_11585);
xor U13317 (N_13317,N_10143,N_9840);
nor U13318 (N_13318,N_10787,N_9387);
and U13319 (N_13319,N_9797,N_11703);
or U13320 (N_13320,N_11873,N_9025);
nor U13321 (N_13321,N_10973,N_11438);
nand U13322 (N_13322,N_11983,N_11345);
or U13323 (N_13323,N_9592,N_11157);
xnor U13324 (N_13324,N_9403,N_10840);
and U13325 (N_13325,N_10832,N_9651);
or U13326 (N_13326,N_10485,N_10976);
or U13327 (N_13327,N_9380,N_9423);
nor U13328 (N_13328,N_10250,N_11976);
xor U13329 (N_13329,N_11751,N_11904);
or U13330 (N_13330,N_11398,N_10475);
nand U13331 (N_13331,N_9180,N_11009);
and U13332 (N_13332,N_10811,N_9619);
nor U13333 (N_13333,N_10453,N_9055);
nor U13334 (N_13334,N_11519,N_10034);
or U13335 (N_13335,N_9570,N_9995);
and U13336 (N_13336,N_11374,N_10996);
xnor U13337 (N_13337,N_11210,N_9817);
xnor U13338 (N_13338,N_11481,N_11958);
nand U13339 (N_13339,N_9892,N_11102);
nand U13340 (N_13340,N_11894,N_11970);
nor U13341 (N_13341,N_9837,N_9772);
xnor U13342 (N_13342,N_9094,N_10358);
or U13343 (N_13343,N_11355,N_11512);
xor U13344 (N_13344,N_11576,N_9738);
or U13345 (N_13345,N_11795,N_9313);
and U13346 (N_13346,N_11492,N_10723);
nand U13347 (N_13347,N_10603,N_9176);
nand U13348 (N_13348,N_9873,N_9085);
nor U13349 (N_13349,N_11912,N_10193);
or U13350 (N_13350,N_10039,N_9796);
xor U13351 (N_13351,N_11864,N_10750);
nor U13352 (N_13352,N_9762,N_9346);
xor U13353 (N_13353,N_11208,N_9706);
and U13354 (N_13354,N_11847,N_10411);
nor U13355 (N_13355,N_9747,N_9526);
nand U13356 (N_13356,N_9966,N_10015);
or U13357 (N_13357,N_9092,N_11145);
nand U13358 (N_13358,N_9070,N_10131);
nand U13359 (N_13359,N_11021,N_9693);
nor U13360 (N_13360,N_10073,N_11386);
and U13361 (N_13361,N_9913,N_11474);
xor U13362 (N_13362,N_10094,N_9990);
nor U13363 (N_13363,N_9826,N_9270);
or U13364 (N_13364,N_10207,N_9131);
nand U13365 (N_13365,N_9236,N_10432);
or U13366 (N_13366,N_10858,N_9761);
nor U13367 (N_13367,N_9984,N_9062);
nand U13368 (N_13368,N_11307,N_11819);
or U13369 (N_13369,N_9465,N_9231);
and U13370 (N_13370,N_9556,N_11403);
and U13371 (N_13371,N_11930,N_10952);
nor U13372 (N_13372,N_9497,N_11450);
and U13373 (N_13373,N_9276,N_11632);
nor U13374 (N_13374,N_9952,N_11118);
nor U13375 (N_13375,N_9599,N_11883);
xnor U13376 (N_13376,N_11754,N_11866);
nand U13377 (N_13377,N_10593,N_11793);
or U13378 (N_13378,N_9733,N_9484);
nor U13379 (N_13379,N_10383,N_11159);
and U13380 (N_13380,N_9157,N_9852);
xnor U13381 (N_13381,N_10922,N_11517);
nor U13382 (N_13382,N_9023,N_11659);
nor U13383 (N_13383,N_11444,N_9268);
and U13384 (N_13384,N_10184,N_10439);
nor U13385 (N_13385,N_9274,N_11314);
nor U13386 (N_13386,N_10702,N_9104);
xnor U13387 (N_13387,N_10884,N_9958);
nor U13388 (N_13388,N_9536,N_11221);
xor U13389 (N_13389,N_10245,N_11476);
xnor U13390 (N_13390,N_11778,N_10125);
and U13391 (N_13391,N_11140,N_10862);
or U13392 (N_13392,N_9206,N_10937);
nor U13393 (N_13393,N_10418,N_9922);
nor U13394 (N_13394,N_10999,N_10205);
nor U13395 (N_13395,N_10074,N_11767);
xnor U13396 (N_13396,N_10931,N_9283);
xnor U13397 (N_13397,N_9851,N_10714);
or U13398 (N_13398,N_11548,N_9878);
or U13399 (N_13399,N_10260,N_9453);
nor U13400 (N_13400,N_11539,N_10625);
nand U13401 (N_13401,N_10901,N_9524);
nor U13402 (N_13402,N_11427,N_11837);
xor U13403 (N_13403,N_9174,N_10903);
or U13404 (N_13404,N_10949,N_10916);
nand U13405 (N_13405,N_11861,N_10407);
and U13406 (N_13406,N_11371,N_9128);
nor U13407 (N_13407,N_10778,N_9395);
or U13408 (N_13408,N_9165,N_11917);
and U13409 (N_13409,N_9224,N_10691);
or U13410 (N_13410,N_10572,N_11259);
or U13411 (N_13411,N_9053,N_11116);
and U13412 (N_13412,N_10048,N_11553);
or U13413 (N_13413,N_9251,N_11237);
and U13414 (N_13414,N_11820,N_9625);
xor U13415 (N_13415,N_9842,N_11203);
and U13416 (N_13416,N_11707,N_11800);
xnor U13417 (N_13417,N_11960,N_10425);
nor U13418 (N_13418,N_11027,N_10045);
nand U13419 (N_13419,N_11780,N_11544);
nor U13420 (N_13420,N_10239,N_11269);
xnor U13421 (N_13421,N_9838,N_11115);
nand U13422 (N_13422,N_9868,N_11459);
nor U13423 (N_13423,N_10277,N_11753);
xor U13424 (N_13424,N_11747,N_11775);
nor U13425 (N_13425,N_11547,N_11191);
nand U13426 (N_13426,N_11788,N_10118);
nor U13427 (N_13427,N_11012,N_9661);
and U13428 (N_13428,N_11302,N_9170);
xnor U13429 (N_13429,N_11823,N_11453);
or U13430 (N_13430,N_10057,N_9921);
nor U13431 (N_13431,N_11416,N_9345);
nor U13432 (N_13432,N_9759,N_9977);
and U13433 (N_13433,N_9169,N_11055);
or U13434 (N_13434,N_9633,N_10695);
xor U13435 (N_13435,N_10320,N_10571);
nand U13436 (N_13436,N_10994,N_10433);
nand U13437 (N_13437,N_10720,N_9024);
xor U13438 (N_13438,N_9755,N_10343);
and U13439 (N_13439,N_10218,N_9173);
or U13440 (N_13440,N_9760,N_11461);
or U13441 (N_13441,N_10807,N_10911);
and U13442 (N_13442,N_11686,N_9324);
xor U13443 (N_13443,N_9948,N_10591);
xor U13444 (N_13444,N_10103,N_10494);
and U13445 (N_13445,N_10208,N_11645);
and U13446 (N_13446,N_10833,N_9907);
or U13447 (N_13447,N_11110,N_10093);
or U13448 (N_13448,N_11737,N_11336);
nor U13449 (N_13449,N_11489,N_11384);
or U13450 (N_13450,N_11774,N_11617);
and U13451 (N_13451,N_10412,N_9279);
nand U13452 (N_13452,N_10292,N_10146);
nor U13453 (N_13453,N_9896,N_9096);
or U13454 (N_13454,N_9245,N_9699);
and U13455 (N_13455,N_9248,N_10424);
nor U13456 (N_13456,N_9278,N_9469);
or U13457 (N_13457,N_10083,N_9700);
nor U13458 (N_13458,N_11106,N_9354);
nand U13459 (N_13459,N_9932,N_10053);
xor U13460 (N_13460,N_10047,N_10470);
nor U13461 (N_13461,N_10230,N_10290);
and U13462 (N_13462,N_9322,N_11376);
nor U13463 (N_13463,N_10263,N_10366);
nor U13464 (N_13464,N_10462,N_11889);
xnor U13465 (N_13465,N_10564,N_11671);
nand U13466 (N_13466,N_10753,N_11469);
or U13467 (N_13467,N_10788,N_10244);
nor U13468 (N_13468,N_11057,N_9255);
xnor U13469 (N_13469,N_10119,N_11546);
nand U13470 (N_13470,N_9850,N_9018);
nand U13471 (N_13471,N_10287,N_11125);
xor U13472 (N_13472,N_9280,N_9615);
xnor U13473 (N_13473,N_10978,N_9452);
xnor U13474 (N_13474,N_11484,N_9953);
nor U13475 (N_13475,N_11235,N_9758);
or U13476 (N_13476,N_9876,N_9945);
and U13477 (N_13477,N_10760,N_10602);
nor U13478 (N_13478,N_11214,N_11891);
nor U13479 (N_13479,N_11749,N_9776);
xnor U13480 (N_13480,N_10367,N_10046);
xor U13481 (N_13481,N_10819,N_11424);
and U13482 (N_13482,N_11752,N_11194);
nand U13483 (N_13483,N_11653,N_11815);
or U13484 (N_13484,N_10346,N_10793);
or U13485 (N_13485,N_11648,N_11668);
or U13486 (N_13486,N_9017,N_9413);
nand U13487 (N_13487,N_10600,N_11759);
nor U13488 (N_13488,N_11486,N_11160);
and U13489 (N_13489,N_9378,N_11448);
nor U13490 (N_13490,N_10604,N_9962);
nand U13491 (N_13491,N_10838,N_10183);
nor U13492 (N_13492,N_9562,N_11325);
and U13493 (N_13493,N_11942,N_11105);
xor U13494 (N_13494,N_10638,N_9375);
xnor U13495 (N_13495,N_9303,N_10569);
nor U13496 (N_13496,N_9122,N_9073);
nor U13497 (N_13497,N_10742,N_9819);
nand U13498 (N_13498,N_11674,N_10071);
xor U13499 (N_13499,N_10241,N_9675);
nor U13500 (N_13500,N_9633,N_11112);
nand U13501 (N_13501,N_10795,N_9070);
xnor U13502 (N_13502,N_9624,N_9808);
and U13503 (N_13503,N_11531,N_11321);
xnor U13504 (N_13504,N_9951,N_9520);
or U13505 (N_13505,N_11352,N_9903);
and U13506 (N_13506,N_11015,N_11203);
and U13507 (N_13507,N_9117,N_10429);
nand U13508 (N_13508,N_11908,N_9091);
or U13509 (N_13509,N_11104,N_10182);
nor U13510 (N_13510,N_10587,N_11253);
and U13511 (N_13511,N_10386,N_11356);
or U13512 (N_13512,N_11662,N_11585);
xor U13513 (N_13513,N_11508,N_9982);
or U13514 (N_13514,N_9595,N_11318);
and U13515 (N_13515,N_10870,N_9010);
nand U13516 (N_13516,N_9043,N_9516);
and U13517 (N_13517,N_10338,N_11741);
nor U13518 (N_13518,N_11129,N_11287);
and U13519 (N_13519,N_11339,N_9133);
nand U13520 (N_13520,N_10873,N_9087);
xnor U13521 (N_13521,N_10112,N_11699);
xor U13522 (N_13522,N_10559,N_9903);
nor U13523 (N_13523,N_10246,N_10962);
xnor U13524 (N_13524,N_11993,N_11820);
nor U13525 (N_13525,N_11860,N_10982);
and U13526 (N_13526,N_11394,N_10626);
nand U13527 (N_13527,N_11254,N_11442);
nor U13528 (N_13528,N_9476,N_9342);
xor U13529 (N_13529,N_10867,N_11107);
xnor U13530 (N_13530,N_11355,N_11277);
xnor U13531 (N_13531,N_11819,N_10947);
and U13532 (N_13532,N_11123,N_10582);
nand U13533 (N_13533,N_11713,N_9397);
xnor U13534 (N_13534,N_10276,N_9719);
or U13535 (N_13535,N_9844,N_9945);
xnor U13536 (N_13536,N_11160,N_9652);
nor U13537 (N_13537,N_10000,N_9736);
or U13538 (N_13538,N_11020,N_10466);
nand U13539 (N_13539,N_10609,N_11423);
or U13540 (N_13540,N_9242,N_11144);
and U13541 (N_13541,N_10940,N_9985);
xnor U13542 (N_13542,N_9474,N_10628);
and U13543 (N_13543,N_9301,N_11493);
nand U13544 (N_13544,N_10658,N_10934);
xor U13545 (N_13545,N_10770,N_10466);
or U13546 (N_13546,N_10438,N_9987);
and U13547 (N_13547,N_11528,N_10480);
nor U13548 (N_13548,N_11931,N_9952);
and U13549 (N_13549,N_10129,N_9109);
and U13550 (N_13550,N_11008,N_10186);
nand U13551 (N_13551,N_9450,N_10250);
nand U13552 (N_13552,N_9144,N_10038);
and U13553 (N_13553,N_10770,N_10293);
or U13554 (N_13554,N_11325,N_9671);
or U13555 (N_13555,N_9094,N_9146);
or U13556 (N_13556,N_11090,N_9971);
nand U13557 (N_13557,N_9989,N_11031);
or U13558 (N_13558,N_11586,N_11458);
nand U13559 (N_13559,N_11593,N_9390);
xor U13560 (N_13560,N_11028,N_11838);
or U13561 (N_13561,N_10029,N_11452);
nor U13562 (N_13562,N_10674,N_9431);
and U13563 (N_13563,N_11573,N_10735);
xor U13564 (N_13564,N_10694,N_10853);
and U13565 (N_13565,N_9304,N_11763);
nor U13566 (N_13566,N_9971,N_10143);
or U13567 (N_13567,N_11218,N_10115);
or U13568 (N_13568,N_9701,N_9562);
nand U13569 (N_13569,N_10565,N_9149);
nor U13570 (N_13570,N_10283,N_10082);
and U13571 (N_13571,N_10452,N_9850);
nand U13572 (N_13572,N_11536,N_9089);
nand U13573 (N_13573,N_10645,N_11828);
nand U13574 (N_13574,N_9616,N_10293);
xnor U13575 (N_13575,N_10151,N_11941);
and U13576 (N_13576,N_10338,N_10751);
and U13577 (N_13577,N_11641,N_9625);
nor U13578 (N_13578,N_9475,N_9199);
nor U13579 (N_13579,N_10686,N_9601);
and U13580 (N_13580,N_10469,N_10601);
or U13581 (N_13581,N_9313,N_10068);
and U13582 (N_13582,N_9382,N_9733);
and U13583 (N_13583,N_9792,N_11536);
or U13584 (N_13584,N_11401,N_11490);
and U13585 (N_13585,N_9651,N_9894);
xor U13586 (N_13586,N_10516,N_10424);
nor U13587 (N_13587,N_10800,N_10802);
or U13588 (N_13588,N_10629,N_9025);
or U13589 (N_13589,N_9950,N_9716);
nor U13590 (N_13590,N_10767,N_9451);
xor U13591 (N_13591,N_11394,N_11832);
or U13592 (N_13592,N_11320,N_10585);
or U13593 (N_13593,N_11865,N_10593);
and U13594 (N_13594,N_10795,N_11178);
xnor U13595 (N_13595,N_10699,N_9374);
nor U13596 (N_13596,N_9192,N_11682);
or U13597 (N_13597,N_11986,N_11809);
nand U13598 (N_13598,N_11481,N_11100);
or U13599 (N_13599,N_11930,N_10660);
and U13600 (N_13600,N_9542,N_11597);
and U13601 (N_13601,N_9543,N_11805);
nor U13602 (N_13602,N_10555,N_10163);
nor U13603 (N_13603,N_10185,N_9306);
nand U13604 (N_13604,N_11599,N_11149);
xnor U13605 (N_13605,N_9934,N_10439);
and U13606 (N_13606,N_9059,N_9425);
xor U13607 (N_13607,N_11011,N_9430);
nor U13608 (N_13608,N_9273,N_9368);
xnor U13609 (N_13609,N_9560,N_10586);
nand U13610 (N_13610,N_9197,N_10786);
xnor U13611 (N_13611,N_11161,N_10502);
nand U13612 (N_13612,N_11602,N_10792);
nand U13613 (N_13613,N_11360,N_11187);
xnor U13614 (N_13614,N_9471,N_9043);
xor U13615 (N_13615,N_11634,N_10195);
nor U13616 (N_13616,N_9301,N_11465);
nor U13617 (N_13617,N_10140,N_10502);
nand U13618 (N_13618,N_10492,N_10372);
or U13619 (N_13619,N_11555,N_10441);
nor U13620 (N_13620,N_10234,N_9800);
and U13621 (N_13621,N_9266,N_11546);
nor U13622 (N_13622,N_10433,N_10722);
or U13623 (N_13623,N_11360,N_11357);
and U13624 (N_13624,N_11282,N_11300);
xor U13625 (N_13625,N_9781,N_10037);
xnor U13626 (N_13626,N_11591,N_11601);
xor U13627 (N_13627,N_10269,N_10184);
and U13628 (N_13628,N_9506,N_11565);
nand U13629 (N_13629,N_11066,N_11844);
nand U13630 (N_13630,N_10612,N_11113);
or U13631 (N_13631,N_10661,N_10084);
and U13632 (N_13632,N_11656,N_11579);
xnor U13633 (N_13633,N_9918,N_11869);
nor U13634 (N_13634,N_11315,N_10604);
xor U13635 (N_13635,N_9033,N_10477);
and U13636 (N_13636,N_11252,N_9824);
or U13637 (N_13637,N_10325,N_11438);
xnor U13638 (N_13638,N_9292,N_9846);
nor U13639 (N_13639,N_11040,N_10002);
nand U13640 (N_13640,N_11419,N_11306);
xor U13641 (N_13641,N_9374,N_9598);
and U13642 (N_13642,N_9899,N_9736);
nor U13643 (N_13643,N_11405,N_11286);
or U13644 (N_13644,N_10879,N_11498);
nor U13645 (N_13645,N_9820,N_11104);
and U13646 (N_13646,N_10723,N_10061);
nand U13647 (N_13647,N_11175,N_9713);
and U13648 (N_13648,N_11729,N_11057);
nor U13649 (N_13649,N_10138,N_11039);
xnor U13650 (N_13650,N_11721,N_11537);
or U13651 (N_13651,N_10214,N_11829);
nand U13652 (N_13652,N_9612,N_10437);
or U13653 (N_13653,N_11531,N_10681);
nor U13654 (N_13654,N_10426,N_9646);
nand U13655 (N_13655,N_9849,N_10560);
nor U13656 (N_13656,N_11628,N_11242);
nor U13657 (N_13657,N_11411,N_11443);
or U13658 (N_13658,N_10019,N_10582);
nand U13659 (N_13659,N_10686,N_9793);
or U13660 (N_13660,N_9114,N_9750);
and U13661 (N_13661,N_10450,N_9547);
or U13662 (N_13662,N_11578,N_9480);
nor U13663 (N_13663,N_10768,N_11190);
nor U13664 (N_13664,N_11751,N_10038);
xor U13665 (N_13665,N_9522,N_9871);
nor U13666 (N_13666,N_11832,N_11850);
xnor U13667 (N_13667,N_10531,N_10372);
xor U13668 (N_13668,N_11526,N_9836);
nor U13669 (N_13669,N_11330,N_10625);
and U13670 (N_13670,N_10455,N_11920);
nor U13671 (N_13671,N_11613,N_9110);
nor U13672 (N_13672,N_10250,N_11801);
xnor U13673 (N_13673,N_9491,N_11906);
nand U13674 (N_13674,N_11098,N_10016);
xor U13675 (N_13675,N_10784,N_9491);
xnor U13676 (N_13676,N_9929,N_9021);
or U13677 (N_13677,N_11715,N_9877);
xnor U13678 (N_13678,N_10350,N_9468);
nand U13679 (N_13679,N_9585,N_10691);
nand U13680 (N_13680,N_10482,N_11143);
nor U13681 (N_13681,N_10103,N_9744);
and U13682 (N_13682,N_11132,N_9859);
nand U13683 (N_13683,N_9296,N_11421);
xor U13684 (N_13684,N_11459,N_9239);
nor U13685 (N_13685,N_9714,N_11965);
or U13686 (N_13686,N_9452,N_9779);
and U13687 (N_13687,N_9297,N_9676);
or U13688 (N_13688,N_9683,N_10328);
or U13689 (N_13689,N_10595,N_9680);
xor U13690 (N_13690,N_11285,N_11474);
nand U13691 (N_13691,N_11657,N_11816);
xor U13692 (N_13692,N_11193,N_11404);
nand U13693 (N_13693,N_9786,N_11003);
nand U13694 (N_13694,N_9793,N_9544);
nor U13695 (N_13695,N_10656,N_11521);
xor U13696 (N_13696,N_11405,N_11610);
or U13697 (N_13697,N_9312,N_11587);
xnor U13698 (N_13698,N_11638,N_10959);
nor U13699 (N_13699,N_9768,N_11808);
nand U13700 (N_13700,N_10775,N_11472);
nor U13701 (N_13701,N_11980,N_9603);
and U13702 (N_13702,N_11300,N_11243);
and U13703 (N_13703,N_10395,N_10920);
xnor U13704 (N_13704,N_9342,N_9694);
nor U13705 (N_13705,N_9353,N_9097);
nand U13706 (N_13706,N_9242,N_10520);
xnor U13707 (N_13707,N_10108,N_9420);
or U13708 (N_13708,N_10414,N_10685);
nor U13709 (N_13709,N_9642,N_9927);
xnor U13710 (N_13710,N_10523,N_11307);
xnor U13711 (N_13711,N_9423,N_10273);
or U13712 (N_13712,N_11693,N_11444);
or U13713 (N_13713,N_10431,N_11155);
or U13714 (N_13714,N_9936,N_11929);
nand U13715 (N_13715,N_9988,N_11250);
or U13716 (N_13716,N_9898,N_9985);
or U13717 (N_13717,N_9595,N_10199);
nor U13718 (N_13718,N_10286,N_11767);
nor U13719 (N_13719,N_11341,N_9992);
or U13720 (N_13720,N_11667,N_10548);
nor U13721 (N_13721,N_9395,N_9345);
nor U13722 (N_13722,N_10224,N_10192);
or U13723 (N_13723,N_9191,N_11251);
nand U13724 (N_13724,N_9576,N_11367);
nand U13725 (N_13725,N_9199,N_11624);
and U13726 (N_13726,N_11632,N_10750);
or U13727 (N_13727,N_9698,N_10884);
or U13728 (N_13728,N_9241,N_10128);
xor U13729 (N_13729,N_9309,N_11192);
nor U13730 (N_13730,N_11388,N_10265);
nand U13731 (N_13731,N_10792,N_9928);
and U13732 (N_13732,N_11602,N_9600);
xor U13733 (N_13733,N_9723,N_11503);
xnor U13734 (N_13734,N_11224,N_9211);
nor U13735 (N_13735,N_9139,N_10945);
and U13736 (N_13736,N_10471,N_9075);
or U13737 (N_13737,N_10578,N_9213);
or U13738 (N_13738,N_11309,N_9077);
nor U13739 (N_13739,N_11357,N_11326);
or U13740 (N_13740,N_10906,N_9906);
nor U13741 (N_13741,N_9669,N_11560);
and U13742 (N_13742,N_9103,N_9526);
nand U13743 (N_13743,N_11489,N_10601);
or U13744 (N_13744,N_9747,N_11661);
and U13745 (N_13745,N_11115,N_10281);
nand U13746 (N_13746,N_9177,N_10185);
nor U13747 (N_13747,N_10449,N_10158);
nor U13748 (N_13748,N_10599,N_10881);
and U13749 (N_13749,N_9676,N_11831);
nor U13750 (N_13750,N_11778,N_10442);
and U13751 (N_13751,N_9870,N_11515);
nand U13752 (N_13752,N_10121,N_9436);
and U13753 (N_13753,N_11418,N_10744);
or U13754 (N_13754,N_9921,N_11344);
or U13755 (N_13755,N_11109,N_9025);
xor U13756 (N_13756,N_10598,N_9875);
xnor U13757 (N_13757,N_11692,N_9324);
nand U13758 (N_13758,N_11624,N_9982);
and U13759 (N_13759,N_9244,N_11625);
nand U13760 (N_13760,N_9707,N_10726);
nor U13761 (N_13761,N_10365,N_10989);
and U13762 (N_13762,N_11559,N_10887);
and U13763 (N_13763,N_10664,N_11260);
xor U13764 (N_13764,N_11779,N_10823);
and U13765 (N_13765,N_10918,N_11725);
xnor U13766 (N_13766,N_9637,N_11676);
xnor U13767 (N_13767,N_11823,N_10625);
and U13768 (N_13768,N_11035,N_9714);
nand U13769 (N_13769,N_11904,N_9684);
nand U13770 (N_13770,N_9031,N_9279);
nor U13771 (N_13771,N_10235,N_9206);
nor U13772 (N_13772,N_11241,N_11955);
and U13773 (N_13773,N_9775,N_10395);
xor U13774 (N_13774,N_11850,N_10141);
nor U13775 (N_13775,N_11209,N_10600);
or U13776 (N_13776,N_10591,N_11945);
nand U13777 (N_13777,N_10229,N_11974);
nor U13778 (N_13778,N_10311,N_9062);
and U13779 (N_13779,N_9701,N_11324);
nor U13780 (N_13780,N_10705,N_11948);
xnor U13781 (N_13781,N_11088,N_9522);
and U13782 (N_13782,N_10057,N_11059);
or U13783 (N_13783,N_9748,N_10700);
nand U13784 (N_13784,N_9381,N_11603);
and U13785 (N_13785,N_9037,N_10811);
nand U13786 (N_13786,N_11895,N_10903);
nand U13787 (N_13787,N_9889,N_11047);
nand U13788 (N_13788,N_11823,N_11656);
and U13789 (N_13789,N_9658,N_10815);
or U13790 (N_13790,N_9494,N_11129);
nor U13791 (N_13791,N_11542,N_9727);
xnor U13792 (N_13792,N_10330,N_9577);
or U13793 (N_13793,N_9319,N_11592);
or U13794 (N_13794,N_10385,N_11953);
nand U13795 (N_13795,N_9069,N_9786);
and U13796 (N_13796,N_9383,N_11916);
xnor U13797 (N_13797,N_9272,N_10132);
or U13798 (N_13798,N_11446,N_11666);
nand U13799 (N_13799,N_10660,N_11323);
and U13800 (N_13800,N_11728,N_11762);
or U13801 (N_13801,N_11937,N_9091);
xnor U13802 (N_13802,N_10446,N_9604);
xor U13803 (N_13803,N_10050,N_10963);
or U13804 (N_13804,N_9021,N_11828);
or U13805 (N_13805,N_9756,N_9227);
and U13806 (N_13806,N_11012,N_10815);
or U13807 (N_13807,N_9523,N_10449);
and U13808 (N_13808,N_11997,N_11409);
and U13809 (N_13809,N_9552,N_11119);
or U13810 (N_13810,N_10047,N_9711);
xnor U13811 (N_13811,N_10765,N_10064);
and U13812 (N_13812,N_9397,N_10900);
nor U13813 (N_13813,N_11173,N_9930);
and U13814 (N_13814,N_9301,N_11229);
nand U13815 (N_13815,N_11406,N_10417);
xor U13816 (N_13816,N_9694,N_9257);
xor U13817 (N_13817,N_9096,N_10790);
xor U13818 (N_13818,N_11961,N_9331);
nand U13819 (N_13819,N_10105,N_11401);
and U13820 (N_13820,N_9491,N_11229);
nand U13821 (N_13821,N_11230,N_9310);
or U13822 (N_13822,N_9047,N_11731);
nor U13823 (N_13823,N_9634,N_11838);
nand U13824 (N_13824,N_11285,N_10684);
or U13825 (N_13825,N_11352,N_9172);
nor U13826 (N_13826,N_9890,N_11078);
and U13827 (N_13827,N_10074,N_10478);
and U13828 (N_13828,N_11152,N_11574);
nor U13829 (N_13829,N_10276,N_11378);
nor U13830 (N_13830,N_9204,N_9605);
xor U13831 (N_13831,N_9360,N_11618);
xnor U13832 (N_13832,N_9715,N_10323);
nand U13833 (N_13833,N_9742,N_10095);
and U13834 (N_13834,N_9765,N_10334);
nor U13835 (N_13835,N_10675,N_9382);
or U13836 (N_13836,N_11316,N_11277);
nor U13837 (N_13837,N_9414,N_9465);
nand U13838 (N_13838,N_11344,N_9729);
nor U13839 (N_13839,N_10318,N_11073);
xnor U13840 (N_13840,N_9641,N_11665);
nand U13841 (N_13841,N_10420,N_11546);
and U13842 (N_13842,N_10071,N_11788);
and U13843 (N_13843,N_10785,N_11689);
or U13844 (N_13844,N_9075,N_11818);
nor U13845 (N_13845,N_11694,N_9913);
nor U13846 (N_13846,N_10392,N_9521);
or U13847 (N_13847,N_9757,N_10466);
xnor U13848 (N_13848,N_9637,N_9639);
and U13849 (N_13849,N_9001,N_10572);
xnor U13850 (N_13850,N_11431,N_9379);
and U13851 (N_13851,N_9116,N_11106);
and U13852 (N_13852,N_9407,N_11883);
nand U13853 (N_13853,N_10609,N_9211);
nor U13854 (N_13854,N_10708,N_10047);
nand U13855 (N_13855,N_11027,N_10124);
and U13856 (N_13856,N_11918,N_9069);
and U13857 (N_13857,N_10966,N_10582);
or U13858 (N_13858,N_11744,N_10792);
xor U13859 (N_13859,N_9479,N_10882);
xnor U13860 (N_13860,N_9101,N_10525);
or U13861 (N_13861,N_11562,N_10404);
xnor U13862 (N_13862,N_11089,N_9170);
nor U13863 (N_13863,N_10176,N_10712);
and U13864 (N_13864,N_10289,N_10792);
nand U13865 (N_13865,N_9871,N_9551);
or U13866 (N_13866,N_10480,N_9582);
or U13867 (N_13867,N_9314,N_10984);
and U13868 (N_13868,N_9778,N_9617);
and U13869 (N_13869,N_11390,N_11926);
xnor U13870 (N_13870,N_10685,N_9096);
or U13871 (N_13871,N_10041,N_10759);
nand U13872 (N_13872,N_10122,N_10615);
or U13873 (N_13873,N_10005,N_10380);
nor U13874 (N_13874,N_11291,N_11485);
nor U13875 (N_13875,N_11312,N_11647);
or U13876 (N_13876,N_11955,N_11002);
nand U13877 (N_13877,N_10848,N_9680);
or U13878 (N_13878,N_9847,N_11324);
or U13879 (N_13879,N_9940,N_11379);
xnor U13880 (N_13880,N_11962,N_10948);
nor U13881 (N_13881,N_11179,N_11281);
nor U13882 (N_13882,N_9579,N_11669);
nor U13883 (N_13883,N_11475,N_10150);
xnor U13884 (N_13884,N_11265,N_9023);
and U13885 (N_13885,N_11156,N_11537);
xor U13886 (N_13886,N_11069,N_10816);
nor U13887 (N_13887,N_11379,N_9629);
or U13888 (N_13888,N_9250,N_9512);
and U13889 (N_13889,N_9902,N_9629);
or U13890 (N_13890,N_10264,N_10856);
nor U13891 (N_13891,N_9872,N_9320);
nand U13892 (N_13892,N_9084,N_11019);
nor U13893 (N_13893,N_9552,N_11293);
and U13894 (N_13894,N_9517,N_10203);
and U13895 (N_13895,N_11836,N_9840);
nand U13896 (N_13896,N_11890,N_10729);
and U13897 (N_13897,N_9362,N_10340);
and U13898 (N_13898,N_9046,N_11759);
nor U13899 (N_13899,N_10111,N_9583);
xor U13900 (N_13900,N_9022,N_11468);
or U13901 (N_13901,N_9127,N_11437);
nand U13902 (N_13902,N_10588,N_9703);
nand U13903 (N_13903,N_10575,N_10685);
nor U13904 (N_13904,N_10652,N_11771);
or U13905 (N_13905,N_10312,N_11390);
or U13906 (N_13906,N_10595,N_9526);
nand U13907 (N_13907,N_11671,N_10645);
nor U13908 (N_13908,N_10776,N_11310);
xor U13909 (N_13909,N_9657,N_11398);
and U13910 (N_13910,N_9131,N_10783);
or U13911 (N_13911,N_11727,N_9143);
or U13912 (N_13912,N_9864,N_11798);
xnor U13913 (N_13913,N_10862,N_10642);
or U13914 (N_13914,N_9883,N_9573);
xor U13915 (N_13915,N_10270,N_11854);
xnor U13916 (N_13916,N_11938,N_9109);
nand U13917 (N_13917,N_10858,N_11199);
or U13918 (N_13918,N_10118,N_10863);
xor U13919 (N_13919,N_10478,N_9467);
nor U13920 (N_13920,N_9916,N_10161);
or U13921 (N_13921,N_9568,N_10585);
xnor U13922 (N_13922,N_11923,N_9868);
and U13923 (N_13923,N_9763,N_10956);
nand U13924 (N_13924,N_10557,N_11709);
nand U13925 (N_13925,N_11030,N_10828);
and U13926 (N_13926,N_11235,N_9391);
xor U13927 (N_13927,N_11346,N_9982);
nand U13928 (N_13928,N_11300,N_9789);
xnor U13929 (N_13929,N_10775,N_9090);
or U13930 (N_13930,N_11895,N_9984);
nor U13931 (N_13931,N_9139,N_11265);
nand U13932 (N_13932,N_11395,N_10634);
or U13933 (N_13933,N_11243,N_10621);
and U13934 (N_13934,N_10487,N_11794);
nand U13935 (N_13935,N_11830,N_10843);
xnor U13936 (N_13936,N_11293,N_10999);
xnor U13937 (N_13937,N_10223,N_9793);
nor U13938 (N_13938,N_9604,N_10452);
nor U13939 (N_13939,N_11014,N_11741);
nor U13940 (N_13940,N_11419,N_10803);
or U13941 (N_13941,N_10089,N_11931);
nand U13942 (N_13942,N_10580,N_9145);
xor U13943 (N_13943,N_9766,N_9978);
xnor U13944 (N_13944,N_11639,N_10027);
and U13945 (N_13945,N_10154,N_10720);
nor U13946 (N_13946,N_9138,N_9763);
or U13947 (N_13947,N_10190,N_10841);
xor U13948 (N_13948,N_9487,N_9902);
nor U13949 (N_13949,N_10963,N_11375);
or U13950 (N_13950,N_11396,N_10207);
xor U13951 (N_13951,N_9276,N_11841);
and U13952 (N_13952,N_11137,N_11868);
and U13953 (N_13953,N_9515,N_10298);
nor U13954 (N_13954,N_10833,N_10955);
and U13955 (N_13955,N_11807,N_11351);
or U13956 (N_13956,N_9745,N_9322);
nor U13957 (N_13957,N_10530,N_11846);
nor U13958 (N_13958,N_9973,N_11198);
or U13959 (N_13959,N_9601,N_10227);
or U13960 (N_13960,N_11667,N_9594);
nor U13961 (N_13961,N_9402,N_9082);
or U13962 (N_13962,N_9127,N_11227);
or U13963 (N_13963,N_11594,N_11244);
nor U13964 (N_13964,N_11365,N_10180);
nand U13965 (N_13965,N_9982,N_10003);
or U13966 (N_13966,N_10405,N_11419);
xor U13967 (N_13967,N_11624,N_11856);
or U13968 (N_13968,N_10803,N_11572);
nor U13969 (N_13969,N_10878,N_10793);
nor U13970 (N_13970,N_9037,N_9646);
nand U13971 (N_13971,N_11502,N_11778);
and U13972 (N_13972,N_10577,N_10037);
nand U13973 (N_13973,N_10416,N_11761);
or U13974 (N_13974,N_9205,N_10871);
nand U13975 (N_13975,N_11163,N_10993);
nand U13976 (N_13976,N_9355,N_9323);
xor U13977 (N_13977,N_10597,N_11771);
nand U13978 (N_13978,N_9377,N_10013);
and U13979 (N_13979,N_11488,N_11764);
nand U13980 (N_13980,N_9719,N_9649);
nor U13981 (N_13981,N_10363,N_10346);
or U13982 (N_13982,N_9151,N_9720);
or U13983 (N_13983,N_9143,N_10361);
nand U13984 (N_13984,N_9983,N_10975);
and U13985 (N_13985,N_10634,N_10533);
and U13986 (N_13986,N_9007,N_9371);
or U13987 (N_13987,N_9151,N_10689);
and U13988 (N_13988,N_9240,N_9308);
xor U13989 (N_13989,N_10688,N_11278);
and U13990 (N_13990,N_11513,N_10213);
and U13991 (N_13991,N_9825,N_9210);
and U13992 (N_13992,N_11156,N_10258);
xnor U13993 (N_13993,N_10652,N_10482);
or U13994 (N_13994,N_11231,N_9885);
and U13995 (N_13995,N_10655,N_9950);
xor U13996 (N_13996,N_11852,N_11526);
nor U13997 (N_13997,N_10204,N_11920);
nor U13998 (N_13998,N_10043,N_10123);
and U13999 (N_13999,N_11591,N_9275);
nand U14000 (N_14000,N_11347,N_10472);
and U14001 (N_14001,N_10156,N_9060);
or U14002 (N_14002,N_10060,N_10918);
nand U14003 (N_14003,N_9501,N_9254);
nor U14004 (N_14004,N_11391,N_11677);
or U14005 (N_14005,N_10523,N_11771);
nand U14006 (N_14006,N_11013,N_11494);
nand U14007 (N_14007,N_11430,N_11934);
nor U14008 (N_14008,N_10367,N_10990);
nand U14009 (N_14009,N_9899,N_9940);
nand U14010 (N_14010,N_10223,N_9564);
nor U14011 (N_14011,N_11754,N_11078);
or U14012 (N_14012,N_9218,N_9295);
or U14013 (N_14013,N_11416,N_10565);
xnor U14014 (N_14014,N_9052,N_11672);
and U14015 (N_14015,N_10348,N_11209);
and U14016 (N_14016,N_11471,N_10355);
nor U14017 (N_14017,N_11747,N_10045);
nor U14018 (N_14018,N_10767,N_11807);
nor U14019 (N_14019,N_11721,N_9535);
nor U14020 (N_14020,N_9412,N_11666);
or U14021 (N_14021,N_10633,N_9189);
nor U14022 (N_14022,N_11480,N_10558);
and U14023 (N_14023,N_11599,N_10760);
xor U14024 (N_14024,N_9164,N_9533);
nand U14025 (N_14025,N_11428,N_11940);
and U14026 (N_14026,N_9007,N_9257);
xor U14027 (N_14027,N_10483,N_10566);
or U14028 (N_14028,N_9525,N_11523);
nand U14029 (N_14029,N_11717,N_10594);
nor U14030 (N_14030,N_11284,N_11705);
or U14031 (N_14031,N_9552,N_10788);
or U14032 (N_14032,N_9656,N_9447);
nand U14033 (N_14033,N_10449,N_10819);
xor U14034 (N_14034,N_10596,N_11668);
and U14035 (N_14035,N_11762,N_9678);
nand U14036 (N_14036,N_11693,N_10597);
nor U14037 (N_14037,N_10416,N_11817);
nand U14038 (N_14038,N_10580,N_10325);
xnor U14039 (N_14039,N_9361,N_9151);
xor U14040 (N_14040,N_11980,N_11280);
xnor U14041 (N_14041,N_10758,N_10695);
or U14042 (N_14042,N_9049,N_9541);
nand U14043 (N_14043,N_9455,N_9123);
xor U14044 (N_14044,N_10772,N_10427);
nand U14045 (N_14045,N_10686,N_10378);
nand U14046 (N_14046,N_10566,N_11286);
xor U14047 (N_14047,N_11641,N_10902);
and U14048 (N_14048,N_11244,N_11750);
nor U14049 (N_14049,N_11401,N_9053);
xnor U14050 (N_14050,N_9385,N_9892);
nor U14051 (N_14051,N_10914,N_11897);
nand U14052 (N_14052,N_9677,N_10866);
xor U14053 (N_14053,N_9120,N_11663);
and U14054 (N_14054,N_11628,N_11435);
nand U14055 (N_14055,N_10848,N_11888);
and U14056 (N_14056,N_11536,N_9331);
xor U14057 (N_14057,N_10768,N_11526);
xor U14058 (N_14058,N_10139,N_9072);
and U14059 (N_14059,N_9074,N_9596);
nand U14060 (N_14060,N_10506,N_11241);
xnor U14061 (N_14061,N_9929,N_10072);
or U14062 (N_14062,N_9060,N_10782);
nor U14063 (N_14063,N_9568,N_10637);
and U14064 (N_14064,N_10152,N_11480);
nor U14065 (N_14065,N_10695,N_10929);
nand U14066 (N_14066,N_9048,N_11310);
and U14067 (N_14067,N_11950,N_9150);
or U14068 (N_14068,N_9350,N_9466);
nor U14069 (N_14069,N_10151,N_9277);
nand U14070 (N_14070,N_10931,N_9067);
or U14071 (N_14071,N_11736,N_11003);
or U14072 (N_14072,N_11929,N_9488);
and U14073 (N_14073,N_9679,N_9879);
and U14074 (N_14074,N_9178,N_11387);
and U14075 (N_14075,N_11158,N_11853);
and U14076 (N_14076,N_9541,N_9223);
and U14077 (N_14077,N_9009,N_11175);
and U14078 (N_14078,N_9207,N_10753);
nand U14079 (N_14079,N_10248,N_9548);
nor U14080 (N_14080,N_11593,N_10299);
nand U14081 (N_14081,N_11807,N_10122);
or U14082 (N_14082,N_9372,N_10158);
or U14083 (N_14083,N_9060,N_11217);
and U14084 (N_14084,N_11945,N_10351);
nand U14085 (N_14085,N_10001,N_10283);
and U14086 (N_14086,N_11268,N_11668);
xor U14087 (N_14087,N_9198,N_11571);
nand U14088 (N_14088,N_10847,N_11435);
and U14089 (N_14089,N_11409,N_11411);
nor U14090 (N_14090,N_10904,N_10763);
and U14091 (N_14091,N_10623,N_9302);
nand U14092 (N_14092,N_9489,N_11334);
xor U14093 (N_14093,N_9055,N_11532);
and U14094 (N_14094,N_11866,N_10238);
nand U14095 (N_14095,N_10082,N_9562);
and U14096 (N_14096,N_10891,N_9103);
nor U14097 (N_14097,N_10106,N_11673);
nand U14098 (N_14098,N_11617,N_10456);
nand U14099 (N_14099,N_11102,N_11649);
nand U14100 (N_14100,N_11585,N_10980);
or U14101 (N_14101,N_9821,N_11928);
xor U14102 (N_14102,N_11425,N_10925);
xnor U14103 (N_14103,N_11017,N_10004);
or U14104 (N_14104,N_10055,N_11060);
or U14105 (N_14105,N_9326,N_10516);
nand U14106 (N_14106,N_9043,N_10379);
nand U14107 (N_14107,N_9265,N_10981);
and U14108 (N_14108,N_11800,N_11431);
and U14109 (N_14109,N_10682,N_11131);
or U14110 (N_14110,N_11006,N_11659);
and U14111 (N_14111,N_11929,N_9687);
nand U14112 (N_14112,N_10687,N_11719);
nand U14113 (N_14113,N_11401,N_10912);
or U14114 (N_14114,N_11553,N_10440);
and U14115 (N_14115,N_10964,N_9419);
and U14116 (N_14116,N_11086,N_9223);
xnor U14117 (N_14117,N_11154,N_11316);
or U14118 (N_14118,N_10858,N_10646);
or U14119 (N_14119,N_9805,N_11852);
or U14120 (N_14120,N_9313,N_10317);
and U14121 (N_14121,N_11329,N_9344);
nand U14122 (N_14122,N_9657,N_9619);
nand U14123 (N_14123,N_9909,N_10096);
nor U14124 (N_14124,N_9330,N_9146);
and U14125 (N_14125,N_10980,N_10852);
and U14126 (N_14126,N_9317,N_9727);
nor U14127 (N_14127,N_9984,N_10880);
nand U14128 (N_14128,N_10816,N_9545);
and U14129 (N_14129,N_11970,N_10058);
xor U14130 (N_14130,N_11176,N_9329);
xnor U14131 (N_14131,N_10184,N_10151);
and U14132 (N_14132,N_11837,N_10120);
or U14133 (N_14133,N_9999,N_11442);
nor U14134 (N_14134,N_10018,N_10622);
nand U14135 (N_14135,N_9661,N_10271);
nand U14136 (N_14136,N_11001,N_9072);
nor U14137 (N_14137,N_10238,N_10188);
nand U14138 (N_14138,N_10201,N_9796);
nand U14139 (N_14139,N_9087,N_11008);
nor U14140 (N_14140,N_9245,N_9189);
nor U14141 (N_14141,N_10967,N_9529);
nor U14142 (N_14142,N_9358,N_11922);
xor U14143 (N_14143,N_10538,N_9702);
nor U14144 (N_14144,N_9754,N_9495);
nand U14145 (N_14145,N_10551,N_9729);
xnor U14146 (N_14146,N_9060,N_9702);
xor U14147 (N_14147,N_9974,N_9306);
and U14148 (N_14148,N_9398,N_9487);
xor U14149 (N_14149,N_11674,N_10588);
and U14150 (N_14150,N_11544,N_11413);
nand U14151 (N_14151,N_9648,N_9306);
nand U14152 (N_14152,N_9935,N_11807);
nor U14153 (N_14153,N_11730,N_10630);
xor U14154 (N_14154,N_10419,N_11373);
or U14155 (N_14155,N_11590,N_10569);
nand U14156 (N_14156,N_10734,N_9360);
nor U14157 (N_14157,N_11756,N_11265);
or U14158 (N_14158,N_9893,N_11264);
or U14159 (N_14159,N_9546,N_11177);
xor U14160 (N_14160,N_9729,N_11124);
and U14161 (N_14161,N_10522,N_11560);
and U14162 (N_14162,N_10790,N_11957);
and U14163 (N_14163,N_11189,N_9701);
or U14164 (N_14164,N_9710,N_11137);
xor U14165 (N_14165,N_11431,N_10360);
nor U14166 (N_14166,N_10348,N_10469);
xnor U14167 (N_14167,N_10586,N_10463);
xnor U14168 (N_14168,N_9455,N_9524);
and U14169 (N_14169,N_10593,N_11102);
nand U14170 (N_14170,N_10465,N_10195);
nand U14171 (N_14171,N_10026,N_9366);
xnor U14172 (N_14172,N_10780,N_11006);
nor U14173 (N_14173,N_10498,N_9086);
or U14174 (N_14174,N_11365,N_9379);
nand U14175 (N_14175,N_11697,N_9317);
xor U14176 (N_14176,N_9392,N_9894);
and U14177 (N_14177,N_9238,N_9431);
and U14178 (N_14178,N_10340,N_9902);
and U14179 (N_14179,N_10073,N_10636);
nand U14180 (N_14180,N_9618,N_11781);
xor U14181 (N_14181,N_11610,N_10333);
nor U14182 (N_14182,N_9680,N_11246);
nand U14183 (N_14183,N_11720,N_11491);
xor U14184 (N_14184,N_10601,N_10201);
or U14185 (N_14185,N_9623,N_11770);
nor U14186 (N_14186,N_9746,N_9780);
nor U14187 (N_14187,N_10770,N_11021);
nand U14188 (N_14188,N_11382,N_9202);
xnor U14189 (N_14189,N_9154,N_10340);
and U14190 (N_14190,N_11158,N_10791);
or U14191 (N_14191,N_11878,N_10075);
and U14192 (N_14192,N_9997,N_10690);
nor U14193 (N_14193,N_11741,N_9794);
or U14194 (N_14194,N_10774,N_9257);
nor U14195 (N_14195,N_9732,N_11553);
or U14196 (N_14196,N_10233,N_10247);
xnor U14197 (N_14197,N_9606,N_11512);
or U14198 (N_14198,N_10922,N_10900);
nand U14199 (N_14199,N_9238,N_11287);
and U14200 (N_14200,N_11408,N_9748);
and U14201 (N_14201,N_10628,N_10849);
or U14202 (N_14202,N_9952,N_11609);
and U14203 (N_14203,N_9392,N_11964);
or U14204 (N_14204,N_9189,N_10826);
xor U14205 (N_14205,N_10490,N_9341);
or U14206 (N_14206,N_9813,N_9001);
nand U14207 (N_14207,N_11715,N_11751);
nand U14208 (N_14208,N_10668,N_9444);
or U14209 (N_14209,N_9137,N_11056);
nand U14210 (N_14210,N_11776,N_11438);
nor U14211 (N_14211,N_9201,N_9705);
nand U14212 (N_14212,N_9672,N_9254);
and U14213 (N_14213,N_11621,N_9114);
and U14214 (N_14214,N_10209,N_9675);
and U14215 (N_14215,N_11623,N_10474);
nor U14216 (N_14216,N_11030,N_10581);
xnor U14217 (N_14217,N_9112,N_10183);
and U14218 (N_14218,N_11116,N_11396);
and U14219 (N_14219,N_10290,N_11399);
xnor U14220 (N_14220,N_11076,N_11468);
nand U14221 (N_14221,N_11249,N_10263);
nor U14222 (N_14222,N_11125,N_9467);
xor U14223 (N_14223,N_10741,N_11547);
nand U14224 (N_14224,N_10510,N_10551);
nand U14225 (N_14225,N_10949,N_9046);
nand U14226 (N_14226,N_10096,N_9226);
nor U14227 (N_14227,N_10091,N_11511);
nor U14228 (N_14228,N_9462,N_9241);
or U14229 (N_14229,N_10526,N_9243);
xor U14230 (N_14230,N_9297,N_10272);
xor U14231 (N_14231,N_9347,N_9911);
nand U14232 (N_14232,N_9518,N_9661);
xor U14233 (N_14233,N_10104,N_11532);
xor U14234 (N_14234,N_10759,N_10664);
or U14235 (N_14235,N_10219,N_10423);
or U14236 (N_14236,N_9609,N_9708);
xnor U14237 (N_14237,N_10275,N_9993);
nor U14238 (N_14238,N_9848,N_11257);
and U14239 (N_14239,N_10981,N_9231);
nor U14240 (N_14240,N_9330,N_10709);
and U14241 (N_14241,N_10367,N_11552);
nor U14242 (N_14242,N_11766,N_9537);
or U14243 (N_14243,N_9796,N_11969);
xor U14244 (N_14244,N_10824,N_11313);
xor U14245 (N_14245,N_11472,N_9883);
nor U14246 (N_14246,N_10987,N_10035);
xor U14247 (N_14247,N_9270,N_11677);
xnor U14248 (N_14248,N_9435,N_11501);
xor U14249 (N_14249,N_10409,N_10263);
xnor U14250 (N_14250,N_9122,N_9149);
or U14251 (N_14251,N_10880,N_11773);
xnor U14252 (N_14252,N_11344,N_9052);
xor U14253 (N_14253,N_11144,N_10652);
nand U14254 (N_14254,N_10765,N_11494);
or U14255 (N_14255,N_9348,N_10288);
nor U14256 (N_14256,N_9816,N_10842);
nand U14257 (N_14257,N_9263,N_11314);
and U14258 (N_14258,N_9896,N_10168);
nand U14259 (N_14259,N_11358,N_11117);
or U14260 (N_14260,N_11878,N_9918);
xnor U14261 (N_14261,N_10112,N_11262);
and U14262 (N_14262,N_10331,N_10362);
or U14263 (N_14263,N_9078,N_10205);
nand U14264 (N_14264,N_10813,N_9938);
and U14265 (N_14265,N_10885,N_9711);
xnor U14266 (N_14266,N_9624,N_11681);
nor U14267 (N_14267,N_11852,N_11191);
and U14268 (N_14268,N_9004,N_9135);
and U14269 (N_14269,N_11704,N_11671);
or U14270 (N_14270,N_11109,N_11947);
and U14271 (N_14271,N_9866,N_11104);
nand U14272 (N_14272,N_9132,N_9063);
nand U14273 (N_14273,N_9248,N_11288);
or U14274 (N_14274,N_9573,N_11848);
or U14275 (N_14275,N_11045,N_11535);
and U14276 (N_14276,N_10500,N_9366);
or U14277 (N_14277,N_9829,N_11419);
and U14278 (N_14278,N_10469,N_10377);
xnor U14279 (N_14279,N_11950,N_10692);
nor U14280 (N_14280,N_9031,N_10275);
or U14281 (N_14281,N_10004,N_11096);
and U14282 (N_14282,N_11725,N_11719);
and U14283 (N_14283,N_11721,N_10172);
and U14284 (N_14284,N_10941,N_9359);
and U14285 (N_14285,N_9399,N_9741);
and U14286 (N_14286,N_9717,N_9972);
nor U14287 (N_14287,N_10353,N_10031);
nor U14288 (N_14288,N_10939,N_10343);
xor U14289 (N_14289,N_11756,N_11289);
and U14290 (N_14290,N_10977,N_9335);
or U14291 (N_14291,N_11443,N_11293);
and U14292 (N_14292,N_9380,N_9178);
nor U14293 (N_14293,N_10755,N_9815);
or U14294 (N_14294,N_9306,N_10105);
nor U14295 (N_14295,N_9574,N_11983);
and U14296 (N_14296,N_10199,N_10459);
and U14297 (N_14297,N_9414,N_11000);
xnor U14298 (N_14298,N_11300,N_10507);
and U14299 (N_14299,N_10038,N_10437);
xor U14300 (N_14300,N_11934,N_11665);
nand U14301 (N_14301,N_9491,N_10025);
nor U14302 (N_14302,N_9291,N_9769);
nand U14303 (N_14303,N_10446,N_11838);
xnor U14304 (N_14304,N_9134,N_11166);
and U14305 (N_14305,N_9488,N_11662);
or U14306 (N_14306,N_9029,N_11452);
nand U14307 (N_14307,N_10078,N_9183);
nor U14308 (N_14308,N_11951,N_9322);
nand U14309 (N_14309,N_10693,N_10942);
nor U14310 (N_14310,N_9912,N_11419);
nor U14311 (N_14311,N_9029,N_11770);
nor U14312 (N_14312,N_9738,N_11042);
or U14313 (N_14313,N_11994,N_9241);
nand U14314 (N_14314,N_9242,N_10305);
nor U14315 (N_14315,N_10413,N_11100);
or U14316 (N_14316,N_10863,N_9170);
nor U14317 (N_14317,N_10373,N_11351);
xor U14318 (N_14318,N_11333,N_11166);
or U14319 (N_14319,N_11616,N_11244);
nor U14320 (N_14320,N_11902,N_11535);
nand U14321 (N_14321,N_9809,N_11624);
nor U14322 (N_14322,N_10915,N_9808);
or U14323 (N_14323,N_10031,N_11917);
nand U14324 (N_14324,N_10904,N_10281);
nor U14325 (N_14325,N_11891,N_10185);
or U14326 (N_14326,N_9071,N_10779);
xor U14327 (N_14327,N_11750,N_10050);
xnor U14328 (N_14328,N_10665,N_11056);
nor U14329 (N_14329,N_9583,N_11912);
xor U14330 (N_14330,N_11320,N_11734);
xnor U14331 (N_14331,N_11085,N_11590);
nor U14332 (N_14332,N_11248,N_10988);
xnor U14333 (N_14333,N_10508,N_10888);
nor U14334 (N_14334,N_9458,N_10901);
nor U14335 (N_14335,N_9416,N_9878);
nand U14336 (N_14336,N_9588,N_10128);
nand U14337 (N_14337,N_10929,N_11776);
nor U14338 (N_14338,N_11543,N_11056);
xnor U14339 (N_14339,N_11889,N_9407);
or U14340 (N_14340,N_10736,N_11623);
xnor U14341 (N_14341,N_10788,N_9270);
and U14342 (N_14342,N_9585,N_10037);
nor U14343 (N_14343,N_11200,N_11239);
nand U14344 (N_14344,N_9110,N_11024);
nand U14345 (N_14345,N_11572,N_10851);
xnor U14346 (N_14346,N_11587,N_10337);
and U14347 (N_14347,N_9713,N_9217);
xnor U14348 (N_14348,N_9292,N_10772);
xor U14349 (N_14349,N_9222,N_9664);
or U14350 (N_14350,N_10465,N_10967);
nand U14351 (N_14351,N_10963,N_11054);
or U14352 (N_14352,N_9673,N_11801);
and U14353 (N_14353,N_9625,N_11751);
nand U14354 (N_14354,N_9498,N_10939);
and U14355 (N_14355,N_10988,N_11272);
xnor U14356 (N_14356,N_11969,N_10190);
xor U14357 (N_14357,N_10137,N_10338);
xnor U14358 (N_14358,N_10981,N_9788);
and U14359 (N_14359,N_9639,N_9647);
nand U14360 (N_14360,N_10270,N_9367);
nor U14361 (N_14361,N_10659,N_11012);
nor U14362 (N_14362,N_11441,N_10999);
xor U14363 (N_14363,N_11304,N_9380);
or U14364 (N_14364,N_11909,N_11973);
xnor U14365 (N_14365,N_9311,N_9149);
or U14366 (N_14366,N_10551,N_9883);
nor U14367 (N_14367,N_11458,N_9137);
or U14368 (N_14368,N_11279,N_10207);
and U14369 (N_14369,N_11806,N_11216);
xor U14370 (N_14370,N_11307,N_9849);
xor U14371 (N_14371,N_10180,N_11853);
xnor U14372 (N_14372,N_10047,N_9981);
nor U14373 (N_14373,N_11937,N_10255);
nor U14374 (N_14374,N_10619,N_10660);
nor U14375 (N_14375,N_10367,N_10801);
xor U14376 (N_14376,N_9592,N_10449);
xnor U14377 (N_14377,N_10232,N_10267);
or U14378 (N_14378,N_10040,N_9875);
and U14379 (N_14379,N_9213,N_9620);
nor U14380 (N_14380,N_9543,N_11718);
nor U14381 (N_14381,N_10218,N_11622);
or U14382 (N_14382,N_11767,N_9168);
nand U14383 (N_14383,N_9802,N_11170);
and U14384 (N_14384,N_10144,N_10077);
nor U14385 (N_14385,N_10278,N_9409);
or U14386 (N_14386,N_11623,N_10479);
or U14387 (N_14387,N_10099,N_11223);
and U14388 (N_14388,N_11849,N_9527);
or U14389 (N_14389,N_9544,N_10049);
nand U14390 (N_14390,N_11124,N_9853);
and U14391 (N_14391,N_9364,N_11523);
or U14392 (N_14392,N_10262,N_10290);
xor U14393 (N_14393,N_9723,N_11141);
nor U14394 (N_14394,N_11724,N_9093);
and U14395 (N_14395,N_9743,N_10672);
nor U14396 (N_14396,N_11580,N_9153);
nand U14397 (N_14397,N_10915,N_9375);
xor U14398 (N_14398,N_9846,N_9981);
nand U14399 (N_14399,N_9250,N_9043);
xor U14400 (N_14400,N_10354,N_10431);
nor U14401 (N_14401,N_10989,N_9268);
and U14402 (N_14402,N_9054,N_10763);
and U14403 (N_14403,N_11220,N_11036);
nand U14404 (N_14404,N_11386,N_9368);
nand U14405 (N_14405,N_11830,N_10041);
nand U14406 (N_14406,N_9469,N_10157);
nor U14407 (N_14407,N_10419,N_11687);
or U14408 (N_14408,N_11787,N_11299);
and U14409 (N_14409,N_11199,N_9777);
nand U14410 (N_14410,N_11492,N_10365);
or U14411 (N_14411,N_9677,N_10516);
and U14412 (N_14412,N_9742,N_11291);
nand U14413 (N_14413,N_9655,N_11305);
xor U14414 (N_14414,N_11236,N_10042);
and U14415 (N_14415,N_11983,N_10128);
nand U14416 (N_14416,N_9270,N_10754);
and U14417 (N_14417,N_11537,N_11421);
nand U14418 (N_14418,N_10976,N_10467);
or U14419 (N_14419,N_11368,N_11500);
nor U14420 (N_14420,N_10181,N_11108);
and U14421 (N_14421,N_9904,N_10245);
nand U14422 (N_14422,N_9990,N_11953);
nand U14423 (N_14423,N_9899,N_11524);
and U14424 (N_14424,N_10145,N_11523);
and U14425 (N_14425,N_11053,N_11934);
nor U14426 (N_14426,N_11672,N_9813);
nor U14427 (N_14427,N_10859,N_10337);
nand U14428 (N_14428,N_9874,N_11440);
nor U14429 (N_14429,N_11916,N_10088);
and U14430 (N_14430,N_9851,N_10756);
nand U14431 (N_14431,N_9097,N_11879);
or U14432 (N_14432,N_10475,N_11139);
xor U14433 (N_14433,N_10261,N_10461);
xnor U14434 (N_14434,N_10518,N_10885);
nand U14435 (N_14435,N_11393,N_9456);
or U14436 (N_14436,N_11622,N_9085);
nand U14437 (N_14437,N_11473,N_10108);
xnor U14438 (N_14438,N_10341,N_11578);
xor U14439 (N_14439,N_9673,N_9067);
and U14440 (N_14440,N_9022,N_11928);
or U14441 (N_14441,N_9310,N_9205);
xor U14442 (N_14442,N_9403,N_10362);
xnor U14443 (N_14443,N_11263,N_11959);
nor U14444 (N_14444,N_9840,N_9978);
nand U14445 (N_14445,N_11626,N_10334);
and U14446 (N_14446,N_10252,N_9474);
nand U14447 (N_14447,N_9955,N_11388);
and U14448 (N_14448,N_10477,N_11475);
and U14449 (N_14449,N_11114,N_9608);
xor U14450 (N_14450,N_10518,N_9609);
or U14451 (N_14451,N_10141,N_9298);
and U14452 (N_14452,N_11473,N_10383);
nand U14453 (N_14453,N_10527,N_9087);
nand U14454 (N_14454,N_10304,N_11670);
nor U14455 (N_14455,N_9945,N_10072);
nor U14456 (N_14456,N_10470,N_10597);
nor U14457 (N_14457,N_9756,N_11488);
nand U14458 (N_14458,N_11868,N_9307);
xnor U14459 (N_14459,N_10656,N_10216);
and U14460 (N_14460,N_11236,N_9070);
nand U14461 (N_14461,N_9142,N_11646);
nand U14462 (N_14462,N_9091,N_11759);
or U14463 (N_14463,N_11974,N_10835);
xnor U14464 (N_14464,N_9973,N_9481);
or U14465 (N_14465,N_9505,N_9501);
nand U14466 (N_14466,N_11545,N_9399);
or U14467 (N_14467,N_9002,N_11815);
nor U14468 (N_14468,N_9773,N_9015);
and U14469 (N_14469,N_11556,N_10777);
nor U14470 (N_14470,N_9818,N_10132);
or U14471 (N_14471,N_10984,N_9310);
nand U14472 (N_14472,N_11710,N_11068);
nand U14473 (N_14473,N_9528,N_9530);
or U14474 (N_14474,N_9553,N_11139);
nand U14475 (N_14475,N_9913,N_11765);
or U14476 (N_14476,N_11534,N_10174);
nor U14477 (N_14477,N_10817,N_11759);
and U14478 (N_14478,N_9542,N_9350);
or U14479 (N_14479,N_10084,N_11710);
or U14480 (N_14480,N_9579,N_10740);
and U14481 (N_14481,N_9121,N_10290);
nand U14482 (N_14482,N_10071,N_9306);
and U14483 (N_14483,N_9273,N_11320);
and U14484 (N_14484,N_9857,N_10255);
or U14485 (N_14485,N_9110,N_9553);
and U14486 (N_14486,N_10431,N_9992);
nand U14487 (N_14487,N_10679,N_9876);
and U14488 (N_14488,N_10635,N_10156);
nand U14489 (N_14489,N_11367,N_9161);
xor U14490 (N_14490,N_9274,N_9268);
and U14491 (N_14491,N_10020,N_9206);
or U14492 (N_14492,N_11487,N_10434);
nand U14493 (N_14493,N_11790,N_10125);
xor U14494 (N_14494,N_11746,N_11358);
nor U14495 (N_14495,N_10468,N_11764);
or U14496 (N_14496,N_11294,N_10221);
and U14497 (N_14497,N_11624,N_11824);
xor U14498 (N_14498,N_10048,N_9945);
nor U14499 (N_14499,N_11899,N_9907);
or U14500 (N_14500,N_10544,N_11135);
or U14501 (N_14501,N_10985,N_10113);
nand U14502 (N_14502,N_10418,N_9395);
nand U14503 (N_14503,N_11873,N_10016);
nand U14504 (N_14504,N_11547,N_9226);
xnor U14505 (N_14505,N_11638,N_11045);
nor U14506 (N_14506,N_10190,N_9183);
or U14507 (N_14507,N_9140,N_9785);
or U14508 (N_14508,N_11802,N_9722);
or U14509 (N_14509,N_11778,N_10368);
or U14510 (N_14510,N_10812,N_10845);
xor U14511 (N_14511,N_9622,N_9671);
nor U14512 (N_14512,N_11403,N_9975);
or U14513 (N_14513,N_9768,N_10630);
nand U14514 (N_14514,N_10741,N_10183);
or U14515 (N_14515,N_11777,N_10210);
xnor U14516 (N_14516,N_9754,N_9092);
and U14517 (N_14517,N_9210,N_11924);
nor U14518 (N_14518,N_11507,N_9718);
or U14519 (N_14519,N_9763,N_9247);
nor U14520 (N_14520,N_11385,N_10808);
nor U14521 (N_14521,N_11483,N_9558);
and U14522 (N_14522,N_11139,N_10735);
xnor U14523 (N_14523,N_10987,N_9192);
or U14524 (N_14524,N_10186,N_10303);
xor U14525 (N_14525,N_11091,N_10085);
or U14526 (N_14526,N_10985,N_11690);
and U14527 (N_14527,N_10827,N_10958);
or U14528 (N_14528,N_9597,N_10158);
nor U14529 (N_14529,N_10267,N_9048);
xnor U14530 (N_14530,N_10344,N_11511);
nor U14531 (N_14531,N_10096,N_11157);
or U14532 (N_14532,N_10112,N_10073);
and U14533 (N_14533,N_11863,N_11678);
xnor U14534 (N_14534,N_9268,N_10548);
and U14535 (N_14535,N_11735,N_11362);
nor U14536 (N_14536,N_9065,N_9735);
or U14537 (N_14537,N_9141,N_10263);
nor U14538 (N_14538,N_9093,N_11322);
and U14539 (N_14539,N_10604,N_10527);
nand U14540 (N_14540,N_11681,N_10028);
and U14541 (N_14541,N_9842,N_9098);
nor U14542 (N_14542,N_11393,N_10489);
nand U14543 (N_14543,N_9749,N_9082);
xnor U14544 (N_14544,N_9874,N_10888);
and U14545 (N_14545,N_11152,N_10671);
and U14546 (N_14546,N_10214,N_9215);
nand U14547 (N_14547,N_9811,N_10277);
nand U14548 (N_14548,N_9583,N_9383);
xor U14549 (N_14549,N_11877,N_10110);
or U14550 (N_14550,N_9166,N_11008);
and U14551 (N_14551,N_10314,N_11501);
xnor U14552 (N_14552,N_10725,N_10123);
and U14553 (N_14553,N_9977,N_10211);
and U14554 (N_14554,N_10087,N_11329);
or U14555 (N_14555,N_11918,N_10956);
nand U14556 (N_14556,N_11572,N_10529);
nor U14557 (N_14557,N_11756,N_10664);
xnor U14558 (N_14558,N_9872,N_9210);
nor U14559 (N_14559,N_9453,N_10565);
and U14560 (N_14560,N_11666,N_10779);
and U14561 (N_14561,N_10095,N_9946);
or U14562 (N_14562,N_9210,N_9326);
nor U14563 (N_14563,N_9484,N_10580);
nor U14564 (N_14564,N_10794,N_10507);
xor U14565 (N_14565,N_9299,N_9942);
or U14566 (N_14566,N_10211,N_9464);
xor U14567 (N_14567,N_11108,N_11806);
nor U14568 (N_14568,N_9462,N_9672);
nand U14569 (N_14569,N_11030,N_10417);
and U14570 (N_14570,N_10050,N_9926);
xor U14571 (N_14571,N_9652,N_9709);
and U14572 (N_14572,N_10061,N_10519);
and U14573 (N_14573,N_9249,N_10295);
nor U14574 (N_14574,N_11459,N_9585);
xor U14575 (N_14575,N_10113,N_9819);
xnor U14576 (N_14576,N_9214,N_10647);
xor U14577 (N_14577,N_11493,N_10771);
xnor U14578 (N_14578,N_9987,N_9196);
nor U14579 (N_14579,N_9747,N_11342);
nand U14580 (N_14580,N_11677,N_11771);
nand U14581 (N_14581,N_9346,N_11320);
nor U14582 (N_14582,N_10551,N_10286);
nor U14583 (N_14583,N_10826,N_9475);
xnor U14584 (N_14584,N_9989,N_9181);
or U14585 (N_14585,N_10321,N_9774);
and U14586 (N_14586,N_9697,N_11717);
and U14587 (N_14587,N_11092,N_10645);
nor U14588 (N_14588,N_11342,N_10572);
xnor U14589 (N_14589,N_10294,N_11871);
nor U14590 (N_14590,N_11374,N_10459);
nor U14591 (N_14591,N_11834,N_10601);
nor U14592 (N_14592,N_11525,N_9911);
xor U14593 (N_14593,N_10562,N_9315);
or U14594 (N_14594,N_11069,N_11528);
xnor U14595 (N_14595,N_10741,N_10457);
and U14596 (N_14596,N_10070,N_9969);
xor U14597 (N_14597,N_11968,N_11598);
and U14598 (N_14598,N_9961,N_11868);
or U14599 (N_14599,N_9405,N_10151);
xor U14600 (N_14600,N_11909,N_9544);
nand U14601 (N_14601,N_10527,N_10649);
xnor U14602 (N_14602,N_10878,N_9666);
nor U14603 (N_14603,N_11364,N_9962);
nor U14604 (N_14604,N_9944,N_10379);
xor U14605 (N_14605,N_9546,N_10132);
nand U14606 (N_14606,N_9947,N_10639);
nand U14607 (N_14607,N_10712,N_10940);
nor U14608 (N_14608,N_9914,N_9227);
nor U14609 (N_14609,N_10077,N_9115);
or U14610 (N_14610,N_9306,N_11030);
or U14611 (N_14611,N_9922,N_10348);
and U14612 (N_14612,N_9193,N_9346);
and U14613 (N_14613,N_9390,N_11548);
nor U14614 (N_14614,N_9164,N_11663);
nand U14615 (N_14615,N_10921,N_9765);
or U14616 (N_14616,N_11910,N_10122);
nand U14617 (N_14617,N_9367,N_10436);
xnor U14618 (N_14618,N_10185,N_11529);
nand U14619 (N_14619,N_11312,N_11223);
or U14620 (N_14620,N_9604,N_11270);
xor U14621 (N_14621,N_10242,N_11714);
xnor U14622 (N_14622,N_11192,N_9283);
or U14623 (N_14623,N_11053,N_9129);
xor U14624 (N_14624,N_11733,N_11365);
nand U14625 (N_14625,N_11863,N_10045);
or U14626 (N_14626,N_11216,N_9762);
or U14627 (N_14627,N_9093,N_10508);
or U14628 (N_14628,N_10009,N_10647);
and U14629 (N_14629,N_9180,N_9346);
nor U14630 (N_14630,N_9613,N_10607);
nand U14631 (N_14631,N_9741,N_10030);
xor U14632 (N_14632,N_10043,N_10405);
nand U14633 (N_14633,N_11944,N_10347);
nand U14634 (N_14634,N_11564,N_11487);
nand U14635 (N_14635,N_10054,N_10096);
nand U14636 (N_14636,N_10861,N_11125);
xnor U14637 (N_14637,N_10678,N_10236);
nand U14638 (N_14638,N_11797,N_9685);
and U14639 (N_14639,N_9195,N_10187);
nand U14640 (N_14640,N_10990,N_10229);
and U14641 (N_14641,N_10162,N_11114);
and U14642 (N_14642,N_11479,N_9135);
and U14643 (N_14643,N_11087,N_9422);
or U14644 (N_14644,N_10245,N_10717);
nor U14645 (N_14645,N_10035,N_11919);
nor U14646 (N_14646,N_11828,N_11467);
nor U14647 (N_14647,N_9497,N_10009);
nor U14648 (N_14648,N_11232,N_10348);
xor U14649 (N_14649,N_10130,N_9348);
and U14650 (N_14650,N_11497,N_11649);
and U14651 (N_14651,N_10875,N_10360);
and U14652 (N_14652,N_11080,N_9226);
nand U14653 (N_14653,N_9028,N_11768);
nand U14654 (N_14654,N_10136,N_11120);
and U14655 (N_14655,N_10177,N_11859);
nor U14656 (N_14656,N_10075,N_11557);
and U14657 (N_14657,N_11620,N_11552);
and U14658 (N_14658,N_11181,N_9837);
xor U14659 (N_14659,N_11017,N_9044);
nor U14660 (N_14660,N_9568,N_10522);
nand U14661 (N_14661,N_10683,N_11032);
or U14662 (N_14662,N_10597,N_9547);
nor U14663 (N_14663,N_10613,N_11969);
nand U14664 (N_14664,N_9609,N_9446);
and U14665 (N_14665,N_9584,N_10712);
nor U14666 (N_14666,N_9786,N_11206);
nand U14667 (N_14667,N_9863,N_10644);
nand U14668 (N_14668,N_11516,N_10358);
or U14669 (N_14669,N_9008,N_11205);
and U14670 (N_14670,N_10310,N_11945);
nand U14671 (N_14671,N_9579,N_9386);
nor U14672 (N_14672,N_9157,N_10729);
and U14673 (N_14673,N_11070,N_9221);
and U14674 (N_14674,N_10865,N_9613);
and U14675 (N_14675,N_11939,N_11400);
xnor U14676 (N_14676,N_9636,N_11466);
or U14677 (N_14677,N_9804,N_11029);
nor U14678 (N_14678,N_9494,N_10454);
and U14679 (N_14679,N_9460,N_9956);
nor U14680 (N_14680,N_11485,N_11941);
nor U14681 (N_14681,N_11901,N_10472);
nand U14682 (N_14682,N_11336,N_9595);
xnor U14683 (N_14683,N_10802,N_9874);
xor U14684 (N_14684,N_11806,N_11836);
nand U14685 (N_14685,N_9385,N_10407);
nand U14686 (N_14686,N_11788,N_10626);
nor U14687 (N_14687,N_10818,N_9611);
nor U14688 (N_14688,N_11566,N_10307);
and U14689 (N_14689,N_11133,N_11093);
xnor U14690 (N_14690,N_11876,N_10358);
or U14691 (N_14691,N_10437,N_9496);
xor U14692 (N_14692,N_9677,N_9879);
nor U14693 (N_14693,N_9149,N_9713);
nand U14694 (N_14694,N_9410,N_9895);
xnor U14695 (N_14695,N_10714,N_11362);
nor U14696 (N_14696,N_10698,N_10936);
and U14697 (N_14697,N_9016,N_10911);
nand U14698 (N_14698,N_11084,N_11550);
nor U14699 (N_14699,N_11979,N_11647);
and U14700 (N_14700,N_10776,N_9766);
nor U14701 (N_14701,N_11633,N_10831);
or U14702 (N_14702,N_9875,N_10983);
or U14703 (N_14703,N_9585,N_9335);
and U14704 (N_14704,N_11576,N_10584);
xnor U14705 (N_14705,N_10993,N_10334);
and U14706 (N_14706,N_9635,N_11342);
or U14707 (N_14707,N_9065,N_11247);
nor U14708 (N_14708,N_9488,N_11470);
nor U14709 (N_14709,N_10643,N_10325);
and U14710 (N_14710,N_10583,N_10641);
nand U14711 (N_14711,N_10742,N_11231);
nor U14712 (N_14712,N_9127,N_11717);
nand U14713 (N_14713,N_10256,N_11241);
or U14714 (N_14714,N_11726,N_10923);
nor U14715 (N_14715,N_11321,N_9741);
and U14716 (N_14716,N_9726,N_11232);
xnor U14717 (N_14717,N_9384,N_10350);
nand U14718 (N_14718,N_9262,N_9658);
nor U14719 (N_14719,N_9555,N_9528);
or U14720 (N_14720,N_10874,N_11128);
or U14721 (N_14721,N_10957,N_11370);
nand U14722 (N_14722,N_10078,N_10799);
nor U14723 (N_14723,N_10784,N_11905);
nand U14724 (N_14724,N_10233,N_10489);
nor U14725 (N_14725,N_11039,N_11257);
and U14726 (N_14726,N_9891,N_11987);
nand U14727 (N_14727,N_10177,N_9558);
or U14728 (N_14728,N_10659,N_11281);
or U14729 (N_14729,N_9840,N_10665);
xnor U14730 (N_14730,N_9715,N_10210);
and U14731 (N_14731,N_11718,N_11311);
and U14732 (N_14732,N_10479,N_10982);
xnor U14733 (N_14733,N_11252,N_10518);
nand U14734 (N_14734,N_9929,N_11472);
or U14735 (N_14735,N_10454,N_9956);
or U14736 (N_14736,N_11599,N_11531);
nor U14737 (N_14737,N_9223,N_9502);
nand U14738 (N_14738,N_11374,N_9303);
and U14739 (N_14739,N_10834,N_9547);
or U14740 (N_14740,N_11809,N_11773);
xor U14741 (N_14741,N_10080,N_10066);
or U14742 (N_14742,N_9551,N_10715);
nand U14743 (N_14743,N_10220,N_11690);
or U14744 (N_14744,N_9884,N_10550);
and U14745 (N_14745,N_11313,N_10249);
or U14746 (N_14746,N_10410,N_10010);
nor U14747 (N_14747,N_10165,N_11741);
or U14748 (N_14748,N_9446,N_11339);
nand U14749 (N_14749,N_9617,N_11501);
nand U14750 (N_14750,N_11702,N_9972);
nor U14751 (N_14751,N_10171,N_10258);
or U14752 (N_14752,N_11960,N_11859);
or U14753 (N_14753,N_11517,N_9555);
nor U14754 (N_14754,N_10994,N_10304);
nor U14755 (N_14755,N_11731,N_11053);
nor U14756 (N_14756,N_11478,N_9984);
xnor U14757 (N_14757,N_10916,N_11672);
nor U14758 (N_14758,N_10998,N_9831);
xor U14759 (N_14759,N_11171,N_10861);
nor U14760 (N_14760,N_9213,N_10999);
or U14761 (N_14761,N_10333,N_11075);
and U14762 (N_14762,N_9213,N_10783);
or U14763 (N_14763,N_10221,N_9762);
and U14764 (N_14764,N_11750,N_11118);
or U14765 (N_14765,N_9296,N_11042);
nor U14766 (N_14766,N_11791,N_10020);
and U14767 (N_14767,N_9608,N_10045);
nor U14768 (N_14768,N_9947,N_9599);
or U14769 (N_14769,N_10198,N_11424);
and U14770 (N_14770,N_9360,N_10825);
nor U14771 (N_14771,N_10332,N_11704);
or U14772 (N_14772,N_9335,N_11603);
xnor U14773 (N_14773,N_10061,N_10787);
nand U14774 (N_14774,N_10982,N_10321);
nand U14775 (N_14775,N_9875,N_9639);
xnor U14776 (N_14776,N_9660,N_11389);
and U14777 (N_14777,N_9236,N_10643);
nand U14778 (N_14778,N_9763,N_9576);
xnor U14779 (N_14779,N_11979,N_10302);
nand U14780 (N_14780,N_10754,N_10648);
nor U14781 (N_14781,N_10972,N_9615);
and U14782 (N_14782,N_9332,N_11958);
nand U14783 (N_14783,N_10235,N_9579);
and U14784 (N_14784,N_9893,N_10252);
or U14785 (N_14785,N_10939,N_11361);
nand U14786 (N_14786,N_9636,N_9347);
or U14787 (N_14787,N_10254,N_9877);
nand U14788 (N_14788,N_10967,N_10884);
nand U14789 (N_14789,N_11954,N_10083);
or U14790 (N_14790,N_11656,N_9884);
xor U14791 (N_14791,N_9986,N_11179);
or U14792 (N_14792,N_11273,N_11536);
nor U14793 (N_14793,N_11048,N_11106);
xnor U14794 (N_14794,N_10658,N_11470);
xnor U14795 (N_14795,N_10034,N_9076);
or U14796 (N_14796,N_9104,N_10357);
nor U14797 (N_14797,N_10976,N_10336);
nand U14798 (N_14798,N_9424,N_11380);
nand U14799 (N_14799,N_10323,N_9725);
and U14800 (N_14800,N_11823,N_10399);
xor U14801 (N_14801,N_9315,N_9103);
xnor U14802 (N_14802,N_10500,N_11014);
nand U14803 (N_14803,N_11967,N_11965);
nand U14804 (N_14804,N_9319,N_11261);
or U14805 (N_14805,N_10278,N_10300);
and U14806 (N_14806,N_9573,N_10083);
nand U14807 (N_14807,N_10428,N_10101);
and U14808 (N_14808,N_9889,N_10973);
or U14809 (N_14809,N_11349,N_11358);
nand U14810 (N_14810,N_11859,N_11537);
xnor U14811 (N_14811,N_10478,N_10760);
nand U14812 (N_14812,N_9201,N_11017);
or U14813 (N_14813,N_11503,N_11803);
xnor U14814 (N_14814,N_10262,N_10753);
and U14815 (N_14815,N_9523,N_9570);
nor U14816 (N_14816,N_11318,N_9417);
nor U14817 (N_14817,N_9659,N_11683);
nor U14818 (N_14818,N_11589,N_10711);
nor U14819 (N_14819,N_11934,N_11021);
xor U14820 (N_14820,N_9835,N_10983);
xnor U14821 (N_14821,N_10719,N_9146);
xor U14822 (N_14822,N_11474,N_9729);
nand U14823 (N_14823,N_11525,N_9800);
nand U14824 (N_14824,N_10869,N_11507);
xor U14825 (N_14825,N_9079,N_11918);
nor U14826 (N_14826,N_10450,N_9096);
and U14827 (N_14827,N_10291,N_9217);
and U14828 (N_14828,N_9503,N_9613);
xor U14829 (N_14829,N_10367,N_10409);
or U14830 (N_14830,N_11318,N_11060);
or U14831 (N_14831,N_11610,N_9253);
nor U14832 (N_14832,N_9633,N_11780);
or U14833 (N_14833,N_9386,N_11421);
or U14834 (N_14834,N_10806,N_11406);
xor U14835 (N_14835,N_11505,N_10931);
and U14836 (N_14836,N_11800,N_9159);
or U14837 (N_14837,N_10776,N_10868);
and U14838 (N_14838,N_11278,N_10904);
xor U14839 (N_14839,N_10682,N_11345);
nor U14840 (N_14840,N_11960,N_10255);
and U14841 (N_14841,N_11210,N_11113);
nand U14842 (N_14842,N_11557,N_11064);
nand U14843 (N_14843,N_9091,N_10770);
xnor U14844 (N_14844,N_11494,N_9410);
and U14845 (N_14845,N_11121,N_11222);
or U14846 (N_14846,N_10925,N_10764);
or U14847 (N_14847,N_9357,N_10277);
nor U14848 (N_14848,N_9756,N_11146);
or U14849 (N_14849,N_10896,N_11732);
nand U14850 (N_14850,N_11734,N_10694);
nor U14851 (N_14851,N_9021,N_10158);
nand U14852 (N_14852,N_9682,N_9889);
xor U14853 (N_14853,N_11173,N_11782);
xnor U14854 (N_14854,N_10726,N_10270);
and U14855 (N_14855,N_10022,N_9075);
or U14856 (N_14856,N_10562,N_10082);
xnor U14857 (N_14857,N_10378,N_9149);
or U14858 (N_14858,N_11547,N_10733);
and U14859 (N_14859,N_11618,N_10302);
nand U14860 (N_14860,N_10331,N_10473);
nor U14861 (N_14861,N_11582,N_11432);
xor U14862 (N_14862,N_9879,N_9874);
or U14863 (N_14863,N_10146,N_11893);
xnor U14864 (N_14864,N_9112,N_9714);
nor U14865 (N_14865,N_11017,N_11047);
xnor U14866 (N_14866,N_10834,N_11204);
and U14867 (N_14867,N_9714,N_11533);
nand U14868 (N_14868,N_11124,N_9568);
xnor U14869 (N_14869,N_9225,N_10054);
nor U14870 (N_14870,N_10081,N_10429);
and U14871 (N_14871,N_11503,N_10219);
nor U14872 (N_14872,N_9579,N_11950);
xor U14873 (N_14873,N_10240,N_10513);
xor U14874 (N_14874,N_11914,N_9358);
nand U14875 (N_14875,N_10682,N_11195);
or U14876 (N_14876,N_11284,N_10082);
nor U14877 (N_14877,N_10481,N_10439);
xnor U14878 (N_14878,N_11027,N_11288);
xnor U14879 (N_14879,N_9564,N_11549);
nor U14880 (N_14880,N_11180,N_10755);
and U14881 (N_14881,N_10167,N_10362);
nand U14882 (N_14882,N_10317,N_10251);
nor U14883 (N_14883,N_10708,N_10120);
xor U14884 (N_14884,N_11500,N_11959);
and U14885 (N_14885,N_11014,N_11543);
xor U14886 (N_14886,N_11016,N_11554);
nor U14887 (N_14887,N_9258,N_9594);
and U14888 (N_14888,N_10982,N_11233);
and U14889 (N_14889,N_11247,N_11808);
or U14890 (N_14890,N_11273,N_9757);
and U14891 (N_14891,N_9949,N_11445);
nand U14892 (N_14892,N_11821,N_9570);
and U14893 (N_14893,N_9602,N_10422);
nor U14894 (N_14894,N_9041,N_10483);
nand U14895 (N_14895,N_9280,N_10767);
and U14896 (N_14896,N_10496,N_11304);
nand U14897 (N_14897,N_10350,N_9298);
nor U14898 (N_14898,N_11036,N_10474);
and U14899 (N_14899,N_9585,N_9046);
xor U14900 (N_14900,N_9483,N_10248);
xor U14901 (N_14901,N_10198,N_9426);
and U14902 (N_14902,N_11458,N_11072);
xor U14903 (N_14903,N_9830,N_11941);
or U14904 (N_14904,N_10522,N_9198);
and U14905 (N_14905,N_11248,N_10322);
or U14906 (N_14906,N_9801,N_10889);
nand U14907 (N_14907,N_11580,N_10392);
or U14908 (N_14908,N_11681,N_9813);
or U14909 (N_14909,N_9384,N_11506);
and U14910 (N_14910,N_11636,N_9404);
and U14911 (N_14911,N_9266,N_10892);
and U14912 (N_14912,N_11241,N_9180);
nor U14913 (N_14913,N_9298,N_10589);
and U14914 (N_14914,N_11056,N_11551);
or U14915 (N_14915,N_9707,N_11362);
or U14916 (N_14916,N_11390,N_11379);
nor U14917 (N_14917,N_11943,N_10434);
and U14918 (N_14918,N_9103,N_11164);
nor U14919 (N_14919,N_10845,N_10380);
or U14920 (N_14920,N_9469,N_11046);
nand U14921 (N_14921,N_9551,N_10864);
xor U14922 (N_14922,N_11000,N_10167);
and U14923 (N_14923,N_11069,N_11841);
nand U14924 (N_14924,N_10246,N_11411);
or U14925 (N_14925,N_9896,N_10403);
and U14926 (N_14926,N_10289,N_9231);
and U14927 (N_14927,N_9482,N_10993);
nor U14928 (N_14928,N_9135,N_10624);
nand U14929 (N_14929,N_9483,N_10070);
xnor U14930 (N_14930,N_11511,N_10566);
and U14931 (N_14931,N_9584,N_10826);
nand U14932 (N_14932,N_9797,N_9524);
and U14933 (N_14933,N_10881,N_11578);
nand U14934 (N_14934,N_10449,N_10603);
or U14935 (N_14935,N_11664,N_9279);
or U14936 (N_14936,N_9903,N_11058);
nor U14937 (N_14937,N_9874,N_9454);
xor U14938 (N_14938,N_11060,N_10655);
or U14939 (N_14939,N_10082,N_10223);
nor U14940 (N_14940,N_10119,N_11227);
or U14941 (N_14941,N_11689,N_11656);
nor U14942 (N_14942,N_11674,N_10960);
and U14943 (N_14943,N_10222,N_11615);
nor U14944 (N_14944,N_10438,N_10870);
or U14945 (N_14945,N_11799,N_11411);
nand U14946 (N_14946,N_9825,N_10404);
xnor U14947 (N_14947,N_10737,N_11821);
nand U14948 (N_14948,N_11312,N_11922);
and U14949 (N_14949,N_10150,N_9917);
xnor U14950 (N_14950,N_11494,N_9326);
nor U14951 (N_14951,N_9903,N_9196);
nand U14952 (N_14952,N_10708,N_10308);
nand U14953 (N_14953,N_11654,N_10525);
nand U14954 (N_14954,N_9676,N_11050);
or U14955 (N_14955,N_11400,N_11418);
or U14956 (N_14956,N_9676,N_10816);
and U14957 (N_14957,N_10285,N_11111);
nor U14958 (N_14958,N_10458,N_10200);
xor U14959 (N_14959,N_9441,N_11160);
xor U14960 (N_14960,N_9121,N_10855);
nor U14961 (N_14961,N_9217,N_11200);
xor U14962 (N_14962,N_11125,N_9931);
xnor U14963 (N_14963,N_10536,N_11377);
and U14964 (N_14964,N_9723,N_10599);
nand U14965 (N_14965,N_11181,N_9532);
nand U14966 (N_14966,N_10448,N_11374);
and U14967 (N_14967,N_9484,N_10285);
and U14968 (N_14968,N_10538,N_9745);
nand U14969 (N_14969,N_10849,N_11317);
xor U14970 (N_14970,N_11111,N_10786);
nor U14971 (N_14971,N_9818,N_11746);
or U14972 (N_14972,N_11582,N_11291);
nor U14973 (N_14973,N_11358,N_9551);
and U14974 (N_14974,N_9473,N_10221);
and U14975 (N_14975,N_9184,N_10115);
nor U14976 (N_14976,N_11921,N_11500);
or U14977 (N_14977,N_9242,N_9359);
or U14978 (N_14978,N_10546,N_9412);
xnor U14979 (N_14979,N_9808,N_9111);
xor U14980 (N_14980,N_11308,N_11509);
and U14981 (N_14981,N_11491,N_11107);
nor U14982 (N_14982,N_10900,N_9963);
nand U14983 (N_14983,N_9770,N_11066);
nand U14984 (N_14984,N_11913,N_10339);
xor U14985 (N_14985,N_9353,N_11889);
or U14986 (N_14986,N_11971,N_9427);
or U14987 (N_14987,N_11266,N_11936);
xor U14988 (N_14988,N_11442,N_9338);
or U14989 (N_14989,N_9813,N_9273);
nand U14990 (N_14990,N_11746,N_11516);
or U14991 (N_14991,N_10132,N_10727);
and U14992 (N_14992,N_11850,N_11301);
nor U14993 (N_14993,N_9460,N_9804);
and U14994 (N_14994,N_11785,N_11735);
nand U14995 (N_14995,N_11414,N_9743);
or U14996 (N_14996,N_9916,N_11309);
nand U14997 (N_14997,N_10039,N_10160);
nor U14998 (N_14998,N_10868,N_11065);
and U14999 (N_14999,N_11984,N_9634);
or UO_0 (O_0,N_13069,N_13802);
nor UO_1 (O_1,N_13732,N_13164);
xnor UO_2 (O_2,N_13443,N_13603);
xnor UO_3 (O_3,N_12481,N_14780);
nor UO_4 (O_4,N_13765,N_13537);
xnor UO_5 (O_5,N_12941,N_14393);
nand UO_6 (O_6,N_14590,N_12128);
or UO_7 (O_7,N_13689,N_13968);
nor UO_8 (O_8,N_12273,N_12446);
nand UO_9 (O_9,N_14748,N_12110);
nor UO_10 (O_10,N_12862,N_14222);
nor UO_11 (O_11,N_13416,N_13769);
nor UO_12 (O_12,N_13155,N_14992);
xnor UO_13 (O_13,N_12838,N_13333);
nor UO_14 (O_14,N_14781,N_13812);
xnor UO_15 (O_15,N_12058,N_14887);
nand UO_16 (O_16,N_14181,N_12097);
nor UO_17 (O_17,N_14046,N_14760);
or UO_18 (O_18,N_14001,N_12482);
and UO_19 (O_19,N_14220,N_14671);
xor UO_20 (O_20,N_14660,N_14014);
xor UO_21 (O_21,N_13612,N_14356);
xnor UO_22 (O_22,N_14951,N_12550);
nor UO_23 (O_23,N_14667,N_12002);
nand UO_24 (O_24,N_14471,N_13144);
nand UO_25 (O_25,N_14280,N_14541);
or UO_26 (O_26,N_13276,N_13924);
and UO_27 (O_27,N_13198,N_12106);
nand UO_28 (O_28,N_14158,N_13727);
xor UO_29 (O_29,N_13264,N_12172);
xor UO_30 (O_30,N_14387,N_14459);
or UO_31 (O_31,N_14658,N_13022);
nand UO_32 (O_32,N_14940,N_14188);
nor UO_33 (O_33,N_12246,N_12994);
nand UO_34 (O_34,N_13967,N_13141);
nand UO_35 (O_35,N_13632,N_14059);
nor UO_36 (O_36,N_13799,N_14576);
nand UO_37 (O_37,N_14410,N_13648);
or UO_38 (O_38,N_14907,N_14699);
and UO_39 (O_39,N_12478,N_14701);
and UO_40 (O_40,N_14479,N_14696);
nand UO_41 (O_41,N_13808,N_13975);
nand UO_42 (O_42,N_14710,N_14661);
xnor UO_43 (O_43,N_14806,N_12056);
nor UO_44 (O_44,N_12256,N_13840);
nand UO_45 (O_45,N_13228,N_14927);
nor UO_46 (O_46,N_13890,N_12865);
nand UO_47 (O_47,N_12803,N_13722);
and UO_48 (O_48,N_13342,N_14881);
and UO_49 (O_49,N_12393,N_12366);
nand UO_50 (O_50,N_12340,N_13123);
and UO_51 (O_51,N_12894,N_14509);
nand UO_52 (O_52,N_14125,N_12285);
xnor UO_53 (O_53,N_13025,N_13281);
or UO_54 (O_54,N_14859,N_13665);
xor UO_55 (O_55,N_12274,N_14982);
or UO_56 (O_56,N_13387,N_13598);
xnor UO_57 (O_57,N_14451,N_13306);
or UO_58 (O_58,N_12013,N_12713);
and UO_59 (O_59,N_14706,N_13704);
nor UO_60 (O_60,N_14104,N_13856);
xor UO_61 (O_61,N_12444,N_12221);
xnor UO_62 (O_62,N_13271,N_14558);
nor UO_63 (O_63,N_14894,N_14013);
xnor UO_64 (O_64,N_14225,N_14552);
or UO_65 (O_65,N_12328,N_12595);
or UO_66 (O_66,N_13922,N_14849);
and UO_67 (O_67,N_14758,N_13772);
nand UO_68 (O_68,N_13724,N_13480);
and UO_69 (O_69,N_12922,N_12122);
xor UO_70 (O_70,N_14553,N_13503);
nand UO_71 (O_71,N_12462,N_13458);
or UO_72 (O_72,N_14350,N_12017);
xor UO_73 (O_73,N_13135,N_13662);
and UO_74 (O_74,N_14914,N_13191);
nor UO_75 (O_75,N_13606,N_12611);
nor UO_76 (O_76,N_12327,N_12660);
and UO_77 (O_77,N_14581,N_14999);
or UO_78 (O_78,N_13292,N_13446);
xnor UO_79 (O_79,N_14926,N_14400);
xnor UO_80 (O_80,N_12488,N_13054);
or UO_81 (O_81,N_12282,N_13422);
nand UO_82 (O_82,N_13705,N_14233);
xor UO_83 (O_83,N_12402,N_12745);
xor UO_84 (O_84,N_14270,N_14729);
nor UO_85 (O_85,N_12010,N_13398);
nand UO_86 (O_86,N_12333,N_13302);
and UO_87 (O_87,N_12014,N_12099);
and UO_88 (O_88,N_12403,N_12652);
xor UO_89 (O_89,N_13644,N_12319);
and UO_90 (O_90,N_12294,N_13110);
and UO_91 (O_91,N_12781,N_12492);
and UO_92 (O_92,N_13921,N_13027);
nor UO_93 (O_93,N_13927,N_14040);
or UO_94 (O_94,N_12170,N_14259);
or UO_95 (O_95,N_13677,N_13592);
xor UO_96 (O_96,N_14353,N_12495);
xor UO_97 (O_97,N_12680,N_14656);
xor UO_98 (O_98,N_12020,N_13622);
or UO_99 (O_99,N_14402,N_13210);
xor UO_100 (O_100,N_14620,N_14885);
xnor UO_101 (O_101,N_12460,N_13623);
and UO_102 (O_102,N_14634,N_12456);
xnor UO_103 (O_103,N_12912,N_12773);
nor UO_104 (O_104,N_13989,N_14812);
nor UO_105 (O_105,N_13279,N_14399);
nand UO_106 (O_106,N_13997,N_13450);
and UO_107 (O_107,N_12578,N_12353);
nor UO_108 (O_108,N_12640,N_14480);
nand UO_109 (O_109,N_12939,N_12078);
nand UO_110 (O_110,N_13148,N_12769);
nand UO_111 (O_111,N_12432,N_13950);
nand UO_112 (O_112,N_14682,N_13243);
nor UO_113 (O_113,N_12793,N_13290);
or UO_114 (O_114,N_12766,N_13096);
nand UO_115 (O_115,N_12591,N_12755);
nor UO_116 (O_116,N_12417,N_13002);
nor UO_117 (O_117,N_12921,N_12301);
nand UO_118 (O_118,N_13958,N_14787);
nand UO_119 (O_119,N_14303,N_13238);
xor UO_120 (O_120,N_13730,N_12725);
or UO_121 (O_121,N_13426,N_14315);
nor UO_122 (O_122,N_12733,N_12396);
nand UO_123 (O_123,N_12180,N_13282);
nor UO_124 (O_124,N_14937,N_12083);
xnor UO_125 (O_125,N_12545,N_14955);
and UO_126 (O_126,N_13520,N_12798);
nor UO_127 (O_127,N_14079,N_12253);
or UO_128 (O_128,N_13587,N_14426);
nand UO_129 (O_129,N_12121,N_12604);
or UO_130 (O_130,N_13857,N_14562);
xnor UO_131 (O_131,N_14377,N_13931);
xor UO_132 (O_132,N_14067,N_14120);
xnor UO_133 (O_133,N_14083,N_12928);
or UO_134 (O_134,N_13378,N_13639);
nor UO_135 (O_135,N_12951,N_12698);
or UO_136 (O_136,N_13809,N_13483);
or UO_137 (O_137,N_12620,N_14271);
and UO_138 (O_138,N_13265,N_14779);
and UO_139 (O_139,N_14853,N_12981);
nor UO_140 (O_140,N_14134,N_12131);
and UO_141 (O_141,N_12592,N_13355);
nand UO_142 (O_142,N_12138,N_14746);
xnor UO_143 (O_143,N_13829,N_14602);
and UO_144 (O_144,N_14476,N_14776);
nor UO_145 (O_145,N_13911,N_13261);
xnor UO_146 (O_146,N_12947,N_12326);
or UO_147 (O_147,N_13330,N_12788);
or UO_148 (O_148,N_13915,N_13147);
nand UO_149 (O_149,N_14938,N_13266);
nor UO_150 (O_150,N_12119,N_13964);
xor UO_151 (O_151,N_14213,N_12305);
nand UO_152 (O_152,N_13115,N_13886);
nor UO_153 (O_153,N_12331,N_12964);
or UO_154 (O_154,N_12452,N_13636);
nand UO_155 (O_155,N_12292,N_13288);
xnor UO_156 (O_156,N_13381,N_12324);
xnor UO_157 (O_157,N_14146,N_12231);
nand UO_158 (O_158,N_13617,N_12001);
nor UO_159 (O_159,N_14441,N_12581);
nand UO_160 (O_160,N_12892,N_13117);
xnor UO_161 (O_161,N_13506,N_13366);
and UO_162 (O_162,N_12323,N_13647);
or UO_163 (O_163,N_14008,N_14644);
xor UO_164 (O_164,N_12734,N_14916);
xor UO_165 (O_165,N_13862,N_12156);
nor UO_166 (O_166,N_14111,N_12743);
or UO_167 (O_167,N_14973,N_13717);
and UO_168 (O_168,N_12489,N_14692);
xor UO_169 (O_169,N_12671,N_12779);
xor UO_170 (O_170,N_14738,N_13373);
and UO_171 (O_171,N_14063,N_14740);
or UO_172 (O_172,N_14736,N_12117);
nor UO_173 (O_173,N_12179,N_14137);
and UO_174 (O_174,N_12057,N_12872);
xor UO_175 (O_175,N_12384,N_13894);
nor UO_176 (O_176,N_14680,N_14767);
or UO_177 (O_177,N_14484,N_13709);
or UO_178 (O_178,N_12206,N_12223);
and UO_179 (O_179,N_14580,N_12435);
xnor UO_180 (O_180,N_12840,N_14338);
xnor UO_181 (O_181,N_12561,N_14604);
nand UO_182 (O_182,N_14172,N_13203);
or UO_183 (O_183,N_14482,N_13309);
and UO_184 (O_184,N_14318,N_13729);
nor UO_185 (O_185,N_12051,N_13254);
and UO_186 (O_186,N_13643,N_12932);
nand UO_187 (O_187,N_13868,N_12351);
nor UO_188 (O_188,N_12350,N_13297);
nor UO_189 (O_189,N_13905,N_12069);
and UO_190 (O_190,N_12505,N_14573);
and UO_191 (O_191,N_13684,N_14783);
xor UO_192 (O_192,N_14336,N_13431);
and UO_193 (O_193,N_13456,N_14072);
nand UO_194 (O_194,N_14022,N_12881);
or UO_195 (O_195,N_12439,N_14769);
nand UO_196 (O_196,N_12919,N_13285);
or UO_197 (O_197,N_12562,N_12100);
xor UO_198 (O_198,N_12085,N_14114);
nand UO_199 (O_199,N_12012,N_13738);
or UO_200 (O_200,N_13143,N_12685);
or UO_201 (O_201,N_12816,N_14249);
and UO_202 (O_202,N_14035,N_13980);
or UO_203 (O_203,N_13269,N_14845);
or UO_204 (O_204,N_12699,N_14086);
xor UO_205 (O_205,N_13917,N_14897);
xnor UO_206 (O_206,N_12307,N_12955);
xnor UO_207 (O_207,N_14678,N_14985);
nor UO_208 (O_208,N_12946,N_14129);
and UO_209 (O_209,N_14613,N_13364);
nand UO_210 (O_210,N_13670,N_13861);
nand UO_211 (O_211,N_13928,N_14852);
nand UO_212 (O_212,N_13409,N_14351);
or UO_213 (O_213,N_13694,N_13523);
xnor UO_214 (O_214,N_14798,N_12169);
xnor UO_215 (O_215,N_13019,N_12015);
or UO_216 (O_216,N_13360,N_13901);
nor UO_217 (O_217,N_14669,N_12686);
nand UO_218 (O_218,N_12414,N_13659);
xor UO_219 (O_219,N_13920,N_13800);
xor UO_220 (O_220,N_13348,N_12244);
nand UO_221 (O_221,N_12287,N_14339);
and UO_222 (O_222,N_14077,N_14737);
xnor UO_223 (O_223,N_14386,N_14851);
and UO_224 (O_224,N_14786,N_12607);
or UO_225 (O_225,N_12860,N_14390);
xnor UO_226 (O_226,N_12339,N_12280);
xnor UO_227 (O_227,N_14159,N_13108);
xnor UO_228 (O_228,N_14878,N_12185);
or UO_229 (O_229,N_13655,N_12814);
or UO_230 (O_230,N_12571,N_13242);
nand UO_231 (O_231,N_13936,N_12893);
nand UO_232 (O_232,N_13516,N_14931);
or UO_233 (O_233,N_14090,N_13500);
xor UO_234 (O_234,N_14643,N_14266);
or UO_235 (O_235,N_14630,N_13628);
or UO_236 (O_236,N_12035,N_14957);
xnor UO_237 (O_237,N_12968,N_13103);
xnor UO_238 (O_238,N_13338,N_12126);
xor UO_239 (O_239,N_12810,N_13011);
and UO_240 (O_240,N_12220,N_12406);
xnor UO_241 (O_241,N_14205,N_12796);
xor UO_242 (O_242,N_13043,N_12942);
nor UO_243 (O_243,N_12885,N_14272);
nor UO_244 (O_244,N_14860,N_13166);
nor UO_245 (O_245,N_13412,N_14969);
and UO_246 (O_246,N_13759,N_13873);
or UO_247 (O_247,N_13579,N_13838);
nor UO_248 (O_248,N_12011,N_13385);
or UO_249 (O_249,N_13491,N_13310);
nor UO_250 (O_250,N_12874,N_13009);
and UO_251 (O_251,N_12768,N_13444);
xor UO_252 (O_252,N_14599,N_12954);
and UO_253 (O_253,N_14516,N_13695);
or UO_254 (O_254,N_14028,N_13651);
xnor UO_255 (O_255,N_12024,N_14385);
and UO_256 (O_256,N_13086,N_13353);
or UO_257 (O_257,N_13082,N_13252);
and UO_258 (O_258,N_14717,N_14942);
nand UO_259 (O_259,N_14713,N_12976);
nand UO_260 (O_260,N_13239,N_14444);
xnor UO_261 (O_261,N_12643,N_12088);
xor UO_262 (O_262,N_12356,N_14021);
nand UO_263 (O_263,N_12689,N_14133);
or UO_264 (O_264,N_14989,N_13566);
xor UO_265 (O_265,N_12225,N_14415);
xor UO_266 (O_266,N_14361,N_12970);
xnor UO_267 (O_267,N_12649,N_14053);
nand UO_268 (O_268,N_12792,N_13347);
xor UO_269 (O_269,N_12802,N_13781);
nor UO_270 (O_270,N_14797,N_13492);
and UO_271 (O_271,N_14827,N_12040);
nor UO_272 (O_272,N_13418,N_14189);
nand UO_273 (O_273,N_12458,N_14847);
or UO_274 (O_274,N_12259,N_13847);
nor UO_275 (O_275,N_14978,N_12050);
nand UO_276 (O_276,N_12383,N_14337);
nand UO_277 (O_277,N_14226,N_13559);
and UO_278 (O_278,N_12746,N_12152);
nand UO_279 (O_279,N_14921,N_12261);
xor UO_280 (O_280,N_12585,N_14378);
xnor UO_281 (O_281,N_13599,N_12335);
and UO_282 (O_282,N_14879,N_14091);
xor UO_283 (O_283,N_13780,N_12381);
nor UO_284 (O_284,N_14347,N_14681);
or UO_285 (O_285,N_13795,N_14081);
xnor UO_286 (O_286,N_14100,N_12778);
and UO_287 (O_287,N_13126,N_14408);
nor UO_288 (O_288,N_13097,N_13206);
or UO_289 (O_289,N_14018,N_12330);
or UO_290 (O_290,N_13919,N_13359);
xnor UO_291 (O_291,N_14200,N_12853);
xor UO_292 (O_292,N_14813,N_13212);
nor UO_293 (O_293,N_12120,N_13748);
and UO_294 (O_294,N_13291,N_12887);
nor UO_295 (O_295,N_14355,N_14504);
nor UO_296 (O_296,N_12210,N_14944);
nor UO_297 (O_297,N_12520,N_13754);
or UO_298 (O_298,N_14398,N_12760);
or UO_299 (O_299,N_12003,N_14301);
and UO_300 (O_300,N_14972,N_12851);
nand UO_301 (O_301,N_14550,N_13014);
and UO_302 (O_302,N_13529,N_12855);
xnor UO_303 (O_303,N_13199,N_14841);
xor UO_304 (O_304,N_12412,N_14169);
nor UO_305 (O_305,N_13033,N_13318);
or UO_306 (O_306,N_12647,N_13156);
and UO_307 (O_307,N_14324,N_12538);
xnor UO_308 (O_308,N_13224,N_13904);
or UO_309 (O_309,N_13358,N_13070);
xnor UO_310 (O_310,N_12199,N_14427);
nor UO_311 (O_311,N_14606,N_12943);
or UO_312 (O_312,N_14011,N_13273);
or UO_313 (O_313,N_12701,N_14262);
nand UO_314 (O_314,N_13395,N_12421);
or UO_315 (O_315,N_12147,N_13442);
xnor UO_316 (O_316,N_12864,N_13549);
nor UO_317 (O_317,N_14207,N_13822);
and UO_318 (O_318,N_13832,N_12343);
nor UO_319 (O_319,N_12009,N_12811);
nor UO_320 (O_320,N_12150,N_12886);
or UO_321 (O_321,N_14099,N_12552);
nor UO_322 (O_322,N_12957,N_12137);
nor UO_323 (O_323,N_13275,N_14264);
nand UO_324 (O_324,N_12518,N_13349);
or UO_325 (O_325,N_14003,N_13787);
xor UO_326 (O_326,N_13059,N_14325);
or UO_327 (O_327,N_13130,N_14561);
nor UO_328 (O_328,N_13714,N_12817);
and UO_329 (O_329,N_13976,N_13413);
and UO_330 (O_330,N_12437,N_14612);
nor UO_331 (O_331,N_13167,N_13757);
nand UO_332 (O_332,N_13843,N_14069);
nand UO_333 (O_333,N_14029,N_14575);
nor UO_334 (O_334,N_12063,N_14138);
nor UO_335 (O_335,N_13060,N_14828);
and UO_336 (O_336,N_14405,N_14292);
and UO_337 (O_337,N_13534,N_13955);
and UO_338 (O_338,N_14322,N_12451);
nand UO_339 (O_339,N_12596,N_12167);
nand UO_340 (O_340,N_13801,N_12399);
nor UO_341 (O_341,N_14755,N_14411);
nand UO_342 (O_342,N_12528,N_12115);
nand UO_343 (O_343,N_13752,N_13380);
xor UO_344 (O_344,N_14278,N_12395);
nand UO_345 (O_345,N_12219,N_14112);
xor UO_346 (O_346,N_13790,N_13956);
xnor UO_347 (O_347,N_13495,N_12633);
or UO_348 (O_348,N_13509,N_12648);
nor UO_349 (O_349,N_14291,N_13184);
nor UO_350 (O_350,N_14815,N_12064);
nor UO_351 (O_351,N_12526,N_12958);
and UO_352 (O_352,N_13369,N_14166);
or UO_353 (O_353,N_14772,N_13240);
nor UO_354 (O_354,N_14539,N_12590);
or UO_355 (O_355,N_14025,N_13233);
nand UO_356 (O_356,N_13341,N_12933);
nand UO_357 (O_357,N_14345,N_13697);
nor UO_358 (O_358,N_14263,N_14413);
xor UO_359 (O_359,N_13823,N_12911);
nand UO_360 (O_360,N_13933,N_13719);
or UO_361 (O_361,N_13107,N_13093);
or UO_362 (O_362,N_13465,N_14705);
and UO_363 (O_363,N_14997,N_13157);
nor UO_364 (O_364,N_13461,N_14060);
and UO_365 (O_365,N_13125,N_14785);
nand UO_366 (O_366,N_14986,N_14799);
nand UO_367 (O_367,N_13187,N_14672);
nor UO_368 (O_368,N_13132,N_14818);
nor UO_369 (O_369,N_13692,N_12971);
xnor UO_370 (O_370,N_13197,N_14858);
nand UO_371 (O_371,N_12850,N_14122);
xnor UO_372 (O_372,N_13981,N_12419);
xor UO_373 (O_373,N_14732,N_14260);
nor UO_374 (O_374,N_12116,N_12747);
xnor UO_375 (O_375,N_13984,N_14055);
nand UO_376 (O_376,N_13401,N_12426);
and UO_377 (O_377,N_12732,N_13083);
xor UO_378 (O_378,N_14420,N_13767);
nor UO_379 (O_379,N_12094,N_13170);
nand UO_380 (O_380,N_12579,N_14589);
and UO_381 (O_381,N_14305,N_12523);
nor UO_382 (O_382,N_14093,N_12107);
nand UO_383 (O_383,N_13760,N_12962);
and UO_384 (O_384,N_12936,N_13718);
nor UO_385 (O_385,N_14326,N_14136);
and UO_386 (O_386,N_13057,N_13740);
or UO_387 (O_387,N_13906,N_12288);
xor UO_388 (O_388,N_14641,N_14275);
or UO_389 (O_389,N_12443,N_14041);
xor UO_390 (O_390,N_14720,N_13026);
xor UO_391 (O_391,N_13930,N_12882);
and UO_392 (O_392,N_14105,N_14614);
nor UO_393 (O_393,N_14979,N_12194);
nand UO_394 (O_394,N_13247,N_12338);
nor UO_395 (O_395,N_13591,N_13755);
nor UO_396 (O_396,N_14636,N_12506);
nand UO_397 (O_397,N_12509,N_13756);
and UO_398 (O_398,N_13547,N_12717);
and UO_399 (O_399,N_12315,N_12915);
and UO_400 (O_400,N_14065,N_14902);
nor UO_401 (O_401,N_13484,N_13877);
nand UO_402 (O_402,N_12142,N_12401);
xnor UO_403 (O_403,N_13517,N_13673);
nor UO_404 (O_404,N_12408,N_13081);
nor UO_405 (O_405,N_14261,N_14566);
or UO_406 (O_406,N_13211,N_13510);
and UO_407 (O_407,N_14952,N_12510);
nor UO_408 (O_408,N_13959,N_14376);
xnor UO_409 (O_409,N_12715,N_13274);
and UO_410 (O_410,N_14267,N_13315);
xnor UO_411 (O_411,N_12457,N_14595);
or UO_412 (O_412,N_13646,N_14174);
xor UO_413 (O_413,N_12672,N_13538);
xor UO_414 (O_414,N_13280,N_14165);
or UO_415 (O_415,N_13219,N_12370);
and UO_416 (O_416,N_14843,N_12547);
xor UO_417 (O_417,N_13848,N_12974);
or UO_418 (O_418,N_14703,N_14341);
nand UO_419 (O_419,N_12512,N_12440);
or UO_420 (O_420,N_12594,N_12880);
nand UO_421 (O_421,N_14373,N_12930);
nand UO_422 (O_422,N_13204,N_14977);
nand UO_423 (O_423,N_13232,N_12876);
nor UO_424 (O_424,N_12471,N_14496);
xnor UO_425 (O_425,N_12372,N_14307);
nand UO_426 (O_426,N_14331,N_14983);
xnor UO_427 (O_427,N_14051,N_13794);
xor UO_428 (O_428,N_13543,N_12308);
or UO_429 (O_429,N_12255,N_14010);
xor UO_430 (O_430,N_13554,N_12599);
xor UO_431 (O_431,N_13879,N_12346);
xor UO_432 (O_432,N_12283,N_12765);
nor UO_433 (O_433,N_14457,N_12422);
xnor UO_434 (O_434,N_13159,N_13565);
xnor UO_435 (O_435,N_13541,N_13186);
nand UO_436 (O_436,N_13272,N_14700);
or UO_437 (O_437,N_14499,N_12151);
nand UO_438 (O_438,N_14214,N_13713);
xor UO_439 (O_439,N_13835,N_13947);
nand UO_440 (O_440,N_14627,N_14932);
nand UO_441 (O_441,N_13526,N_12631);
nor UO_442 (O_442,N_14153,N_12425);
nor UO_443 (O_443,N_14628,N_13152);
nor UO_444 (O_444,N_12830,N_12867);
nand UO_445 (O_445,N_13452,N_12197);
xnor UO_446 (O_446,N_14753,N_12797);
nor UO_447 (O_447,N_13678,N_14768);
nand UO_448 (O_448,N_12977,N_13635);
or UO_449 (O_449,N_13440,N_14468);
nand UO_450 (O_450,N_14635,N_14493);
xnor UO_451 (O_451,N_12312,N_12804);
nand UO_452 (O_452,N_12985,N_12527);
nand UO_453 (O_453,N_12663,N_13568);
nor UO_454 (O_454,N_13319,N_13683);
nand UO_455 (O_455,N_13831,N_14330);
and UO_456 (O_456,N_14893,N_14505);
nand UO_457 (O_457,N_13542,N_13007);
nand UO_458 (O_458,N_14358,N_14287);
or UO_459 (O_459,N_13001,N_13163);
and UO_460 (O_460,N_12418,N_13171);
or UO_461 (O_461,N_12230,N_13698);
xor UO_462 (O_462,N_14936,N_14431);
xnor UO_463 (O_463,N_13467,N_12770);
and UO_464 (O_464,N_13903,N_14142);
or UO_465 (O_465,N_12560,N_13501);
nand UO_466 (O_466,N_12473,N_14362);
and UO_467 (O_467,N_14102,N_13720);
and UO_468 (O_468,N_14794,N_13177);
and UO_469 (O_469,N_13995,N_13574);
or UO_470 (O_470,N_12271,N_14619);
nor UO_471 (O_471,N_12600,N_13737);
and UO_472 (O_472,N_14494,N_13098);
or UO_473 (O_473,N_14147,N_12483);
xor UO_474 (O_474,N_14803,N_13588);
nand UO_475 (O_475,N_14929,N_12272);
nand UO_476 (O_476,N_14250,N_12098);
nor UO_477 (O_477,N_12365,N_12187);
nor UO_478 (O_478,N_13596,N_13268);
nor UO_479 (O_479,N_13601,N_13470);
and UO_480 (O_480,N_12763,N_12320);
nor UO_481 (O_481,N_12025,N_14559);
and UO_482 (O_482,N_12409,N_14583);
or UO_483 (O_483,N_14107,N_13257);
and UO_484 (O_484,N_14175,N_14934);
nor UO_485 (O_485,N_12837,N_14309);
xor UO_486 (O_486,N_14255,N_13154);
nand UO_487 (O_487,N_13352,N_14108);
and UO_488 (O_488,N_13608,N_12113);
and UO_489 (O_489,N_12758,N_14958);
nor UO_490 (O_490,N_13853,N_14877);
nand UO_491 (O_491,N_13788,N_12352);
nand UO_492 (O_492,N_12250,N_12163);
xor UO_493 (O_493,N_12575,N_12790);
or UO_494 (O_494,N_13746,N_13558);
nand UO_495 (O_495,N_14766,N_13656);
and UO_496 (O_496,N_13251,N_13750);
or UO_497 (O_497,N_12313,N_12924);
nand UO_498 (O_498,N_12400,N_12714);
nor UO_499 (O_499,N_14469,N_12177);
nor UO_500 (O_500,N_12683,N_14313);
or UO_501 (O_501,N_13663,N_14585);
xnor UO_502 (O_502,N_13102,N_13575);
nand UO_503 (O_503,N_13084,N_13405);
nor UO_504 (O_504,N_13003,N_13045);
xor UO_505 (O_505,N_12679,N_13842);
nor UO_506 (O_506,N_14749,N_14835);
nand UO_507 (O_507,N_12966,N_13284);
and UO_508 (O_508,N_12903,N_13996);
xor UO_509 (O_509,N_14912,N_14012);
or UO_510 (O_510,N_14097,N_12606);
nand UO_511 (O_511,N_13642,N_14208);
or UO_512 (O_512,N_14597,N_13881);
nand UO_513 (O_513,N_13188,N_14546);
nor UO_514 (O_514,N_14052,N_12027);
nand UO_515 (O_515,N_13336,N_14126);
nor UO_516 (O_516,N_14075,N_13028);
xor UO_517 (O_517,N_14687,N_14409);
and UO_518 (O_518,N_13897,N_12783);
nor UO_519 (O_519,N_14962,N_14368);
xor UO_520 (O_520,N_12262,N_14395);
and UO_521 (O_521,N_13784,N_14913);
and UO_522 (O_522,N_12030,N_13020);
and UO_523 (O_523,N_12666,N_14911);
xnor UO_524 (O_524,N_12669,N_12202);
and UO_525 (O_525,N_14131,N_14447);
nor UO_526 (O_526,N_13455,N_13560);
xor UO_527 (O_527,N_13221,N_13016);
xnor UO_528 (O_528,N_14118,N_13669);
nand UO_529 (O_529,N_13476,N_13650);
or UO_530 (O_530,N_12028,N_14149);
xor UO_531 (O_531,N_12815,N_14564);
or UO_532 (O_532,N_12228,N_13998);
xor UO_533 (O_533,N_12940,N_14370);
nand UO_534 (O_534,N_14603,N_13667);
or UO_535 (O_535,N_14731,N_12929);
and UO_536 (O_536,N_12780,N_14042);
or UO_537 (O_537,N_13039,N_14920);
and UO_538 (O_538,N_14555,N_14068);
nor UO_539 (O_539,N_12037,N_14823);
or UO_540 (O_540,N_13753,N_14950);
nand UO_541 (O_541,N_14430,N_12777);
or UO_542 (O_542,N_12245,N_14229);
and UO_543 (O_543,N_14437,N_12470);
and UO_544 (O_544,N_12508,N_13438);
nor UO_545 (O_545,N_14295,N_14503);
xor UO_546 (O_546,N_14498,N_14196);
xor UO_547 (O_547,N_13397,N_13585);
nor UO_548 (O_548,N_12155,N_14819);
or UO_549 (O_549,N_14542,N_13408);
nor UO_550 (O_550,N_13439,N_13023);
xor UO_551 (O_551,N_14971,N_12361);
nand UO_552 (O_552,N_13111,N_13485);
xnor UO_553 (O_553,N_14332,N_13231);
or UO_554 (O_554,N_12431,N_12682);
and UO_555 (O_555,N_13192,N_12501);
nor UO_556 (O_556,N_13131,N_13255);
nand UO_557 (O_557,N_14891,N_12000);
xor UO_558 (O_558,N_13138,N_13024);
nor UO_559 (O_559,N_12897,N_12953);
xor UO_560 (O_560,N_14714,N_12848);
and UO_561 (O_561,N_12318,N_12175);
xnor UO_562 (O_562,N_12619,N_12914);
nand UO_563 (O_563,N_13085,N_14961);
xnor UO_564 (O_564,N_12466,N_12222);
nand UO_565 (O_565,N_12143,N_14177);
xnor UO_566 (O_566,N_12467,N_14963);
and UO_567 (O_567,N_12289,N_13441);
and UO_568 (O_568,N_14246,N_13258);
or UO_569 (O_569,N_12438,N_12720);
nand UO_570 (O_570,N_12238,N_14556);
nor UO_571 (O_571,N_13926,N_12153);
or UO_572 (O_572,N_12521,N_14547);
nor UO_573 (O_573,N_12587,N_14683);
or UO_574 (O_574,N_14218,N_12908);
nand UO_575 (O_575,N_13365,N_12691);
xor UO_576 (O_576,N_12843,N_14078);
nand UO_577 (O_577,N_13042,N_14689);
or UO_578 (O_578,N_12563,N_13893);
or UO_579 (O_579,N_14056,N_14299);
nand UO_580 (O_580,N_14201,N_12716);
or UO_581 (O_581,N_12515,N_12812);
nand UO_582 (O_582,N_12178,N_13489);
nor UO_583 (O_583,N_13572,N_12364);
nor UO_584 (O_584,N_12926,N_13726);
xor UO_585 (O_585,N_13849,N_12844);
xnor UO_586 (O_586,N_14702,N_12543);
and UO_587 (O_587,N_12712,N_13844);
nor UO_588 (O_588,N_13226,N_12826);
or UO_589 (O_589,N_12574,N_12907);
and UO_590 (O_590,N_14084,N_12196);
and UO_591 (O_591,N_13374,N_12173);
nor UO_592 (O_592,N_12854,N_14892);
nor UO_593 (O_593,N_13518,N_14862);
xnor UO_594 (O_594,N_13813,N_14923);
nand UO_595 (O_595,N_12375,N_13428);
and UO_596 (O_596,N_12183,N_14005);
nor UO_597 (O_597,N_13350,N_13320);
and UO_598 (O_598,N_13396,N_12148);
or UO_599 (O_599,N_14764,N_14281);
nand UO_600 (O_600,N_14381,N_14728);
xor UO_601 (O_601,N_12124,N_12045);
or UO_602 (O_602,N_13447,N_14115);
nor UO_603 (O_603,N_14639,N_13985);
and UO_604 (O_604,N_13776,N_14511);
nor UO_605 (O_605,N_12309,N_13423);
or UO_606 (O_606,N_13721,N_12065);
and UO_607 (O_607,N_14535,N_12293);
nand UO_608 (O_608,N_13473,N_14477);
and UO_609 (O_609,N_13878,N_14624);
nor UO_610 (O_610,N_12710,N_14928);
or UO_611 (O_611,N_12593,N_13624);
nor UO_612 (O_612,N_12625,N_14707);
nand UO_613 (O_613,N_12092,N_14652);
nand UO_614 (O_614,N_14579,N_12664);
xnor UO_615 (O_615,N_13691,N_12111);
and UO_616 (O_616,N_12637,N_14501);
nand UO_617 (O_617,N_14664,N_14141);
nand UO_618 (O_618,N_13777,N_13627);
nor UO_619 (O_619,N_14015,N_12468);
xor UO_620 (O_620,N_13837,N_13814);
xor UO_621 (O_621,N_14533,N_13715);
xnor UO_622 (O_622,N_12558,N_14334);
nor UO_623 (O_623,N_14327,N_14677);
and UO_624 (O_624,N_12380,N_14993);
nand UO_625 (O_625,N_12901,N_12251);
or UO_626 (O_626,N_12822,N_14199);
nor UO_627 (O_627,N_14917,N_13230);
xor UO_628 (O_628,N_14185,N_12890);
nand UO_629 (O_629,N_12007,N_13322);
xnor UO_630 (O_630,N_12411,N_13420);
nand UO_631 (O_631,N_12961,N_13965);
and UO_632 (O_632,N_13189,N_14626);
nor UO_633 (O_633,N_14663,N_14066);
nor UO_634 (O_634,N_12049,N_13524);
nor UO_635 (O_635,N_12654,N_12615);
or UO_636 (O_636,N_13142,N_14792);
and UO_637 (O_637,N_13012,N_12950);
xor UO_638 (O_638,N_12295,N_14238);
nor UO_639 (O_639,N_14863,N_12090);
or UO_640 (O_640,N_13762,N_12052);
xor UO_641 (O_641,N_13270,N_14321);
xor UO_642 (O_642,N_12948,N_13421);
nand UO_643 (O_643,N_13414,N_13816);
or UO_644 (O_644,N_12978,N_12741);
nor UO_645 (O_645,N_14694,N_12477);
nand UO_646 (O_646,N_14591,N_14082);
xor UO_647 (O_647,N_13957,N_14446);
or UO_648 (O_648,N_13519,N_14209);
nand UO_649 (O_649,N_12580,N_14735);
or UO_650 (O_650,N_14007,N_13326);
nand UO_651 (O_651,N_13314,N_14502);
nand UO_652 (O_652,N_13248,N_12764);
and UO_653 (O_653,N_14357,N_14421);
or UO_654 (O_654,N_12572,N_12551);
nor UO_655 (O_655,N_12134,N_13583);
nand UO_656 (O_656,N_14623,N_14953);
xnor UO_657 (O_657,N_14933,N_12494);
nor UO_658 (O_658,N_13613,N_14340);
nand UO_659 (O_659,N_14532,N_14784);
or UO_660 (O_660,N_14964,N_13078);
nor UO_661 (O_661,N_13679,N_14106);
xor UO_662 (O_662,N_13939,N_14530);
or UO_663 (O_663,N_13390,N_14221);
xor UO_664 (O_664,N_12232,N_13654);
xnor UO_665 (O_665,N_14486,N_14124);
and UO_666 (O_666,N_14164,N_14618);
nand UO_667 (O_667,N_14026,N_14582);
and UO_668 (O_668,N_13448,N_12442);
xnor UO_669 (O_669,N_13317,N_12805);
nand UO_670 (O_670,N_14049,N_12559);
and UO_671 (O_671,N_12789,N_12428);
nor UO_672 (O_672,N_14465,N_12612);
nand UO_673 (O_673,N_14888,N_13778);
and UO_674 (O_674,N_13640,N_13151);
or UO_675 (O_675,N_13564,N_12900);
nand UO_676 (O_676,N_14414,N_13545);
nor UO_677 (O_677,N_12449,N_12472);
and UO_678 (O_678,N_12059,N_12602);
or UO_679 (O_679,N_14460,N_14850);
xor UO_680 (O_680,N_12856,N_14000);
nand UO_681 (O_681,N_12989,N_13741);
and UO_682 (O_682,N_13546,N_13463);
or UO_683 (O_683,N_13690,N_14695);
nand UO_684 (O_684,N_14302,N_12441);
nand UO_685 (O_685,N_14244,N_13969);
xnor UO_686 (O_686,N_13471,N_12371);
and UO_687 (O_687,N_13136,N_13015);
xnor UO_688 (O_688,N_12731,N_12405);
and UO_689 (O_689,N_12709,N_13190);
xnor UO_690 (O_690,N_14311,N_12201);
and UO_691 (O_691,N_12931,N_12992);
nor UO_692 (O_692,N_13818,N_13095);
xnor UO_693 (O_693,N_13340,N_13514);
xnor UO_694 (O_694,N_12388,N_12146);
xor UO_695 (O_695,N_14076,N_12818);
xnor UO_696 (O_696,N_13196,N_13122);
nor UO_697 (O_697,N_14730,N_14173);
xor UO_698 (O_698,N_12479,N_12430);
or UO_699 (O_699,N_12358,N_14490);
or UO_700 (O_700,N_14223,N_13259);
and UO_701 (O_701,N_14320,N_12761);
nand UO_702 (O_702,N_13345,N_13666);
xnor UO_703 (O_703,N_12321,N_13792);
nor UO_704 (O_704,N_12986,N_13499);
nand UO_705 (O_705,N_13368,N_14711);
xor UO_706 (O_706,N_12357,N_12999);
nand UO_707 (O_707,N_13978,N_12070);
xnor UO_708 (O_708,N_14773,N_12360);
or UO_709 (O_709,N_13594,N_12891);
nor UO_710 (O_710,N_12684,N_14243);
xor UO_711 (O_711,N_14708,N_13064);
nand UO_712 (O_712,N_12791,N_14882);
and UO_713 (O_713,N_12485,N_12645);
xnor UO_714 (O_714,N_13649,N_14840);
nand UO_715 (O_715,N_13552,N_12218);
xor UO_716 (O_716,N_14103,N_14514);
xor UO_717 (O_717,N_12841,N_13490);
nor UO_718 (O_718,N_12207,N_13764);
and UO_719 (O_719,N_14210,N_14567);
and UO_720 (O_720,N_14167,N_14765);
and UO_721 (O_721,N_14148,N_14211);
and UO_722 (O_722,N_13174,N_14363);
xnor UO_723 (O_723,N_14425,N_14328);
xnor UO_724 (O_724,N_12870,N_13830);
or UO_725 (O_725,N_13382,N_12598);
nand UO_726 (O_726,N_14528,N_13072);
nand UO_727 (O_727,N_14422,N_13860);
nor UO_728 (O_728,N_13631,N_14632);
and UO_729 (O_729,N_14922,N_14654);
and UO_730 (O_730,N_12852,N_13567);
and UO_731 (O_731,N_14517,N_14467);
and UO_732 (O_732,N_12835,N_13992);
or UO_733 (O_733,N_12540,N_14873);
nand UO_734 (O_734,N_12299,N_13701);
nand UO_735 (O_735,N_12123,N_13889);
xnor UO_736 (O_736,N_12748,N_12888);
nand UO_737 (O_737,N_13411,N_13680);
nor UO_738 (O_738,N_13327,N_13207);
nor UO_739 (O_739,N_12374,N_12248);
xnor UO_740 (O_740,N_12514,N_14508);
xor UO_741 (O_741,N_14061,N_13324);
nand UO_742 (O_742,N_12609,N_14691);
or UO_743 (O_743,N_14587,N_14830);
nor UO_744 (O_744,N_12242,N_12447);
xor UO_745 (O_745,N_13427,N_13236);
nor UO_746 (O_746,N_14157,N_12184);
nand UO_747 (O_747,N_14163,N_14043);
nand UO_748 (O_748,N_12500,N_12135);
and UO_749 (O_749,N_14253,N_14904);
xnor UO_750 (O_750,N_12385,N_13256);
nand UO_751 (O_751,N_14745,N_13706);
and UO_752 (O_752,N_12268,N_12636);
or UO_753 (O_753,N_13791,N_14824);
xor UO_754 (O_754,N_12317,N_13050);
nor UO_755 (O_755,N_14019,N_12249);
nor UO_756 (O_756,N_12519,N_12567);
or UO_757 (O_757,N_12820,N_13977);
xnor UO_758 (O_758,N_14155,N_12476);
and UO_759 (O_759,N_12601,N_14686);
or UO_760 (O_760,N_13953,N_13951);
or UO_761 (O_761,N_12493,N_14389);
xor UO_762 (O_762,N_13134,N_12993);
nand UO_763 (O_763,N_12605,N_12808);
nor UO_764 (O_764,N_12708,N_12681);
and UO_765 (O_765,N_14719,N_13293);
xnor UO_766 (O_766,N_12077,N_13605);
nand UO_767 (O_767,N_12089,N_12603);
xor UO_768 (O_768,N_12080,N_13652);
xnor UO_769 (O_769,N_12846,N_13841);
xor UO_770 (O_770,N_14293,N_13307);
xnor UO_771 (O_771,N_12736,N_12697);
or UO_772 (O_772,N_14116,N_13884);
nand UO_773 (O_773,N_13052,N_12744);
and UO_774 (O_774,N_14359,N_13562);
nand UO_775 (O_775,N_13041,N_12502);
xor UO_776 (O_776,N_14416,N_13749);
nor UO_777 (O_777,N_12093,N_14544);
and UO_778 (O_778,N_14870,N_14642);
and UO_779 (O_779,N_13744,N_13040);
xnor UO_780 (O_780,N_12074,N_12016);
nor UO_781 (O_781,N_12533,N_13331);
nor UO_782 (O_782,N_12639,N_12145);
xor UO_783 (O_783,N_13782,N_14057);
nor UO_784 (O_784,N_12516,N_13357);
xor UO_785 (O_785,N_14162,N_14466);
xnor UO_786 (O_786,N_14252,N_13018);
or UO_787 (O_787,N_14306,N_14833);
xnor UO_788 (O_788,N_14609,N_12832);
and UO_789 (O_789,N_12095,N_13165);
xor UO_790 (O_790,N_13668,N_14924);
nand UO_791 (O_791,N_14569,N_12982);
nor UO_792 (O_792,N_13035,N_12569);
nor UO_793 (O_793,N_12047,N_14855);
or UO_794 (O_794,N_13734,N_14369);
nor UO_795 (O_795,N_14796,N_14991);
xnor UO_796 (O_796,N_12622,N_12749);
nor UO_797 (O_797,N_13653,N_12008);
nor UO_798 (O_798,N_13301,N_13090);
and UO_799 (O_799,N_12129,N_12101);
nor UO_800 (O_800,N_12022,N_14622);
nand UO_801 (O_801,N_12589,N_14607);
nor UO_802 (O_802,N_13645,N_14215);
and UO_803 (O_803,N_13445,N_12062);
and UO_804 (O_804,N_14715,N_12258);
or UO_805 (O_805,N_13569,N_14452);
or UO_806 (O_806,N_13934,N_13308);
nand UO_807 (O_807,N_12784,N_12191);
nor UO_808 (O_808,N_13183,N_14757);
nor UO_809 (O_809,N_12433,N_12858);
and UO_810 (O_810,N_14854,N_14941);
nor UO_811 (O_811,N_13245,N_14443);
and UO_812 (O_812,N_12524,N_14909);
nand UO_813 (O_813,N_13971,N_13892);
nand UO_814 (O_814,N_13325,N_13488);
nor UO_815 (O_815,N_13676,N_13071);
and UO_816 (O_816,N_14195,N_13923);
nor UO_817 (O_817,N_13941,N_13218);
xor UO_818 (O_818,N_13335,N_13145);
or UO_819 (O_819,N_12549,N_12038);
nor UO_820 (O_820,N_14679,N_13637);
nand UO_821 (O_821,N_14834,N_13209);
xor UO_822 (O_822,N_13863,N_12208);
and UO_823 (O_823,N_12916,N_12475);
xnor UO_824 (O_824,N_12076,N_12387);
xor UO_825 (O_825,N_13429,N_12678);
nor UO_826 (O_826,N_12019,N_12772);
or UO_827 (O_827,N_14442,N_12542);
and UO_828 (O_828,N_13539,N_13323);
nand UO_829 (O_829,N_12036,N_13660);
or UO_830 (O_830,N_14523,N_13508);
xor UO_831 (O_831,N_13505,N_14698);
or UO_832 (O_832,N_13377,N_13597);
nor UO_833 (O_833,N_12742,N_13087);
or UO_834 (O_834,N_12081,N_12539);
xnor UO_835 (O_835,N_13089,N_14176);
nor UO_836 (O_836,N_13885,N_13305);
nand UO_837 (O_837,N_13817,N_14388);
or UO_838 (O_838,N_12023,N_14178);
nand UO_839 (O_839,N_12461,N_13876);
xnor UO_840 (O_840,N_13682,N_14478);
xor UO_841 (O_841,N_14294,N_14009);
and UO_842 (O_842,N_12072,N_13774);
xnor UO_843 (O_843,N_13437,N_13571);
nor UO_844 (O_844,N_12531,N_14071);
xor UO_845 (O_845,N_14127,N_13337);
or UO_846 (O_846,N_14864,N_12237);
nor UO_847 (O_847,N_13589,N_12005);
xor UO_848 (O_848,N_12641,N_12737);
nor UO_849 (O_849,N_14551,N_14289);
xor UO_850 (O_850,N_14161,N_13899);
and UO_851 (O_851,N_13112,N_13852);
and UO_852 (O_852,N_14203,N_14033);
and UO_853 (O_853,N_12203,N_14743);
nor UO_854 (O_854,N_14419,N_13182);
nor UO_855 (O_855,N_12597,N_14394);
or UO_856 (O_856,N_12198,N_12021);
and UO_857 (O_857,N_14364,N_14890);
nor UO_858 (O_858,N_12877,N_12270);
or UO_859 (O_859,N_12226,N_14734);
or UO_860 (O_860,N_13530,N_12827);
nor UO_861 (O_861,N_14856,N_14500);
and UO_862 (O_862,N_14807,N_13766);
xor UO_863 (O_863,N_13295,N_13056);
xor UO_864 (O_864,N_14640,N_12795);
nand UO_865 (O_865,N_12952,N_12286);
nand UO_866 (O_866,N_14095,N_13775);
nand UO_867 (O_867,N_14407,N_12166);
or UO_868 (O_868,N_14098,N_14770);
and UO_869 (O_869,N_12109,N_12348);
xor UO_870 (O_870,N_12800,N_14192);
or UO_871 (O_871,N_13063,N_13481);
xnor UO_872 (O_872,N_14727,N_14085);
nand UO_873 (O_873,N_14296,N_13051);
and UO_874 (O_874,N_13810,N_14424);
nand UO_875 (O_875,N_12190,N_12487);
or UO_876 (O_876,N_14586,N_13161);
or UO_877 (O_877,N_12875,N_12486);
xor UO_878 (O_878,N_13604,N_13386);
xnor UO_879 (O_879,N_12427,N_12967);
or UO_880 (O_880,N_13372,N_12066);
nor UO_881 (O_881,N_14721,N_14655);
nand UO_882 (O_882,N_13819,N_14242);
xor UO_883 (O_883,N_14352,N_12263);
or UO_884 (O_884,N_14132,N_14608);
xor UO_885 (O_885,N_14239,N_14954);
xor UO_886 (O_886,N_14506,N_12171);
nand UO_887 (O_887,N_13987,N_13149);
xnor UO_888 (O_888,N_13858,N_12265);
and UO_889 (O_889,N_12668,N_13262);
xor UO_890 (O_890,N_13962,N_13763);
nand UO_891 (O_891,N_12503,N_14811);
and UO_892 (O_892,N_13477,N_12556);
xor UO_893 (O_893,N_12463,N_14284);
and UO_894 (O_894,N_12665,N_12048);
xor UO_895 (O_895,N_13948,N_14526);
xnor UO_896 (O_896,N_13786,N_12923);
xnor UO_897 (O_897,N_14967,N_13294);
or UO_898 (O_898,N_13216,N_13871);
nor UO_899 (O_899,N_13590,N_14485);
and UO_900 (O_900,N_14565,N_14908);
nor UO_901 (O_901,N_14073,N_14842);
xnor UO_902 (O_902,N_13246,N_12061);
nor UO_903 (O_903,N_12136,N_13283);
or UO_904 (O_904,N_14461,N_12046);
or UO_905 (O_905,N_13686,N_14070);
nor UO_906 (O_906,N_14383,N_13945);
and UO_907 (O_907,N_12869,N_13457);
nand UO_908 (O_908,N_12842,N_14522);
nor UO_909 (O_909,N_14088,N_13770);
nand UO_910 (O_910,N_12379,N_14236);
nand UO_911 (O_911,N_13882,N_12674);
or UO_912 (O_912,N_14435,N_13496);
and UO_913 (O_913,N_13296,N_13745);
nand UO_914 (O_914,N_13469,N_13533);
and UO_915 (O_915,N_14367,N_13961);
or UO_916 (O_916,N_14254,N_13553);
nor UO_917 (O_917,N_12694,N_13399);
nand UO_918 (O_918,N_14880,N_12845);
or UO_919 (O_919,N_14406,N_12125);
and UO_920 (O_920,N_12608,N_14959);
or UO_921 (O_921,N_12534,N_14876);
nor UO_922 (O_922,N_14816,N_13902);
or UO_923 (O_923,N_14802,N_13176);
and UO_924 (O_924,N_12157,N_13214);
nor UO_925 (O_925,N_14456,N_13581);
xor UO_926 (O_926,N_13910,N_14247);
nor UO_927 (O_927,N_13952,N_14031);
xnor UO_928 (O_928,N_13938,N_13304);
or UO_929 (O_929,N_12140,N_13068);
and UO_930 (O_930,N_13511,N_13038);
nor UO_931 (O_931,N_13907,N_13963);
nand UO_932 (O_932,N_12158,N_14557);
xnor UO_933 (O_933,N_12944,N_14900);
nand UO_934 (O_934,N_14481,N_13993);
xor UO_935 (O_935,N_13113,N_14212);
and UO_936 (O_936,N_12229,N_14121);
or UO_937 (O_937,N_14895,N_13960);
nor UO_938 (O_938,N_13556,N_14775);
xnor UO_939 (O_939,N_14659,N_14791);
nand UO_940 (O_940,N_12673,N_13370);
and UO_941 (O_941,N_13332,N_13334);
nand UO_942 (O_942,N_12341,N_14987);
xnor UO_943 (O_943,N_13811,N_13392);
nand UO_944 (O_944,N_12314,N_13925);
or UO_945 (O_945,N_12499,N_12662);
or UO_946 (O_946,N_14810,N_14397);
nor UO_947 (O_947,N_14935,N_14617);
and UO_948 (O_948,N_14910,N_14030);
or UO_949 (O_949,N_14335,N_13073);
xnor UO_950 (O_950,N_14723,N_14319);
nand UO_951 (O_951,N_13515,N_13486);
or UO_952 (O_952,N_14650,N_13615);
nor UO_953 (O_953,N_13688,N_14906);
xor UO_954 (O_954,N_12079,N_13460);
nor UO_955 (O_955,N_14143,N_14439);
xor UO_956 (O_956,N_13609,N_13079);
and UO_957 (O_957,N_13133,N_12909);
nor UO_958 (O_958,N_12276,N_13114);
xor UO_959 (O_959,N_13005,N_12264);
nor UO_960 (O_960,N_13158,N_14540);
nor UO_961 (O_961,N_12834,N_12656);
and UO_962 (O_962,N_12344,N_12991);
nand UO_963 (O_963,N_12905,N_14804);
or UO_964 (O_964,N_14577,N_12234);
nor UO_965 (O_965,N_13241,N_14762);
and UO_966 (O_966,N_12159,N_14379);
nor UO_967 (O_967,N_13181,N_14463);
nor UO_968 (O_968,N_12404,N_12275);
xor UO_969 (O_969,N_14930,N_12075);
xor UO_970 (O_970,N_12188,N_13806);
nor UO_971 (O_971,N_13195,N_12651);
or UO_972 (O_972,N_12965,N_12459);
nor UO_973 (O_973,N_12910,N_13633);
xor UO_974 (O_974,N_14662,N_14288);
or UO_975 (O_975,N_12536,N_12573);
nor UO_976 (O_976,N_12809,N_14754);
or UO_977 (O_977,N_12363,N_14343);
nor UO_978 (O_978,N_12990,N_13436);
and UO_979 (O_979,N_12511,N_13032);
and UO_980 (O_980,N_14039,N_14574);
or UO_981 (O_981,N_12067,N_12239);
xnor UO_982 (O_982,N_14123,N_13940);
or UO_983 (O_983,N_13424,N_14193);
nand UO_984 (O_984,N_12692,N_13303);
and UO_985 (O_985,N_13173,N_14673);
and UO_986 (O_986,N_12450,N_14554);
and UO_987 (O_987,N_13178,N_14371);
or UO_988 (O_988,N_12160,N_12705);
nor UO_989 (O_989,N_13826,N_13037);
and UO_990 (O_990,N_13661,N_14360);
nor UO_991 (O_991,N_14171,N_12711);
or UO_992 (O_992,N_13498,N_13105);
or UO_993 (O_993,N_12621,N_13250);
nand UO_994 (O_994,N_13531,N_13493);
nand UO_995 (O_995,N_12785,N_14947);
or UO_996 (O_996,N_13946,N_14685);
nor UO_997 (O_997,N_12703,N_12721);
and UO_998 (O_998,N_14697,N_12799);
and UO_999 (O_999,N_14901,N_14844);
nor UO_1000 (O_1000,N_14918,N_12771);
or UO_1001 (O_1001,N_13536,N_14300);
and UO_1002 (O_1002,N_14837,N_14832);
nor UO_1003 (O_1003,N_14217,N_14633);
and UO_1004 (O_1004,N_13010,N_13908);
nor UO_1005 (O_1005,N_13747,N_12376);
xnor UO_1006 (O_1006,N_14884,N_13736);
or UO_1007 (O_1007,N_13641,N_13815);
xor UO_1008 (O_1008,N_13106,N_14495);
nor UO_1009 (O_1009,N_14240,N_14448);
xor UO_1010 (O_1010,N_12532,N_13394);
xor UO_1011 (O_1011,N_14998,N_12445);
and UO_1012 (O_1012,N_13118,N_12866);
and UO_1013 (O_1013,N_13472,N_12034);
xor UO_1014 (O_1014,N_12868,N_13062);
xor UO_1015 (O_1015,N_12390,N_12243);
and UO_1016 (O_1016,N_13404,N_14529);
nand UO_1017 (O_1017,N_14487,N_12655);
or UO_1018 (O_1018,N_12448,N_14693);
nor UO_1019 (O_1019,N_13031,N_13419);
nand UO_1020 (O_1020,N_14128,N_13943);
or UO_1021 (O_1021,N_14228,N_13935);
and UO_1022 (O_1022,N_13478,N_14790);
xnor UO_1023 (O_1023,N_14144,N_13723);
xnor UO_1024 (O_1024,N_14744,N_12306);
or UO_1025 (O_1025,N_14593,N_13201);
nand UO_1026 (O_1026,N_12836,N_13918);
or UO_1027 (O_1027,N_13367,N_12302);
or UO_1028 (O_1028,N_13312,N_13870);
nand UO_1029 (O_1029,N_14563,N_14184);
nor UO_1030 (O_1030,N_13127,N_12041);
and UO_1031 (O_1031,N_14342,N_12553);
xor UO_1032 (O_1032,N_13479,N_13354);
or UO_1033 (O_1033,N_14531,N_12752);
or UO_1034 (O_1034,N_13779,N_13913);
and UO_1035 (O_1035,N_13119,N_13611);
nor UO_1036 (O_1036,N_14194,N_13146);
nand UO_1037 (O_1037,N_12627,N_14674);
nor UO_1038 (O_1038,N_13388,N_12628);
nand UO_1039 (O_1039,N_14515,N_12391);
xnor UO_1040 (O_1040,N_13100,N_14216);
nand UO_1041 (O_1041,N_14269,N_13761);
xnor UO_1042 (O_1042,N_14970,N_13343);
nor UO_1043 (O_1043,N_12316,N_12382);
and UO_1044 (O_1044,N_13880,N_12774);
or UO_1045 (O_1045,N_13577,N_14308);
xor UO_1046 (O_1046,N_12667,N_13850);
and UO_1047 (O_1047,N_13561,N_14282);
nand UO_1048 (O_1048,N_12610,N_13169);
xnor UO_1049 (O_1049,N_14256,N_13521);
or UO_1050 (O_1050,N_13217,N_12267);
or UO_1051 (O_1051,N_14024,N_12269);
and UO_1052 (O_1052,N_12857,N_13891);
nor UO_1053 (O_1053,N_14925,N_13048);
or UO_1054 (O_1054,N_12727,N_13916);
nor UO_1055 (O_1055,N_12706,N_13430);
nor UO_1056 (O_1056,N_13685,N_13932);
xnor UO_1057 (O_1057,N_12548,N_12564);
and UO_1058 (O_1058,N_14570,N_14145);
or UO_1059 (O_1059,N_14826,N_13616);
and UO_1060 (O_1060,N_14191,N_14578);
and UO_1061 (O_1061,N_14808,N_13099);
and UO_1062 (O_1062,N_14518,N_13036);
xor UO_1063 (O_1063,N_14601,N_14537);
xor UO_1064 (O_1064,N_14657,N_13454);
or UO_1065 (O_1065,N_14645,N_12429);
nand UO_1066 (O_1066,N_12896,N_12616);
and UO_1067 (O_1067,N_14625,N_12103);
or UO_1068 (O_1068,N_12565,N_13797);
xnor UO_1069 (O_1069,N_13711,N_13168);
nand UO_1070 (O_1070,N_13638,N_12026);
nor UO_1071 (O_1071,N_14946,N_14183);
nor UO_1072 (O_1072,N_12979,N_14464);
nor UO_1073 (O_1073,N_13550,N_14889);
or UO_1074 (O_1074,N_12168,N_14227);
and UO_1075 (O_1075,N_13540,N_13425);
nor UO_1076 (O_1076,N_12304,N_13664);
or UO_1077 (O_1077,N_13657,N_13725);
nor UO_1078 (O_1078,N_12700,N_12413);
and UO_1079 (O_1079,N_13828,N_14429);
or UO_1080 (O_1080,N_12638,N_14455);
xnor UO_1081 (O_1081,N_14317,N_12033);
and UO_1082 (O_1082,N_14616,N_12029);
and UO_1083 (O_1083,N_14170,N_13548);
nor UO_1084 (O_1084,N_13895,N_13739);
xor UO_1085 (O_1085,N_12537,N_12566);
and UO_1086 (O_1086,N_14087,N_14265);
and UO_1087 (O_1087,N_12904,N_13434);
nand UO_1088 (O_1088,N_12044,N_13384);
nand UO_1089 (O_1089,N_12465,N_14610);
xnor UO_1090 (O_1090,N_14568,N_12935);
or UO_1091 (O_1091,N_13586,N_14788);
xor UO_1092 (O_1092,N_12517,N_12729);
and UO_1093 (O_1093,N_13433,N_13728);
or UO_1094 (O_1094,N_14450,N_13580);
and UO_1095 (O_1095,N_13593,N_14483);
and UO_1096 (O_1096,N_14417,N_14690);
or UO_1097 (O_1097,N_12211,N_14198);
nor UO_1098 (O_1098,N_14825,N_14676);
or UO_1099 (O_1099,N_14273,N_13013);
and UO_1100 (O_1100,N_13502,N_14838);
nand UO_1101 (O_1101,N_12332,N_13834);
or UO_1102 (O_1102,N_14666,N_13708);
nand UO_1103 (O_1103,N_14062,N_13287);
nor UO_1104 (O_1104,N_13785,N_12584);
or UO_1105 (O_1105,N_12227,N_12728);
nand UO_1106 (O_1106,N_14534,N_12960);
or UO_1107 (O_1107,N_13527,N_12192);
nor UO_1108 (O_1108,N_12833,N_13621);
nand UO_1109 (O_1109,N_14965,N_12723);
and UO_1110 (O_1110,N_14032,N_12161);
nor UO_1111 (O_1111,N_12849,N_12861);
or UO_1112 (O_1112,N_14782,N_12899);
nand UO_1113 (O_1113,N_13137,N_14915);
nor UO_1114 (O_1114,N_14080,N_14572);
or UO_1115 (O_1115,N_12291,N_14638);
nand UO_1116 (O_1116,N_13929,N_12963);
nand UO_1117 (O_1117,N_13825,N_14489);
or UO_1118 (O_1118,N_14805,N_14763);
or UO_1119 (O_1119,N_13839,N_12252);
and UO_1120 (O_1120,N_14795,N_13047);
xnor UO_1121 (O_1121,N_13869,N_14751);
nor UO_1122 (O_1122,N_12278,N_13512);
and UO_1123 (O_1123,N_14323,N_12902);
and UO_1124 (O_1124,N_12453,N_13820);
or UO_1125 (O_1125,N_14536,N_12632);
nor UO_1126 (O_1126,N_12336,N_13403);
nand UO_1127 (O_1127,N_14139,N_14709);
and UO_1128 (O_1128,N_14034,N_14919);
and UO_1129 (O_1129,N_14374,N_12878);
or UO_1130 (O_1130,N_12829,N_13875);
nor UO_1131 (O_1131,N_14440,N_14665);
or UO_1132 (O_1132,N_13208,N_14202);
or UO_1133 (O_1133,N_13299,N_14432);
xnor UO_1134 (O_1134,N_14054,N_12801);
xor UO_1135 (O_1135,N_13974,N_12416);
nor UO_1136 (O_1136,N_13311,N_14778);
and UO_1137 (O_1137,N_14151,N_12756);
xor UO_1138 (O_1138,N_13222,N_12434);
nand UO_1139 (O_1139,N_12055,N_13410);
and UO_1140 (O_1140,N_14458,N_13618);
and UO_1141 (O_1141,N_13803,N_14867);
and UO_1142 (O_1142,N_13990,N_12873);
nor UO_1143 (O_1143,N_12039,N_12004);
and UO_1144 (O_1144,N_13584,N_12658);
nand UO_1145 (O_1145,N_13898,N_14454);
and UO_1146 (O_1146,N_13393,N_12224);
xnor UO_1147 (O_1147,N_12209,N_14939);
nor UO_1148 (O_1148,N_13735,N_12189);
and UO_1149 (O_1149,N_12825,N_13004);
nand UO_1150 (O_1150,N_14733,N_14316);
nor UO_1151 (O_1151,N_13091,N_14472);
xnor UO_1152 (O_1152,N_12623,N_12831);
xnor UO_1153 (O_1153,N_12661,N_14996);
nor UO_1154 (O_1154,N_12053,N_14739);
and UO_1155 (O_1155,N_13798,N_12676);
nand UO_1156 (O_1156,N_12776,N_14020);
nor UO_1157 (O_1157,N_13972,N_12215);
nor UO_1158 (O_1158,N_13200,N_12392);
and UO_1159 (O_1159,N_12349,N_14670);
nand UO_1160 (O_1160,N_13865,N_14219);
xor UO_1161 (O_1161,N_12925,N_12216);
xnor UO_1162 (O_1162,N_12144,N_12504);
xor UO_1163 (O_1163,N_13213,N_14726);
xnor UO_1164 (O_1164,N_12889,N_14412);
nor UO_1165 (O_1165,N_13344,N_13731);
or UO_1166 (O_1166,N_14945,N_13225);
nand UO_1167 (O_1167,N_14949,N_13046);
nor UO_1168 (O_1168,N_13733,N_14438);
or UO_1169 (O_1169,N_13573,N_12650);
xor UO_1170 (O_1170,N_14423,N_13887);
or UO_1171 (O_1171,N_12529,N_13693);
nor UO_1172 (O_1172,N_12257,N_14868);
nor UO_1173 (O_1173,N_14462,N_13021);
xor UO_1174 (O_1174,N_13227,N_12133);
and UO_1175 (O_1175,N_14814,N_13836);
xor UO_1176 (O_1176,N_14817,N_14470);
or UO_1177 (O_1177,N_14434,N_13215);
nor UO_1178 (O_1178,N_12496,N_12497);
nor UO_1179 (O_1179,N_13487,N_12895);
or UO_1180 (O_1180,N_12972,N_12530);
xnor UO_1181 (O_1181,N_13094,N_14647);
xor UO_1182 (O_1182,N_12217,N_14898);
nand UO_1183 (O_1183,N_14036,N_12290);
nand UO_1184 (O_1184,N_12277,N_12568);
or UO_1185 (O_1185,N_12498,N_13700);
nor UO_1186 (O_1186,N_13153,N_13162);
and UO_1187 (O_1187,N_12006,N_14875);
xor UO_1188 (O_1188,N_12724,N_14197);
or UO_1189 (O_1189,N_12247,N_12718);
xnor UO_1190 (O_1190,N_12310,N_12738);
nand UO_1191 (O_1191,N_14948,N_13432);
or UO_1192 (O_1192,N_12750,N_13563);
or UO_1193 (O_1193,N_14473,N_12644);
or UO_1194 (O_1194,N_13607,N_12949);
nand UO_1195 (O_1195,N_14396,N_14241);
nand UO_1196 (O_1196,N_14857,N_12054);
and UO_1197 (O_1197,N_12464,N_12104);
xnor UO_1198 (O_1198,N_12635,N_13061);
xor UO_1199 (O_1199,N_13053,N_12410);
nor UO_1200 (O_1200,N_13179,N_13845);
xnor UO_1201 (O_1201,N_14600,N_12775);
or UO_1202 (O_1202,N_14044,N_14348);
nor UO_1203 (O_1203,N_13681,N_14276);
or UO_1204 (O_1204,N_14871,N_14899);
or UO_1205 (O_1205,N_14488,N_12646);
and UO_1206 (O_1206,N_13080,N_12544);
and UO_1207 (O_1207,N_12325,N_12576);
nor UO_1208 (O_1208,N_13058,N_13300);
nor UO_1209 (O_1209,N_14759,N_12823);
nor UO_1210 (O_1210,N_14777,N_14047);
xor UO_1211 (O_1211,N_12082,N_14279);
xnor UO_1212 (O_1212,N_13851,N_12959);
nor UO_1213 (O_1213,N_12726,N_12132);
xor UO_1214 (O_1214,N_12469,N_13101);
xnor UO_1215 (O_1215,N_13375,N_14831);
nand UO_1216 (O_1216,N_14310,N_12642);
nor UO_1217 (O_1217,N_14135,N_12819);
and UO_1218 (O_1218,N_12630,N_12127);
or UO_1219 (O_1219,N_12917,N_14257);
nand UO_1220 (O_1220,N_12165,N_14150);
and UO_1221 (O_1221,N_13773,N_13570);
or UO_1222 (O_1222,N_14548,N_13391);
nand UO_1223 (O_1223,N_14741,N_13703);
nand UO_1224 (O_1224,N_12254,N_14436);
nor UO_1225 (O_1225,N_12983,N_12130);
nor UO_1226 (O_1226,N_14750,N_13400);
nand UO_1227 (O_1227,N_12695,N_13494);
xnor UO_1228 (O_1228,N_12762,N_12345);
xnor UO_1229 (O_1229,N_14475,N_12347);
xnor UO_1230 (O_1230,N_12806,N_13937);
and UO_1231 (O_1231,N_14372,N_12614);
nor UO_1232 (O_1232,N_12677,N_14392);
or UO_1233 (O_1233,N_12073,N_14002);
and UO_1234 (O_1234,N_13824,N_13557);
nand UO_1235 (O_1235,N_12214,N_12730);
or UO_1236 (O_1236,N_12657,N_12355);
xor UO_1237 (O_1237,N_12424,N_12687);
nand UO_1238 (O_1238,N_14285,N_14771);
and UO_1239 (O_1239,N_14333,N_13497);
nor UO_1240 (O_1240,N_12883,N_14976);
and UO_1241 (O_1241,N_12322,N_13532);
or UO_1242 (O_1242,N_12342,N_14704);
nand UO_1243 (O_1243,N_14224,N_13034);
or UO_1244 (O_1244,N_12807,N_14839);
nor UO_1245 (O_1245,N_13595,N_12634);
nand UO_1246 (O_1246,N_14512,N_12670);
nand UO_1247 (O_1247,N_14023,N_13077);
or UO_1248 (O_1248,N_14064,N_12407);
nand UO_1249 (O_1249,N_13006,N_12205);
or UO_1250 (O_1250,N_14980,N_14521);
and UO_1251 (O_1251,N_14716,N_14829);
xnor UO_1252 (O_1252,N_14329,N_12987);
or UO_1253 (O_1253,N_12722,N_13914);
nand UO_1254 (O_1254,N_13909,N_14800);
xor UO_1255 (O_1255,N_12490,N_12995);
xor UO_1256 (O_1256,N_13768,N_14119);
xor UO_1257 (O_1257,N_12368,N_14571);
nor UO_1258 (O_1258,N_13827,N_12956);
nand UO_1259 (O_1259,N_12373,N_14251);
or UO_1260 (O_1260,N_12554,N_14836);
or UO_1261 (O_1261,N_13966,N_13263);
xnor UO_1262 (O_1262,N_14180,N_14524);
or UO_1263 (O_1263,N_12423,N_14156);
nor UO_1264 (O_1264,N_13864,N_14507);
xor UO_1265 (O_1265,N_12787,N_12690);
and UO_1266 (O_1266,N_14187,N_14453);
nor UO_1267 (O_1267,N_12329,N_13600);
xnor UO_1268 (O_1268,N_13970,N_12629);
nand UO_1269 (O_1269,N_14045,N_13109);
and UO_1270 (O_1270,N_13351,N_12906);
or UO_1271 (O_1271,N_13435,N_13371);
nand UO_1272 (O_1272,N_12617,N_12369);
nor UO_1273 (O_1273,N_12707,N_13859);
or UO_1274 (O_1274,N_14404,N_13286);
and UO_1275 (O_1275,N_13846,N_13277);
xor UO_1276 (O_1276,N_12359,N_13278);
xor UO_1277 (O_1277,N_14848,N_13313);
and UO_1278 (O_1278,N_12068,N_14354);
nand UO_1279 (O_1279,N_13406,N_13260);
and UO_1280 (O_1280,N_12555,N_13049);
and UO_1281 (O_1281,N_12060,N_14545);
and UO_1282 (O_1282,N_14883,N_14237);
nor UO_1283 (O_1283,N_13253,N_14006);
or UO_1284 (O_1284,N_12740,N_12084);
or UO_1285 (O_1285,N_12759,N_13696);
nor UO_1286 (O_1286,N_12583,N_14594);
nand UO_1287 (O_1287,N_12112,N_13716);
and UO_1288 (O_1288,N_13008,N_14391);
or UO_1289 (O_1289,N_14896,N_13244);
xnor UO_1290 (O_1290,N_13172,N_14204);
xor UO_1291 (O_1291,N_12154,N_13888);
nor UO_1292 (O_1292,N_14027,N_13758);
nor UO_1293 (O_1293,N_12934,N_14975);
nor UO_1294 (O_1294,N_13954,N_13139);
and UO_1295 (O_1295,N_14865,N_14096);
nor UO_1296 (O_1296,N_13356,N_13576);
and UO_1297 (O_1297,N_14543,N_12767);
nor UO_1298 (O_1298,N_12863,N_12181);
or UO_1299 (O_1299,N_12193,N_13328);
xor UO_1300 (O_1300,N_14401,N_14886);
and UO_1301 (O_1301,N_14290,N_13074);
or UO_1302 (O_1302,N_13459,N_13900);
xnor UO_1303 (O_1303,N_12898,N_12415);
nand UO_1304 (O_1304,N_14789,N_12186);
and UO_1305 (O_1305,N_13675,N_12311);
xor UO_1306 (O_1306,N_13602,N_14722);
xor UO_1307 (O_1307,N_13793,N_14675);
or UO_1308 (O_1308,N_12297,N_12546);
nand UO_1309 (O_1309,N_13474,N_14117);
or UO_1310 (O_1310,N_12296,N_12279);
xnor UO_1311 (O_1311,N_14943,N_12389);
nor UO_1312 (O_1312,N_12149,N_13507);
or UO_1313 (O_1313,N_12281,N_14231);
or UO_1314 (O_1314,N_14380,N_12996);
and UO_1315 (O_1315,N_12377,N_12235);
nand UO_1316 (O_1316,N_12212,N_14869);
xnor UO_1317 (O_1317,N_12300,N_14611);
and UO_1318 (O_1318,N_13120,N_12298);
or UO_1319 (O_1319,N_13522,N_14668);
and UO_1320 (O_1320,N_13066,N_14968);
nor UO_1321 (O_1321,N_13513,N_14349);
and UO_1322 (O_1322,N_13417,N_13629);
xnor UO_1323 (O_1323,N_14110,N_13634);
nand UO_1324 (O_1324,N_12735,N_14584);
xnor UO_1325 (O_1325,N_12474,N_12937);
or UO_1326 (O_1326,N_12087,N_13029);
or UO_1327 (O_1327,N_14637,N_13614);
nand UO_1328 (O_1328,N_13687,N_13983);
or UO_1329 (O_1329,N_12164,N_12204);
nor UO_1330 (O_1330,N_12043,N_13202);
and UO_1331 (O_1331,N_13389,N_12195);
and UO_1332 (O_1332,N_12018,N_12200);
xor UO_1333 (O_1333,N_14525,N_13855);
or UO_1334 (O_1334,N_13065,N_12920);
or UO_1335 (O_1335,N_14793,N_13979);
nor UO_1336 (O_1336,N_13528,N_13658);
nand UO_1337 (O_1337,N_14520,N_14418);
or UO_1338 (O_1338,N_13316,N_13249);
and UO_1339 (O_1339,N_14433,N_14994);
or UO_1340 (O_1340,N_13462,N_14752);
and UO_1341 (O_1341,N_12236,N_13912);
or UO_1342 (O_1342,N_12975,N_14631);
and UO_1343 (O_1343,N_14995,N_12988);
nor UO_1344 (O_1344,N_13555,N_13379);
xor UO_1345 (O_1345,N_12241,N_14966);
nor UO_1346 (O_1346,N_12071,N_14809);
nand UO_1347 (O_1347,N_13710,N_12624);
nand UO_1348 (O_1348,N_14874,N_12782);
nor UO_1349 (O_1349,N_12139,N_12918);
or UO_1350 (O_1350,N_14245,N_13067);
nor UO_1351 (O_1351,N_12378,N_14048);
and UO_1352 (O_1352,N_14761,N_14960);
nand UO_1353 (O_1353,N_14268,N_13205);
nor UO_1354 (O_1354,N_14510,N_12980);
xnor UO_1355 (O_1355,N_14050,N_14872);
nand UO_1356 (O_1356,N_14190,N_13743);
xor UO_1357 (O_1357,N_13116,N_13464);
xor UO_1358 (O_1358,N_13949,N_13699);
nor UO_1359 (O_1359,N_13504,N_14684);
nand UO_1360 (O_1360,N_12367,N_13175);
xnor UO_1361 (O_1361,N_13329,N_12613);
and UO_1362 (O_1362,N_14718,N_14688);
nand UO_1363 (O_1363,N_14186,N_14724);
nor UO_1364 (O_1364,N_12704,N_12354);
and UO_1365 (O_1365,N_14905,N_12871);
nand UO_1366 (O_1366,N_12938,N_14314);
xnor UO_1367 (O_1367,N_13988,N_12386);
nand UO_1368 (O_1368,N_12303,N_14538);
and UO_1369 (O_1369,N_12588,N_13578);
nand UO_1370 (O_1370,N_13535,N_13140);
and UO_1371 (O_1371,N_14037,N_14258);
nand UO_1372 (O_1372,N_14956,N_14445);
and UO_1373 (O_1373,N_13194,N_13150);
xor UO_1374 (O_1374,N_13789,N_12114);
xnor UO_1375 (O_1375,N_13702,N_13712);
xor UO_1376 (O_1376,N_14866,N_14304);
and UO_1377 (O_1377,N_12491,N_13672);
xor UO_1378 (O_1378,N_14089,N_14101);
nand UO_1379 (O_1379,N_12484,N_13298);
or UO_1380 (O_1380,N_12577,N_13999);
nor UO_1381 (O_1381,N_13674,N_13854);
nand UO_1382 (O_1382,N_13991,N_14822);
or UO_1383 (O_1383,N_13055,N_14074);
xnor UO_1384 (O_1384,N_14298,N_13402);
and UO_1385 (O_1385,N_13551,N_13234);
nand UO_1386 (O_1386,N_13088,N_12839);
nor UO_1387 (O_1387,N_13124,N_13475);
nand UO_1388 (O_1388,N_12813,N_14774);
xnor UO_1389 (O_1389,N_14648,N_13121);
nand UO_1390 (O_1390,N_12884,N_12847);
nor UO_1391 (O_1391,N_14449,N_13076);
or UO_1392 (O_1392,N_14474,N_13807);
nand UO_1393 (O_1393,N_12420,N_12480);
and UO_1394 (O_1394,N_13783,N_13751);
nor UO_1395 (O_1395,N_12557,N_14491);
nor UO_1396 (O_1396,N_14615,N_13129);
nor UO_1397 (O_1397,N_12096,N_12174);
and UO_1398 (O_1398,N_12032,N_14981);
xor UO_1399 (O_1399,N_14629,N_13104);
nand UO_1400 (O_1400,N_14230,N_14653);
xor UO_1401 (O_1401,N_14903,N_13874);
and UO_1402 (O_1402,N_14605,N_14235);
or UO_1403 (O_1403,N_13525,N_12945);
xnor UO_1404 (O_1404,N_14596,N_12927);
xnor UO_1405 (O_1405,N_14179,N_12337);
and UO_1406 (O_1406,N_13582,N_13771);
nand UO_1407 (O_1407,N_14182,N_12141);
or UO_1408 (O_1408,N_14113,N_14168);
and UO_1409 (O_1409,N_13804,N_13030);
or UO_1410 (O_1410,N_13942,N_14560);
nor UO_1411 (O_1411,N_12108,N_13482);
xor UO_1412 (O_1412,N_12879,N_13044);
xnor UO_1413 (O_1413,N_13376,N_14346);
or UO_1414 (O_1414,N_12786,N_12398);
nor UO_1415 (O_1415,N_14283,N_12719);
or UO_1416 (O_1416,N_14058,N_14206);
nand UO_1417 (O_1417,N_12859,N_12821);
nor UO_1418 (O_1418,N_12794,N_14274);
or UO_1419 (O_1419,N_13180,N_12828);
nor UO_1420 (O_1420,N_13383,N_14974);
or UO_1421 (O_1421,N_13867,N_14092);
and UO_1422 (O_1422,N_12513,N_13468);
nand UO_1423 (O_1423,N_13986,N_13671);
nor UO_1424 (O_1424,N_12653,N_13339);
xor UO_1425 (O_1425,N_14820,N_14004);
xor UO_1426 (O_1426,N_13883,N_12454);
or UO_1427 (O_1427,N_12973,N_12334);
xor UO_1428 (O_1428,N_13944,N_14513);
nand UO_1429 (O_1429,N_13866,N_12260);
nor UO_1430 (O_1430,N_14519,N_12913);
xor UO_1431 (O_1431,N_12233,N_14621);
or UO_1432 (O_1432,N_14297,N_14990);
xor UO_1433 (O_1433,N_14712,N_12436);
nor UO_1434 (O_1434,N_13185,N_12102);
or UO_1435 (O_1435,N_13289,N_13362);
nor UO_1436 (O_1436,N_14742,N_12525);
xor UO_1437 (O_1437,N_14846,N_13346);
nor UO_1438 (O_1438,N_14130,N_14527);
xnor UO_1439 (O_1439,N_14861,N_14598);
and UO_1440 (O_1440,N_12091,N_14747);
xnor UO_1441 (O_1441,N_13805,N_14286);
xnor UO_1442 (O_1442,N_13363,N_14403);
nor UO_1443 (O_1443,N_13453,N_12626);
xnor UO_1444 (O_1444,N_13544,N_14592);
nand UO_1445 (O_1445,N_12753,N_14801);
nand UO_1446 (O_1446,N_14384,N_12522);
or UO_1447 (O_1447,N_13896,N_12162);
xor UO_1448 (O_1448,N_12031,N_12586);
and UO_1449 (O_1449,N_12541,N_12213);
nand UO_1450 (O_1450,N_13223,N_12042);
xnor UO_1451 (O_1451,N_14756,N_12182);
or UO_1452 (O_1452,N_13451,N_13626);
and UO_1453 (O_1453,N_13449,N_12397);
or UO_1454 (O_1454,N_13619,N_13321);
or UO_1455 (O_1455,N_12739,N_12284);
or UO_1456 (O_1456,N_13994,N_13630);
nor UO_1457 (O_1457,N_14649,N_13000);
or UO_1458 (O_1458,N_12984,N_14094);
nor UO_1459 (O_1459,N_14154,N_14375);
xnor UO_1460 (O_1460,N_13220,N_13625);
xor UO_1461 (O_1461,N_14038,N_13361);
nor UO_1462 (O_1462,N_13017,N_13415);
nor UO_1463 (O_1463,N_13229,N_13796);
xnor UO_1464 (O_1464,N_12570,N_14109);
and UO_1465 (O_1465,N_14344,N_12659);
nand UO_1466 (O_1466,N_12696,N_14588);
nor UO_1467 (O_1467,N_13466,N_12105);
nor UO_1468 (O_1468,N_13267,N_14277);
and UO_1469 (O_1469,N_13075,N_14152);
or UO_1470 (O_1470,N_14646,N_13620);
or UO_1471 (O_1471,N_12240,N_14140);
or UO_1472 (O_1472,N_14497,N_14234);
or UO_1473 (O_1473,N_13237,N_13160);
nand UO_1474 (O_1474,N_12086,N_12118);
nand UO_1475 (O_1475,N_12754,N_14232);
nand UO_1476 (O_1476,N_13610,N_14017);
nor UO_1477 (O_1477,N_12507,N_12824);
nand UO_1478 (O_1478,N_14016,N_12394);
xnor UO_1479 (O_1479,N_14725,N_12997);
xnor UO_1480 (O_1480,N_13193,N_12618);
xor UO_1481 (O_1481,N_14366,N_12751);
and UO_1482 (O_1482,N_12535,N_14312);
or UO_1483 (O_1483,N_14492,N_13833);
nand UO_1484 (O_1484,N_12688,N_13872);
and UO_1485 (O_1485,N_12675,N_12969);
nand UO_1486 (O_1486,N_12998,N_13821);
and UO_1487 (O_1487,N_12266,N_13982);
nand UO_1488 (O_1488,N_12702,N_14382);
xor UO_1489 (O_1489,N_13407,N_13235);
nand UO_1490 (O_1490,N_14248,N_14549);
xnor UO_1491 (O_1491,N_13128,N_12362);
nor UO_1492 (O_1492,N_14988,N_14365);
nand UO_1493 (O_1493,N_12176,N_14160);
xnor UO_1494 (O_1494,N_14984,N_14821);
xnor UO_1495 (O_1495,N_13707,N_12693);
nor UO_1496 (O_1496,N_12582,N_13973);
xor UO_1497 (O_1497,N_13742,N_13092);
nor UO_1498 (O_1498,N_12757,N_12455);
and UO_1499 (O_1499,N_14651,N_14428);
xor UO_1500 (O_1500,N_14354,N_14734);
nor UO_1501 (O_1501,N_13929,N_12544);
xor UO_1502 (O_1502,N_14443,N_14685);
xor UO_1503 (O_1503,N_12968,N_12246);
or UO_1504 (O_1504,N_14110,N_14454);
nor UO_1505 (O_1505,N_14950,N_14519);
nor UO_1506 (O_1506,N_13099,N_12558);
xnor UO_1507 (O_1507,N_12032,N_14021);
nand UO_1508 (O_1508,N_14393,N_12108);
nand UO_1509 (O_1509,N_14006,N_12862);
xor UO_1510 (O_1510,N_12000,N_14412);
nand UO_1511 (O_1511,N_13847,N_13230);
or UO_1512 (O_1512,N_14822,N_13398);
or UO_1513 (O_1513,N_13323,N_13296);
xnor UO_1514 (O_1514,N_13000,N_13206);
nor UO_1515 (O_1515,N_14277,N_13748);
and UO_1516 (O_1516,N_12923,N_14024);
nor UO_1517 (O_1517,N_13916,N_12918);
nand UO_1518 (O_1518,N_12744,N_14019);
nor UO_1519 (O_1519,N_13617,N_12920);
nand UO_1520 (O_1520,N_14957,N_12884);
nor UO_1521 (O_1521,N_13321,N_12038);
xor UO_1522 (O_1522,N_14031,N_14407);
nand UO_1523 (O_1523,N_12591,N_14901);
nor UO_1524 (O_1524,N_13789,N_14666);
xnor UO_1525 (O_1525,N_12467,N_12290);
or UO_1526 (O_1526,N_13212,N_12428);
or UO_1527 (O_1527,N_14972,N_12763);
xnor UO_1528 (O_1528,N_13566,N_14138);
or UO_1529 (O_1529,N_14854,N_14424);
nor UO_1530 (O_1530,N_12179,N_13857);
xnor UO_1531 (O_1531,N_13783,N_12849);
xnor UO_1532 (O_1532,N_12557,N_14395);
nor UO_1533 (O_1533,N_14638,N_12633);
or UO_1534 (O_1534,N_12587,N_12299);
and UO_1535 (O_1535,N_14948,N_14294);
and UO_1536 (O_1536,N_13622,N_14034);
nand UO_1537 (O_1537,N_14315,N_14567);
or UO_1538 (O_1538,N_13303,N_12470);
nand UO_1539 (O_1539,N_14732,N_14898);
and UO_1540 (O_1540,N_13943,N_12152);
xor UO_1541 (O_1541,N_13320,N_14595);
xnor UO_1542 (O_1542,N_13158,N_14223);
nor UO_1543 (O_1543,N_14385,N_12766);
or UO_1544 (O_1544,N_14758,N_12107);
nand UO_1545 (O_1545,N_13598,N_12444);
or UO_1546 (O_1546,N_12984,N_14078);
or UO_1547 (O_1547,N_12082,N_12966);
xor UO_1548 (O_1548,N_14215,N_13449);
nor UO_1549 (O_1549,N_12763,N_12732);
and UO_1550 (O_1550,N_13250,N_13374);
or UO_1551 (O_1551,N_12001,N_13712);
nand UO_1552 (O_1552,N_14887,N_14861);
nand UO_1553 (O_1553,N_14744,N_14757);
or UO_1554 (O_1554,N_12656,N_14299);
xor UO_1555 (O_1555,N_12692,N_14436);
nor UO_1556 (O_1556,N_13839,N_13844);
nor UO_1557 (O_1557,N_14363,N_14687);
nand UO_1558 (O_1558,N_12908,N_12367);
nand UO_1559 (O_1559,N_14846,N_14310);
xor UO_1560 (O_1560,N_13414,N_14703);
xor UO_1561 (O_1561,N_12320,N_13788);
and UO_1562 (O_1562,N_13165,N_13573);
or UO_1563 (O_1563,N_14978,N_14899);
or UO_1564 (O_1564,N_12116,N_12260);
nand UO_1565 (O_1565,N_14625,N_12436);
nand UO_1566 (O_1566,N_13492,N_14730);
or UO_1567 (O_1567,N_12526,N_14373);
nor UO_1568 (O_1568,N_12097,N_12816);
nand UO_1569 (O_1569,N_12046,N_14859);
nand UO_1570 (O_1570,N_12419,N_12277);
xor UO_1571 (O_1571,N_12788,N_13555);
or UO_1572 (O_1572,N_14801,N_13645);
xor UO_1573 (O_1573,N_12803,N_12826);
or UO_1574 (O_1574,N_13801,N_13756);
nand UO_1575 (O_1575,N_14704,N_13550);
nand UO_1576 (O_1576,N_12215,N_14694);
xnor UO_1577 (O_1577,N_12961,N_13897);
nand UO_1578 (O_1578,N_13653,N_12085);
and UO_1579 (O_1579,N_12062,N_14614);
nor UO_1580 (O_1580,N_14449,N_13007);
nor UO_1581 (O_1581,N_13872,N_12848);
nor UO_1582 (O_1582,N_12537,N_13935);
xor UO_1583 (O_1583,N_13119,N_12374);
nand UO_1584 (O_1584,N_12885,N_12373);
xnor UO_1585 (O_1585,N_12103,N_12226);
nor UO_1586 (O_1586,N_14446,N_13593);
nor UO_1587 (O_1587,N_14689,N_14010);
nor UO_1588 (O_1588,N_12150,N_14336);
nand UO_1589 (O_1589,N_12534,N_12267);
and UO_1590 (O_1590,N_12785,N_13351);
and UO_1591 (O_1591,N_14492,N_13336);
nor UO_1592 (O_1592,N_14095,N_13185);
xnor UO_1593 (O_1593,N_12822,N_13613);
and UO_1594 (O_1594,N_14064,N_12727);
nand UO_1595 (O_1595,N_14602,N_13115);
nor UO_1596 (O_1596,N_13054,N_12992);
or UO_1597 (O_1597,N_14931,N_13439);
nor UO_1598 (O_1598,N_14420,N_14081);
nand UO_1599 (O_1599,N_12961,N_13102);
nor UO_1600 (O_1600,N_12715,N_14398);
nand UO_1601 (O_1601,N_14146,N_12071);
and UO_1602 (O_1602,N_12881,N_13452);
xnor UO_1603 (O_1603,N_14039,N_14487);
xor UO_1604 (O_1604,N_12458,N_12409);
and UO_1605 (O_1605,N_12403,N_12145);
or UO_1606 (O_1606,N_13812,N_12946);
nand UO_1607 (O_1607,N_12998,N_12507);
and UO_1608 (O_1608,N_14325,N_13191);
xnor UO_1609 (O_1609,N_13310,N_14862);
and UO_1610 (O_1610,N_14329,N_14122);
or UO_1611 (O_1611,N_13787,N_14245);
nor UO_1612 (O_1612,N_14213,N_12292);
nor UO_1613 (O_1613,N_14033,N_14120);
nand UO_1614 (O_1614,N_13457,N_14376);
and UO_1615 (O_1615,N_12372,N_14514);
nor UO_1616 (O_1616,N_13655,N_14515);
or UO_1617 (O_1617,N_14635,N_12994);
xor UO_1618 (O_1618,N_12636,N_12689);
or UO_1619 (O_1619,N_12529,N_13959);
xnor UO_1620 (O_1620,N_14328,N_12350);
xor UO_1621 (O_1621,N_13780,N_14473);
and UO_1622 (O_1622,N_14487,N_12647);
xor UO_1623 (O_1623,N_12818,N_14399);
or UO_1624 (O_1624,N_14657,N_14571);
or UO_1625 (O_1625,N_13215,N_13667);
nand UO_1626 (O_1626,N_13254,N_13304);
and UO_1627 (O_1627,N_14545,N_13021);
nand UO_1628 (O_1628,N_14744,N_12210);
nand UO_1629 (O_1629,N_13599,N_14082);
nand UO_1630 (O_1630,N_13194,N_14057);
xor UO_1631 (O_1631,N_14745,N_12231);
and UO_1632 (O_1632,N_12230,N_12122);
xor UO_1633 (O_1633,N_14258,N_14636);
or UO_1634 (O_1634,N_12961,N_14021);
or UO_1635 (O_1635,N_12345,N_14087);
or UO_1636 (O_1636,N_13454,N_13763);
nor UO_1637 (O_1637,N_13227,N_14960);
nand UO_1638 (O_1638,N_12059,N_13808);
or UO_1639 (O_1639,N_14006,N_14168);
or UO_1640 (O_1640,N_12651,N_13423);
and UO_1641 (O_1641,N_12796,N_12533);
nor UO_1642 (O_1642,N_13638,N_13325);
xnor UO_1643 (O_1643,N_13426,N_13496);
nor UO_1644 (O_1644,N_13278,N_12788);
nor UO_1645 (O_1645,N_12034,N_14742);
nand UO_1646 (O_1646,N_13937,N_13367);
and UO_1647 (O_1647,N_13185,N_13739);
and UO_1648 (O_1648,N_12756,N_13275);
or UO_1649 (O_1649,N_12016,N_12716);
nand UO_1650 (O_1650,N_14784,N_14186);
or UO_1651 (O_1651,N_13471,N_13894);
xnor UO_1652 (O_1652,N_14217,N_12418);
nand UO_1653 (O_1653,N_12278,N_13004);
and UO_1654 (O_1654,N_12445,N_13520);
nand UO_1655 (O_1655,N_14186,N_14402);
and UO_1656 (O_1656,N_12405,N_14448);
or UO_1657 (O_1657,N_12619,N_12897);
nor UO_1658 (O_1658,N_13288,N_12980);
nand UO_1659 (O_1659,N_14789,N_12110);
nor UO_1660 (O_1660,N_14857,N_13958);
or UO_1661 (O_1661,N_12011,N_12398);
nand UO_1662 (O_1662,N_12217,N_14463);
or UO_1663 (O_1663,N_13048,N_14214);
or UO_1664 (O_1664,N_13813,N_13579);
nor UO_1665 (O_1665,N_14467,N_13215);
nand UO_1666 (O_1666,N_14599,N_13804);
nor UO_1667 (O_1667,N_12486,N_14761);
xor UO_1668 (O_1668,N_14717,N_12902);
xnor UO_1669 (O_1669,N_12456,N_12761);
and UO_1670 (O_1670,N_12919,N_13697);
nor UO_1671 (O_1671,N_13807,N_14852);
and UO_1672 (O_1672,N_13487,N_14259);
or UO_1673 (O_1673,N_13593,N_12850);
and UO_1674 (O_1674,N_14782,N_12562);
or UO_1675 (O_1675,N_12844,N_12866);
nand UO_1676 (O_1676,N_12691,N_12106);
nor UO_1677 (O_1677,N_12999,N_14576);
nand UO_1678 (O_1678,N_13521,N_13787);
and UO_1679 (O_1679,N_12228,N_14642);
nand UO_1680 (O_1680,N_14994,N_13707);
nand UO_1681 (O_1681,N_14578,N_13968);
xor UO_1682 (O_1682,N_14682,N_14647);
nand UO_1683 (O_1683,N_13449,N_12814);
nand UO_1684 (O_1684,N_12155,N_12665);
nor UO_1685 (O_1685,N_14973,N_13919);
and UO_1686 (O_1686,N_12866,N_13289);
and UO_1687 (O_1687,N_13082,N_14805);
nor UO_1688 (O_1688,N_14070,N_14780);
xor UO_1689 (O_1689,N_14197,N_13809);
xnor UO_1690 (O_1690,N_14705,N_14400);
and UO_1691 (O_1691,N_14624,N_14406);
or UO_1692 (O_1692,N_13145,N_12463);
and UO_1693 (O_1693,N_12628,N_14899);
nand UO_1694 (O_1694,N_13778,N_12511);
xnor UO_1695 (O_1695,N_14518,N_12511);
nand UO_1696 (O_1696,N_14984,N_13889);
nor UO_1697 (O_1697,N_13772,N_14174);
xnor UO_1698 (O_1698,N_13783,N_14128);
xnor UO_1699 (O_1699,N_14674,N_12421);
nand UO_1700 (O_1700,N_13550,N_12772);
xnor UO_1701 (O_1701,N_13839,N_14320);
nor UO_1702 (O_1702,N_14320,N_12669);
or UO_1703 (O_1703,N_13043,N_12248);
nor UO_1704 (O_1704,N_12816,N_14236);
and UO_1705 (O_1705,N_14660,N_13832);
xor UO_1706 (O_1706,N_12982,N_14101);
nor UO_1707 (O_1707,N_13036,N_12971);
xor UO_1708 (O_1708,N_14841,N_14267);
or UO_1709 (O_1709,N_14196,N_13502);
or UO_1710 (O_1710,N_13357,N_13702);
nor UO_1711 (O_1711,N_14241,N_12906);
nor UO_1712 (O_1712,N_14168,N_13263);
nor UO_1713 (O_1713,N_13186,N_14587);
nor UO_1714 (O_1714,N_13328,N_12992);
nand UO_1715 (O_1715,N_12955,N_13977);
or UO_1716 (O_1716,N_13682,N_14019);
xnor UO_1717 (O_1717,N_14236,N_14009);
and UO_1718 (O_1718,N_12268,N_13237);
nor UO_1719 (O_1719,N_13291,N_13948);
and UO_1720 (O_1720,N_12628,N_13873);
nand UO_1721 (O_1721,N_12256,N_12491);
nor UO_1722 (O_1722,N_12156,N_14417);
or UO_1723 (O_1723,N_14685,N_13106);
nand UO_1724 (O_1724,N_13914,N_13089);
xnor UO_1725 (O_1725,N_13033,N_14125);
nand UO_1726 (O_1726,N_13489,N_12570);
nand UO_1727 (O_1727,N_13267,N_14246);
xnor UO_1728 (O_1728,N_12600,N_13391);
and UO_1729 (O_1729,N_14813,N_13478);
and UO_1730 (O_1730,N_13272,N_13241);
and UO_1731 (O_1731,N_14887,N_12932);
xor UO_1732 (O_1732,N_12875,N_12382);
xnor UO_1733 (O_1733,N_12920,N_14934);
or UO_1734 (O_1734,N_12135,N_14339);
and UO_1735 (O_1735,N_12157,N_13355);
nand UO_1736 (O_1736,N_12315,N_12135);
or UO_1737 (O_1737,N_13800,N_14693);
or UO_1738 (O_1738,N_12600,N_14848);
nand UO_1739 (O_1739,N_13472,N_13892);
nor UO_1740 (O_1740,N_14155,N_14994);
nand UO_1741 (O_1741,N_12475,N_12634);
nand UO_1742 (O_1742,N_14162,N_12823);
and UO_1743 (O_1743,N_13740,N_13207);
nor UO_1744 (O_1744,N_13085,N_14153);
xor UO_1745 (O_1745,N_13817,N_14215);
or UO_1746 (O_1746,N_14242,N_14815);
nor UO_1747 (O_1747,N_14536,N_13485);
xor UO_1748 (O_1748,N_12460,N_14874);
xor UO_1749 (O_1749,N_12898,N_12036);
nand UO_1750 (O_1750,N_14491,N_14629);
nor UO_1751 (O_1751,N_13320,N_12341);
xor UO_1752 (O_1752,N_13559,N_14691);
or UO_1753 (O_1753,N_13385,N_13177);
nand UO_1754 (O_1754,N_12359,N_13779);
xor UO_1755 (O_1755,N_13309,N_13996);
nor UO_1756 (O_1756,N_12112,N_13486);
and UO_1757 (O_1757,N_14005,N_14143);
nand UO_1758 (O_1758,N_12236,N_14595);
or UO_1759 (O_1759,N_14031,N_13043);
xor UO_1760 (O_1760,N_12131,N_14504);
and UO_1761 (O_1761,N_12775,N_12281);
xnor UO_1762 (O_1762,N_12864,N_14431);
nor UO_1763 (O_1763,N_14172,N_13833);
nand UO_1764 (O_1764,N_14577,N_14229);
nor UO_1765 (O_1765,N_14046,N_13920);
and UO_1766 (O_1766,N_13112,N_13454);
or UO_1767 (O_1767,N_12347,N_13295);
nor UO_1768 (O_1768,N_13736,N_13447);
and UO_1769 (O_1769,N_13410,N_13338);
and UO_1770 (O_1770,N_13166,N_14151);
xnor UO_1771 (O_1771,N_13559,N_14225);
or UO_1772 (O_1772,N_13818,N_12914);
xnor UO_1773 (O_1773,N_12754,N_13840);
and UO_1774 (O_1774,N_14979,N_14638);
or UO_1775 (O_1775,N_12659,N_13351);
nor UO_1776 (O_1776,N_14773,N_14436);
xor UO_1777 (O_1777,N_14885,N_12572);
nor UO_1778 (O_1778,N_14282,N_12079);
and UO_1779 (O_1779,N_12661,N_12124);
xnor UO_1780 (O_1780,N_12420,N_14881);
nor UO_1781 (O_1781,N_14270,N_12977);
xnor UO_1782 (O_1782,N_13909,N_13977);
xnor UO_1783 (O_1783,N_13852,N_14720);
xnor UO_1784 (O_1784,N_13004,N_14369);
nand UO_1785 (O_1785,N_12902,N_14033);
xnor UO_1786 (O_1786,N_12549,N_14588);
nand UO_1787 (O_1787,N_13279,N_14648);
nand UO_1788 (O_1788,N_14138,N_12018);
nand UO_1789 (O_1789,N_14601,N_12243);
nand UO_1790 (O_1790,N_14875,N_14033);
or UO_1791 (O_1791,N_13956,N_13330);
and UO_1792 (O_1792,N_12146,N_12075);
nor UO_1793 (O_1793,N_14713,N_12156);
nand UO_1794 (O_1794,N_13432,N_14442);
or UO_1795 (O_1795,N_14427,N_12278);
and UO_1796 (O_1796,N_12130,N_13062);
and UO_1797 (O_1797,N_13881,N_12417);
xor UO_1798 (O_1798,N_12677,N_13994);
xor UO_1799 (O_1799,N_14368,N_14830);
nand UO_1800 (O_1800,N_12839,N_14372);
nor UO_1801 (O_1801,N_13446,N_14321);
nand UO_1802 (O_1802,N_14814,N_14943);
or UO_1803 (O_1803,N_12790,N_14943);
xor UO_1804 (O_1804,N_12714,N_12330);
and UO_1805 (O_1805,N_14339,N_14897);
or UO_1806 (O_1806,N_12198,N_12568);
nand UO_1807 (O_1807,N_12267,N_13138);
nor UO_1808 (O_1808,N_13844,N_13462);
xnor UO_1809 (O_1809,N_14637,N_14995);
nand UO_1810 (O_1810,N_13775,N_13654);
xor UO_1811 (O_1811,N_14575,N_13690);
nand UO_1812 (O_1812,N_12960,N_14332);
xnor UO_1813 (O_1813,N_14129,N_13049);
nor UO_1814 (O_1814,N_12976,N_12754);
nand UO_1815 (O_1815,N_13709,N_14536);
nor UO_1816 (O_1816,N_13098,N_14236);
nor UO_1817 (O_1817,N_13234,N_14183);
xor UO_1818 (O_1818,N_13085,N_12064);
or UO_1819 (O_1819,N_14181,N_14028);
nand UO_1820 (O_1820,N_14489,N_13109);
nand UO_1821 (O_1821,N_12836,N_13513);
xor UO_1822 (O_1822,N_13462,N_14525);
nor UO_1823 (O_1823,N_13559,N_14258);
nand UO_1824 (O_1824,N_14519,N_12819);
and UO_1825 (O_1825,N_12999,N_13420);
and UO_1826 (O_1826,N_14717,N_14223);
and UO_1827 (O_1827,N_13861,N_14992);
nor UO_1828 (O_1828,N_13178,N_12516);
or UO_1829 (O_1829,N_13089,N_14567);
nand UO_1830 (O_1830,N_13329,N_14563);
and UO_1831 (O_1831,N_14666,N_12408);
or UO_1832 (O_1832,N_12599,N_12162);
nor UO_1833 (O_1833,N_13885,N_12356);
xnor UO_1834 (O_1834,N_13409,N_12277);
nor UO_1835 (O_1835,N_12508,N_12155);
or UO_1836 (O_1836,N_13942,N_14002);
nand UO_1837 (O_1837,N_13396,N_13442);
and UO_1838 (O_1838,N_13608,N_12357);
nor UO_1839 (O_1839,N_12230,N_14933);
xnor UO_1840 (O_1840,N_12692,N_12976);
xor UO_1841 (O_1841,N_14319,N_12714);
or UO_1842 (O_1842,N_12290,N_12641);
nor UO_1843 (O_1843,N_14973,N_14502);
or UO_1844 (O_1844,N_12368,N_12817);
or UO_1845 (O_1845,N_14196,N_12639);
xnor UO_1846 (O_1846,N_12289,N_13510);
nand UO_1847 (O_1847,N_13897,N_14962);
nor UO_1848 (O_1848,N_12474,N_12979);
and UO_1849 (O_1849,N_14467,N_14411);
and UO_1850 (O_1850,N_13129,N_12355);
nand UO_1851 (O_1851,N_13145,N_12813);
or UO_1852 (O_1852,N_14568,N_13687);
and UO_1853 (O_1853,N_13038,N_14454);
nand UO_1854 (O_1854,N_14856,N_13939);
nor UO_1855 (O_1855,N_12817,N_13124);
nand UO_1856 (O_1856,N_14846,N_12937);
xnor UO_1857 (O_1857,N_13039,N_14323);
or UO_1858 (O_1858,N_14014,N_12516);
nand UO_1859 (O_1859,N_14346,N_13428);
or UO_1860 (O_1860,N_14142,N_12316);
and UO_1861 (O_1861,N_14441,N_13468);
xor UO_1862 (O_1862,N_12270,N_13602);
xor UO_1863 (O_1863,N_12334,N_14939);
and UO_1864 (O_1864,N_14983,N_14362);
xnor UO_1865 (O_1865,N_12399,N_12727);
nand UO_1866 (O_1866,N_14772,N_13803);
xnor UO_1867 (O_1867,N_13211,N_14070);
and UO_1868 (O_1868,N_12554,N_12457);
nor UO_1869 (O_1869,N_14466,N_14573);
nand UO_1870 (O_1870,N_14474,N_14974);
xor UO_1871 (O_1871,N_14880,N_14443);
and UO_1872 (O_1872,N_14315,N_13785);
and UO_1873 (O_1873,N_13211,N_12879);
nor UO_1874 (O_1874,N_12654,N_13084);
or UO_1875 (O_1875,N_14226,N_13605);
xor UO_1876 (O_1876,N_13465,N_14623);
xor UO_1877 (O_1877,N_13086,N_14437);
nand UO_1878 (O_1878,N_13967,N_13277);
xnor UO_1879 (O_1879,N_12300,N_14690);
nand UO_1880 (O_1880,N_13467,N_13652);
xnor UO_1881 (O_1881,N_14119,N_12467);
nor UO_1882 (O_1882,N_13708,N_13237);
nand UO_1883 (O_1883,N_12846,N_14641);
nor UO_1884 (O_1884,N_13812,N_13218);
nor UO_1885 (O_1885,N_13107,N_13990);
nor UO_1886 (O_1886,N_12314,N_13100);
xnor UO_1887 (O_1887,N_13409,N_13646);
or UO_1888 (O_1888,N_13481,N_12820);
or UO_1889 (O_1889,N_14676,N_13233);
or UO_1890 (O_1890,N_14488,N_14844);
or UO_1891 (O_1891,N_13214,N_12729);
nand UO_1892 (O_1892,N_14519,N_13647);
xnor UO_1893 (O_1893,N_12926,N_14915);
nand UO_1894 (O_1894,N_13526,N_12817);
or UO_1895 (O_1895,N_13208,N_13095);
or UO_1896 (O_1896,N_13833,N_13912);
nor UO_1897 (O_1897,N_12794,N_13698);
and UO_1898 (O_1898,N_14051,N_14254);
nand UO_1899 (O_1899,N_14049,N_12137);
nand UO_1900 (O_1900,N_14955,N_14695);
xnor UO_1901 (O_1901,N_12855,N_13625);
xor UO_1902 (O_1902,N_12616,N_13725);
nand UO_1903 (O_1903,N_14065,N_13018);
nor UO_1904 (O_1904,N_13369,N_14562);
and UO_1905 (O_1905,N_12742,N_12300);
or UO_1906 (O_1906,N_14592,N_12672);
xnor UO_1907 (O_1907,N_13713,N_14437);
nor UO_1908 (O_1908,N_14574,N_13434);
or UO_1909 (O_1909,N_14253,N_14881);
nor UO_1910 (O_1910,N_14061,N_12551);
nor UO_1911 (O_1911,N_12525,N_12023);
and UO_1912 (O_1912,N_14590,N_13178);
nor UO_1913 (O_1913,N_13697,N_13860);
and UO_1914 (O_1914,N_12996,N_14271);
xor UO_1915 (O_1915,N_12453,N_13162);
nand UO_1916 (O_1916,N_13620,N_14558);
and UO_1917 (O_1917,N_12488,N_14019);
nor UO_1918 (O_1918,N_14071,N_12943);
or UO_1919 (O_1919,N_14458,N_12261);
nor UO_1920 (O_1920,N_12028,N_12816);
xor UO_1921 (O_1921,N_12497,N_13412);
xnor UO_1922 (O_1922,N_13347,N_12510);
xnor UO_1923 (O_1923,N_12506,N_12318);
and UO_1924 (O_1924,N_13755,N_12530);
and UO_1925 (O_1925,N_14517,N_12945);
and UO_1926 (O_1926,N_13836,N_13721);
and UO_1927 (O_1927,N_13846,N_13824);
and UO_1928 (O_1928,N_12179,N_12589);
or UO_1929 (O_1929,N_14255,N_12785);
nor UO_1930 (O_1930,N_13213,N_12330);
or UO_1931 (O_1931,N_14569,N_12772);
nor UO_1932 (O_1932,N_14789,N_12781);
or UO_1933 (O_1933,N_14004,N_14084);
nor UO_1934 (O_1934,N_12827,N_13348);
xor UO_1935 (O_1935,N_13344,N_12369);
or UO_1936 (O_1936,N_14671,N_12761);
xor UO_1937 (O_1937,N_14431,N_13600);
xnor UO_1938 (O_1938,N_14432,N_14628);
xor UO_1939 (O_1939,N_12517,N_14736);
xnor UO_1940 (O_1940,N_13856,N_13467);
and UO_1941 (O_1941,N_12268,N_14875);
or UO_1942 (O_1942,N_12114,N_14978);
or UO_1943 (O_1943,N_13753,N_13215);
and UO_1944 (O_1944,N_12986,N_13420);
nand UO_1945 (O_1945,N_12409,N_13391);
or UO_1946 (O_1946,N_13938,N_14759);
and UO_1947 (O_1947,N_13814,N_12422);
xnor UO_1948 (O_1948,N_13827,N_13423);
nand UO_1949 (O_1949,N_12331,N_13548);
or UO_1950 (O_1950,N_13965,N_12417);
or UO_1951 (O_1951,N_14952,N_14045);
or UO_1952 (O_1952,N_13072,N_14380);
or UO_1953 (O_1953,N_12968,N_14095);
and UO_1954 (O_1954,N_14000,N_14552);
xor UO_1955 (O_1955,N_12272,N_13627);
xnor UO_1956 (O_1956,N_12985,N_13453);
nand UO_1957 (O_1957,N_12229,N_14571);
and UO_1958 (O_1958,N_13284,N_14987);
and UO_1959 (O_1959,N_14358,N_13491);
xnor UO_1960 (O_1960,N_12214,N_12757);
and UO_1961 (O_1961,N_13363,N_13093);
or UO_1962 (O_1962,N_13131,N_12418);
or UO_1963 (O_1963,N_12420,N_13462);
and UO_1964 (O_1964,N_12804,N_14069);
or UO_1965 (O_1965,N_13120,N_13228);
xnor UO_1966 (O_1966,N_14087,N_14999);
nand UO_1967 (O_1967,N_14525,N_14087);
and UO_1968 (O_1968,N_14704,N_13965);
nor UO_1969 (O_1969,N_14325,N_14547);
or UO_1970 (O_1970,N_14774,N_12199);
and UO_1971 (O_1971,N_14874,N_13767);
nor UO_1972 (O_1972,N_13321,N_13491);
nor UO_1973 (O_1973,N_12967,N_13564);
xnor UO_1974 (O_1974,N_14703,N_14149);
xor UO_1975 (O_1975,N_12595,N_13921);
nor UO_1976 (O_1976,N_14098,N_12821);
nor UO_1977 (O_1977,N_13127,N_12007);
xnor UO_1978 (O_1978,N_13402,N_14110);
and UO_1979 (O_1979,N_14668,N_13364);
or UO_1980 (O_1980,N_13818,N_14176);
nor UO_1981 (O_1981,N_14731,N_14063);
xor UO_1982 (O_1982,N_14469,N_14546);
xor UO_1983 (O_1983,N_13870,N_13224);
xnor UO_1984 (O_1984,N_14665,N_13477);
xnor UO_1985 (O_1985,N_12946,N_14875);
nand UO_1986 (O_1986,N_12081,N_13307);
nand UO_1987 (O_1987,N_12278,N_14871);
or UO_1988 (O_1988,N_12396,N_13782);
and UO_1989 (O_1989,N_14938,N_13533);
nor UO_1990 (O_1990,N_13272,N_12478);
nor UO_1991 (O_1991,N_13182,N_12929);
xor UO_1992 (O_1992,N_12303,N_13833);
xnor UO_1993 (O_1993,N_14628,N_14454);
xor UO_1994 (O_1994,N_13994,N_12522);
and UO_1995 (O_1995,N_13376,N_13469);
xor UO_1996 (O_1996,N_13041,N_13702);
nor UO_1997 (O_1997,N_12284,N_12625);
and UO_1998 (O_1998,N_13953,N_12606);
or UO_1999 (O_1999,N_12965,N_14400);
endmodule