module basic_2500_25000_3000_10_levels_5xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
nor U0 (N_0,In_1118,In_416);
or U1 (N_1,In_1114,In_1812);
nand U2 (N_2,In_1699,In_2424);
nor U3 (N_3,In_1564,In_1456);
or U4 (N_4,In_1794,In_755);
nor U5 (N_5,In_2190,In_2053);
and U6 (N_6,In_502,In_596);
nor U7 (N_7,In_268,In_429);
nor U8 (N_8,In_967,In_1679);
or U9 (N_9,In_537,In_506);
nand U10 (N_10,In_911,In_2057);
nor U11 (N_11,In_1582,In_2295);
nand U12 (N_12,In_1144,In_783);
and U13 (N_13,In_585,In_1662);
nor U14 (N_14,In_1408,In_570);
nor U15 (N_15,In_1871,In_970);
and U16 (N_16,In_568,In_30);
nor U17 (N_17,In_2299,In_2391);
nor U18 (N_18,In_533,In_554);
nand U19 (N_19,In_224,In_255);
or U20 (N_20,In_2138,In_1826);
or U21 (N_21,In_1062,In_808);
nor U22 (N_22,In_751,In_2064);
and U23 (N_23,In_2346,In_857);
or U24 (N_24,In_275,In_689);
nand U25 (N_25,In_158,In_241);
xnor U26 (N_26,In_192,In_1804);
nor U27 (N_27,In_1563,In_1148);
nor U28 (N_28,In_1467,In_1844);
or U29 (N_29,In_398,In_238);
or U30 (N_30,In_1536,In_1676);
nor U31 (N_31,In_166,In_627);
nor U32 (N_32,In_2278,In_1483);
or U33 (N_33,In_344,In_648);
nand U34 (N_34,In_61,In_2326);
and U35 (N_35,In_2469,In_1675);
or U36 (N_36,In_1103,In_744);
or U37 (N_37,In_2217,In_2117);
nand U38 (N_38,In_769,In_991);
nor U39 (N_39,In_2102,In_280);
or U40 (N_40,In_1452,In_287);
nand U41 (N_41,In_1228,In_993);
nor U42 (N_42,In_2353,In_294);
nand U43 (N_43,In_274,In_386);
or U44 (N_44,In_1460,In_408);
xor U45 (N_45,In_1601,In_1386);
nand U46 (N_46,In_181,In_1901);
nand U47 (N_47,In_367,In_950);
nand U48 (N_48,In_2001,In_1082);
nor U49 (N_49,In_578,In_413);
nor U50 (N_50,In_1323,In_361);
xor U51 (N_51,In_104,In_1372);
nor U52 (N_52,In_433,In_2047);
nand U53 (N_53,In_2262,In_1077);
xor U54 (N_54,In_604,In_851);
nand U55 (N_55,In_440,In_813);
or U56 (N_56,In_197,In_2071);
or U57 (N_57,In_2442,In_904);
nand U58 (N_58,In_1809,In_2386);
or U59 (N_59,In_1501,In_853);
or U60 (N_60,In_544,In_52);
nand U61 (N_61,In_639,In_2192);
nor U62 (N_62,In_491,In_1015);
and U63 (N_63,In_592,In_2499);
or U64 (N_64,In_2125,In_1146);
and U65 (N_65,In_2062,In_1224);
or U66 (N_66,In_373,In_2183);
and U67 (N_67,In_757,In_272);
nand U68 (N_68,In_459,In_1576);
or U69 (N_69,In_1722,In_2477);
or U70 (N_70,In_2006,In_2007);
xor U71 (N_71,In_2449,In_1530);
or U72 (N_72,In_1936,In_80);
nor U73 (N_73,In_850,In_27);
nor U74 (N_74,In_362,In_1924);
nor U75 (N_75,In_2033,In_2372);
nor U76 (N_76,In_2294,In_1898);
or U77 (N_77,In_636,In_1332);
nand U78 (N_78,In_2093,In_1657);
nor U79 (N_79,In_2446,In_2286);
or U80 (N_80,In_2384,In_2281);
nand U81 (N_81,In_267,In_1014);
nand U82 (N_82,In_436,In_2152);
and U83 (N_83,In_253,In_1);
nor U84 (N_84,In_1199,In_2454);
or U85 (N_85,In_1239,In_1990);
and U86 (N_86,In_133,In_256);
nor U87 (N_87,In_2284,In_624);
or U88 (N_88,In_1234,In_1738);
nor U89 (N_89,In_726,In_2277);
and U90 (N_90,In_1375,In_2336);
xnor U91 (N_91,In_2272,In_1207);
nand U92 (N_92,In_1002,In_1472);
or U93 (N_93,In_1449,In_244);
nor U94 (N_94,In_1714,In_2309);
and U95 (N_95,In_269,In_2388);
and U96 (N_96,In_1208,In_1997);
nand U97 (N_97,In_1238,In_2396);
nor U98 (N_98,In_1448,In_883);
nand U99 (N_99,In_2400,In_1878);
nor U100 (N_100,In_2123,In_1379);
and U101 (N_101,In_1399,In_1130);
nor U102 (N_102,In_358,In_737);
nor U103 (N_103,In_1250,In_637);
nor U104 (N_104,In_1097,In_829);
nand U105 (N_105,In_2169,In_2279);
nand U106 (N_106,In_1565,In_750);
xnor U107 (N_107,In_1293,In_2034);
nor U108 (N_108,In_1435,In_2359);
or U109 (N_109,In_2099,In_2023);
nor U110 (N_110,In_305,In_1227);
nor U111 (N_111,In_2362,In_1217);
xnor U112 (N_112,In_1249,In_277);
xor U113 (N_113,In_558,In_1173);
nor U114 (N_114,In_1661,In_2214);
nor U115 (N_115,In_380,In_1696);
xor U116 (N_116,In_780,In_487);
or U117 (N_117,In_410,In_577);
nand U118 (N_118,In_1307,In_2110);
or U119 (N_119,In_1761,In_1656);
and U120 (N_120,In_1628,In_526);
xnor U121 (N_121,In_308,In_1469);
and U122 (N_122,In_1065,In_708);
or U123 (N_123,In_259,In_1621);
nor U124 (N_124,In_1337,In_196);
nor U125 (N_125,In_70,In_2076);
nor U126 (N_126,In_620,In_2453);
and U127 (N_127,In_1038,In_67);
or U128 (N_128,In_1382,In_1504);
xor U129 (N_129,In_1949,In_836);
or U130 (N_130,In_1063,In_388);
xor U131 (N_131,In_1300,In_2228);
or U132 (N_132,In_1478,In_151);
xnor U133 (N_133,In_250,In_2283);
nor U134 (N_134,In_1983,In_2486);
nand U135 (N_135,In_1213,In_34);
nor U136 (N_136,In_1919,In_1795);
nor U137 (N_137,In_1683,In_1996);
and U138 (N_138,In_296,In_975);
and U139 (N_139,In_679,In_276);
nor U140 (N_140,In_1098,In_1974);
xnor U141 (N_141,In_1183,In_842);
nor U142 (N_142,In_111,In_715);
and U143 (N_143,In_1774,In_1653);
nor U144 (N_144,In_1368,In_317);
and U145 (N_145,In_573,In_1182);
or U146 (N_146,In_1432,In_306);
or U147 (N_147,In_472,In_2221);
nor U148 (N_148,In_1736,In_13);
nor U149 (N_149,In_1214,In_1269);
and U150 (N_150,In_1578,In_49);
or U151 (N_151,In_2105,In_858);
nand U152 (N_152,In_763,In_2095);
nand U153 (N_153,In_157,In_2434);
or U154 (N_154,In_616,In_201);
nand U155 (N_155,In_411,In_1988);
and U156 (N_156,In_374,In_1150);
or U157 (N_157,In_1111,In_2098);
nor U158 (N_158,In_873,In_610);
xor U159 (N_159,In_2307,In_234);
nand U160 (N_160,In_1244,In_939);
and U161 (N_161,In_901,In_2244);
nor U162 (N_162,In_2136,In_476);
xnor U163 (N_163,In_1003,In_442);
xnor U164 (N_164,In_35,In_1594);
nand U165 (N_165,In_1407,In_1781);
nand U166 (N_166,In_657,In_579);
and U167 (N_167,In_886,In_2412);
nand U168 (N_168,In_2389,In_1821);
and U169 (N_169,In_712,In_915);
nor U170 (N_170,In_2259,In_177);
nand U171 (N_171,In_1485,In_134);
nand U172 (N_172,In_1907,In_371);
xnor U173 (N_173,In_36,In_2418);
and U174 (N_174,In_147,In_1700);
and U175 (N_175,In_123,In_1680);
xnor U176 (N_176,In_717,In_2414);
nand U177 (N_177,In_795,In_1664);
nor U178 (N_178,In_2457,In_1330);
or U179 (N_179,In_927,In_1768);
nand U180 (N_180,In_703,In_840);
or U181 (N_181,In_1954,In_72);
and U182 (N_182,In_1817,In_926);
and U183 (N_183,In_1885,In_1253);
or U184 (N_184,In_1721,In_1490);
nand U185 (N_185,In_377,In_81);
and U186 (N_186,In_891,In_1906);
and U187 (N_187,In_1868,In_525);
or U188 (N_188,In_1393,In_711);
nor U189 (N_189,In_95,In_527);
nand U190 (N_190,In_1373,In_800);
nand U191 (N_191,In_1270,In_879);
nor U192 (N_192,In_2492,In_1987);
nor U193 (N_193,In_190,In_1273);
nand U194 (N_194,In_1262,In_794);
nor U195 (N_195,In_1569,In_1566);
nor U196 (N_196,In_141,In_1808);
nand U197 (N_197,In_1806,In_1494);
nand U198 (N_198,In_530,In_2364);
and U199 (N_199,In_687,In_1415);
and U200 (N_200,In_2480,In_540);
nand U201 (N_201,In_496,In_1554);
nor U202 (N_202,In_793,In_2276);
nand U203 (N_203,In_1994,In_1685);
and U204 (N_204,In_435,In_2288);
xnor U205 (N_205,In_1004,In_2489);
or U206 (N_206,In_1682,In_1663);
and U207 (N_207,In_1265,In_1887);
nor U208 (N_208,In_273,In_1650);
and U209 (N_209,In_1807,In_206);
nor U210 (N_210,In_194,In_1541);
nor U211 (N_211,In_2014,In_2111);
nor U212 (N_212,In_1986,In_1836);
nand U213 (N_213,In_167,In_1880);
and U214 (N_214,In_1294,In_2450);
nand U215 (N_215,In_567,In_1785);
nand U216 (N_216,In_816,In_292);
nor U217 (N_217,In_2074,In_1588);
nand U218 (N_218,In_528,In_1903);
and U219 (N_219,In_2328,In_2160);
nor U220 (N_220,In_548,In_90);
nand U221 (N_221,In_1652,In_2493);
or U222 (N_222,In_1403,In_1544);
nand U223 (N_223,In_1391,In_2425);
or U224 (N_224,In_187,In_1838);
nor U225 (N_225,In_1215,In_576);
and U226 (N_226,In_2205,In_1600);
and U227 (N_227,In_1510,In_835);
nor U228 (N_228,In_2091,In_1428);
nand U229 (N_229,In_503,In_565);
or U230 (N_230,In_881,In_1922);
xnor U231 (N_231,In_178,In_588);
xnor U232 (N_232,In_2049,In_2464);
nand U233 (N_233,In_1477,In_401);
and U234 (N_234,In_675,In_14);
nand U235 (N_235,In_1025,In_2269);
and U236 (N_236,In_59,In_659);
or U237 (N_237,In_1728,In_217);
xor U238 (N_238,In_647,In_2432);
or U239 (N_239,In_803,In_1989);
or U240 (N_240,In_1669,In_2306);
nor U241 (N_241,In_907,In_1952);
nor U242 (N_242,In_2310,In_339);
nor U243 (N_243,In_71,In_2227);
nand U244 (N_244,In_784,In_1513);
nand U245 (N_245,In_895,In_1170);
and U246 (N_246,In_2089,In_1048);
xnor U247 (N_247,In_2218,In_204);
or U248 (N_248,In_311,In_1495);
or U249 (N_249,In_428,In_1869);
or U250 (N_250,In_1445,In_841);
or U251 (N_251,In_446,In_1316);
or U252 (N_252,In_2246,In_2041);
and U253 (N_253,In_210,In_329);
and U254 (N_254,In_1101,In_2422);
and U255 (N_255,In_1404,In_1387);
nand U256 (N_256,In_266,In_600);
or U257 (N_257,In_22,In_1427);
nor U258 (N_258,In_1525,In_254);
nand U259 (N_259,In_1848,In_1290);
and U260 (N_260,In_2251,In_1859);
and U261 (N_261,In_1532,In_1455);
and U262 (N_262,In_366,In_1672);
or U263 (N_263,In_1678,In_2213);
and U264 (N_264,In_1166,In_326);
and U265 (N_265,In_1789,In_1094);
nand U266 (N_266,In_2385,In_1598);
and U267 (N_267,In_38,In_1967);
xor U268 (N_268,In_1295,In_2050);
and U269 (N_269,In_1342,In_370);
xor U270 (N_270,In_1202,In_766);
nand U271 (N_271,In_1610,In_1458);
xor U272 (N_272,In_82,In_231);
or U273 (N_273,In_2380,In_710);
or U274 (N_274,In_1646,In_574);
and U275 (N_275,In_1523,In_2456);
and U276 (N_276,In_43,In_1134);
nand U277 (N_277,In_729,In_1557);
nand U278 (N_278,In_1626,In_124);
nor U279 (N_279,In_1897,In_1831);
nor U280 (N_280,In_348,In_2265);
nor U281 (N_281,In_1964,In_245);
nand U282 (N_282,In_1059,In_1767);
and U283 (N_283,In_2255,In_1645);
nand U284 (N_284,In_1978,In_2161);
and U285 (N_285,In_1298,In_1210);
and U286 (N_286,In_1963,In_168);
nand U287 (N_287,In_1279,In_477);
nand U288 (N_288,In_466,In_91);
nor U289 (N_289,In_84,In_1629);
nor U290 (N_290,In_1140,In_1374);
or U291 (N_291,In_2333,In_1322);
nand U292 (N_292,In_1827,In_922);
nor U293 (N_293,In_660,In_1890);
and U294 (N_294,In_1036,In_559);
or U295 (N_295,In_2484,In_867);
nand U296 (N_296,In_1231,In_6);
and U297 (N_297,In_1151,In_1357);
nor U298 (N_298,In_1479,In_137);
and U299 (N_299,In_58,In_1046);
nor U300 (N_300,In_1092,In_2379);
nor U301 (N_301,In_1260,In_174);
and U302 (N_302,In_1892,In_1266);
nor U303 (N_303,In_847,In_2168);
xor U304 (N_304,In_1198,In_498);
and U305 (N_305,In_1017,In_1693);
or U306 (N_306,In_332,In_1889);
or U307 (N_307,In_2285,In_789);
nand U308 (N_308,In_223,In_623);
nand U309 (N_309,In_962,In_475);
and U310 (N_310,In_790,In_2035);
nand U311 (N_311,In_2229,In_66);
nor U312 (N_312,In_1232,In_488);
nand U313 (N_313,In_334,In_243);
and U314 (N_314,In_644,In_2483);
nand U315 (N_315,In_731,In_1287);
nor U316 (N_316,In_412,In_2417);
nor U317 (N_317,In_979,In_382);
or U318 (N_318,In_1715,In_2462);
or U319 (N_319,In_892,In_2323);
and U320 (N_320,In_323,In_233);
and U321 (N_321,In_1691,In_2438);
or U322 (N_322,In_1457,In_1546);
and U323 (N_323,In_1481,In_2458);
and U324 (N_324,In_493,In_2239);
xor U325 (N_325,In_112,In_2381);
nand U326 (N_326,In_365,In_291);
xnor U327 (N_327,In_1591,In_299);
nor U328 (N_328,In_1087,In_2476);
nor U329 (N_329,In_953,In_1473);
nor U330 (N_330,In_607,In_1786);
xnor U331 (N_331,In_2119,In_1589);
nand U332 (N_332,In_1982,In_1943);
nor U333 (N_333,In_692,In_1620);
nor U334 (N_334,In_2191,In_664);
nand U335 (N_335,In_2000,In_806);
nand U336 (N_336,In_100,In_2487);
nand U337 (N_337,In_129,In_1158);
nor U338 (N_338,In_239,In_987);
nand U339 (N_339,In_102,In_1815);
and U340 (N_340,In_2497,In_745);
or U341 (N_341,In_2009,In_1074);
nand U342 (N_342,In_2366,In_1751);
nand U343 (N_343,In_1820,In_2070);
nor U344 (N_344,In_2056,In_1181);
or U345 (N_345,In_2471,In_1008);
or U346 (N_346,In_768,In_2357);
and U347 (N_347,In_1431,In_1032);
or U348 (N_348,In_1798,In_1968);
and U349 (N_349,In_357,In_2025);
nor U350 (N_350,In_1649,In_738);
or U351 (N_351,In_2491,In_1306);
xor U352 (N_352,In_749,In_782);
nor U353 (N_353,In_1753,In_593);
and U354 (N_354,In_2097,In_517);
or U355 (N_355,In_1367,In_1389);
nor U356 (N_356,In_106,In_1673);
or U357 (N_357,In_1475,In_1519);
nand U358 (N_358,In_1313,In_1430);
and U359 (N_359,In_1631,In_1258);
nor U360 (N_360,In_1778,In_2167);
nand U361 (N_361,In_2054,In_2201);
or U362 (N_362,In_747,In_676);
nand U363 (N_363,In_566,In_1230);
or U364 (N_364,In_2066,In_1618);
or U365 (N_365,In_897,In_1980);
or U366 (N_366,In_2126,In_1770);
or U367 (N_367,In_369,In_638);
xnor U368 (N_368,In_1297,In_2081);
or U369 (N_369,In_1834,In_1052);
nor U370 (N_370,In_1701,In_1528);
or U371 (N_371,In_2027,In_810);
and U372 (N_372,In_1762,In_471);
nand U373 (N_373,In_2003,In_1910);
nor U374 (N_374,In_1507,In_824);
and U375 (N_375,In_958,In_1694);
nand U376 (N_376,In_1927,In_48);
and U377 (N_377,In_595,In_2116);
xnor U378 (N_378,In_760,In_1965);
and U379 (N_379,In_336,In_1969);
or U380 (N_380,In_26,In_1086);
xnor U381 (N_381,In_1687,In_1886);
nor U382 (N_382,In_1744,In_295);
and U383 (N_383,In_246,In_1168);
nand U384 (N_384,In_191,In_748);
nor U385 (N_385,In_462,In_1291);
and U386 (N_386,In_919,In_603);
and U387 (N_387,In_2065,In_700);
nand U388 (N_388,In_1587,In_2202);
or U389 (N_389,In_2315,In_545);
xnor U390 (N_390,In_85,In_916);
nor U391 (N_391,In_150,In_2382);
nand U392 (N_392,In_1951,In_118);
and U393 (N_393,In_438,In_2236);
nand U394 (N_394,In_684,In_47);
or U395 (N_395,In_2036,In_2475);
nor U396 (N_396,In_1309,In_896);
nor U397 (N_397,In_89,In_889);
nor U398 (N_398,In_2005,In_667);
or U399 (N_399,In_1212,In_2094);
nand U400 (N_400,In_1275,In_1724);
and U401 (N_401,In_165,In_1196);
nor U402 (N_402,In_302,In_1139);
or U403 (N_403,In_832,In_1000);
or U404 (N_404,In_1613,In_1045);
xnor U405 (N_405,In_2242,In_1350);
nand U406 (N_406,In_826,In_467);
and U407 (N_407,In_218,In_449);
xor U408 (N_408,In_316,In_184);
and U409 (N_409,In_2485,In_2247);
nand U410 (N_410,In_57,In_2208);
nor U411 (N_411,In_1902,In_1850);
or U412 (N_412,In_2447,In_2374);
or U413 (N_413,In_2122,In_955);
and U414 (N_414,In_2332,In_3);
nand U415 (N_415,In_1125,In_1156);
and U416 (N_416,In_1285,In_2189);
nor U417 (N_417,In_343,In_289);
nor U418 (N_418,In_680,In_1264);
xor U419 (N_419,In_2340,In_1200);
and U420 (N_420,In_1896,In_2437);
nand U421 (N_421,In_222,In_868);
and U422 (N_422,In_1705,In_482);
nand U423 (N_423,In_779,In_2423);
or U424 (N_424,In_1338,In_2107);
nand U425 (N_425,In_930,In_354);
and U426 (N_426,In_2377,In_1937);
nand U427 (N_427,In_2029,In_1899);
and U428 (N_428,In_240,In_2134);
and U429 (N_429,In_1042,In_1740);
nor U430 (N_430,In_2378,In_1348);
and U431 (N_431,In_913,In_2271);
xor U432 (N_432,In_1935,In_2182);
and U433 (N_433,In_2352,In_1341);
xnor U434 (N_434,In_1846,In_1075);
nand U435 (N_435,In_172,In_655);
nor U436 (N_436,In_1378,In_2226);
and U437 (N_437,In_1559,In_1277);
and U438 (N_438,In_1873,In_1602);
or U439 (N_439,In_894,In_481);
and U440 (N_440,In_2390,In_2211);
nand U441 (N_441,In_115,In_2143);
and U442 (N_442,In_282,In_1520);
nand U443 (N_443,In_1141,In_805);
or U444 (N_444,In_945,In_1135);
and U445 (N_445,In_846,In_531);
nand U446 (N_446,In_934,In_2282);
and U447 (N_447,In_1057,In_1888);
nand U448 (N_448,In_1426,In_1604);
or U449 (N_449,In_8,In_621);
and U450 (N_450,In_468,In_1521);
or U451 (N_451,In_929,In_1671);
xor U452 (N_452,In_772,In_1344);
or U453 (N_453,In_2341,In_1115);
or U454 (N_454,In_2090,In_2488);
nor U455 (N_455,In_2124,In_1371);
nor U456 (N_456,In_2348,In_1369);
and U457 (N_457,In_265,In_1073);
xnor U458 (N_458,In_418,In_1558);
and U459 (N_459,In_1962,In_387);
nor U460 (N_460,In_866,In_1484);
and U461 (N_461,In_54,In_1875);
or U462 (N_462,In_843,In_582);
nor U463 (N_463,In_1654,In_1939);
nor U464 (N_464,In_1787,In_2360);
xor U465 (N_465,In_226,In_1777);
xnor U466 (N_466,In_1047,In_2319);
nor U467 (N_467,In_2305,In_562);
nor U468 (N_468,In_2210,In_1284);
nand U469 (N_469,In_1858,In_490);
nor U470 (N_470,In_791,In_335);
nor U471 (N_471,In_2067,In_640);
and U472 (N_472,In_415,In_2460);
and U473 (N_473,In_1051,In_1425);
nor U474 (N_474,In_469,In_1319);
nand U475 (N_475,In_2403,In_855);
and U476 (N_476,In_538,In_1766);
or U477 (N_477,In_88,In_1992);
or U478 (N_478,In_1058,In_1184);
or U479 (N_479,In_1211,In_252);
and U480 (N_480,In_862,In_1945);
and U481 (N_481,In_1776,In_149);
nand U482 (N_482,In_1677,In_1792);
or U483 (N_483,In_1934,In_63);
nand U484 (N_484,In_1105,In_2237);
xnor U485 (N_485,In_678,In_138);
nand U486 (N_486,In_143,In_1499);
or U487 (N_487,In_126,In_536);
nand U488 (N_488,In_1138,In_1551);
nor U489 (N_489,In_2154,In_876);
and U490 (N_490,In_767,In_1019);
nor U491 (N_491,In_2465,In_1735);
nand U492 (N_492,In_2174,In_1667);
xnor U493 (N_493,In_227,In_2101);
nand U494 (N_494,In_1424,In_912);
or U495 (N_495,In_1511,In_2164);
nor U496 (N_496,In_1153,In_812);
or U497 (N_497,In_765,In_1923);
nand U498 (N_498,In_2399,In_2235);
nor U499 (N_499,In_1802,In_125);
nor U500 (N_500,In_1957,In_818);
nand U501 (N_501,In_445,In_1966);
and U502 (N_502,In_423,In_98);
nor U503 (N_503,In_698,In_1380);
and U504 (N_504,In_198,In_1145);
or U505 (N_505,In_2397,In_1276);
nand U506 (N_506,In_170,In_1644);
and U507 (N_507,In_448,In_1328);
nor U508 (N_508,In_699,In_1418);
nor U509 (N_509,In_2401,In_480);
and U510 (N_510,In_457,In_686);
or U511 (N_511,In_1692,In_1837);
nor U512 (N_512,In_941,In_833);
or U513 (N_513,In_541,In_2061);
or U514 (N_514,In_1007,In_1849);
xnor U515 (N_515,In_509,In_1854);
nand U516 (N_516,In_279,In_515);
nor U517 (N_517,In_696,In_505);
or U518 (N_518,In_1535,In_909);
or U519 (N_519,In_969,In_893);
or U520 (N_520,In_1959,In_1717);
nor U521 (N_521,In_1155,In_1233);
nor U522 (N_522,In_2429,In_2274);
nand U523 (N_523,In_914,In_706);
nand U524 (N_524,In_1642,In_1979);
or U525 (N_525,In_212,In_1027);
nor U526 (N_526,In_2215,In_1188);
and U527 (N_527,In_2494,In_984);
xnor U528 (N_528,In_2075,In_2017);
xor U529 (N_529,In_1084,In_1660);
nand U530 (N_530,In_1863,In_632);
and U531 (N_531,In_1526,In_2083);
nor U532 (N_532,In_1496,In_670);
nor U533 (N_533,In_2142,In_1572);
nor U534 (N_534,In_2149,In_2445);
xor U535 (N_535,In_1303,In_653);
xor U536 (N_536,In_2369,In_630);
or U537 (N_537,In_1608,In_2495);
or U538 (N_538,In_1471,In_397);
nand U539 (N_539,In_546,In_330);
nor U540 (N_540,In_2051,In_1248);
nand U541 (N_541,In_1719,In_383);
or U542 (N_542,In_1716,In_1900);
or U543 (N_543,In_1944,In_2166);
and U544 (N_544,In_142,In_1772);
nand U545 (N_545,In_2461,In_203);
or U546 (N_546,In_1197,In_2459);
or U547 (N_547,In_671,In_580);
or U548 (N_548,In_2141,In_1235);
nand U549 (N_549,In_1189,In_1491);
or U550 (N_550,In_1615,In_1593);
or U551 (N_551,In_718,In_1339);
and U552 (N_552,In_1162,In_1548);
and U553 (N_553,In_1121,In_441);
or U554 (N_554,In_7,In_781);
nand U555 (N_555,In_1024,In_1315);
nor U556 (N_556,In_626,In_1713);
nand U557 (N_557,In_978,In_734);
xnor U558 (N_558,In_1710,In_1131);
xor U559 (N_559,In_1750,In_1940);
nor U560 (N_560,In_1033,In_2024);
nor U561 (N_561,In_2371,In_1972);
xnor U562 (N_562,In_4,In_1123);
or U563 (N_563,In_2108,In_1128);
and U564 (N_564,In_1816,In_854);
xor U565 (N_565,In_2304,In_1670);
nor U566 (N_566,In_1078,In_1261);
nand U567 (N_567,In_2347,In_2343);
nand U568 (N_568,In_645,In_838);
xnor U569 (N_569,In_823,In_649);
nand U570 (N_570,In_673,In_654);
nand U571 (N_571,In_2433,In_1413);
and U572 (N_572,In_2203,In_611);
or U573 (N_573,In_792,In_2022);
nand U574 (N_574,In_2128,In_2406);
xnor U575 (N_575,In_1814,In_1622);
and U576 (N_576,In_1414,In_2018);
nand U577 (N_577,In_739,In_1028);
nand U578 (N_578,In_628,In_614);
nand U579 (N_579,In_510,In_553);
and U580 (N_580,In_1852,In_2151);
nand U581 (N_581,In_961,In_2361);
or U582 (N_582,In_622,In_1113);
nor U583 (N_583,In_2129,In_1366);
and U584 (N_584,In_798,In_285);
and U585 (N_585,In_1818,In_404);
and U586 (N_586,In_1085,In_2021);
nor U587 (N_587,In_309,In_152);
and U588 (N_588,In_2132,In_450);
nor U589 (N_589,In_1447,In_1577);
xor U590 (N_590,In_10,In_730);
and U591 (N_591,In_248,In_29);
nand U592 (N_592,In_1488,In_1246);
nor U593 (N_593,In_1124,In_2498);
or U594 (N_594,In_427,In_392);
or U595 (N_595,In_2220,In_1866);
nand U596 (N_596,In_31,In_2028);
or U597 (N_597,In_1606,In_1882);
xnor U598 (N_598,In_1788,In_1872);
and U599 (N_599,In_2197,In_1707);
xnor U600 (N_600,In_1474,In_2039);
nand U601 (N_601,In_1185,In_396);
or U602 (N_602,In_727,In_924);
nor U603 (N_603,In_1981,In_740);
nand U604 (N_604,In_1851,In_495);
nor U605 (N_605,In_2478,In_2118);
nand U606 (N_606,In_188,In_1267);
or U607 (N_607,In_145,In_2426);
or U608 (N_608,In_2430,In_403);
nand U609 (N_609,In_483,In_860);
nand U610 (N_610,In_1651,In_463);
nand U611 (N_611,In_1026,In_68);
and U612 (N_612,In_2207,In_92);
xnor U613 (N_613,In_561,In_1975);
nor U614 (N_614,In_590,In_1632);
xor U615 (N_615,In_1659,In_669);
nand U616 (N_616,In_589,In_107);
nor U617 (N_617,In_557,In_5);
or U618 (N_618,In_1462,In_2367);
xnor U619 (N_619,In_736,In_1704);
nand U620 (N_620,In_2421,In_931);
or U621 (N_621,In_1929,In_965);
nor U622 (N_622,In_2355,In_284);
nand U623 (N_623,In_1648,In_1783);
nor U624 (N_624,In_1921,In_1305);
nand U625 (N_625,In_1603,In_324);
nand U626 (N_626,In_159,In_825);
nor U627 (N_627,In_584,In_1567);
or U628 (N_628,In_2268,In_1365);
nor U629 (N_629,In_1023,In_724);
nand U630 (N_630,In_1941,In_321);
xnor U631 (N_631,In_923,In_2230);
or U632 (N_632,In_1206,In_2026);
or U633 (N_633,In_874,In_1636);
nor U634 (N_634,In_1773,In_1698);
or U635 (N_635,In_1638,In_2470);
nand U636 (N_636,In_1668,In_127);
nor U637 (N_637,In_1020,In_1219);
nor U638 (N_638,In_1555,In_2144);
nand U639 (N_639,In_1920,In_1742);
or U640 (N_640,In_186,In_2114);
nand U641 (N_641,In_1089,In_349);
or U642 (N_642,In_1720,In_185);
nand U643 (N_643,In_1394,In_1829);
xor U644 (N_644,In_345,In_2296);
nand U645 (N_645,In_2209,In_1072);
xor U646 (N_646,In_944,In_802);
nand U647 (N_647,In_1596,In_28);
nand U648 (N_648,In_633,In_1973);
xnor U649 (N_649,In_37,In_2335);
and U650 (N_650,In_2216,In_1830);
nand U651 (N_651,In_775,In_1493);
nor U652 (N_652,In_677,In_2302);
xnor U653 (N_653,In_1165,In_1463);
nand U654 (N_654,In_1916,In_2325);
nand U655 (N_655,In_1450,In_1327);
and U656 (N_656,In_391,In_819);
nand U657 (N_657,In_1611,In_451);
or U658 (N_658,In_318,In_1917);
nor U659 (N_659,In_205,In_1116);
nor U660 (N_660,In_1446,In_1406);
or U661 (N_661,In_1503,In_2073);
nor U662 (N_662,In_2139,In_2320);
and U663 (N_663,In_301,In_1018);
xor U664 (N_664,In_148,In_473);
or U665 (N_665,In_1529,In_434);
or U666 (N_666,In_988,In_17);
nand U667 (N_667,In_1946,In_2212);
and U668 (N_668,In_656,In_946);
nor U669 (N_669,In_2416,In_1860);
nand U670 (N_670,In_839,In_132);
nand U671 (N_671,In_2427,In_1580);
nand U672 (N_672,In_1272,In_1175);
or U673 (N_673,In_733,In_350);
nand U674 (N_674,In_863,In_2474);
or U675 (N_675,In_720,In_2313);
or U676 (N_676,In_776,In_864);
nand U677 (N_677,In_372,In_1392);
and U678 (N_678,In_756,In_2087);
or U679 (N_679,In_1152,In_163);
or U680 (N_680,In_2200,In_2435);
xor U681 (N_681,In_1090,In_1022);
xor U682 (N_682,In_2156,In_709);
and U683 (N_683,In_572,In_641);
and U684 (N_684,In_2109,In_1088);
and U685 (N_685,In_1254,In_1204);
nor U686 (N_686,In_1695,In_417);
nor U687 (N_687,In_2339,In_534);
and U688 (N_688,In_105,In_1746);
nand U689 (N_689,In_1358,In_1542);
or U690 (N_690,In_2231,In_690);
and U691 (N_691,In_1711,In_114);
or U692 (N_692,In_1739,In_1451);
nand U693 (N_693,In_431,In_1352);
and U694 (N_694,In_208,In_1302);
or U695 (N_695,In_1537,In_966);
or U696 (N_696,In_651,In_2222);
nor U697 (N_697,In_1531,In_591);
or U698 (N_698,In_615,In_2481);
nor U699 (N_699,In_1274,In_65);
and U700 (N_700,In_1609,In_1955);
or U701 (N_701,In_1703,In_2356);
and U702 (N_702,In_2238,In_2292);
and U703 (N_703,In_1221,In_1370);
xnor U704 (N_704,In_214,In_1257);
or U705 (N_705,In_1381,In_1799);
or U706 (N_706,In_424,In_1349);
nand U707 (N_707,In_1666,In_2052);
nor U708 (N_708,In_156,In_880);
nand U709 (N_709,In_53,In_774);
nor U710 (N_710,In_2206,In_1833);
and U711 (N_711,In_2198,In_1355);
and U712 (N_712,In_164,In_447);
or U713 (N_713,In_247,In_1324);
or U714 (N_714,In_452,In_497);
and U715 (N_715,In_1194,In_2408);
and U716 (N_716,In_986,In_1726);
and U717 (N_717,In_1252,In_146);
or U718 (N_718,In_674,In_56);
and U719 (N_719,In_402,In_16);
nand U720 (N_720,In_2224,In_2318);
or U721 (N_721,In_1522,In_2466);
and U722 (N_722,In_2019,In_455);
nand U723 (N_723,In_1894,In_1747);
and U724 (N_724,In_1035,In_1579);
and U725 (N_725,In_1049,In_1126);
or U726 (N_726,In_2162,In_379);
xnor U727 (N_727,In_1486,In_960);
and U728 (N_728,In_762,In_693);
or U729 (N_729,In_25,In_1926);
nand U730 (N_730,In_1690,In_1112);
nor U731 (N_731,In_281,In_1190);
and U732 (N_732,In_1209,In_815);
nand U733 (N_733,In_2455,In_385);
and U734 (N_734,In_1314,In_327);
nor U735 (N_735,In_2358,In_796);
nor U736 (N_736,In_1730,In_1616);
or U737 (N_737,In_1684,In_1040);
nor U738 (N_738,In_1416,In_2184);
nand U739 (N_739,In_1819,In_11);
and U740 (N_740,In_1803,In_1993);
nor U741 (N_741,In_1304,In_1487);
xnor U742 (N_742,In_2300,In_33);
nor U743 (N_743,In_598,In_1712);
or U744 (N_744,In_1641,In_875);
xnor U745 (N_745,In_236,In_947);
nand U746 (N_746,In_2431,In_2148);
nor U747 (N_747,In_2248,In_1263);
and U748 (N_748,In_229,In_353);
and U749 (N_749,In_207,In_44);
and U750 (N_750,In_980,In_550);
nor U751 (N_751,In_2331,In_837);
and U752 (N_752,In_1737,In_2223);
nand U753 (N_753,In_508,In_1440);
nor U754 (N_754,In_786,In_555);
nand U755 (N_755,In_341,In_682);
or U756 (N_756,In_2140,In_1960);
xor U757 (N_757,In_2303,In_20);
and U758 (N_758,In_1056,In_964);
and U759 (N_759,In_2080,In_342);
nand U760 (N_760,In_337,In_2257);
nand U761 (N_761,In_1255,In_785);
nand U762 (N_762,In_171,In_642);
xnor U763 (N_763,In_1093,In_113);
nand U764 (N_764,In_906,In_2298);
xor U765 (N_765,In_182,In_933);
xnor U766 (N_766,In_900,In_2468);
nand U767 (N_767,In_518,In_869);
or U768 (N_768,In_1482,In_1914);
xnor U769 (N_769,In_1397,In_453);
or U770 (N_770,In_613,In_634);
xor U771 (N_771,In_1010,In_520);
nor U772 (N_772,In_1764,In_1343);
or U773 (N_773,In_1760,In_209);
or U774 (N_774,In_2439,In_261);
xor U775 (N_775,In_2137,In_2293);
or U776 (N_776,In_375,In_1061);
and U777 (N_777,In_2013,In_2443);
or U778 (N_778,In_176,In_1856);
and U779 (N_779,In_552,In_1351);
xnor U780 (N_780,In_771,In_1453);
nand U781 (N_781,In_1067,In_96);
xnor U782 (N_782,In_1731,In_1161);
nor U783 (N_783,In_270,In_230);
xor U784 (N_784,In_1571,In_1154);
nor U785 (N_785,In_1709,In_575);
nor U786 (N_786,In_646,In_2085);
or U787 (N_787,In_1508,In_1396);
nand U788 (N_788,In_2415,In_144);
or U789 (N_789,In_1725,In_605);
and U790 (N_790,In_820,In_959);
xnor U791 (N_791,In_283,In_1741);
and U792 (N_792,In_882,In_97);
or U793 (N_793,In_2405,In_1915);
nor U794 (N_794,In_489,In_405);
and U795 (N_795,In_1755,In_601);
nor U796 (N_796,In_542,In_1122);
nor U797 (N_797,In_1805,In_1060);
and U798 (N_798,In_2349,In_2155);
xnor U799 (N_799,In_722,In_1634);
xnor U800 (N_800,In_688,In_293);
xnor U801 (N_801,In_2146,In_1583);
nand U802 (N_802,In_985,In_2199);
and U803 (N_803,In_618,In_79);
xor U804 (N_804,In_1053,In_1241);
or U805 (N_805,In_1464,In_631);
nand U806 (N_806,In_1064,In_1100);
and U807 (N_807,In_663,In_635);
nand U808 (N_808,In_1395,In_461);
nor U809 (N_809,In_1203,In_691);
and U810 (N_810,In_1647,In_968);
or U811 (N_811,In_1353,In_474);
xor U812 (N_812,In_1334,In_310);
xor U813 (N_813,In_753,In_1665);
or U814 (N_814,In_643,In_1796);
nor U815 (N_815,In_1771,In_136);
xor U816 (N_816,In_352,In_797);
nor U817 (N_817,In_1054,In_2176);
or U818 (N_818,In_972,In_1627);
and U819 (N_819,In_1039,In_2100);
nand U820 (N_820,In_1318,In_1079);
nor U821 (N_821,In_139,In_1842);
nor U822 (N_822,In_390,In_1108);
and U823 (N_823,In_949,In_856);
or U824 (N_824,In_547,In_1133);
and U825 (N_825,In_2338,In_1991);
nand U826 (N_826,In_1727,In_60);
and U827 (N_827,In_2370,In_2096);
nand U828 (N_828,In_407,In_828);
and U829 (N_829,In_1547,In_1434);
nand U830 (N_830,In_1931,In_2241);
or U831 (N_831,In_1441,In_1938);
nand U832 (N_832,In_1470,In_1195);
xor U833 (N_833,In_1752,In_1468);
nand U834 (N_834,In_1005,In_422);
nor U835 (N_835,In_101,In_2350);
and U836 (N_836,In_1825,In_1091);
and U837 (N_837,In_834,In_2258);
or U838 (N_838,In_381,In_764);
or U839 (N_839,In_787,In_376);
nand U840 (N_840,In_921,In_1016);
xor U841 (N_841,In_956,In_938);
nor U842 (N_842,In_2275,In_135);
nand U843 (N_843,In_1590,In_1874);
nand U844 (N_844,In_702,In_2103);
or U845 (N_845,In_1689,In_1617);
and U846 (N_846,In_870,In_2245);
xnor U847 (N_847,In_551,In_2186);
nor U848 (N_848,In_1055,In_1877);
nand U849 (N_849,In_1688,In_1839);
or U850 (N_850,In_2410,In_479);
or U851 (N_851,In_2330,In_2150);
nand U852 (N_852,In_257,In_2344);
xor U853 (N_853,In_1841,In_87);
and U854 (N_854,In_877,In_2181);
or U855 (N_855,In_1127,In_501);
nand U856 (N_856,In_1192,In_258);
and U857 (N_857,In_1186,In_2368);
nor U858 (N_858,In_237,In_2171);
or U859 (N_859,In_770,In_122);
xor U860 (N_860,In_1364,In_903);
nor U861 (N_861,In_1331,In_1534);
or U862 (N_862,In_2072,In_831);
or U863 (N_863,In_1918,In_1797);
nand U864 (N_864,In_1625,In_1999);
or U865 (N_865,In_1614,In_773);
and U866 (N_866,In_990,In_1346);
xor U867 (N_867,In_2172,In_1041);
nand U868 (N_868,In_18,In_905);
xnor U869 (N_869,In_1556,In_2127);
nor U870 (N_870,In_2031,In_23);
and U871 (N_871,In_1813,In_1225);
or U872 (N_872,In_1743,In_951);
or U873 (N_873,In_40,In_1597);
and U874 (N_874,In_179,In_235);
nand U875 (N_875,In_1942,In_865);
and U876 (N_876,In_1009,In_1612);
or U877 (N_877,In_120,In_1220);
xor U878 (N_878,In_777,In_1779);
and U879 (N_879,In_1524,In_346);
or U880 (N_880,In_1256,In_543);
xnor U881 (N_881,In_319,In_1461);
or U882 (N_882,In_2250,In_2145);
or U883 (N_883,In_1623,In_1505);
and U884 (N_884,In_221,In_1769);
xor U885 (N_885,In_2078,In_1681);
or U886 (N_886,In_220,In_2020);
nor U887 (N_887,In_935,In_173);
and U888 (N_888,In_2037,In_2266);
nand U889 (N_889,In_523,In_2496);
and U890 (N_890,In_1037,In_262);
nor U891 (N_891,In_2011,In_1568);
xor U892 (N_892,In_1540,In_2042);
and U893 (N_893,In_1925,In_1268);
nor U894 (N_894,In_697,In_1076);
nand U895 (N_895,In_1466,In_701);
or U896 (N_896,In_2261,In_117);
nand U897 (N_897,In_563,In_355);
or U898 (N_898,In_549,In_602);
nand U899 (N_899,In_499,In_1226);
nor U900 (N_900,In_1905,In_1345);
nand U901 (N_901,In_50,In_811);
nand U902 (N_902,In_2482,In_827);
nor U903 (N_903,In_1282,In_884);
or U904 (N_904,In_1171,In_1066);
nand U905 (N_905,In_1498,In_976);
nor U906 (N_906,In_1405,In_1283);
or U907 (N_907,In_1436,In_2113);
nor U908 (N_908,In_2308,In_2392);
nand U909 (N_909,In_1867,In_606);
nor U910 (N_910,In_1748,In_721);
or U911 (N_911,In_845,In_485);
xnor U912 (N_912,In_2317,In_594);
nand U913 (N_913,In_1706,In_1500);
nand U914 (N_914,In_1801,In_658);
nand U915 (N_915,In_928,In_1947);
and U916 (N_916,In_2351,In_160);
nand U917 (N_917,In_821,In_1518);
and U918 (N_918,In_1732,In_1096);
nor U919 (N_919,In_228,In_2204);
and U920 (N_920,In_571,In_1893);
or U921 (N_921,In_1423,In_1102);
nand U922 (N_922,In_2409,In_608);
and U923 (N_923,In_351,In_581);
nand U924 (N_924,In_1984,In_1635);
xnor U925 (N_925,In_2032,In_2383);
xor U926 (N_926,In_1029,In_1857);
nand U927 (N_927,In_1179,In_2329);
nor U928 (N_928,In_2287,In_1071);
and U929 (N_929,In_2043,In_504);
nor U930 (N_930,In_421,In_1237);
and U931 (N_931,In_426,In_925);
nor U932 (N_932,In_723,In_464);
xnor U933 (N_933,In_957,In_2030);
nor U934 (N_934,In_529,In_619);
or U935 (N_935,In_887,In_1909);
or U936 (N_936,In_1422,In_2069);
and U937 (N_937,In_74,In_494);
xnor U938 (N_938,In_1639,In_1674);
or U939 (N_939,In_297,In_219);
and U940 (N_940,In_2419,In_761);
nand U941 (N_941,In_46,In_1359);
and U942 (N_942,In_2121,In_1281);
xnor U943 (N_943,In_213,In_1976);
and U944 (N_944,In_1081,In_2015);
nor U945 (N_945,In_1958,In_286);
and U946 (N_946,In_2084,In_1506);
xor U947 (N_947,In_492,In_2440);
or U948 (N_948,In_1402,In_2157);
nand U949 (N_949,In_1176,In_1733);
or U950 (N_950,In_1104,In_1044);
and U951 (N_951,In_1354,In_193);
xor U952 (N_952,In_1780,In_859);
and U953 (N_953,In_1317,In_338);
xnor U954 (N_954,In_849,In_1749);
and U955 (N_955,In_1296,In_1147);
and U956 (N_956,In_211,In_2158);
nor U957 (N_957,In_460,In_313);
nor U958 (N_958,In_1050,In_1895);
xor U959 (N_959,In_1843,In_2376);
or U960 (N_960,In_719,In_9);
or U961 (N_961,In_1242,In_1259);
nor U962 (N_962,In_1791,In_668);
and U963 (N_963,In_2420,In_1998);
nand U964 (N_964,In_2322,In_300);
or U965 (N_965,In_1340,In_1229);
or U966 (N_966,In_1476,In_2472);
or U967 (N_967,In_1607,In_2280);
and U968 (N_968,In_1883,In_1708);
and U969 (N_969,In_175,In_1163);
or U970 (N_970,In_1001,In_45);
nor U971 (N_971,In_997,In_1411);
nand U972 (N_972,In_1325,In_1509);
or U973 (N_973,In_804,In_333);
nand U974 (N_974,In_822,In_1759);
or U975 (N_975,In_1030,In_1655);
xnor U976 (N_976,In_908,In_1137);
nor U977 (N_977,In_918,In_1110);
xor U978 (N_978,In_569,In_1417);
and U979 (N_979,In_1543,In_131);
nor U980 (N_980,In_1985,In_948);
nand U981 (N_981,In_1658,In_2060);
nand U982 (N_982,In_1553,In_290);
and U983 (N_983,In_216,In_1419);
or U984 (N_984,In_1884,In_1388);
or U985 (N_985,In_1326,In_2402);
and U986 (N_986,In_817,In_564);
or U987 (N_987,In_2411,In_121);
or U988 (N_988,In_512,In_2297);
nand U989 (N_989,In_2187,In_2104);
or U990 (N_990,In_288,In_2314);
and U991 (N_991,In_2086,In_898);
nor U992 (N_992,In_1444,In_2068);
nor U993 (N_993,In_2264,In_249);
and U994 (N_994,In_19,In_456);
nand U995 (N_995,In_2324,In_183);
or U996 (N_996,In_890,In_2301);
nand U997 (N_997,In_532,In_2448);
or U998 (N_998,In_1136,In_2321);
nor U999 (N_999,In_2016,In_1360);
xnor U1000 (N_1000,In_1174,In_1757);
or U1001 (N_1001,In_1119,In_1361);
nor U1002 (N_1002,In_2365,In_524);
or U1003 (N_1003,In_778,In_394);
nand U1004 (N_1004,In_340,In_597);
nor U1005 (N_1005,In_844,In_2196);
nor U1006 (N_1006,In_1729,In_2316);
nand U1007 (N_1007,In_1069,In_1545);
or U1008 (N_1008,In_2398,In_1172);
nand U1009 (N_1009,In_1312,In_799);
and U1010 (N_1010,In_368,In_486);
or U1011 (N_1011,In_278,In_2479);
nor U1012 (N_1012,In_1383,In_1308);
nor U1013 (N_1013,In_1624,In_360);
and U1014 (N_1014,In_625,In_1637);
nand U1015 (N_1015,In_2311,In_1157);
or U1016 (N_1016,In_1400,In_2363);
nand U1017 (N_1017,In_2058,In_556);
or U1018 (N_1018,In_454,In_1271);
or U1019 (N_1019,In_662,In_2404);
nor U1020 (N_1020,In_1592,In_996);
or U1021 (N_1021,In_1574,In_425);
nand U1022 (N_1022,In_809,In_1828);
nor U1023 (N_1023,In_320,In_1497);
or U1024 (N_1024,In_1117,In_725);
and U1025 (N_1025,In_713,In_1149);
nand U1026 (N_1026,In_2273,In_2345);
or U1027 (N_1027,In_2436,In_1193);
nand U1028 (N_1028,In_1021,In_998);
nor U1029 (N_1029,In_1971,In_2252);
nand U1030 (N_1030,In_1527,In_169);
nand U1031 (N_1031,In_2120,In_1800);
or U1032 (N_1032,In_1480,In_1109);
nand U1033 (N_1033,In_1908,In_1433);
or U1034 (N_1034,In_963,In_861);
nand U1035 (N_1035,In_1575,In_1201);
or U1036 (N_1036,In_1356,In_1538);
nand U1037 (N_1037,In_39,In_1398);
nor U1038 (N_1038,In_444,In_1756);
or U1039 (N_1039,In_315,In_1376);
and U1040 (N_1040,In_94,In_1533);
nand U1041 (N_1041,In_260,In_2290);
nand U1042 (N_1042,In_1401,In_1784);
nor U1043 (N_1043,In_872,In_1489);
or U1044 (N_1044,In_2428,In_189);
or U1045 (N_1045,In_1697,In_2467);
nor U1046 (N_1046,In_1099,In_2267);
and U1047 (N_1047,In_419,In_162);
xor U1048 (N_1048,In_539,In_1847);
and U1049 (N_1049,In_1222,In_1385);
nand U1050 (N_1050,In_62,In_1167);
nand U1051 (N_1051,In_977,In_2082);
and U1052 (N_1052,In_2194,In_1956);
nand U1053 (N_1053,In_1409,In_15);
xor U1054 (N_1054,In_1492,In_2395);
and U1055 (N_1055,In_2088,In_2165);
and U1056 (N_1056,In_1120,In_741);
nand U1057 (N_1057,In_2387,In_1243);
xor U1058 (N_1058,In_560,In_936);
nand U1059 (N_1059,In_1421,In_2441);
and U1060 (N_1060,In_1950,In_399);
nand U1061 (N_1061,In_981,In_406);
nand U1062 (N_1062,In_1961,In_484);
nor U1063 (N_1063,In_1581,In_110);
nor U1064 (N_1064,In_271,In_180);
or U1065 (N_1065,In_704,In_2048);
nand U1066 (N_1066,In_1643,In_99);
nand U1067 (N_1067,In_754,In_2040);
or U1068 (N_1068,In_999,In_1013);
nand U1069 (N_1069,In_75,In_661);
nor U1070 (N_1070,In_1881,In_1723);
or U1071 (N_1071,In_2173,In_200);
nor U1072 (N_1072,In_1251,In_871);
nand U1073 (N_1073,In_732,In_1811);
or U1074 (N_1074,In_465,In_470);
nor U1075 (N_1075,In_507,In_759);
or U1076 (N_1076,In_1586,In_2046);
nor U1077 (N_1077,In_1454,In_1106);
nor U1078 (N_1078,In_583,In_1561);
nand U1079 (N_1079,In_1459,In_1321);
nand U1080 (N_1080,In_1223,In_1216);
and U1081 (N_1081,In_1288,In_2253);
xnor U1082 (N_1082,In_1429,In_2291);
nor U1083 (N_1083,In_2249,In_1347);
or U1084 (N_1084,In_458,In_1143);
nand U1085 (N_1085,In_2178,In_2452);
nand U1086 (N_1086,In_378,In_409);
and U1087 (N_1087,In_1278,In_1970);
nor U1088 (N_1088,In_746,In_119);
nor U1089 (N_1089,In_1822,In_1336);
xnor U1090 (N_1090,In_1160,In_1006);
and U1091 (N_1091,In_1465,In_1745);
nand U1092 (N_1092,In_1169,In_1862);
or U1093 (N_1093,In_2106,In_989);
nand U1094 (N_1094,In_420,In_78);
xor U1095 (N_1095,In_516,In_1823);
nand U1096 (N_1096,In_443,In_705);
xor U1097 (N_1097,In_331,In_263);
nand U1098 (N_1098,In_1205,In_672);
nor U1099 (N_1099,In_1177,In_752);
nor U1100 (N_1100,In_2188,In_1550);
nand U1101 (N_1101,In_2256,In_384);
and U1102 (N_1102,In_155,In_1034);
and U1103 (N_1103,In_1333,In_1605);
and U1104 (N_1104,In_312,In_974);
and U1105 (N_1105,In_942,In_2232);
xnor U1106 (N_1106,In_325,In_1142);
xor U1107 (N_1107,In_995,In_77);
and U1108 (N_1108,In_2394,In_1437);
nor U1109 (N_1109,In_1977,In_2010);
or U1110 (N_1110,In_430,In_2375);
nand U1111 (N_1111,In_666,In_1904);
nand U1112 (N_1112,In_2092,In_902);
or U1113 (N_1113,In_2059,In_1832);
or U1114 (N_1114,In_695,In_1810);
nor U1115 (N_1115,In_2337,In_535);
nand U1116 (N_1116,In_1584,In_1995);
nand U1117 (N_1117,In_652,In_1599);
nor U1118 (N_1118,In_943,In_1377);
or U1119 (N_1119,In_920,In_393);
nor U1120 (N_1120,In_1335,In_2133);
or U1121 (N_1121,In_314,In_728);
or U1122 (N_1122,In_1280,In_742);
and U1123 (N_1123,In_1573,In_1299);
nor U1124 (N_1124,In_1329,In_24);
nand U1125 (N_1125,In_1129,In_586);
and U1126 (N_1126,In_888,In_500);
or U1127 (N_1127,In_1782,In_685);
and U1128 (N_1128,In_1516,In_1630);
and U1129 (N_1129,In_665,In_707);
and U1130 (N_1130,In_940,In_328);
xor U1131 (N_1131,In_1539,In_64);
or U1132 (N_1132,In_973,In_437);
nor U1133 (N_1133,In_994,In_298);
nand U1134 (N_1134,In_363,In_2112);
or U1135 (N_1135,In_2240,In_195);
nor U1136 (N_1136,In_432,In_2393);
nor U1137 (N_1137,In_1870,In_2045);
or U1138 (N_1138,In_814,In_128);
nor U1139 (N_1139,In_599,In_93);
and U1140 (N_1140,In_1068,In_21);
and U1141 (N_1141,In_2444,In_1932);
xnor U1142 (N_1142,In_2234,In_1390);
nand U1143 (N_1143,In_1512,In_1443);
nand U1144 (N_1144,In_1953,In_2254);
nand U1145 (N_1145,In_1245,In_917);
nor U1146 (N_1146,In_1420,In_982);
and U1147 (N_1147,In_2038,In_1549);
nor U1148 (N_1148,In_609,In_32);
nor U1149 (N_1149,In_1080,In_2373);
nor U1150 (N_1150,In_1845,In_103);
and U1151 (N_1151,In_1853,In_1911);
or U1152 (N_1152,In_1236,In_1891);
nor U1153 (N_1153,In_1439,In_1865);
or U1154 (N_1154,In_414,In_242);
or U1155 (N_1155,In_1310,In_788);
nand U1156 (N_1156,In_322,In_51);
nand U1157 (N_1157,In_1095,In_694);
nor U1158 (N_1158,In_650,In_954);
nor U1159 (N_1159,In_86,In_1384);
or U1160 (N_1160,In_154,In_714);
nand U1161 (N_1161,In_109,In_1913);
xnor U1162 (N_1162,In_2451,In_2044);
and U1163 (N_1163,In_2115,In_1933);
or U1164 (N_1164,In_2175,In_2147);
nor U1165 (N_1165,In_612,In_2263);
and U1166 (N_1166,In_1132,In_807);
and U1167 (N_1167,In_307,In_629);
xnor U1168 (N_1168,In_0,In_1718);
or U1169 (N_1169,In_910,In_1928);
nor U1170 (N_1170,In_2179,In_1514);
or U1171 (N_1171,In_69,In_1835);
nand U1172 (N_1172,In_2131,In_1552);
or U1173 (N_1173,In_2225,In_2185);
nand U1174 (N_1174,In_2063,In_2012);
and U1175 (N_1175,In_735,In_514);
nand U1176 (N_1176,In_2270,In_251);
or U1177 (N_1177,In_12,In_359);
or U1178 (N_1178,In_1948,In_2243);
nand U1179 (N_1179,In_2180,In_2490);
xor U1180 (N_1180,In_1240,In_140);
nand U1181 (N_1181,In_1320,In_1187);
nor U1182 (N_1182,In_830,In_130);
or U1183 (N_1183,In_1311,In_801);
nor U1184 (N_1184,In_364,In_1247);
and U1185 (N_1185,In_617,In_2055);
or U1186 (N_1186,In_937,In_1410);
nand U1187 (N_1187,In_1793,In_76);
xor U1188 (N_1188,In_2219,In_1560);
nand U1189 (N_1189,In_519,In_1515);
or U1190 (N_1190,In_1754,In_758);
nor U1191 (N_1191,In_116,In_521);
nand U1192 (N_1192,In_1758,In_983);
nand U1193 (N_1193,In_1912,In_2413);
nand U1194 (N_1194,In_1790,In_2008);
or U1195 (N_1195,In_2159,In_587);
nand U1196 (N_1196,In_1363,In_1734);
nand U1197 (N_1197,In_478,In_389);
or U1198 (N_1198,In_1879,In_2354);
xor U1199 (N_1199,In_1070,In_1765);
nor U1200 (N_1200,In_1412,In_852);
nand U1201 (N_1201,In_400,In_1562);
and U1202 (N_1202,In_108,In_232);
nor U1203 (N_1203,In_2004,In_2079);
and U1204 (N_1204,In_1840,In_2170);
and U1205 (N_1205,In_73,In_513);
nand U1206 (N_1206,In_395,In_2193);
and U1207 (N_1207,In_1159,In_1289);
and U1208 (N_1208,In_2177,In_2233);
or U1209 (N_1209,In_1083,In_1876);
and U1210 (N_1210,In_83,In_42);
or U1211 (N_1211,In_971,In_1442);
xnor U1212 (N_1212,In_1043,In_1864);
xnor U1213 (N_1213,In_1502,In_1011);
xor U1214 (N_1214,In_2153,In_215);
and U1215 (N_1215,In_1178,In_1438);
and U1216 (N_1216,In_2260,In_2289);
nand U1217 (N_1217,In_716,In_2407);
or U1218 (N_1218,In_1855,In_2473);
nor U1219 (N_1219,In_153,In_1164);
nand U1220 (N_1220,In_1218,In_1570);
xnor U1221 (N_1221,In_55,In_1362);
nor U1222 (N_1222,In_952,In_1292);
nor U1223 (N_1223,In_439,In_303);
nand U1224 (N_1224,In_2195,In_511);
xor U1225 (N_1225,In_932,In_899);
nand U1226 (N_1226,In_885,In_356);
nor U1227 (N_1227,In_161,In_522);
xor U1228 (N_1228,In_199,In_2342);
nand U1229 (N_1229,In_1585,In_1619);
and U1230 (N_1230,In_992,In_347);
nand U1231 (N_1231,In_1286,In_1031);
and U1232 (N_1232,In_2312,In_2);
nor U1233 (N_1233,In_1824,In_1595);
or U1234 (N_1234,In_848,In_878);
nand U1235 (N_1235,In_2163,In_681);
nand U1236 (N_1236,In_1702,In_2077);
and U1237 (N_1237,In_264,In_1517);
nand U1238 (N_1238,In_683,In_2463);
and U1239 (N_1239,In_1640,In_41);
nand U1240 (N_1240,In_743,In_304);
or U1241 (N_1241,In_1633,In_1686);
or U1242 (N_1242,In_1861,In_2334);
or U1243 (N_1243,In_1180,In_1012);
nor U1244 (N_1244,In_1763,In_225);
or U1245 (N_1245,In_202,In_1107);
or U1246 (N_1246,In_2002,In_2135);
or U1247 (N_1247,In_2327,In_1930);
xor U1248 (N_1248,In_1301,In_2130);
nor U1249 (N_1249,In_1775,In_1191);
xnor U1250 (N_1250,In_135,In_1742);
and U1251 (N_1251,In_210,In_2120);
or U1252 (N_1252,In_177,In_1852);
nor U1253 (N_1253,In_550,In_2094);
and U1254 (N_1254,In_1392,In_834);
and U1255 (N_1255,In_285,In_1622);
and U1256 (N_1256,In_2241,In_1040);
nand U1257 (N_1257,In_811,In_1892);
or U1258 (N_1258,In_253,In_1356);
nor U1259 (N_1259,In_381,In_2403);
nand U1260 (N_1260,In_863,In_802);
nand U1261 (N_1261,In_2375,In_1385);
xor U1262 (N_1262,In_1367,In_497);
and U1263 (N_1263,In_766,In_1212);
xnor U1264 (N_1264,In_134,In_1487);
or U1265 (N_1265,In_2145,In_811);
nor U1266 (N_1266,In_245,In_1932);
or U1267 (N_1267,In_981,In_89);
or U1268 (N_1268,In_1655,In_2188);
xnor U1269 (N_1269,In_544,In_1079);
nor U1270 (N_1270,In_1831,In_1976);
nand U1271 (N_1271,In_148,In_439);
or U1272 (N_1272,In_121,In_1931);
nand U1273 (N_1273,In_1305,In_1306);
or U1274 (N_1274,In_699,In_1711);
nand U1275 (N_1275,In_821,In_605);
xnor U1276 (N_1276,In_2449,In_306);
and U1277 (N_1277,In_2377,In_349);
and U1278 (N_1278,In_44,In_101);
nand U1279 (N_1279,In_288,In_1322);
nor U1280 (N_1280,In_1504,In_255);
and U1281 (N_1281,In_446,In_1632);
or U1282 (N_1282,In_1864,In_201);
or U1283 (N_1283,In_1438,In_1436);
nand U1284 (N_1284,In_2174,In_1935);
nand U1285 (N_1285,In_1255,In_1488);
xor U1286 (N_1286,In_2131,In_823);
and U1287 (N_1287,In_856,In_411);
and U1288 (N_1288,In_1580,In_1088);
and U1289 (N_1289,In_2288,In_88);
and U1290 (N_1290,In_1758,In_1122);
or U1291 (N_1291,In_2474,In_680);
nand U1292 (N_1292,In_30,In_1859);
or U1293 (N_1293,In_2194,In_1714);
nand U1294 (N_1294,In_782,In_2195);
and U1295 (N_1295,In_1929,In_1871);
nand U1296 (N_1296,In_1200,In_2166);
xnor U1297 (N_1297,In_704,In_1697);
or U1298 (N_1298,In_837,In_2376);
nor U1299 (N_1299,In_712,In_765);
and U1300 (N_1300,In_176,In_1768);
nand U1301 (N_1301,In_1388,In_2139);
xnor U1302 (N_1302,In_1783,In_1791);
or U1303 (N_1303,In_814,In_1321);
xor U1304 (N_1304,In_457,In_392);
nand U1305 (N_1305,In_2034,In_200);
or U1306 (N_1306,In_2216,In_1227);
nor U1307 (N_1307,In_1980,In_100);
nor U1308 (N_1308,In_1638,In_1970);
and U1309 (N_1309,In_537,In_1698);
or U1310 (N_1310,In_1379,In_464);
nor U1311 (N_1311,In_590,In_2369);
and U1312 (N_1312,In_2336,In_1783);
nor U1313 (N_1313,In_2076,In_272);
or U1314 (N_1314,In_779,In_251);
or U1315 (N_1315,In_1029,In_1482);
nor U1316 (N_1316,In_1723,In_615);
or U1317 (N_1317,In_360,In_375);
and U1318 (N_1318,In_523,In_2409);
nor U1319 (N_1319,In_2215,In_1467);
and U1320 (N_1320,In_2165,In_576);
nor U1321 (N_1321,In_1184,In_339);
nor U1322 (N_1322,In_394,In_1416);
and U1323 (N_1323,In_1727,In_883);
xor U1324 (N_1324,In_1850,In_1576);
and U1325 (N_1325,In_442,In_1955);
and U1326 (N_1326,In_1918,In_1381);
nor U1327 (N_1327,In_270,In_973);
and U1328 (N_1328,In_541,In_1702);
xnor U1329 (N_1329,In_2032,In_711);
nor U1330 (N_1330,In_342,In_1087);
nand U1331 (N_1331,In_1288,In_1611);
nor U1332 (N_1332,In_1457,In_1540);
nor U1333 (N_1333,In_1579,In_140);
and U1334 (N_1334,In_2454,In_1559);
and U1335 (N_1335,In_1150,In_1036);
nor U1336 (N_1336,In_471,In_1351);
or U1337 (N_1337,In_2205,In_31);
nor U1338 (N_1338,In_1477,In_97);
nand U1339 (N_1339,In_1202,In_580);
xor U1340 (N_1340,In_292,In_2446);
and U1341 (N_1341,In_2077,In_723);
and U1342 (N_1342,In_1957,In_626);
nand U1343 (N_1343,In_111,In_749);
or U1344 (N_1344,In_978,In_238);
nand U1345 (N_1345,In_1473,In_2124);
or U1346 (N_1346,In_1497,In_803);
and U1347 (N_1347,In_2388,In_596);
nor U1348 (N_1348,In_1787,In_1761);
nor U1349 (N_1349,In_2202,In_2095);
or U1350 (N_1350,In_1957,In_46);
and U1351 (N_1351,In_2227,In_1624);
or U1352 (N_1352,In_447,In_1754);
nand U1353 (N_1353,In_631,In_2105);
and U1354 (N_1354,In_1002,In_2013);
and U1355 (N_1355,In_178,In_787);
nand U1356 (N_1356,In_1638,In_751);
nor U1357 (N_1357,In_141,In_612);
or U1358 (N_1358,In_998,In_1905);
nor U1359 (N_1359,In_1309,In_401);
or U1360 (N_1360,In_2416,In_743);
and U1361 (N_1361,In_2079,In_1270);
nand U1362 (N_1362,In_1853,In_433);
nor U1363 (N_1363,In_827,In_1272);
nor U1364 (N_1364,In_861,In_1416);
or U1365 (N_1365,In_1324,In_428);
nand U1366 (N_1366,In_1479,In_937);
or U1367 (N_1367,In_1079,In_521);
nand U1368 (N_1368,In_937,In_2471);
xnor U1369 (N_1369,In_1777,In_270);
or U1370 (N_1370,In_1754,In_1327);
nor U1371 (N_1371,In_2092,In_2110);
and U1372 (N_1372,In_76,In_2381);
and U1373 (N_1373,In_1891,In_2333);
nand U1374 (N_1374,In_2412,In_1591);
nand U1375 (N_1375,In_924,In_1427);
or U1376 (N_1376,In_678,In_2189);
or U1377 (N_1377,In_1089,In_1095);
nor U1378 (N_1378,In_1288,In_1232);
or U1379 (N_1379,In_1270,In_871);
or U1380 (N_1380,In_1806,In_442);
nand U1381 (N_1381,In_2060,In_796);
nand U1382 (N_1382,In_1626,In_1265);
or U1383 (N_1383,In_1211,In_1643);
or U1384 (N_1384,In_986,In_1297);
and U1385 (N_1385,In_838,In_1569);
xnor U1386 (N_1386,In_603,In_2392);
or U1387 (N_1387,In_742,In_1251);
nor U1388 (N_1388,In_312,In_1986);
or U1389 (N_1389,In_1746,In_2255);
nor U1390 (N_1390,In_1226,In_1234);
nand U1391 (N_1391,In_1044,In_46);
and U1392 (N_1392,In_192,In_2110);
or U1393 (N_1393,In_2413,In_1353);
nand U1394 (N_1394,In_1486,In_842);
xnor U1395 (N_1395,In_1799,In_122);
nor U1396 (N_1396,In_1218,In_2056);
and U1397 (N_1397,In_1988,In_863);
xnor U1398 (N_1398,In_1088,In_1040);
nand U1399 (N_1399,In_525,In_1836);
nor U1400 (N_1400,In_2294,In_979);
nand U1401 (N_1401,In_1317,In_1221);
nand U1402 (N_1402,In_1905,In_951);
and U1403 (N_1403,In_2447,In_1258);
and U1404 (N_1404,In_1678,In_1185);
nand U1405 (N_1405,In_2003,In_221);
and U1406 (N_1406,In_1254,In_57);
nand U1407 (N_1407,In_1961,In_561);
or U1408 (N_1408,In_1486,In_2098);
or U1409 (N_1409,In_1838,In_1592);
or U1410 (N_1410,In_1539,In_638);
and U1411 (N_1411,In_239,In_706);
nor U1412 (N_1412,In_1756,In_363);
or U1413 (N_1413,In_1434,In_705);
and U1414 (N_1414,In_1326,In_1118);
nand U1415 (N_1415,In_631,In_287);
and U1416 (N_1416,In_754,In_912);
nand U1417 (N_1417,In_152,In_1693);
xnor U1418 (N_1418,In_664,In_1619);
xnor U1419 (N_1419,In_2304,In_1193);
or U1420 (N_1420,In_2481,In_2031);
nand U1421 (N_1421,In_2277,In_1320);
and U1422 (N_1422,In_2469,In_1363);
nand U1423 (N_1423,In_494,In_2264);
nor U1424 (N_1424,In_477,In_478);
nor U1425 (N_1425,In_12,In_490);
xor U1426 (N_1426,In_746,In_2113);
or U1427 (N_1427,In_1434,In_1945);
nand U1428 (N_1428,In_1720,In_1492);
nor U1429 (N_1429,In_1999,In_1193);
nand U1430 (N_1430,In_1714,In_565);
or U1431 (N_1431,In_200,In_828);
xor U1432 (N_1432,In_1627,In_1112);
nor U1433 (N_1433,In_1093,In_212);
and U1434 (N_1434,In_2316,In_449);
nand U1435 (N_1435,In_1473,In_507);
nor U1436 (N_1436,In_1109,In_840);
nor U1437 (N_1437,In_1913,In_1995);
nand U1438 (N_1438,In_940,In_686);
nand U1439 (N_1439,In_926,In_2456);
nor U1440 (N_1440,In_1405,In_956);
and U1441 (N_1441,In_1590,In_1076);
xnor U1442 (N_1442,In_1585,In_2409);
or U1443 (N_1443,In_617,In_376);
nor U1444 (N_1444,In_2277,In_507);
and U1445 (N_1445,In_1989,In_106);
nand U1446 (N_1446,In_975,In_1446);
or U1447 (N_1447,In_552,In_670);
and U1448 (N_1448,In_1449,In_2316);
nand U1449 (N_1449,In_87,In_2006);
or U1450 (N_1450,In_469,In_2019);
nor U1451 (N_1451,In_1121,In_2241);
and U1452 (N_1452,In_1352,In_121);
nor U1453 (N_1453,In_1805,In_2270);
or U1454 (N_1454,In_909,In_1572);
nor U1455 (N_1455,In_1531,In_2421);
nor U1456 (N_1456,In_152,In_734);
nor U1457 (N_1457,In_809,In_430);
nor U1458 (N_1458,In_780,In_1756);
nor U1459 (N_1459,In_2186,In_227);
and U1460 (N_1460,In_1057,In_862);
or U1461 (N_1461,In_764,In_355);
nand U1462 (N_1462,In_1750,In_1380);
nand U1463 (N_1463,In_2422,In_2248);
nand U1464 (N_1464,In_665,In_1448);
or U1465 (N_1465,In_514,In_1566);
nand U1466 (N_1466,In_583,In_1004);
or U1467 (N_1467,In_1983,In_1191);
or U1468 (N_1468,In_925,In_1704);
nor U1469 (N_1469,In_222,In_1492);
or U1470 (N_1470,In_1213,In_980);
or U1471 (N_1471,In_1092,In_1798);
or U1472 (N_1472,In_576,In_1930);
and U1473 (N_1473,In_405,In_994);
nand U1474 (N_1474,In_1643,In_968);
nand U1475 (N_1475,In_1334,In_2396);
nand U1476 (N_1476,In_846,In_2075);
nor U1477 (N_1477,In_1072,In_419);
and U1478 (N_1478,In_430,In_705);
or U1479 (N_1479,In_1288,In_260);
or U1480 (N_1480,In_1700,In_1992);
or U1481 (N_1481,In_301,In_337);
and U1482 (N_1482,In_1279,In_1437);
nor U1483 (N_1483,In_873,In_1592);
or U1484 (N_1484,In_825,In_510);
or U1485 (N_1485,In_1908,In_1378);
nor U1486 (N_1486,In_2108,In_1258);
nand U1487 (N_1487,In_2142,In_1259);
and U1488 (N_1488,In_1384,In_674);
and U1489 (N_1489,In_923,In_764);
or U1490 (N_1490,In_2132,In_1351);
and U1491 (N_1491,In_1919,In_1606);
nor U1492 (N_1492,In_2027,In_1253);
and U1493 (N_1493,In_225,In_69);
and U1494 (N_1494,In_237,In_760);
nor U1495 (N_1495,In_2186,In_1865);
nand U1496 (N_1496,In_685,In_2391);
xor U1497 (N_1497,In_2420,In_1924);
and U1498 (N_1498,In_2036,In_1643);
or U1499 (N_1499,In_1291,In_221);
xnor U1500 (N_1500,In_211,In_2093);
nor U1501 (N_1501,In_1369,In_1341);
or U1502 (N_1502,In_1664,In_451);
and U1503 (N_1503,In_595,In_1346);
nand U1504 (N_1504,In_768,In_2432);
and U1505 (N_1505,In_2033,In_1174);
nor U1506 (N_1506,In_31,In_329);
or U1507 (N_1507,In_1961,In_1057);
xor U1508 (N_1508,In_352,In_920);
or U1509 (N_1509,In_1525,In_1017);
nor U1510 (N_1510,In_23,In_755);
or U1511 (N_1511,In_1994,In_1683);
nand U1512 (N_1512,In_594,In_1862);
nand U1513 (N_1513,In_506,In_1102);
and U1514 (N_1514,In_596,In_1816);
nand U1515 (N_1515,In_311,In_744);
xor U1516 (N_1516,In_369,In_420);
and U1517 (N_1517,In_2492,In_658);
nand U1518 (N_1518,In_20,In_1140);
and U1519 (N_1519,In_1265,In_1245);
or U1520 (N_1520,In_848,In_1004);
xor U1521 (N_1521,In_296,In_66);
nor U1522 (N_1522,In_592,In_412);
nand U1523 (N_1523,In_887,In_1129);
xor U1524 (N_1524,In_1380,In_1962);
and U1525 (N_1525,In_1616,In_680);
nor U1526 (N_1526,In_2258,In_2030);
nand U1527 (N_1527,In_1536,In_1200);
xor U1528 (N_1528,In_2341,In_524);
xor U1529 (N_1529,In_1208,In_1382);
and U1530 (N_1530,In_1649,In_472);
and U1531 (N_1531,In_1207,In_2045);
or U1532 (N_1532,In_1201,In_1333);
nand U1533 (N_1533,In_2315,In_1179);
and U1534 (N_1534,In_2418,In_755);
nand U1535 (N_1535,In_222,In_1524);
nor U1536 (N_1536,In_1772,In_341);
and U1537 (N_1537,In_890,In_1913);
nand U1538 (N_1538,In_1977,In_702);
nor U1539 (N_1539,In_1629,In_653);
nand U1540 (N_1540,In_358,In_2358);
xor U1541 (N_1541,In_2193,In_1325);
nand U1542 (N_1542,In_300,In_2108);
nor U1543 (N_1543,In_1689,In_1811);
xor U1544 (N_1544,In_2342,In_2422);
or U1545 (N_1545,In_1657,In_428);
nor U1546 (N_1546,In_1135,In_2075);
or U1547 (N_1547,In_567,In_1365);
and U1548 (N_1548,In_1334,In_1373);
nand U1549 (N_1549,In_616,In_2227);
or U1550 (N_1550,In_1768,In_2120);
or U1551 (N_1551,In_2182,In_1691);
nand U1552 (N_1552,In_493,In_2040);
and U1553 (N_1553,In_63,In_169);
or U1554 (N_1554,In_5,In_1971);
nor U1555 (N_1555,In_905,In_213);
nor U1556 (N_1556,In_1243,In_1525);
nand U1557 (N_1557,In_198,In_879);
nand U1558 (N_1558,In_1392,In_71);
and U1559 (N_1559,In_2146,In_1996);
and U1560 (N_1560,In_1803,In_609);
nand U1561 (N_1561,In_2151,In_397);
or U1562 (N_1562,In_657,In_2350);
or U1563 (N_1563,In_785,In_2147);
nand U1564 (N_1564,In_856,In_971);
nor U1565 (N_1565,In_526,In_751);
nand U1566 (N_1566,In_1636,In_771);
and U1567 (N_1567,In_1067,In_591);
nand U1568 (N_1568,In_1736,In_1160);
nand U1569 (N_1569,In_1949,In_1994);
nand U1570 (N_1570,In_647,In_1965);
nand U1571 (N_1571,In_977,In_241);
nand U1572 (N_1572,In_712,In_503);
and U1573 (N_1573,In_1039,In_2417);
and U1574 (N_1574,In_1983,In_2403);
nand U1575 (N_1575,In_1770,In_1742);
nor U1576 (N_1576,In_918,In_688);
xor U1577 (N_1577,In_868,In_762);
and U1578 (N_1578,In_1233,In_1069);
and U1579 (N_1579,In_2096,In_580);
nor U1580 (N_1580,In_878,In_1133);
nor U1581 (N_1581,In_1623,In_1443);
nand U1582 (N_1582,In_107,In_115);
nand U1583 (N_1583,In_204,In_993);
nor U1584 (N_1584,In_2072,In_111);
nor U1585 (N_1585,In_472,In_2040);
or U1586 (N_1586,In_2449,In_1417);
nand U1587 (N_1587,In_1624,In_309);
or U1588 (N_1588,In_151,In_2413);
xor U1589 (N_1589,In_1727,In_1075);
nor U1590 (N_1590,In_1891,In_792);
and U1591 (N_1591,In_1423,In_1569);
or U1592 (N_1592,In_2368,In_109);
nor U1593 (N_1593,In_1406,In_1828);
nor U1594 (N_1594,In_1012,In_915);
nand U1595 (N_1595,In_2014,In_1126);
and U1596 (N_1596,In_1682,In_1908);
nor U1597 (N_1597,In_1379,In_837);
and U1598 (N_1598,In_1154,In_1734);
nand U1599 (N_1599,In_2314,In_2366);
and U1600 (N_1600,In_1734,In_2230);
or U1601 (N_1601,In_159,In_1443);
nand U1602 (N_1602,In_1157,In_844);
nand U1603 (N_1603,In_977,In_2483);
or U1604 (N_1604,In_667,In_1084);
nor U1605 (N_1605,In_2319,In_1703);
or U1606 (N_1606,In_1438,In_2036);
and U1607 (N_1607,In_1921,In_1338);
nor U1608 (N_1608,In_1107,In_1980);
nand U1609 (N_1609,In_1284,In_404);
nor U1610 (N_1610,In_1790,In_2322);
or U1611 (N_1611,In_13,In_1113);
and U1612 (N_1612,In_805,In_486);
xnor U1613 (N_1613,In_1186,In_2115);
or U1614 (N_1614,In_762,In_389);
nand U1615 (N_1615,In_2340,In_2144);
and U1616 (N_1616,In_64,In_2129);
nand U1617 (N_1617,In_1295,In_2241);
and U1618 (N_1618,In_1765,In_1888);
nand U1619 (N_1619,In_527,In_1584);
and U1620 (N_1620,In_859,In_584);
and U1621 (N_1621,In_630,In_75);
or U1622 (N_1622,In_1748,In_2005);
and U1623 (N_1623,In_1496,In_1884);
nor U1624 (N_1624,In_2404,In_192);
xor U1625 (N_1625,In_2026,In_580);
and U1626 (N_1626,In_1486,In_992);
and U1627 (N_1627,In_2342,In_1598);
or U1628 (N_1628,In_1629,In_2450);
nand U1629 (N_1629,In_949,In_604);
or U1630 (N_1630,In_2278,In_1342);
and U1631 (N_1631,In_1525,In_2422);
or U1632 (N_1632,In_7,In_1105);
nand U1633 (N_1633,In_731,In_1536);
nor U1634 (N_1634,In_1335,In_660);
or U1635 (N_1635,In_1298,In_1722);
nand U1636 (N_1636,In_161,In_240);
nor U1637 (N_1637,In_1259,In_383);
or U1638 (N_1638,In_172,In_2289);
or U1639 (N_1639,In_1789,In_428);
nor U1640 (N_1640,In_2381,In_692);
nor U1641 (N_1641,In_1920,In_1725);
and U1642 (N_1642,In_523,In_2020);
and U1643 (N_1643,In_2386,In_1538);
nor U1644 (N_1644,In_2008,In_104);
and U1645 (N_1645,In_2468,In_754);
nor U1646 (N_1646,In_1432,In_2473);
xor U1647 (N_1647,In_1860,In_421);
nand U1648 (N_1648,In_169,In_1580);
nand U1649 (N_1649,In_897,In_2290);
and U1650 (N_1650,In_1956,In_464);
nand U1651 (N_1651,In_341,In_1097);
nor U1652 (N_1652,In_353,In_1708);
nor U1653 (N_1653,In_726,In_1989);
nor U1654 (N_1654,In_2098,In_1683);
nor U1655 (N_1655,In_2267,In_908);
nand U1656 (N_1656,In_160,In_1935);
xor U1657 (N_1657,In_1430,In_1079);
nor U1658 (N_1658,In_2434,In_357);
xor U1659 (N_1659,In_98,In_529);
nand U1660 (N_1660,In_425,In_899);
nor U1661 (N_1661,In_1670,In_1867);
nand U1662 (N_1662,In_1662,In_984);
and U1663 (N_1663,In_1125,In_892);
nor U1664 (N_1664,In_114,In_933);
or U1665 (N_1665,In_475,In_61);
nor U1666 (N_1666,In_2393,In_2056);
nand U1667 (N_1667,In_2259,In_612);
and U1668 (N_1668,In_1956,In_1194);
nor U1669 (N_1669,In_2297,In_654);
nand U1670 (N_1670,In_829,In_1981);
xnor U1671 (N_1671,In_877,In_135);
and U1672 (N_1672,In_1553,In_939);
or U1673 (N_1673,In_2266,In_2288);
nand U1674 (N_1674,In_301,In_1037);
nor U1675 (N_1675,In_1160,In_2018);
nor U1676 (N_1676,In_1269,In_668);
nand U1677 (N_1677,In_2247,In_1402);
and U1678 (N_1678,In_373,In_1046);
or U1679 (N_1679,In_1312,In_1968);
or U1680 (N_1680,In_1448,In_1111);
xnor U1681 (N_1681,In_807,In_2055);
nor U1682 (N_1682,In_1777,In_935);
or U1683 (N_1683,In_90,In_2315);
nor U1684 (N_1684,In_1141,In_448);
nand U1685 (N_1685,In_2016,In_732);
xnor U1686 (N_1686,In_1779,In_1676);
and U1687 (N_1687,In_2356,In_800);
and U1688 (N_1688,In_1819,In_376);
xor U1689 (N_1689,In_1496,In_1162);
nor U1690 (N_1690,In_1545,In_264);
or U1691 (N_1691,In_207,In_1675);
or U1692 (N_1692,In_1174,In_77);
nand U1693 (N_1693,In_1413,In_1015);
or U1694 (N_1694,In_542,In_1109);
nand U1695 (N_1695,In_406,In_924);
or U1696 (N_1696,In_235,In_63);
and U1697 (N_1697,In_899,In_1928);
and U1698 (N_1698,In_2258,In_1517);
and U1699 (N_1699,In_231,In_947);
or U1700 (N_1700,In_1865,In_1966);
nor U1701 (N_1701,In_2179,In_1161);
nor U1702 (N_1702,In_1097,In_1716);
and U1703 (N_1703,In_917,In_1373);
nand U1704 (N_1704,In_1328,In_9);
or U1705 (N_1705,In_716,In_216);
xnor U1706 (N_1706,In_1653,In_1660);
and U1707 (N_1707,In_1203,In_2484);
or U1708 (N_1708,In_1869,In_2426);
nor U1709 (N_1709,In_861,In_1053);
or U1710 (N_1710,In_2135,In_906);
or U1711 (N_1711,In_1825,In_1411);
xor U1712 (N_1712,In_107,In_1026);
xnor U1713 (N_1713,In_2221,In_811);
nand U1714 (N_1714,In_415,In_2043);
or U1715 (N_1715,In_1734,In_1959);
nand U1716 (N_1716,In_147,In_281);
or U1717 (N_1717,In_976,In_2102);
nor U1718 (N_1718,In_5,In_66);
nor U1719 (N_1719,In_775,In_1886);
nor U1720 (N_1720,In_1034,In_26);
nor U1721 (N_1721,In_507,In_1243);
nor U1722 (N_1722,In_1239,In_612);
or U1723 (N_1723,In_13,In_529);
nor U1724 (N_1724,In_1782,In_335);
nor U1725 (N_1725,In_1202,In_257);
and U1726 (N_1726,In_1648,In_208);
nor U1727 (N_1727,In_940,In_1267);
and U1728 (N_1728,In_320,In_37);
or U1729 (N_1729,In_1481,In_1599);
or U1730 (N_1730,In_752,In_1548);
nand U1731 (N_1731,In_791,In_1931);
nor U1732 (N_1732,In_789,In_2316);
and U1733 (N_1733,In_1122,In_333);
and U1734 (N_1734,In_1265,In_1478);
and U1735 (N_1735,In_1309,In_848);
and U1736 (N_1736,In_1232,In_821);
xnor U1737 (N_1737,In_1846,In_55);
or U1738 (N_1738,In_2278,In_679);
nor U1739 (N_1739,In_864,In_2055);
or U1740 (N_1740,In_284,In_184);
or U1741 (N_1741,In_652,In_87);
xnor U1742 (N_1742,In_249,In_1343);
or U1743 (N_1743,In_570,In_1767);
nor U1744 (N_1744,In_451,In_983);
nand U1745 (N_1745,In_934,In_1596);
nand U1746 (N_1746,In_1441,In_697);
xor U1747 (N_1747,In_64,In_1887);
and U1748 (N_1748,In_1108,In_357);
or U1749 (N_1749,In_2294,In_250);
nand U1750 (N_1750,In_1700,In_2234);
nor U1751 (N_1751,In_2010,In_1473);
or U1752 (N_1752,In_602,In_1810);
and U1753 (N_1753,In_233,In_1070);
or U1754 (N_1754,In_1320,In_2184);
nand U1755 (N_1755,In_2406,In_2018);
and U1756 (N_1756,In_1057,In_1911);
and U1757 (N_1757,In_2289,In_880);
nor U1758 (N_1758,In_759,In_38);
and U1759 (N_1759,In_31,In_493);
nor U1760 (N_1760,In_1102,In_1237);
nand U1761 (N_1761,In_1716,In_2014);
xor U1762 (N_1762,In_285,In_2153);
or U1763 (N_1763,In_2498,In_2129);
or U1764 (N_1764,In_2114,In_1073);
xor U1765 (N_1765,In_1898,In_1165);
and U1766 (N_1766,In_2078,In_1486);
nand U1767 (N_1767,In_1817,In_2306);
nand U1768 (N_1768,In_985,In_417);
nor U1769 (N_1769,In_1378,In_997);
and U1770 (N_1770,In_360,In_270);
and U1771 (N_1771,In_2385,In_2407);
and U1772 (N_1772,In_2305,In_871);
and U1773 (N_1773,In_2358,In_1663);
or U1774 (N_1774,In_2243,In_4);
nor U1775 (N_1775,In_1286,In_886);
and U1776 (N_1776,In_455,In_899);
nand U1777 (N_1777,In_1835,In_1883);
nand U1778 (N_1778,In_1570,In_762);
nor U1779 (N_1779,In_1662,In_1813);
and U1780 (N_1780,In_2303,In_331);
or U1781 (N_1781,In_641,In_2140);
or U1782 (N_1782,In_1142,In_1278);
nor U1783 (N_1783,In_249,In_95);
or U1784 (N_1784,In_1072,In_107);
or U1785 (N_1785,In_2479,In_40);
or U1786 (N_1786,In_2253,In_2079);
nor U1787 (N_1787,In_1783,In_2042);
or U1788 (N_1788,In_879,In_211);
nand U1789 (N_1789,In_496,In_715);
and U1790 (N_1790,In_90,In_105);
xor U1791 (N_1791,In_2499,In_1376);
nand U1792 (N_1792,In_1955,In_1605);
nor U1793 (N_1793,In_335,In_1777);
xnor U1794 (N_1794,In_1524,In_2488);
nor U1795 (N_1795,In_2461,In_2445);
or U1796 (N_1796,In_345,In_370);
nand U1797 (N_1797,In_2363,In_1906);
nand U1798 (N_1798,In_1563,In_124);
nor U1799 (N_1799,In_2296,In_905);
and U1800 (N_1800,In_2456,In_642);
xor U1801 (N_1801,In_2051,In_1650);
nor U1802 (N_1802,In_1716,In_2072);
nor U1803 (N_1803,In_854,In_1163);
nand U1804 (N_1804,In_716,In_79);
and U1805 (N_1805,In_199,In_1016);
and U1806 (N_1806,In_2278,In_804);
nand U1807 (N_1807,In_770,In_684);
nor U1808 (N_1808,In_1208,In_579);
nand U1809 (N_1809,In_310,In_1379);
and U1810 (N_1810,In_1140,In_177);
nand U1811 (N_1811,In_1526,In_1538);
or U1812 (N_1812,In_2456,In_1506);
and U1813 (N_1813,In_297,In_526);
nand U1814 (N_1814,In_1433,In_521);
nand U1815 (N_1815,In_32,In_697);
or U1816 (N_1816,In_1256,In_830);
or U1817 (N_1817,In_552,In_1279);
xnor U1818 (N_1818,In_433,In_834);
and U1819 (N_1819,In_523,In_2295);
nand U1820 (N_1820,In_1567,In_412);
nor U1821 (N_1821,In_1739,In_1619);
nor U1822 (N_1822,In_1161,In_199);
nor U1823 (N_1823,In_1414,In_1334);
nand U1824 (N_1824,In_1488,In_2025);
or U1825 (N_1825,In_1608,In_1216);
xnor U1826 (N_1826,In_2214,In_1581);
nand U1827 (N_1827,In_1590,In_2390);
nor U1828 (N_1828,In_1535,In_1725);
or U1829 (N_1829,In_2243,In_1712);
and U1830 (N_1830,In_1131,In_639);
or U1831 (N_1831,In_881,In_583);
and U1832 (N_1832,In_2281,In_1425);
nand U1833 (N_1833,In_2495,In_2030);
and U1834 (N_1834,In_811,In_21);
nor U1835 (N_1835,In_1456,In_612);
nand U1836 (N_1836,In_573,In_1421);
or U1837 (N_1837,In_1973,In_1583);
nand U1838 (N_1838,In_2047,In_1887);
or U1839 (N_1839,In_1499,In_870);
nor U1840 (N_1840,In_1145,In_66);
and U1841 (N_1841,In_237,In_1332);
nor U1842 (N_1842,In_1943,In_1436);
nand U1843 (N_1843,In_1994,In_1858);
and U1844 (N_1844,In_2253,In_2303);
nand U1845 (N_1845,In_760,In_1427);
and U1846 (N_1846,In_505,In_1888);
nor U1847 (N_1847,In_452,In_107);
xnor U1848 (N_1848,In_1342,In_936);
nand U1849 (N_1849,In_711,In_1941);
and U1850 (N_1850,In_2048,In_922);
nor U1851 (N_1851,In_687,In_961);
nand U1852 (N_1852,In_172,In_145);
nand U1853 (N_1853,In_2296,In_1474);
nand U1854 (N_1854,In_822,In_2441);
or U1855 (N_1855,In_857,In_1847);
xnor U1856 (N_1856,In_942,In_463);
xor U1857 (N_1857,In_1012,In_1445);
and U1858 (N_1858,In_1063,In_1848);
or U1859 (N_1859,In_1096,In_2490);
nand U1860 (N_1860,In_1085,In_201);
nand U1861 (N_1861,In_1936,In_1719);
nand U1862 (N_1862,In_1184,In_970);
nand U1863 (N_1863,In_1663,In_1015);
or U1864 (N_1864,In_2213,In_688);
nand U1865 (N_1865,In_698,In_2098);
nor U1866 (N_1866,In_1791,In_704);
and U1867 (N_1867,In_29,In_785);
or U1868 (N_1868,In_1284,In_2140);
nand U1869 (N_1869,In_1873,In_1002);
nand U1870 (N_1870,In_1015,In_1782);
nor U1871 (N_1871,In_2360,In_667);
and U1872 (N_1872,In_2472,In_413);
nand U1873 (N_1873,In_1149,In_2050);
nand U1874 (N_1874,In_1111,In_183);
or U1875 (N_1875,In_894,In_154);
and U1876 (N_1876,In_2353,In_2208);
xor U1877 (N_1877,In_243,In_791);
nor U1878 (N_1878,In_287,In_827);
nand U1879 (N_1879,In_2155,In_2143);
or U1880 (N_1880,In_1754,In_1766);
nor U1881 (N_1881,In_2289,In_496);
nand U1882 (N_1882,In_2246,In_370);
or U1883 (N_1883,In_993,In_2083);
and U1884 (N_1884,In_298,In_1260);
xnor U1885 (N_1885,In_1494,In_1137);
and U1886 (N_1886,In_1218,In_1248);
nand U1887 (N_1887,In_323,In_2086);
nor U1888 (N_1888,In_1571,In_1058);
or U1889 (N_1889,In_603,In_2391);
and U1890 (N_1890,In_167,In_2027);
nor U1891 (N_1891,In_426,In_28);
nor U1892 (N_1892,In_902,In_814);
and U1893 (N_1893,In_1782,In_59);
and U1894 (N_1894,In_1009,In_461);
nor U1895 (N_1895,In_1511,In_2172);
or U1896 (N_1896,In_2343,In_1199);
and U1897 (N_1897,In_295,In_1763);
or U1898 (N_1898,In_2195,In_6);
and U1899 (N_1899,In_209,In_778);
and U1900 (N_1900,In_531,In_738);
nor U1901 (N_1901,In_1072,In_39);
nor U1902 (N_1902,In_2143,In_1719);
or U1903 (N_1903,In_1303,In_297);
and U1904 (N_1904,In_2155,In_1054);
or U1905 (N_1905,In_1576,In_1237);
and U1906 (N_1906,In_1720,In_252);
or U1907 (N_1907,In_932,In_1387);
nor U1908 (N_1908,In_1862,In_919);
nor U1909 (N_1909,In_374,In_2104);
or U1910 (N_1910,In_2385,In_1076);
and U1911 (N_1911,In_291,In_2312);
nand U1912 (N_1912,In_634,In_417);
nand U1913 (N_1913,In_551,In_1234);
nand U1914 (N_1914,In_2396,In_1687);
nand U1915 (N_1915,In_167,In_2382);
nand U1916 (N_1916,In_1482,In_1383);
and U1917 (N_1917,In_141,In_1787);
or U1918 (N_1918,In_2494,In_100);
and U1919 (N_1919,In_1421,In_637);
and U1920 (N_1920,In_787,In_680);
nand U1921 (N_1921,In_1592,In_2321);
nand U1922 (N_1922,In_2046,In_653);
nand U1923 (N_1923,In_395,In_1780);
and U1924 (N_1924,In_2166,In_701);
or U1925 (N_1925,In_1371,In_2055);
xnor U1926 (N_1926,In_1259,In_268);
nor U1927 (N_1927,In_1843,In_448);
nand U1928 (N_1928,In_2360,In_1129);
and U1929 (N_1929,In_1884,In_1293);
nor U1930 (N_1930,In_886,In_285);
or U1931 (N_1931,In_935,In_2086);
nor U1932 (N_1932,In_938,In_1713);
nor U1933 (N_1933,In_1775,In_1270);
nor U1934 (N_1934,In_639,In_283);
nand U1935 (N_1935,In_217,In_1760);
or U1936 (N_1936,In_334,In_2157);
nand U1937 (N_1937,In_2061,In_637);
nor U1938 (N_1938,In_2110,In_1103);
and U1939 (N_1939,In_1178,In_1709);
or U1940 (N_1940,In_990,In_833);
xnor U1941 (N_1941,In_1680,In_793);
nand U1942 (N_1942,In_2463,In_2088);
or U1943 (N_1943,In_2134,In_1926);
and U1944 (N_1944,In_1360,In_1143);
and U1945 (N_1945,In_346,In_90);
nor U1946 (N_1946,In_32,In_867);
and U1947 (N_1947,In_242,In_1733);
and U1948 (N_1948,In_1980,In_971);
and U1949 (N_1949,In_372,In_2368);
or U1950 (N_1950,In_2272,In_1111);
or U1951 (N_1951,In_2400,In_569);
and U1952 (N_1952,In_257,In_509);
or U1953 (N_1953,In_2090,In_389);
or U1954 (N_1954,In_1497,In_182);
nor U1955 (N_1955,In_148,In_1385);
or U1956 (N_1956,In_628,In_358);
nor U1957 (N_1957,In_1514,In_218);
nand U1958 (N_1958,In_1840,In_841);
and U1959 (N_1959,In_2105,In_664);
nand U1960 (N_1960,In_1896,In_739);
nand U1961 (N_1961,In_1228,In_1614);
and U1962 (N_1962,In_184,In_838);
or U1963 (N_1963,In_276,In_876);
nor U1964 (N_1964,In_1000,In_2300);
or U1965 (N_1965,In_765,In_456);
nand U1966 (N_1966,In_620,In_647);
or U1967 (N_1967,In_1131,In_2169);
nand U1968 (N_1968,In_423,In_2237);
nand U1969 (N_1969,In_829,In_845);
and U1970 (N_1970,In_560,In_2174);
nand U1971 (N_1971,In_1798,In_1689);
nor U1972 (N_1972,In_974,In_491);
nand U1973 (N_1973,In_635,In_1855);
nand U1974 (N_1974,In_854,In_307);
nor U1975 (N_1975,In_729,In_747);
nor U1976 (N_1976,In_1060,In_947);
nor U1977 (N_1977,In_838,In_1801);
nand U1978 (N_1978,In_560,In_1945);
nor U1979 (N_1979,In_341,In_2403);
and U1980 (N_1980,In_1280,In_1068);
and U1981 (N_1981,In_100,In_2385);
and U1982 (N_1982,In_933,In_874);
nor U1983 (N_1983,In_171,In_1652);
and U1984 (N_1984,In_1273,In_170);
nand U1985 (N_1985,In_2048,In_1593);
nor U1986 (N_1986,In_2041,In_2243);
or U1987 (N_1987,In_307,In_2209);
nor U1988 (N_1988,In_1841,In_1460);
nand U1989 (N_1989,In_1783,In_608);
nand U1990 (N_1990,In_1738,In_686);
or U1991 (N_1991,In_587,In_117);
nand U1992 (N_1992,In_195,In_1360);
and U1993 (N_1993,In_1230,In_2428);
or U1994 (N_1994,In_2305,In_2060);
nand U1995 (N_1995,In_823,In_1286);
nand U1996 (N_1996,In_711,In_2353);
nand U1997 (N_1997,In_440,In_416);
or U1998 (N_1998,In_1452,In_482);
nor U1999 (N_1999,In_39,In_2110);
and U2000 (N_2000,In_1224,In_2356);
and U2001 (N_2001,In_1702,In_1133);
or U2002 (N_2002,In_1661,In_1485);
xnor U2003 (N_2003,In_1146,In_2061);
nand U2004 (N_2004,In_2142,In_2294);
nand U2005 (N_2005,In_1940,In_1521);
or U2006 (N_2006,In_1862,In_540);
or U2007 (N_2007,In_1288,In_583);
and U2008 (N_2008,In_310,In_2254);
nand U2009 (N_2009,In_284,In_1058);
nand U2010 (N_2010,In_1252,In_1921);
and U2011 (N_2011,In_2399,In_2032);
nor U2012 (N_2012,In_541,In_2179);
and U2013 (N_2013,In_2404,In_882);
nor U2014 (N_2014,In_963,In_1379);
and U2015 (N_2015,In_2098,In_228);
and U2016 (N_2016,In_565,In_2491);
and U2017 (N_2017,In_1339,In_1788);
nor U2018 (N_2018,In_590,In_2126);
nand U2019 (N_2019,In_1784,In_1177);
nand U2020 (N_2020,In_2107,In_2000);
nand U2021 (N_2021,In_1112,In_1870);
nand U2022 (N_2022,In_1422,In_1425);
nand U2023 (N_2023,In_249,In_1380);
nand U2024 (N_2024,In_16,In_77);
nand U2025 (N_2025,In_1364,In_2498);
nand U2026 (N_2026,In_1671,In_589);
nor U2027 (N_2027,In_1354,In_266);
nand U2028 (N_2028,In_319,In_2172);
and U2029 (N_2029,In_1117,In_1915);
or U2030 (N_2030,In_615,In_15);
and U2031 (N_2031,In_2269,In_1169);
or U2032 (N_2032,In_2386,In_704);
nand U2033 (N_2033,In_1396,In_1137);
nor U2034 (N_2034,In_374,In_133);
or U2035 (N_2035,In_680,In_850);
and U2036 (N_2036,In_805,In_1444);
and U2037 (N_2037,In_1620,In_1666);
nand U2038 (N_2038,In_1415,In_1775);
nor U2039 (N_2039,In_919,In_2291);
or U2040 (N_2040,In_1296,In_2264);
nor U2041 (N_2041,In_1177,In_974);
nor U2042 (N_2042,In_1655,In_168);
or U2043 (N_2043,In_472,In_445);
nand U2044 (N_2044,In_2324,In_1934);
nand U2045 (N_2045,In_129,In_576);
nor U2046 (N_2046,In_1265,In_1818);
nor U2047 (N_2047,In_2417,In_804);
and U2048 (N_2048,In_95,In_2126);
and U2049 (N_2049,In_522,In_1801);
nor U2050 (N_2050,In_2201,In_46);
and U2051 (N_2051,In_1118,In_1382);
nor U2052 (N_2052,In_1901,In_1373);
nand U2053 (N_2053,In_867,In_937);
nor U2054 (N_2054,In_698,In_753);
nor U2055 (N_2055,In_1467,In_802);
nand U2056 (N_2056,In_1432,In_1128);
nand U2057 (N_2057,In_2063,In_98);
or U2058 (N_2058,In_1553,In_1295);
xor U2059 (N_2059,In_1158,In_943);
nor U2060 (N_2060,In_626,In_79);
nor U2061 (N_2061,In_1624,In_1679);
and U2062 (N_2062,In_1913,In_930);
and U2063 (N_2063,In_1688,In_937);
or U2064 (N_2064,In_1801,In_842);
and U2065 (N_2065,In_1968,In_335);
and U2066 (N_2066,In_379,In_2179);
and U2067 (N_2067,In_204,In_954);
nor U2068 (N_2068,In_2009,In_1253);
xnor U2069 (N_2069,In_644,In_1372);
nor U2070 (N_2070,In_2322,In_954);
nor U2071 (N_2071,In_1734,In_2048);
nor U2072 (N_2072,In_2295,In_2270);
nor U2073 (N_2073,In_406,In_1860);
and U2074 (N_2074,In_1840,In_923);
nand U2075 (N_2075,In_789,In_2492);
nand U2076 (N_2076,In_1860,In_1506);
nand U2077 (N_2077,In_1291,In_2133);
or U2078 (N_2078,In_446,In_894);
or U2079 (N_2079,In_2008,In_1272);
nor U2080 (N_2080,In_614,In_1916);
or U2081 (N_2081,In_1437,In_1547);
xor U2082 (N_2082,In_2220,In_535);
nand U2083 (N_2083,In_1239,In_378);
or U2084 (N_2084,In_1386,In_1637);
and U2085 (N_2085,In_403,In_1943);
nand U2086 (N_2086,In_1044,In_1024);
or U2087 (N_2087,In_735,In_864);
or U2088 (N_2088,In_1237,In_2319);
nor U2089 (N_2089,In_1444,In_944);
and U2090 (N_2090,In_80,In_458);
and U2091 (N_2091,In_729,In_860);
nor U2092 (N_2092,In_2294,In_2082);
nand U2093 (N_2093,In_1859,In_2063);
nand U2094 (N_2094,In_422,In_2246);
nor U2095 (N_2095,In_1353,In_2139);
nor U2096 (N_2096,In_2008,In_95);
and U2097 (N_2097,In_2120,In_2381);
and U2098 (N_2098,In_1544,In_753);
nor U2099 (N_2099,In_899,In_97);
or U2100 (N_2100,In_1603,In_1071);
nand U2101 (N_2101,In_686,In_1387);
nand U2102 (N_2102,In_761,In_126);
nand U2103 (N_2103,In_2418,In_1575);
nand U2104 (N_2104,In_752,In_1647);
or U2105 (N_2105,In_1395,In_570);
nor U2106 (N_2106,In_791,In_379);
or U2107 (N_2107,In_2066,In_1294);
and U2108 (N_2108,In_723,In_1404);
nand U2109 (N_2109,In_1231,In_1413);
nor U2110 (N_2110,In_517,In_360);
or U2111 (N_2111,In_575,In_2015);
nor U2112 (N_2112,In_141,In_1408);
and U2113 (N_2113,In_1243,In_870);
and U2114 (N_2114,In_709,In_1893);
or U2115 (N_2115,In_1461,In_68);
nor U2116 (N_2116,In_77,In_1007);
nand U2117 (N_2117,In_25,In_948);
nor U2118 (N_2118,In_2285,In_910);
or U2119 (N_2119,In_1759,In_488);
nor U2120 (N_2120,In_634,In_126);
nand U2121 (N_2121,In_2440,In_263);
or U2122 (N_2122,In_181,In_1466);
nor U2123 (N_2123,In_574,In_240);
nand U2124 (N_2124,In_417,In_2294);
xnor U2125 (N_2125,In_294,In_1732);
xor U2126 (N_2126,In_124,In_532);
nand U2127 (N_2127,In_2424,In_1954);
or U2128 (N_2128,In_773,In_1705);
nand U2129 (N_2129,In_674,In_1977);
nor U2130 (N_2130,In_2228,In_1093);
or U2131 (N_2131,In_1656,In_2473);
or U2132 (N_2132,In_1224,In_596);
nor U2133 (N_2133,In_1868,In_1651);
and U2134 (N_2134,In_2181,In_1654);
or U2135 (N_2135,In_905,In_1684);
or U2136 (N_2136,In_1963,In_2153);
and U2137 (N_2137,In_1299,In_1307);
xor U2138 (N_2138,In_2043,In_172);
and U2139 (N_2139,In_1412,In_613);
or U2140 (N_2140,In_179,In_1854);
nand U2141 (N_2141,In_636,In_1827);
or U2142 (N_2142,In_1428,In_2499);
and U2143 (N_2143,In_2289,In_1899);
or U2144 (N_2144,In_532,In_2158);
or U2145 (N_2145,In_667,In_1869);
or U2146 (N_2146,In_407,In_1266);
nor U2147 (N_2147,In_495,In_968);
or U2148 (N_2148,In_625,In_608);
nand U2149 (N_2149,In_1248,In_410);
or U2150 (N_2150,In_2342,In_98);
and U2151 (N_2151,In_1721,In_174);
nor U2152 (N_2152,In_700,In_240);
nor U2153 (N_2153,In_1700,In_560);
nand U2154 (N_2154,In_332,In_2367);
and U2155 (N_2155,In_1393,In_1977);
nand U2156 (N_2156,In_1075,In_1215);
nor U2157 (N_2157,In_1141,In_2358);
nor U2158 (N_2158,In_2025,In_2410);
nor U2159 (N_2159,In_2219,In_2063);
and U2160 (N_2160,In_2263,In_1103);
or U2161 (N_2161,In_291,In_370);
nor U2162 (N_2162,In_1839,In_56);
and U2163 (N_2163,In_1442,In_960);
nor U2164 (N_2164,In_2051,In_189);
or U2165 (N_2165,In_1664,In_395);
xor U2166 (N_2166,In_2124,In_101);
nand U2167 (N_2167,In_469,In_1788);
nor U2168 (N_2168,In_588,In_1865);
nor U2169 (N_2169,In_1775,In_949);
nor U2170 (N_2170,In_744,In_1455);
and U2171 (N_2171,In_1149,In_237);
or U2172 (N_2172,In_1795,In_1768);
nand U2173 (N_2173,In_1257,In_685);
or U2174 (N_2174,In_420,In_2269);
or U2175 (N_2175,In_259,In_131);
nand U2176 (N_2176,In_1492,In_244);
and U2177 (N_2177,In_2448,In_810);
nand U2178 (N_2178,In_548,In_560);
nand U2179 (N_2179,In_218,In_1968);
nand U2180 (N_2180,In_935,In_548);
xor U2181 (N_2181,In_2254,In_1686);
and U2182 (N_2182,In_2399,In_747);
or U2183 (N_2183,In_205,In_1401);
nor U2184 (N_2184,In_104,In_913);
and U2185 (N_2185,In_1713,In_1693);
or U2186 (N_2186,In_2151,In_1510);
and U2187 (N_2187,In_881,In_1045);
nand U2188 (N_2188,In_707,In_1912);
xor U2189 (N_2189,In_912,In_1260);
nand U2190 (N_2190,In_677,In_1818);
nor U2191 (N_2191,In_1428,In_1849);
nand U2192 (N_2192,In_1786,In_970);
and U2193 (N_2193,In_272,In_1613);
xnor U2194 (N_2194,In_1156,In_207);
nor U2195 (N_2195,In_2381,In_2146);
and U2196 (N_2196,In_813,In_1921);
and U2197 (N_2197,In_2233,In_855);
nand U2198 (N_2198,In_951,In_1414);
or U2199 (N_2199,In_419,In_216);
and U2200 (N_2200,In_249,In_1431);
and U2201 (N_2201,In_1140,In_1710);
and U2202 (N_2202,In_1762,In_1101);
nor U2203 (N_2203,In_888,In_1188);
nor U2204 (N_2204,In_1787,In_2217);
nor U2205 (N_2205,In_682,In_631);
xnor U2206 (N_2206,In_1975,In_1976);
or U2207 (N_2207,In_806,In_1144);
nor U2208 (N_2208,In_51,In_1376);
nand U2209 (N_2209,In_1698,In_2209);
or U2210 (N_2210,In_2455,In_272);
or U2211 (N_2211,In_1201,In_1488);
and U2212 (N_2212,In_127,In_195);
nand U2213 (N_2213,In_1028,In_259);
nor U2214 (N_2214,In_808,In_226);
and U2215 (N_2215,In_2137,In_360);
or U2216 (N_2216,In_2375,In_445);
and U2217 (N_2217,In_680,In_2045);
nand U2218 (N_2218,In_1438,In_990);
xnor U2219 (N_2219,In_1864,In_2150);
or U2220 (N_2220,In_485,In_1264);
or U2221 (N_2221,In_1084,In_441);
and U2222 (N_2222,In_1837,In_932);
nor U2223 (N_2223,In_2256,In_1193);
and U2224 (N_2224,In_6,In_1949);
nor U2225 (N_2225,In_726,In_2217);
and U2226 (N_2226,In_1772,In_1199);
nor U2227 (N_2227,In_1223,In_1556);
nor U2228 (N_2228,In_2394,In_1285);
nor U2229 (N_2229,In_1243,In_1301);
nand U2230 (N_2230,In_1915,In_1868);
xnor U2231 (N_2231,In_808,In_1054);
or U2232 (N_2232,In_357,In_644);
nor U2233 (N_2233,In_2339,In_674);
and U2234 (N_2234,In_50,In_1389);
nor U2235 (N_2235,In_60,In_2173);
nand U2236 (N_2236,In_1408,In_2173);
and U2237 (N_2237,In_1050,In_184);
or U2238 (N_2238,In_1177,In_1508);
xor U2239 (N_2239,In_1869,In_391);
nor U2240 (N_2240,In_378,In_2212);
or U2241 (N_2241,In_986,In_2104);
nor U2242 (N_2242,In_606,In_715);
and U2243 (N_2243,In_1134,In_1847);
or U2244 (N_2244,In_1236,In_526);
and U2245 (N_2245,In_388,In_1670);
nand U2246 (N_2246,In_775,In_1228);
xor U2247 (N_2247,In_1415,In_1690);
and U2248 (N_2248,In_1128,In_1495);
nor U2249 (N_2249,In_2164,In_2125);
or U2250 (N_2250,In_1309,In_992);
or U2251 (N_2251,In_165,In_2199);
nor U2252 (N_2252,In_664,In_1368);
nand U2253 (N_2253,In_1489,In_581);
nor U2254 (N_2254,In_1865,In_873);
or U2255 (N_2255,In_117,In_1844);
and U2256 (N_2256,In_1268,In_867);
and U2257 (N_2257,In_1295,In_2069);
nor U2258 (N_2258,In_1406,In_1142);
nor U2259 (N_2259,In_1243,In_1882);
and U2260 (N_2260,In_1925,In_1881);
nand U2261 (N_2261,In_2141,In_390);
nor U2262 (N_2262,In_336,In_1988);
and U2263 (N_2263,In_1324,In_575);
nor U2264 (N_2264,In_884,In_376);
nand U2265 (N_2265,In_1914,In_1054);
nor U2266 (N_2266,In_1859,In_2031);
xnor U2267 (N_2267,In_2476,In_890);
or U2268 (N_2268,In_1611,In_2147);
or U2269 (N_2269,In_347,In_1256);
or U2270 (N_2270,In_1564,In_2162);
or U2271 (N_2271,In_1667,In_1110);
and U2272 (N_2272,In_1721,In_1421);
and U2273 (N_2273,In_1938,In_11);
nand U2274 (N_2274,In_2191,In_2422);
nor U2275 (N_2275,In_2091,In_726);
xor U2276 (N_2276,In_680,In_419);
or U2277 (N_2277,In_939,In_901);
nand U2278 (N_2278,In_879,In_1302);
nor U2279 (N_2279,In_1300,In_2231);
and U2280 (N_2280,In_2133,In_2494);
or U2281 (N_2281,In_2024,In_2048);
and U2282 (N_2282,In_1689,In_408);
nand U2283 (N_2283,In_1154,In_320);
nand U2284 (N_2284,In_1265,In_2172);
and U2285 (N_2285,In_1302,In_865);
nand U2286 (N_2286,In_307,In_2380);
nor U2287 (N_2287,In_1462,In_1645);
and U2288 (N_2288,In_1426,In_190);
nand U2289 (N_2289,In_1748,In_1274);
and U2290 (N_2290,In_660,In_755);
nand U2291 (N_2291,In_160,In_968);
nor U2292 (N_2292,In_371,In_429);
nor U2293 (N_2293,In_1615,In_1983);
nor U2294 (N_2294,In_451,In_959);
nor U2295 (N_2295,In_655,In_1057);
and U2296 (N_2296,In_830,In_630);
nor U2297 (N_2297,In_1937,In_1171);
or U2298 (N_2298,In_2477,In_2402);
and U2299 (N_2299,In_1194,In_401);
nand U2300 (N_2300,In_1833,In_1478);
nor U2301 (N_2301,In_1866,In_285);
xor U2302 (N_2302,In_2256,In_935);
and U2303 (N_2303,In_451,In_2465);
xor U2304 (N_2304,In_1623,In_1203);
nor U2305 (N_2305,In_1059,In_1912);
nand U2306 (N_2306,In_1228,In_1083);
nor U2307 (N_2307,In_2035,In_1400);
nand U2308 (N_2308,In_1582,In_1519);
and U2309 (N_2309,In_1794,In_1838);
xnor U2310 (N_2310,In_876,In_1452);
nand U2311 (N_2311,In_1959,In_2335);
or U2312 (N_2312,In_122,In_299);
xnor U2313 (N_2313,In_927,In_8);
nor U2314 (N_2314,In_889,In_286);
nand U2315 (N_2315,In_11,In_1181);
or U2316 (N_2316,In_372,In_2457);
nor U2317 (N_2317,In_472,In_809);
and U2318 (N_2318,In_1076,In_1621);
nor U2319 (N_2319,In_1493,In_1376);
and U2320 (N_2320,In_21,In_2090);
or U2321 (N_2321,In_1644,In_1045);
or U2322 (N_2322,In_1329,In_193);
or U2323 (N_2323,In_235,In_281);
or U2324 (N_2324,In_601,In_1525);
and U2325 (N_2325,In_840,In_1667);
or U2326 (N_2326,In_2222,In_878);
and U2327 (N_2327,In_2405,In_135);
and U2328 (N_2328,In_621,In_264);
nand U2329 (N_2329,In_2126,In_682);
and U2330 (N_2330,In_2411,In_1792);
and U2331 (N_2331,In_2151,In_2487);
nor U2332 (N_2332,In_263,In_89);
nand U2333 (N_2333,In_1432,In_1221);
and U2334 (N_2334,In_1645,In_761);
xor U2335 (N_2335,In_1490,In_1804);
or U2336 (N_2336,In_515,In_1668);
nor U2337 (N_2337,In_1098,In_2439);
nand U2338 (N_2338,In_8,In_792);
and U2339 (N_2339,In_2259,In_397);
nor U2340 (N_2340,In_1689,In_1112);
or U2341 (N_2341,In_14,In_1058);
and U2342 (N_2342,In_778,In_1606);
or U2343 (N_2343,In_586,In_650);
and U2344 (N_2344,In_817,In_504);
nand U2345 (N_2345,In_598,In_803);
and U2346 (N_2346,In_1924,In_350);
and U2347 (N_2347,In_702,In_2134);
or U2348 (N_2348,In_514,In_448);
or U2349 (N_2349,In_1317,In_1435);
and U2350 (N_2350,In_896,In_2056);
nor U2351 (N_2351,In_2161,In_2377);
or U2352 (N_2352,In_1314,In_202);
nor U2353 (N_2353,In_2118,In_966);
and U2354 (N_2354,In_1880,In_740);
nor U2355 (N_2355,In_2189,In_381);
or U2356 (N_2356,In_1195,In_1273);
and U2357 (N_2357,In_1505,In_942);
and U2358 (N_2358,In_2308,In_1801);
and U2359 (N_2359,In_2015,In_1223);
or U2360 (N_2360,In_1752,In_1285);
nor U2361 (N_2361,In_143,In_1799);
nor U2362 (N_2362,In_1340,In_1182);
nand U2363 (N_2363,In_2287,In_676);
nand U2364 (N_2364,In_2038,In_2104);
nand U2365 (N_2365,In_1229,In_1143);
xnor U2366 (N_2366,In_1079,In_1254);
and U2367 (N_2367,In_2263,In_1194);
or U2368 (N_2368,In_39,In_2208);
nand U2369 (N_2369,In_2193,In_823);
nor U2370 (N_2370,In_300,In_2353);
nor U2371 (N_2371,In_2323,In_1722);
or U2372 (N_2372,In_1504,In_2202);
or U2373 (N_2373,In_1469,In_1967);
or U2374 (N_2374,In_1695,In_347);
nand U2375 (N_2375,In_2447,In_2182);
xnor U2376 (N_2376,In_2328,In_1752);
nor U2377 (N_2377,In_1581,In_2433);
and U2378 (N_2378,In_2294,In_1956);
nand U2379 (N_2379,In_418,In_626);
and U2380 (N_2380,In_1052,In_1724);
xnor U2381 (N_2381,In_748,In_525);
and U2382 (N_2382,In_166,In_1802);
and U2383 (N_2383,In_759,In_258);
and U2384 (N_2384,In_2142,In_822);
or U2385 (N_2385,In_727,In_1802);
nand U2386 (N_2386,In_704,In_1521);
nor U2387 (N_2387,In_1072,In_849);
xor U2388 (N_2388,In_1655,In_102);
xor U2389 (N_2389,In_2390,In_1173);
xnor U2390 (N_2390,In_1595,In_407);
xor U2391 (N_2391,In_1635,In_2096);
xor U2392 (N_2392,In_1041,In_520);
nor U2393 (N_2393,In_2422,In_1247);
nand U2394 (N_2394,In_165,In_21);
and U2395 (N_2395,In_438,In_1720);
or U2396 (N_2396,In_818,In_1666);
nand U2397 (N_2397,In_668,In_2035);
and U2398 (N_2398,In_1236,In_780);
nor U2399 (N_2399,In_1208,In_1615);
xor U2400 (N_2400,In_900,In_1978);
nand U2401 (N_2401,In_2097,In_1061);
nor U2402 (N_2402,In_803,In_476);
nand U2403 (N_2403,In_874,In_1886);
nand U2404 (N_2404,In_856,In_1445);
nand U2405 (N_2405,In_2390,In_1745);
nand U2406 (N_2406,In_1569,In_2499);
nand U2407 (N_2407,In_2414,In_667);
nand U2408 (N_2408,In_1972,In_3);
xor U2409 (N_2409,In_1714,In_894);
nand U2410 (N_2410,In_278,In_957);
nand U2411 (N_2411,In_1400,In_453);
and U2412 (N_2412,In_862,In_1232);
nor U2413 (N_2413,In_1113,In_2474);
or U2414 (N_2414,In_1340,In_1048);
nor U2415 (N_2415,In_611,In_2435);
nor U2416 (N_2416,In_977,In_1029);
nor U2417 (N_2417,In_1706,In_892);
nand U2418 (N_2418,In_696,In_1733);
nand U2419 (N_2419,In_2400,In_2085);
or U2420 (N_2420,In_2460,In_803);
or U2421 (N_2421,In_1620,In_1256);
nand U2422 (N_2422,In_1665,In_1333);
and U2423 (N_2423,In_2419,In_1864);
and U2424 (N_2424,In_1616,In_1585);
nor U2425 (N_2425,In_826,In_1389);
nand U2426 (N_2426,In_1024,In_1395);
nand U2427 (N_2427,In_1024,In_1223);
xor U2428 (N_2428,In_749,In_1276);
nor U2429 (N_2429,In_148,In_779);
xnor U2430 (N_2430,In_1938,In_1325);
nor U2431 (N_2431,In_957,In_1359);
and U2432 (N_2432,In_2080,In_430);
or U2433 (N_2433,In_1228,In_288);
nand U2434 (N_2434,In_2473,In_550);
nand U2435 (N_2435,In_1887,In_1782);
nand U2436 (N_2436,In_1981,In_1195);
nor U2437 (N_2437,In_207,In_2126);
or U2438 (N_2438,In_1956,In_780);
and U2439 (N_2439,In_1080,In_86);
and U2440 (N_2440,In_1961,In_1691);
nor U2441 (N_2441,In_2099,In_1572);
or U2442 (N_2442,In_1050,In_1010);
nand U2443 (N_2443,In_1622,In_2305);
and U2444 (N_2444,In_2284,In_1476);
or U2445 (N_2445,In_1265,In_913);
nor U2446 (N_2446,In_2407,In_1636);
nand U2447 (N_2447,In_455,In_1305);
or U2448 (N_2448,In_729,In_2353);
nor U2449 (N_2449,In_2230,In_2384);
and U2450 (N_2450,In_621,In_2200);
and U2451 (N_2451,In_1639,In_2257);
and U2452 (N_2452,In_1405,In_451);
or U2453 (N_2453,In_41,In_12);
and U2454 (N_2454,In_784,In_1073);
or U2455 (N_2455,In_198,In_484);
nand U2456 (N_2456,In_1970,In_772);
nor U2457 (N_2457,In_449,In_345);
nand U2458 (N_2458,In_717,In_1946);
or U2459 (N_2459,In_70,In_2055);
nor U2460 (N_2460,In_2094,In_2344);
xnor U2461 (N_2461,In_2368,In_502);
nor U2462 (N_2462,In_464,In_1159);
or U2463 (N_2463,In_138,In_226);
xnor U2464 (N_2464,In_1260,In_2299);
nand U2465 (N_2465,In_1195,In_721);
nor U2466 (N_2466,In_1209,In_255);
xor U2467 (N_2467,In_1668,In_2338);
nor U2468 (N_2468,In_1392,In_2332);
xor U2469 (N_2469,In_1279,In_1891);
xnor U2470 (N_2470,In_1071,In_1448);
nand U2471 (N_2471,In_128,In_1210);
nor U2472 (N_2472,In_1664,In_1092);
nand U2473 (N_2473,In_937,In_1282);
nor U2474 (N_2474,In_1109,In_24);
nor U2475 (N_2475,In_2261,In_2152);
or U2476 (N_2476,In_1854,In_1447);
nor U2477 (N_2477,In_490,In_2163);
or U2478 (N_2478,In_2307,In_2405);
or U2479 (N_2479,In_1851,In_2293);
nand U2480 (N_2480,In_158,In_1935);
nand U2481 (N_2481,In_371,In_1543);
or U2482 (N_2482,In_722,In_591);
nor U2483 (N_2483,In_2283,In_1051);
or U2484 (N_2484,In_1608,In_1279);
nor U2485 (N_2485,In_850,In_1669);
and U2486 (N_2486,In_1641,In_656);
and U2487 (N_2487,In_421,In_544);
nand U2488 (N_2488,In_824,In_1503);
or U2489 (N_2489,In_2236,In_1153);
nor U2490 (N_2490,In_2478,In_296);
nand U2491 (N_2491,In_1063,In_923);
and U2492 (N_2492,In_2048,In_1756);
xnor U2493 (N_2493,In_1031,In_117);
nand U2494 (N_2494,In_410,In_740);
nand U2495 (N_2495,In_2204,In_987);
or U2496 (N_2496,In_1486,In_795);
nand U2497 (N_2497,In_952,In_877);
nand U2498 (N_2498,In_2359,In_765);
or U2499 (N_2499,In_258,In_370);
or U2500 (N_2500,N_2456,N_892);
xor U2501 (N_2501,N_1085,N_1942);
and U2502 (N_2502,N_2121,N_1781);
xnor U2503 (N_2503,N_253,N_1151);
nand U2504 (N_2504,N_1928,N_885);
nand U2505 (N_2505,N_1845,N_365);
nor U2506 (N_2506,N_2046,N_1498);
nor U2507 (N_2507,N_837,N_1792);
and U2508 (N_2508,N_1200,N_46);
and U2509 (N_2509,N_567,N_2250);
or U2510 (N_2510,N_91,N_1473);
xnor U2511 (N_2511,N_438,N_718);
or U2512 (N_2512,N_244,N_785);
and U2513 (N_2513,N_2099,N_2461);
or U2514 (N_2514,N_2203,N_650);
and U2515 (N_2515,N_385,N_2404);
xnor U2516 (N_2516,N_345,N_1884);
or U2517 (N_2517,N_1423,N_1376);
nor U2518 (N_2518,N_1240,N_1970);
and U2519 (N_2519,N_1869,N_443);
and U2520 (N_2520,N_80,N_2395);
nand U2521 (N_2521,N_2268,N_762);
nor U2522 (N_2522,N_1474,N_790);
or U2523 (N_2523,N_2146,N_1715);
xnor U2524 (N_2524,N_208,N_423);
or U2525 (N_2525,N_2154,N_1433);
or U2526 (N_2526,N_2051,N_301);
nor U2527 (N_2527,N_842,N_479);
and U2528 (N_2528,N_2297,N_2366);
nand U2529 (N_2529,N_2439,N_461);
nor U2530 (N_2530,N_867,N_1176);
or U2531 (N_2531,N_865,N_1594);
nand U2532 (N_2532,N_1686,N_1401);
nor U2533 (N_2533,N_2091,N_1698);
xor U2534 (N_2534,N_2306,N_575);
or U2535 (N_2535,N_84,N_2227);
xnor U2536 (N_2536,N_2024,N_2133);
nor U2537 (N_2537,N_1757,N_1952);
or U2538 (N_2538,N_2440,N_994);
and U2539 (N_2539,N_1231,N_529);
nor U2540 (N_2540,N_145,N_1770);
or U2541 (N_2541,N_116,N_1662);
nor U2542 (N_2542,N_69,N_1491);
nand U2543 (N_2543,N_792,N_1724);
xor U2544 (N_2544,N_1890,N_760);
nand U2545 (N_2545,N_2428,N_176);
xnor U2546 (N_2546,N_2073,N_452);
or U2547 (N_2547,N_2482,N_2271);
nor U2548 (N_2548,N_1456,N_36);
or U2549 (N_2549,N_1917,N_808);
and U2550 (N_2550,N_1935,N_2067);
xnor U2551 (N_2551,N_2446,N_696);
xnor U2552 (N_2552,N_2131,N_2334);
xnor U2553 (N_2553,N_2122,N_1650);
and U2554 (N_2554,N_1112,N_511);
nand U2555 (N_2555,N_197,N_1824);
nor U2556 (N_2556,N_802,N_94);
and U2557 (N_2557,N_1398,N_1145);
and U2558 (N_2558,N_2052,N_1087);
xnor U2559 (N_2559,N_1056,N_1199);
nand U2560 (N_2560,N_150,N_2264);
or U2561 (N_2561,N_75,N_1697);
nand U2562 (N_2562,N_2295,N_1225);
nand U2563 (N_2563,N_24,N_2350);
nand U2564 (N_2564,N_1572,N_1321);
nor U2565 (N_2565,N_630,N_2090);
and U2566 (N_2566,N_1033,N_49);
nor U2567 (N_2567,N_2173,N_1064);
and U2568 (N_2568,N_106,N_1124);
or U2569 (N_2569,N_1834,N_1731);
and U2570 (N_2570,N_1624,N_68);
or U2571 (N_2571,N_1946,N_1180);
or U2572 (N_2572,N_1341,N_1072);
or U2573 (N_2573,N_1214,N_196);
nor U2574 (N_2574,N_2362,N_1611);
or U2575 (N_2575,N_499,N_1919);
nand U2576 (N_2576,N_2465,N_2151);
or U2577 (N_2577,N_535,N_1162);
nand U2578 (N_2578,N_974,N_1999);
nand U2579 (N_2579,N_1493,N_2347);
nand U2580 (N_2580,N_2088,N_1931);
nand U2581 (N_2581,N_1837,N_1522);
xnor U2582 (N_2582,N_912,N_827);
or U2583 (N_2583,N_1796,N_891);
nor U2584 (N_2584,N_305,N_829);
nor U2585 (N_2585,N_192,N_336);
nand U2586 (N_2586,N_218,N_1964);
nor U2587 (N_2587,N_2235,N_262);
nand U2588 (N_2588,N_360,N_2008);
or U2589 (N_2589,N_991,N_1872);
nand U2590 (N_2590,N_1562,N_2269);
or U2591 (N_2591,N_772,N_163);
and U2592 (N_2592,N_662,N_77);
or U2593 (N_2593,N_520,N_1722);
and U2594 (N_2594,N_430,N_1909);
nand U2595 (N_2595,N_1308,N_2244);
or U2596 (N_2596,N_623,N_694);
nand U2597 (N_2597,N_1971,N_1404);
nor U2598 (N_2598,N_1568,N_1143);
nand U2599 (N_2599,N_1218,N_1879);
or U2600 (N_2600,N_1868,N_1209);
nand U2601 (N_2601,N_1313,N_1523);
nor U2602 (N_2602,N_2260,N_2400);
or U2603 (N_2603,N_126,N_1735);
or U2604 (N_2604,N_228,N_1860);
and U2605 (N_2605,N_844,N_55);
or U2606 (N_2606,N_560,N_1179);
and U2607 (N_2607,N_2031,N_1476);
nand U2608 (N_2608,N_45,N_321);
nand U2609 (N_2609,N_1751,N_1047);
nor U2610 (N_2610,N_731,N_1853);
nand U2611 (N_2611,N_841,N_801);
nor U2612 (N_2612,N_1488,N_803);
or U2613 (N_2613,N_564,N_2246);
nand U2614 (N_2614,N_1628,N_2323);
xor U2615 (N_2615,N_516,N_21);
nor U2616 (N_2616,N_1435,N_2174);
and U2617 (N_2617,N_328,N_750);
nor U2618 (N_2618,N_298,N_1670);
nand U2619 (N_2619,N_1227,N_1621);
nor U2620 (N_2620,N_971,N_99);
nor U2621 (N_2621,N_189,N_1497);
nor U2622 (N_2622,N_1323,N_2191);
and U2623 (N_2623,N_1627,N_2218);
or U2624 (N_2624,N_2374,N_763);
and U2625 (N_2625,N_20,N_2201);
nand U2626 (N_2626,N_2460,N_166);
nand U2627 (N_2627,N_1986,N_645);
or U2628 (N_2628,N_775,N_1876);
and U2629 (N_2629,N_1635,N_1017);
or U2630 (N_2630,N_2365,N_1472);
nor U2631 (N_2631,N_471,N_2345);
nor U2632 (N_2632,N_1893,N_1446);
nand U2633 (N_2633,N_528,N_2305);
nand U2634 (N_2634,N_181,N_1949);
xor U2635 (N_2635,N_1267,N_1338);
or U2636 (N_2636,N_275,N_1190);
and U2637 (N_2637,N_2050,N_1330);
nor U2638 (N_2638,N_437,N_1120);
nand U2639 (N_2639,N_2065,N_2022);
nand U2640 (N_2640,N_691,N_1492);
or U2641 (N_2641,N_723,N_389);
nor U2642 (N_2642,N_463,N_727);
and U2643 (N_2643,N_2032,N_2125);
nor U2644 (N_2644,N_911,N_935);
nand U2645 (N_2645,N_2495,N_513);
nand U2646 (N_2646,N_2445,N_2005);
nor U2647 (N_2647,N_2221,N_507);
nand U2648 (N_2648,N_2182,N_2128);
or U2649 (N_2649,N_919,N_120);
nand U2650 (N_2650,N_2288,N_669);
nand U2651 (N_2651,N_473,N_2381);
nor U2652 (N_2652,N_561,N_2416);
nor U2653 (N_2653,N_1546,N_1383);
or U2654 (N_2654,N_1743,N_2123);
nor U2655 (N_2655,N_2393,N_647);
and U2656 (N_2656,N_1694,N_2486);
nor U2657 (N_2657,N_2226,N_1010);
nor U2658 (N_2658,N_558,N_1082);
or U2659 (N_2659,N_586,N_810);
xor U2660 (N_2660,N_1977,N_1263);
and U2661 (N_2661,N_619,N_825);
and U2662 (N_2662,N_2037,N_1244);
nand U2663 (N_2663,N_1726,N_285);
and U2664 (N_2664,N_1517,N_1717);
nand U2665 (N_2665,N_2144,N_2292);
xor U2666 (N_2666,N_362,N_428);
or U2667 (N_2667,N_973,N_2224);
xor U2668 (N_2668,N_1030,N_1987);
nand U2669 (N_2669,N_703,N_514);
nand U2670 (N_2670,N_2443,N_1885);
and U2671 (N_2671,N_1141,N_1235);
nor U2672 (N_2672,N_1891,N_2337);
nand U2673 (N_2673,N_2136,N_1956);
nand U2674 (N_2674,N_2296,N_308);
nor U2675 (N_2675,N_1318,N_533);
or U2676 (N_2676,N_1560,N_2332);
or U2677 (N_2677,N_933,N_1291);
and U2678 (N_2678,N_1368,N_1453);
nor U2679 (N_2679,N_554,N_927);
nor U2680 (N_2680,N_1671,N_2220);
xor U2681 (N_2681,N_1927,N_313);
or U2682 (N_2682,N_1565,N_241);
or U2683 (N_2683,N_2243,N_877);
nor U2684 (N_2684,N_2336,N_2259);
and U2685 (N_2685,N_1979,N_141);
or U2686 (N_2686,N_1596,N_2343);
nor U2687 (N_2687,N_777,N_1312);
and U2688 (N_2688,N_1669,N_1302);
nand U2689 (N_2689,N_483,N_1035);
nor U2690 (N_2690,N_1096,N_331);
and U2691 (N_2691,N_980,N_1349);
nand U2692 (N_2692,N_2496,N_2265);
or U2693 (N_2693,N_1483,N_913);
or U2694 (N_2694,N_2326,N_127);
or U2695 (N_2695,N_1679,N_2459);
xnor U2696 (N_2696,N_422,N_1823);
and U2697 (N_2697,N_782,N_118);
or U2698 (N_2698,N_2000,N_171);
and U2699 (N_2699,N_1363,N_2344);
nor U2700 (N_2700,N_1486,N_323);
or U2701 (N_2701,N_491,N_43);
nor U2702 (N_2702,N_311,N_314);
nand U2703 (N_2703,N_569,N_322);
or U2704 (N_2704,N_1926,N_2442);
nand U2705 (N_2705,N_229,N_5);
nand U2706 (N_2706,N_1672,N_713);
nand U2707 (N_2707,N_1236,N_1591);
and U2708 (N_2708,N_1391,N_2255);
and U2709 (N_2709,N_1829,N_1188);
and U2710 (N_2710,N_294,N_2066);
xnor U2711 (N_2711,N_1393,N_690);
nand U2712 (N_2712,N_1520,N_2383);
and U2713 (N_2713,N_1646,N_636);
xor U2714 (N_2714,N_1347,N_2029);
nand U2715 (N_2715,N_901,N_1582);
nand U2716 (N_2716,N_699,N_1097);
and U2717 (N_2717,N_888,N_532);
nor U2718 (N_2718,N_2207,N_1642);
or U2719 (N_2719,N_2248,N_125);
and U2720 (N_2720,N_1693,N_1816);
nor U2721 (N_2721,N_194,N_917);
nor U2722 (N_2722,N_361,N_1502);
xnor U2723 (N_2723,N_2168,N_2150);
nand U2724 (N_2724,N_1563,N_185);
or U2725 (N_2725,N_1873,N_993);
nand U2726 (N_2726,N_2450,N_540);
nor U2727 (N_2727,N_2223,N_269);
nor U2728 (N_2728,N_642,N_2233);
xor U2729 (N_2729,N_2194,N_1586);
or U2730 (N_2730,N_905,N_245);
nor U2731 (N_2731,N_2072,N_1471);
nand U2732 (N_2732,N_2256,N_2078);
nor U2733 (N_2733,N_1083,N_1864);
xnor U2734 (N_2734,N_859,N_1791);
nor U2735 (N_2735,N_2307,N_1988);
nand U2736 (N_2736,N_1299,N_2373);
and U2737 (N_2737,N_136,N_1108);
nor U2738 (N_2738,N_498,N_286);
and U2739 (N_2739,N_1754,N_1602);
nand U2740 (N_2740,N_338,N_2308);
xor U2741 (N_2741,N_2097,N_1265);
or U2742 (N_2742,N_793,N_488);
xor U2743 (N_2743,N_2143,N_1548);
and U2744 (N_2744,N_1392,N_1929);
nor U2745 (N_2745,N_2180,N_1610);
nand U2746 (N_2746,N_2270,N_644);
xnor U2747 (N_2747,N_1232,N_129);
nor U2748 (N_2748,N_2464,N_969);
xnor U2749 (N_2749,N_2011,N_661);
nor U2750 (N_2750,N_109,N_1794);
nand U2751 (N_2751,N_1266,N_555);
or U2752 (N_2752,N_2145,N_2274);
or U2753 (N_2753,N_640,N_1558);
or U2754 (N_2754,N_697,N_2363);
or U2755 (N_2755,N_755,N_2176);
or U2756 (N_2756,N_1273,N_2367);
xor U2757 (N_2757,N_1215,N_1477);
and U2758 (N_2758,N_392,N_1380);
or U2759 (N_2759,N_1793,N_1003);
and U2760 (N_2760,N_2184,N_1783);
and U2761 (N_2761,N_1128,N_909);
or U2762 (N_2762,N_942,N_1555);
nand U2763 (N_2763,N_930,N_907);
or U2764 (N_2764,N_2245,N_273);
nor U2765 (N_2765,N_603,N_1766);
nor U2766 (N_2766,N_1556,N_17);
nor U2767 (N_2767,N_1101,N_387);
nor U2768 (N_2768,N_1311,N_455);
nand U2769 (N_2769,N_578,N_850);
or U2770 (N_2770,N_1482,N_964);
and U2771 (N_2771,N_1746,N_303);
nand U2772 (N_2772,N_626,N_2009);
and U2773 (N_2773,N_2480,N_284);
or U2774 (N_2774,N_1198,N_1216);
nor U2775 (N_2775,N_27,N_340);
nor U2776 (N_2776,N_2441,N_2199);
or U2777 (N_2777,N_468,N_620);
nor U2778 (N_2778,N_503,N_610);
and U2779 (N_2779,N_960,N_1584);
or U2780 (N_2780,N_482,N_18);
nand U2781 (N_2781,N_710,N_1489);
nand U2782 (N_2782,N_724,N_2198);
xor U2783 (N_2783,N_2148,N_2010);
nand U2784 (N_2784,N_1664,N_799);
and U2785 (N_2785,N_958,N_193);
and U2786 (N_2786,N_1786,N_306);
nand U2787 (N_2787,N_1161,N_2474);
nor U2788 (N_2788,N_735,N_1090);
or U2789 (N_2789,N_2061,N_1840);
nand U2790 (N_2790,N_1408,N_2408);
nand U2791 (N_2791,N_1171,N_2215);
or U2792 (N_2792,N_1126,N_1674);
xor U2793 (N_2793,N_2386,N_998);
xnor U2794 (N_2794,N_824,N_131);
xnor U2795 (N_2795,N_725,N_1819);
and U2796 (N_2796,N_490,N_1593);
nand U2797 (N_2797,N_769,N_2102);
and U2798 (N_2798,N_1666,N_1057);
nand U2799 (N_2799,N_2453,N_1012);
xor U2800 (N_2800,N_1682,N_233);
and U2801 (N_2801,N_231,N_1177);
nor U2802 (N_2802,N_1278,N_265);
nor U2803 (N_2803,N_1098,N_2272);
or U2804 (N_2804,N_1881,N_652);
nor U2805 (N_2805,N_1129,N_1851);
nand U2806 (N_2806,N_1982,N_2411);
nand U2807 (N_2807,N_1071,N_1470);
nor U2808 (N_2808,N_1677,N_1613);
nor U2809 (N_2809,N_1619,N_1510);
and U2810 (N_2810,N_1153,N_1737);
nor U2811 (N_2811,N_2019,N_874);
nor U2812 (N_2812,N_2045,N_1902);
nor U2813 (N_2813,N_1683,N_472);
or U2814 (N_2814,N_1822,N_1925);
nand U2815 (N_2815,N_58,N_2396);
nand U2816 (N_2816,N_604,N_2406);
xnor U2817 (N_2817,N_1078,N_1243);
or U2818 (N_2818,N_1248,N_870);
or U2819 (N_2819,N_1695,N_1196);
nand U2820 (N_2820,N_1821,N_665);
and U2821 (N_2821,N_315,N_1798);
or U2822 (N_2822,N_2415,N_133);
nor U2823 (N_2823,N_2095,N_2462);
or U2824 (N_2824,N_1575,N_1343);
or U2825 (N_2825,N_2432,N_2290);
or U2826 (N_2826,N_1040,N_1849);
or U2827 (N_2827,N_948,N_1833);
or U2828 (N_2828,N_41,N_1967);
xnor U2829 (N_2829,N_2025,N_1797);
nand U2830 (N_2830,N_2322,N_2285);
nand U2831 (N_2831,N_419,N_809);
nand U2832 (N_2832,N_2401,N_1385);
nand U2833 (N_2833,N_97,N_148);
or U2834 (N_2834,N_481,N_325);
nor U2835 (N_2835,N_2457,N_1533);
nand U2836 (N_2836,N_119,N_2124);
or U2837 (N_2837,N_2298,N_1888);
or U2838 (N_2838,N_796,N_1194);
xnor U2839 (N_2839,N_74,N_289);
and U2840 (N_2840,N_749,N_344);
or U2841 (N_2841,N_2449,N_952);
nor U2842 (N_2842,N_2080,N_1300);
nand U2843 (N_2843,N_582,N_847);
and U2844 (N_2844,N_932,N_2049);
nand U2845 (N_2845,N_547,N_153);
nand U2846 (N_2846,N_1687,N_7);
nand U2847 (N_2847,N_1808,N_1142);
or U2848 (N_2848,N_2166,N_202);
nand U2849 (N_2849,N_1675,N_2488);
nand U2850 (N_2850,N_1564,N_1720);
and U2851 (N_2851,N_2342,N_2360);
or U2852 (N_2852,N_538,N_2284);
nand U2853 (N_2853,N_1636,N_2351);
nand U2854 (N_2854,N_967,N_895);
nor U2855 (N_2855,N_1855,N_266);
or U2856 (N_2856,N_54,N_1756);
xnor U2857 (N_2857,N_1105,N_2093);
nand U2858 (N_2858,N_1629,N_134);
nand U2859 (N_2859,N_62,N_1782);
nand U2860 (N_2860,N_1414,N_1282);
and U2861 (N_2861,N_786,N_754);
nor U2862 (N_2862,N_1723,N_254);
and U2863 (N_2863,N_2179,N_82);
nor U2864 (N_2864,N_1478,N_649);
nand U2865 (N_2865,N_2079,N_2013);
and U2866 (N_2866,N_409,N_343);
nor U2867 (N_2867,N_878,N_648);
nand U2868 (N_2868,N_217,N_1961);
nand U2869 (N_2869,N_1053,N_383);
nand U2870 (N_2870,N_1966,N_34);
nor U2871 (N_2871,N_1883,N_1760);
nor U2872 (N_2872,N_1689,N_2289);
xnor U2873 (N_2873,N_1043,N_1547);
nor U2874 (N_2874,N_1439,N_1137);
or U2875 (N_2875,N_2325,N_168);
nand U2876 (N_2876,N_2472,N_2071);
nor U2877 (N_2877,N_1789,N_2254);
xor U2878 (N_2878,N_2475,N_1277);
xor U2879 (N_2879,N_130,N_1415);
and U2880 (N_2880,N_1866,N_2253);
and U2881 (N_2881,N_1981,N_248);
and U2882 (N_2882,N_1202,N_203);
or U2883 (N_2883,N_819,N_1984);
and U2884 (N_2884,N_820,N_549);
nor U2885 (N_2885,N_1023,N_2109);
nand U2886 (N_2886,N_1444,N_1150);
and U2887 (N_2887,N_1131,N_397);
nor U2888 (N_2888,N_1660,N_1752);
xor U2889 (N_2889,N_1940,N_2170);
nor U2890 (N_2890,N_1634,N_2329);
and U2891 (N_2891,N_1577,N_2320);
or U2892 (N_2892,N_2476,N_2229);
and U2893 (N_2893,N_2007,N_707);
or U2894 (N_2894,N_1711,N_2435);
nand U2895 (N_2895,N_2081,N_92);
or U2896 (N_2896,N_377,N_413);
nand U2897 (N_2897,N_295,N_530);
or U2898 (N_2898,N_1146,N_1951);
nand U2899 (N_2899,N_2478,N_1750);
or U2900 (N_2900,N_1088,N_950);
or U2901 (N_2901,N_1309,N_87);
xnor U2902 (N_2902,N_2068,N_276);
or U2903 (N_2903,N_962,N_210);
and U2904 (N_2904,N_704,N_2135);
and U2905 (N_2905,N_2370,N_1348);
nor U2906 (N_2906,N_287,N_559);
or U2907 (N_2907,N_1425,N_1732);
and U2908 (N_2908,N_1136,N_2479);
nand U2909 (N_2909,N_1827,N_1799);
or U2910 (N_2910,N_1297,N_386);
and U2911 (N_2911,N_519,N_988);
and U2912 (N_2912,N_1587,N_326);
nor U2913 (N_2913,N_1405,N_711);
nor U2914 (N_2914,N_271,N_444);
nand U2915 (N_2915,N_467,N_2222);
or U2916 (N_2916,N_2341,N_931);
or U2917 (N_2917,N_897,N_348);
nor U2918 (N_2918,N_2043,N_1595);
nor U2919 (N_2919,N_631,N_1241);
nor U2920 (N_2920,N_2156,N_2056);
or U2921 (N_2921,N_251,N_2277);
and U2922 (N_2922,N_1490,N_1164);
nor U2923 (N_2923,N_1997,N_596);
nor U2924 (N_2924,N_1815,N_1653);
and U2925 (N_2925,N_1597,N_1549);
nor U2926 (N_2926,N_651,N_2487);
nand U2927 (N_2927,N_140,N_476);
nor U2928 (N_2928,N_1804,N_1052);
nor U2929 (N_2929,N_1173,N_1361);
nand U2930 (N_2930,N_702,N_427);
nand U2931 (N_2931,N_1411,N_2282);
nand U2932 (N_2932,N_2060,N_2369);
or U2933 (N_2933,N_1109,N_22);
xor U2934 (N_2934,N_436,N_1734);
or U2935 (N_2935,N_291,N_1514);
nand U2936 (N_2936,N_42,N_1197);
nand U2937 (N_2937,N_2177,N_599);
nor U2938 (N_2938,N_4,N_1485);
nand U2939 (N_2939,N_2437,N_65);
nand U2940 (N_2940,N_2020,N_2433);
nor U2941 (N_2941,N_128,N_2152);
or U2942 (N_2942,N_1065,N_1328);
nor U2943 (N_2943,N_1279,N_102);
nand U2944 (N_2944,N_1592,N_1692);
and U2945 (N_2945,N_2448,N_1989);
nor U2946 (N_2946,N_1887,N_910);
and U2947 (N_2947,N_545,N_2267);
or U2948 (N_2948,N_1326,N_1727);
nor U2949 (N_2949,N_1460,N_791);
and U2950 (N_2950,N_1357,N_678);
xor U2951 (N_2951,N_180,N_1443);
or U2952 (N_2952,N_274,N_1008);
nand U2953 (N_2953,N_2236,N_66);
xor U2954 (N_2954,N_2263,N_2249);
or U2955 (N_2955,N_454,N_1095);
or U2956 (N_2956,N_1973,N_2202);
nor U2957 (N_2957,N_1974,N_1283);
nand U2958 (N_2958,N_399,N_671);
nor U2959 (N_2959,N_2162,N_1748);
nand U2960 (N_2960,N_1422,N_637);
nand U2961 (N_2961,N_435,N_1285);
or U2962 (N_2962,N_990,N_811);
and U2963 (N_2963,N_2064,N_469);
and U2964 (N_2964,N_903,N_2075);
nand U2965 (N_2965,N_1599,N_470);
and U2966 (N_2966,N_961,N_1813);
or U2967 (N_2967,N_239,N_1707);
or U2968 (N_2968,N_1479,N_687);
nand U2969 (N_2969,N_450,N_812);
nand U2970 (N_2970,N_2252,N_1573);
nor U2971 (N_2971,N_1980,N_542);
and U2972 (N_2972,N_1219,N_2210);
nand U2973 (N_2973,N_2158,N_981);
and U2974 (N_2974,N_936,N_999);
and U2975 (N_2975,N_400,N_926);
xnor U2976 (N_2976,N_915,N_105);
nand U2977 (N_2977,N_1144,N_833);
or U2978 (N_2978,N_822,N_283);
and U2979 (N_2979,N_2407,N_807);
nor U2980 (N_2980,N_1969,N_2193);
or U2981 (N_2981,N_2103,N_1696);
nor U2982 (N_2982,N_12,N_924);
nor U2983 (N_2983,N_746,N_1284);
xor U2984 (N_2984,N_1544,N_366);
or U2985 (N_2985,N_1432,N_453);
or U2986 (N_2986,N_162,N_1644);
nand U2987 (N_2987,N_868,N_235);
nand U2988 (N_2988,N_568,N_351);
nand U2989 (N_2989,N_1738,N_573);
nand U2990 (N_2990,N_714,N_508);
nor U2991 (N_2991,N_1749,N_2016);
xnor U2992 (N_2992,N_1509,N_712);
nor U2993 (N_2993,N_541,N_206);
and U2994 (N_2994,N_1086,N_609);
xor U2995 (N_2995,N_2074,N_1907);
nand U2996 (N_2996,N_1805,N_2012);
and U2997 (N_2997,N_1863,N_1739);
nand U2998 (N_2998,N_159,N_1512);
nand U2999 (N_2999,N_302,N_641);
or U3000 (N_3000,N_2028,N_737);
and U3001 (N_3001,N_2409,N_2498);
and U3002 (N_3002,N_494,N_738);
and U3003 (N_3003,N_1647,N_462);
or U3004 (N_3004,N_989,N_1138);
or U3005 (N_3005,N_686,N_1388);
nand U3006 (N_3006,N_1015,N_2317);
nor U3007 (N_3007,N_2328,N_869);
or U3008 (N_3008,N_184,N_1645);
nor U3009 (N_3009,N_1480,N_904);
and U3010 (N_3010,N_2262,N_247);
xnor U3011 (N_3011,N_615,N_1002);
and U3012 (N_3012,N_1776,N_1220);
and U3013 (N_3013,N_1615,N_1788);
or U3014 (N_3014,N_2331,N_1113);
and U3015 (N_3015,N_67,N_1367);
or U3016 (N_3016,N_855,N_527);
and U3017 (N_3017,N_2116,N_584);
nand U3018 (N_3018,N_589,N_2057);
nand U3019 (N_3019,N_2380,N_1046);
or U3020 (N_3020,N_766,N_1036);
and U3021 (N_3021,N_1747,N_2276);
or U3022 (N_3022,N_1933,N_1920);
or U3023 (N_3023,N_618,N_779);
or U3024 (N_3024,N_2107,N_2055);
and U3025 (N_3025,N_838,N_595);
nor U3026 (N_3026,N_149,N_174);
and U3027 (N_3027,N_1571,N_621);
and U3028 (N_3028,N_1018,N_451);
and U3029 (N_3029,N_384,N_975);
nand U3030 (N_3030,N_299,N_2159);
and U3031 (N_3031,N_622,N_200);
or U3032 (N_3032,N_1580,N_1614);
and U3033 (N_3033,N_2204,N_1945);
nand U3034 (N_3034,N_1254,N_1331);
xor U3035 (N_3035,N_222,N_1184);
nor U3036 (N_3036,N_2291,N_466);
xnor U3037 (N_3037,N_1908,N_2033);
nand U3038 (N_3038,N_1317,N_2197);
nand U3039 (N_3039,N_2161,N_2398);
or U3040 (N_3040,N_2117,N_401);
and U3041 (N_3041,N_590,N_1000);
or U3042 (N_3042,N_1394,N_2104);
nor U3043 (N_3043,N_272,N_729);
nor U3044 (N_3044,N_1778,N_2063);
or U3045 (N_3045,N_1539,N_976);
xor U3046 (N_3046,N_278,N_1042);
xor U3047 (N_3047,N_259,N_2232);
and U3048 (N_3048,N_1402,N_30);
nand U3049 (N_3049,N_6,N_1532);
and U3050 (N_3050,N_744,N_2038);
and U3051 (N_3051,N_1685,N_534);
xor U3052 (N_3052,N_1772,N_591);
nand U3053 (N_3053,N_487,N_236);
and U3054 (N_3054,N_1941,N_1237);
nand U3055 (N_3055,N_1839,N_525);
xor U3056 (N_3056,N_633,N_1238);
and U3057 (N_3057,N_495,N_937);
nor U3058 (N_3058,N_1775,N_550);
or U3059 (N_3059,N_1178,N_1205);
and U3060 (N_3060,N_398,N_164);
nand U3061 (N_3061,N_1431,N_363);
nor U3062 (N_3062,N_318,N_2083);
nand U3063 (N_3063,N_1167,N_2466);
or U3064 (N_3064,N_64,N_390);
or U3065 (N_3065,N_1354,N_1276);
and U3066 (N_3066,N_1079,N_380);
xor U3067 (N_3067,N_1475,N_1352);
nand U3068 (N_3068,N_1574,N_1700);
or U3069 (N_3069,N_370,N_2169);
and U3070 (N_3070,N_1350,N_2389);
and U3071 (N_3071,N_38,N_660);
nand U3072 (N_3072,N_1430,N_1160);
nand U3073 (N_3073,N_1260,N_611);
and U3074 (N_3074,N_1007,N_155);
nor U3075 (N_3075,N_1044,N_195);
and U3076 (N_3076,N_1608,N_2413);
or U3077 (N_3077,N_979,N_115);
and U3078 (N_3078,N_1419,N_1806);
and U3079 (N_3079,N_339,N_1857);
or U3080 (N_3080,N_1356,N_682);
or U3081 (N_3081,N_1561,N_1742);
nand U3082 (N_3082,N_1364,N_1487);
nor U3083 (N_3083,N_316,N_2436);
and U3084 (N_3084,N_1985,N_448);
xnor U3085 (N_3085,N_1820,N_1800);
nor U3086 (N_3086,N_1875,N_941);
nand U3087 (N_3087,N_1690,N_743);
xnor U3088 (N_3088,N_656,N_393);
xor U3089 (N_3089,N_261,N_1346);
or U3090 (N_3090,N_1631,N_1027);
and U3091 (N_3091,N_212,N_1758);
xnor U3092 (N_3092,N_1972,N_290);
and U3093 (N_3093,N_138,N_2340);
xnor U3094 (N_3094,N_681,N_1515);
and U3095 (N_3095,N_1465,N_970);
nand U3096 (N_3096,N_2452,N_2094);
nor U3097 (N_3097,N_1089,N_1080);
nor U3098 (N_3098,N_1858,N_1103);
and U3099 (N_3099,N_783,N_689);
nand U3100 (N_3100,N_1421,N_402);
and U3101 (N_3101,N_1484,N_854);
or U3102 (N_3102,N_1626,N_396);
or U3103 (N_3103,N_2394,N_2257);
nand U3104 (N_3104,N_2178,N_2004);
nand U3105 (N_3105,N_1084,N_1074);
and U3106 (N_3106,N_1763,N_814);
and U3107 (N_3107,N_2149,N_280);
xnor U3108 (N_3108,N_882,N_794);
nand U3109 (N_3109,N_858,N_597);
xnor U3110 (N_3110,N_2120,N_1247);
or U3111 (N_3111,N_581,N_110);
nor U3112 (N_3112,N_182,N_983);
xor U3113 (N_3113,N_2412,N_307);
and U3114 (N_3114,N_1125,N_2467);
nand U3115 (N_3115,N_2247,N_2217);
nand U3116 (N_3116,N_1287,N_2077);
nand U3117 (N_3117,N_1332,N_1428);
and U3118 (N_3118,N_2132,N_1104);
and U3119 (N_3119,N_1665,N_433);
and U3120 (N_3120,N_1950,N_417);
and U3121 (N_3121,N_1803,N_1680);
nor U3122 (N_3122,N_740,N_1191);
nand U3123 (N_3123,N_2208,N_1990);
or U3124 (N_3124,N_1229,N_1550);
or U3125 (N_3125,N_949,N_2147);
nand U3126 (N_3126,N_1704,N_1617);
nand U3127 (N_3127,N_943,N_2183);
or U3128 (N_3128,N_1259,N_1452);
nor U3129 (N_3129,N_408,N_373);
nand U3130 (N_3130,N_1850,N_1921);
nor U3131 (N_3131,N_1506,N_1169);
nor U3132 (N_3132,N_161,N_679);
or U3133 (N_3133,N_2027,N_632);
and U3134 (N_3134,N_492,N_1944);
or U3135 (N_3135,N_1451,N_1228);
or U3136 (N_3136,N_1068,N_1848);
or U3137 (N_3137,N_1516,N_1832);
or U3138 (N_3138,N_918,N_1659);
or U3139 (N_3139,N_1947,N_1802);
and U3140 (N_3140,N_288,N_557);
nor U3141 (N_3141,N_57,N_101);
nand U3142 (N_3142,N_1269,N_1306);
or U3143 (N_3143,N_1959,N_925);
nand U3144 (N_3144,N_1154,N_1390);
and U3145 (N_3145,N_281,N_122);
or U3146 (N_3146,N_1301,N_1272);
nor U3147 (N_3147,N_1339,N_1994);
and U3148 (N_3148,N_2089,N_2110);
xnor U3149 (N_3149,N_2304,N_2481);
and U3150 (N_3150,N_353,N_1569);
nor U3151 (N_3151,N_1050,N_1530);
nor U3152 (N_3152,N_1825,N_1983);
or U3153 (N_3153,N_173,N_1359);
and U3154 (N_3154,N_2405,N_172);
xnor U3155 (N_3155,N_2001,N_889);
nor U3156 (N_3156,N_2364,N_1609);
xor U3157 (N_3157,N_226,N_627);
and U3158 (N_3158,N_1384,N_1355);
xnor U3159 (N_3159,N_188,N_1566);
xor U3160 (N_3160,N_2115,N_14);
or U3161 (N_3161,N_426,N_2113);
or U3162 (N_3162,N_79,N_83);
xnor U3163 (N_3163,N_745,N_1434);
or U3164 (N_3164,N_1537,N_2108);
nand U3165 (N_3165,N_685,N_152);
and U3166 (N_3166,N_2041,N_2098);
and U3167 (N_3167,N_1705,N_376);
nor U3168 (N_3168,N_1324,N_672);
xnor U3169 (N_3169,N_1841,N_1930);
or U3170 (N_3170,N_1242,N_391);
xor U3171 (N_3171,N_1127,N_350);
or U3172 (N_3172,N_1004,N_898);
nor U3173 (N_3173,N_2356,N_310);
and U3174 (N_3174,N_1133,N_1761);
xnor U3175 (N_3175,N_2188,N_2181);
xor U3176 (N_3176,N_1632,N_1641);
nor U3177 (N_3177,N_853,N_2358);
nor U3178 (N_3178,N_1344,N_1892);
nand U3179 (N_3179,N_953,N_1462);
or U3180 (N_3180,N_985,N_1836);
nand U3181 (N_3181,N_670,N_1026);
nand U3182 (N_3182,N_593,N_178);
nand U3183 (N_3183,N_170,N_1389);
nor U3184 (N_3184,N_59,N_1094);
and U3185 (N_3185,N_1261,N_1831);
or U3186 (N_3186,N_1396,N_583);
and U3187 (N_3187,N_1045,N_135);
xor U3188 (N_3188,N_1441,N_1454);
nor U3189 (N_3189,N_2126,N_1062);
nand U3190 (N_3190,N_404,N_548);
nor U3191 (N_3191,N_1013,N_1115);
nand U3192 (N_3192,N_1406,N_1852);
or U3193 (N_3193,N_566,N_2421);
or U3194 (N_3194,N_705,N_1304);
nor U3195 (N_3195,N_861,N_938);
xor U3196 (N_3196,N_412,N_1871);
xor U3197 (N_3197,N_612,N_2138);
nor U3198 (N_3198,N_250,N_1811);
nor U3199 (N_3199,N_2458,N_1867);
nand U3200 (N_3200,N_1449,N_571);
xnor U3201 (N_3201,N_1499,N_249);
nand U3202 (N_3202,N_1135,N_2361);
and U3203 (N_3203,N_50,N_506);
or U3204 (N_3204,N_81,N_922);
and U3205 (N_3205,N_332,N_562);
xnor U3206 (N_3206,N_1965,N_716);
xor U3207 (N_3207,N_1440,N_1870);
nand U3208 (N_3208,N_420,N_2251);
and U3209 (N_3209,N_977,N_1102);
nor U3210 (N_3210,N_337,N_1733);
or U3211 (N_3211,N_800,N_1365);
nor U3212 (N_3212,N_165,N_1121);
nand U3213 (N_3213,N_1897,N_1729);
and U3214 (N_3214,N_1336,N_1787);
nand U3215 (N_3215,N_1777,N_2266);
nand U3216 (N_3216,N_1320,N_1536);
or U3217 (N_3217,N_1256,N_515);
nand U3218 (N_3218,N_536,N_722);
or U3219 (N_3219,N_658,N_186);
and U3220 (N_3220,N_369,N_663);
or U3221 (N_3221,N_1643,N_778);
nand U3222 (N_3222,N_1651,N_1149);
nor U3223 (N_3223,N_1899,N_1077);
xor U3224 (N_3224,N_1362,N_355);
or U3225 (N_3225,N_2273,N_899);
or U3226 (N_3226,N_282,N_1996);
xnor U3227 (N_3227,N_1063,N_939);
and U3228 (N_3228,N_2420,N_1024);
and U3229 (N_3229,N_2294,N_367);
or U3230 (N_3230,N_2348,N_2239);
nand U3231 (N_3231,N_2359,N_1122);
or U3232 (N_3232,N_1880,N_1542);
xnor U3233 (N_3233,N_2048,N_2002);
and U3234 (N_3234,N_1172,N_459);
nor U3235 (N_3235,N_876,N_496);
nand U3236 (N_3236,N_613,N_570);
nand U3237 (N_3237,N_10,N_2310);
nand U3238 (N_3238,N_1213,N_1603);
xor U3239 (N_3239,N_460,N_327);
nand U3240 (N_3240,N_764,N_2084);
and U3241 (N_3241,N_1006,N_2209);
xor U3242 (N_3242,N_742,N_1412);
nor U3243 (N_3243,N_1842,N_35);
or U3244 (N_3244,N_243,N_1463);
nor U3245 (N_3245,N_955,N_1814);
nor U3246 (N_3246,N_480,N_219);
or U3247 (N_3247,N_1387,N_432);
and U3248 (N_3248,N_1255,N_1652);
nand U3249 (N_3249,N_1319,N_1107);
nor U3250 (N_3250,N_2053,N_1139);
nor U3251 (N_3251,N_1607,N_757);
nand U3252 (N_3252,N_2300,N_872);
and U3253 (N_3253,N_1570,N_2186);
nand U3254 (N_3254,N_1067,N_821);
xor U3255 (N_3255,N_509,N_85);
or U3256 (N_3256,N_968,N_1576);
nor U3257 (N_3257,N_1337,N_1936);
or U3258 (N_3258,N_1372,N_719);
nor U3259 (N_3259,N_1620,N_628);
or U3260 (N_3260,N_70,N_1281);
nor U3261 (N_3261,N_1862,N_415);
xor U3262 (N_3262,N_920,N_1250);
nor U3263 (N_3263,N_2485,N_1910);
nor U3264 (N_3264,N_223,N_1906);
nor U3265 (N_3265,N_880,N_1923);
nand U3266 (N_3266,N_1457,N_502);
and U3267 (N_3267,N_1668,N_2023);
nor U3268 (N_3268,N_1874,N_606);
and U3269 (N_3269,N_2231,N_654);
nor U3270 (N_3270,N_1581,N_709);
or U3271 (N_3271,N_832,N_446);
nor U3272 (N_3272,N_923,N_1625);
xor U3273 (N_3273,N_1953,N_1699);
and U3274 (N_3274,N_1111,N_292);
nand U3275 (N_3275,N_1011,N_485);
xnor U3276 (N_3276,N_379,N_2444);
and U3277 (N_3277,N_770,N_2237);
nor U3278 (N_3278,N_78,N_123);
nor U3279 (N_3279,N_177,N_768);
nand U3280 (N_3280,N_1785,N_2425);
or U3281 (N_3281,N_1500,N_1903);
nand U3282 (N_3282,N_1623,N_137);
and U3283 (N_3283,N_823,N_1716);
nor U3284 (N_3284,N_2230,N_1051);
or U3285 (N_3285,N_2484,N_673);
or U3286 (N_3286,N_2403,N_1764);
and U3287 (N_3287,N_151,N_2499);
or U3288 (N_3288,N_1504,N_1790);
and U3289 (N_3289,N_230,N_2014);
nor U3290 (N_3290,N_835,N_1329);
or U3291 (N_3291,N_1784,N_879);
or U3292 (N_3292,N_1706,N_978);
nand U3293 (N_3293,N_252,N_1501);
xor U3294 (N_3294,N_902,N_2390);
nor U3295 (N_3295,N_1262,N_1889);
and U3296 (N_3296,N_1397,N_945);
and U3297 (N_3297,N_634,N_15);
nand U3298 (N_3298,N_2212,N_518);
or U3299 (N_3299,N_1991,N_2003);
xor U3300 (N_3300,N_2018,N_954);
xor U3301 (N_3301,N_258,N_237);
nor U3302 (N_3302,N_1511,N_1211);
or U3303 (N_3303,N_2127,N_1995);
or U3304 (N_3304,N_1130,N_580);
and U3305 (N_3305,N_60,N_1410);
nor U3306 (N_3306,N_146,N_1416);
nor U3307 (N_3307,N_587,N_356);
and U3308 (N_3308,N_1020,N_767);
nor U3309 (N_3309,N_826,N_2167);
or U3310 (N_3310,N_431,N_929);
nor U3311 (N_3311,N_198,N_8);
and U3312 (N_3312,N_594,N_1809);
nor U3313 (N_3313,N_1826,N_816);
nand U3314 (N_3314,N_956,N_1310);
nor U3315 (N_3315,N_565,N_753);
nor U3316 (N_3316,N_1676,N_117);
xor U3317 (N_3317,N_1771,N_2062);
and U3318 (N_3318,N_639,N_2286);
and U3319 (N_3319,N_1295,N_2185);
and U3320 (N_3320,N_1637,N_175);
and U3321 (N_3321,N_1847,N_1333);
or U3322 (N_3322,N_501,N_1147);
or U3323 (N_3323,N_700,N_1186);
and U3324 (N_3324,N_1765,N_475);
xnor U3325 (N_3325,N_1271,N_1535);
nand U3326 (N_3326,N_875,N_1189);
and U3327 (N_3327,N_1655,N_1426);
nand U3328 (N_3328,N_2402,N_1774);
nand U3329 (N_3329,N_784,N_1203);
and U3330 (N_3330,N_124,N_588);
or U3331 (N_3331,N_1345,N_1325);
or U3332 (N_3332,N_407,N_424);
and U3333 (N_3333,N_32,N_143);
and U3334 (N_3334,N_1315,N_86);
nor U3335 (N_3335,N_1274,N_1590);
and U3336 (N_3336,N_664,N_16);
nor U3337 (N_3337,N_1519,N_1258);
nand U3338 (N_3338,N_1038,N_2241);
or U3339 (N_3339,N_1148,N_29);
xor U3340 (N_3340,N_2034,N_61);
or U3341 (N_3341,N_2302,N_1206);
nand U3342 (N_3342,N_2303,N_2357);
and U3343 (N_3343,N_2371,N_2316);
or U3344 (N_3344,N_2355,N_1767);
or U3345 (N_3345,N_668,N_625);
xnor U3346 (N_3346,N_1381,N_997);
nand U3347 (N_3347,N_577,N_0);
and U3348 (N_3348,N_132,N_341);
xor U3349 (N_3349,N_1379,N_1245);
and U3350 (N_3350,N_410,N_1579);
or U3351 (N_3351,N_893,N_88);
or U3352 (N_3352,N_1865,N_2426);
nor U3353 (N_3353,N_1598,N_1551);
or U3354 (N_3354,N_414,N_1296);
and U3355 (N_3355,N_2085,N_1725);
xor U3356 (N_3356,N_1290,N_1962);
nor U3357 (N_3357,N_300,N_2318);
nand U3358 (N_3358,N_2153,N_982);
or U3359 (N_3359,N_2082,N_2493);
and U3360 (N_3360,N_2339,N_1222);
and U3361 (N_3361,N_1588,N_1132);
nor U3362 (N_3362,N_1975,N_1916);
and U3363 (N_3363,N_2387,N_26);
nor U3364 (N_3364,N_439,N_908);
nor U3365 (N_3365,N_1378,N_2058);
nor U3366 (N_3366,N_1552,N_883);
or U3367 (N_3367,N_2319,N_296);
nand U3368 (N_3368,N_2160,N_1968);
xnor U3369 (N_3369,N_1630,N_1249);
or U3370 (N_3370,N_1957,N_2214);
or U3371 (N_3371,N_1648,N_425);
and U3372 (N_3372,N_2275,N_2134);
and U3373 (N_3373,N_1667,N_457);
or U3374 (N_3374,N_2189,N_23);
and U3375 (N_3375,N_2491,N_1894);
nor U3376 (N_3376,N_720,N_2192);
nor U3377 (N_3377,N_2293,N_1307);
or U3378 (N_3378,N_2054,N_1048);
nand U3379 (N_3379,N_1838,N_2190);
or U3380 (N_3380,N_465,N_238);
xor U3381 (N_3381,N_2385,N_1022);
or U3382 (N_3382,N_213,N_1905);
nand U3383 (N_3383,N_486,N_1503);
and U3384 (N_3384,N_774,N_2399);
nand U3385 (N_3385,N_329,N_1755);
nand U3386 (N_3386,N_2106,N_758);
nand U3387 (N_3387,N_1545,N_445);
nand U3388 (N_3388,N_2388,N_1192);
nand U3389 (N_3389,N_643,N_1055);
nor U3390 (N_3390,N_1016,N_2324);
nand U3391 (N_3391,N_1157,N_2382);
nand U3392 (N_3392,N_232,N_815);
nor U3393 (N_3393,N_1656,N_1039);
and U3394 (N_3394,N_884,N_1270);
nand U3395 (N_3395,N_2410,N_1369);
and U3396 (N_3396,N_403,N_781);
or U3397 (N_3397,N_2492,N_2349);
xnor U3398 (N_3398,N_635,N_1467);
nor U3399 (N_3399,N_1713,N_1638);
or U3400 (N_3400,N_1622,N_972);
and U3401 (N_3401,N_411,N_187);
and U3402 (N_3402,N_1688,N_537);
or U3403 (N_3403,N_2463,N_730);
nor U3404 (N_3404,N_579,N_2047);
xnor U3405 (N_3405,N_1437,N_839);
nand U3406 (N_3406,N_771,N_368);
nand U3407 (N_3407,N_100,N_1618);
xnor U3408 (N_3408,N_2451,N_890);
nand U3409 (N_3409,N_1233,N_1069);
or U3410 (N_3410,N_1034,N_1251);
nor U3411 (N_3411,N_2015,N_851);
nand U3412 (N_3412,N_1684,N_2111);
or U3413 (N_3413,N_1316,N_1058);
and U3414 (N_3414,N_940,N_2187);
nand U3415 (N_3415,N_2069,N_9);
and U3416 (N_3416,N_1559,N_524);
nor U3417 (N_3417,N_157,N_2112);
and U3418 (N_3418,N_456,N_551);
and U3419 (N_3419,N_887,N_1123);
and U3420 (N_3420,N_2137,N_1230);
nor U3421 (N_3421,N_220,N_546);
or U3422 (N_3422,N_352,N_504);
nand U3423 (N_3423,N_2469,N_1681);
or U3424 (N_3424,N_1264,N_1066);
nor U3425 (N_3425,N_934,N_1529);
nor U3426 (N_3426,N_1710,N_2424);
and U3427 (N_3427,N_1041,N_523);
nand U3428 (N_3428,N_1450,N_984);
or U3429 (N_3429,N_293,N_359);
nand U3430 (N_3430,N_156,N_13);
nand U3431 (N_3431,N_1709,N_1464);
and U3432 (N_3432,N_1915,N_442);
and U3433 (N_3433,N_1678,N_692);
and U3434 (N_3434,N_1289,N_1524);
or U3435 (N_3435,N_98,N_2280);
and U3436 (N_3436,N_966,N_2101);
and U3437 (N_3437,N_574,N_944);
or U3438 (N_3438,N_335,N_517);
nand U3439 (N_3439,N_598,N_39);
nand U3440 (N_3440,N_629,N_388);
xnor U3441 (N_3441,N_1753,N_204);
or U3442 (N_3442,N_317,N_1640);
nor U3443 (N_3443,N_2141,N_1812);
or U3444 (N_3444,N_1691,N_1400);
xor U3445 (N_3445,N_963,N_2076);
xor U3446 (N_3446,N_1856,N_207);
nor U3447 (N_3447,N_2040,N_1854);
nand U3448 (N_3448,N_2234,N_552);
or U3449 (N_3449,N_510,N_371);
and U3450 (N_3450,N_1061,N_539);
nor U3451 (N_3451,N_1461,N_405);
nand U3452 (N_3452,N_846,N_1938);
nor U3453 (N_3453,N_234,N_1117);
nand U3454 (N_3454,N_817,N_2301);
nand U3455 (N_3455,N_28,N_1934);
nor U3456 (N_3456,N_946,N_2427);
or U3457 (N_3457,N_2070,N_154);
xnor U3458 (N_3458,N_309,N_47);
nand U3459 (N_3459,N_2278,N_2281);
nand U3460 (N_3460,N_320,N_1708);
nand U3461 (N_3461,N_1922,N_1001);
and U3462 (N_3462,N_1481,N_1557);
and U3463 (N_3463,N_334,N_144);
xnor U3464 (N_3464,N_2419,N_1436);
nand U3465 (N_3465,N_2368,N_1661);
nand U3466 (N_3466,N_183,N_1835);
nand U3467 (N_3467,N_3,N_107);
and U3468 (N_3468,N_2434,N_1649);
or U3469 (N_3469,N_1303,N_2418);
nor U3470 (N_3470,N_458,N_267);
nor U3471 (N_3471,N_1494,N_199);
nand U3472 (N_3472,N_1518,N_544);
and U3473 (N_3473,N_1939,N_2309);
nor U3474 (N_3474,N_2035,N_1861);
nor U3475 (N_3475,N_2200,N_1807);
nand U3476 (N_3476,N_1583,N_1877);
or U3477 (N_3477,N_1882,N_894);
nor U3478 (N_3478,N_375,N_776);
or U3479 (N_3479,N_1185,N_806);
nor U3480 (N_3480,N_1224,N_76);
and U3481 (N_3481,N_675,N_221);
nor U3482 (N_3482,N_1195,N_1817);
nor U3483 (N_3483,N_1878,N_607);
xor U3484 (N_3484,N_1152,N_1508);
and U3485 (N_3485,N_349,N_279);
nor U3486 (N_3486,N_2314,N_986);
and U3487 (N_3487,N_1210,N_95);
or U3488 (N_3488,N_1118,N_2490);
and U3489 (N_3489,N_1059,N_1073);
or U3490 (N_3490,N_19,N_2086);
and U3491 (N_3491,N_1534,N_688);
and U3492 (N_3492,N_1589,N_1600);
nand U3493 (N_3493,N_653,N_40);
and U3494 (N_3494,N_1028,N_995);
or U3495 (N_3495,N_900,N_2471);
nand U3496 (N_3496,N_167,N_2219);
nand U3497 (N_3497,N_698,N_357);
and U3498 (N_3498,N_1616,N_242);
xnor U3499 (N_3499,N_1896,N_1843);
and U3500 (N_3500,N_104,N_2335);
nor U3501 (N_3501,N_576,N_1342);
or U3502 (N_3502,N_857,N_1768);
nor U3503 (N_3503,N_1540,N_505);
nor U3504 (N_3504,N_1217,N_2312);
nand U3505 (N_3505,N_728,N_103);
xnor U3506 (N_3506,N_992,N_1382);
nor U3507 (N_3507,N_521,N_2299);
xor U3508 (N_3508,N_512,N_896);
nor U3509 (N_3509,N_1846,N_1091);
nor U3510 (N_3510,N_90,N_1730);
xor U3511 (N_3511,N_270,N_813);
nor U3512 (N_3512,N_2142,N_214);
or U3513 (N_3513,N_706,N_1447);
nor U3514 (N_3514,N_1187,N_1049);
and U3515 (N_3515,N_965,N_493);
nor U3516 (N_3516,N_2238,N_324);
nand U3517 (N_3517,N_1911,N_1322);
nor U3518 (N_3518,N_1403,N_1413);
nor U3519 (N_3519,N_1585,N_2092);
and U3520 (N_3520,N_268,N_862);
xor U3521 (N_3521,N_2417,N_1606);
nand U3522 (N_3522,N_1657,N_1578);
or U3523 (N_3523,N_1395,N_1818);
or U3524 (N_3524,N_592,N_364);
and U3525 (N_3525,N_1293,N_227);
and U3526 (N_3526,N_2372,N_1455);
and U3527 (N_3527,N_2378,N_526);
and U3528 (N_3528,N_2497,N_1913);
and U3529 (N_3529,N_834,N_614);
or U3530 (N_3530,N_828,N_63);
nor U3531 (N_3531,N_2477,N_1009);
nand U3532 (N_3532,N_205,N_655);
nand U3533 (N_3533,N_1366,N_1168);
or U3534 (N_3534,N_1360,N_1275);
nor U3535 (N_3535,N_1924,N_1918);
nor U3536 (N_3536,N_788,N_996);
and U3537 (N_3537,N_429,N_1021);
and U3538 (N_3538,N_638,N_1458);
or U3539 (N_3539,N_674,N_139);
nor U3540 (N_3540,N_25,N_1958);
or U3541 (N_3541,N_1943,N_169);
or U3542 (N_3542,N_1375,N_449);
nor U3543 (N_3543,N_37,N_2118);
nor U3544 (N_3544,N_677,N_255);
and U3545 (N_3545,N_1528,N_1201);
and U3546 (N_3546,N_346,N_1468);
nor U3547 (N_3547,N_1092,N_381);
nand U3548 (N_3548,N_484,N_111);
nand U3549 (N_3549,N_843,N_1305);
nand U3550 (N_3550,N_225,N_1525);
or U3551 (N_3551,N_1658,N_2026);
and U3552 (N_3552,N_1159,N_1370);
nand U3553 (N_3553,N_2414,N_1810);
nor U3554 (N_3554,N_871,N_33);
or U3555 (N_3555,N_2017,N_1170);
and U3556 (N_3556,N_1663,N_2242);
or U3557 (N_3557,N_695,N_1937);
and U3558 (N_3558,N_2397,N_751);
and U3559 (N_3559,N_1234,N_1093);
and U3560 (N_3560,N_1538,N_1759);
xor U3561 (N_3561,N_2333,N_2352);
nor U3562 (N_3562,N_416,N_715);
xnor U3563 (N_3563,N_2216,N_1744);
nand U3564 (N_3564,N_693,N_2130);
nor U3565 (N_3565,N_657,N_1714);
or U3566 (N_3566,N_805,N_752);
nand U3567 (N_3567,N_1166,N_2030);
or U3568 (N_3568,N_211,N_2163);
or U3569 (N_3569,N_2021,N_2036);
nand U3570 (N_3570,N_1373,N_1100);
nand U3571 (N_3571,N_734,N_1553);
and U3572 (N_3572,N_1377,N_354);
nand U3573 (N_3573,N_1106,N_1418);
or U3574 (N_3574,N_616,N_795);
and U3575 (N_3575,N_1221,N_676);
or U3576 (N_3576,N_1032,N_2114);
or U3577 (N_3577,N_1900,N_1037);
nand U3578 (N_3578,N_921,N_147);
nor U3579 (N_3579,N_1601,N_1099);
or U3580 (N_3580,N_2100,N_2261);
nor U3581 (N_3581,N_2129,N_2213);
xor U3582 (N_3582,N_1955,N_916);
and U3583 (N_3583,N_1459,N_1427);
nor U3584 (N_3584,N_1780,N_264);
nand U3585 (N_3585,N_2283,N_158);
nand U3586 (N_3586,N_224,N_873);
nor U3587 (N_3587,N_1407,N_659);
nand U3588 (N_3588,N_863,N_1954);
xnor U3589 (N_3589,N_840,N_2438);
nand U3590 (N_3590,N_304,N_48);
nor U3591 (N_3591,N_142,N_2379);
nor U3592 (N_3592,N_112,N_342);
nor U3593 (N_3593,N_1204,N_947);
and U3594 (N_3594,N_2164,N_2454);
nor U3595 (N_3595,N_2139,N_1424);
and U3596 (N_3596,N_1496,N_741);
nor U3597 (N_3597,N_72,N_1268);
nor U3598 (N_3598,N_756,N_2377);
xor U3599 (N_3599,N_1181,N_2119);
and U3600 (N_3600,N_464,N_1193);
nor U3601 (N_3601,N_2346,N_2);
xnor U3602 (N_3602,N_1567,N_2338);
and U3603 (N_3603,N_2391,N_2165);
or U3604 (N_3604,N_51,N_683);
and U3605 (N_3605,N_563,N_2258);
nor U3606 (N_3606,N_1769,N_1448);
nand U3607 (N_3607,N_2211,N_2140);
nand U3608 (N_3608,N_2483,N_497);
xnor U3609 (N_3609,N_477,N_1801);
nor U3610 (N_3610,N_2039,N_1844);
and U3611 (N_3611,N_1155,N_1978);
nor U3612 (N_3612,N_864,N_1223);
and U3613 (N_3613,N_421,N_1612);
nor U3614 (N_3614,N_1156,N_2171);
nor U3615 (N_3615,N_1163,N_1014);
nand U3616 (N_3616,N_2225,N_845);
or U3617 (N_3617,N_1353,N_1779);
nor U3618 (N_3618,N_2228,N_1116);
nand U3619 (N_3619,N_543,N_798);
nand U3620 (N_3620,N_721,N_2287);
xnor U3621 (N_3621,N_1417,N_1895);
or U3622 (N_3622,N_1605,N_2494);
or U3623 (N_3623,N_2375,N_765);
xnor U3624 (N_3624,N_2447,N_1207);
or U3625 (N_3625,N_1246,N_849);
nor U3626 (N_3626,N_1466,N_608);
nor U3627 (N_3627,N_684,N_1298);
and U3628 (N_3628,N_89,N_478);
nor U3629 (N_3629,N_1948,N_2330);
nor U3630 (N_3630,N_263,N_881);
nor U3631 (N_3631,N_747,N_708);
nand U3632 (N_3632,N_2240,N_2455);
nand U3633 (N_3633,N_1076,N_2279);
and U3634 (N_3634,N_1399,N_2422);
and U3635 (N_3635,N_1351,N_2175);
and U3636 (N_3636,N_2353,N_1292);
xnor U3637 (N_3637,N_1374,N_2087);
and U3638 (N_3638,N_601,N_1912);
nand U3639 (N_3639,N_333,N_789);
nand U3640 (N_3640,N_209,N_2006);
nand U3641 (N_3641,N_2430,N_886);
and U3642 (N_3642,N_374,N_1420);
nand U3643 (N_3643,N_1702,N_1280);
nand U3644 (N_3644,N_836,N_297);
nor U3645 (N_3645,N_1513,N_1976);
xnor U3646 (N_3646,N_2470,N_73);
and U3647 (N_3647,N_394,N_928);
nand U3648 (N_3648,N_2206,N_957);
nand U3649 (N_3649,N_556,N_1226);
or U3650 (N_3650,N_121,N_2155);
or U3651 (N_3651,N_1314,N_56);
or U3652 (N_3652,N_395,N_1386);
nor U3653 (N_3653,N_1960,N_447);
or U3654 (N_3654,N_240,N_434);
nand U3655 (N_3655,N_1673,N_617);
nand U3656 (N_3656,N_2096,N_717);
nor U3657 (N_3657,N_1701,N_347);
or U3658 (N_3658,N_1294,N_1438);
nand U3659 (N_3659,N_1252,N_866);
nand U3660 (N_3660,N_2431,N_1541);
and U3661 (N_3661,N_1,N_1932);
and U3662 (N_3662,N_2321,N_2205);
or U3663 (N_3663,N_1531,N_2489);
nand U3664 (N_3664,N_818,N_260);
nor U3665 (N_3665,N_2423,N_2042);
nor U3666 (N_3666,N_1114,N_378);
or U3667 (N_3667,N_2044,N_1719);
xnor U3668 (N_3668,N_959,N_246);
nand U3669 (N_3669,N_1886,N_830);
xor U3670 (N_3670,N_1963,N_108);
nor U3671 (N_3671,N_1998,N_190);
or U3672 (N_3672,N_71,N_914);
nand U3673 (N_3673,N_773,N_761);
or U3674 (N_3674,N_2384,N_680);
nor U3675 (N_3675,N_1081,N_602);
nor U3676 (N_3676,N_1208,N_31);
and U3677 (N_3677,N_1070,N_860);
nand U3678 (N_3678,N_666,N_1604);
nand U3679 (N_3679,N_256,N_2172);
or U3680 (N_3680,N_1745,N_1505);
or U3681 (N_3681,N_96,N_216);
nand U3682 (N_3682,N_1110,N_1442);
nor U3683 (N_3683,N_1175,N_906);
or U3684 (N_3684,N_1158,N_624);
nor U3685 (N_3685,N_1029,N_11);
xnor U3686 (N_3686,N_1371,N_179);
and U3687 (N_3687,N_2315,N_1445);
nor U3688 (N_3688,N_489,N_201);
or U3689 (N_3689,N_1140,N_1773);
and U3690 (N_3690,N_1031,N_215);
xnor U3691 (N_3691,N_1741,N_160);
xor U3692 (N_3692,N_440,N_1253);
or U3693 (N_3693,N_1859,N_1358);
nand U3694 (N_3694,N_1721,N_1762);
nand U3695 (N_3695,N_1019,N_1075);
and U3696 (N_3696,N_1060,N_2196);
nor U3697 (N_3697,N_1795,N_531);
nor U3698 (N_3698,N_1165,N_1340);
or U3699 (N_3699,N_2157,N_572);
nor U3700 (N_3700,N_2327,N_2354);
nor U3701 (N_3701,N_1543,N_951);
and U3702 (N_3702,N_113,N_733);
and U3703 (N_3703,N_441,N_831);
nor U3704 (N_3704,N_1830,N_2468);
nor U3705 (N_3705,N_2195,N_44);
nand U3706 (N_3706,N_1639,N_1288);
xnor U3707 (N_3707,N_1429,N_585);
xor U3708 (N_3708,N_1495,N_2376);
nor U3709 (N_3709,N_1507,N_277);
or U3710 (N_3710,N_2392,N_1005);
or U3711 (N_3711,N_1054,N_2105);
nor U3712 (N_3712,N_1335,N_1728);
nor U3713 (N_3713,N_797,N_1992);
xnor U3714 (N_3714,N_1703,N_787);
nand U3715 (N_3715,N_406,N_1527);
and U3716 (N_3716,N_804,N_1327);
nand U3717 (N_3717,N_330,N_312);
nand U3718 (N_3718,N_848,N_522);
nor U3719 (N_3719,N_418,N_605);
and U3720 (N_3720,N_2473,N_987);
xnor U3721 (N_3721,N_1134,N_1901);
nor U3722 (N_3722,N_852,N_1633);
nor U3723 (N_3723,N_1712,N_358);
nor U3724 (N_3724,N_736,N_382);
or U3725 (N_3725,N_1554,N_114);
and U3726 (N_3726,N_1409,N_1257);
xnor U3727 (N_3727,N_1025,N_1286);
and U3728 (N_3728,N_1736,N_1183);
nand U3729 (N_3729,N_319,N_257);
or U3730 (N_3730,N_191,N_726);
or U3731 (N_3731,N_1469,N_1119);
xnor U3732 (N_3732,N_93,N_701);
or U3733 (N_3733,N_1526,N_2429);
nor U3734 (N_3734,N_1182,N_748);
or U3735 (N_3735,N_856,N_1828);
nand U3736 (N_3736,N_600,N_1718);
and U3737 (N_3737,N_1521,N_553);
nand U3738 (N_3738,N_1212,N_52);
xor U3739 (N_3739,N_1334,N_1654);
and U3740 (N_3740,N_1993,N_500);
xnor U3741 (N_3741,N_780,N_759);
nand U3742 (N_3742,N_53,N_1239);
nand U3743 (N_3743,N_732,N_2059);
nor U3744 (N_3744,N_667,N_1904);
nand U3745 (N_3745,N_646,N_2311);
nand U3746 (N_3746,N_1914,N_372);
or U3747 (N_3747,N_739,N_474);
or U3748 (N_3748,N_1174,N_2313);
or U3749 (N_3749,N_1898,N_1740);
and U3750 (N_3750,N_1864,N_2419);
and U3751 (N_3751,N_1909,N_536);
nor U3752 (N_3752,N_237,N_1845);
and U3753 (N_3753,N_945,N_1012);
nand U3754 (N_3754,N_1690,N_383);
nand U3755 (N_3755,N_1266,N_2179);
nand U3756 (N_3756,N_2446,N_2404);
and U3757 (N_3757,N_2084,N_252);
or U3758 (N_3758,N_103,N_2492);
or U3759 (N_3759,N_139,N_1878);
xor U3760 (N_3760,N_1642,N_2106);
nor U3761 (N_3761,N_850,N_1445);
and U3762 (N_3762,N_595,N_1595);
or U3763 (N_3763,N_1792,N_825);
and U3764 (N_3764,N_2369,N_96);
nor U3765 (N_3765,N_1707,N_675);
or U3766 (N_3766,N_1331,N_752);
or U3767 (N_3767,N_606,N_2095);
nor U3768 (N_3768,N_216,N_202);
xor U3769 (N_3769,N_1626,N_382);
and U3770 (N_3770,N_2307,N_1323);
and U3771 (N_3771,N_1843,N_1197);
nand U3772 (N_3772,N_1890,N_908);
and U3773 (N_3773,N_234,N_663);
and U3774 (N_3774,N_2344,N_1521);
and U3775 (N_3775,N_221,N_2008);
or U3776 (N_3776,N_1951,N_1771);
or U3777 (N_3777,N_2347,N_1956);
xnor U3778 (N_3778,N_1281,N_2365);
and U3779 (N_3779,N_1911,N_895);
nand U3780 (N_3780,N_2069,N_1237);
xnor U3781 (N_3781,N_1069,N_1920);
and U3782 (N_3782,N_2195,N_1788);
xnor U3783 (N_3783,N_1762,N_1380);
xor U3784 (N_3784,N_719,N_1494);
or U3785 (N_3785,N_326,N_2249);
and U3786 (N_3786,N_1827,N_1989);
nand U3787 (N_3787,N_2260,N_2036);
nand U3788 (N_3788,N_1207,N_2119);
nor U3789 (N_3789,N_481,N_1189);
nand U3790 (N_3790,N_750,N_788);
and U3791 (N_3791,N_1205,N_2436);
or U3792 (N_3792,N_572,N_1106);
and U3793 (N_3793,N_2190,N_655);
nor U3794 (N_3794,N_1790,N_1320);
and U3795 (N_3795,N_1514,N_2204);
xor U3796 (N_3796,N_1906,N_1421);
nand U3797 (N_3797,N_2164,N_721);
nor U3798 (N_3798,N_1897,N_675);
and U3799 (N_3799,N_1934,N_2188);
and U3800 (N_3800,N_8,N_589);
nand U3801 (N_3801,N_59,N_21);
nor U3802 (N_3802,N_483,N_1278);
nand U3803 (N_3803,N_1171,N_2172);
nor U3804 (N_3804,N_1029,N_130);
or U3805 (N_3805,N_2203,N_820);
nor U3806 (N_3806,N_1235,N_1739);
xor U3807 (N_3807,N_2289,N_2125);
and U3808 (N_3808,N_2263,N_1828);
nand U3809 (N_3809,N_22,N_1946);
nand U3810 (N_3810,N_641,N_115);
nor U3811 (N_3811,N_2277,N_2136);
nand U3812 (N_3812,N_2051,N_1620);
nor U3813 (N_3813,N_1335,N_13);
or U3814 (N_3814,N_1219,N_1886);
xor U3815 (N_3815,N_1811,N_1857);
nand U3816 (N_3816,N_891,N_1338);
nor U3817 (N_3817,N_1192,N_495);
and U3818 (N_3818,N_371,N_136);
or U3819 (N_3819,N_2132,N_990);
and U3820 (N_3820,N_1809,N_811);
or U3821 (N_3821,N_2319,N_1373);
nand U3822 (N_3822,N_1865,N_1597);
nand U3823 (N_3823,N_1228,N_113);
nor U3824 (N_3824,N_1055,N_229);
nor U3825 (N_3825,N_2176,N_1493);
nor U3826 (N_3826,N_495,N_1053);
and U3827 (N_3827,N_663,N_1925);
nand U3828 (N_3828,N_1377,N_1391);
xnor U3829 (N_3829,N_250,N_178);
nand U3830 (N_3830,N_2469,N_148);
and U3831 (N_3831,N_230,N_1910);
nor U3832 (N_3832,N_2100,N_129);
or U3833 (N_3833,N_954,N_1254);
xor U3834 (N_3834,N_918,N_2184);
nand U3835 (N_3835,N_494,N_1210);
or U3836 (N_3836,N_766,N_1119);
and U3837 (N_3837,N_2449,N_356);
and U3838 (N_3838,N_967,N_344);
or U3839 (N_3839,N_1096,N_1856);
xnor U3840 (N_3840,N_1447,N_1874);
nand U3841 (N_3841,N_31,N_889);
and U3842 (N_3842,N_2185,N_1454);
and U3843 (N_3843,N_257,N_2271);
or U3844 (N_3844,N_848,N_750);
nor U3845 (N_3845,N_842,N_2238);
and U3846 (N_3846,N_2139,N_123);
nor U3847 (N_3847,N_67,N_2373);
nand U3848 (N_3848,N_1708,N_2399);
nand U3849 (N_3849,N_1427,N_419);
nand U3850 (N_3850,N_1682,N_299);
xnor U3851 (N_3851,N_91,N_147);
and U3852 (N_3852,N_569,N_1753);
and U3853 (N_3853,N_1627,N_771);
xor U3854 (N_3854,N_1137,N_2427);
nand U3855 (N_3855,N_848,N_137);
and U3856 (N_3856,N_424,N_2448);
nand U3857 (N_3857,N_945,N_1857);
nand U3858 (N_3858,N_837,N_2326);
and U3859 (N_3859,N_1375,N_820);
nand U3860 (N_3860,N_579,N_2064);
nor U3861 (N_3861,N_1304,N_223);
nor U3862 (N_3862,N_1882,N_592);
or U3863 (N_3863,N_2271,N_686);
or U3864 (N_3864,N_2230,N_1116);
nor U3865 (N_3865,N_2488,N_1439);
and U3866 (N_3866,N_479,N_1111);
nand U3867 (N_3867,N_1539,N_1055);
or U3868 (N_3868,N_2015,N_45);
and U3869 (N_3869,N_541,N_134);
or U3870 (N_3870,N_1994,N_2467);
nand U3871 (N_3871,N_280,N_2118);
or U3872 (N_3872,N_1900,N_1517);
and U3873 (N_3873,N_1258,N_591);
nor U3874 (N_3874,N_91,N_1996);
nor U3875 (N_3875,N_1974,N_331);
and U3876 (N_3876,N_1210,N_1287);
nand U3877 (N_3877,N_1018,N_879);
and U3878 (N_3878,N_940,N_593);
or U3879 (N_3879,N_237,N_523);
nand U3880 (N_3880,N_1905,N_2249);
nand U3881 (N_3881,N_2419,N_727);
nand U3882 (N_3882,N_477,N_876);
nand U3883 (N_3883,N_1868,N_1643);
and U3884 (N_3884,N_1390,N_1739);
and U3885 (N_3885,N_1185,N_944);
and U3886 (N_3886,N_47,N_1024);
nand U3887 (N_3887,N_403,N_1191);
and U3888 (N_3888,N_864,N_1305);
nor U3889 (N_3889,N_756,N_1297);
xor U3890 (N_3890,N_2424,N_824);
nand U3891 (N_3891,N_784,N_751);
and U3892 (N_3892,N_2395,N_493);
nand U3893 (N_3893,N_2087,N_312);
nand U3894 (N_3894,N_2256,N_1050);
nor U3895 (N_3895,N_229,N_2464);
nor U3896 (N_3896,N_2263,N_668);
nand U3897 (N_3897,N_1105,N_2009);
nand U3898 (N_3898,N_1049,N_1794);
xnor U3899 (N_3899,N_123,N_1649);
nor U3900 (N_3900,N_1123,N_762);
nand U3901 (N_3901,N_1944,N_189);
nand U3902 (N_3902,N_746,N_40);
nand U3903 (N_3903,N_770,N_706);
and U3904 (N_3904,N_2253,N_1635);
xnor U3905 (N_3905,N_2199,N_603);
nor U3906 (N_3906,N_19,N_2048);
nand U3907 (N_3907,N_1549,N_929);
nand U3908 (N_3908,N_668,N_2144);
nand U3909 (N_3909,N_1092,N_619);
or U3910 (N_3910,N_1738,N_971);
xnor U3911 (N_3911,N_1881,N_641);
or U3912 (N_3912,N_862,N_915);
and U3913 (N_3913,N_2466,N_337);
and U3914 (N_3914,N_154,N_857);
nand U3915 (N_3915,N_347,N_1785);
nand U3916 (N_3916,N_1074,N_233);
nor U3917 (N_3917,N_2100,N_183);
and U3918 (N_3918,N_881,N_1629);
or U3919 (N_3919,N_2044,N_531);
nor U3920 (N_3920,N_710,N_545);
xnor U3921 (N_3921,N_2346,N_1237);
and U3922 (N_3922,N_1508,N_1306);
xnor U3923 (N_3923,N_358,N_264);
nor U3924 (N_3924,N_1684,N_1078);
or U3925 (N_3925,N_1456,N_177);
and U3926 (N_3926,N_2396,N_686);
or U3927 (N_3927,N_622,N_1661);
nand U3928 (N_3928,N_1015,N_1439);
nor U3929 (N_3929,N_1254,N_805);
or U3930 (N_3930,N_1826,N_1188);
and U3931 (N_3931,N_2141,N_868);
or U3932 (N_3932,N_281,N_2000);
xnor U3933 (N_3933,N_2152,N_1410);
nand U3934 (N_3934,N_1978,N_1068);
or U3935 (N_3935,N_624,N_781);
xor U3936 (N_3936,N_1060,N_603);
xnor U3937 (N_3937,N_838,N_1937);
or U3938 (N_3938,N_1714,N_2053);
and U3939 (N_3939,N_466,N_2281);
or U3940 (N_3940,N_2288,N_2024);
nor U3941 (N_3941,N_1077,N_132);
and U3942 (N_3942,N_788,N_1766);
nor U3943 (N_3943,N_212,N_1705);
and U3944 (N_3944,N_1531,N_597);
and U3945 (N_3945,N_2496,N_1532);
nand U3946 (N_3946,N_1470,N_33);
and U3947 (N_3947,N_1288,N_1955);
nor U3948 (N_3948,N_1242,N_382);
xor U3949 (N_3949,N_2123,N_1187);
nand U3950 (N_3950,N_73,N_2240);
and U3951 (N_3951,N_2016,N_169);
and U3952 (N_3952,N_7,N_700);
nand U3953 (N_3953,N_1815,N_1834);
xor U3954 (N_3954,N_2458,N_1078);
nor U3955 (N_3955,N_1177,N_281);
or U3956 (N_3956,N_2012,N_1809);
xor U3957 (N_3957,N_510,N_356);
nor U3958 (N_3958,N_2393,N_1827);
or U3959 (N_3959,N_897,N_1089);
and U3960 (N_3960,N_217,N_511);
xnor U3961 (N_3961,N_1367,N_282);
and U3962 (N_3962,N_2157,N_2056);
and U3963 (N_3963,N_498,N_1010);
and U3964 (N_3964,N_912,N_1822);
or U3965 (N_3965,N_136,N_997);
or U3966 (N_3966,N_611,N_949);
and U3967 (N_3967,N_814,N_746);
nand U3968 (N_3968,N_1289,N_1400);
or U3969 (N_3969,N_2199,N_1500);
and U3970 (N_3970,N_1749,N_330);
nand U3971 (N_3971,N_2053,N_1675);
xnor U3972 (N_3972,N_1101,N_2381);
and U3973 (N_3973,N_387,N_1063);
nand U3974 (N_3974,N_327,N_832);
and U3975 (N_3975,N_1227,N_1985);
nand U3976 (N_3976,N_2149,N_1072);
nor U3977 (N_3977,N_1009,N_1210);
nand U3978 (N_3978,N_2442,N_2445);
or U3979 (N_3979,N_1872,N_700);
nand U3980 (N_3980,N_731,N_1492);
nor U3981 (N_3981,N_1918,N_1935);
or U3982 (N_3982,N_1171,N_687);
nor U3983 (N_3983,N_44,N_1515);
nand U3984 (N_3984,N_581,N_1231);
or U3985 (N_3985,N_393,N_1391);
xor U3986 (N_3986,N_1279,N_2047);
or U3987 (N_3987,N_1784,N_2337);
xor U3988 (N_3988,N_2185,N_2270);
xor U3989 (N_3989,N_1084,N_2107);
nand U3990 (N_3990,N_1298,N_180);
or U3991 (N_3991,N_1575,N_341);
nand U3992 (N_3992,N_632,N_2191);
nand U3993 (N_3993,N_460,N_1736);
nand U3994 (N_3994,N_98,N_195);
nor U3995 (N_3995,N_238,N_2468);
and U3996 (N_3996,N_1559,N_1080);
nor U3997 (N_3997,N_1448,N_1532);
and U3998 (N_3998,N_1427,N_2119);
nor U3999 (N_3999,N_1215,N_45);
or U4000 (N_4000,N_2322,N_752);
xor U4001 (N_4001,N_645,N_2366);
and U4002 (N_4002,N_2220,N_455);
and U4003 (N_4003,N_1448,N_1720);
nor U4004 (N_4004,N_1642,N_1054);
xnor U4005 (N_4005,N_2154,N_1819);
nand U4006 (N_4006,N_943,N_497);
and U4007 (N_4007,N_1957,N_2237);
nor U4008 (N_4008,N_866,N_1106);
or U4009 (N_4009,N_1651,N_2492);
and U4010 (N_4010,N_2285,N_1339);
or U4011 (N_4011,N_789,N_322);
nor U4012 (N_4012,N_956,N_1848);
and U4013 (N_4013,N_2109,N_553);
nand U4014 (N_4014,N_360,N_736);
or U4015 (N_4015,N_1709,N_53);
nor U4016 (N_4016,N_2009,N_1228);
xnor U4017 (N_4017,N_1325,N_2215);
or U4018 (N_4018,N_1366,N_1979);
and U4019 (N_4019,N_485,N_635);
nand U4020 (N_4020,N_956,N_1625);
or U4021 (N_4021,N_535,N_1842);
or U4022 (N_4022,N_41,N_1078);
and U4023 (N_4023,N_55,N_2286);
nand U4024 (N_4024,N_1949,N_1075);
nand U4025 (N_4025,N_1825,N_12);
or U4026 (N_4026,N_965,N_423);
nor U4027 (N_4027,N_2309,N_728);
or U4028 (N_4028,N_1537,N_1686);
or U4029 (N_4029,N_2241,N_1694);
xor U4030 (N_4030,N_970,N_2291);
or U4031 (N_4031,N_158,N_2360);
nand U4032 (N_4032,N_2191,N_334);
nor U4033 (N_4033,N_2232,N_202);
and U4034 (N_4034,N_1627,N_1899);
nand U4035 (N_4035,N_2447,N_607);
nand U4036 (N_4036,N_978,N_1896);
nand U4037 (N_4037,N_1580,N_202);
and U4038 (N_4038,N_367,N_1674);
xor U4039 (N_4039,N_134,N_607);
nor U4040 (N_4040,N_78,N_778);
or U4041 (N_4041,N_1313,N_1373);
and U4042 (N_4042,N_795,N_1632);
nand U4043 (N_4043,N_1381,N_570);
xor U4044 (N_4044,N_2008,N_1936);
or U4045 (N_4045,N_2072,N_2359);
and U4046 (N_4046,N_478,N_104);
nand U4047 (N_4047,N_1268,N_1852);
and U4048 (N_4048,N_2498,N_2373);
nor U4049 (N_4049,N_1606,N_1348);
nor U4050 (N_4050,N_1654,N_16);
nor U4051 (N_4051,N_2085,N_1139);
or U4052 (N_4052,N_1984,N_868);
or U4053 (N_4053,N_1709,N_1558);
nor U4054 (N_4054,N_1895,N_307);
nor U4055 (N_4055,N_1255,N_1788);
or U4056 (N_4056,N_1250,N_1174);
or U4057 (N_4057,N_1218,N_2461);
nor U4058 (N_4058,N_1182,N_802);
nand U4059 (N_4059,N_250,N_1598);
nor U4060 (N_4060,N_47,N_162);
or U4061 (N_4061,N_1511,N_2232);
nand U4062 (N_4062,N_372,N_613);
and U4063 (N_4063,N_448,N_256);
and U4064 (N_4064,N_122,N_2462);
nor U4065 (N_4065,N_1513,N_1244);
or U4066 (N_4066,N_2464,N_1701);
nand U4067 (N_4067,N_1625,N_750);
or U4068 (N_4068,N_1988,N_1235);
and U4069 (N_4069,N_1774,N_966);
nand U4070 (N_4070,N_2258,N_1052);
or U4071 (N_4071,N_1651,N_492);
nand U4072 (N_4072,N_1737,N_1546);
or U4073 (N_4073,N_2494,N_56);
nor U4074 (N_4074,N_1154,N_994);
nor U4075 (N_4075,N_335,N_710);
or U4076 (N_4076,N_228,N_2416);
xor U4077 (N_4077,N_114,N_1722);
nor U4078 (N_4078,N_1501,N_2059);
nand U4079 (N_4079,N_367,N_2389);
nor U4080 (N_4080,N_1460,N_2265);
nand U4081 (N_4081,N_1730,N_2072);
nor U4082 (N_4082,N_1107,N_2124);
or U4083 (N_4083,N_727,N_262);
nor U4084 (N_4084,N_2418,N_378);
and U4085 (N_4085,N_913,N_227);
nor U4086 (N_4086,N_1702,N_1198);
nand U4087 (N_4087,N_1490,N_2294);
nor U4088 (N_4088,N_2330,N_672);
nand U4089 (N_4089,N_508,N_554);
nand U4090 (N_4090,N_190,N_1218);
and U4091 (N_4091,N_671,N_1099);
xnor U4092 (N_4092,N_625,N_293);
or U4093 (N_4093,N_2016,N_619);
xnor U4094 (N_4094,N_2257,N_1600);
and U4095 (N_4095,N_1135,N_1395);
nor U4096 (N_4096,N_590,N_258);
nand U4097 (N_4097,N_612,N_933);
or U4098 (N_4098,N_168,N_529);
or U4099 (N_4099,N_2406,N_170);
nand U4100 (N_4100,N_1598,N_736);
nand U4101 (N_4101,N_1333,N_225);
xnor U4102 (N_4102,N_847,N_709);
and U4103 (N_4103,N_832,N_2380);
nand U4104 (N_4104,N_268,N_2370);
nor U4105 (N_4105,N_545,N_2271);
nor U4106 (N_4106,N_2019,N_285);
and U4107 (N_4107,N_1331,N_110);
nor U4108 (N_4108,N_310,N_1855);
nand U4109 (N_4109,N_2357,N_1342);
and U4110 (N_4110,N_1578,N_2294);
nand U4111 (N_4111,N_1497,N_609);
and U4112 (N_4112,N_2107,N_844);
and U4113 (N_4113,N_615,N_249);
nor U4114 (N_4114,N_529,N_108);
nor U4115 (N_4115,N_994,N_2418);
nor U4116 (N_4116,N_2275,N_537);
or U4117 (N_4117,N_211,N_1619);
or U4118 (N_4118,N_74,N_1424);
nand U4119 (N_4119,N_1201,N_575);
or U4120 (N_4120,N_1253,N_2029);
nor U4121 (N_4121,N_1843,N_1007);
nand U4122 (N_4122,N_1566,N_1928);
and U4123 (N_4123,N_1704,N_330);
and U4124 (N_4124,N_1100,N_2031);
xnor U4125 (N_4125,N_594,N_212);
and U4126 (N_4126,N_2249,N_1680);
xor U4127 (N_4127,N_339,N_1206);
nor U4128 (N_4128,N_2198,N_2269);
and U4129 (N_4129,N_141,N_425);
or U4130 (N_4130,N_1690,N_1231);
xor U4131 (N_4131,N_1675,N_1420);
and U4132 (N_4132,N_803,N_339);
or U4133 (N_4133,N_2107,N_183);
nor U4134 (N_4134,N_465,N_782);
and U4135 (N_4135,N_1823,N_1673);
nor U4136 (N_4136,N_2363,N_758);
nor U4137 (N_4137,N_685,N_1880);
nand U4138 (N_4138,N_2129,N_2292);
and U4139 (N_4139,N_1269,N_2392);
and U4140 (N_4140,N_1490,N_501);
xor U4141 (N_4141,N_964,N_1260);
or U4142 (N_4142,N_2376,N_1973);
or U4143 (N_4143,N_2497,N_1697);
or U4144 (N_4144,N_1656,N_2089);
nand U4145 (N_4145,N_139,N_1318);
nor U4146 (N_4146,N_235,N_1150);
nand U4147 (N_4147,N_251,N_84);
nor U4148 (N_4148,N_1067,N_1076);
and U4149 (N_4149,N_833,N_2455);
and U4150 (N_4150,N_1067,N_1964);
nand U4151 (N_4151,N_26,N_2303);
or U4152 (N_4152,N_444,N_1608);
and U4153 (N_4153,N_1836,N_2193);
nand U4154 (N_4154,N_1922,N_617);
or U4155 (N_4155,N_1189,N_880);
and U4156 (N_4156,N_1896,N_1212);
and U4157 (N_4157,N_242,N_1298);
nor U4158 (N_4158,N_2431,N_401);
nor U4159 (N_4159,N_537,N_1028);
nand U4160 (N_4160,N_2368,N_1199);
and U4161 (N_4161,N_2059,N_1560);
nand U4162 (N_4162,N_1169,N_1967);
or U4163 (N_4163,N_2155,N_22);
xor U4164 (N_4164,N_907,N_375);
nor U4165 (N_4165,N_1671,N_1206);
nor U4166 (N_4166,N_1061,N_2083);
nand U4167 (N_4167,N_2332,N_2215);
and U4168 (N_4168,N_1642,N_851);
nand U4169 (N_4169,N_1427,N_1939);
nand U4170 (N_4170,N_2447,N_843);
or U4171 (N_4171,N_330,N_702);
nand U4172 (N_4172,N_1608,N_640);
nand U4173 (N_4173,N_2215,N_790);
nor U4174 (N_4174,N_30,N_623);
nand U4175 (N_4175,N_1553,N_1339);
nor U4176 (N_4176,N_1156,N_278);
and U4177 (N_4177,N_1046,N_1278);
or U4178 (N_4178,N_1515,N_1928);
xor U4179 (N_4179,N_1814,N_2367);
nand U4180 (N_4180,N_1813,N_2318);
and U4181 (N_4181,N_2343,N_2026);
nand U4182 (N_4182,N_1332,N_2011);
nor U4183 (N_4183,N_735,N_2409);
nor U4184 (N_4184,N_2245,N_1902);
nand U4185 (N_4185,N_2237,N_480);
nor U4186 (N_4186,N_2355,N_343);
nand U4187 (N_4187,N_2320,N_761);
or U4188 (N_4188,N_1030,N_302);
nand U4189 (N_4189,N_436,N_821);
nor U4190 (N_4190,N_1329,N_307);
and U4191 (N_4191,N_1560,N_91);
or U4192 (N_4192,N_451,N_1385);
nor U4193 (N_4193,N_2045,N_1839);
and U4194 (N_4194,N_1306,N_2);
nand U4195 (N_4195,N_1098,N_898);
and U4196 (N_4196,N_1188,N_451);
or U4197 (N_4197,N_874,N_2395);
and U4198 (N_4198,N_1717,N_1224);
and U4199 (N_4199,N_2387,N_2346);
xnor U4200 (N_4200,N_289,N_460);
and U4201 (N_4201,N_2263,N_901);
xnor U4202 (N_4202,N_1189,N_1339);
nor U4203 (N_4203,N_2054,N_1496);
and U4204 (N_4204,N_1426,N_806);
and U4205 (N_4205,N_2015,N_49);
nor U4206 (N_4206,N_1584,N_2025);
and U4207 (N_4207,N_669,N_1691);
nor U4208 (N_4208,N_1562,N_2490);
nor U4209 (N_4209,N_711,N_571);
and U4210 (N_4210,N_1478,N_471);
and U4211 (N_4211,N_203,N_1718);
nor U4212 (N_4212,N_733,N_1501);
xor U4213 (N_4213,N_990,N_1539);
nor U4214 (N_4214,N_2025,N_92);
nand U4215 (N_4215,N_1260,N_1196);
or U4216 (N_4216,N_2313,N_1579);
nor U4217 (N_4217,N_783,N_1422);
nor U4218 (N_4218,N_1440,N_1160);
and U4219 (N_4219,N_1686,N_2347);
nand U4220 (N_4220,N_2059,N_1115);
nand U4221 (N_4221,N_1494,N_1903);
nor U4222 (N_4222,N_550,N_1080);
or U4223 (N_4223,N_1739,N_1803);
nand U4224 (N_4224,N_16,N_42);
nand U4225 (N_4225,N_1290,N_434);
nand U4226 (N_4226,N_788,N_1311);
nand U4227 (N_4227,N_708,N_461);
or U4228 (N_4228,N_2483,N_2381);
and U4229 (N_4229,N_1495,N_765);
xor U4230 (N_4230,N_1603,N_579);
or U4231 (N_4231,N_616,N_835);
xor U4232 (N_4232,N_668,N_216);
xor U4233 (N_4233,N_1871,N_2196);
or U4234 (N_4234,N_2448,N_387);
nor U4235 (N_4235,N_918,N_1460);
and U4236 (N_4236,N_1791,N_1835);
nand U4237 (N_4237,N_1590,N_1246);
nand U4238 (N_4238,N_313,N_2388);
or U4239 (N_4239,N_381,N_791);
xnor U4240 (N_4240,N_2172,N_1783);
nand U4241 (N_4241,N_1916,N_1358);
nand U4242 (N_4242,N_2035,N_520);
and U4243 (N_4243,N_2326,N_2319);
nand U4244 (N_4244,N_2378,N_2219);
xnor U4245 (N_4245,N_1538,N_1092);
or U4246 (N_4246,N_2185,N_1027);
or U4247 (N_4247,N_986,N_284);
or U4248 (N_4248,N_1255,N_406);
and U4249 (N_4249,N_2272,N_1740);
and U4250 (N_4250,N_1470,N_450);
or U4251 (N_4251,N_435,N_776);
nor U4252 (N_4252,N_2212,N_2441);
or U4253 (N_4253,N_829,N_1910);
or U4254 (N_4254,N_704,N_2371);
nor U4255 (N_4255,N_2146,N_531);
or U4256 (N_4256,N_2360,N_1837);
nor U4257 (N_4257,N_1525,N_1345);
or U4258 (N_4258,N_1672,N_1048);
or U4259 (N_4259,N_659,N_2113);
and U4260 (N_4260,N_377,N_381);
nor U4261 (N_4261,N_193,N_1424);
or U4262 (N_4262,N_1883,N_891);
nand U4263 (N_4263,N_116,N_1515);
nand U4264 (N_4264,N_1460,N_1255);
and U4265 (N_4265,N_2057,N_56);
nor U4266 (N_4266,N_51,N_146);
or U4267 (N_4267,N_2265,N_1727);
nand U4268 (N_4268,N_1394,N_168);
nor U4269 (N_4269,N_844,N_1325);
xor U4270 (N_4270,N_2333,N_15);
nand U4271 (N_4271,N_2441,N_1337);
nand U4272 (N_4272,N_1569,N_468);
and U4273 (N_4273,N_596,N_511);
nand U4274 (N_4274,N_276,N_538);
or U4275 (N_4275,N_986,N_1701);
or U4276 (N_4276,N_2350,N_2161);
and U4277 (N_4277,N_1636,N_1236);
or U4278 (N_4278,N_710,N_1005);
xor U4279 (N_4279,N_874,N_865);
and U4280 (N_4280,N_2080,N_2353);
or U4281 (N_4281,N_1858,N_1270);
and U4282 (N_4282,N_316,N_2400);
or U4283 (N_4283,N_1864,N_1472);
nor U4284 (N_4284,N_520,N_710);
and U4285 (N_4285,N_1157,N_1858);
nor U4286 (N_4286,N_2415,N_775);
nand U4287 (N_4287,N_1606,N_1158);
nand U4288 (N_4288,N_752,N_2275);
nor U4289 (N_4289,N_999,N_207);
nand U4290 (N_4290,N_2125,N_14);
and U4291 (N_4291,N_948,N_601);
nor U4292 (N_4292,N_1561,N_2250);
nand U4293 (N_4293,N_855,N_778);
xor U4294 (N_4294,N_531,N_1542);
nand U4295 (N_4295,N_126,N_1229);
nand U4296 (N_4296,N_1741,N_2161);
nand U4297 (N_4297,N_1592,N_349);
and U4298 (N_4298,N_1821,N_752);
and U4299 (N_4299,N_2345,N_2317);
nand U4300 (N_4300,N_2107,N_380);
nor U4301 (N_4301,N_228,N_2293);
nor U4302 (N_4302,N_304,N_1678);
nor U4303 (N_4303,N_2425,N_1783);
or U4304 (N_4304,N_27,N_216);
xnor U4305 (N_4305,N_2262,N_2021);
and U4306 (N_4306,N_83,N_104);
and U4307 (N_4307,N_124,N_863);
nand U4308 (N_4308,N_1850,N_1322);
nor U4309 (N_4309,N_357,N_2169);
xor U4310 (N_4310,N_887,N_2198);
nor U4311 (N_4311,N_1568,N_1861);
xor U4312 (N_4312,N_1206,N_874);
or U4313 (N_4313,N_1287,N_1184);
nor U4314 (N_4314,N_295,N_1735);
and U4315 (N_4315,N_1504,N_609);
nor U4316 (N_4316,N_1484,N_903);
or U4317 (N_4317,N_2344,N_73);
or U4318 (N_4318,N_1897,N_1819);
nor U4319 (N_4319,N_402,N_1863);
or U4320 (N_4320,N_2318,N_1872);
or U4321 (N_4321,N_2069,N_1883);
nor U4322 (N_4322,N_1480,N_202);
xnor U4323 (N_4323,N_1574,N_600);
and U4324 (N_4324,N_1125,N_2211);
or U4325 (N_4325,N_772,N_1676);
nand U4326 (N_4326,N_1795,N_2140);
nor U4327 (N_4327,N_419,N_1249);
nand U4328 (N_4328,N_1461,N_1134);
and U4329 (N_4329,N_581,N_1979);
nand U4330 (N_4330,N_2392,N_2274);
nand U4331 (N_4331,N_369,N_38);
nor U4332 (N_4332,N_1911,N_595);
or U4333 (N_4333,N_1974,N_1663);
nor U4334 (N_4334,N_1975,N_2357);
nor U4335 (N_4335,N_386,N_1186);
nor U4336 (N_4336,N_2039,N_2210);
and U4337 (N_4337,N_1127,N_1331);
xor U4338 (N_4338,N_517,N_1071);
and U4339 (N_4339,N_17,N_608);
nor U4340 (N_4340,N_1218,N_1459);
or U4341 (N_4341,N_2397,N_1060);
or U4342 (N_4342,N_646,N_1566);
nor U4343 (N_4343,N_200,N_1014);
xnor U4344 (N_4344,N_421,N_1211);
and U4345 (N_4345,N_2028,N_507);
nand U4346 (N_4346,N_292,N_530);
or U4347 (N_4347,N_1151,N_7);
or U4348 (N_4348,N_1920,N_1213);
or U4349 (N_4349,N_2070,N_1454);
and U4350 (N_4350,N_2172,N_1546);
nor U4351 (N_4351,N_2261,N_926);
or U4352 (N_4352,N_311,N_711);
and U4353 (N_4353,N_681,N_200);
nor U4354 (N_4354,N_2094,N_1251);
nor U4355 (N_4355,N_1938,N_1244);
nand U4356 (N_4356,N_863,N_1517);
nor U4357 (N_4357,N_1274,N_2283);
xor U4358 (N_4358,N_2425,N_621);
and U4359 (N_4359,N_271,N_354);
or U4360 (N_4360,N_2088,N_1726);
or U4361 (N_4361,N_935,N_1436);
nand U4362 (N_4362,N_1609,N_1763);
nor U4363 (N_4363,N_1939,N_1736);
nand U4364 (N_4364,N_760,N_1610);
nand U4365 (N_4365,N_822,N_475);
xor U4366 (N_4366,N_1959,N_222);
nand U4367 (N_4367,N_1021,N_632);
or U4368 (N_4368,N_337,N_2312);
xor U4369 (N_4369,N_1756,N_1934);
nand U4370 (N_4370,N_637,N_1138);
nand U4371 (N_4371,N_689,N_1022);
nand U4372 (N_4372,N_1819,N_1691);
nand U4373 (N_4373,N_736,N_519);
and U4374 (N_4374,N_2355,N_2161);
nand U4375 (N_4375,N_1842,N_775);
and U4376 (N_4376,N_1557,N_2290);
and U4377 (N_4377,N_2166,N_290);
nand U4378 (N_4378,N_625,N_598);
nor U4379 (N_4379,N_916,N_1043);
nor U4380 (N_4380,N_1328,N_1266);
nand U4381 (N_4381,N_1881,N_1988);
and U4382 (N_4382,N_2079,N_1062);
xnor U4383 (N_4383,N_1854,N_2);
or U4384 (N_4384,N_853,N_890);
and U4385 (N_4385,N_1450,N_494);
nor U4386 (N_4386,N_573,N_1531);
nand U4387 (N_4387,N_2380,N_351);
xnor U4388 (N_4388,N_1120,N_209);
or U4389 (N_4389,N_923,N_1285);
or U4390 (N_4390,N_2328,N_887);
and U4391 (N_4391,N_495,N_1720);
nand U4392 (N_4392,N_1589,N_1428);
or U4393 (N_4393,N_712,N_1105);
xnor U4394 (N_4394,N_1089,N_728);
and U4395 (N_4395,N_959,N_1929);
nand U4396 (N_4396,N_1354,N_2027);
or U4397 (N_4397,N_451,N_1473);
nand U4398 (N_4398,N_477,N_268);
nor U4399 (N_4399,N_2184,N_1379);
nor U4400 (N_4400,N_952,N_1038);
nand U4401 (N_4401,N_56,N_713);
nand U4402 (N_4402,N_886,N_386);
or U4403 (N_4403,N_2243,N_368);
nor U4404 (N_4404,N_1626,N_1305);
xor U4405 (N_4405,N_719,N_35);
or U4406 (N_4406,N_138,N_377);
and U4407 (N_4407,N_875,N_1071);
nand U4408 (N_4408,N_576,N_1988);
nor U4409 (N_4409,N_673,N_1932);
or U4410 (N_4410,N_354,N_2087);
nand U4411 (N_4411,N_2179,N_1696);
nand U4412 (N_4412,N_1798,N_2115);
nand U4413 (N_4413,N_434,N_1849);
and U4414 (N_4414,N_1115,N_2079);
nand U4415 (N_4415,N_1885,N_1434);
or U4416 (N_4416,N_986,N_1841);
and U4417 (N_4417,N_830,N_853);
nor U4418 (N_4418,N_934,N_238);
nor U4419 (N_4419,N_675,N_1494);
nor U4420 (N_4420,N_2139,N_731);
nor U4421 (N_4421,N_1724,N_1920);
and U4422 (N_4422,N_994,N_1781);
nor U4423 (N_4423,N_732,N_1297);
and U4424 (N_4424,N_981,N_896);
or U4425 (N_4425,N_1005,N_1601);
nand U4426 (N_4426,N_269,N_67);
and U4427 (N_4427,N_1261,N_2274);
xnor U4428 (N_4428,N_2212,N_2269);
nand U4429 (N_4429,N_174,N_1731);
and U4430 (N_4430,N_1432,N_2299);
and U4431 (N_4431,N_1274,N_1446);
nand U4432 (N_4432,N_1215,N_1802);
or U4433 (N_4433,N_715,N_301);
and U4434 (N_4434,N_822,N_164);
or U4435 (N_4435,N_947,N_1178);
xnor U4436 (N_4436,N_1030,N_1699);
nor U4437 (N_4437,N_220,N_237);
nand U4438 (N_4438,N_2410,N_24);
nand U4439 (N_4439,N_95,N_2065);
nor U4440 (N_4440,N_312,N_1207);
nor U4441 (N_4441,N_1593,N_1021);
and U4442 (N_4442,N_981,N_219);
and U4443 (N_4443,N_1961,N_421);
and U4444 (N_4444,N_809,N_488);
nor U4445 (N_4445,N_2495,N_458);
nor U4446 (N_4446,N_2456,N_1872);
nand U4447 (N_4447,N_952,N_1136);
nand U4448 (N_4448,N_486,N_82);
nand U4449 (N_4449,N_2090,N_451);
and U4450 (N_4450,N_1629,N_276);
or U4451 (N_4451,N_1988,N_1031);
and U4452 (N_4452,N_1954,N_2307);
and U4453 (N_4453,N_930,N_12);
nand U4454 (N_4454,N_345,N_1532);
or U4455 (N_4455,N_1561,N_758);
nor U4456 (N_4456,N_1691,N_1155);
nor U4457 (N_4457,N_1430,N_87);
or U4458 (N_4458,N_716,N_943);
or U4459 (N_4459,N_1395,N_97);
xor U4460 (N_4460,N_1915,N_1280);
and U4461 (N_4461,N_1009,N_125);
nor U4462 (N_4462,N_902,N_2257);
or U4463 (N_4463,N_2172,N_2023);
nand U4464 (N_4464,N_2082,N_1732);
nand U4465 (N_4465,N_2146,N_1410);
and U4466 (N_4466,N_1102,N_849);
and U4467 (N_4467,N_2401,N_196);
and U4468 (N_4468,N_2187,N_274);
and U4469 (N_4469,N_585,N_329);
nor U4470 (N_4470,N_283,N_1907);
and U4471 (N_4471,N_1989,N_2111);
and U4472 (N_4472,N_482,N_1111);
nor U4473 (N_4473,N_1990,N_1109);
xor U4474 (N_4474,N_1781,N_701);
nor U4475 (N_4475,N_1747,N_2451);
nand U4476 (N_4476,N_756,N_1949);
nand U4477 (N_4477,N_1494,N_1706);
and U4478 (N_4478,N_1555,N_1323);
nor U4479 (N_4479,N_1045,N_1003);
xnor U4480 (N_4480,N_1843,N_861);
xnor U4481 (N_4481,N_907,N_582);
nor U4482 (N_4482,N_2372,N_1168);
and U4483 (N_4483,N_1604,N_265);
or U4484 (N_4484,N_2294,N_1956);
nor U4485 (N_4485,N_125,N_1278);
or U4486 (N_4486,N_2299,N_1233);
xor U4487 (N_4487,N_257,N_700);
or U4488 (N_4488,N_1830,N_1234);
nor U4489 (N_4489,N_523,N_1429);
nand U4490 (N_4490,N_1553,N_1112);
nand U4491 (N_4491,N_515,N_740);
nand U4492 (N_4492,N_2031,N_895);
nor U4493 (N_4493,N_2279,N_749);
and U4494 (N_4494,N_1225,N_1058);
nand U4495 (N_4495,N_1795,N_138);
nor U4496 (N_4496,N_1716,N_84);
nand U4497 (N_4497,N_2485,N_1729);
nand U4498 (N_4498,N_1617,N_1633);
nand U4499 (N_4499,N_2099,N_1636);
nand U4500 (N_4500,N_371,N_1797);
or U4501 (N_4501,N_1589,N_1120);
nor U4502 (N_4502,N_2265,N_324);
nand U4503 (N_4503,N_866,N_656);
nor U4504 (N_4504,N_125,N_464);
nand U4505 (N_4505,N_42,N_2454);
nor U4506 (N_4506,N_951,N_1333);
nand U4507 (N_4507,N_2195,N_550);
nand U4508 (N_4508,N_1894,N_708);
nand U4509 (N_4509,N_600,N_46);
and U4510 (N_4510,N_1568,N_967);
nand U4511 (N_4511,N_1243,N_26);
and U4512 (N_4512,N_2345,N_2004);
nor U4513 (N_4513,N_633,N_1218);
nand U4514 (N_4514,N_1649,N_1739);
or U4515 (N_4515,N_847,N_993);
nor U4516 (N_4516,N_631,N_1117);
nor U4517 (N_4517,N_1758,N_2078);
or U4518 (N_4518,N_2270,N_333);
nand U4519 (N_4519,N_361,N_2188);
and U4520 (N_4520,N_1941,N_2287);
nor U4521 (N_4521,N_1317,N_1214);
nand U4522 (N_4522,N_283,N_452);
and U4523 (N_4523,N_1486,N_2131);
and U4524 (N_4524,N_2217,N_564);
nand U4525 (N_4525,N_2454,N_1509);
nor U4526 (N_4526,N_1053,N_2132);
and U4527 (N_4527,N_933,N_2358);
nand U4528 (N_4528,N_1883,N_2335);
and U4529 (N_4529,N_2154,N_2329);
nor U4530 (N_4530,N_262,N_909);
nand U4531 (N_4531,N_154,N_1631);
xnor U4532 (N_4532,N_1760,N_2089);
and U4533 (N_4533,N_1648,N_1628);
and U4534 (N_4534,N_1309,N_195);
nand U4535 (N_4535,N_1607,N_2318);
or U4536 (N_4536,N_1397,N_732);
and U4537 (N_4537,N_2369,N_483);
nor U4538 (N_4538,N_738,N_1925);
nor U4539 (N_4539,N_2318,N_2122);
nand U4540 (N_4540,N_1735,N_612);
nor U4541 (N_4541,N_616,N_2495);
nor U4542 (N_4542,N_1705,N_2167);
or U4543 (N_4543,N_1714,N_214);
xnor U4544 (N_4544,N_499,N_2006);
nand U4545 (N_4545,N_451,N_718);
or U4546 (N_4546,N_1916,N_1713);
or U4547 (N_4547,N_1238,N_312);
nor U4548 (N_4548,N_1885,N_161);
or U4549 (N_4549,N_1325,N_70);
nor U4550 (N_4550,N_1257,N_2288);
nor U4551 (N_4551,N_2300,N_899);
nand U4552 (N_4552,N_627,N_2085);
nand U4553 (N_4553,N_1183,N_1657);
xor U4554 (N_4554,N_1615,N_1746);
nor U4555 (N_4555,N_255,N_623);
or U4556 (N_4556,N_1083,N_2313);
nand U4557 (N_4557,N_607,N_1324);
and U4558 (N_4558,N_565,N_1145);
and U4559 (N_4559,N_1782,N_1930);
nand U4560 (N_4560,N_2167,N_2173);
or U4561 (N_4561,N_780,N_516);
or U4562 (N_4562,N_1566,N_1916);
nor U4563 (N_4563,N_48,N_224);
and U4564 (N_4564,N_2429,N_665);
nand U4565 (N_4565,N_1164,N_52);
nor U4566 (N_4566,N_1834,N_470);
nor U4567 (N_4567,N_2290,N_213);
nor U4568 (N_4568,N_1985,N_428);
or U4569 (N_4569,N_1366,N_2000);
nor U4570 (N_4570,N_966,N_124);
nand U4571 (N_4571,N_2067,N_467);
and U4572 (N_4572,N_1080,N_884);
nand U4573 (N_4573,N_391,N_1458);
nand U4574 (N_4574,N_2143,N_2391);
xor U4575 (N_4575,N_1515,N_1301);
and U4576 (N_4576,N_2013,N_1172);
or U4577 (N_4577,N_984,N_817);
xnor U4578 (N_4578,N_1073,N_2032);
or U4579 (N_4579,N_1865,N_834);
or U4580 (N_4580,N_2360,N_708);
nor U4581 (N_4581,N_2044,N_555);
xnor U4582 (N_4582,N_1144,N_310);
nand U4583 (N_4583,N_1806,N_741);
xor U4584 (N_4584,N_1282,N_1123);
nor U4585 (N_4585,N_41,N_1572);
nand U4586 (N_4586,N_242,N_1599);
or U4587 (N_4587,N_665,N_2445);
nand U4588 (N_4588,N_558,N_992);
nor U4589 (N_4589,N_126,N_912);
nand U4590 (N_4590,N_221,N_524);
and U4591 (N_4591,N_2095,N_790);
nor U4592 (N_4592,N_2061,N_1045);
or U4593 (N_4593,N_637,N_2187);
nand U4594 (N_4594,N_1073,N_442);
nor U4595 (N_4595,N_31,N_700);
or U4596 (N_4596,N_2283,N_715);
and U4597 (N_4597,N_58,N_298);
and U4598 (N_4598,N_1337,N_1095);
xor U4599 (N_4599,N_234,N_1010);
or U4600 (N_4600,N_1610,N_516);
and U4601 (N_4601,N_1872,N_1298);
nand U4602 (N_4602,N_474,N_1305);
or U4603 (N_4603,N_933,N_60);
nor U4604 (N_4604,N_1079,N_156);
nor U4605 (N_4605,N_963,N_142);
xnor U4606 (N_4606,N_2222,N_1861);
nor U4607 (N_4607,N_2327,N_891);
xnor U4608 (N_4608,N_2185,N_2276);
nand U4609 (N_4609,N_1826,N_1565);
nor U4610 (N_4610,N_1489,N_999);
or U4611 (N_4611,N_1746,N_2306);
nand U4612 (N_4612,N_1770,N_2309);
or U4613 (N_4613,N_452,N_260);
or U4614 (N_4614,N_13,N_895);
nor U4615 (N_4615,N_1697,N_2401);
and U4616 (N_4616,N_2392,N_1300);
xnor U4617 (N_4617,N_939,N_2268);
nor U4618 (N_4618,N_551,N_27);
xnor U4619 (N_4619,N_1354,N_2447);
and U4620 (N_4620,N_2441,N_1716);
nor U4621 (N_4621,N_2361,N_2275);
or U4622 (N_4622,N_132,N_0);
or U4623 (N_4623,N_56,N_1961);
xor U4624 (N_4624,N_2173,N_45);
or U4625 (N_4625,N_2261,N_2469);
xnor U4626 (N_4626,N_648,N_670);
or U4627 (N_4627,N_2335,N_1794);
nand U4628 (N_4628,N_2029,N_2239);
and U4629 (N_4629,N_904,N_2035);
and U4630 (N_4630,N_1170,N_60);
nand U4631 (N_4631,N_285,N_2224);
nor U4632 (N_4632,N_1734,N_2353);
or U4633 (N_4633,N_362,N_210);
nand U4634 (N_4634,N_1236,N_451);
nand U4635 (N_4635,N_1965,N_1386);
nand U4636 (N_4636,N_264,N_118);
or U4637 (N_4637,N_1053,N_2161);
or U4638 (N_4638,N_974,N_632);
or U4639 (N_4639,N_1339,N_154);
xor U4640 (N_4640,N_1093,N_1913);
nor U4641 (N_4641,N_134,N_1209);
nor U4642 (N_4642,N_752,N_1029);
and U4643 (N_4643,N_1213,N_575);
and U4644 (N_4644,N_1293,N_2279);
nor U4645 (N_4645,N_2259,N_270);
and U4646 (N_4646,N_974,N_408);
and U4647 (N_4647,N_735,N_1348);
and U4648 (N_4648,N_2188,N_1600);
nor U4649 (N_4649,N_717,N_780);
xor U4650 (N_4650,N_192,N_2287);
xnor U4651 (N_4651,N_1519,N_33);
and U4652 (N_4652,N_1586,N_1019);
nor U4653 (N_4653,N_1960,N_694);
and U4654 (N_4654,N_1441,N_1222);
or U4655 (N_4655,N_639,N_528);
nand U4656 (N_4656,N_763,N_579);
nand U4657 (N_4657,N_1983,N_1217);
or U4658 (N_4658,N_1383,N_875);
nor U4659 (N_4659,N_142,N_1290);
nand U4660 (N_4660,N_914,N_2453);
or U4661 (N_4661,N_312,N_1546);
or U4662 (N_4662,N_254,N_2305);
xnor U4663 (N_4663,N_610,N_377);
nand U4664 (N_4664,N_43,N_637);
or U4665 (N_4665,N_1566,N_712);
nand U4666 (N_4666,N_502,N_2410);
and U4667 (N_4667,N_128,N_1703);
nand U4668 (N_4668,N_1207,N_1677);
nand U4669 (N_4669,N_1909,N_524);
nor U4670 (N_4670,N_1504,N_1318);
and U4671 (N_4671,N_2252,N_473);
or U4672 (N_4672,N_139,N_279);
nand U4673 (N_4673,N_2214,N_547);
nand U4674 (N_4674,N_2169,N_1523);
nor U4675 (N_4675,N_797,N_1254);
nor U4676 (N_4676,N_1873,N_1441);
and U4677 (N_4677,N_1816,N_107);
nand U4678 (N_4678,N_688,N_706);
or U4679 (N_4679,N_569,N_1502);
and U4680 (N_4680,N_420,N_94);
nor U4681 (N_4681,N_1305,N_171);
or U4682 (N_4682,N_945,N_1741);
nor U4683 (N_4683,N_2087,N_1708);
or U4684 (N_4684,N_588,N_617);
nor U4685 (N_4685,N_844,N_1527);
xnor U4686 (N_4686,N_1457,N_365);
nor U4687 (N_4687,N_804,N_764);
and U4688 (N_4688,N_1168,N_1613);
or U4689 (N_4689,N_1429,N_884);
or U4690 (N_4690,N_1154,N_2285);
nand U4691 (N_4691,N_594,N_2327);
or U4692 (N_4692,N_64,N_783);
nor U4693 (N_4693,N_2255,N_88);
or U4694 (N_4694,N_961,N_1112);
or U4695 (N_4695,N_2170,N_677);
and U4696 (N_4696,N_2266,N_2275);
and U4697 (N_4697,N_1353,N_569);
and U4698 (N_4698,N_1417,N_48);
nor U4699 (N_4699,N_645,N_797);
nand U4700 (N_4700,N_2200,N_844);
xor U4701 (N_4701,N_2321,N_575);
and U4702 (N_4702,N_2262,N_1288);
and U4703 (N_4703,N_675,N_957);
xnor U4704 (N_4704,N_2150,N_147);
and U4705 (N_4705,N_230,N_36);
and U4706 (N_4706,N_538,N_961);
nor U4707 (N_4707,N_2391,N_1575);
nor U4708 (N_4708,N_1077,N_2141);
nand U4709 (N_4709,N_1734,N_69);
or U4710 (N_4710,N_385,N_1209);
nand U4711 (N_4711,N_798,N_847);
nand U4712 (N_4712,N_179,N_1159);
nor U4713 (N_4713,N_487,N_1816);
nor U4714 (N_4714,N_72,N_1666);
and U4715 (N_4715,N_270,N_95);
xor U4716 (N_4716,N_1822,N_703);
nor U4717 (N_4717,N_1562,N_1063);
nand U4718 (N_4718,N_591,N_1301);
and U4719 (N_4719,N_419,N_1740);
nor U4720 (N_4720,N_2082,N_1021);
or U4721 (N_4721,N_1379,N_2478);
nor U4722 (N_4722,N_694,N_906);
nor U4723 (N_4723,N_571,N_625);
or U4724 (N_4724,N_250,N_926);
xnor U4725 (N_4725,N_1977,N_2165);
nor U4726 (N_4726,N_2015,N_1672);
and U4727 (N_4727,N_1505,N_1185);
nor U4728 (N_4728,N_1721,N_1192);
or U4729 (N_4729,N_242,N_1825);
nor U4730 (N_4730,N_1198,N_1465);
and U4731 (N_4731,N_1489,N_827);
xnor U4732 (N_4732,N_1399,N_1940);
nand U4733 (N_4733,N_36,N_2411);
or U4734 (N_4734,N_2073,N_2002);
nor U4735 (N_4735,N_1728,N_1750);
or U4736 (N_4736,N_2044,N_1473);
and U4737 (N_4737,N_1804,N_1434);
nor U4738 (N_4738,N_1235,N_2357);
and U4739 (N_4739,N_1851,N_1224);
or U4740 (N_4740,N_1406,N_341);
xnor U4741 (N_4741,N_1422,N_1567);
xor U4742 (N_4742,N_1387,N_2313);
or U4743 (N_4743,N_1708,N_1111);
and U4744 (N_4744,N_1015,N_2135);
nand U4745 (N_4745,N_1001,N_2392);
nor U4746 (N_4746,N_1980,N_1218);
and U4747 (N_4747,N_2337,N_1038);
nor U4748 (N_4748,N_42,N_1234);
or U4749 (N_4749,N_772,N_1982);
nand U4750 (N_4750,N_138,N_442);
and U4751 (N_4751,N_1009,N_566);
nand U4752 (N_4752,N_61,N_918);
nand U4753 (N_4753,N_168,N_2446);
nand U4754 (N_4754,N_820,N_2447);
nand U4755 (N_4755,N_1377,N_2095);
and U4756 (N_4756,N_774,N_1091);
and U4757 (N_4757,N_1501,N_474);
or U4758 (N_4758,N_2345,N_8);
nor U4759 (N_4759,N_818,N_400);
or U4760 (N_4760,N_1170,N_11);
and U4761 (N_4761,N_1239,N_2432);
nand U4762 (N_4762,N_1755,N_1796);
nor U4763 (N_4763,N_583,N_481);
or U4764 (N_4764,N_1098,N_1591);
and U4765 (N_4765,N_842,N_1259);
xnor U4766 (N_4766,N_2153,N_2020);
or U4767 (N_4767,N_1692,N_1771);
or U4768 (N_4768,N_1094,N_993);
nor U4769 (N_4769,N_1938,N_1808);
or U4770 (N_4770,N_2380,N_1099);
and U4771 (N_4771,N_311,N_2148);
nor U4772 (N_4772,N_547,N_617);
nand U4773 (N_4773,N_905,N_842);
and U4774 (N_4774,N_1293,N_17);
and U4775 (N_4775,N_281,N_1194);
xnor U4776 (N_4776,N_1822,N_600);
and U4777 (N_4777,N_1332,N_1875);
and U4778 (N_4778,N_1427,N_1982);
nand U4779 (N_4779,N_230,N_2135);
and U4780 (N_4780,N_2091,N_1142);
and U4781 (N_4781,N_2223,N_564);
and U4782 (N_4782,N_2201,N_1305);
and U4783 (N_4783,N_2257,N_647);
and U4784 (N_4784,N_558,N_1673);
nor U4785 (N_4785,N_2269,N_2315);
or U4786 (N_4786,N_2188,N_1478);
and U4787 (N_4787,N_486,N_2262);
or U4788 (N_4788,N_89,N_1980);
nand U4789 (N_4789,N_1363,N_2274);
or U4790 (N_4790,N_2151,N_1045);
nor U4791 (N_4791,N_1736,N_1404);
nand U4792 (N_4792,N_879,N_2081);
nor U4793 (N_4793,N_999,N_1994);
nor U4794 (N_4794,N_2035,N_166);
nor U4795 (N_4795,N_1909,N_765);
and U4796 (N_4796,N_1749,N_1187);
and U4797 (N_4797,N_1877,N_1880);
and U4798 (N_4798,N_315,N_1110);
nor U4799 (N_4799,N_563,N_1208);
and U4800 (N_4800,N_74,N_1542);
nor U4801 (N_4801,N_819,N_2049);
nand U4802 (N_4802,N_925,N_1004);
and U4803 (N_4803,N_677,N_1112);
nand U4804 (N_4804,N_1531,N_563);
nand U4805 (N_4805,N_1809,N_409);
xor U4806 (N_4806,N_1101,N_1055);
or U4807 (N_4807,N_1534,N_985);
or U4808 (N_4808,N_1398,N_2179);
nor U4809 (N_4809,N_45,N_970);
nor U4810 (N_4810,N_141,N_1813);
xor U4811 (N_4811,N_169,N_2101);
nand U4812 (N_4812,N_1349,N_44);
xor U4813 (N_4813,N_1541,N_2085);
nor U4814 (N_4814,N_42,N_1792);
and U4815 (N_4815,N_2062,N_1373);
nor U4816 (N_4816,N_1655,N_1028);
nand U4817 (N_4817,N_1276,N_1382);
nand U4818 (N_4818,N_209,N_746);
nor U4819 (N_4819,N_1820,N_516);
nor U4820 (N_4820,N_1632,N_1871);
or U4821 (N_4821,N_271,N_1289);
nand U4822 (N_4822,N_1472,N_1847);
or U4823 (N_4823,N_769,N_437);
and U4824 (N_4824,N_298,N_1234);
nor U4825 (N_4825,N_308,N_952);
or U4826 (N_4826,N_430,N_1493);
nor U4827 (N_4827,N_2047,N_648);
nand U4828 (N_4828,N_1263,N_1008);
nand U4829 (N_4829,N_256,N_453);
and U4830 (N_4830,N_2181,N_167);
nand U4831 (N_4831,N_1214,N_108);
nand U4832 (N_4832,N_1733,N_32);
nand U4833 (N_4833,N_1945,N_2379);
nor U4834 (N_4834,N_1256,N_717);
or U4835 (N_4835,N_469,N_776);
or U4836 (N_4836,N_310,N_1731);
nor U4837 (N_4837,N_1952,N_1607);
xor U4838 (N_4838,N_1523,N_930);
and U4839 (N_4839,N_2084,N_1429);
nand U4840 (N_4840,N_1419,N_24);
and U4841 (N_4841,N_1306,N_1282);
nand U4842 (N_4842,N_1056,N_1720);
nand U4843 (N_4843,N_1183,N_2497);
nand U4844 (N_4844,N_2011,N_839);
and U4845 (N_4845,N_2369,N_1247);
and U4846 (N_4846,N_1759,N_958);
nor U4847 (N_4847,N_884,N_2290);
nand U4848 (N_4848,N_301,N_2060);
nand U4849 (N_4849,N_1475,N_759);
and U4850 (N_4850,N_683,N_2357);
nor U4851 (N_4851,N_1928,N_2318);
or U4852 (N_4852,N_1298,N_1211);
nor U4853 (N_4853,N_1412,N_606);
and U4854 (N_4854,N_1599,N_2357);
nand U4855 (N_4855,N_2028,N_233);
and U4856 (N_4856,N_2312,N_1225);
nor U4857 (N_4857,N_829,N_1907);
or U4858 (N_4858,N_2379,N_570);
or U4859 (N_4859,N_342,N_578);
nand U4860 (N_4860,N_288,N_442);
nand U4861 (N_4861,N_521,N_1180);
nor U4862 (N_4862,N_1652,N_2419);
nor U4863 (N_4863,N_634,N_1319);
and U4864 (N_4864,N_1458,N_2195);
or U4865 (N_4865,N_2020,N_1904);
nor U4866 (N_4866,N_331,N_1710);
nand U4867 (N_4867,N_827,N_969);
and U4868 (N_4868,N_619,N_2423);
nor U4869 (N_4869,N_692,N_112);
nand U4870 (N_4870,N_43,N_1412);
and U4871 (N_4871,N_1445,N_1592);
and U4872 (N_4872,N_135,N_77);
or U4873 (N_4873,N_1789,N_1795);
and U4874 (N_4874,N_1583,N_2208);
xor U4875 (N_4875,N_2334,N_1411);
nand U4876 (N_4876,N_2431,N_2266);
and U4877 (N_4877,N_730,N_1528);
or U4878 (N_4878,N_67,N_1910);
nor U4879 (N_4879,N_1127,N_2314);
nand U4880 (N_4880,N_270,N_1689);
nor U4881 (N_4881,N_61,N_1508);
nand U4882 (N_4882,N_1785,N_1524);
nor U4883 (N_4883,N_128,N_481);
nand U4884 (N_4884,N_2418,N_1191);
and U4885 (N_4885,N_2303,N_874);
and U4886 (N_4886,N_446,N_1623);
and U4887 (N_4887,N_322,N_1148);
xnor U4888 (N_4888,N_2493,N_1843);
and U4889 (N_4889,N_1590,N_388);
nor U4890 (N_4890,N_2441,N_2011);
nor U4891 (N_4891,N_1956,N_239);
nand U4892 (N_4892,N_967,N_2499);
nand U4893 (N_4893,N_1695,N_1699);
or U4894 (N_4894,N_540,N_2398);
or U4895 (N_4895,N_494,N_816);
or U4896 (N_4896,N_429,N_1452);
and U4897 (N_4897,N_1668,N_1301);
or U4898 (N_4898,N_560,N_691);
nand U4899 (N_4899,N_1167,N_302);
xnor U4900 (N_4900,N_2492,N_2167);
nor U4901 (N_4901,N_1219,N_1242);
or U4902 (N_4902,N_1579,N_1551);
and U4903 (N_4903,N_784,N_2370);
xor U4904 (N_4904,N_291,N_1349);
nand U4905 (N_4905,N_1735,N_1574);
nand U4906 (N_4906,N_2399,N_1558);
nor U4907 (N_4907,N_1110,N_803);
or U4908 (N_4908,N_542,N_911);
or U4909 (N_4909,N_1831,N_257);
and U4910 (N_4910,N_2450,N_2019);
nand U4911 (N_4911,N_123,N_1222);
and U4912 (N_4912,N_406,N_1167);
nor U4913 (N_4913,N_719,N_673);
nand U4914 (N_4914,N_414,N_713);
or U4915 (N_4915,N_1874,N_123);
nand U4916 (N_4916,N_2044,N_396);
nor U4917 (N_4917,N_832,N_1037);
or U4918 (N_4918,N_1373,N_90);
xnor U4919 (N_4919,N_1025,N_1802);
and U4920 (N_4920,N_2229,N_2078);
xnor U4921 (N_4921,N_602,N_978);
or U4922 (N_4922,N_1630,N_2075);
and U4923 (N_4923,N_2026,N_1364);
or U4924 (N_4924,N_1129,N_1447);
nand U4925 (N_4925,N_64,N_350);
nor U4926 (N_4926,N_2449,N_1730);
nand U4927 (N_4927,N_296,N_812);
or U4928 (N_4928,N_1184,N_2401);
nand U4929 (N_4929,N_164,N_35);
and U4930 (N_4930,N_2122,N_2493);
nand U4931 (N_4931,N_2147,N_1197);
and U4932 (N_4932,N_1506,N_933);
nand U4933 (N_4933,N_222,N_512);
nor U4934 (N_4934,N_94,N_2099);
or U4935 (N_4935,N_1826,N_1307);
nand U4936 (N_4936,N_1994,N_258);
nor U4937 (N_4937,N_678,N_926);
nor U4938 (N_4938,N_2401,N_806);
nand U4939 (N_4939,N_1635,N_677);
nand U4940 (N_4940,N_1344,N_1284);
nand U4941 (N_4941,N_66,N_76);
xnor U4942 (N_4942,N_688,N_2443);
or U4943 (N_4943,N_1973,N_1645);
or U4944 (N_4944,N_1211,N_1048);
nand U4945 (N_4945,N_1730,N_11);
or U4946 (N_4946,N_2468,N_1214);
and U4947 (N_4947,N_933,N_2185);
and U4948 (N_4948,N_165,N_2068);
or U4949 (N_4949,N_1618,N_467);
or U4950 (N_4950,N_1996,N_766);
or U4951 (N_4951,N_1862,N_1386);
or U4952 (N_4952,N_2306,N_1014);
nand U4953 (N_4953,N_894,N_212);
and U4954 (N_4954,N_1152,N_32);
nand U4955 (N_4955,N_1976,N_115);
nor U4956 (N_4956,N_1004,N_2204);
or U4957 (N_4957,N_65,N_2049);
nor U4958 (N_4958,N_759,N_562);
nor U4959 (N_4959,N_2499,N_766);
nor U4960 (N_4960,N_666,N_1731);
and U4961 (N_4961,N_560,N_1852);
xnor U4962 (N_4962,N_80,N_1951);
nand U4963 (N_4963,N_1145,N_2044);
xnor U4964 (N_4964,N_750,N_2218);
nor U4965 (N_4965,N_263,N_2461);
nand U4966 (N_4966,N_1824,N_1382);
nor U4967 (N_4967,N_1762,N_137);
nor U4968 (N_4968,N_307,N_758);
nand U4969 (N_4969,N_1318,N_1526);
nand U4970 (N_4970,N_2139,N_518);
xnor U4971 (N_4971,N_491,N_1802);
nand U4972 (N_4972,N_1956,N_1080);
nand U4973 (N_4973,N_1888,N_1959);
or U4974 (N_4974,N_169,N_1038);
xnor U4975 (N_4975,N_2415,N_2159);
xnor U4976 (N_4976,N_1604,N_637);
or U4977 (N_4977,N_1033,N_1316);
nor U4978 (N_4978,N_1983,N_130);
or U4979 (N_4979,N_1995,N_1916);
and U4980 (N_4980,N_1177,N_1909);
nor U4981 (N_4981,N_1590,N_1442);
and U4982 (N_4982,N_1804,N_87);
and U4983 (N_4983,N_1357,N_473);
and U4984 (N_4984,N_2338,N_1604);
or U4985 (N_4985,N_1911,N_938);
or U4986 (N_4986,N_1038,N_1278);
or U4987 (N_4987,N_1613,N_999);
nand U4988 (N_4988,N_22,N_1340);
nand U4989 (N_4989,N_1871,N_92);
nor U4990 (N_4990,N_315,N_2499);
nor U4991 (N_4991,N_1150,N_2227);
or U4992 (N_4992,N_1816,N_1012);
or U4993 (N_4993,N_721,N_997);
and U4994 (N_4994,N_1547,N_1041);
nor U4995 (N_4995,N_834,N_1391);
nor U4996 (N_4996,N_960,N_2007);
or U4997 (N_4997,N_799,N_576);
and U4998 (N_4998,N_566,N_1837);
and U4999 (N_4999,N_2027,N_249);
nor U5000 (N_5000,N_3275,N_4202);
and U5001 (N_5001,N_3007,N_2883);
or U5002 (N_5002,N_3186,N_3977);
nand U5003 (N_5003,N_3245,N_4056);
and U5004 (N_5004,N_3589,N_4276);
nor U5005 (N_5005,N_3322,N_4092);
nand U5006 (N_5006,N_3013,N_3765);
nor U5007 (N_5007,N_2755,N_3266);
nor U5008 (N_5008,N_3848,N_4689);
and U5009 (N_5009,N_3874,N_3548);
nand U5010 (N_5010,N_2833,N_3715);
or U5011 (N_5011,N_4782,N_4046);
and U5012 (N_5012,N_4924,N_3429);
nand U5013 (N_5013,N_3815,N_2630);
nand U5014 (N_5014,N_4960,N_2684);
nand U5015 (N_5015,N_2825,N_4641);
xnor U5016 (N_5016,N_2893,N_3226);
nand U5017 (N_5017,N_3210,N_3242);
and U5018 (N_5018,N_2814,N_3495);
or U5019 (N_5019,N_2939,N_3507);
nand U5020 (N_5020,N_4721,N_4470);
or U5021 (N_5021,N_3239,N_4115);
or U5022 (N_5022,N_4569,N_4726);
and U5023 (N_5023,N_4822,N_4579);
and U5024 (N_5024,N_3697,N_2777);
xor U5025 (N_5025,N_3571,N_3097);
and U5026 (N_5026,N_4733,N_4356);
nand U5027 (N_5027,N_3936,N_3469);
and U5028 (N_5028,N_2556,N_4362);
and U5029 (N_5029,N_4748,N_4526);
or U5030 (N_5030,N_4973,N_4433);
nand U5031 (N_5031,N_2666,N_3684);
or U5032 (N_5032,N_3636,N_4232);
or U5033 (N_5033,N_4511,N_4057);
nor U5034 (N_5034,N_4919,N_4141);
nand U5035 (N_5035,N_4675,N_4869);
nand U5036 (N_5036,N_3385,N_4576);
and U5037 (N_5037,N_3817,N_3247);
nor U5038 (N_5038,N_2846,N_4347);
nor U5039 (N_5039,N_2652,N_4738);
and U5040 (N_5040,N_4472,N_3283);
and U5041 (N_5041,N_2534,N_3623);
and U5042 (N_5042,N_2874,N_4586);
or U5043 (N_5043,N_3327,N_4997);
nand U5044 (N_5044,N_3798,N_3331);
nand U5045 (N_5045,N_3150,N_4102);
nor U5046 (N_5046,N_2856,N_2980);
nand U5047 (N_5047,N_3596,N_3086);
and U5048 (N_5048,N_4030,N_2806);
and U5049 (N_5049,N_4329,N_2665);
or U5050 (N_5050,N_2809,N_3124);
and U5051 (N_5051,N_4215,N_3825);
and U5052 (N_5052,N_3843,N_4468);
and U5053 (N_5053,N_4193,N_4669);
nand U5054 (N_5054,N_3888,N_2632);
and U5055 (N_5055,N_4553,N_4364);
and U5056 (N_5056,N_3037,N_2798);
nand U5057 (N_5057,N_3199,N_2711);
and U5058 (N_5058,N_3502,N_4596);
and U5059 (N_5059,N_3712,N_4983);
nand U5060 (N_5060,N_4194,N_2881);
or U5061 (N_5061,N_3774,N_3728);
nand U5062 (N_5062,N_3736,N_3145);
nor U5063 (N_5063,N_3036,N_3750);
or U5064 (N_5064,N_2906,N_4004);
nor U5065 (N_5065,N_2947,N_2959);
xor U5066 (N_5066,N_4652,N_3497);
nor U5067 (N_5067,N_3442,N_3237);
nand U5068 (N_5068,N_4839,N_2918);
nand U5069 (N_5069,N_2697,N_2862);
or U5070 (N_5070,N_3346,N_3466);
nor U5071 (N_5071,N_2553,N_4899);
and U5072 (N_5072,N_4577,N_2827);
nand U5073 (N_5073,N_2935,N_3216);
nand U5074 (N_5074,N_3930,N_4547);
or U5075 (N_5075,N_4161,N_3972);
and U5076 (N_5076,N_4771,N_2640);
nand U5077 (N_5077,N_2960,N_3742);
nor U5078 (N_5078,N_4758,N_4851);
or U5079 (N_5079,N_2545,N_3441);
nor U5080 (N_5080,N_2708,N_3414);
nor U5081 (N_5081,N_4327,N_3209);
xnor U5082 (N_5082,N_2966,N_4411);
nor U5083 (N_5083,N_3514,N_3382);
nor U5084 (N_5084,N_3876,N_3590);
or U5085 (N_5085,N_3775,N_2706);
or U5086 (N_5086,N_4500,N_4808);
xor U5087 (N_5087,N_3938,N_2989);
and U5088 (N_5088,N_4506,N_4306);
nand U5089 (N_5089,N_3787,N_2804);
or U5090 (N_5090,N_4213,N_3871);
and U5091 (N_5091,N_4481,N_2902);
or U5092 (N_5092,N_4156,N_3043);
or U5093 (N_5093,N_2657,N_3383);
and U5094 (N_5094,N_3010,N_4892);
nand U5095 (N_5095,N_4795,N_4316);
and U5096 (N_5096,N_3979,N_4012);
or U5097 (N_5097,N_3842,N_3272);
or U5098 (N_5098,N_4251,N_4660);
nor U5099 (N_5099,N_2735,N_2532);
xor U5100 (N_5100,N_3838,N_4204);
nor U5101 (N_5101,N_3473,N_4431);
and U5102 (N_5102,N_3225,N_3480);
nand U5103 (N_5103,N_3873,N_2780);
nor U5104 (N_5104,N_4637,N_2816);
xor U5105 (N_5105,N_4437,N_3082);
nor U5106 (N_5106,N_4461,N_4580);
or U5107 (N_5107,N_2639,N_3986);
and U5108 (N_5108,N_2982,N_4099);
nand U5109 (N_5109,N_2547,N_3132);
or U5110 (N_5110,N_3500,N_3601);
nor U5111 (N_5111,N_2509,N_4294);
nor U5112 (N_5112,N_2851,N_4295);
nand U5113 (N_5113,N_4659,N_3376);
nand U5114 (N_5114,N_2857,N_3880);
and U5115 (N_5115,N_4516,N_3947);
or U5116 (N_5116,N_4959,N_4556);
and U5117 (N_5117,N_3749,N_3129);
and U5118 (N_5118,N_3546,N_2681);
nand U5119 (N_5119,N_4858,N_3030);
nor U5120 (N_5120,N_4107,N_4503);
or U5121 (N_5121,N_4904,N_2572);
nand U5122 (N_5122,N_4015,N_4941);
and U5123 (N_5123,N_2507,N_3791);
xnor U5124 (N_5124,N_4911,N_2835);
nand U5125 (N_5125,N_4163,N_3118);
xor U5126 (N_5126,N_3444,N_4802);
or U5127 (N_5127,N_4335,N_4272);
nor U5128 (N_5128,N_3326,N_3528);
xor U5129 (N_5129,N_2736,N_3052);
nand U5130 (N_5130,N_2828,N_3660);
xor U5131 (N_5131,N_4151,N_2739);
nand U5132 (N_5132,N_2717,N_3300);
or U5133 (N_5133,N_4860,N_4914);
nand U5134 (N_5134,N_4706,N_3181);
xnor U5135 (N_5135,N_4908,N_3614);
or U5136 (N_5136,N_2931,N_3851);
nand U5137 (N_5137,N_4633,N_4837);
and U5138 (N_5138,N_4832,N_3014);
or U5139 (N_5139,N_4751,N_3869);
nand U5140 (N_5140,N_3709,N_2559);
and U5141 (N_5141,N_4293,N_3359);
nand U5142 (N_5142,N_3690,N_3317);
or U5143 (N_5143,N_2970,N_4769);
nor U5144 (N_5144,N_3374,N_3924);
or U5145 (N_5145,N_4289,N_2557);
and U5146 (N_5146,N_4268,N_3185);
xor U5147 (N_5147,N_2675,N_4760);
and U5148 (N_5148,N_3106,N_3920);
nand U5149 (N_5149,N_3021,N_4302);
nand U5150 (N_5150,N_3421,N_4352);
nand U5151 (N_5151,N_4361,N_3723);
or U5152 (N_5152,N_3913,N_3306);
nor U5153 (N_5153,N_2913,N_4666);
xor U5154 (N_5154,N_3609,N_4820);
and U5155 (N_5155,N_3653,N_3779);
nor U5156 (N_5156,N_3987,N_3463);
nor U5157 (N_5157,N_2741,N_4985);
nor U5158 (N_5158,N_4138,N_3948);
xor U5159 (N_5159,N_2868,N_3515);
nor U5160 (N_5160,N_4389,N_2535);
or U5161 (N_5161,N_4703,N_2818);
xnor U5162 (N_5162,N_4891,N_3789);
nand U5163 (N_5163,N_2709,N_4342);
nor U5164 (N_5164,N_4994,N_4608);
or U5165 (N_5165,N_2945,N_3155);
or U5166 (N_5166,N_4429,N_3436);
nor U5167 (N_5167,N_3470,N_4290);
nand U5168 (N_5168,N_3627,N_4281);
and U5169 (N_5169,N_4712,N_3137);
or U5170 (N_5170,N_3751,N_3767);
nor U5171 (N_5171,N_4585,N_3064);
xnor U5172 (N_5172,N_4300,N_3070);
and U5173 (N_5173,N_3719,N_3868);
nand U5174 (N_5174,N_3941,N_4076);
and U5175 (N_5175,N_4118,N_4385);
nand U5176 (N_5176,N_4223,N_3567);
or U5177 (N_5177,N_4113,N_4021);
and U5178 (N_5178,N_3015,N_4693);
nand U5179 (N_5179,N_3020,N_3380);
and U5180 (N_5180,N_4010,N_3295);
and U5181 (N_5181,N_2569,N_4977);
or U5182 (N_5182,N_4520,N_3762);
nor U5183 (N_5183,N_3487,N_2589);
xor U5184 (N_5184,N_4862,N_2979);
nand U5185 (N_5185,N_3333,N_2936);
nor U5186 (N_5186,N_4797,N_2949);
or U5187 (N_5187,N_4307,N_3356);
nand U5188 (N_5188,N_3364,N_3894);
nand U5189 (N_5189,N_4403,N_4685);
and U5190 (N_5190,N_4755,N_3416);
nand U5191 (N_5191,N_4578,N_3363);
xnor U5192 (N_5192,N_3864,N_4691);
nand U5193 (N_5193,N_3622,N_2585);
nand U5194 (N_5194,N_3286,N_2648);
or U5195 (N_5195,N_3565,N_4589);
or U5196 (N_5196,N_2552,N_2571);
or U5197 (N_5197,N_4388,N_4286);
nand U5198 (N_5198,N_4434,N_3800);
nand U5199 (N_5199,N_2782,N_3566);
nand U5200 (N_5200,N_4939,N_4753);
nor U5201 (N_5201,N_2996,N_4047);
nor U5202 (N_5202,N_4765,N_4148);
or U5203 (N_5203,N_4786,N_4273);
or U5204 (N_5204,N_2712,N_3157);
and U5205 (N_5205,N_3475,N_3974);
and U5206 (N_5206,N_2933,N_4017);
nand U5207 (N_5207,N_3462,N_4773);
or U5208 (N_5208,N_3555,N_4331);
nand U5209 (N_5209,N_2824,N_4700);
nand U5210 (N_5210,N_4583,N_4390);
nor U5211 (N_5211,N_2616,N_4261);
nor U5212 (N_5212,N_2749,N_3572);
or U5213 (N_5213,N_4709,N_2978);
and U5214 (N_5214,N_2500,N_4715);
or U5215 (N_5215,N_3320,N_2638);
xnor U5216 (N_5216,N_3553,N_2860);
or U5217 (N_5217,N_4681,N_4146);
or U5218 (N_5218,N_2529,N_3193);
or U5219 (N_5219,N_3141,N_3588);
and U5220 (N_5220,N_4916,N_4640);
or U5221 (N_5221,N_3189,N_4946);
nand U5222 (N_5222,N_4512,N_4953);
xor U5223 (N_5223,N_4182,N_4925);
and U5224 (N_5224,N_4680,N_2718);
nand U5225 (N_5225,N_4843,N_3091);
or U5226 (N_5226,N_3178,N_3228);
nor U5227 (N_5227,N_3928,N_4616);
and U5228 (N_5228,N_4117,N_3744);
nand U5229 (N_5229,N_3362,N_4764);
nand U5230 (N_5230,N_2924,N_2727);
or U5231 (N_5231,N_3998,N_4311);
xor U5232 (N_5232,N_3665,N_4699);
nor U5233 (N_5233,N_4610,N_3618);
or U5234 (N_5234,N_3695,N_2597);
xnor U5235 (N_5235,N_4000,N_3780);
and U5236 (N_5236,N_4452,N_3822);
and U5237 (N_5237,N_3630,N_3398);
xnor U5238 (N_5238,N_4915,N_2864);
or U5239 (N_5239,N_2591,N_3976);
nand U5240 (N_5240,N_4372,N_3373);
nand U5241 (N_5241,N_3926,N_3093);
nand U5242 (N_5242,N_2668,N_3856);
nand U5243 (N_5243,N_4741,N_4631);
or U5244 (N_5244,N_3901,N_2691);
nor U5245 (N_5245,N_4657,N_2546);
nand U5246 (N_5246,N_4127,N_2513);
or U5247 (N_5247,N_3907,N_3872);
or U5248 (N_5248,N_4150,N_4999);
or U5249 (N_5249,N_3525,N_4386);
xor U5250 (N_5250,N_3580,N_2839);
nand U5251 (N_5251,N_3975,N_2633);
nand U5252 (N_5252,N_3646,N_3532);
and U5253 (N_5253,N_4479,N_3425);
nand U5254 (N_5254,N_4776,N_4188);
or U5255 (N_5255,N_3121,N_4662);
nor U5256 (N_5256,N_4745,N_2976);
or U5257 (N_5257,N_3077,N_3598);
xor U5258 (N_5258,N_3533,N_4038);
or U5259 (N_5259,N_3810,N_3116);
nand U5260 (N_5260,N_2897,N_2821);
and U5261 (N_5261,N_4237,N_4510);
nand U5262 (N_5262,N_4068,N_3246);
and U5263 (N_5263,N_2713,N_2795);
nand U5264 (N_5264,N_4857,N_3814);
xor U5265 (N_5265,N_4049,N_3278);
xnor U5266 (N_5266,N_3995,N_4739);
nor U5267 (N_5267,N_2984,N_4383);
nor U5268 (N_5268,N_3467,N_4285);
nor U5269 (N_5269,N_3659,N_4720);
nand U5270 (N_5270,N_2650,N_4676);
nand U5271 (N_5271,N_3739,N_3248);
and U5272 (N_5272,N_3277,N_4072);
nor U5273 (N_5273,N_3252,N_4957);
nor U5274 (N_5274,N_3329,N_3102);
or U5275 (N_5275,N_3845,N_4852);
nor U5276 (N_5276,N_2937,N_2905);
nand U5277 (N_5277,N_4458,N_2954);
xnor U5278 (N_5278,N_4169,N_3403);
and U5279 (N_5279,N_2987,N_4257);
nor U5280 (N_5280,N_4724,N_4874);
nand U5281 (N_5281,N_4630,N_4514);
or U5282 (N_5282,N_4210,N_3893);
nor U5283 (N_5283,N_3075,N_4153);
nor U5284 (N_5284,N_2578,N_3722);
nand U5285 (N_5285,N_4218,N_3732);
xnor U5286 (N_5286,N_3044,N_2636);
and U5287 (N_5287,N_4829,N_3549);
or U5288 (N_5288,N_4574,N_3761);
nor U5289 (N_5289,N_4673,N_4848);
nand U5290 (N_5290,N_3217,N_4325);
nand U5291 (N_5291,N_4473,N_2623);
or U5292 (N_5292,N_3029,N_4853);
xnor U5293 (N_5293,N_3144,N_4743);
nand U5294 (N_5294,N_3877,N_4014);
xor U5295 (N_5295,N_3677,N_3531);
nor U5296 (N_5296,N_2956,N_3018);
nand U5297 (N_5297,N_2761,N_4996);
nor U5298 (N_5298,N_4492,N_4626);
xnor U5299 (N_5299,N_3633,N_3159);
or U5300 (N_5300,N_3508,N_4634);
and U5301 (N_5301,N_4591,N_4958);
and U5302 (N_5302,N_4040,N_4597);
nor U5303 (N_5303,N_3233,N_2844);
nand U5304 (N_5304,N_3424,N_3294);
and U5305 (N_5305,N_4836,N_3343);
nand U5306 (N_5306,N_3235,N_2587);
nor U5307 (N_5307,N_3956,N_3691);
nand U5308 (N_5308,N_2516,N_4821);
and U5309 (N_5309,N_4165,N_4435);
or U5310 (N_5310,N_3912,N_4909);
and U5311 (N_5311,N_2667,N_3041);
nand U5312 (N_5312,N_3692,N_3784);
nand U5313 (N_5313,N_3156,N_4444);
nand U5314 (N_5314,N_3164,N_4546);
nand U5315 (N_5315,N_4493,N_2505);
nand U5316 (N_5316,N_3316,N_2619);
nor U5317 (N_5317,N_3154,N_3683);
or U5318 (N_5318,N_4376,N_2922);
and U5319 (N_5319,N_4628,N_4519);
nor U5320 (N_5320,N_4894,N_2624);
or U5321 (N_5321,N_4581,N_2929);
nand U5322 (N_5322,N_3619,N_3599);
or U5323 (N_5323,N_3196,N_3918);
and U5324 (N_5324,N_4031,N_3391);
or U5325 (N_5325,N_3954,N_3131);
xnor U5326 (N_5326,N_2768,N_2873);
or U5327 (N_5327,N_3153,N_4001);
nand U5328 (N_5328,N_3152,N_3165);
or U5329 (N_5329,N_3937,N_4918);
and U5330 (N_5330,N_4587,N_3017);
or U5331 (N_5331,N_3831,N_4058);
nand U5332 (N_5332,N_3142,N_4934);
xor U5333 (N_5333,N_3504,N_2600);
and U5334 (N_5334,N_3870,N_2593);
nand U5335 (N_5335,N_2610,N_4677);
or U5336 (N_5336,N_3778,N_3056);
nor U5337 (N_5337,N_4353,N_4684);
nand U5338 (N_5338,N_2703,N_3305);
nand U5339 (N_5339,N_2676,N_4968);
or U5340 (N_5340,N_4978,N_3001);
or U5341 (N_5341,N_3944,N_3940);
or U5342 (N_5342,N_2672,N_2891);
nor U5343 (N_5343,N_4088,N_4318);
nor U5344 (N_5344,N_3647,N_3335);
nand U5345 (N_5345,N_3881,N_4100);
and U5346 (N_5346,N_3483,N_4243);
nand U5347 (N_5347,N_2679,N_2888);
xor U5348 (N_5348,N_4246,N_3108);
nor U5349 (N_5349,N_4219,N_2934);
xnor U5350 (N_5350,N_4486,N_4871);
nand U5351 (N_5351,N_3369,N_2807);
or U5352 (N_5352,N_4085,N_4487);
nor U5353 (N_5353,N_4650,N_3114);
nand U5354 (N_5354,N_4398,N_2991);
nand U5355 (N_5355,N_3349,N_3241);
or U5356 (N_5356,N_3770,N_4540);
and U5357 (N_5357,N_4560,N_4471);
and U5358 (N_5358,N_4255,N_3388);
xor U5359 (N_5359,N_3726,N_3667);
nor U5360 (N_5360,N_4439,N_2762);
and U5361 (N_5361,N_4599,N_4949);
nand U5362 (N_5362,N_3439,N_4780);
xnor U5363 (N_5363,N_4930,N_3971);
nor U5364 (N_5364,N_2886,N_4746);
nand U5365 (N_5365,N_2948,N_3417);
and U5366 (N_5366,N_4618,N_2927);
xnor U5367 (N_5367,N_3109,N_4499);
and U5368 (N_5368,N_4196,N_2889);
or U5369 (N_5369,N_3341,N_2656);
and U5370 (N_5370,N_4686,N_4212);
and U5371 (N_5371,N_4078,N_4341);
or U5372 (N_5372,N_3348,N_2654);
xor U5373 (N_5373,N_3451,N_3119);
and U5374 (N_5374,N_3190,N_3909);
and U5375 (N_5375,N_3575,N_3428);
xnor U5376 (N_5376,N_4734,N_4834);
nor U5377 (N_5377,N_3564,N_3758);
nor U5378 (N_5378,N_2830,N_4947);
or U5379 (N_5379,N_3128,N_3895);
nor U5380 (N_5380,N_4615,N_3731);
and U5381 (N_5381,N_4060,N_4263);
or U5382 (N_5382,N_3650,N_3671);
and U5383 (N_5383,N_2800,N_2701);
nand U5384 (N_5384,N_3195,N_4338);
and U5385 (N_5385,N_2582,N_4737);
nor U5386 (N_5386,N_4988,N_4873);
nor U5387 (N_5387,N_3557,N_2799);
and U5388 (N_5388,N_3517,N_3518);
nand U5389 (N_5389,N_2618,N_3570);
and U5390 (N_5390,N_4671,N_4077);
nor U5391 (N_5391,N_3812,N_4954);
xor U5392 (N_5392,N_4421,N_4125);
nor U5393 (N_5393,N_2729,N_3768);
nor U5394 (N_5394,N_3801,N_4467);
xor U5395 (N_5395,N_4523,N_3016);
xor U5396 (N_5396,N_4785,N_3587);
and U5397 (N_5397,N_3088,N_3892);
nand U5398 (N_5398,N_3796,N_3919);
nand U5399 (N_5399,N_4980,N_4174);
nand U5400 (N_5400,N_3127,N_2673);
nand U5401 (N_5401,N_3631,N_3766);
and U5402 (N_5402,N_2865,N_2627);
and U5403 (N_5403,N_3311,N_3586);
and U5404 (N_5404,N_3049,N_4164);
or U5405 (N_5405,N_3850,N_4402);
nand U5406 (N_5406,N_3748,N_4238);
xor U5407 (N_5407,N_4594,N_2564);
or U5408 (N_5408,N_4705,N_2565);
nor U5409 (N_5409,N_4695,N_3835);
nor U5410 (N_5410,N_3496,N_2907);
nor U5411 (N_5411,N_3224,N_3964);
and U5412 (N_5412,N_2520,N_4016);
or U5413 (N_5413,N_4424,N_3027);
xnor U5414 (N_5414,N_4927,N_4887);
nand U5415 (N_5415,N_2548,N_4967);
or U5416 (N_5416,N_3457,N_3446);
or U5417 (N_5417,N_4239,N_3973);
nor U5418 (N_5418,N_4639,N_4866);
and U5419 (N_5419,N_4043,N_4299);
or U5420 (N_5420,N_3280,N_4106);
or U5421 (N_5421,N_2805,N_4450);
and U5422 (N_5422,N_3803,N_3392);
xnor U5423 (N_5423,N_4466,N_3218);
xor U5424 (N_5424,N_3524,N_3889);
and U5425 (N_5425,N_4382,N_3632);
or U5426 (N_5426,N_2992,N_4441);
nor U5427 (N_5427,N_3769,N_3509);
nor U5428 (N_5428,N_2751,N_2542);
and U5429 (N_5429,N_2784,N_4074);
nand U5430 (N_5430,N_2525,N_3427);
xor U5431 (N_5431,N_4815,N_3503);
and U5432 (N_5432,N_3053,N_3288);
nor U5433 (N_5433,N_3071,N_4635);
nor U5434 (N_5434,N_2871,N_2748);
nor U5435 (N_5435,N_4687,N_3999);
and U5436 (N_5436,N_3897,N_4132);
or U5437 (N_5437,N_2872,N_4917);
xor U5438 (N_5438,N_2826,N_4698);
nand U5439 (N_5439,N_2659,N_4418);
nor U5440 (N_5440,N_2953,N_4661);
nand U5441 (N_5441,N_4998,N_3257);
nand U5442 (N_5442,N_3984,N_4199);
or U5443 (N_5443,N_2621,N_4969);
and U5444 (N_5444,N_3962,N_2859);
or U5445 (N_5445,N_2614,N_3811);
nand U5446 (N_5446,N_4475,N_3841);
nor U5447 (N_5447,N_3797,N_4093);
xnor U5448 (N_5448,N_3148,N_4707);
or U5449 (N_5449,N_3299,N_3404);
or U5450 (N_5450,N_3371,N_3182);
and U5451 (N_5451,N_2921,N_4536);
nor U5452 (N_5452,N_4323,N_3642);
nor U5453 (N_5453,N_4962,N_3420);
xnor U5454 (N_5454,N_4789,N_3465);
xor U5455 (N_5455,N_2919,N_3094);
nand U5456 (N_5456,N_3012,N_4087);
nand U5457 (N_5457,N_3578,N_4137);
and U5458 (N_5458,N_4886,N_3201);
or U5459 (N_5459,N_4090,N_4678);
xnor U5460 (N_5460,N_3621,N_2887);
or U5461 (N_5461,N_3191,N_3304);
or U5462 (N_5462,N_3231,N_3125);
or U5463 (N_5463,N_4710,N_2834);
or U5464 (N_5464,N_3925,N_2812);
xor U5465 (N_5465,N_4966,N_2950);
or U5466 (N_5466,N_3763,N_4474);
and U5467 (N_5467,N_2977,N_3558);
xor U5468 (N_5468,N_2951,N_3965);
or U5469 (N_5469,N_2752,N_3522);
nor U5470 (N_5470,N_4575,N_3639);
nand U5471 (N_5471,N_2778,N_3935);
xnor U5472 (N_5472,N_3551,N_3287);
xnor U5473 (N_5473,N_4665,N_3205);
nor U5474 (N_5474,N_3471,N_4480);
nand U5475 (N_5475,N_4177,N_3161);
xor U5476 (N_5476,N_4613,N_4013);
or U5477 (N_5477,N_4736,N_3172);
xor U5478 (N_5478,N_3584,N_3040);
nor U5479 (N_5479,N_2998,N_2620);
or U5480 (N_5480,N_3354,N_2775);
nor U5481 (N_5481,N_2588,N_4082);
nor U5482 (N_5482,N_4477,N_3932);
nor U5483 (N_5483,N_3651,N_2724);
nor U5484 (N_5484,N_2958,N_3721);
xnor U5485 (N_5485,N_4766,N_4620);
and U5486 (N_5486,N_3661,N_4426);
nor U5487 (N_5487,N_4778,N_3492);
or U5488 (N_5488,N_4226,N_3802);
nand U5489 (N_5489,N_2747,N_3338);
or U5490 (N_5490,N_3673,N_3535);
nor U5491 (N_5491,N_4701,N_3577);
or U5492 (N_5492,N_4184,N_4876);
nor U5493 (N_5493,N_2766,N_3556);
nor U5494 (N_5494,N_4761,N_4233);
or U5495 (N_5495,N_2803,N_4945);
or U5496 (N_5496,N_3607,N_2661);
nor U5497 (N_5497,N_4079,N_2995);
xor U5498 (N_5498,N_4982,N_4309);
or U5499 (N_5499,N_4539,N_3711);
nor U5500 (N_5500,N_3261,N_4339);
nand U5501 (N_5501,N_4344,N_3753);
and U5502 (N_5502,N_3640,N_4910);
nand U5503 (N_5503,N_3561,N_3134);
nor U5504 (N_5504,N_4956,N_2715);
or U5505 (N_5505,N_2943,N_2732);
nand U5506 (N_5506,N_4882,N_3777);
or U5507 (N_5507,N_4777,N_4220);
nor U5508 (N_5508,N_4207,N_2563);
nand U5509 (N_5509,N_4841,N_4315);
nand U5510 (N_5510,N_2605,N_3076);
xnor U5511 (N_5511,N_2915,N_4845);
nand U5512 (N_5512,N_4534,N_3955);
nor U5513 (N_5513,N_2754,N_4679);
xnor U5514 (N_5514,N_3934,N_2704);
nand U5515 (N_5515,N_2813,N_3068);
and U5516 (N_5516,N_2794,N_4494);
and U5517 (N_5517,N_4515,N_3297);
and U5518 (N_5518,N_3818,N_3291);
nor U5519 (N_5519,N_4951,N_4026);
nor U5520 (N_5520,N_4029,N_3808);
and U5521 (N_5521,N_4926,N_3963);
nand U5522 (N_5522,N_4649,N_4807);
nand U5523 (N_5523,N_2721,N_3066);
or U5524 (N_5524,N_4897,N_3072);
or U5525 (N_5525,N_3318,N_3401);
nand U5526 (N_5526,N_3519,N_4230);
nor U5527 (N_5527,N_3323,N_2745);
and U5528 (N_5528,N_2940,N_4394);
nand U5529 (N_5529,N_4267,N_3813);
xnor U5530 (N_5530,N_2845,N_2700);
or U5531 (N_5531,N_2581,N_4136);
and U5532 (N_5532,N_3652,N_3741);
xor U5533 (N_5533,N_4279,N_2682);
and U5534 (N_5534,N_3171,N_2926);
or U5535 (N_5535,N_3550,N_4728);
or U5536 (N_5536,N_2734,N_3585);
nand U5537 (N_5537,N_3537,N_3698);
nand U5538 (N_5538,N_3900,N_2764);
or U5539 (N_5539,N_3685,N_3206);
nand U5540 (N_5540,N_4938,N_3649);
or U5541 (N_5541,N_4357,N_2670);
and U5542 (N_5542,N_2823,N_3807);
or U5543 (N_5543,N_2738,N_4354);
or U5544 (N_5544,N_2750,N_4044);
nor U5545 (N_5545,N_4572,N_3705);
and U5546 (N_5546,N_3055,N_3100);
or U5547 (N_5547,N_2728,N_3175);
nor U5548 (N_5548,N_4097,N_4120);
xnor U5549 (N_5549,N_3764,N_4647);
nand U5550 (N_5550,N_4369,N_3755);
or U5551 (N_5551,N_2696,N_4993);
nor U5552 (N_5552,N_4225,N_3303);
nand U5553 (N_5553,N_3756,N_4241);
nand U5554 (N_5554,N_3710,N_4855);
nor U5555 (N_5555,N_2957,N_4343);
or U5556 (N_5556,N_3208,N_3752);
nand U5557 (N_5557,N_4818,N_3875);
xnor U5558 (N_5558,N_4823,N_4683);
or U5559 (N_5559,N_4692,N_4195);
or U5560 (N_5560,N_4222,N_3992);
or U5561 (N_5561,N_3905,N_4933);
or U5562 (N_5562,N_3223,N_3099);
or U5563 (N_5563,N_4502,N_3419);
xnor U5564 (N_5564,N_4907,N_3696);
nor U5565 (N_5565,N_3635,N_4787);
and U5566 (N_5566,N_2602,N_4094);
or U5567 (N_5567,N_4149,N_2743);
or U5568 (N_5568,N_4391,N_4645);
nor U5569 (N_5569,N_4612,N_2543);
nand U5570 (N_5570,N_4065,N_3629);
xor U5571 (N_5571,N_2916,N_4825);
and U5572 (N_5572,N_4425,N_4719);
and U5573 (N_5573,N_2692,N_2963);
or U5574 (N_5574,N_4448,N_4172);
or U5575 (N_5575,N_3703,N_4742);
nor U5576 (N_5576,N_2853,N_4071);
nor U5577 (N_5577,N_3267,N_4242);
and U5578 (N_5578,N_2796,N_2802);
nand U5579 (N_5579,N_3350,N_4066);
or U5580 (N_5580,N_3289,N_2645);
or U5581 (N_5581,N_4644,N_3330);
nor U5582 (N_5582,N_3902,N_3282);
nor U5583 (N_5583,N_2837,N_3961);
and U5584 (N_5584,N_2688,N_4443);
xor U5585 (N_5585,N_4168,N_4989);
nand U5586 (N_5586,N_4224,N_2994);
nor U5587 (N_5587,N_2733,N_4397);
and U5588 (N_5588,N_4532,N_3293);
nand U5589 (N_5589,N_2567,N_2983);
or U5590 (N_5590,N_4627,N_4240);
nand U5591 (N_5591,N_4654,N_3151);
or U5592 (N_5592,N_4880,N_3911);
nand U5593 (N_5593,N_4784,N_3443);
and U5594 (N_5594,N_3034,N_3849);
nand U5595 (N_5595,N_4370,N_4763);
or U5596 (N_5596,N_4260,N_3253);
or U5597 (N_5597,N_4531,N_4408);
nor U5598 (N_5598,N_3521,N_2858);
nand U5599 (N_5599,N_4740,N_3552);
nand U5600 (N_5600,N_4140,N_2849);
xnor U5601 (N_5601,N_4459,N_2925);
nand U5602 (N_5602,N_3122,N_4105);
or U5603 (N_5603,N_3981,N_2695);
or U5604 (N_5604,N_4131,N_4216);
and U5605 (N_5605,N_4624,N_4875);
or U5606 (N_5606,N_4508,N_4108);
or U5607 (N_5607,N_4826,N_3644);
xnor U5608 (N_5608,N_3626,N_4593);
or U5609 (N_5609,N_3445,N_3396);
and U5610 (N_5610,N_3433,N_3236);
or U5611 (N_5611,N_2544,N_3340);
or U5612 (N_5612,N_4170,N_2810);
or U5613 (N_5613,N_3861,N_4971);
or U5614 (N_5614,N_4582,N_3003);
xnor U5615 (N_5615,N_3951,N_4896);
nand U5616 (N_5616,N_4833,N_3285);
nor U5617 (N_5617,N_3177,N_4653);
nor U5618 (N_5618,N_3339,N_3167);
or U5619 (N_5619,N_3232,N_3855);
or U5620 (N_5620,N_4929,N_3526);
or U5621 (N_5621,N_4902,N_3059);
and U5622 (N_5622,N_4250,N_2758);
and U5623 (N_5623,N_4128,N_2892);
or U5624 (N_5624,N_3468,N_3418);
xnor U5625 (N_5625,N_3019,N_3545);
and U5626 (N_5626,N_3336,N_3591);
and U5627 (N_5627,N_4249,N_3678);
or U5628 (N_5628,N_4544,N_2819);
nand U5629 (N_5629,N_3050,N_4943);
or U5630 (N_5630,N_2531,N_4718);
or U5631 (N_5631,N_3735,N_3953);
nor U5632 (N_5632,N_3945,N_3670);
and U5633 (N_5633,N_4670,N_2690);
nand U5634 (N_5634,N_4573,N_3309);
and U5635 (N_5635,N_2694,N_2861);
and U5636 (N_5636,N_3747,N_3783);
nand U5637 (N_5637,N_4095,N_3746);
or U5638 (N_5638,N_3455,N_4550);
or U5639 (N_5639,N_3188,N_3098);
nor U5640 (N_5640,N_4312,N_3576);
nand U5641 (N_5641,N_3760,N_3269);
nand U5642 (N_5642,N_3506,N_3166);
nand U5643 (N_5643,N_3024,N_2866);
nand U5644 (N_5644,N_3505,N_3222);
and U5645 (N_5645,N_4447,N_3542);
nor U5646 (N_5646,N_3516,N_3456);
and U5647 (N_5647,N_3538,N_4297);
and U5648 (N_5648,N_4584,N_3194);
nand U5649 (N_5649,N_2504,N_3308);
or U5650 (N_5650,N_3840,N_4032);
xor U5651 (N_5651,N_3713,N_3062);
or U5652 (N_5652,N_4023,N_3022);
or U5653 (N_5653,N_4410,N_3804);
nand U5654 (N_5654,N_2642,N_4422);
nor U5655 (N_5655,N_4463,N_3169);
xor U5656 (N_5656,N_4940,N_3654);
and U5657 (N_5657,N_4696,N_4067);
nand U5658 (N_5658,N_3170,N_2612);
and U5659 (N_5659,N_3273,N_2767);
xnor U5660 (N_5660,N_3104,N_4133);
or U5661 (N_5661,N_3090,N_2855);
nor U5662 (N_5662,N_4143,N_3402);
or U5663 (N_5663,N_3637,N_4256);
and U5664 (N_5664,N_3069,N_4555);
or U5665 (N_5665,N_4221,N_3583);
and U5666 (N_5666,N_3574,N_2787);
nor U5667 (N_5667,N_4646,N_3460);
nand U5668 (N_5668,N_4495,N_4704);
nand U5669 (N_5669,N_2669,N_2637);
xor U5670 (N_5670,N_4611,N_2683);
nor U5671 (N_5671,N_3816,N_4912);
nor U5672 (N_5672,N_3000,N_2574);
nor U5673 (N_5673,N_4349,N_3544);
and U5674 (N_5674,N_4380,N_3704);
nor U5675 (N_5675,N_4528,N_4602);
and U5676 (N_5676,N_2575,N_3967);
or U5677 (N_5677,N_4537,N_2899);
and U5678 (N_5678,N_3743,N_3790);
and U5679 (N_5679,N_2566,N_4336);
and U5680 (N_5680,N_2607,N_4180);
nand U5681 (N_5681,N_4827,N_3794);
nand U5682 (N_5682,N_3957,N_3686);
or U5683 (N_5683,N_3847,N_4371);
nor U5684 (N_5684,N_4186,N_4846);
or U5685 (N_5685,N_4183,N_2843);
nor U5686 (N_5686,N_3357,N_2774);
and U5687 (N_5687,N_2658,N_3260);
and U5688 (N_5688,N_3060,N_4759);
or U5689 (N_5689,N_4490,N_2519);
or U5690 (N_5690,N_4176,N_4171);
nand U5691 (N_5691,N_3087,N_2533);
or U5692 (N_5692,N_4053,N_2685);
nor U5693 (N_5693,N_3078,N_3573);
or U5694 (N_5694,N_3244,N_4619);
and U5695 (N_5695,N_3033,N_3716);
nor U5696 (N_5696,N_3884,N_4535);
and U5697 (N_5697,N_3879,N_3234);
nor U5698 (N_5698,N_2836,N_3543);
nand U5699 (N_5699,N_4144,N_4792);
xnor U5700 (N_5700,N_2643,N_2549);
xor U5701 (N_5701,N_4275,N_4788);
and U5702 (N_5702,N_2938,N_3628);
xor U5703 (N_5703,N_2974,N_3219);
xnor U5704 (N_5704,N_3643,N_3826);
nand U5705 (N_5705,N_4725,N_4301);
nor U5706 (N_5706,N_3689,N_3488);
nand U5707 (N_5707,N_3493,N_4932);
nand U5708 (N_5708,N_3276,N_3958);
and U5709 (N_5709,N_3828,N_4990);
nand U5710 (N_5710,N_3249,N_4674);
and U5711 (N_5711,N_3908,N_3270);
nand U5712 (N_5712,N_3426,N_4191);
and U5713 (N_5713,N_3387,N_3725);
and U5714 (N_5714,N_4449,N_2955);
nor U5715 (N_5715,N_2961,N_4570);
xnor U5716 (N_5716,N_3680,N_3009);
xor U5717 (N_5717,N_4900,N_3982);
nor U5718 (N_5718,N_3328,N_4881);
nand U5719 (N_5719,N_4166,N_4901);
nor U5720 (N_5720,N_4824,N_2530);
or U5721 (N_5721,N_4414,N_3284);
or U5722 (N_5722,N_4181,N_3702);
nand U5723 (N_5723,N_3809,N_4070);
nand U5724 (N_5724,N_4811,N_4889);
and U5725 (N_5725,N_3061,N_2655);
xor U5726 (N_5726,N_4340,N_3501);
and U5727 (N_5727,N_3727,N_3315);
nand U5728 (N_5728,N_2890,N_4955);
nand U5729 (N_5729,N_3023,N_3898);
nand U5730 (N_5730,N_2631,N_4245);
or U5731 (N_5731,N_3658,N_4147);
nand U5732 (N_5732,N_4817,N_4850);
or U5733 (N_5733,N_2601,N_4682);
xnor U5734 (N_5734,N_4022,N_2594);
nand U5735 (N_5735,N_3085,N_3740);
xnor U5736 (N_5736,N_3450,N_3612);
and U5737 (N_5737,N_3681,N_3679);
nor U5738 (N_5738,N_4605,N_4754);
nor U5739 (N_5739,N_3606,N_4355);
or U5740 (N_5740,N_4774,N_2898);
or U5741 (N_5741,N_4277,N_2677);
nand U5742 (N_5742,N_2608,N_3891);
and U5743 (N_5743,N_3969,N_4020);
nor U5744 (N_5744,N_4055,N_4545);
and U5745 (N_5745,N_4121,N_4606);
nor U5746 (N_5746,N_2971,N_4298);
nand U5747 (N_5747,N_3634,N_2882);
nor U5748 (N_5748,N_4375,N_2576);
and U5749 (N_5749,N_3243,N_4112);
or U5750 (N_5750,N_3454,N_4542);
xor U5751 (N_5751,N_3858,N_4800);
nor U5752 (N_5752,N_2562,N_3367);
and U5753 (N_5753,N_4231,N_4935);
nand U5754 (N_5754,N_4206,N_3994);
or U5755 (N_5755,N_4135,N_3988);
or U5756 (N_5756,N_4831,N_3559);
and U5757 (N_5757,N_3324,N_4623);
nand U5758 (N_5758,N_4395,N_3792);
nor U5759 (N_5759,N_3980,N_2876);
nor U5760 (N_5760,N_4440,N_4566);
and U5761 (N_5761,N_2908,N_2797);
and U5762 (N_5762,N_3203,N_4007);
or U5763 (N_5763,N_4114,N_4314);
nor U5764 (N_5764,N_3378,N_4805);
nor U5765 (N_5765,N_3915,N_2964);
or U5766 (N_5766,N_4209,N_3568);
nor U5767 (N_5767,N_2952,N_4050);
nand U5768 (N_5768,N_4278,N_2920);
xor U5769 (N_5769,N_2928,N_3890);
and U5770 (N_5770,N_2792,N_4189);
or U5771 (N_5771,N_3389,N_3386);
and U5772 (N_5772,N_2719,N_3883);
nor U5773 (N_5773,N_3950,N_2895);
xor U5774 (N_5774,N_3541,N_3602);
or U5775 (N_5775,N_2801,N_3922);
or U5776 (N_5776,N_2629,N_4861);
and U5777 (N_5777,N_4304,N_3133);
and U5778 (N_5778,N_3112,N_3865);
nand U5779 (N_5779,N_4104,N_4961);
nand U5780 (N_5780,N_4816,N_3408);
or U5781 (N_5781,N_3176,N_4005);
and U5782 (N_5782,N_2880,N_4664);
nand U5783 (N_5783,N_4485,N_4110);
xnor U5784 (N_5784,N_3296,N_3149);
and U5785 (N_5785,N_3666,N_4658);
nand U5786 (N_5786,N_4870,N_4937);
nor U5787 (N_5787,N_2863,N_4697);
or U5788 (N_5788,N_3032,N_4756);
or U5789 (N_5789,N_2702,N_4702);
or U5790 (N_5790,N_3539,N_4142);
nand U5791 (N_5791,N_3491,N_2884);
nand U5792 (N_5792,N_3939,N_4423);
nor U5793 (N_5793,N_3611,N_4505);
nand U5794 (N_5794,N_4454,N_4772);
nand U5795 (N_5795,N_3510,N_4155);
nand U5796 (N_5796,N_4548,N_4888);
xnor U5797 (N_5797,N_3413,N_3412);
or U5798 (N_5798,N_4694,N_3668);
and U5799 (N_5799,N_2634,N_4358);
nand U5800 (N_5800,N_4964,N_3569);
nand U5801 (N_5801,N_3896,N_3754);
and U5802 (N_5802,N_2737,N_4750);
and U5803 (N_5803,N_3111,N_4793);
and U5804 (N_5804,N_4086,N_4979);
and U5805 (N_5805,N_3047,N_3478);
or U5806 (N_5806,N_2611,N_4571);
and U5807 (N_5807,N_3793,N_4235);
nor U5808 (N_5808,N_4783,N_4590);
nand U5809 (N_5809,N_3334,N_3821);
or U5810 (N_5810,N_2558,N_4965);
and U5811 (N_5811,N_4723,N_4781);
or U5812 (N_5812,N_3985,N_2962);
nand U5813 (N_5813,N_2941,N_4600);
nor U5814 (N_5814,N_4809,N_3990);
nor U5815 (N_5815,N_2720,N_3130);
nor U5816 (N_5816,N_3852,N_3139);
xor U5817 (N_5817,N_3251,N_2901);
nor U5818 (N_5818,N_4288,N_4252);
nand U5819 (N_5819,N_2793,N_4236);
and U5820 (N_5820,N_3214,N_3459);
nor U5821 (N_5821,N_3782,N_4614);
or U5822 (N_5822,N_3405,N_4812);
nor U5823 (N_5823,N_3472,N_4509);
and U5824 (N_5824,N_4379,N_3372);
or U5825 (N_5825,N_4381,N_3435);
nand U5826 (N_5826,N_4399,N_3083);
or U5827 (N_5827,N_4752,N_3603);
and U5828 (N_5828,N_3259,N_3434);
or U5829 (N_5829,N_3342,N_4442);
and U5830 (N_5830,N_3238,N_2820);
and U5831 (N_5831,N_3207,N_2541);
and U5832 (N_5832,N_4462,N_3688);
and U5833 (N_5833,N_3949,N_3440);
nor U5834 (N_5834,N_3904,N_4415);
nand U5835 (N_5835,N_2710,N_3540);
nand U5836 (N_5836,N_2832,N_3337);
nor U5837 (N_5837,N_3989,N_3042);
or U5838 (N_5838,N_2502,N_3978);
nand U5839 (N_5839,N_3714,N_4091);
nor U5840 (N_5840,N_3301,N_3885);
nor U5841 (N_5841,N_4280,N_2686);
nor U5842 (N_5842,N_4069,N_2662);
nand U5843 (N_5843,N_3117,N_3163);
nor U5844 (N_5844,N_4214,N_3422);
or U5845 (N_5845,N_3162,N_2997);
and U5846 (N_5846,N_4558,N_3833);
nand U5847 (N_5847,N_4310,N_4974);
and U5848 (N_5848,N_4073,N_4478);
or U5849 (N_5849,N_2512,N_2515);
or U5850 (N_5850,N_3474,N_3486);
nor U5851 (N_5851,N_3563,N_4436);
or U5852 (N_5852,N_3250,N_4363);
or U5853 (N_5853,N_4404,N_3837);
xor U5854 (N_5854,N_2613,N_3931);
nand U5855 (N_5855,N_3264,N_4187);
and U5856 (N_5856,N_2975,N_2625);
and U5857 (N_5857,N_3447,N_4794);
nor U5858 (N_5858,N_3830,N_4019);
nor U5859 (N_5859,N_3863,N_4033);
nor U5860 (N_5860,N_4089,N_4360);
and U5861 (N_5861,N_4621,N_4796);
nor U5862 (N_5862,N_3407,N_4460);
nand U5863 (N_5863,N_3310,N_4865);
and U5864 (N_5864,N_2765,N_4830);
and U5865 (N_5865,N_4009,N_3008);
xnor U5866 (N_5866,N_4098,N_4563);
or U5867 (N_5867,N_3105,N_4729);
xnor U5868 (N_5868,N_4308,N_4541);
and U5869 (N_5869,N_2759,N_3215);
and U5870 (N_5870,N_4885,N_4877);
nand U5871 (N_5871,N_4334,N_3063);
nor U5872 (N_5872,N_3672,N_3927);
or U5873 (N_5873,N_3120,N_3397);
nor U5874 (N_5874,N_3110,N_4234);
or U5875 (N_5875,N_4406,N_2840);
nand U5876 (N_5876,N_3258,N_3693);
and U5877 (N_5877,N_3878,N_4711);
xor U5878 (N_5878,N_3657,N_4498);
or U5879 (N_5879,N_4775,N_3806);
xor U5880 (N_5880,N_4160,N_3820);
nor U5881 (N_5881,N_4322,N_2896);
or U5882 (N_5882,N_4024,N_3882);
nand U5883 (N_5883,N_4457,N_2885);
nand U5884 (N_5884,N_4849,N_4203);
nor U5885 (N_5885,N_3554,N_4884);
and U5886 (N_5886,N_4420,N_4476);
or U5887 (N_5887,N_3624,N_4247);
xnor U5888 (N_5888,N_4651,N_4655);
nor U5889 (N_5889,N_4326,N_2769);
nor U5890 (N_5890,N_4749,N_3379);
nor U5891 (N_5891,N_2596,N_4906);
xor U5892 (N_5892,N_3321,N_4292);
and U5893 (N_5893,N_2986,N_2687);
and U5894 (N_5894,N_4413,N_3004);
nand U5895 (N_5895,N_3430,N_4258);
and U5896 (N_5896,N_2999,N_3687);
nor U5897 (N_5897,N_3996,N_4152);
nor U5898 (N_5898,N_3997,N_3344);
and U5899 (N_5899,N_3617,N_2550);
nor U5900 (N_5900,N_4629,N_3381);
nand U5901 (N_5901,N_2817,N_3263);
nor U5902 (N_5902,N_2877,N_4976);
or U5903 (N_5903,N_4008,N_4913);
nor U5904 (N_5904,N_3126,N_4197);
nor U5905 (N_5905,N_3074,N_4714);
xnor U5906 (N_5906,N_2707,N_3917);
nor U5907 (N_5907,N_4264,N_4801);
nand U5908 (N_5908,N_4345,N_4656);
and U5909 (N_5909,N_4116,N_3655);
and U5910 (N_5910,N_4770,N_4762);
nand U5911 (N_5911,N_4819,N_4928);
and U5912 (N_5912,N_4359,N_4200);
nand U5913 (N_5913,N_3365,N_2829);
nor U5914 (N_5914,N_3597,N_4842);
nor U5915 (N_5915,N_3255,N_4101);
nor U5916 (N_5916,N_2521,N_2912);
or U5917 (N_5917,N_2615,N_3302);
or U5918 (N_5918,N_2900,N_4190);
nor U5919 (N_5919,N_4942,N_3610);
nor U5920 (N_5920,N_3096,N_3140);
nand U5921 (N_5921,N_3370,N_3933);
nand U5922 (N_5922,N_2554,N_4284);
nand U5923 (N_5923,N_3307,N_3844);
nand U5924 (N_5924,N_3536,N_3274);
nand U5925 (N_5925,N_4844,N_3827);
nand U5926 (N_5926,N_4804,N_3481);
and U5927 (N_5927,N_3795,N_4400);
and U5928 (N_5928,N_3184,N_3256);
nand U5929 (N_5929,N_4732,N_2854);
nand U5930 (N_5930,N_4893,N_3757);
and U5931 (N_5931,N_3485,N_4923);
nor U5932 (N_5932,N_3415,N_4522);
or U5933 (N_5933,N_3708,N_4052);
or U5934 (N_5934,N_2698,N_4981);
nand U5935 (N_5935,N_4348,N_4179);
xnor U5936 (N_5936,N_4521,N_3527);
and U5937 (N_5937,N_2560,N_3476);
nor U5938 (N_5938,N_4828,N_2555);
and U5939 (N_5939,N_3929,N_2523);
and U5940 (N_5940,N_4059,N_3674);
or U5941 (N_5941,N_4405,N_2604);
and U5942 (N_5942,N_4972,N_2822);
and U5943 (N_5943,N_3616,N_4373);
or U5944 (N_5944,N_3738,N_4167);
or U5945 (N_5945,N_3410,N_2689);
and U5946 (N_5946,N_2942,N_3313);
or U5947 (N_5947,N_3592,N_4350);
nand U5948 (N_5948,N_3080,N_3737);
nor U5949 (N_5949,N_4731,N_4201);
or U5950 (N_5950,N_2911,N_3839);
nand U5951 (N_5951,N_3158,N_3530);
and U5952 (N_5952,N_4564,N_4387);
or U5953 (N_5953,N_3625,N_4672);
and U5954 (N_5954,N_3512,N_4632);
nand U5955 (N_5955,N_3641,N_2592);
or U5956 (N_5956,N_2815,N_2503);
and U5957 (N_5957,N_2763,N_4254);
and U5958 (N_5958,N_4518,N_4963);
nand U5959 (N_5959,N_4037,N_3562);
and U5960 (N_5960,N_4446,N_4139);
or U5961 (N_5961,N_4465,N_4324);
or U5962 (N_5962,N_2968,N_2644);
or U5963 (N_5963,N_4080,N_3265);
and U5964 (N_5964,N_3773,N_4028);
and U5965 (N_5965,N_4838,N_2879);
nor U5966 (N_5966,N_3377,N_4663);
and U5967 (N_5967,N_3921,N_4598);
or U5968 (N_5968,N_4921,N_4497);
xor U5969 (N_5969,N_3160,N_3788);
and U5970 (N_5970,N_3079,N_3862);
nand U5971 (N_5971,N_3707,N_4559);
nand U5972 (N_5972,N_4244,N_4482);
nor U5973 (N_5973,N_4096,N_2785);
xor U5974 (N_5974,N_2617,N_2914);
or U5975 (N_5975,N_4636,N_4330);
and U5976 (N_5976,N_2842,N_3458);
xnor U5977 (N_5977,N_3092,N_2923);
nand U5978 (N_5978,N_4248,N_4747);
nand U5979 (N_5979,N_3123,N_4625);
and U5980 (N_5980,N_3136,N_4717);
and U5981 (N_5981,N_3846,N_4259);
nand U5982 (N_5982,N_3292,N_2789);
nand U5983 (N_5983,N_2909,N_3319);
and U5984 (N_5984,N_3211,N_2783);
or U5985 (N_5985,N_4305,N_2847);
xnor U5986 (N_5986,N_2510,N_4525);
nand U5987 (N_5987,N_3395,N_3581);
nor U5988 (N_5988,N_3393,N_3819);
and U5989 (N_5989,N_3970,N_2731);
nor U5990 (N_5990,N_4757,N_4567);
nor U5991 (N_5991,N_4504,N_3452);
nor U5992 (N_5992,N_4863,N_3648);
nor U5993 (N_5993,N_4124,N_4456);
or U5994 (N_5994,N_4543,N_3461);
nand U5995 (N_5995,N_2967,N_2985);
and U5996 (N_5996,N_4283,N_3745);
or U5997 (N_5997,N_3039,N_3366);
and U5998 (N_5998,N_4595,N_2878);
nand U5999 (N_5999,N_3916,N_4313);
and U6000 (N_6000,N_4270,N_3011);
nand U6001 (N_6001,N_2730,N_2517);
or U6002 (N_6002,N_4062,N_3054);
nor U6003 (N_6003,N_2904,N_2746);
and U6004 (N_6004,N_2838,N_3547);
or U6005 (N_6005,N_2850,N_4205);
and U6006 (N_6006,N_3204,N_4713);
or U6007 (N_6007,N_3089,N_4123);
and U6008 (N_6008,N_4501,N_4002);
xnor U6009 (N_6009,N_3180,N_3494);
nor U6010 (N_6010,N_3227,N_2990);
nand U6011 (N_6011,N_4407,N_3347);
or U6012 (N_6012,N_3361,N_4768);
or U6013 (N_6013,N_4192,N_3853);
or U6014 (N_6014,N_4368,N_4533);
nor U6015 (N_6015,N_4835,N_4321);
nand U6016 (N_6016,N_4366,N_2903);
and U6017 (N_6017,N_4064,N_3613);
xnor U6018 (N_6018,N_4922,N_3638);
and U6019 (N_6019,N_2722,N_4430);
or U6020 (N_6020,N_3513,N_4491);
and U6021 (N_6021,N_2723,N_4287);
nand U6022 (N_6022,N_4617,N_3390);
and U6023 (N_6023,N_3290,N_4018);
and U6024 (N_6024,N_3399,N_4688);
nor U6025 (N_6025,N_4557,N_3262);
nand U6026 (N_6026,N_3173,N_4803);
xnor U6027 (N_6027,N_3067,N_4061);
nor U6028 (N_6028,N_3400,N_2944);
or U6029 (N_6029,N_4995,N_4274);
nor U6030 (N_6030,N_3966,N_2773);
and U6031 (N_6031,N_3057,N_2726);
nor U6032 (N_6032,N_4806,N_4432);
nand U6033 (N_6033,N_4496,N_3230);
or U6034 (N_6034,N_4337,N_3051);
or U6035 (N_6035,N_4034,N_2770);
nand U6036 (N_6036,N_3776,N_3676);
or U6037 (N_6037,N_4271,N_2649);
nand U6038 (N_6038,N_4856,N_2776);
or U6039 (N_6039,N_4011,N_3991);
and U6040 (N_6040,N_4730,N_4905);
or U6041 (N_6041,N_2831,N_3867);
nand U6042 (N_6042,N_4690,N_3394);
nand U6043 (N_6043,N_2501,N_3384);
xor U6044 (N_6044,N_3368,N_3006);
xor U6045 (N_6045,N_2779,N_4799);
and U6046 (N_6046,N_4208,N_3595);
nor U6047 (N_6047,N_2506,N_4333);
nand U6048 (N_6048,N_4412,N_4944);
nand U6049 (N_6049,N_3101,N_3608);
nor U6050 (N_6050,N_4872,N_4552);
nor U6051 (N_6051,N_4568,N_4119);
or U6052 (N_6052,N_4455,N_3923);
and U6053 (N_6053,N_4048,N_4178);
nor U6054 (N_6054,N_4484,N_3669);
and U6055 (N_6055,N_3045,N_4948);
nand U6056 (N_6056,N_4282,N_4984);
or U6057 (N_6057,N_2848,N_2867);
nand U6058 (N_6058,N_4109,N_3656);
nor U6059 (N_6059,N_3187,N_2511);
nand U6060 (N_6060,N_2917,N_3772);
nand U6061 (N_6061,N_2538,N_3899);
or U6062 (N_6062,N_3866,N_3694);
or U6063 (N_6063,N_3600,N_4722);
nand U6064 (N_6064,N_4638,N_4438);
nor U6065 (N_6065,N_2790,N_4303);
nand U6066 (N_6066,N_3718,N_4603);
xor U6067 (N_6067,N_3682,N_4291);
nand U6068 (N_6068,N_3146,N_4367);
xnor U6069 (N_6069,N_3534,N_3479);
and U6070 (N_6070,N_2781,N_2788);
nor U6071 (N_6071,N_3115,N_4158);
nand U6072 (N_6072,N_2771,N_3268);
nand U6073 (N_6073,N_3832,N_3664);
or U6074 (N_6074,N_2946,N_4970);
nor U6075 (N_6075,N_4991,N_3829);
or U6076 (N_6076,N_4975,N_3734);
and U6077 (N_6077,N_2852,N_4319);
and U6078 (N_6078,N_3781,N_2753);
or U6079 (N_6079,N_4145,N_4173);
and U6080 (N_6080,N_4527,N_4217);
nor U6081 (N_6081,N_2757,N_2540);
or U6082 (N_6082,N_4469,N_2570);
or U6083 (N_6083,N_3663,N_2725);
xor U6084 (N_6084,N_4453,N_4642);
and U6085 (N_6085,N_4296,N_3886);
or U6086 (N_6086,N_4716,N_3065);
nor U6087 (N_6087,N_2599,N_2527);
and U6088 (N_6088,N_3729,N_3179);
nand U6089 (N_6089,N_3887,N_4365);
or U6090 (N_6090,N_3200,N_2522);
xnor U6091 (N_6091,N_2663,N_2760);
or U6092 (N_6092,N_2628,N_4903);
nor U6093 (N_6093,N_4103,N_3854);
nand U6094 (N_6094,N_3498,N_2742);
nand U6095 (N_6095,N_4041,N_3805);
nand U6096 (N_6096,N_2678,N_2786);
and U6097 (N_6097,N_4320,N_3490);
or U6098 (N_6098,N_3942,N_2539);
xnor U6099 (N_6099,N_3910,N_2568);
nand U6100 (N_6100,N_3183,N_3449);
and U6101 (N_6101,N_4409,N_2660);
nand U6102 (N_6102,N_4211,N_4006);
nor U6103 (N_6103,N_3113,N_2870);
or U6104 (N_6104,N_3615,N_4986);
and U6105 (N_6105,N_3084,N_3859);
and U6106 (N_6106,N_2714,N_2606);
or U6107 (N_6107,N_3511,N_3240);
and U6108 (N_6108,N_3720,N_3174);
nor U6109 (N_6109,N_4895,N_3448);
xor U6110 (N_6110,N_4035,N_3312);
or U6111 (N_6111,N_2969,N_3906);
nor U6112 (N_6112,N_4427,N_2875);
xnor U6113 (N_6113,N_2622,N_4393);
and U6114 (N_6114,N_2756,N_2537);
nand U6115 (N_6115,N_3799,N_3983);
nand U6116 (N_6116,N_4392,N_3520);
xor U6117 (N_6117,N_4262,N_2744);
nand U6118 (N_6118,N_4883,N_2869);
nand U6119 (N_6119,N_3353,N_2595);
and U6120 (N_6120,N_3107,N_3081);
or U6121 (N_6121,N_4524,N_3352);
or U6122 (N_6122,N_4451,N_4445);
and U6123 (N_6123,N_4003,N_4648);
xnor U6124 (N_6124,N_3073,N_4859);
or U6125 (N_6125,N_2965,N_2583);
xnor U6126 (N_6126,N_2573,N_4643);
and U6127 (N_6127,N_4562,N_4489);
and U6128 (N_6128,N_3579,N_4840);
nand U6129 (N_6129,N_4779,N_2584);
nand U6130 (N_6130,N_3605,N_4810);
or U6131 (N_6131,N_4867,N_4122);
nand U6132 (N_6132,N_3058,N_4266);
nor U6133 (N_6133,N_2664,N_3857);
and U6134 (N_6134,N_3717,N_3423);
nor U6135 (N_6135,N_3046,N_3147);
nor U6136 (N_6136,N_3197,N_4417);
nor U6137 (N_6137,N_3523,N_4609);
nor U6138 (N_6138,N_4936,N_2740);
nand U6139 (N_6139,N_4084,N_3332);
nand U6140 (N_6140,N_3221,N_3834);
nand U6141 (N_6141,N_4332,N_4507);
nand U6142 (N_6142,N_4162,N_3325);
and U6143 (N_6143,N_4111,N_3706);
and U6144 (N_6144,N_2528,N_4529);
or U6145 (N_6145,N_4735,N_4384);
nor U6146 (N_6146,N_3836,N_3482);
or U6147 (N_6147,N_2993,N_3786);
and U6148 (N_6148,N_2988,N_3002);
xor U6149 (N_6149,N_3701,N_4269);
nand U6150 (N_6150,N_3254,N_3229);
nor U6151 (N_6151,N_4814,N_2626);
nand U6152 (N_6152,N_4987,N_4622);
or U6153 (N_6153,N_3355,N_3582);
nand U6154 (N_6154,N_4538,N_4227);
nor U6155 (N_6155,N_3437,N_2699);
nor U6156 (N_6156,N_4039,N_2561);
and U6157 (N_6157,N_3993,N_3560);
nand U6158 (N_6158,N_2841,N_4604);
or U6159 (N_6159,N_2693,N_4054);
or U6160 (N_6160,N_3431,N_3031);
or U6161 (N_6161,N_2894,N_3499);
nand U6162 (N_6162,N_4864,N_4228);
or U6163 (N_6163,N_4154,N_3192);
nand U6164 (N_6164,N_2716,N_3952);
nand U6165 (N_6165,N_4561,N_4992);
nand U6166 (N_6166,N_4159,N_4931);
nor U6167 (N_6167,N_3699,N_2647);
nor U6168 (N_6168,N_3028,N_4042);
nor U6169 (N_6169,N_2514,N_4253);
nor U6170 (N_6170,N_3005,N_4920);
nor U6171 (N_6171,N_4950,N_3594);
or U6172 (N_6172,N_4668,N_3143);
and U6173 (N_6173,N_3675,N_2671);
nand U6174 (N_6174,N_3360,N_3345);
and U6175 (N_6175,N_2651,N_3375);
xnor U6176 (N_6176,N_4396,N_4081);
nand U6177 (N_6177,N_3135,N_4854);
nand U6178 (N_6178,N_3035,N_4083);
or U6179 (N_6179,N_3095,N_4126);
or U6180 (N_6180,N_4767,N_4328);
nand U6181 (N_6181,N_2586,N_2811);
or U6182 (N_6182,N_2598,N_3771);
nor U6183 (N_6183,N_2674,N_3662);
and U6184 (N_6184,N_3220,N_4428);
nand U6185 (N_6185,N_2536,N_4051);
nor U6186 (N_6186,N_4517,N_3271);
nor U6187 (N_6187,N_4667,N_3358);
and U6188 (N_6188,N_4744,N_3968);
or U6189 (N_6189,N_3409,N_4868);
nor U6190 (N_6190,N_2641,N_3298);
and U6191 (N_6191,N_4588,N_3484);
nor U6192 (N_6192,N_3213,N_2932);
or U6193 (N_6193,N_4488,N_2609);
and U6194 (N_6194,N_4890,N_2972);
nand U6195 (N_6195,N_3914,N_3438);
or U6196 (N_6196,N_4708,N_3025);
and U6197 (N_6197,N_3314,N_4416);
or U6198 (N_6198,N_3489,N_3477);
and U6199 (N_6199,N_4554,N_3730);
nand U6200 (N_6200,N_3824,N_3946);
and U6201 (N_6201,N_3453,N_3138);
nand U6202 (N_6202,N_2518,N_3860);
nand U6203 (N_6203,N_3351,N_4565);
and U6204 (N_6204,N_3168,N_3529);
nor U6205 (N_6205,N_4130,N_3620);
nor U6206 (N_6206,N_3406,N_4346);
or U6207 (N_6207,N_3411,N_2930);
nor U6208 (N_6208,N_2680,N_2772);
and U6209 (N_6209,N_2646,N_4847);
nand U6210 (N_6210,N_2705,N_2508);
and U6211 (N_6211,N_2808,N_2579);
nor U6212 (N_6212,N_3464,N_4464);
nand U6213 (N_6213,N_4791,N_4798);
nor U6214 (N_6214,N_4378,N_4952);
nor U6215 (N_6215,N_4063,N_4198);
or U6216 (N_6216,N_4129,N_3645);
nor U6217 (N_6217,N_4607,N_4374);
nand U6218 (N_6218,N_3785,N_3593);
nand U6219 (N_6219,N_4025,N_2580);
and U6220 (N_6220,N_3048,N_3279);
and U6221 (N_6221,N_3198,N_2590);
xor U6222 (N_6222,N_4551,N_4419);
and U6223 (N_6223,N_3103,N_4790);
or U6224 (N_6224,N_4879,N_4036);
and U6225 (N_6225,N_4175,N_4513);
nor U6226 (N_6226,N_4265,N_3724);
nand U6227 (N_6227,N_2973,N_4401);
or U6228 (N_6228,N_2551,N_3943);
and U6229 (N_6229,N_3212,N_2524);
or U6230 (N_6230,N_4530,N_2981);
and U6231 (N_6231,N_3432,N_2635);
nand U6232 (N_6232,N_2791,N_4549);
or U6233 (N_6233,N_3823,N_4045);
or U6234 (N_6234,N_3038,N_3903);
nand U6235 (N_6235,N_4157,N_4898);
or U6236 (N_6236,N_4229,N_3960);
nor U6237 (N_6237,N_4377,N_3026);
or U6238 (N_6238,N_4134,N_4727);
nor U6239 (N_6239,N_4317,N_4813);
nand U6240 (N_6240,N_4075,N_2526);
or U6241 (N_6241,N_3202,N_4483);
nor U6242 (N_6242,N_3759,N_4601);
nor U6243 (N_6243,N_3733,N_2910);
or U6244 (N_6244,N_2603,N_3604);
and U6245 (N_6245,N_3281,N_4185);
nor U6246 (N_6246,N_3959,N_4878);
nand U6247 (N_6247,N_4351,N_3700);
and U6248 (N_6248,N_4592,N_4027);
or U6249 (N_6249,N_2577,N_2653);
or U6250 (N_6250,N_4788,N_3997);
and U6251 (N_6251,N_3334,N_3785);
nor U6252 (N_6252,N_2826,N_2817);
xnor U6253 (N_6253,N_4312,N_3713);
or U6254 (N_6254,N_3869,N_2547);
nor U6255 (N_6255,N_2817,N_3837);
nor U6256 (N_6256,N_2666,N_4967);
nor U6257 (N_6257,N_2697,N_4262);
nor U6258 (N_6258,N_4072,N_4635);
nor U6259 (N_6259,N_4865,N_4560);
nand U6260 (N_6260,N_3130,N_4019);
or U6261 (N_6261,N_2684,N_4436);
nand U6262 (N_6262,N_2676,N_4936);
xnor U6263 (N_6263,N_3046,N_2978);
nor U6264 (N_6264,N_4064,N_2706);
nand U6265 (N_6265,N_4556,N_3615);
xor U6266 (N_6266,N_3608,N_3030);
xor U6267 (N_6267,N_2926,N_3739);
or U6268 (N_6268,N_4597,N_3134);
or U6269 (N_6269,N_2830,N_2622);
and U6270 (N_6270,N_4060,N_2878);
and U6271 (N_6271,N_3346,N_4577);
and U6272 (N_6272,N_4083,N_4895);
and U6273 (N_6273,N_2624,N_4853);
nor U6274 (N_6274,N_2620,N_3461);
nand U6275 (N_6275,N_3224,N_4377);
nand U6276 (N_6276,N_4218,N_3940);
or U6277 (N_6277,N_4831,N_2651);
and U6278 (N_6278,N_4035,N_4959);
nor U6279 (N_6279,N_3906,N_4051);
nand U6280 (N_6280,N_3439,N_3253);
nor U6281 (N_6281,N_2894,N_3604);
and U6282 (N_6282,N_2959,N_4431);
nand U6283 (N_6283,N_3642,N_2563);
nand U6284 (N_6284,N_4565,N_3050);
or U6285 (N_6285,N_4357,N_3949);
nor U6286 (N_6286,N_4186,N_2791);
xor U6287 (N_6287,N_2619,N_4562);
nor U6288 (N_6288,N_4365,N_4451);
and U6289 (N_6289,N_4061,N_4076);
nor U6290 (N_6290,N_4501,N_3864);
and U6291 (N_6291,N_4419,N_2761);
nor U6292 (N_6292,N_3782,N_4836);
nand U6293 (N_6293,N_3785,N_2870);
or U6294 (N_6294,N_4151,N_4779);
nand U6295 (N_6295,N_3447,N_4882);
nand U6296 (N_6296,N_4065,N_3330);
nor U6297 (N_6297,N_4480,N_3189);
or U6298 (N_6298,N_3659,N_2697);
nor U6299 (N_6299,N_2956,N_3507);
and U6300 (N_6300,N_4469,N_4983);
nor U6301 (N_6301,N_2510,N_3356);
nand U6302 (N_6302,N_3842,N_4079);
and U6303 (N_6303,N_3180,N_3499);
nand U6304 (N_6304,N_2671,N_4999);
nand U6305 (N_6305,N_3408,N_3812);
xnor U6306 (N_6306,N_4611,N_4929);
or U6307 (N_6307,N_3519,N_4473);
xnor U6308 (N_6308,N_2669,N_3760);
nor U6309 (N_6309,N_4513,N_2554);
or U6310 (N_6310,N_4961,N_4681);
xnor U6311 (N_6311,N_3506,N_4211);
and U6312 (N_6312,N_2639,N_4676);
xor U6313 (N_6313,N_4623,N_3580);
or U6314 (N_6314,N_3959,N_4455);
and U6315 (N_6315,N_3922,N_4409);
nor U6316 (N_6316,N_4467,N_4015);
and U6317 (N_6317,N_4299,N_2763);
nor U6318 (N_6318,N_4555,N_4197);
nand U6319 (N_6319,N_3076,N_2866);
or U6320 (N_6320,N_4203,N_3728);
or U6321 (N_6321,N_2620,N_4923);
and U6322 (N_6322,N_4403,N_4364);
or U6323 (N_6323,N_3204,N_3702);
and U6324 (N_6324,N_3153,N_4050);
and U6325 (N_6325,N_4561,N_3735);
and U6326 (N_6326,N_2643,N_4775);
xor U6327 (N_6327,N_4580,N_3562);
nand U6328 (N_6328,N_3110,N_3287);
and U6329 (N_6329,N_3886,N_3199);
nor U6330 (N_6330,N_2615,N_4425);
and U6331 (N_6331,N_4657,N_2978);
nor U6332 (N_6332,N_3425,N_3396);
or U6333 (N_6333,N_4200,N_2698);
nor U6334 (N_6334,N_4977,N_3667);
nand U6335 (N_6335,N_2969,N_4229);
nor U6336 (N_6336,N_4333,N_4343);
and U6337 (N_6337,N_3703,N_3324);
or U6338 (N_6338,N_4358,N_2836);
or U6339 (N_6339,N_4686,N_3523);
nand U6340 (N_6340,N_3162,N_3947);
nand U6341 (N_6341,N_3892,N_3962);
nand U6342 (N_6342,N_4586,N_3912);
or U6343 (N_6343,N_4356,N_2961);
nand U6344 (N_6344,N_2834,N_2916);
nor U6345 (N_6345,N_3262,N_3667);
and U6346 (N_6346,N_2631,N_4439);
nand U6347 (N_6347,N_3075,N_3661);
and U6348 (N_6348,N_2690,N_4236);
nand U6349 (N_6349,N_3318,N_3952);
nor U6350 (N_6350,N_3414,N_4972);
or U6351 (N_6351,N_3278,N_3028);
or U6352 (N_6352,N_3544,N_4302);
nor U6353 (N_6353,N_4546,N_4502);
nand U6354 (N_6354,N_3445,N_4569);
xnor U6355 (N_6355,N_4651,N_3998);
and U6356 (N_6356,N_3754,N_2871);
xor U6357 (N_6357,N_4577,N_4103);
nor U6358 (N_6358,N_4419,N_3435);
and U6359 (N_6359,N_2877,N_4619);
nor U6360 (N_6360,N_4286,N_4487);
nand U6361 (N_6361,N_4213,N_3319);
nand U6362 (N_6362,N_4626,N_4365);
and U6363 (N_6363,N_3928,N_3109);
or U6364 (N_6364,N_2714,N_2633);
or U6365 (N_6365,N_3968,N_4335);
nor U6366 (N_6366,N_3955,N_4958);
nand U6367 (N_6367,N_3251,N_4900);
nand U6368 (N_6368,N_4637,N_4765);
and U6369 (N_6369,N_4381,N_4097);
nor U6370 (N_6370,N_4885,N_4914);
nand U6371 (N_6371,N_2912,N_2900);
and U6372 (N_6372,N_4370,N_4590);
or U6373 (N_6373,N_3364,N_3884);
xor U6374 (N_6374,N_2785,N_3818);
nand U6375 (N_6375,N_3081,N_3921);
nor U6376 (N_6376,N_3633,N_3011);
nand U6377 (N_6377,N_2960,N_3449);
nand U6378 (N_6378,N_4563,N_4001);
nor U6379 (N_6379,N_3786,N_4106);
nor U6380 (N_6380,N_3896,N_3905);
nor U6381 (N_6381,N_3830,N_2708);
or U6382 (N_6382,N_3517,N_2938);
and U6383 (N_6383,N_4769,N_3034);
nand U6384 (N_6384,N_3465,N_4409);
nand U6385 (N_6385,N_4538,N_2925);
nor U6386 (N_6386,N_2720,N_2809);
xor U6387 (N_6387,N_2630,N_4480);
nor U6388 (N_6388,N_4557,N_4495);
and U6389 (N_6389,N_4203,N_2514);
nor U6390 (N_6390,N_3058,N_3459);
and U6391 (N_6391,N_4376,N_4931);
nand U6392 (N_6392,N_4110,N_3147);
xnor U6393 (N_6393,N_2711,N_4057);
and U6394 (N_6394,N_3892,N_3716);
or U6395 (N_6395,N_4845,N_3748);
nor U6396 (N_6396,N_4552,N_4228);
nand U6397 (N_6397,N_4083,N_4439);
or U6398 (N_6398,N_4326,N_4199);
or U6399 (N_6399,N_3302,N_3969);
and U6400 (N_6400,N_4717,N_3806);
or U6401 (N_6401,N_2980,N_2630);
nand U6402 (N_6402,N_2878,N_4122);
or U6403 (N_6403,N_4277,N_3807);
nand U6404 (N_6404,N_4199,N_3396);
and U6405 (N_6405,N_4428,N_4582);
or U6406 (N_6406,N_2733,N_3383);
xnor U6407 (N_6407,N_3634,N_4751);
or U6408 (N_6408,N_3214,N_3457);
nor U6409 (N_6409,N_4627,N_4070);
nand U6410 (N_6410,N_4737,N_4661);
nand U6411 (N_6411,N_4507,N_4731);
xnor U6412 (N_6412,N_3094,N_3651);
and U6413 (N_6413,N_4998,N_4861);
nand U6414 (N_6414,N_3763,N_2547);
nand U6415 (N_6415,N_3072,N_4396);
or U6416 (N_6416,N_3004,N_3611);
and U6417 (N_6417,N_4672,N_2764);
nand U6418 (N_6418,N_3791,N_4936);
nor U6419 (N_6419,N_3796,N_4277);
nor U6420 (N_6420,N_2628,N_4169);
or U6421 (N_6421,N_4879,N_4270);
or U6422 (N_6422,N_4761,N_2559);
or U6423 (N_6423,N_3041,N_3114);
nand U6424 (N_6424,N_4997,N_3414);
or U6425 (N_6425,N_4136,N_3463);
or U6426 (N_6426,N_3492,N_4856);
and U6427 (N_6427,N_4351,N_3520);
or U6428 (N_6428,N_4999,N_4920);
xor U6429 (N_6429,N_2572,N_4049);
or U6430 (N_6430,N_4634,N_3801);
or U6431 (N_6431,N_3167,N_3667);
nor U6432 (N_6432,N_4039,N_2731);
nor U6433 (N_6433,N_3037,N_4559);
or U6434 (N_6434,N_3238,N_3532);
and U6435 (N_6435,N_3000,N_4357);
or U6436 (N_6436,N_3206,N_2881);
and U6437 (N_6437,N_4791,N_2790);
nand U6438 (N_6438,N_3148,N_4149);
nor U6439 (N_6439,N_2604,N_3753);
and U6440 (N_6440,N_4981,N_4918);
and U6441 (N_6441,N_2545,N_2835);
nor U6442 (N_6442,N_3597,N_3017);
xor U6443 (N_6443,N_4820,N_2791);
or U6444 (N_6444,N_4896,N_4859);
nor U6445 (N_6445,N_3262,N_2887);
nor U6446 (N_6446,N_3039,N_4618);
nand U6447 (N_6447,N_4760,N_4498);
nand U6448 (N_6448,N_4368,N_4334);
nor U6449 (N_6449,N_2988,N_3068);
or U6450 (N_6450,N_3820,N_4974);
nor U6451 (N_6451,N_4451,N_4020);
nand U6452 (N_6452,N_4785,N_4311);
or U6453 (N_6453,N_4631,N_4780);
nor U6454 (N_6454,N_2725,N_3031);
or U6455 (N_6455,N_4025,N_3979);
and U6456 (N_6456,N_4552,N_3911);
nand U6457 (N_6457,N_4591,N_3402);
or U6458 (N_6458,N_4535,N_4796);
xor U6459 (N_6459,N_2652,N_3963);
nand U6460 (N_6460,N_3013,N_4672);
nand U6461 (N_6461,N_4886,N_3243);
nand U6462 (N_6462,N_4077,N_4432);
and U6463 (N_6463,N_2579,N_2716);
and U6464 (N_6464,N_4873,N_4884);
nand U6465 (N_6465,N_4384,N_4813);
and U6466 (N_6466,N_4790,N_4966);
xnor U6467 (N_6467,N_3588,N_2962);
and U6468 (N_6468,N_3415,N_4152);
and U6469 (N_6469,N_3462,N_4876);
nand U6470 (N_6470,N_3281,N_3625);
or U6471 (N_6471,N_4967,N_3422);
and U6472 (N_6472,N_3799,N_3626);
and U6473 (N_6473,N_3817,N_3167);
or U6474 (N_6474,N_4888,N_4097);
nor U6475 (N_6475,N_4487,N_4478);
or U6476 (N_6476,N_3141,N_3718);
nand U6477 (N_6477,N_3064,N_3491);
and U6478 (N_6478,N_2650,N_3078);
xnor U6479 (N_6479,N_4068,N_3531);
or U6480 (N_6480,N_3724,N_4860);
and U6481 (N_6481,N_4914,N_2718);
nand U6482 (N_6482,N_4248,N_3119);
and U6483 (N_6483,N_4514,N_4553);
nor U6484 (N_6484,N_3083,N_3675);
nor U6485 (N_6485,N_4219,N_3092);
or U6486 (N_6486,N_3259,N_3987);
xnor U6487 (N_6487,N_2623,N_2710);
and U6488 (N_6488,N_4227,N_3429);
nand U6489 (N_6489,N_3535,N_4274);
nand U6490 (N_6490,N_3243,N_4407);
or U6491 (N_6491,N_2879,N_4559);
and U6492 (N_6492,N_3426,N_2595);
and U6493 (N_6493,N_4568,N_4967);
and U6494 (N_6494,N_3178,N_4687);
or U6495 (N_6495,N_3819,N_4819);
nand U6496 (N_6496,N_4727,N_4231);
and U6497 (N_6497,N_3936,N_4627);
and U6498 (N_6498,N_3538,N_3176);
nand U6499 (N_6499,N_3314,N_3554);
nand U6500 (N_6500,N_3908,N_4102);
or U6501 (N_6501,N_2933,N_2767);
nand U6502 (N_6502,N_4661,N_4272);
nor U6503 (N_6503,N_4034,N_2940);
xnor U6504 (N_6504,N_2607,N_3939);
or U6505 (N_6505,N_2720,N_4638);
nor U6506 (N_6506,N_4610,N_4268);
or U6507 (N_6507,N_3629,N_3203);
nor U6508 (N_6508,N_4539,N_3894);
nand U6509 (N_6509,N_3572,N_4271);
or U6510 (N_6510,N_2830,N_3304);
nand U6511 (N_6511,N_3303,N_2847);
nor U6512 (N_6512,N_3763,N_4201);
nand U6513 (N_6513,N_3407,N_2954);
or U6514 (N_6514,N_4258,N_4359);
nand U6515 (N_6515,N_2827,N_3150);
nor U6516 (N_6516,N_4451,N_3276);
or U6517 (N_6517,N_4057,N_4808);
or U6518 (N_6518,N_2760,N_4182);
and U6519 (N_6519,N_4513,N_3020);
and U6520 (N_6520,N_3131,N_3151);
nor U6521 (N_6521,N_4916,N_3394);
or U6522 (N_6522,N_2564,N_4025);
and U6523 (N_6523,N_4693,N_3688);
xor U6524 (N_6524,N_2510,N_3674);
or U6525 (N_6525,N_4064,N_3442);
nor U6526 (N_6526,N_3129,N_3788);
nand U6527 (N_6527,N_3516,N_2585);
nand U6528 (N_6528,N_4430,N_2915);
xnor U6529 (N_6529,N_3214,N_3194);
or U6530 (N_6530,N_2978,N_4916);
and U6531 (N_6531,N_4103,N_4774);
nand U6532 (N_6532,N_3423,N_4259);
nor U6533 (N_6533,N_3360,N_2987);
nor U6534 (N_6534,N_4064,N_2501);
or U6535 (N_6535,N_2549,N_4251);
nand U6536 (N_6536,N_3347,N_2995);
or U6537 (N_6537,N_3241,N_3668);
nand U6538 (N_6538,N_3132,N_2732);
or U6539 (N_6539,N_4039,N_4947);
or U6540 (N_6540,N_4584,N_4057);
and U6541 (N_6541,N_2967,N_2566);
nand U6542 (N_6542,N_3419,N_2642);
nor U6543 (N_6543,N_3680,N_4240);
nand U6544 (N_6544,N_4984,N_4919);
nor U6545 (N_6545,N_4257,N_4733);
nand U6546 (N_6546,N_2587,N_3484);
nand U6547 (N_6547,N_3169,N_4725);
nand U6548 (N_6548,N_2619,N_2627);
or U6549 (N_6549,N_3958,N_2700);
nand U6550 (N_6550,N_3774,N_2620);
and U6551 (N_6551,N_4655,N_4596);
and U6552 (N_6552,N_4019,N_2968);
nand U6553 (N_6553,N_3612,N_4256);
xor U6554 (N_6554,N_3919,N_2804);
nor U6555 (N_6555,N_3359,N_3522);
nor U6556 (N_6556,N_3585,N_4143);
nor U6557 (N_6557,N_4170,N_4064);
or U6558 (N_6558,N_3730,N_4530);
and U6559 (N_6559,N_3661,N_3257);
or U6560 (N_6560,N_3441,N_2730);
and U6561 (N_6561,N_2647,N_4330);
and U6562 (N_6562,N_4786,N_3698);
nand U6563 (N_6563,N_3676,N_3861);
nand U6564 (N_6564,N_3813,N_2705);
nand U6565 (N_6565,N_2940,N_3695);
and U6566 (N_6566,N_2787,N_3527);
and U6567 (N_6567,N_4580,N_3656);
nand U6568 (N_6568,N_4154,N_4195);
xnor U6569 (N_6569,N_3580,N_4664);
nand U6570 (N_6570,N_4933,N_3270);
nand U6571 (N_6571,N_4333,N_4072);
or U6572 (N_6572,N_2663,N_4711);
nand U6573 (N_6573,N_4950,N_4180);
nand U6574 (N_6574,N_4513,N_4926);
and U6575 (N_6575,N_4859,N_3689);
or U6576 (N_6576,N_4374,N_3702);
and U6577 (N_6577,N_3438,N_2963);
xor U6578 (N_6578,N_3123,N_4187);
nor U6579 (N_6579,N_2529,N_2520);
xor U6580 (N_6580,N_2834,N_2858);
and U6581 (N_6581,N_2938,N_3208);
xor U6582 (N_6582,N_3088,N_3507);
nor U6583 (N_6583,N_3042,N_3498);
nand U6584 (N_6584,N_4463,N_4391);
and U6585 (N_6585,N_2837,N_3791);
nor U6586 (N_6586,N_3537,N_4766);
nor U6587 (N_6587,N_3839,N_3052);
nand U6588 (N_6588,N_2972,N_4338);
or U6589 (N_6589,N_3872,N_3153);
and U6590 (N_6590,N_2735,N_4619);
nand U6591 (N_6591,N_2725,N_4480);
and U6592 (N_6592,N_4005,N_2667);
nor U6593 (N_6593,N_3103,N_4239);
nand U6594 (N_6594,N_2528,N_2896);
nor U6595 (N_6595,N_4344,N_4111);
nand U6596 (N_6596,N_3737,N_4046);
and U6597 (N_6597,N_4113,N_2868);
or U6598 (N_6598,N_4929,N_4233);
or U6599 (N_6599,N_3100,N_3192);
nand U6600 (N_6600,N_2684,N_3819);
and U6601 (N_6601,N_4127,N_4948);
nor U6602 (N_6602,N_3282,N_3650);
xor U6603 (N_6603,N_4913,N_2958);
nand U6604 (N_6604,N_3851,N_2575);
nor U6605 (N_6605,N_3512,N_3835);
nand U6606 (N_6606,N_4149,N_2586);
and U6607 (N_6607,N_3206,N_4009);
or U6608 (N_6608,N_4190,N_2627);
xor U6609 (N_6609,N_4443,N_3219);
and U6610 (N_6610,N_2607,N_3508);
and U6611 (N_6611,N_2538,N_4972);
or U6612 (N_6612,N_4313,N_3618);
nor U6613 (N_6613,N_4766,N_2544);
and U6614 (N_6614,N_4031,N_4928);
nand U6615 (N_6615,N_4449,N_4930);
or U6616 (N_6616,N_4058,N_3341);
nor U6617 (N_6617,N_4244,N_2796);
nor U6618 (N_6618,N_3142,N_2910);
nor U6619 (N_6619,N_2982,N_4591);
or U6620 (N_6620,N_2667,N_2563);
nor U6621 (N_6621,N_3368,N_4023);
xor U6622 (N_6622,N_4567,N_3204);
and U6623 (N_6623,N_3403,N_4593);
nor U6624 (N_6624,N_3074,N_4861);
nand U6625 (N_6625,N_4931,N_3132);
and U6626 (N_6626,N_4394,N_4220);
or U6627 (N_6627,N_4114,N_3566);
or U6628 (N_6628,N_3587,N_3162);
nor U6629 (N_6629,N_3504,N_4516);
and U6630 (N_6630,N_3340,N_3500);
or U6631 (N_6631,N_4124,N_3404);
or U6632 (N_6632,N_3931,N_3514);
xor U6633 (N_6633,N_4623,N_4056);
and U6634 (N_6634,N_2922,N_3060);
nand U6635 (N_6635,N_2732,N_4168);
or U6636 (N_6636,N_2505,N_4518);
or U6637 (N_6637,N_4010,N_4603);
or U6638 (N_6638,N_2606,N_3621);
and U6639 (N_6639,N_2786,N_4461);
and U6640 (N_6640,N_4536,N_2728);
nor U6641 (N_6641,N_2536,N_4343);
nand U6642 (N_6642,N_4153,N_4899);
nand U6643 (N_6643,N_4472,N_2522);
nor U6644 (N_6644,N_4430,N_4795);
xor U6645 (N_6645,N_4363,N_4829);
nor U6646 (N_6646,N_2835,N_4507);
xor U6647 (N_6647,N_4733,N_2593);
or U6648 (N_6648,N_2682,N_3683);
and U6649 (N_6649,N_3435,N_4572);
and U6650 (N_6650,N_3484,N_3254);
or U6651 (N_6651,N_3304,N_3940);
nand U6652 (N_6652,N_4349,N_2698);
nand U6653 (N_6653,N_2738,N_3801);
and U6654 (N_6654,N_3053,N_4545);
nand U6655 (N_6655,N_4712,N_3779);
nor U6656 (N_6656,N_4430,N_2604);
or U6657 (N_6657,N_4615,N_3070);
xnor U6658 (N_6658,N_4600,N_3037);
nor U6659 (N_6659,N_2848,N_4133);
nor U6660 (N_6660,N_3090,N_2949);
nor U6661 (N_6661,N_4642,N_3394);
xnor U6662 (N_6662,N_3487,N_4089);
nor U6663 (N_6663,N_3381,N_2757);
nor U6664 (N_6664,N_4373,N_4302);
nand U6665 (N_6665,N_3746,N_2771);
nand U6666 (N_6666,N_4956,N_3026);
and U6667 (N_6667,N_4891,N_3286);
nor U6668 (N_6668,N_4872,N_4740);
or U6669 (N_6669,N_3492,N_3715);
nand U6670 (N_6670,N_2681,N_3418);
or U6671 (N_6671,N_3873,N_3025);
and U6672 (N_6672,N_4040,N_3575);
xor U6673 (N_6673,N_4956,N_3264);
or U6674 (N_6674,N_4106,N_3434);
nand U6675 (N_6675,N_4673,N_4544);
nand U6676 (N_6676,N_2796,N_2672);
or U6677 (N_6677,N_2879,N_4700);
nand U6678 (N_6678,N_4410,N_4472);
nand U6679 (N_6679,N_3493,N_4618);
or U6680 (N_6680,N_4458,N_4217);
and U6681 (N_6681,N_3469,N_4903);
xnor U6682 (N_6682,N_2859,N_4588);
or U6683 (N_6683,N_2511,N_3971);
and U6684 (N_6684,N_3013,N_3678);
and U6685 (N_6685,N_3371,N_4668);
and U6686 (N_6686,N_3997,N_3952);
or U6687 (N_6687,N_2609,N_3951);
and U6688 (N_6688,N_3254,N_2771);
nand U6689 (N_6689,N_2524,N_3750);
nand U6690 (N_6690,N_3614,N_3640);
nand U6691 (N_6691,N_2702,N_4935);
xnor U6692 (N_6692,N_2708,N_3232);
nand U6693 (N_6693,N_2710,N_4524);
nor U6694 (N_6694,N_4319,N_3194);
or U6695 (N_6695,N_4467,N_2549);
and U6696 (N_6696,N_4681,N_3542);
or U6697 (N_6697,N_3575,N_3310);
nand U6698 (N_6698,N_3645,N_3445);
nand U6699 (N_6699,N_3982,N_4214);
and U6700 (N_6700,N_3439,N_2886);
nand U6701 (N_6701,N_3797,N_4081);
nor U6702 (N_6702,N_3633,N_4585);
nor U6703 (N_6703,N_4753,N_4839);
nand U6704 (N_6704,N_4446,N_4056);
nand U6705 (N_6705,N_3325,N_2969);
nand U6706 (N_6706,N_2744,N_4035);
and U6707 (N_6707,N_3525,N_4517);
or U6708 (N_6708,N_4777,N_3625);
nand U6709 (N_6709,N_4366,N_2753);
nand U6710 (N_6710,N_3249,N_2526);
nor U6711 (N_6711,N_3590,N_4617);
or U6712 (N_6712,N_2911,N_3898);
nand U6713 (N_6713,N_3917,N_3671);
or U6714 (N_6714,N_3312,N_3953);
and U6715 (N_6715,N_4625,N_3238);
nor U6716 (N_6716,N_3962,N_4581);
and U6717 (N_6717,N_2773,N_4298);
and U6718 (N_6718,N_2829,N_2994);
nand U6719 (N_6719,N_2667,N_3526);
and U6720 (N_6720,N_3000,N_4850);
nand U6721 (N_6721,N_2521,N_3990);
nand U6722 (N_6722,N_3223,N_4833);
or U6723 (N_6723,N_3579,N_4218);
nor U6724 (N_6724,N_4754,N_3219);
or U6725 (N_6725,N_3771,N_4479);
nand U6726 (N_6726,N_4034,N_2912);
xnor U6727 (N_6727,N_3450,N_3462);
and U6728 (N_6728,N_4604,N_4702);
xnor U6729 (N_6729,N_3081,N_2992);
nand U6730 (N_6730,N_2702,N_4514);
nor U6731 (N_6731,N_4971,N_3714);
and U6732 (N_6732,N_3227,N_3215);
xor U6733 (N_6733,N_4940,N_3429);
or U6734 (N_6734,N_3426,N_3725);
or U6735 (N_6735,N_3920,N_4874);
or U6736 (N_6736,N_4062,N_4748);
and U6737 (N_6737,N_4064,N_2810);
nor U6738 (N_6738,N_3745,N_4738);
nand U6739 (N_6739,N_3639,N_3111);
xor U6740 (N_6740,N_3188,N_4415);
and U6741 (N_6741,N_3857,N_2609);
xnor U6742 (N_6742,N_3461,N_3880);
and U6743 (N_6743,N_4441,N_2878);
nand U6744 (N_6744,N_3413,N_4990);
or U6745 (N_6745,N_2952,N_4889);
nand U6746 (N_6746,N_3011,N_4334);
nor U6747 (N_6747,N_4485,N_4622);
or U6748 (N_6748,N_3790,N_2900);
or U6749 (N_6749,N_2937,N_3481);
or U6750 (N_6750,N_3167,N_2994);
or U6751 (N_6751,N_3564,N_3836);
nor U6752 (N_6752,N_4217,N_3337);
nor U6753 (N_6753,N_2891,N_2968);
nor U6754 (N_6754,N_2500,N_4614);
and U6755 (N_6755,N_4970,N_4746);
nand U6756 (N_6756,N_4504,N_3609);
nor U6757 (N_6757,N_4552,N_3579);
or U6758 (N_6758,N_2781,N_3406);
nor U6759 (N_6759,N_4471,N_2667);
nor U6760 (N_6760,N_4282,N_3922);
nor U6761 (N_6761,N_4163,N_2736);
nand U6762 (N_6762,N_4800,N_3904);
nand U6763 (N_6763,N_3283,N_4563);
nor U6764 (N_6764,N_4695,N_4725);
xnor U6765 (N_6765,N_2838,N_3112);
xor U6766 (N_6766,N_4352,N_4368);
nand U6767 (N_6767,N_4466,N_3501);
and U6768 (N_6768,N_2580,N_3762);
nand U6769 (N_6769,N_4575,N_4644);
or U6770 (N_6770,N_4369,N_2665);
nor U6771 (N_6771,N_4649,N_3995);
nand U6772 (N_6772,N_3820,N_2784);
xor U6773 (N_6773,N_2897,N_4554);
and U6774 (N_6774,N_3662,N_3725);
and U6775 (N_6775,N_4379,N_2833);
nand U6776 (N_6776,N_2944,N_2941);
nand U6777 (N_6777,N_4520,N_2856);
nor U6778 (N_6778,N_3848,N_4446);
xor U6779 (N_6779,N_4059,N_4380);
nand U6780 (N_6780,N_4616,N_4287);
and U6781 (N_6781,N_3397,N_2670);
nand U6782 (N_6782,N_4895,N_4441);
nor U6783 (N_6783,N_4926,N_2736);
or U6784 (N_6784,N_3142,N_4362);
or U6785 (N_6785,N_3495,N_3882);
nand U6786 (N_6786,N_3428,N_4007);
nand U6787 (N_6787,N_4003,N_3259);
xnor U6788 (N_6788,N_4592,N_3603);
and U6789 (N_6789,N_4570,N_3287);
and U6790 (N_6790,N_2862,N_2657);
and U6791 (N_6791,N_4382,N_2960);
and U6792 (N_6792,N_3564,N_4521);
and U6793 (N_6793,N_3319,N_2906);
nand U6794 (N_6794,N_2924,N_3596);
nor U6795 (N_6795,N_3518,N_3880);
xor U6796 (N_6796,N_2547,N_4663);
nor U6797 (N_6797,N_3138,N_4146);
nand U6798 (N_6798,N_3898,N_4020);
nor U6799 (N_6799,N_3473,N_2879);
nor U6800 (N_6800,N_3150,N_4971);
or U6801 (N_6801,N_3906,N_4393);
nand U6802 (N_6802,N_3892,N_2671);
or U6803 (N_6803,N_4885,N_3487);
nor U6804 (N_6804,N_4890,N_4721);
nor U6805 (N_6805,N_3609,N_3418);
nand U6806 (N_6806,N_2705,N_3894);
or U6807 (N_6807,N_3732,N_3409);
and U6808 (N_6808,N_4836,N_4744);
or U6809 (N_6809,N_3464,N_2997);
or U6810 (N_6810,N_4946,N_3016);
nor U6811 (N_6811,N_4903,N_3532);
nand U6812 (N_6812,N_4318,N_3481);
nor U6813 (N_6813,N_4203,N_3506);
or U6814 (N_6814,N_2963,N_3914);
or U6815 (N_6815,N_3026,N_3621);
or U6816 (N_6816,N_4877,N_3989);
or U6817 (N_6817,N_4383,N_3366);
or U6818 (N_6818,N_4375,N_2574);
xnor U6819 (N_6819,N_3584,N_3102);
or U6820 (N_6820,N_3843,N_4775);
xnor U6821 (N_6821,N_4774,N_4093);
xnor U6822 (N_6822,N_4972,N_2770);
xor U6823 (N_6823,N_4961,N_4913);
or U6824 (N_6824,N_3954,N_2644);
and U6825 (N_6825,N_4609,N_3477);
and U6826 (N_6826,N_4161,N_3511);
and U6827 (N_6827,N_4897,N_3534);
or U6828 (N_6828,N_3006,N_4906);
and U6829 (N_6829,N_4015,N_3217);
or U6830 (N_6830,N_4969,N_3126);
nor U6831 (N_6831,N_4944,N_3393);
nor U6832 (N_6832,N_3380,N_3991);
xor U6833 (N_6833,N_4172,N_3432);
nand U6834 (N_6834,N_4482,N_4270);
nor U6835 (N_6835,N_4512,N_4186);
or U6836 (N_6836,N_4498,N_4601);
or U6837 (N_6837,N_3962,N_4869);
nor U6838 (N_6838,N_2670,N_3096);
and U6839 (N_6839,N_3393,N_4312);
and U6840 (N_6840,N_3818,N_2670);
and U6841 (N_6841,N_2974,N_2803);
nand U6842 (N_6842,N_2969,N_3429);
nand U6843 (N_6843,N_2524,N_3680);
nand U6844 (N_6844,N_2543,N_4915);
nand U6845 (N_6845,N_4568,N_2508);
or U6846 (N_6846,N_4257,N_3382);
and U6847 (N_6847,N_4137,N_3106);
nor U6848 (N_6848,N_3466,N_4398);
and U6849 (N_6849,N_3128,N_3612);
and U6850 (N_6850,N_3091,N_4584);
nor U6851 (N_6851,N_3129,N_3347);
nor U6852 (N_6852,N_2846,N_4091);
or U6853 (N_6853,N_4625,N_2979);
or U6854 (N_6854,N_3833,N_3059);
or U6855 (N_6855,N_2961,N_3807);
nand U6856 (N_6856,N_2764,N_4940);
or U6857 (N_6857,N_4624,N_3714);
and U6858 (N_6858,N_4971,N_4695);
nand U6859 (N_6859,N_3718,N_2645);
xor U6860 (N_6860,N_4655,N_4543);
xnor U6861 (N_6861,N_3785,N_4087);
nor U6862 (N_6862,N_3405,N_3222);
nor U6863 (N_6863,N_4133,N_4554);
nand U6864 (N_6864,N_3618,N_3836);
and U6865 (N_6865,N_4442,N_4584);
nor U6866 (N_6866,N_4372,N_4172);
or U6867 (N_6867,N_4519,N_4289);
nand U6868 (N_6868,N_4602,N_4438);
and U6869 (N_6869,N_3420,N_4921);
or U6870 (N_6870,N_4001,N_4570);
and U6871 (N_6871,N_4273,N_3351);
and U6872 (N_6872,N_2738,N_3345);
nor U6873 (N_6873,N_3637,N_3222);
xor U6874 (N_6874,N_3230,N_3961);
and U6875 (N_6875,N_2607,N_2984);
or U6876 (N_6876,N_4984,N_4229);
nand U6877 (N_6877,N_2972,N_4420);
and U6878 (N_6878,N_2933,N_4812);
or U6879 (N_6879,N_3819,N_3519);
and U6880 (N_6880,N_2720,N_3505);
nand U6881 (N_6881,N_4211,N_3002);
nand U6882 (N_6882,N_3242,N_2842);
or U6883 (N_6883,N_3327,N_2913);
nand U6884 (N_6884,N_4368,N_3189);
and U6885 (N_6885,N_4030,N_4053);
xnor U6886 (N_6886,N_3729,N_3217);
nor U6887 (N_6887,N_3785,N_3649);
xor U6888 (N_6888,N_4728,N_3811);
nand U6889 (N_6889,N_2808,N_2992);
or U6890 (N_6890,N_4660,N_2774);
nand U6891 (N_6891,N_3014,N_3095);
or U6892 (N_6892,N_2527,N_2846);
nand U6893 (N_6893,N_3449,N_3063);
or U6894 (N_6894,N_2926,N_4372);
and U6895 (N_6895,N_3575,N_2984);
and U6896 (N_6896,N_3835,N_4768);
nand U6897 (N_6897,N_3639,N_4667);
nor U6898 (N_6898,N_4408,N_3188);
and U6899 (N_6899,N_3252,N_3241);
nand U6900 (N_6900,N_3457,N_4438);
xor U6901 (N_6901,N_4786,N_2505);
or U6902 (N_6902,N_3720,N_3281);
nand U6903 (N_6903,N_3234,N_4065);
and U6904 (N_6904,N_4300,N_2859);
nand U6905 (N_6905,N_3955,N_3381);
nand U6906 (N_6906,N_3285,N_3186);
nor U6907 (N_6907,N_2562,N_4570);
and U6908 (N_6908,N_2541,N_4864);
or U6909 (N_6909,N_2529,N_3196);
or U6910 (N_6910,N_3498,N_4600);
or U6911 (N_6911,N_4849,N_4538);
nor U6912 (N_6912,N_4283,N_3254);
xnor U6913 (N_6913,N_4808,N_4663);
nand U6914 (N_6914,N_2550,N_3782);
nand U6915 (N_6915,N_2790,N_4120);
nor U6916 (N_6916,N_3084,N_3248);
and U6917 (N_6917,N_3713,N_3079);
nand U6918 (N_6918,N_2501,N_3619);
xnor U6919 (N_6919,N_2546,N_4251);
and U6920 (N_6920,N_2780,N_3395);
nand U6921 (N_6921,N_4506,N_3997);
and U6922 (N_6922,N_3517,N_3692);
xnor U6923 (N_6923,N_3897,N_2987);
xor U6924 (N_6924,N_2757,N_3738);
nor U6925 (N_6925,N_2524,N_4487);
or U6926 (N_6926,N_3019,N_3597);
nand U6927 (N_6927,N_2911,N_4381);
or U6928 (N_6928,N_3220,N_2944);
and U6929 (N_6929,N_3010,N_4572);
or U6930 (N_6930,N_4862,N_2991);
or U6931 (N_6931,N_3510,N_2592);
and U6932 (N_6932,N_3561,N_4939);
and U6933 (N_6933,N_4091,N_3063);
and U6934 (N_6934,N_4875,N_3005);
nor U6935 (N_6935,N_4370,N_3595);
nor U6936 (N_6936,N_3900,N_4800);
and U6937 (N_6937,N_4184,N_4937);
and U6938 (N_6938,N_3615,N_3737);
nand U6939 (N_6939,N_4749,N_2807);
or U6940 (N_6940,N_3174,N_4392);
xor U6941 (N_6941,N_4364,N_4166);
nand U6942 (N_6942,N_2816,N_4806);
xnor U6943 (N_6943,N_3292,N_3198);
or U6944 (N_6944,N_4539,N_4027);
or U6945 (N_6945,N_4696,N_4844);
xnor U6946 (N_6946,N_2540,N_3552);
nor U6947 (N_6947,N_4555,N_4312);
xor U6948 (N_6948,N_3193,N_3772);
and U6949 (N_6949,N_4314,N_2755);
xnor U6950 (N_6950,N_3262,N_4009);
nor U6951 (N_6951,N_2742,N_4688);
nor U6952 (N_6952,N_4619,N_4755);
or U6953 (N_6953,N_4412,N_4061);
nand U6954 (N_6954,N_3786,N_4056);
xor U6955 (N_6955,N_3680,N_3259);
and U6956 (N_6956,N_2571,N_3062);
or U6957 (N_6957,N_3529,N_2807);
nor U6958 (N_6958,N_3148,N_4816);
or U6959 (N_6959,N_4925,N_4547);
and U6960 (N_6960,N_2693,N_4490);
nand U6961 (N_6961,N_2522,N_2561);
or U6962 (N_6962,N_2625,N_3653);
nor U6963 (N_6963,N_3312,N_3532);
and U6964 (N_6964,N_3634,N_3323);
nand U6965 (N_6965,N_4638,N_3291);
nand U6966 (N_6966,N_3004,N_4240);
nand U6967 (N_6967,N_2979,N_2742);
xnor U6968 (N_6968,N_3471,N_4991);
or U6969 (N_6969,N_4417,N_4978);
nand U6970 (N_6970,N_4644,N_4198);
nand U6971 (N_6971,N_4152,N_2720);
and U6972 (N_6972,N_3357,N_3401);
or U6973 (N_6973,N_3477,N_3770);
xor U6974 (N_6974,N_3369,N_4890);
and U6975 (N_6975,N_2986,N_2592);
nand U6976 (N_6976,N_4473,N_4048);
or U6977 (N_6977,N_3369,N_3958);
or U6978 (N_6978,N_4508,N_4500);
and U6979 (N_6979,N_3554,N_3943);
or U6980 (N_6980,N_4754,N_4850);
nor U6981 (N_6981,N_3691,N_4283);
nand U6982 (N_6982,N_2764,N_2599);
xnor U6983 (N_6983,N_4096,N_4477);
and U6984 (N_6984,N_4503,N_3747);
nand U6985 (N_6985,N_4319,N_4519);
nand U6986 (N_6986,N_3980,N_3110);
nor U6987 (N_6987,N_3773,N_3122);
or U6988 (N_6988,N_4066,N_4750);
nand U6989 (N_6989,N_2573,N_4861);
and U6990 (N_6990,N_3710,N_3531);
or U6991 (N_6991,N_3196,N_2724);
or U6992 (N_6992,N_2797,N_4171);
nand U6993 (N_6993,N_2740,N_4613);
xnor U6994 (N_6994,N_4353,N_2646);
nand U6995 (N_6995,N_3307,N_4904);
and U6996 (N_6996,N_2555,N_4970);
or U6997 (N_6997,N_3064,N_3737);
nor U6998 (N_6998,N_3722,N_3435);
or U6999 (N_6999,N_4425,N_4633);
xnor U7000 (N_7000,N_2962,N_4405);
nor U7001 (N_7001,N_4446,N_4404);
or U7002 (N_7002,N_4160,N_4777);
nor U7003 (N_7003,N_3166,N_2849);
and U7004 (N_7004,N_3046,N_4735);
xnor U7005 (N_7005,N_4628,N_2937);
and U7006 (N_7006,N_2519,N_3000);
and U7007 (N_7007,N_4956,N_3709);
nor U7008 (N_7008,N_3366,N_3205);
or U7009 (N_7009,N_3588,N_3478);
nand U7010 (N_7010,N_4468,N_4711);
nor U7011 (N_7011,N_4811,N_3732);
or U7012 (N_7012,N_4176,N_2672);
or U7013 (N_7013,N_3760,N_2962);
xnor U7014 (N_7014,N_2819,N_4632);
xor U7015 (N_7015,N_3818,N_4606);
nor U7016 (N_7016,N_3075,N_4784);
and U7017 (N_7017,N_2817,N_4361);
nor U7018 (N_7018,N_4920,N_3065);
xnor U7019 (N_7019,N_2556,N_3816);
nand U7020 (N_7020,N_4554,N_4650);
or U7021 (N_7021,N_3864,N_3535);
or U7022 (N_7022,N_4445,N_3643);
nor U7023 (N_7023,N_4500,N_4245);
nor U7024 (N_7024,N_3909,N_4664);
nor U7025 (N_7025,N_3480,N_2545);
and U7026 (N_7026,N_3972,N_4499);
xor U7027 (N_7027,N_3757,N_2776);
and U7028 (N_7028,N_4963,N_2630);
nand U7029 (N_7029,N_4908,N_2628);
xor U7030 (N_7030,N_2909,N_3660);
nand U7031 (N_7031,N_4680,N_4457);
nor U7032 (N_7032,N_4519,N_4738);
and U7033 (N_7033,N_4768,N_3257);
and U7034 (N_7034,N_3094,N_4739);
and U7035 (N_7035,N_4256,N_4875);
and U7036 (N_7036,N_2706,N_3481);
and U7037 (N_7037,N_2689,N_2749);
and U7038 (N_7038,N_3590,N_4975);
nand U7039 (N_7039,N_4090,N_4216);
nor U7040 (N_7040,N_4013,N_4204);
nand U7041 (N_7041,N_2659,N_3667);
or U7042 (N_7042,N_4660,N_4811);
or U7043 (N_7043,N_4341,N_2705);
nor U7044 (N_7044,N_4898,N_4198);
nand U7045 (N_7045,N_4811,N_3576);
or U7046 (N_7046,N_2854,N_3951);
and U7047 (N_7047,N_3029,N_3031);
nor U7048 (N_7048,N_3285,N_4270);
nand U7049 (N_7049,N_4593,N_3671);
and U7050 (N_7050,N_4834,N_3004);
and U7051 (N_7051,N_3009,N_3040);
nor U7052 (N_7052,N_4133,N_4083);
nor U7053 (N_7053,N_4798,N_2608);
nor U7054 (N_7054,N_3533,N_4761);
and U7055 (N_7055,N_3367,N_4061);
or U7056 (N_7056,N_4224,N_4569);
or U7057 (N_7057,N_3027,N_3558);
or U7058 (N_7058,N_3434,N_2997);
nand U7059 (N_7059,N_3169,N_3635);
and U7060 (N_7060,N_2896,N_4589);
nor U7061 (N_7061,N_3989,N_4723);
nand U7062 (N_7062,N_3723,N_3087);
nor U7063 (N_7063,N_4296,N_2823);
nor U7064 (N_7064,N_3466,N_2573);
and U7065 (N_7065,N_3333,N_3572);
nor U7066 (N_7066,N_4727,N_3067);
nor U7067 (N_7067,N_3469,N_2826);
and U7068 (N_7068,N_3013,N_2733);
nand U7069 (N_7069,N_4207,N_2567);
nand U7070 (N_7070,N_4560,N_4542);
nand U7071 (N_7071,N_3678,N_4187);
nand U7072 (N_7072,N_4399,N_3246);
nand U7073 (N_7073,N_4781,N_4821);
or U7074 (N_7074,N_2939,N_3276);
nand U7075 (N_7075,N_3127,N_3062);
nor U7076 (N_7076,N_3177,N_4214);
nor U7077 (N_7077,N_3582,N_4277);
and U7078 (N_7078,N_4797,N_3838);
nand U7079 (N_7079,N_4011,N_4791);
and U7080 (N_7080,N_3805,N_2799);
or U7081 (N_7081,N_4969,N_3812);
nor U7082 (N_7082,N_2863,N_3167);
nor U7083 (N_7083,N_3403,N_4468);
nor U7084 (N_7084,N_4778,N_2945);
and U7085 (N_7085,N_3230,N_4202);
xor U7086 (N_7086,N_3750,N_4528);
and U7087 (N_7087,N_3966,N_3450);
or U7088 (N_7088,N_2743,N_2728);
nor U7089 (N_7089,N_3351,N_4469);
nand U7090 (N_7090,N_2907,N_4598);
nand U7091 (N_7091,N_3268,N_3693);
or U7092 (N_7092,N_4268,N_3644);
or U7093 (N_7093,N_4185,N_4120);
nand U7094 (N_7094,N_3843,N_3529);
nand U7095 (N_7095,N_2595,N_3250);
and U7096 (N_7096,N_3907,N_4138);
nand U7097 (N_7097,N_3967,N_3276);
and U7098 (N_7098,N_2758,N_4730);
nand U7099 (N_7099,N_4301,N_4950);
nor U7100 (N_7100,N_3521,N_3357);
xnor U7101 (N_7101,N_2705,N_3149);
nand U7102 (N_7102,N_4303,N_3319);
and U7103 (N_7103,N_2513,N_3732);
nand U7104 (N_7104,N_4741,N_3559);
nand U7105 (N_7105,N_3999,N_3560);
xnor U7106 (N_7106,N_3885,N_4685);
and U7107 (N_7107,N_3534,N_4407);
xor U7108 (N_7108,N_4867,N_2571);
nor U7109 (N_7109,N_4926,N_2839);
nor U7110 (N_7110,N_2924,N_3843);
and U7111 (N_7111,N_3429,N_3440);
or U7112 (N_7112,N_3108,N_3637);
xnor U7113 (N_7113,N_2674,N_3583);
or U7114 (N_7114,N_3827,N_3812);
nand U7115 (N_7115,N_2772,N_2892);
and U7116 (N_7116,N_4807,N_2921);
and U7117 (N_7117,N_4838,N_3743);
and U7118 (N_7118,N_3098,N_4331);
nand U7119 (N_7119,N_2551,N_3627);
and U7120 (N_7120,N_4849,N_4559);
and U7121 (N_7121,N_3131,N_3995);
or U7122 (N_7122,N_4626,N_4327);
nand U7123 (N_7123,N_3150,N_3351);
and U7124 (N_7124,N_3827,N_3990);
xor U7125 (N_7125,N_3012,N_4792);
and U7126 (N_7126,N_2970,N_2986);
nand U7127 (N_7127,N_3854,N_3340);
or U7128 (N_7128,N_2684,N_3116);
nand U7129 (N_7129,N_3667,N_2716);
xor U7130 (N_7130,N_4483,N_4523);
nand U7131 (N_7131,N_2940,N_4494);
or U7132 (N_7132,N_3775,N_3072);
nand U7133 (N_7133,N_4173,N_4981);
nor U7134 (N_7134,N_4675,N_2576);
nand U7135 (N_7135,N_4299,N_3192);
nand U7136 (N_7136,N_3590,N_4841);
nor U7137 (N_7137,N_3707,N_4640);
or U7138 (N_7138,N_4432,N_4877);
nor U7139 (N_7139,N_3881,N_2509);
or U7140 (N_7140,N_4734,N_3513);
nand U7141 (N_7141,N_4342,N_4791);
or U7142 (N_7142,N_4185,N_2887);
or U7143 (N_7143,N_2733,N_3976);
or U7144 (N_7144,N_4610,N_3892);
or U7145 (N_7145,N_2951,N_3587);
nand U7146 (N_7146,N_2701,N_3130);
xor U7147 (N_7147,N_3200,N_3925);
nor U7148 (N_7148,N_4336,N_4482);
or U7149 (N_7149,N_3766,N_3187);
nor U7150 (N_7150,N_3008,N_3272);
and U7151 (N_7151,N_4327,N_2909);
and U7152 (N_7152,N_4873,N_4749);
xnor U7153 (N_7153,N_2755,N_3975);
and U7154 (N_7154,N_3532,N_3398);
nand U7155 (N_7155,N_4277,N_4862);
xnor U7156 (N_7156,N_3219,N_4179);
or U7157 (N_7157,N_3968,N_4008);
nand U7158 (N_7158,N_3888,N_2566);
nor U7159 (N_7159,N_4071,N_2826);
or U7160 (N_7160,N_2662,N_4018);
and U7161 (N_7161,N_4150,N_4128);
or U7162 (N_7162,N_4539,N_3752);
or U7163 (N_7163,N_4000,N_3132);
nand U7164 (N_7164,N_4046,N_4432);
nand U7165 (N_7165,N_4908,N_4744);
nor U7166 (N_7166,N_3466,N_3718);
or U7167 (N_7167,N_3228,N_2837);
nand U7168 (N_7168,N_4772,N_3688);
xnor U7169 (N_7169,N_4022,N_2800);
nor U7170 (N_7170,N_2740,N_2877);
nor U7171 (N_7171,N_3782,N_4699);
or U7172 (N_7172,N_4351,N_3471);
nor U7173 (N_7173,N_3395,N_3983);
and U7174 (N_7174,N_2511,N_2586);
nor U7175 (N_7175,N_3494,N_2535);
nor U7176 (N_7176,N_4715,N_4053);
and U7177 (N_7177,N_3336,N_3461);
and U7178 (N_7178,N_3669,N_2758);
and U7179 (N_7179,N_2550,N_4033);
or U7180 (N_7180,N_4071,N_3691);
nor U7181 (N_7181,N_2714,N_2922);
nand U7182 (N_7182,N_3679,N_4008);
and U7183 (N_7183,N_3529,N_2577);
nor U7184 (N_7184,N_4333,N_3964);
or U7185 (N_7185,N_3737,N_4381);
nor U7186 (N_7186,N_4136,N_4248);
and U7187 (N_7187,N_2851,N_2625);
or U7188 (N_7188,N_3196,N_3515);
or U7189 (N_7189,N_3441,N_4259);
or U7190 (N_7190,N_3063,N_2963);
xor U7191 (N_7191,N_4598,N_2577);
or U7192 (N_7192,N_4887,N_4922);
and U7193 (N_7193,N_2916,N_2687);
nor U7194 (N_7194,N_3182,N_3971);
nand U7195 (N_7195,N_3375,N_2895);
and U7196 (N_7196,N_2698,N_4587);
or U7197 (N_7197,N_3044,N_2926);
or U7198 (N_7198,N_4258,N_3702);
nand U7199 (N_7199,N_3416,N_3189);
nor U7200 (N_7200,N_3609,N_4697);
and U7201 (N_7201,N_3056,N_4260);
and U7202 (N_7202,N_4758,N_2521);
or U7203 (N_7203,N_4446,N_3005);
or U7204 (N_7204,N_3082,N_3058);
xnor U7205 (N_7205,N_4113,N_2908);
nor U7206 (N_7206,N_4206,N_2590);
nand U7207 (N_7207,N_3684,N_3920);
nor U7208 (N_7208,N_3897,N_2757);
nand U7209 (N_7209,N_3090,N_4560);
or U7210 (N_7210,N_3085,N_2734);
or U7211 (N_7211,N_4283,N_3152);
nor U7212 (N_7212,N_4466,N_3191);
nand U7213 (N_7213,N_4516,N_4486);
nor U7214 (N_7214,N_4357,N_3732);
or U7215 (N_7215,N_3132,N_4296);
or U7216 (N_7216,N_4954,N_2852);
nand U7217 (N_7217,N_4787,N_4690);
and U7218 (N_7218,N_4962,N_2737);
or U7219 (N_7219,N_2554,N_4488);
xnor U7220 (N_7220,N_2508,N_3453);
or U7221 (N_7221,N_2524,N_3481);
and U7222 (N_7222,N_2761,N_2668);
or U7223 (N_7223,N_4821,N_4863);
or U7224 (N_7224,N_3277,N_2589);
or U7225 (N_7225,N_4597,N_4937);
xnor U7226 (N_7226,N_3875,N_4445);
and U7227 (N_7227,N_2758,N_4889);
nand U7228 (N_7228,N_4540,N_2764);
or U7229 (N_7229,N_4853,N_2668);
nor U7230 (N_7230,N_4439,N_3403);
xor U7231 (N_7231,N_3692,N_3218);
nand U7232 (N_7232,N_4031,N_4835);
nand U7233 (N_7233,N_3154,N_3302);
nand U7234 (N_7234,N_4685,N_2786);
or U7235 (N_7235,N_3090,N_3028);
nor U7236 (N_7236,N_3367,N_4983);
nor U7237 (N_7237,N_4975,N_4309);
nand U7238 (N_7238,N_3315,N_4390);
nand U7239 (N_7239,N_4593,N_4402);
and U7240 (N_7240,N_3084,N_3453);
nand U7241 (N_7241,N_2793,N_4458);
or U7242 (N_7242,N_3647,N_3007);
xnor U7243 (N_7243,N_4165,N_3871);
xor U7244 (N_7244,N_4260,N_4459);
xor U7245 (N_7245,N_2568,N_2753);
nor U7246 (N_7246,N_4372,N_2901);
or U7247 (N_7247,N_2818,N_4119);
nand U7248 (N_7248,N_3265,N_4943);
or U7249 (N_7249,N_4960,N_3067);
or U7250 (N_7250,N_4982,N_4772);
xnor U7251 (N_7251,N_4979,N_2944);
nand U7252 (N_7252,N_3157,N_2668);
or U7253 (N_7253,N_2650,N_4046);
or U7254 (N_7254,N_4872,N_3065);
and U7255 (N_7255,N_3664,N_3598);
or U7256 (N_7256,N_4667,N_4162);
nor U7257 (N_7257,N_3940,N_4207);
nor U7258 (N_7258,N_3691,N_4487);
xor U7259 (N_7259,N_3130,N_3417);
xnor U7260 (N_7260,N_2995,N_3252);
nand U7261 (N_7261,N_3211,N_3934);
and U7262 (N_7262,N_3849,N_4437);
or U7263 (N_7263,N_3254,N_4806);
nor U7264 (N_7264,N_4785,N_4239);
xor U7265 (N_7265,N_2778,N_4098);
or U7266 (N_7266,N_4485,N_3477);
or U7267 (N_7267,N_2891,N_4645);
nand U7268 (N_7268,N_4489,N_3686);
and U7269 (N_7269,N_4526,N_2708);
or U7270 (N_7270,N_3162,N_4581);
and U7271 (N_7271,N_2579,N_3022);
nor U7272 (N_7272,N_2930,N_4228);
nand U7273 (N_7273,N_3894,N_3610);
nor U7274 (N_7274,N_4091,N_3830);
nor U7275 (N_7275,N_2798,N_3670);
or U7276 (N_7276,N_4298,N_2918);
nor U7277 (N_7277,N_4019,N_2502);
xor U7278 (N_7278,N_3570,N_4138);
xor U7279 (N_7279,N_3585,N_4968);
and U7280 (N_7280,N_2559,N_3402);
nor U7281 (N_7281,N_3766,N_2796);
or U7282 (N_7282,N_3904,N_4268);
and U7283 (N_7283,N_3777,N_2772);
or U7284 (N_7284,N_2529,N_3312);
xnor U7285 (N_7285,N_2855,N_2819);
or U7286 (N_7286,N_2568,N_3933);
xnor U7287 (N_7287,N_4912,N_2790);
or U7288 (N_7288,N_4653,N_3836);
nand U7289 (N_7289,N_3542,N_3319);
or U7290 (N_7290,N_4257,N_4612);
and U7291 (N_7291,N_3435,N_4033);
nor U7292 (N_7292,N_3888,N_3926);
nand U7293 (N_7293,N_4126,N_2816);
xnor U7294 (N_7294,N_3203,N_4679);
and U7295 (N_7295,N_4410,N_3209);
xnor U7296 (N_7296,N_4391,N_4359);
nor U7297 (N_7297,N_4862,N_2968);
and U7298 (N_7298,N_4599,N_3754);
and U7299 (N_7299,N_4740,N_3956);
nand U7300 (N_7300,N_3394,N_2776);
nand U7301 (N_7301,N_2982,N_4014);
or U7302 (N_7302,N_2572,N_2586);
or U7303 (N_7303,N_4617,N_3894);
xor U7304 (N_7304,N_2817,N_3977);
nor U7305 (N_7305,N_4178,N_3050);
xor U7306 (N_7306,N_4126,N_2946);
nand U7307 (N_7307,N_2923,N_3384);
and U7308 (N_7308,N_3195,N_3911);
or U7309 (N_7309,N_4223,N_4822);
xor U7310 (N_7310,N_4488,N_4393);
or U7311 (N_7311,N_2994,N_4666);
nand U7312 (N_7312,N_4566,N_3259);
or U7313 (N_7313,N_3280,N_3815);
nand U7314 (N_7314,N_3533,N_2530);
nor U7315 (N_7315,N_4390,N_3748);
and U7316 (N_7316,N_4076,N_3650);
and U7317 (N_7317,N_2764,N_4416);
and U7318 (N_7318,N_3749,N_4899);
nor U7319 (N_7319,N_4125,N_4307);
xor U7320 (N_7320,N_4835,N_4006);
nand U7321 (N_7321,N_2689,N_3987);
or U7322 (N_7322,N_3914,N_4971);
and U7323 (N_7323,N_4745,N_4307);
and U7324 (N_7324,N_2977,N_2685);
nand U7325 (N_7325,N_4566,N_3367);
or U7326 (N_7326,N_3262,N_3926);
or U7327 (N_7327,N_4838,N_4917);
or U7328 (N_7328,N_4536,N_4723);
nor U7329 (N_7329,N_4349,N_4208);
nand U7330 (N_7330,N_4870,N_3515);
nand U7331 (N_7331,N_4219,N_4474);
nor U7332 (N_7332,N_3196,N_2837);
nand U7333 (N_7333,N_2927,N_4905);
and U7334 (N_7334,N_3546,N_4960);
nand U7335 (N_7335,N_2609,N_2748);
nand U7336 (N_7336,N_4297,N_2992);
or U7337 (N_7337,N_3024,N_3744);
nor U7338 (N_7338,N_2732,N_3658);
and U7339 (N_7339,N_4533,N_2679);
nand U7340 (N_7340,N_4839,N_2923);
nand U7341 (N_7341,N_3649,N_3339);
nand U7342 (N_7342,N_4919,N_4902);
nand U7343 (N_7343,N_2811,N_3620);
nor U7344 (N_7344,N_4385,N_4106);
and U7345 (N_7345,N_3860,N_4747);
or U7346 (N_7346,N_4955,N_3665);
nand U7347 (N_7347,N_4469,N_3458);
or U7348 (N_7348,N_4456,N_3986);
and U7349 (N_7349,N_4710,N_4321);
xor U7350 (N_7350,N_3071,N_4366);
nand U7351 (N_7351,N_4041,N_3801);
xnor U7352 (N_7352,N_2990,N_3858);
or U7353 (N_7353,N_2811,N_3721);
or U7354 (N_7354,N_3571,N_3160);
or U7355 (N_7355,N_2803,N_4126);
nor U7356 (N_7356,N_3094,N_2732);
and U7357 (N_7357,N_3483,N_4198);
nor U7358 (N_7358,N_4558,N_3948);
or U7359 (N_7359,N_4500,N_4591);
nor U7360 (N_7360,N_4351,N_3795);
nand U7361 (N_7361,N_3077,N_3121);
nor U7362 (N_7362,N_2753,N_4989);
and U7363 (N_7363,N_4398,N_3486);
nor U7364 (N_7364,N_4498,N_3888);
nor U7365 (N_7365,N_3077,N_4888);
nor U7366 (N_7366,N_4108,N_4732);
and U7367 (N_7367,N_4140,N_2611);
nor U7368 (N_7368,N_4130,N_4494);
and U7369 (N_7369,N_2683,N_3650);
nand U7370 (N_7370,N_3039,N_3455);
and U7371 (N_7371,N_4587,N_2870);
or U7372 (N_7372,N_2550,N_4346);
nand U7373 (N_7373,N_3201,N_2993);
xnor U7374 (N_7374,N_2965,N_4922);
xor U7375 (N_7375,N_4398,N_2704);
nand U7376 (N_7376,N_2794,N_3954);
nand U7377 (N_7377,N_4586,N_3445);
nand U7378 (N_7378,N_4527,N_3167);
and U7379 (N_7379,N_3389,N_3858);
and U7380 (N_7380,N_2987,N_3900);
nand U7381 (N_7381,N_4020,N_4527);
or U7382 (N_7382,N_4138,N_2784);
or U7383 (N_7383,N_4545,N_4266);
or U7384 (N_7384,N_4194,N_2945);
xor U7385 (N_7385,N_2580,N_2594);
or U7386 (N_7386,N_3675,N_2560);
nand U7387 (N_7387,N_3673,N_4093);
or U7388 (N_7388,N_4576,N_3801);
and U7389 (N_7389,N_4178,N_3416);
nor U7390 (N_7390,N_4326,N_2510);
nand U7391 (N_7391,N_4874,N_4531);
or U7392 (N_7392,N_3898,N_4141);
nor U7393 (N_7393,N_4501,N_3237);
or U7394 (N_7394,N_4750,N_3640);
nand U7395 (N_7395,N_3581,N_3087);
or U7396 (N_7396,N_2638,N_3436);
or U7397 (N_7397,N_4584,N_4650);
xor U7398 (N_7398,N_3619,N_4100);
nor U7399 (N_7399,N_4096,N_4752);
nor U7400 (N_7400,N_3136,N_3793);
nand U7401 (N_7401,N_2882,N_3916);
nand U7402 (N_7402,N_3786,N_3517);
nor U7403 (N_7403,N_4023,N_4540);
nand U7404 (N_7404,N_4364,N_3682);
or U7405 (N_7405,N_2890,N_3897);
nand U7406 (N_7406,N_4111,N_4305);
and U7407 (N_7407,N_3690,N_4042);
nand U7408 (N_7408,N_3775,N_2901);
and U7409 (N_7409,N_2858,N_4349);
or U7410 (N_7410,N_4823,N_3653);
or U7411 (N_7411,N_3003,N_4481);
nand U7412 (N_7412,N_3730,N_4028);
nor U7413 (N_7413,N_3054,N_4013);
and U7414 (N_7414,N_4374,N_4973);
or U7415 (N_7415,N_3817,N_4849);
and U7416 (N_7416,N_3936,N_3908);
nor U7417 (N_7417,N_3343,N_4550);
nor U7418 (N_7418,N_2750,N_4775);
or U7419 (N_7419,N_3317,N_4924);
xor U7420 (N_7420,N_3028,N_3477);
nand U7421 (N_7421,N_2575,N_3470);
or U7422 (N_7422,N_3244,N_4053);
nand U7423 (N_7423,N_3404,N_2846);
nor U7424 (N_7424,N_3500,N_3290);
and U7425 (N_7425,N_3088,N_3138);
nor U7426 (N_7426,N_3297,N_3972);
nand U7427 (N_7427,N_2857,N_3320);
and U7428 (N_7428,N_3717,N_3920);
nor U7429 (N_7429,N_4378,N_4299);
and U7430 (N_7430,N_4094,N_4487);
and U7431 (N_7431,N_3657,N_4632);
and U7432 (N_7432,N_3077,N_3830);
nand U7433 (N_7433,N_4099,N_3901);
nor U7434 (N_7434,N_2899,N_3322);
nor U7435 (N_7435,N_4215,N_4183);
xnor U7436 (N_7436,N_4089,N_3897);
nand U7437 (N_7437,N_3765,N_4742);
nand U7438 (N_7438,N_3038,N_4002);
or U7439 (N_7439,N_4666,N_3716);
nor U7440 (N_7440,N_3070,N_2814);
xnor U7441 (N_7441,N_4690,N_4242);
nand U7442 (N_7442,N_3487,N_3643);
xor U7443 (N_7443,N_2681,N_3909);
nor U7444 (N_7444,N_4558,N_2774);
and U7445 (N_7445,N_2799,N_2671);
or U7446 (N_7446,N_2911,N_2750);
and U7447 (N_7447,N_2970,N_3698);
or U7448 (N_7448,N_2579,N_3547);
nor U7449 (N_7449,N_3817,N_4703);
or U7450 (N_7450,N_4691,N_4475);
nor U7451 (N_7451,N_3061,N_4048);
and U7452 (N_7452,N_4295,N_4103);
and U7453 (N_7453,N_2794,N_4904);
nor U7454 (N_7454,N_4256,N_3512);
nand U7455 (N_7455,N_4380,N_3306);
and U7456 (N_7456,N_4616,N_3168);
or U7457 (N_7457,N_4106,N_2639);
and U7458 (N_7458,N_3007,N_4693);
and U7459 (N_7459,N_4752,N_4005);
nand U7460 (N_7460,N_3195,N_4696);
nor U7461 (N_7461,N_4894,N_4495);
nand U7462 (N_7462,N_3423,N_3504);
nor U7463 (N_7463,N_4043,N_4028);
and U7464 (N_7464,N_4825,N_4893);
and U7465 (N_7465,N_2914,N_3201);
or U7466 (N_7466,N_2737,N_4400);
nand U7467 (N_7467,N_3828,N_4134);
nand U7468 (N_7468,N_2976,N_3291);
and U7469 (N_7469,N_3070,N_3646);
xnor U7470 (N_7470,N_4999,N_2546);
or U7471 (N_7471,N_3071,N_3380);
nand U7472 (N_7472,N_4437,N_3605);
or U7473 (N_7473,N_3921,N_3787);
and U7474 (N_7474,N_4831,N_3443);
nor U7475 (N_7475,N_4194,N_3702);
nor U7476 (N_7476,N_4827,N_3109);
nor U7477 (N_7477,N_4468,N_3423);
and U7478 (N_7478,N_3746,N_4098);
and U7479 (N_7479,N_4011,N_3858);
or U7480 (N_7480,N_3029,N_2899);
or U7481 (N_7481,N_3479,N_3005);
nor U7482 (N_7482,N_3732,N_3334);
nand U7483 (N_7483,N_4464,N_3619);
nor U7484 (N_7484,N_4935,N_2893);
nor U7485 (N_7485,N_2672,N_2938);
or U7486 (N_7486,N_2726,N_2853);
or U7487 (N_7487,N_3036,N_3026);
nand U7488 (N_7488,N_4928,N_4097);
or U7489 (N_7489,N_4089,N_4327);
nor U7490 (N_7490,N_2713,N_2816);
or U7491 (N_7491,N_2938,N_3080);
or U7492 (N_7492,N_3946,N_2973);
nand U7493 (N_7493,N_4010,N_4815);
xor U7494 (N_7494,N_4754,N_2507);
and U7495 (N_7495,N_4864,N_4291);
nand U7496 (N_7496,N_4755,N_3856);
nand U7497 (N_7497,N_3701,N_3757);
or U7498 (N_7498,N_3254,N_3592);
xnor U7499 (N_7499,N_4284,N_4447);
nand U7500 (N_7500,N_6322,N_7250);
xor U7501 (N_7501,N_7104,N_6925);
nand U7502 (N_7502,N_5792,N_6977);
nor U7503 (N_7503,N_5812,N_6495);
or U7504 (N_7504,N_7024,N_5154);
or U7505 (N_7505,N_5900,N_6484);
nor U7506 (N_7506,N_6889,N_6671);
and U7507 (N_7507,N_6319,N_5361);
nor U7508 (N_7508,N_5916,N_6173);
xnor U7509 (N_7509,N_7483,N_6140);
nor U7510 (N_7510,N_6865,N_7429);
nand U7511 (N_7511,N_5710,N_6784);
nand U7512 (N_7512,N_6523,N_5715);
nor U7513 (N_7513,N_6618,N_6378);
or U7514 (N_7514,N_7372,N_7439);
and U7515 (N_7515,N_7327,N_7394);
or U7516 (N_7516,N_6046,N_5537);
and U7517 (N_7517,N_6213,N_5991);
nand U7518 (N_7518,N_5031,N_6829);
and U7519 (N_7519,N_7242,N_5511);
or U7520 (N_7520,N_5906,N_5822);
and U7521 (N_7521,N_5249,N_6045);
nand U7522 (N_7522,N_6540,N_5513);
nor U7523 (N_7523,N_5211,N_6556);
and U7524 (N_7524,N_7435,N_6089);
nor U7525 (N_7525,N_7017,N_5394);
nand U7526 (N_7526,N_5516,N_7197);
nand U7527 (N_7527,N_6757,N_6419);
nand U7528 (N_7528,N_5193,N_6962);
nor U7529 (N_7529,N_7166,N_5437);
nand U7530 (N_7530,N_7055,N_6694);
and U7531 (N_7531,N_6225,N_6490);
and U7532 (N_7532,N_6305,N_7345);
nor U7533 (N_7533,N_6166,N_6281);
and U7534 (N_7534,N_6496,N_6760);
and U7535 (N_7535,N_6672,N_5555);
or U7536 (N_7536,N_5178,N_7083);
and U7537 (N_7537,N_7335,N_6425);
xnor U7538 (N_7538,N_5327,N_5163);
or U7539 (N_7539,N_6176,N_5568);
xnor U7540 (N_7540,N_6600,N_5374);
nand U7541 (N_7541,N_6428,N_6786);
or U7542 (N_7542,N_7387,N_6218);
nor U7543 (N_7543,N_7040,N_6666);
nand U7544 (N_7544,N_6697,N_6973);
nand U7545 (N_7545,N_6685,N_5399);
nand U7546 (N_7546,N_6152,N_5586);
nand U7547 (N_7547,N_5821,N_7234);
nand U7548 (N_7548,N_5818,N_5425);
nor U7549 (N_7549,N_6242,N_5848);
nor U7550 (N_7550,N_5451,N_6871);
and U7551 (N_7551,N_5474,N_5306);
and U7552 (N_7552,N_5933,N_6433);
or U7553 (N_7553,N_6071,N_5939);
or U7554 (N_7554,N_6261,N_6082);
nand U7555 (N_7555,N_6588,N_7023);
nor U7556 (N_7556,N_7231,N_5053);
or U7557 (N_7557,N_5096,N_5747);
and U7558 (N_7558,N_5033,N_5109);
and U7559 (N_7559,N_5161,N_6712);
nand U7560 (N_7560,N_6078,N_5532);
xor U7561 (N_7561,N_7337,N_5844);
nand U7562 (N_7562,N_6307,N_5930);
and U7563 (N_7563,N_6640,N_5221);
or U7564 (N_7564,N_6996,N_6407);
xnor U7565 (N_7565,N_7046,N_6581);
nand U7566 (N_7566,N_5722,N_6975);
nand U7567 (N_7567,N_6596,N_5853);
or U7568 (N_7568,N_5379,N_6853);
nand U7569 (N_7569,N_6347,N_5291);
nor U7570 (N_7570,N_6849,N_7299);
and U7571 (N_7571,N_7235,N_5522);
nor U7572 (N_7572,N_6919,N_5423);
or U7573 (N_7573,N_7244,N_6524);
nand U7574 (N_7574,N_7045,N_7262);
or U7575 (N_7575,N_6668,N_7436);
nor U7576 (N_7576,N_7370,N_6563);
nand U7577 (N_7577,N_5799,N_5765);
and U7578 (N_7578,N_5877,N_6498);
nand U7579 (N_7579,N_6435,N_7000);
or U7580 (N_7580,N_7119,N_6793);
nand U7581 (N_7581,N_7216,N_6687);
and U7582 (N_7582,N_5119,N_6650);
and U7583 (N_7583,N_7125,N_6880);
and U7584 (N_7584,N_7034,N_5776);
nor U7585 (N_7585,N_5354,N_5478);
nor U7586 (N_7586,N_6280,N_6591);
xor U7587 (N_7587,N_5226,N_6300);
or U7588 (N_7588,N_5116,N_6177);
or U7589 (N_7589,N_5064,N_5772);
nand U7590 (N_7590,N_6724,N_6288);
or U7591 (N_7591,N_5349,N_5688);
nand U7592 (N_7592,N_6249,N_6284);
and U7593 (N_7593,N_5364,N_5059);
and U7594 (N_7594,N_6681,N_6748);
nand U7595 (N_7595,N_5040,N_6135);
and U7596 (N_7596,N_6903,N_6890);
nor U7597 (N_7597,N_5597,N_7389);
and U7598 (N_7598,N_7332,N_6478);
or U7599 (N_7599,N_6796,N_6172);
nor U7600 (N_7600,N_5131,N_6623);
xnor U7601 (N_7601,N_5655,N_5563);
nand U7602 (N_7602,N_5908,N_6544);
and U7603 (N_7603,N_7316,N_5001);
and U7604 (N_7604,N_6874,N_6682);
or U7605 (N_7605,N_7217,N_5144);
or U7606 (N_7606,N_6129,N_6402);
or U7607 (N_7607,N_6550,N_5248);
or U7608 (N_7608,N_5920,N_6301);
and U7609 (N_7609,N_6103,N_7373);
nor U7610 (N_7610,N_5781,N_5223);
and U7611 (N_7611,N_5443,N_6987);
nand U7612 (N_7612,N_5907,N_6802);
nand U7613 (N_7613,N_7246,N_7494);
nor U7614 (N_7614,N_5889,N_5758);
or U7615 (N_7615,N_6960,N_6018);
nor U7616 (N_7616,N_5703,N_5992);
and U7617 (N_7617,N_6990,N_6616);
and U7618 (N_7618,N_6329,N_6265);
nand U7619 (N_7619,N_5837,N_6233);
nor U7620 (N_7620,N_6891,N_5551);
and U7621 (N_7621,N_6610,N_7012);
nor U7622 (N_7622,N_5460,N_6794);
or U7623 (N_7623,N_6215,N_6223);
and U7624 (N_7624,N_5305,N_7148);
and U7625 (N_7625,N_6426,N_5285);
and U7626 (N_7626,N_5684,N_5525);
or U7627 (N_7627,N_6159,N_6745);
or U7628 (N_7628,N_5762,N_5990);
or U7629 (N_7629,N_6455,N_6287);
xor U7630 (N_7630,N_5442,N_7186);
or U7631 (N_7631,N_6232,N_6959);
nand U7632 (N_7632,N_5069,N_5888);
nor U7633 (N_7633,N_5810,N_5387);
nor U7634 (N_7634,N_6744,N_6943);
xnor U7635 (N_7635,N_7444,N_6612);
nor U7636 (N_7636,N_6942,N_6528);
nor U7637 (N_7637,N_6441,N_6816);
and U7638 (N_7638,N_6838,N_6150);
and U7639 (N_7639,N_7098,N_6310);
nand U7640 (N_7640,N_7112,N_6795);
nand U7641 (N_7641,N_7448,N_5052);
or U7642 (N_7642,N_6229,N_5179);
xor U7643 (N_7643,N_6345,N_6812);
xnor U7644 (N_7644,N_5599,N_5768);
nand U7645 (N_7645,N_6655,N_6151);
nor U7646 (N_7646,N_6298,N_5011);
or U7647 (N_7647,N_5791,N_6139);
or U7648 (N_7648,N_6214,N_5608);
nor U7649 (N_7649,N_5921,N_6438);
or U7650 (N_7650,N_6790,N_7154);
nor U7651 (N_7651,N_5659,N_6081);
nor U7652 (N_7652,N_5543,N_6955);
and U7653 (N_7653,N_5074,N_7451);
and U7654 (N_7654,N_7086,N_5487);
and U7655 (N_7655,N_7093,N_5104);
and U7656 (N_7656,N_6134,N_5197);
nand U7657 (N_7657,N_5459,N_6217);
and U7658 (N_7658,N_5167,N_5883);
nand U7659 (N_7659,N_7028,N_5072);
or U7660 (N_7660,N_5376,N_7264);
nand U7661 (N_7661,N_6130,N_5700);
nand U7662 (N_7662,N_5704,N_5773);
nor U7663 (N_7663,N_5689,N_6083);
or U7664 (N_7664,N_6270,N_5686);
nor U7665 (N_7665,N_5878,N_6916);
nor U7666 (N_7666,N_5635,N_5742);
and U7667 (N_7667,N_5493,N_5547);
nand U7668 (N_7668,N_6917,N_6657);
xnor U7669 (N_7669,N_7014,N_5673);
nor U7670 (N_7670,N_6936,N_6226);
nand U7671 (N_7671,N_6377,N_6572);
nand U7672 (N_7672,N_5067,N_6359);
or U7673 (N_7673,N_5785,N_5189);
or U7674 (N_7674,N_6695,N_6782);
and U7675 (N_7675,N_5216,N_6734);
and U7676 (N_7676,N_5819,N_6797);
or U7677 (N_7677,N_6541,N_5574);
nor U7678 (N_7678,N_6351,N_5447);
or U7679 (N_7679,N_5606,N_6028);
xnor U7680 (N_7680,N_7110,N_6380);
xnor U7681 (N_7681,N_5220,N_7386);
or U7682 (N_7682,N_5389,N_5807);
xnor U7683 (N_7683,N_5491,N_6978);
nand U7684 (N_7684,N_7171,N_7411);
and U7685 (N_7685,N_6315,N_5965);
nand U7686 (N_7686,N_6843,N_7041);
or U7687 (N_7687,N_7209,N_5232);
or U7688 (N_7688,N_6532,N_5101);
xnor U7689 (N_7689,N_6900,N_6907);
nand U7690 (N_7690,N_5676,N_5118);
and U7691 (N_7691,N_7390,N_6014);
and U7692 (N_7692,N_7427,N_7224);
xnor U7693 (N_7693,N_7275,N_5887);
and U7694 (N_7694,N_7450,N_6465);
or U7695 (N_7695,N_6393,N_7274);
or U7696 (N_7696,N_6905,N_7457);
or U7697 (N_7697,N_5899,N_7117);
and U7698 (N_7698,N_5174,N_5417);
nand U7699 (N_7699,N_6066,N_6160);
xor U7700 (N_7700,N_7477,N_5165);
nor U7701 (N_7701,N_5669,N_5200);
and U7702 (N_7702,N_5088,N_7067);
or U7703 (N_7703,N_6112,N_6503);
nand U7704 (N_7704,N_6461,N_5158);
nand U7705 (N_7705,N_7290,N_6914);
or U7706 (N_7706,N_6183,N_7184);
and U7707 (N_7707,N_7406,N_5569);
nor U7708 (N_7708,N_5971,N_6957);
nand U7709 (N_7709,N_7367,N_5029);
xnor U7710 (N_7710,N_5126,N_6479);
and U7711 (N_7711,N_6920,N_5912);
xor U7712 (N_7712,N_6374,N_7047);
or U7713 (N_7713,N_5308,N_5218);
nor U7714 (N_7714,N_5868,N_6124);
and U7715 (N_7715,N_5637,N_5470);
nand U7716 (N_7716,N_6677,N_5619);
nand U7717 (N_7717,N_6911,N_5277);
and U7718 (N_7718,N_6201,N_6637);
nor U7719 (N_7719,N_5759,N_6448);
xnor U7720 (N_7720,N_5296,N_6709);
and U7721 (N_7721,N_5648,N_5601);
nand U7722 (N_7722,N_5754,N_5488);
and U7723 (N_7723,N_5527,N_5505);
nor U7724 (N_7724,N_5661,N_6883);
nand U7725 (N_7725,N_5806,N_6042);
or U7726 (N_7726,N_7140,N_5658);
nand U7727 (N_7727,N_5646,N_7421);
xnor U7728 (N_7728,N_6371,N_5894);
nand U7729 (N_7729,N_6335,N_5398);
nand U7730 (N_7730,N_5645,N_5872);
or U7731 (N_7731,N_7095,N_5852);
and U7732 (N_7732,N_7350,N_7304);
or U7733 (N_7733,N_5098,N_5610);
nor U7734 (N_7734,N_5050,N_6778);
nor U7735 (N_7735,N_6069,N_7205);
nand U7736 (N_7736,N_6404,N_6624);
xnor U7737 (N_7737,N_7079,N_6779);
and U7738 (N_7738,N_5611,N_6488);
and U7739 (N_7739,N_7283,N_6231);
nor U7740 (N_7740,N_6759,N_7252);
nor U7741 (N_7741,N_5430,N_6946);
or U7742 (N_7742,N_6326,N_7393);
and U7743 (N_7743,N_6508,N_5018);
nor U7744 (N_7744,N_7378,N_5795);
or U7745 (N_7745,N_6728,N_7100);
nor U7746 (N_7746,N_5042,N_5647);
or U7747 (N_7747,N_7156,N_6399);
nor U7748 (N_7748,N_5782,N_5203);
nor U7749 (N_7749,N_5466,N_5958);
nor U7750 (N_7750,N_7097,N_5030);
nor U7751 (N_7751,N_7422,N_6257);
or U7752 (N_7752,N_6125,N_5699);
nand U7753 (N_7753,N_5738,N_5651);
and U7754 (N_7754,N_6539,N_5632);
nand U7755 (N_7755,N_6851,N_6391);
nor U7756 (N_7756,N_6023,N_7414);
or U7757 (N_7757,N_6247,N_6516);
nor U7758 (N_7758,N_6956,N_5805);
and U7759 (N_7759,N_5885,N_5713);
nand U7760 (N_7760,N_5280,N_5078);
nand U7761 (N_7761,N_5953,N_5368);
nor U7762 (N_7762,N_5186,N_5204);
and U7763 (N_7763,N_5335,N_7385);
xor U7764 (N_7764,N_5902,N_5656);
nand U7765 (N_7765,N_5183,N_6645);
or U7766 (N_7766,N_6717,N_6923);
nor U7767 (N_7767,N_6867,N_6100);
and U7768 (N_7768,N_6210,N_6458);
xor U7769 (N_7769,N_6334,N_5784);
nor U7770 (N_7770,N_5037,N_7431);
nand U7771 (N_7771,N_5314,N_6161);
or U7772 (N_7772,N_5624,N_5633);
nand U7773 (N_7773,N_6593,N_5681);
or U7774 (N_7774,N_7308,N_5051);
or U7775 (N_7775,N_6510,N_6573);
or U7776 (N_7776,N_5978,N_5347);
nor U7777 (N_7777,N_5485,N_7134);
nor U7778 (N_7778,N_5435,N_6167);
xor U7779 (N_7779,N_6630,N_7059);
or U7780 (N_7780,N_7094,N_5181);
nor U7781 (N_7781,N_6240,N_5561);
and U7782 (N_7782,N_7286,N_6120);
nor U7783 (N_7783,N_5892,N_6352);
nand U7784 (N_7784,N_7305,N_7215);
nand U7785 (N_7785,N_7163,N_7452);
nand U7786 (N_7786,N_6897,N_6235);
and U7787 (N_7787,N_5917,N_6641);
nand U7788 (N_7788,N_6447,N_7175);
nand U7789 (N_7789,N_7049,N_7297);
or U7790 (N_7790,N_6767,N_5631);
xnor U7791 (N_7791,N_5025,N_5842);
xor U7792 (N_7792,N_7035,N_7314);
or U7793 (N_7793,N_5424,N_5039);
nor U7794 (N_7794,N_6821,N_5140);
and U7795 (N_7795,N_6466,N_5392);
and U7796 (N_7796,N_7392,N_5084);
xnor U7797 (N_7797,N_5458,N_5496);
nor U7798 (N_7798,N_6730,N_6627);
or U7799 (N_7799,N_7063,N_5514);
and U7800 (N_7800,N_6169,N_6250);
nor U7801 (N_7801,N_5915,N_6144);
or U7802 (N_7802,N_5304,N_7238);
or U7803 (N_7803,N_5506,N_7398);
nand U7804 (N_7804,N_6570,N_5589);
and U7805 (N_7805,N_7182,N_7053);
and U7806 (N_7806,N_6686,N_5247);
nor U7807 (N_7807,N_6893,N_7311);
xnor U7808 (N_7808,N_5986,N_6025);
and U7809 (N_7809,N_6171,N_5663);
and U7810 (N_7810,N_6274,N_5567);
or U7811 (N_7811,N_5698,N_6780);
nor U7812 (N_7812,N_6613,N_7167);
or U7813 (N_7813,N_6077,N_6947);
nand U7814 (N_7814,N_5279,N_7396);
nor U7815 (N_7815,N_7129,N_6758);
xnor U7816 (N_7816,N_6678,N_5855);
nor U7817 (N_7817,N_5767,N_5185);
nand U7818 (N_7818,N_5969,N_6245);
xnor U7819 (N_7819,N_7263,N_5278);
xor U7820 (N_7820,N_6755,N_6105);
nand U7821 (N_7821,N_6847,N_5966);
or U7822 (N_7822,N_5393,N_5061);
xnor U7823 (N_7823,N_6592,N_5217);
nor U7824 (N_7824,N_6088,N_5508);
or U7825 (N_7825,N_6002,N_7213);
or U7826 (N_7826,N_6848,N_5929);
or U7827 (N_7827,N_7251,N_6775);
nor U7828 (N_7828,N_5225,N_7267);
xor U7829 (N_7829,N_6004,N_5503);
nor U7830 (N_7830,N_7441,N_6789);
and U7831 (N_7831,N_6965,N_6387);
nand U7832 (N_7832,N_6453,N_6255);
and U7833 (N_7833,N_5310,N_5509);
and U7834 (N_7834,N_5985,N_5679);
nand U7835 (N_7835,N_6859,N_6625);
nand U7836 (N_7836,N_5881,N_7257);
nor U7837 (N_7837,N_5636,N_6132);
or U7838 (N_7838,N_7006,N_7228);
nand U7839 (N_7839,N_6571,N_6228);
nand U7840 (N_7840,N_7176,N_5639);
nand U7841 (N_7841,N_6111,N_5056);
nor U7842 (N_7842,N_5467,N_7223);
nand U7843 (N_7843,N_6554,N_7447);
nand U7844 (N_7844,N_6041,N_6826);
xor U7845 (N_7845,N_6884,N_6713);
and U7846 (N_7846,N_6719,N_7091);
or U7847 (N_7847,N_6649,N_5114);
and U7848 (N_7848,N_5886,N_7432);
xor U7849 (N_7849,N_5272,N_6175);
or U7850 (N_7850,N_7058,N_6459);
and U7851 (N_7851,N_6189,N_5453);
and U7852 (N_7852,N_5489,N_6499);
or U7853 (N_7853,N_5951,N_6328);
nand U7854 (N_7854,N_6485,N_7070);
xnor U7855 (N_7855,N_5823,N_6044);
or U7856 (N_7856,N_6259,N_7072);
and U7857 (N_7857,N_5261,N_6267);
and U7858 (N_7858,N_6746,N_5613);
or U7859 (N_7859,N_5143,N_7199);
nand U7860 (N_7860,N_5627,N_6675);
and U7861 (N_7861,N_5097,N_5519);
nor U7862 (N_7862,N_6230,N_5949);
nand U7863 (N_7863,N_7075,N_5022);
nand U7864 (N_7864,N_6862,N_6358);
and U7865 (N_7865,N_6211,N_5919);
or U7866 (N_7866,N_5816,N_7342);
nor U7867 (N_7867,N_5145,N_5290);
and U7868 (N_7868,N_5734,N_7181);
or U7869 (N_7869,N_7031,N_5122);
nand U7870 (N_7870,N_6047,N_5446);
xor U7871 (N_7871,N_5450,N_5021);
xor U7872 (N_7872,N_6684,N_6639);
nor U7873 (N_7873,N_7124,N_5857);
and U7874 (N_7874,N_5346,N_5706);
and U7875 (N_7875,N_5826,N_5370);
or U7876 (N_7876,N_6136,N_6238);
xor U7877 (N_7877,N_6716,N_5115);
xor U7878 (N_7878,N_6057,N_7408);
or U7879 (N_7879,N_7418,N_5432);
and U7880 (N_7880,N_6423,N_5012);
or U7881 (N_7881,N_6060,N_7484);
and U7882 (N_7882,N_7320,N_7381);
and U7883 (N_7883,N_7210,N_6852);
xor U7884 (N_7884,N_5156,N_7004);
and U7885 (N_7885,N_5191,N_7021);
nand U7886 (N_7886,N_6578,N_7255);
nand U7887 (N_7887,N_5128,N_7227);
and U7888 (N_7888,N_5884,N_7177);
and U7889 (N_7889,N_5457,N_5546);
or U7890 (N_7890,N_7201,N_5438);
and U7891 (N_7891,N_6579,N_5764);
and U7892 (N_7892,N_6086,N_6308);
xor U7893 (N_7893,N_6054,N_7464);
and U7894 (N_7894,N_6379,N_5770);
and U7895 (N_7895,N_7225,N_5644);
and U7896 (N_7896,N_6019,N_5210);
or U7897 (N_7897,N_5132,N_7138);
xnor U7898 (N_7898,N_6765,N_7476);
and U7899 (N_7899,N_7145,N_6314);
nand U7900 (N_7900,N_6791,N_6414);
nand U7901 (N_7901,N_5922,N_6918);
nor U7902 (N_7902,N_6087,N_7336);
and U7903 (N_7903,N_6034,N_5517);
or U7904 (N_7904,N_5668,N_5494);
or U7905 (N_7905,N_5250,N_5413);
nor U7906 (N_7906,N_6986,N_6291);
or U7907 (N_7907,N_6582,N_7382);
or U7908 (N_7908,N_5572,N_7278);
nor U7909 (N_7909,N_6013,N_7380);
or U7910 (N_7910,N_6405,N_6706);
or U7911 (N_7911,N_5177,N_7168);
nand U7912 (N_7912,N_7276,N_6262);
or U7913 (N_7913,N_7042,N_6137);
xor U7914 (N_7914,N_5797,N_5623);
xnor U7915 (N_7915,N_6622,N_7366);
and U7916 (N_7916,N_5521,N_6673);
nand U7917 (N_7917,N_6584,N_5542);
nand U7918 (N_7918,N_5192,N_5827);
nor U7919 (N_7919,N_6783,N_6756);
nor U7920 (N_7920,N_6559,N_7349);
and U7921 (N_7921,N_6729,N_6036);
or U7922 (N_7922,N_5461,N_6055);
and U7923 (N_7923,N_7153,N_6770);
and U7924 (N_7924,N_6222,N_5076);
nor U7925 (N_7925,N_6564,N_6339);
nand U7926 (N_7926,N_7268,N_6953);
nand U7927 (N_7927,N_6850,N_6832);
or U7928 (N_7928,N_7245,N_6792);
xnor U7929 (N_7929,N_7008,N_5263);
nor U7930 (N_7930,N_5238,N_7434);
nor U7931 (N_7931,N_5495,N_5110);
xnor U7932 (N_7932,N_5545,N_5977);
nand U7933 (N_7933,N_7022,N_5600);
nand U7934 (N_7934,N_6306,N_6062);
nor U7935 (N_7935,N_7229,N_7056);
nand U7936 (N_7936,N_6431,N_5345);
nor U7937 (N_7937,N_5988,N_6493);
and U7938 (N_7938,N_7020,N_5405);
xnor U7939 (N_7939,N_6708,N_5719);
xor U7940 (N_7940,N_5146,N_5800);
xor U7941 (N_7941,N_5909,N_6654);
and U7942 (N_7942,N_6609,N_6170);
nor U7943 (N_7943,N_7218,N_7188);
or U7944 (N_7944,N_6147,N_6881);
xnor U7945 (N_7945,N_6075,N_5214);
or U7946 (N_7946,N_6445,N_5242);
and U7947 (N_7947,N_6670,N_5295);
nand U7948 (N_7948,N_5880,N_6619);
and U7949 (N_7949,N_6661,N_6133);
or U7950 (N_7950,N_7488,N_5316);
and U7951 (N_7951,N_7437,N_6991);
nor U7952 (N_7952,N_6094,N_6952);
or U7953 (N_7953,N_6735,N_5979);
or U7954 (N_7954,N_6800,N_6737);
and U7955 (N_7955,N_6363,N_6254);
nor U7956 (N_7956,N_5381,N_5160);
nand U7957 (N_7957,N_6383,N_7438);
and U7958 (N_7958,N_5580,N_6084);
nor U7959 (N_7959,N_5923,N_5950);
or U7960 (N_7960,N_6754,N_6092);
and U7961 (N_7961,N_5241,N_5409);
nand U7962 (N_7962,N_6527,N_6015);
and U7963 (N_7963,N_7473,N_5483);
or U7964 (N_7964,N_6356,N_5386);
or U7965 (N_7965,N_7127,N_5326);
nand U7966 (N_7966,N_7160,N_6669);
or U7967 (N_7967,N_6753,N_6148);
nand U7968 (N_7968,N_6409,N_6174);
and U7969 (N_7969,N_5691,N_6557);
nand U7970 (N_7970,N_7497,N_7064);
nor U7971 (N_7971,N_7352,N_7496);
and U7972 (N_7972,N_7016,N_5869);
and U7973 (N_7973,N_6195,N_6104);
or U7974 (N_7974,N_7123,N_7403);
nor U7975 (N_7975,N_5720,N_5402);
or U7976 (N_7976,N_6003,N_6586);
nor U7977 (N_7977,N_6194,N_6598);
and U7978 (N_7978,N_6472,N_5803);
or U7979 (N_7979,N_5371,N_5288);
nand U7980 (N_7980,N_5998,N_6497);
and U7981 (N_7981,N_5257,N_6841);
nand U7982 (N_7982,N_5340,N_7165);
xnor U7983 (N_7983,N_5105,N_6569);
and U7984 (N_7984,N_7121,N_7354);
and U7985 (N_7985,N_6412,N_6456);
nor U7986 (N_7986,N_6938,N_6185);
xnor U7987 (N_7987,N_5850,N_5712);
nor U7988 (N_7988,N_7061,N_6626);
or U7989 (N_7989,N_7480,N_6408);
and U7990 (N_7990,N_5865,N_6033);
nand U7991 (N_7991,N_6517,N_5879);
nand U7992 (N_7992,N_6869,N_5390);
nor U7993 (N_7993,N_7458,N_5594);
and U7994 (N_7994,N_5337,N_6926);
nand U7995 (N_7995,N_6806,N_7080);
nand U7996 (N_7996,N_5871,N_7193);
nor U7997 (N_7997,N_5338,N_5016);
nand U7998 (N_7998,N_5541,N_6933);
and U7999 (N_7999,N_6357,N_6511);
or U8000 (N_8000,N_5587,N_6417);
nand U8001 (N_8001,N_5728,N_5297);
nand U8002 (N_8002,N_6266,N_6879);
xnor U8003 (N_8003,N_5617,N_5400);
nor U8004 (N_8004,N_6436,N_5520);
nand U8005 (N_8005,N_5783,N_6894);
xnor U8006 (N_8006,N_6864,N_5766);
xnor U8007 (N_8007,N_5421,N_5838);
xnor U8008 (N_8008,N_7142,N_5149);
or U8009 (N_8009,N_6721,N_6396);
xor U8010 (N_8010,N_6482,N_6958);
and U8011 (N_8011,N_5976,N_6921);
and U8012 (N_8012,N_5813,N_6204);
nand U8013 (N_8013,N_5073,N_5092);
nor U8014 (N_8014,N_6704,N_6590);
nand U8015 (N_8015,N_6674,N_6154);
or U8016 (N_8016,N_5804,N_7253);
nand U8017 (N_8017,N_7365,N_6809);
and U8018 (N_8018,N_7298,N_5725);
and U8019 (N_8019,N_5476,N_7471);
nand U8020 (N_8020,N_5705,N_6886);
or U8021 (N_8021,N_5188,N_5660);
nand U8022 (N_8022,N_5693,N_6644);
nand U8023 (N_8023,N_5695,N_7334);
xnor U8024 (N_8024,N_7226,N_6574);
or U8025 (N_8025,N_6442,N_6543);
and U8026 (N_8026,N_5536,N_7377);
nor U8027 (N_8027,N_5955,N_6220);
or U8028 (N_8028,N_6143,N_6067);
nor U8029 (N_8029,N_6562,N_6703);
nor U8030 (N_8030,N_6449,N_5544);
nand U8031 (N_8031,N_6389,N_5331);
nand U8032 (N_8032,N_5367,N_6727);
or U8033 (N_8033,N_7001,N_5168);
or U8034 (N_8034,N_5987,N_6763);
or U8035 (N_8035,N_6248,N_5935);
nor U8036 (N_8036,N_6974,N_6258);
nor U8037 (N_8037,N_6801,N_5618);
nor U8038 (N_8038,N_7328,N_6361);
nand U8039 (N_8039,N_7324,N_5463);
and U8040 (N_8040,N_5891,N_7137);
nor U8041 (N_8041,N_6983,N_5983);
xnor U8042 (N_8042,N_5283,N_5436);
nand U8043 (N_8043,N_5219,N_6477);
nor U8044 (N_8044,N_7077,N_5412);
or U8045 (N_8045,N_6576,N_5206);
nor U8046 (N_8046,N_5380,N_6464);
or U8047 (N_8047,N_5269,N_7400);
nand U8048 (N_8048,N_6691,N_6992);
nand U8049 (N_8049,N_5584,N_6536);
nor U8050 (N_8050,N_5213,N_7107);
nand U8051 (N_8051,N_5847,N_7482);
or U8052 (N_8052,N_6317,N_6416);
nor U8053 (N_8053,N_5017,N_6949);
and U8054 (N_8054,N_5187,N_5448);
or U8055 (N_8055,N_6922,N_7212);
and U8056 (N_8056,N_6440,N_6944);
nand U8057 (N_8057,N_5339,N_7287);
or U8058 (N_8058,N_7492,N_5993);
or U8059 (N_8059,N_6007,N_7085);
and U8060 (N_8060,N_6048,N_6040);
nand U8061 (N_8061,N_6773,N_7048);
or U8062 (N_8062,N_7424,N_7037);
nand U8063 (N_8063,N_6252,N_6056);
nand U8064 (N_8064,N_5026,N_7189);
or U8065 (N_8065,N_5615,N_6418);
or U8066 (N_8066,N_5369,N_5091);
or U8067 (N_8067,N_5103,N_6312);
nor U8068 (N_8068,N_5596,N_5311);
or U8069 (N_8069,N_5948,N_6263);
or U8070 (N_8070,N_5938,N_7420);
or U8071 (N_8071,N_5325,N_6652);
xor U8072 (N_8072,N_7289,N_5654);
xor U8073 (N_8073,N_5102,N_5240);
and U8074 (N_8074,N_5642,N_6998);
and U8075 (N_8075,N_7198,N_7306);
or U8076 (N_8076,N_5535,N_5426);
or U8077 (N_8077,N_5129,N_5787);
and U8078 (N_8078,N_5864,N_5260);
and U8079 (N_8079,N_6787,N_6366);
and U8080 (N_8080,N_6268,N_6446);
or U8081 (N_8081,N_5529,N_7487);
nand U8082 (N_8082,N_7146,N_5538);
or U8083 (N_8083,N_7194,N_5150);
and U8084 (N_8084,N_6606,N_5138);
and U8085 (N_8085,N_5931,N_6321);
nand U8086 (N_8086,N_7109,N_6052);
and U8087 (N_8087,N_5049,N_6665);
and U8088 (N_8088,N_6885,N_6241);
or U8089 (N_8089,N_5256,N_5717);
nand U8090 (N_8090,N_6193,N_5507);
nand U8091 (N_8091,N_5275,N_7440);
nor U8092 (N_8092,N_5205,N_5528);
xnor U8093 (N_8093,N_6187,N_5863);
or U8094 (N_8094,N_6401,N_6732);
nor U8095 (N_8095,N_5043,N_7060);
and U8096 (N_8096,N_6750,N_6355);
nor U8097 (N_8097,N_6474,N_7013);
nor U8098 (N_8098,N_5397,N_5472);
or U8099 (N_8099,N_6629,N_6537);
or U8100 (N_8100,N_5484,N_6785);
nand U8101 (N_8101,N_7346,N_5385);
nand U8102 (N_8102,N_5997,N_5531);
or U8103 (N_8103,N_7187,N_5708);
nor U8104 (N_8104,N_5482,N_6823);
and U8105 (N_8105,N_5775,N_6017);
nand U8106 (N_8106,N_7362,N_6696);
nor U8107 (N_8107,N_6932,N_6299);
or U8108 (N_8108,N_5779,N_7051);
or U8109 (N_8109,N_5771,N_6289);
nand U8110 (N_8110,N_6179,N_7130);
and U8111 (N_8111,N_7409,N_5180);
nand U8112 (N_8112,N_6877,N_5559);
xor U8113 (N_8113,N_5023,N_5774);
nor U8114 (N_8114,N_5422,N_7033);
nor U8115 (N_8115,N_5077,N_5287);
nand U8116 (N_8116,N_6191,N_6032);
nor U8117 (N_8117,N_5107,N_6710);
nor U8118 (N_8118,N_6181,N_7151);
and U8119 (N_8119,N_5047,N_7183);
nor U8120 (N_8120,N_6365,N_6831);
or U8121 (N_8121,N_6460,N_7159);
and U8122 (N_8122,N_7347,N_6138);
and U8123 (N_8123,N_7169,N_5100);
nor U8124 (N_8124,N_5682,N_5239);
nor U8125 (N_8125,N_6788,N_7485);
nor U8126 (N_8126,N_7490,N_6123);
or U8127 (N_8127,N_7486,N_6692);
and U8128 (N_8128,N_5913,N_6846);
nor U8129 (N_8129,N_6607,N_6116);
and U8130 (N_8130,N_6061,N_5723);
or U8131 (N_8131,N_5497,N_5961);
nand U8132 (N_8132,N_5745,N_6835);
nor U8133 (N_8133,N_6469,N_6106);
nand U8134 (N_8134,N_5141,N_6659);
or U8135 (N_8135,N_7003,N_6997);
or U8136 (N_8136,N_5898,N_6839);
and U8137 (N_8137,N_6514,N_5411);
nor U8138 (N_8138,N_6275,N_6875);
and U8139 (N_8139,N_6109,N_7397);
and U8140 (N_8140,N_7233,N_6899);
nand U8141 (N_8141,N_6707,N_5079);
nand U8142 (N_8142,N_5622,N_6739);
and U8143 (N_8143,N_6122,N_5106);
and U8144 (N_8144,N_5044,N_5652);
nor U8145 (N_8145,N_7295,N_6725);
nor U8146 (N_8146,N_5013,N_6827);
or U8147 (N_8147,N_6994,N_6117);
nand U8148 (N_8148,N_6454,N_5841);
nand U8149 (N_8149,N_7073,N_5360);
nor U8150 (N_8150,N_6102,N_6908);
nor U8151 (N_8151,N_6237,N_7236);
nand U8152 (N_8152,N_7491,N_5970);
nor U8153 (N_8153,N_5640,N_5836);
or U8154 (N_8154,N_7472,N_5996);
nor U8155 (N_8155,N_6080,N_7413);
and U8156 (N_8156,N_6747,N_5322);
nand U8157 (N_8157,N_5946,N_5905);
xnor U8158 (N_8158,N_5199,N_5566);
or U8159 (N_8159,N_5741,N_6546);
and U8160 (N_8160,N_5477,N_5634);
nand U8161 (N_8161,N_5066,N_6985);
nor U8162 (N_8162,N_6752,N_5224);
xnor U8163 (N_8163,N_7344,N_6279);
nand U8164 (N_8164,N_6825,N_6020);
and U8165 (N_8165,N_6993,N_5750);
nor U8166 (N_8166,N_7232,N_6731);
nand U8167 (N_8167,N_5408,N_5373);
nand U8168 (N_8168,N_5271,N_6483);
nand U8169 (N_8169,N_5897,N_5416);
xor U8170 (N_8170,N_5010,N_6188);
and U8171 (N_8171,N_5914,N_7241);
xnor U8172 (N_8172,N_6615,N_5048);
or U8173 (N_8173,N_6542,N_7239);
xor U8174 (N_8174,N_7384,N_5267);
and U8175 (N_8175,N_6395,N_6585);
or U8176 (N_8176,N_6037,N_5124);
nor U8177 (N_8177,N_7402,N_5604);
or U8178 (N_8178,N_7074,N_5270);
or U8179 (N_8179,N_5231,N_5515);
nand U8180 (N_8180,N_5840,N_5918);
or U8181 (N_8181,N_5343,N_5388);
and U8182 (N_8182,N_5502,N_5714);
or U8183 (N_8183,N_6774,N_6979);
nand U8184 (N_8184,N_5968,N_5924);
or U8185 (N_8185,N_7260,N_6385);
and U8186 (N_8186,N_5135,N_5558);
or U8187 (N_8187,N_7459,N_7461);
or U8188 (N_8188,N_6676,N_5954);
or U8189 (N_8189,N_6901,N_5824);
nand U8190 (N_8190,N_5182,N_5866);
or U8191 (N_8191,N_6705,N_6068);
or U8192 (N_8192,N_6534,N_6165);
nor U8193 (N_8193,N_6803,N_7087);
and U8194 (N_8194,N_6273,N_6058);
and U8195 (N_8195,N_5228,N_5329);
nor U8196 (N_8196,N_5638,N_5730);
or U8197 (N_8197,N_6568,N_6182);
or U8198 (N_8198,N_6163,N_5382);
nand U8199 (N_8199,N_5258,N_7259);
and U8200 (N_8200,N_7416,N_6545);
nand U8201 (N_8201,N_6384,N_6558);
nor U8202 (N_8202,N_5972,N_6085);
or U8203 (N_8203,N_6323,N_6762);
nor U8204 (N_8204,N_6295,N_7284);
and U8205 (N_8205,N_5490,N_6035);
xor U8206 (N_8206,N_6221,N_6413);
nand U8207 (N_8207,N_7162,N_6244);
nand U8208 (N_8208,N_7371,N_6309);
nand U8209 (N_8209,N_6145,N_5831);
or U8210 (N_8210,N_7065,N_5032);
or U8211 (N_8211,N_6663,N_5697);
and U8212 (N_8212,N_5653,N_6012);
nand U8213 (N_8213,N_7321,N_7428);
or U8214 (N_8214,N_7222,N_6642);
nand U8215 (N_8215,N_5620,N_6439);
nand U8216 (N_8216,N_6243,N_5628);
xnor U8217 (N_8217,N_5294,N_7454);
xnor U8218 (N_8218,N_5579,N_5212);
xor U8219 (N_8219,N_7133,N_7192);
and U8220 (N_8220,N_5330,N_7407);
nor U8221 (N_8221,N_6761,N_6451);
or U8222 (N_8222,N_7415,N_7313);
or U8223 (N_8223,N_6989,N_7135);
and U8224 (N_8224,N_5510,N_6475);
nor U8225 (N_8225,N_7330,N_6502);
or U8226 (N_8226,N_5609,N_6804);
nor U8227 (N_8227,N_6239,N_5229);
or U8228 (N_8228,N_7068,N_5117);
or U8229 (N_8229,N_6271,N_5406);
nor U8230 (N_8230,N_5276,N_6362);
and U8231 (N_8231,N_5670,N_7310);
xnor U8232 (N_8232,N_5328,N_5756);
nor U8233 (N_8233,N_6648,N_5299);
and U8234 (N_8234,N_6063,N_5778);
nand U8235 (N_8235,N_6525,N_5082);
nor U8236 (N_8236,N_6098,N_5383);
nand U8237 (N_8237,N_5737,N_7489);
nor U8238 (N_8238,N_5678,N_5761);
and U8239 (N_8239,N_6980,N_6207);
and U8240 (N_8240,N_5870,N_5058);
nor U8241 (N_8241,N_6010,N_5081);
or U8242 (N_8242,N_6567,N_5744);
nand U8243 (N_8243,N_7118,N_7339);
and U8244 (N_8244,N_6810,N_6205);
nand U8245 (N_8245,N_5208,N_6972);
and U8246 (N_8246,N_7469,N_7089);
nand U8247 (N_8247,N_7271,N_7139);
or U8248 (N_8248,N_7190,N_7150);
nand U8249 (N_8249,N_5882,N_5995);
nand U8250 (N_8250,N_5825,N_6101);
and U8251 (N_8251,N_6382,N_6861);
nand U8252 (N_8252,N_5378,N_5274);
nand U8253 (N_8253,N_5355,N_5602);
and U8254 (N_8254,N_5469,N_5975);
nand U8255 (N_8255,N_6364,N_5662);
nand U8256 (N_8256,N_5262,N_6341);
nand U8257 (N_8257,N_5711,N_5575);
nor U8258 (N_8258,N_5875,N_6072);
or U8259 (N_8259,N_6354,N_7301);
nand U8260 (N_8260,N_6196,N_5480);
nor U8261 (N_8261,N_5099,N_6001);
nand U8262 (N_8262,N_6906,N_7360);
or U8263 (N_8263,N_5874,N_5598);
nand U8264 (N_8264,N_5675,N_5989);
and U8265 (N_8265,N_6486,N_6689);
xor U8266 (N_8266,N_7364,N_6680);
or U8267 (N_8267,N_5928,N_6197);
and U8268 (N_8268,N_5829,N_6327);
xor U8269 (N_8269,N_5616,N_6856);
and U8270 (N_8270,N_6961,N_5147);
nand U8271 (N_8271,N_6376,N_7466);
or U8272 (N_8272,N_5006,N_6303);
nor U8273 (N_8273,N_5222,N_5570);
and U8274 (N_8274,N_6599,N_6507);
and U8275 (N_8275,N_6693,N_5940);
and U8276 (N_8276,N_5336,N_6966);
or U8277 (N_8277,N_5152,N_6030);
nor U8278 (N_8278,N_6024,N_6011);
nand U8279 (N_8279,N_5504,N_5253);
nor U8280 (N_8280,N_6264,N_7391);
nand U8281 (N_8281,N_5843,N_6814);
nand U8282 (N_8282,N_6282,N_5614);
nor U8283 (N_8283,N_5501,N_7164);
or U8284 (N_8284,N_6533,N_7481);
xnor U8285 (N_8285,N_5148,N_5649);
and U8286 (N_8286,N_7005,N_5724);
and U8287 (N_8287,N_6555,N_5157);
nand U8288 (N_8288,N_6928,N_7078);
nor U8289 (N_8289,N_5817,N_5418);
or U8290 (N_8290,N_6688,N_5350);
and U8291 (N_8291,N_7149,N_6079);
nand U8292 (N_8292,N_5499,N_7174);
nand U8293 (N_8293,N_7052,N_6764);
nand U8294 (N_8294,N_6601,N_6715);
xor U8295 (N_8295,N_6343,N_5000);
xor U8296 (N_8296,N_5981,N_6740);
or U8297 (N_8297,N_5071,N_6611);
nand U8298 (N_8298,N_5757,N_6866);
or U8299 (N_8299,N_6471,N_7106);
and U8300 (N_8300,N_5665,N_6350);
nor U8301 (N_8301,N_6813,N_6494);
and U8302 (N_8302,N_5342,N_6272);
or U8303 (N_8303,N_6348,N_6406);
nand U8304 (N_8304,N_6070,N_7309);
nor U8305 (N_8305,N_6519,N_6180);
xor U8306 (N_8306,N_6522,N_7030);
xor U8307 (N_8307,N_7143,N_7318);
and U8308 (N_8308,N_5273,N_6219);
or U8309 (N_8309,N_7088,N_5359);
or U8310 (N_8310,N_6913,N_6614);
xor U8311 (N_8311,N_6121,N_5733);
and U8312 (N_8312,N_6833,N_6807);
and U8313 (N_8313,N_5927,N_7114);
and U8314 (N_8314,N_6234,N_6489);
and U8315 (N_8315,N_5019,N_5171);
and U8316 (N_8316,N_6006,N_7206);
nand U8317 (N_8317,N_5629,N_5356);
xnor U8318 (N_8318,N_5313,N_5123);
or U8319 (N_8319,N_6547,N_6506);
and U8320 (N_8320,N_5366,N_7027);
nand U8321 (N_8321,N_7026,N_6679);
and U8322 (N_8322,N_6766,N_7355);
nor U8323 (N_8323,N_5244,N_6701);
nor U8324 (N_8324,N_6420,N_6162);
nand U8325 (N_8325,N_5353,N_6256);
nor U8326 (N_8326,N_5038,N_6108);
xor U8327 (N_8327,N_5420,N_5552);
or U8328 (N_8328,N_5687,N_6837);
or U8329 (N_8329,N_5731,N_6811);
xor U8330 (N_8330,N_7279,N_5903);
nand U8331 (N_8331,N_5321,N_7273);
nor U8332 (N_8332,N_6929,N_5952);
xnor U8333 (N_8333,N_6260,N_6538);
nor U8334 (N_8334,N_5065,N_6518);
nor U8335 (N_8335,N_7307,N_6353);
nor U8336 (N_8336,N_5301,N_5282);
xor U8337 (N_8337,N_6940,N_5755);
nor U8338 (N_8338,N_6840,N_7249);
and U8339 (N_8339,N_5943,N_6656);
or U8340 (N_8340,N_6203,N_7478);
and U8341 (N_8341,N_7128,N_7101);
nor U8342 (N_8342,N_6898,N_6039);
and U8343 (N_8343,N_6690,N_5184);
and U8344 (N_8344,N_6501,N_5677);
nand U8345 (N_8345,N_5377,N_7057);
and U8346 (N_8346,N_5583,N_5352);
or U8347 (N_8347,N_5410,N_7272);
and U8348 (N_8348,N_6022,N_5384);
nand U8349 (N_8349,N_6126,N_5581);
and U8350 (N_8350,N_6421,N_5592);
nand U8351 (N_8351,N_5401,N_6369);
xor U8352 (N_8352,N_6184,N_5320);
or U8353 (N_8353,N_7062,N_7433);
or U8354 (N_8354,N_7388,N_6470);
nand U8355 (N_8355,N_7015,N_5358);
nor U8356 (N_8356,N_7296,N_5121);
nor U8357 (N_8357,N_5034,N_5585);
or U8358 (N_8358,N_7261,N_6156);
nor U8359 (N_8359,N_7322,N_6186);
nand U8360 (N_8360,N_7265,N_6430);
nand U8361 (N_8361,N_5014,N_5999);
nand U8362 (N_8362,N_5630,N_7280);
and U8363 (N_8363,N_6253,N_5334);
nor U8364 (N_8364,N_5808,N_5234);
nand U8365 (N_8365,N_5593,N_5454);
nand U8366 (N_8366,N_5846,N_7084);
nand U8367 (N_8367,N_7247,N_6090);
or U8368 (N_8368,N_6324,N_7446);
nor U8369 (N_8369,N_7300,N_7375);
nand U8370 (N_8370,N_6021,N_7499);
or U8371 (N_8371,N_7426,N_6375);
nand U8372 (N_8372,N_7425,N_6722);
or U8373 (N_8373,N_5486,N_6664);
nand U8374 (N_8374,N_6505,N_7423);
xor U8375 (N_8375,N_5395,N_6158);
nor U8376 (N_8376,N_5243,N_5130);
nand U8377 (N_8377,N_6995,N_5798);
nor U8378 (N_8378,N_5667,N_5317);
and U8379 (N_8379,N_6437,N_5173);
or U8380 (N_8380,N_6597,N_6799);
nor U8381 (N_8381,N_5994,N_5556);
or U8382 (N_8382,N_7453,N_5562);
nand U8383 (N_8383,N_5315,N_5539);
or U8384 (N_8384,N_6168,N_5571);
and U8385 (N_8385,N_5028,N_5582);
or U8386 (N_8386,N_6954,N_5252);
or U8387 (N_8387,N_5434,N_5672);
xnor U8388 (N_8388,N_5643,N_5080);
nand U8389 (N_8389,N_7288,N_5202);
and U8390 (N_8390,N_5498,N_7081);
and U8391 (N_8391,N_6198,N_5024);
and U8392 (N_8392,N_5303,N_5237);
and U8393 (N_8393,N_6491,N_5657);
or U8394 (N_8394,N_6860,N_7449);
and U8395 (N_8395,N_5777,N_6738);
nor U8396 (N_8396,N_7019,N_6373);
and U8397 (N_8397,N_7011,N_5834);
nor U8398 (N_8398,N_5605,N_6930);
nor U8399 (N_8399,N_6526,N_6400);
nor U8400 (N_8400,N_6492,N_7207);
or U8401 (N_8401,N_6450,N_5045);
or U8402 (N_8402,N_7002,N_6699);
and U8403 (N_8403,N_6051,N_7460);
and U8404 (N_8404,N_5573,N_5007);
or U8405 (N_8405,N_6820,N_6155);
nor U8406 (N_8406,N_5591,N_6937);
and U8407 (N_8407,N_7341,N_6236);
nand U8408 (N_8408,N_7348,N_5934);
or U8409 (N_8409,N_7358,N_7498);
and U8410 (N_8410,N_5151,N_5462);
nor U8411 (N_8411,N_6512,N_5512);
nand U8412 (N_8412,N_6857,N_5780);
nor U8413 (N_8413,N_6934,N_5086);
and U8414 (N_8414,N_5440,N_5890);
or U8415 (N_8415,N_5003,N_5944);
nand U8416 (N_8416,N_6834,N_5054);
nand U8417 (N_8417,N_7410,N_7326);
xnor U8418 (N_8418,N_6815,N_7363);
or U8419 (N_8419,N_5319,N_5087);
or U8420 (N_8420,N_5333,N_6605);
or U8421 (N_8421,N_5859,N_7111);
and U8422 (N_8422,N_6902,N_6026);
nor U8423 (N_8423,N_5113,N_6698);
or U8424 (N_8424,N_5534,N_5739);
nand U8425 (N_8425,N_7120,N_6390);
or U8426 (N_8426,N_5468,N_7122);
nand U8427 (N_8427,N_7369,N_6604);
nor U8428 (N_8428,N_6065,N_5790);
nor U8429 (N_8429,N_6038,N_5942);
or U8430 (N_8430,N_5576,N_6113);
nand U8431 (N_8431,N_6192,N_7191);
and U8432 (N_8432,N_5404,N_5941);
or U8433 (N_8433,N_5020,N_6781);
or U8434 (N_8434,N_6473,N_5763);
xor U8435 (N_8435,N_5726,N_7430);
nor U8436 (N_8436,N_5577,N_6772);
or U8437 (N_8437,N_5732,N_7069);
nor U8438 (N_8438,N_7220,N_5127);
nor U8439 (N_8439,N_6029,N_7195);
or U8440 (N_8440,N_5230,N_5895);
xor U8441 (N_8441,N_6342,N_5947);
or U8442 (N_8442,N_6463,N_5901);
or U8443 (N_8443,N_6633,N_5284);
and U8444 (N_8444,N_6128,N_5548);
or U8445 (N_8445,N_6149,N_5255);
nand U8446 (N_8446,N_7071,N_5433);
nor U8447 (N_8447,N_5707,N_5814);
nor U8448 (N_8448,N_5603,N_5062);
and U8449 (N_8449,N_5578,N_5341);
and U8450 (N_8450,N_6304,N_6720);
nand U8451 (N_8451,N_6895,N_6742);
and U8452 (N_8452,N_5083,N_5962);
and U8453 (N_8453,N_5142,N_5002);
nand U8454 (N_8454,N_5060,N_6206);
xnor U8455 (N_8455,N_7282,N_6771);
and U8456 (N_8456,N_5554,N_7479);
or U8457 (N_8457,N_5351,N_6381);
nand U8458 (N_8458,N_6099,N_6662);
nand U8459 (N_8459,N_5664,N_5526);
and U8460 (N_8460,N_6982,N_5264);
or U8461 (N_8461,N_6349,N_5911);
and U8462 (N_8462,N_6005,N_5198);
and U8463 (N_8463,N_5960,N_6318);
or U8464 (N_8464,N_6504,N_7180);
and U8465 (N_8465,N_6457,N_5407);
and U8466 (N_8466,N_5251,N_5560);
nand U8467 (N_8467,N_6963,N_7090);
and U8468 (N_8468,N_5292,N_6636);
nand U8469 (N_8469,N_6509,N_6976);
nand U8470 (N_8470,N_5849,N_5625);
nand U8471 (N_8471,N_6939,N_5005);
or U8472 (N_8472,N_6114,N_7325);
nand U8473 (N_8473,N_6200,N_6016);
or U8474 (N_8474,N_7240,N_6776);
or U8475 (N_8475,N_5815,N_5786);
nor U8476 (N_8476,N_7147,N_5027);
nand U8477 (N_8477,N_5749,N_5694);
or U8478 (N_8478,N_7395,N_7179);
and U8479 (N_8479,N_7405,N_5873);
or U8480 (N_8480,N_5414,N_6110);
nor U8481 (N_8481,N_6091,N_5746);
and U8482 (N_8482,N_6638,N_7126);
nor U8483 (N_8483,N_5565,N_6587);
or U8484 (N_8484,N_5428,N_6031);
nand U8485 (N_8485,N_7131,N_5500);
nand U8486 (N_8486,N_5743,N_5456);
or U8487 (N_8487,N_6876,N_6286);
and U8488 (N_8488,N_6325,N_5403);
nand U8489 (N_8489,N_6798,N_6398);
xor U8490 (N_8490,N_6950,N_5736);
or U8491 (N_8491,N_5041,N_6153);
and U8492 (N_8492,N_7292,N_6411);
nor U8493 (N_8493,N_5365,N_6209);
nand U8494 (N_8494,N_6530,N_7379);
and U8495 (N_8495,N_5851,N_6822);
nand U8496 (N_8496,N_6768,N_5936);
or U8497 (N_8497,N_5479,N_5164);
or U8498 (N_8498,N_5789,N_6277);
nor U8499 (N_8499,N_6863,N_6316);
and U8500 (N_8500,N_7099,N_7303);
nand U8501 (N_8501,N_7455,N_6311);
and U8502 (N_8502,N_5925,N_5166);
or U8503 (N_8503,N_5957,N_6830);
or U8504 (N_8504,N_5445,N_5439);
and U8505 (N_8505,N_6845,N_5449);
and U8506 (N_8506,N_7493,N_6878);
and U8507 (N_8507,N_7412,N_7474);
and U8508 (N_8508,N_6646,N_6658);
nand U8509 (N_8509,N_5641,N_7357);
xor U8510 (N_8510,N_6050,N_7383);
or U8511 (N_8511,N_6059,N_7144);
nand U8512 (N_8512,N_5473,N_6027);
and U8513 (N_8513,N_6910,N_7401);
and U8514 (N_8514,N_7333,N_5035);
and U8515 (N_8515,N_6513,N_5125);
nor U8516 (N_8516,N_6580,N_6634);
and U8517 (N_8517,N_6093,N_5727);
or U8518 (N_8518,N_5155,N_7039);
nand U8519 (N_8519,N_5195,N_6452);
or U8520 (N_8520,N_6429,N_5540);
and U8521 (N_8521,N_5716,N_5959);
xnor U8522 (N_8522,N_5533,N_6337);
and U8523 (N_8523,N_6076,N_7132);
and U8524 (N_8524,N_5932,N_6873);
and U8525 (N_8525,N_7353,N_5134);
or U8526 (N_8526,N_7443,N_6855);
or U8527 (N_8527,N_7319,N_7317);
xor U8528 (N_8528,N_5590,N_7076);
and U8529 (N_8529,N_5788,N_6667);
nor U8530 (N_8530,N_6951,N_5830);
nor U8531 (N_8531,N_5286,N_7141);
nand U8532 (N_8532,N_7243,N_5169);
and U8533 (N_8533,N_6000,N_5362);
or U8534 (N_8534,N_6340,N_5095);
or U8535 (N_8535,N_5524,N_7376);
and U8536 (N_8536,N_6711,N_5984);
nand U8537 (N_8537,N_5227,N_5068);
nor U8538 (N_8538,N_5794,N_6246);
and U8539 (N_8539,N_5111,N_6520);
and U8540 (N_8540,N_5057,N_5607);
nand U8541 (N_8541,N_6285,N_6566);
or U8542 (N_8542,N_6935,N_7161);
nand U8543 (N_8543,N_5557,N_6653);
nand U8544 (N_8544,N_7417,N_6118);
nand U8545 (N_8545,N_6468,N_5481);
nor U8546 (N_8546,N_6212,N_6631);
nand U8547 (N_8547,N_6008,N_5008);
or U8548 (N_8548,N_5215,N_6146);
nor U8549 (N_8549,N_6331,N_6620);
or U8550 (N_8550,N_7158,N_6999);
or U8551 (N_8551,N_6608,N_5004);
nand U8552 (N_8552,N_6141,N_7399);
or U8553 (N_8553,N_6971,N_6199);
nand U8554 (N_8554,N_5452,N_5518);
and U8555 (N_8555,N_7152,N_5289);
nor U8556 (N_8556,N_5937,N_7445);
nor U8557 (N_8557,N_5415,N_6073);
or U8558 (N_8558,N_6415,N_5926);
and U8559 (N_8559,N_5974,N_7208);
nand U8560 (N_8560,N_5809,N_5235);
nand U8561 (N_8561,N_5861,N_5170);
xnor U8562 (N_8562,N_5671,N_6190);
xor U8563 (N_8563,N_7468,N_7018);
xnor U8564 (N_8564,N_6320,N_7172);
or U8565 (N_8565,N_5910,N_7258);
nand U8566 (N_8566,N_7230,N_5372);
or U8567 (N_8567,N_6868,N_6660);
and U8568 (N_8568,N_6346,N_7103);
nor U8569 (N_8569,N_6733,N_7155);
or U8570 (N_8570,N_7329,N_6870);
nand U8571 (N_8571,N_7343,N_7203);
xor U8572 (N_8572,N_5588,N_7293);
nor U8573 (N_8573,N_6551,N_5323);
nor U8574 (N_8574,N_7082,N_6632);
or U8575 (N_8575,N_7115,N_5595);
and U8576 (N_8576,N_6372,N_6096);
and U8577 (N_8577,N_5201,N_5523);
or U8578 (N_8578,N_6964,N_5427);
nand U8579 (N_8579,N_5980,N_7044);
and U8580 (N_8580,N_6332,N_6565);
nor U8581 (N_8581,N_5190,N_6941);
nand U8582 (N_8582,N_6628,N_5302);
nand U8583 (N_8583,N_5621,N_5307);
nor U8584 (N_8584,N_5701,N_5015);
and U8585 (N_8585,N_6945,N_6808);
or U8586 (N_8586,N_5293,N_7248);
nand U8587 (N_8587,N_7096,N_7043);
xnor U8588 (N_8588,N_5796,N_5751);
or U8589 (N_8589,N_6142,N_5419);
nor U8590 (N_8590,N_5858,N_5839);
and U8591 (N_8591,N_5833,N_5956);
or U8592 (N_8592,N_6700,N_7211);
nor U8593 (N_8593,N_6476,N_5236);
xor U8594 (N_8594,N_7202,N_6726);
nor U8595 (N_8595,N_6515,N_7281);
nor U8596 (N_8596,N_6278,N_5802);
nand U8597 (N_8597,N_6386,N_6292);
nor U8598 (N_8598,N_7323,N_6531);
or U8599 (N_8599,N_5904,N_5492);
and U8600 (N_8600,N_7442,N_7302);
nand U8601 (N_8601,N_7196,N_7185);
and U8602 (N_8602,N_5564,N_5854);
nand U8603 (N_8603,N_6276,N_7291);
or U8604 (N_8604,N_6904,N_7029);
or U8605 (N_8605,N_7465,N_6403);
and U8606 (N_8606,N_5046,N_6424);
and U8607 (N_8607,N_6769,N_6948);
or U8608 (N_8608,N_6817,N_6053);
or U8609 (N_8609,N_6924,N_7470);
nand U8610 (N_8610,N_5108,N_5265);
xor U8611 (N_8611,N_6432,N_6635);
or U8612 (N_8612,N_7204,N_5760);
nor U8613 (N_8613,N_6290,N_7254);
and U8614 (N_8614,N_5721,N_6560);
nor U8615 (N_8615,N_6896,N_6434);
or U8616 (N_8616,N_5094,N_7136);
or U8617 (N_8617,N_5832,N_5009);
and U8618 (N_8618,N_6561,N_7219);
nor U8619 (N_8619,N_6836,N_7105);
and U8620 (N_8620,N_7456,N_5441);
nand U8621 (N_8621,N_6751,N_6500);
nand U8622 (N_8622,N_6842,N_6981);
and U8623 (N_8623,N_6577,N_6931);
nor U8624 (N_8624,N_6549,N_6216);
xnor U8625 (N_8625,N_5431,N_5729);
nand U8626 (N_8626,N_7010,N_6736);
nor U8627 (N_8627,N_5674,N_5666);
nor U8628 (N_8628,N_7331,N_6009);
xnor U8629 (N_8629,N_6444,N_7463);
nand U8630 (N_8630,N_5391,N_5444);
and U8631 (N_8631,N_7404,N_6621);
or U8632 (N_8632,N_7312,N_7368);
and U8633 (N_8633,N_5964,N_5475);
xor U8634 (N_8634,N_7009,N_7270);
or U8635 (N_8635,N_5176,N_6888);
or U8636 (N_8636,N_7054,N_7032);
nand U8637 (N_8637,N_6462,N_6467);
or U8638 (N_8638,N_6119,N_6819);
and U8639 (N_8639,N_5828,N_5835);
or U8640 (N_8640,N_6043,N_6595);
xnor U8641 (N_8641,N_5465,N_5139);
or U8642 (N_8642,N_7102,N_5626);
and U8643 (N_8643,N_5811,N_5085);
nor U8644 (N_8644,N_6552,N_5172);
xor U8645 (N_8645,N_5324,N_7025);
and U8646 (N_8646,N_5162,N_6967);
or U8647 (N_8647,N_5550,N_7113);
nand U8648 (N_8648,N_6302,N_5036);
or U8649 (N_8649,N_6602,N_6202);
or U8650 (N_8650,N_5860,N_6589);
and U8651 (N_8651,N_5793,N_6392);
nor U8652 (N_8652,N_5175,N_7361);
nand U8653 (N_8653,N_6164,N_6283);
or U8654 (N_8654,N_5464,N_6422);
and U8655 (N_8655,N_6296,N_5876);
nor U8656 (N_8656,N_6968,N_7351);
or U8657 (N_8657,N_6107,N_6872);
and U8658 (N_8658,N_6487,N_5982);
nand U8659 (N_8659,N_6892,N_5209);
xnor U8660 (N_8660,N_5455,N_6617);
or U8661 (N_8661,N_6074,N_6224);
or U8662 (N_8662,N_5196,N_6651);
or U8663 (N_8663,N_6157,N_5769);
xnor U8664 (N_8664,N_5685,N_6481);
nor U8665 (N_8665,N_5553,N_6397);
nor U8666 (N_8666,N_5696,N_5375);
nor U8667 (N_8667,N_5254,N_5055);
nor U8668 (N_8668,N_7221,N_6367);
or U8669 (N_8669,N_6127,N_7315);
nand U8670 (N_8670,N_5348,N_5268);
and U8671 (N_8671,N_6909,N_6360);
nand U8672 (N_8672,N_6844,N_5967);
or U8673 (N_8673,N_7066,N_6521);
nor U8674 (N_8674,N_6330,N_7277);
nor U8675 (N_8675,N_5963,N_6741);
xnor U8676 (N_8676,N_7475,N_7092);
and U8677 (N_8677,N_5090,N_6912);
and U8678 (N_8678,N_5683,N_5862);
or U8679 (N_8679,N_5344,N_5748);
or U8680 (N_8680,N_6575,N_5740);
and U8681 (N_8681,N_6824,N_5845);
nand U8682 (N_8682,N_6368,N_5820);
nor U8683 (N_8683,N_6594,N_6269);
or U8684 (N_8684,N_7007,N_7116);
or U8685 (N_8685,N_6293,N_5530);
and U8686 (N_8686,N_5298,N_5896);
or U8687 (N_8687,N_7374,N_5093);
nand U8688 (N_8688,N_6410,N_6251);
nand U8689 (N_8689,N_5300,N_6749);
and U8690 (N_8690,N_5680,N_7157);
nor U8691 (N_8691,N_5893,N_6583);
or U8692 (N_8692,N_5281,N_7050);
xnor U8693 (N_8693,N_6208,N_5266);
and U8694 (N_8694,N_6443,N_6297);
xor U8695 (N_8695,N_6818,N_6344);
nor U8696 (N_8696,N_7467,N_5318);
or U8697 (N_8697,N_7237,N_6388);
nor U8698 (N_8698,N_7108,N_5867);
nor U8699 (N_8699,N_5120,N_6915);
nand U8700 (N_8700,N_5363,N_7338);
nand U8701 (N_8701,N_5207,N_6743);
nor U8702 (N_8702,N_5136,N_6828);
nand U8703 (N_8703,N_6882,N_5137);
nor U8704 (N_8704,N_5063,N_7495);
nand U8705 (N_8705,N_6984,N_6049);
nand U8706 (N_8706,N_5332,N_6683);
or U8707 (N_8707,N_7178,N_5309);
nand U8708 (N_8708,N_5709,N_6777);
xnor U8709 (N_8709,N_6095,N_6427);
and U8710 (N_8710,N_7356,N_5246);
and U8711 (N_8711,N_6603,N_5233);
or U8712 (N_8712,N_6064,N_6294);
or U8713 (N_8713,N_5690,N_7266);
nand U8714 (N_8714,N_6927,N_5612);
and U8715 (N_8715,N_6535,N_5945);
and U8716 (N_8716,N_5112,N_6643);
xnor U8717 (N_8717,N_6394,N_5075);
nor U8718 (N_8718,N_7269,N_5735);
nor U8719 (N_8719,N_6336,N_5753);
or U8720 (N_8720,N_6988,N_6313);
and U8721 (N_8721,N_7462,N_5133);
nand U8722 (N_8722,N_6969,N_6131);
nor U8723 (N_8723,N_7285,N_5429);
xnor U8724 (N_8724,N_6178,N_7036);
nand U8725 (N_8725,N_6647,N_7170);
and U8726 (N_8726,N_5396,N_6858);
and U8727 (N_8727,N_5752,N_7256);
and U8728 (N_8728,N_6702,N_5471);
nor U8729 (N_8729,N_5549,N_7173);
and U8730 (N_8730,N_7214,N_7200);
nand U8731 (N_8731,N_6887,N_6718);
or U8732 (N_8732,N_5856,N_6097);
xor U8733 (N_8733,N_7359,N_5070);
or U8734 (N_8734,N_6333,N_5194);
nand U8735 (N_8735,N_6548,N_5718);
or U8736 (N_8736,N_5357,N_6854);
xnor U8737 (N_8737,N_6529,N_6480);
nor U8738 (N_8738,N_5692,N_5089);
nor U8739 (N_8739,N_5702,N_6553);
or U8740 (N_8740,N_7294,N_5153);
and U8741 (N_8741,N_6714,N_6115);
or U8742 (N_8742,N_6970,N_6805);
and U8743 (N_8743,N_7038,N_6723);
and U8744 (N_8744,N_5245,N_5801);
xnor U8745 (N_8745,N_6227,N_6338);
nand U8746 (N_8746,N_5159,N_7340);
and U8747 (N_8747,N_5312,N_5259);
nand U8748 (N_8748,N_6370,N_5650);
and U8749 (N_8749,N_7419,N_5973);
xor U8750 (N_8750,N_7225,N_5531);
and U8751 (N_8751,N_6806,N_6876);
or U8752 (N_8752,N_5940,N_6695);
and U8753 (N_8753,N_5558,N_7318);
and U8754 (N_8754,N_6911,N_6713);
nand U8755 (N_8755,N_5959,N_7133);
nor U8756 (N_8756,N_6319,N_7033);
or U8757 (N_8757,N_5421,N_6380);
and U8758 (N_8758,N_6852,N_5943);
nand U8759 (N_8759,N_6722,N_6423);
xnor U8760 (N_8760,N_5121,N_7017);
or U8761 (N_8761,N_5072,N_5987);
or U8762 (N_8762,N_5836,N_5588);
and U8763 (N_8763,N_7439,N_6397);
and U8764 (N_8764,N_6377,N_7053);
nand U8765 (N_8765,N_6124,N_6156);
nor U8766 (N_8766,N_7204,N_6899);
nor U8767 (N_8767,N_5112,N_7283);
xor U8768 (N_8768,N_6803,N_5621);
or U8769 (N_8769,N_6125,N_5424);
nand U8770 (N_8770,N_6771,N_7283);
nor U8771 (N_8771,N_5204,N_6427);
nand U8772 (N_8772,N_6709,N_5066);
and U8773 (N_8773,N_6614,N_5620);
nand U8774 (N_8774,N_5166,N_7177);
and U8775 (N_8775,N_6485,N_6161);
or U8776 (N_8776,N_7008,N_6416);
nand U8777 (N_8777,N_5662,N_5663);
and U8778 (N_8778,N_5546,N_7123);
nand U8779 (N_8779,N_6112,N_5837);
nor U8780 (N_8780,N_5859,N_6540);
nand U8781 (N_8781,N_5485,N_5040);
nand U8782 (N_8782,N_6737,N_5865);
nor U8783 (N_8783,N_6567,N_6911);
or U8784 (N_8784,N_6873,N_7037);
nand U8785 (N_8785,N_5165,N_5119);
nor U8786 (N_8786,N_6946,N_5606);
nand U8787 (N_8787,N_5381,N_5294);
and U8788 (N_8788,N_6323,N_5809);
nand U8789 (N_8789,N_6078,N_5206);
or U8790 (N_8790,N_6614,N_6074);
or U8791 (N_8791,N_7402,N_5622);
or U8792 (N_8792,N_6917,N_6121);
nor U8793 (N_8793,N_5380,N_5560);
nor U8794 (N_8794,N_7126,N_7090);
or U8795 (N_8795,N_7109,N_7386);
nor U8796 (N_8796,N_6153,N_5003);
nand U8797 (N_8797,N_6711,N_6656);
nand U8798 (N_8798,N_7492,N_6324);
xor U8799 (N_8799,N_6557,N_5619);
nand U8800 (N_8800,N_6013,N_6869);
nor U8801 (N_8801,N_5863,N_7169);
and U8802 (N_8802,N_6512,N_5713);
nand U8803 (N_8803,N_6405,N_6726);
and U8804 (N_8804,N_6855,N_6962);
or U8805 (N_8805,N_6734,N_6747);
nand U8806 (N_8806,N_7213,N_7445);
or U8807 (N_8807,N_5450,N_7362);
and U8808 (N_8808,N_5459,N_5422);
or U8809 (N_8809,N_6032,N_6181);
xor U8810 (N_8810,N_7127,N_6350);
nand U8811 (N_8811,N_6793,N_6880);
xnor U8812 (N_8812,N_6823,N_7435);
nor U8813 (N_8813,N_5108,N_5951);
or U8814 (N_8814,N_6425,N_6107);
and U8815 (N_8815,N_5539,N_7260);
nand U8816 (N_8816,N_6521,N_7150);
nand U8817 (N_8817,N_7427,N_5677);
xor U8818 (N_8818,N_7117,N_7259);
nor U8819 (N_8819,N_5995,N_5702);
and U8820 (N_8820,N_5516,N_7176);
nand U8821 (N_8821,N_6431,N_7385);
nor U8822 (N_8822,N_5612,N_7046);
nor U8823 (N_8823,N_5251,N_6509);
xor U8824 (N_8824,N_5505,N_5455);
or U8825 (N_8825,N_6725,N_6768);
xor U8826 (N_8826,N_6815,N_6978);
and U8827 (N_8827,N_6430,N_6055);
or U8828 (N_8828,N_6253,N_6272);
nand U8829 (N_8829,N_6320,N_5015);
xor U8830 (N_8830,N_6362,N_7111);
and U8831 (N_8831,N_6473,N_6658);
xnor U8832 (N_8832,N_6241,N_6250);
nand U8833 (N_8833,N_7388,N_6752);
nor U8834 (N_8834,N_6314,N_5438);
and U8835 (N_8835,N_7267,N_6550);
and U8836 (N_8836,N_6724,N_6638);
nor U8837 (N_8837,N_5737,N_6562);
nor U8838 (N_8838,N_7027,N_7130);
nand U8839 (N_8839,N_5293,N_6680);
or U8840 (N_8840,N_7439,N_6061);
or U8841 (N_8841,N_7433,N_6896);
and U8842 (N_8842,N_7388,N_7176);
and U8843 (N_8843,N_5042,N_5485);
and U8844 (N_8844,N_5431,N_7474);
xor U8845 (N_8845,N_7247,N_5948);
or U8846 (N_8846,N_7326,N_6248);
and U8847 (N_8847,N_5129,N_5270);
xnor U8848 (N_8848,N_7070,N_6385);
nor U8849 (N_8849,N_6625,N_7133);
nor U8850 (N_8850,N_5059,N_5095);
nand U8851 (N_8851,N_6032,N_5696);
nor U8852 (N_8852,N_5911,N_5037);
and U8853 (N_8853,N_5519,N_5377);
nor U8854 (N_8854,N_7410,N_7463);
nand U8855 (N_8855,N_6402,N_6253);
nor U8856 (N_8856,N_5603,N_6270);
xnor U8857 (N_8857,N_6774,N_5874);
or U8858 (N_8858,N_6972,N_6781);
nand U8859 (N_8859,N_5149,N_5179);
or U8860 (N_8860,N_5489,N_5730);
nor U8861 (N_8861,N_7056,N_5907);
or U8862 (N_8862,N_6028,N_6822);
or U8863 (N_8863,N_7360,N_5708);
nand U8864 (N_8864,N_7454,N_5510);
nand U8865 (N_8865,N_5308,N_5422);
xor U8866 (N_8866,N_5994,N_6907);
and U8867 (N_8867,N_7065,N_6688);
and U8868 (N_8868,N_6600,N_7350);
nor U8869 (N_8869,N_5137,N_5270);
nor U8870 (N_8870,N_5936,N_7385);
xnor U8871 (N_8871,N_6796,N_5716);
nand U8872 (N_8872,N_7002,N_5229);
nand U8873 (N_8873,N_5758,N_7447);
nand U8874 (N_8874,N_7330,N_5642);
and U8875 (N_8875,N_7138,N_6037);
nor U8876 (N_8876,N_7294,N_6193);
or U8877 (N_8877,N_7469,N_6839);
and U8878 (N_8878,N_6779,N_5619);
and U8879 (N_8879,N_7012,N_7452);
nor U8880 (N_8880,N_6598,N_5322);
and U8881 (N_8881,N_7026,N_6421);
nor U8882 (N_8882,N_5927,N_5019);
nand U8883 (N_8883,N_6245,N_5223);
nand U8884 (N_8884,N_5521,N_5497);
and U8885 (N_8885,N_5512,N_6089);
xor U8886 (N_8886,N_5003,N_6314);
nand U8887 (N_8887,N_6627,N_6167);
nor U8888 (N_8888,N_5213,N_7100);
nor U8889 (N_8889,N_7345,N_6239);
or U8890 (N_8890,N_6461,N_7480);
or U8891 (N_8891,N_6277,N_5000);
nor U8892 (N_8892,N_7036,N_6927);
xor U8893 (N_8893,N_6336,N_7473);
nor U8894 (N_8894,N_5274,N_6077);
nor U8895 (N_8895,N_5308,N_5281);
xnor U8896 (N_8896,N_6316,N_5967);
and U8897 (N_8897,N_7490,N_5904);
or U8898 (N_8898,N_6527,N_5027);
and U8899 (N_8899,N_7326,N_6285);
or U8900 (N_8900,N_7220,N_5321);
or U8901 (N_8901,N_5105,N_6940);
and U8902 (N_8902,N_6477,N_5770);
and U8903 (N_8903,N_5804,N_6728);
nor U8904 (N_8904,N_5938,N_5743);
and U8905 (N_8905,N_5816,N_6739);
nand U8906 (N_8906,N_7196,N_7320);
and U8907 (N_8907,N_6975,N_5210);
or U8908 (N_8908,N_5749,N_5325);
or U8909 (N_8909,N_5131,N_7287);
nand U8910 (N_8910,N_5921,N_5901);
nand U8911 (N_8911,N_7226,N_6061);
nor U8912 (N_8912,N_5126,N_5398);
nand U8913 (N_8913,N_6653,N_6405);
nand U8914 (N_8914,N_7183,N_6043);
nor U8915 (N_8915,N_5896,N_6852);
and U8916 (N_8916,N_6471,N_5583);
and U8917 (N_8917,N_7150,N_6737);
and U8918 (N_8918,N_6870,N_7283);
and U8919 (N_8919,N_5699,N_5924);
or U8920 (N_8920,N_6555,N_7300);
nor U8921 (N_8921,N_6861,N_6465);
nor U8922 (N_8922,N_5769,N_5931);
nand U8923 (N_8923,N_6312,N_7094);
xnor U8924 (N_8924,N_6909,N_5040);
and U8925 (N_8925,N_6373,N_7340);
nand U8926 (N_8926,N_7363,N_6299);
and U8927 (N_8927,N_5505,N_7409);
nand U8928 (N_8928,N_6420,N_5317);
and U8929 (N_8929,N_7013,N_7477);
and U8930 (N_8930,N_6378,N_5259);
nor U8931 (N_8931,N_6254,N_5688);
and U8932 (N_8932,N_6255,N_5837);
nor U8933 (N_8933,N_5634,N_5548);
xnor U8934 (N_8934,N_7484,N_6132);
xor U8935 (N_8935,N_6398,N_5186);
nand U8936 (N_8936,N_6675,N_6782);
or U8937 (N_8937,N_5614,N_6243);
nor U8938 (N_8938,N_5123,N_6235);
and U8939 (N_8939,N_7441,N_7254);
nand U8940 (N_8940,N_6361,N_5909);
nor U8941 (N_8941,N_7031,N_7261);
nand U8942 (N_8942,N_6252,N_6876);
and U8943 (N_8943,N_5161,N_6935);
xor U8944 (N_8944,N_6690,N_6612);
nand U8945 (N_8945,N_5918,N_5661);
nor U8946 (N_8946,N_5344,N_6473);
and U8947 (N_8947,N_5741,N_7210);
nor U8948 (N_8948,N_6447,N_5968);
or U8949 (N_8949,N_6689,N_6373);
or U8950 (N_8950,N_5612,N_5411);
nand U8951 (N_8951,N_5544,N_6275);
or U8952 (N_8952,N_5630,N_6908);
nand U8953 (N_8953,N_5147,N_5531);
nand U8954 (N_8954,N_5502,N_6706);
and U8955 (N_8955,N_5763,N_5703);
xor U8956 (N_8956,N_5591,N_6885);
or U8957 (N_8957,N_6034,N_6615);
nand U8958 (N_8958,N_6937,N_5117);
xnor U8959 (N_8959,N_5645,N_7239);
xnor U8960 (N_8960,N_6202,N_7086);
or U8961 (N_8961,N_6165,N_6951);
and U8962 (N_8962,N_5525,N_6875);
and U8963 (N_8963,N_5576,N_6018);
nor U8964 (N_8964,N_6078,N_5944);
nand U8965 (N_8965,N_7427,N_6228);
or U8966 (N_8966,N_5428,N_5273);
or U8967 (N_8967,N_5306,N_5568);
xor U8968 (N_8968,N_7401,N_5069);
or U8969 (N_8969,N_6647,N_7144);
nand U8970 (N_8970,N_6526,N_7156);
and U8971 (N_8971,N_6172,N_6611);
and U8972 (N_8972,N_6705,N_5367);
nor U8973 (N_8973,N_6844,N_5291);
nor U8974 (N_8974,N_5153,N_6207);
or U8975 (N_8975,N_6222,N_7277);
or U8976 (N_8976,N_5858,N_7120);
nor U8977 (N_8977,N_5158,N_6613);
nor U8978 (N_8978,N_5788,N_7060);
nand U8979 (N_8979,N_6368,N_6979);
nand U8980 (N_8980,N_7474,N_6375);
xor U8981 (N_8981,N_5809,N_5598);
nor U8982 (N_8982,N_5997,N_6765);
nor U8983 (N_8983,N_7234,N_6645);
or U8984 (N_8984,N_6953,N_6644);
or U8985 (N_8985,N_7217,N_6593);
nand U8986 (N_8986,N_5566,N_5001);
or U8987 (N_8987,N_5307,N_6481);
xor U8988 (N_8988,N_6373,N_7111);
nor U8989 (N_8989,N_5212,N_7321);
or U8990 (N_8990,N_5470,N_6167);
and U8991 (N_8991,N_5457,N_5388);
or U8992 (N_8992,N_7095,N_5980);
or U8993 (N_8993,N_6853,N_6014);
nand U8994 (N_8994,N_7277,N_6482);
nor U8995 (N_8995,N_6908,N_6119);
nor U8996 (N_8996,N_6069,N_5496);
nand U8997 (N_8997,N_6499,N_5443);
nor U8998 (N_8998,N_7069,N_7386);
xnor U8999 (N_8999,N_5924,N_6659);
nand U9000 (N_9000,N_5988,N_5894);
nand U9001 (N_9001,N_5871,N_6113);
nand U9002 (N_9002,N_5757,N_7203);
nor U9003 (N_9003,N_5946,N_7252);
nand U9004 (N_9004,N_7033,N_6291);
and U9005 (N_9005,N_6315,N_6143);
nor U9006 (N_9006,N_7488,N_6708);
or U9007 (N_9007,N_5718,N_5701);
nor U9008 (N_9008,N_6919,N_6937);
or U9009 (N_9009,N_5423,N_5369);
nand U9010 (N_9010,N_6083,N_6413);
nor U9011 (N_9011,N_6002,N_5344);
nor U9012 (N_9012,N_5449,N_5607);
nor U9013 (N_9013,N_5221,N_6010);
nand U9014 (N_9014,N_6411,N_5806);
or U9015 (N_9015,N_5608,N_7400);
and U9016 (N_9016,N_6095,N_5384);
or U9017 (N_9017,N_5960,N_6598);
nor U9018 (N_9018,N_6730,N_5141);
nand U9019 (N_9019,N_5271,N_5253);
and U9020 (N_9020,N_5842,N_6203);
and U9021 (N_9021,N_7281,N_6128);
or U9022 (N_9022,N_5872,N_6005);
and U9023 (N_9023,N_7092,N_5208);
or U9024 (N_9024,N_6533,N_5894);
nor U9025 (N_9025,N_6260,N_5776);
nand U9026 (N_9026,N_6458,N_6019);
and U9027 (N_9027,N_6675,N_6865);
or U9028 (N_9028,N_5860,N_6190);
or U9029 (N_9029,N_5690,N_5655);
or U9030 (N_9030,N_7161,N_6826);
nor U9031 (N_9031,N_6448,N_6411);
nand U9032 (N_9032,N_6297,N_6526);
nand U9033 (N_9033,N_6326,N_6481);
nor U9034 (N_9034,N_5651,N_6872);
nor U9035 (N_9035,N_6674,N_6204);
nor U9036 (N_9036,N_6346,N_5630);
nand U9037 (N_9037,N_5612,N_6111);
nand U9038 (N_9038,N_6741,N_5496);
or U9039 (N_9039,N_6178,N_6358);
and U9040 (N_9040,N_5489,N_5075);
or U9041 (N_9041,N_6628,N_6694);
or U9042 (N_9042,N_7059,N_5066);
nor U9043 (N_9043,N_5577,N_5816);
nor U9044 (N_9044,N_7218,N_6112);
nand U9045 (N_9045,N_5523,N_6135);
nor U9046 (N_9046,N_7418,N_5413);
nand U9047 (N_9047,N_5170,N_5758);
nand U9048 (N_9048,N_6623,N_5309);
nand U9049 (N_9049,N_5672,N_6423);
nand U9050 (N_9050,N_7248,N_6508);
or U9051 (N_9051,N_7203,N_6746);
or U9052 (N_9052,N_7204,N_6919);
and U9053 (N_9053,N_5055,N_5111);
or U9054 (N_9054,N_6124,N_6607);
nor U9055 (N_9055,N_5926,N_5076);
nand U9056 (N_9056,N_5174,N_5667);
nor U9057 (N_9057,N_7265,N_6360);
nand U9058 (N_9058,N_6847,N_5230);
and U9059 (N_9059,N_5384,N_6082);
nand U9060 (N_9060,N_5557,N_6800);
and U9061 (N_9061,N_6499,N_7379);
and U9062 (N_9062,N_6737,N_5860);
nand U9063 (N_9063,N_5352,N_6015);
nor U9064 (N_9064,N_5399,N_5262);
or U9065 (N_9065,N_5372,N_7428);
and U9066 (N_9066,N_6028,N_5966);
nor U9067 (N_9067,N_6040,N_7229);
and U9068 (N_9068,N_6128,N_7156);
or U9069 (N_9069,N_7330,N_6213);
nor U9070 (N_9070,N_7164,N_5282);
nand U9071 (N_9071,N_5975,N_5394);
or U9072 (N_9072,N_7478,N_6465);
nand U9073 (N_9073,N_6309,N_6223);
nor U9074 (N_9074,N_5450,N_6755);
and U9075 (N_9075,N_6389,N_5386);
or U9076 (N_9076,N_6728,N_5159);
nor U9077 (N_9077,N_6412,N_6996);
or U9078 (N_9078,N_6353,N_7477);
nand U9079 (N_9079,N_7054,N_5162);
nor U9080 (N_9080,N_6978,N_5891);
or U9081 (N_9081,N_6217,N_5527);
and U9082 (N_9082,N_5632,N_7247);
or U9083 (N_9083,N_6627,N_5556);
nand U9084 (N_9084,N_6831,N_6727);
and U9085 (N_9085,N_6809,N_5848);
xor U9086 (N_9086,N_6620,N_6457);
and U9087 (N_9087,N_5901,N_5236);
or U9088 (N_9088,N_5639,N_7053);
or U9089 (N_9089,N_6672,N_6160);
and U9090 (N_9090,N_7084,N_5468);
or U9091 (N_9091,N_5192,N_5257);
nor U9092 (N_9092,N_5889,N_6641);
nand U9093 (N_9093,N_6387,N_7062);
nor U9094 (N_9094,N_6346,N_5489);
nand U9095 (N_9095,N_7407,N_5976);
and U9096 (N_9096,N_6411,N_5054);
nor U9097 (N_9097,N_6008,N_7100);
nor U9098 (N_9098,N_6459,N_7457);
nand U9099 (N_9099,N_6723,N_6653);
and U9100 (N_9100,N_6405,N_6437);
nand U9101 (N_9101,N_6394,N_6937);
and U9102 (N_9102,N_5103,N_7440);
and U9103 (N_9103,N_5860,N_7485);
nand U9104 (N_9104,N_5414,N_6243);
nand U9105 (N_9105,N_6497,N_7002);
xor U9106 (N_9106,N_6172,N_6090);
and U9107 (N_9107,N_5169,N_6698);
and U9108 (N_9108,N_5884,N_6475);
nand U9109 (N_9109,N_6949,N_7392);
xnor U9110 (N_9110,N_5083,N_6338);
xnor U9111 (N_9111,N_5562,N_7141);
nand U9112 (N_9112,N_7336,N_6170);
xnor U9113 (N_9113,N_5421,N_5383);
and U9114 (N_9114,N_7412,N_5573);
nor U9115 (N_9115,N_6213,N_7063);
nor U9116 (N_9116,N_5636,N_5135);
or U9117 (N_9117,N_6557,N_6470);
nor U9118 (N_9118,N_5800,N_6412);
nor U9119 (N_9119,N_5877,N_6273);
nand U9120 (N_9120,N_6456,N_5321);
nand U9121 (N_9121,N_6325,N_6764);
nor U9122 (N_9122,N_6151,N_7313);
and U9123 (N_9123,N_6950,N_5519);
nor U9124 (N_9124,N_5663,N_5590);
xnor U9125 (N_9125,N_6119,N_5686);
or U9126 (N_9126,N_6740,N_6210);
nand U9127 (N_9127,N_6719,N_5414);
or U9128 (N_9128,N_6849,N_7337);
nand U9129 (N_9129,N_6396,N_6742);
and U9130 (N_9130,N_5991,N_6870);
nand U9131 (N_9131,N_6661,N_5701);
nor U9132 (N_9132,N_5367,N_5694);
or U9133 (N_9133,N_6459,N_5543);
and U9134 (N_9134,N_7499,N_6267);
nor U9135 (N_9135,N_6860,N_5092);
and U9136 (N_9136,N_6999,N_6988);
or U9137 (N_9137,N_7240,N_6448);
and U9138 (N_9138,N_6693,N_6327);
nand U9139 (N_9139,N_6880,N_7444);
nand U9140 (N_9140,N_6216,N_5738);
nand U9141 (N_9141,N_5782,N_6673);
and U9142 (N_9142,N_6010,N_6713);
nand U9143 (N_9143,N_7360,N_7065);
nand U9144 (N_9144,N_7258,N_6382);
nand U9145 (N_9145,N_5873,N_5164);
xnor U9146 (N_9146,N_6576,N_7060);
or U9147 (N_9147,N_5331,N_5124);
nor U9148 (N_9148,N_7315,N_6344);
and U9149 (N_9149,N_7400,N_5145);
nand U9150 (N_9150,N_7466,N_7189);
xnor U9151 (N_9151,N_7061,N_5859);
and U9152 (N_9152,N_5610,N_7414);
nand U9153 (N_9153,N_6938,N_6175);
nand U9154 (N_9154,N_7187,N_6037);
nand U9155 (N_9155,N_5093,N_7052);
nand U9156 (N_9156,N_7037,N_5710);
nor U9157 (N_9157,N_6531,N_6609);
and U9158 (N_9158,N_6818,N_5892);
and U9159 (N_9159,N_7183,N_5311);
and U9160 (N_9160,N_6846,N_5946);
nand U9161 (N_9161,N_6294,N_5509);
nand U9162 (N_9162,N_6685,N_5320);
or U9163 (N_9163,N_5912,N_5949);
nand U9164 (N_9164,N_6201,N_7077);
nor U9165 (N_9165,N_5075,N_5123);
nor U9166 (N_9166,N_5749,N_7462);
or U9167 (N_9167,N_5439,N_5584);
nor U9168 (N_9168,N_6957,N_6533);
or U9169 (N_9169,N_6530,N_5693);
nand U9170 (N_9170,N_5291,N_5896);
or U9171 (N_9171,N_6664,N_7216);
and U9172 (N_9172,N_6464,N_6091);
nand U9173 (N_9173,N_5861,N_5715);
or U9174 (N_9174,N_5229,N_7184);
nand U9175 (N_9175,N_6531,N_7328);
and U9176 (N_9176,N_5955,N_5045);
nor U9177 (N_9177,N_5108,N_5324);
nor U9178 (N_9178,N_7492,N_5814);
and U9179 (N_9179,N_6430,N_6747);
nor U9180 (N_9180,N_5423,N_6286);
xnor U9181 (N_9181,N_5088,N_7013);
or U9182 (N_9182,N_6056,N_5962);
xor U9183 (N_9183,N_7381,N_5666);
nand U9184 (N_9184,N_7260,N_5419);
or U9185 (N_9185,N_5527,N_5671);
nand U9186 (N_9186,N_6779,N_6738);
nand U9187 (N_9187,N_5373,N_5084);
and U9188 (N_9188,N_7109,N_5994);
nand U9189 (N_9189,N_6728,N_6161);
nand U9190 (N_9190,N_5920,N_7360);
xor U9191 (N_9191,N_6918,N_6956);
xnor U9192 (N_9192,N_6358,N_7111);
nand U9193 (N_9193,N_7143,N_6556);
and U9194 (N_9194,N_5398,N_6519);
and U9195 (N_9195,N_7377,N_5189);
nor U9196 (N_9196,N_6098,N_5713);
and U9197 (N_9197,N_5618,N_7407);
xor U9198 (N_9198,N_6162,N_5324);
or U9199 (N_9199,N_5089,N_5847);
nand U9200 (N_9200,N_6859,N_6143);
or U9201 (N_9201,N_7300,N_7317);
or U9202 (N_9202,N_5032,N_5906);
and U9203 (N_9203,N_6574,N_6501);
or U9204 (N_9204,N_6397,N_5622);
or U9205 (N_9205,N_6617,N_7135);
or U9206 (N_9206,N_5028,N_5994);
nand U9207 (N_9207,N_5804,N_5924);
nand U9208 (N_9208,N_6226,N_6819);
or U9209 (N_9209,N_6231,N_5290);
or U9210 (N_9210,N_6724,N_6560);
nand U9211 (N_9211,N_6549,N_5903);
or U9212 (N_9212,N_5788,N_5188);
and U9213 (N_9213,N_5012,N_5531);
xnor U9214 (N_9214,N_6699,N_5489);
and U9215 (N_9215,N_5920,N_5522);
and U9216 (N_9216,N_7058,N_6965);
nor U9217 (N_9217,N_5031,N_6475);
nand U9218 (N_9218,N_6822,N_5765);
nor U9219 (N_9219,N_6735,N_6707);
and U9220 (N_9220,N_7249,N_5750);
nor U9221 (N_9221,N_5973,N_6612);
and U9222 (N_9222,N_6230,N_6609);
or U9223 (N_9223,N_5602,N_6635);
nand U9224 (N_9224,N_6779,N_7021);
nor U9225 (N_9225,N_5640,N_6166);
nor U9226 (N_9226,N_5804,N_6407);
or U9227 (N_9227,N_6253,N_5000);
and U9228 (N_9228,N_6039,N_6529);
and U9229 (N_9229,N_6722,N_6897);
and U9230 (N_9230,N_6373,N_5190);
nand U9231 (N_9231,N_5932,N_7202);
and U9232 (N_9232,N_5825,N_6198);
or U9233 (N_9233,N_5373,N_6390);
nor U9234 (N_9234,N_5856,N_5290);
nand U9235 (N_9235,N_5537,N_5057);
nor U9236 (N_9236,N_6958,N_6733);
nor U9237 (N_9237,N_6148,N_5488);
nor U9238 (N_9238,N_6561,N_6856);
nor U9239 (N_9239,N_5803,N_6235);
or U9240 (N_9240,N_7301,N_5635);
and U9241 (N_9241,N_6214,N_5576);
nand U9242 (N_9242,N_6589,N_5759);
nor U9243 (N_9243,N_7398,N_5938);
nor U9244 (N_9244,N_5593,N_6935);
nor U9245 (N_9245,N_6053,N_5438);
nor U9246 (N_9246,N_7389,N_6747);
and U9247 (N_9247,N_5425,N_5264);
nor U9248 (N_9248,N_6294,N_5398);
nor U9249 (N_9249,N_5282,N_7379);
nor U9250 (N_9250,N_5188,N_7375);
nor U9251 (N_9251,N_5520,N_6091);
or U9252 (N_9252,N_7445,N_6994);
or U9253 (N_9253,N_7421,N_5030);
and U9254 (N_9254,N_6559,N_6318);
or U9255 (N_9255,N_7186,N_5571);
nor U9256 (N_9256,N_6179,N_7481);
or U9257 (N_9257,N_6036,N_6853);
or U9258 (N_9258,N_5484,N_6197);
nor U9259 (N_9259,N_6858,N_5838);
or U9260 (N_9260,N_7283,N_6115);
or U9261 (N_9261,N_6009,N_5480);
or U9262 (N_9262,N_7191,N_5249);
xor U9263 (N_9263,N_5231,N_5865);
nor U9264 (N_9264,N_7001,N_7229);
nand U9265 (N_9265,N_5787,N_6457);
xnor U9266 (N_9266,N_5769,N_5506);
nor U9267 (N_9267,N_6802,N_6758);
or U9268 (N_9268,N_5595,N_5431);
nand U9269 (N_9269,N_5092,N_5763);
and U9270 (N_9270,N_7419,N_6465);
or U9271 (N_9271,N_5810,N_6917);
and U9272 (N_9272,N_5359,N_5235);
nand U9273 (N_9273,N_5454,N_6671);
or U9274 (N_9274,N_5875,N_5512);
nand U9275 (N_9275,N_6891,N_6486);
nor U9276 (N_9276,N_6911,N_5931);
or U9277 (N_9277,N_5647,N_6324);
and U9278 (N_9278,N_5033,N_5513);
and U9279 (N_9279,N_5432,N_5656);
nor U9280 (N_9280,N_6510,N_5387);
or U9281 (N_9281,N_6203,N_7282);
xnor U9282 (N_9282,N_5754,N_5034);
nand U9283 (N_9283,N_7249,N_6768);
xnor U9284 (N_9284,N_6986,N_7301);
and U9285 (N_9285,N_5595,N_6170);
nand U9286 (N_9286,N_6934,N_7460);
and U9287 (N_9287,N_6674,N_5942);
or U9288 (N_9288,N_5148,N_6573);
xor U9289 (N_9289,N_7253,N_6008);
nand U9290 (N_9290,N_7266,N_6047);
nor U9291 (N_9291,N_6226,N_7439);
xnor U9292 (N_9292,N_7414,N_7063);
nand U9293 (N_9293,N_6231,N_5654);
xor U9294 (N_9294,N_5288,N_6279);
and U9295 (N_9295,N_5982,N_6905);
and U9296 (N_9296,N_6386,N_6913);
nand U9297 (N_9297,N_6788,N_5236);
and U9298 (N_9298,N_6002,N_7193);
and U9299 (N_9299,N_7330,N_5752);
and U9300 (N_9300,N_5702,N_6600);
or U9301 (N_9301,N_5062,N_7103);
nand U9302 (N_9302,N_5535,N_7203);
or U9303 (N_9303,N_6274,N_5154);
and U9304 (N_9304,N_7159,N_5138);
or U9305 (N_9305,N_6353,N_5849);
and U9306 (N_9306,N_5647,N_5833);
xnor U9307 (N_9307,N_5906,N_6551);
xnor U9308 (N_9308,N_6058,N_7434);
and U9309 (N_9309,N_5647,N_6540);
xnor U9310 (N_9310,N_6322,N_7263);
and U9311 (N_9311,N_5934,N_5085);
nand U9312 (N_9312,N_5184,N_6846);
or U9313 (N_9313,N_7052,N_7170);
or U9314 (N_9314,N_5127,N_5327);
xnor U9315 (N_9315,N_7243,N_6707);
nor U9316 (N_9316,N_7375,N_6317);
nor U9317 (N_9317,N_7220,N_7342);
and U9318 (N_9318,N_5908,N_5210);
nor U9319 (N_9319,N_5609,N_7114);
and U9320 (N_9320,N_5474,N_5650);
nor U9321 (N_9321,N_6890,N_6984);
nor U9322 (N_9322,N_5510,N_5832);
nor U9323 (N_9323,N_5392,N_7074);
and U9324 (N_9324,N_5513,N_7491);
nor U9325 (N_9325,N_6778,N_6743);
and U9326 (N_9326,N_6232,N_7396);
nand U9327 (N_9327,N_6799,N_7288);
nor U9328 (N_9328,N_6000,N_7444);
nor U9329 (N_9329,N_6276,N_5478);
or U9330 (N_9330,N_6749,N_6138);
or U9331 (N_9331,N_5490,N_6643);
nand U9332 (N_9332,N_5953,N_7002);
nor U9333 (N_9333,N_6578,N_5325);
or U9334 (N_9334,N_6849,N_7080);
and U9335 (N_9335,N_6276,N_5204);
and U9336 (N_9336,N_5737,N_5968);
nand U9337 (N_9337,N_7353,N_5041);
and U9338 (N_9338,N_5190,N_5894);
and U9339 (N_9339,N_5614,N_5716);
or U9340 (N_9340,N_7365,N_7439);
or U9341 (N_9341,N_7317,N_5613);
xnor U9342 (N_9342,N_5680,N_6559);
or U9343 (N_9343,N_6480,N_6196);
nor U9344 (N_9344,N_6016,N_7358);
xor U9345 (N_9345,N_7131,N_5510);
nand U9346 (N_9346,N_6917,N_6772);
or U9347 (N_9347,N_6888,N_6134);
xnor U9348 (N_9348,N_6162,N_6399);
nor U9349 (N_9349,N_5973,N_7045);
nand U9350 (N_9350,N_6130,N_5642);
xnor U9351 (N_9351,N_5731,N_5502);
xor U9352 (N_9352,N_5694,N_5696);
and U9353 (N_9353,N_7271,N_5755);
nand U9354 (N_9354,N_5593,N_7115);
nor U9355 (N_9355,N_7183,N_6967);
or U9356 (N_9356,N_6087,N_7372);
nor U9357 (N_9357,N_6624,N_6009);
xnor U9358 (N_9358,N_6220,N_6383);
or U9359 (N_9359,N_7114,N_6154);
or U9360 (N_9360,N_6540,N_5403);
nor U9361 (N_9361,N_6590,N_5229);
nor U9362 (N_9362,N_5604,N_5631);
or U9363 (N_9363,N_5509,N_5813);
or U9364 (N_9364,N_5599,N_7086);
nand U9365 (N_9365,N_5549,N_6976);
nor U9366 (N_9366,N_7365,N_7181);
nor U9367 (N_9367,N_5098,N_5602);
nand U9368 (N_9368,N_5007,N_7099);
or U9369 (N_9369,N_7022,N_5948);
or U9370 (N_9370,N_6326,N_6704);
nand U9371 (N_9371,N_6924,N_6591);
and U9372 (N_9372,N_7000,N_6075);
nand U9373 (N_9373,N_7416,N_6655);
nor U9374 (N_9374,N_7070,N_6513);
or U9375 (N_9375,N_7061,N_6446);
and U9376 (N_9376,N_7459,N_7222);
and U9377 (N_9377,N_6616,N_6068);
nor U9378 (N_9378,N_6146,N_6160);
nor U9379 (N_9379,N_7062,N_5256);
nor U9380 (N_9380,N_6992,N_5634);
and U9381 (N_9381,N_7237,N_5311);
and U9382 (N_9382,N_5026,N_6594);
or U9383 (N_9383,N_7357,N_7251);
and U9384 (N_9384,N_6682,N_5337);
nand U9385 (N_9385,N_6711,N_6556);
nor U9386 (N_9386,N_6728,N_6627);
or U9387 (N_9387,N_5721,N_5379);
nor U9388 (N_9388,N_6567,N_6056);
nor U9389 (N_9389,N_5591,N_5946);
xor U9390 (N_9390,N_5912,N_6304);
or U9391 (N_9391,N_6926,N_5772);
nand U9392 (N_9392,N_6704,N_7249);
and U9393 (N_9393,N_6128,N_7320);
nand U9394 (N_9394,N_6301,N_5686);
nor U9395 (N_9395,N_6773,N_5059);
xor U9396 (N_9396,N_7281,N_5903);
nor U9397 (N_9397,N_7236,N_6977);
nor U9398 (N_9398,N_5844,N_5615);
and U9399 (N_9399,N_6125,N_7066);
nand U9400 (N_9400,N_5763,N_7084);
or U9401 (N_9401,N_5480,N_6019);
and U9402 (N_9402,N_6932,N_6621);
nand U9403 (N_9403,N_6114,N_5328);
nand U9404 (N_9404,N_6630,N_5624);
and U9405 (N_9405,N_6451,N_5047);
nor U9406 (N_9406,N_6583,N_5180);
nor U9407 (N_9407,N_6971,N_5059);
xnor U9408 (N_9408,N_5770,N_7234);
or U9409 (N_9409,N_5853,N_6857);
and U9410 (N_9410,N_6280,N_5192);
and U9411 (N_9411,N_5604,N_7182);
or U9412 (N_9412,N_5059,N_7276);
nand U9413 (N_9413,N_7171,N_5990);
and U9414 (N_9414,N_6571,N_5001);
or U9415 (N_9415,N_6893,N_6873);
nand U9416 (N_9416,N_7217,N_5153);
nand U9417 (N_9417,N_7308,N_5293);
nand U9418 (N_9418,N_7068,N_5324);
nand U9419 (N_9419,N_6989,N_7149);
and U9420 (N_9420,N_7006,N_6057);
or U9421 (N_9421,N_7117,N_7361);
or U9422 (N_9422,N_5178,N_5513);
and U9423 (N_9423,N_5667,N_5711);
nor U9424 (N_9424,N_6834,N_5955);
or U9425 (N_9425,N_7017,N_6715);
nand U9426 (N_9426,N_7495,N_7106);
nand U9427 (N_9427,N_6126,N_6930);
or U9428 (N_9428,N_6416,N_7269);
and U9429 (N_9429,N_6029,N_7122);
nand U9430 (N_9430,N_6774,N_7253);
nor U9431 (N_9431,N_7289,N_6540);
or U9432 (N_9432,N_6460,N_5837);
or U9433 (N_9433,N_6541,N_5048);
nor U9434 (N_9434,N_5678,N_6093);
nand U9435 (N_9435,N_5013,N_5231);
or U9436 (N_9436,N_7197,N_5890);
nand U9437 (N_9437,N_7362,N_7489);
or U9438 (N_9438,N_5207,N_5694);
or U9439 (N_9439,N_6388,N_6422);
and U9440 (N_9440,N_6852,N_6249);
or U9441 (N_9441,N_5386,N_6475);
or U9442 (N_9442,N_5784,N_7122);
nor U9443 (N_9443,N_7492,N_7434);
and U9444 (N_9444,N_5578,N_6297);
nand U9445 (N_9445,N_5670,N_6347);
nor U9446 (N_9446,N_5028,N_6057);
and U9447 (N_9447,N_7009,N_6839);
nor U9448 (N_9448,N_7145,N_5715);
nand U9449 (N_9449,N_5884,N_7253);
nor U9450 (N_9450,N_5036,N_5089);
xnor U9451 (N_9451,N_7068,N_5146);
or U9452 (N_9452,N_5689,N_5055);
or U9453 (N_9453,N_5526,N_5955);
or U9454 (N_9454,N_7462,N_6829);
nand U9455 (N_9455,N_7421,N_5944);
nor U9456 (N_9456,N_7363,N_5704);
nand U9457 (N_9457,N_7333,N_6049);
and U9458 (N_9458,N_5876,N_6645);
xor U9459 (N_9459,N_5535,N_7173);
nor U9460 (N_9460,N_6738,N_5881);
or U9461 (N_9461,N_6722,N_6533);
or U9462 (N_9462,N_6318,N_7110);
and U9463 (N_9463,N_7271,N_7376);
and U9464 (N_9464,N_5252,N_5302);
nor U9465 (N_9465,N_5327,N_6261);
nand U9466 (N_9466,N_5032,N_6599);
xor U9467 (N_9467,N_5945,N_5984);
and U9468 (N_9468,N_6434,N_7329);
and U9469 (N_9469,N_5185,N_6596);
and U9470 (N_9470,N_6955,N_5368);
nor U9471 (N_9471,N_5156,N_6054);
nand U9472 (N_9472,N_5951,N_5721);
nor U9473 (N_9473,N_7259,N_6353);
or U9474 (N_9474,N_6919,N_5072);
and U9475 (N_9475,N_5653,N_7418);
nand U9476 (N_9476,N_6188,N_7157);
or U9477 (N_9477,N_7263,N_6351);
nand U9478 (N_9478,N_5730,N_5852);
and U9479 (N_9479,N_7451,N_5018);
and U9480 (N_9480,N_5808,N_5058);
nand U9481 (N_9481,N_5805,N_5258);
nor U9482 (N_9482,N_7227,N_6245);
nand U9483 (N_9483,N_6461,N_5434);
nand U9484 (N_9484,N_5612,N_6648);
nor U9485 (N_9485,N_5111,N_6734);
or U9486 (N_9486,N_6548,N_6796);
xor U9487 (N_9487,N_7428,N_5384);
or U9488 (N_9488,N_6363,N_6293);
nor U9489 (N_9489,N_5967,N_5416);
nor U9490 (N_9490,N_6348,N_7023);
xor U9491 (N_9491,N_5305,N_5584);
xnor U9492 (N_9492,N_5439,N_6095);
nand U9493 (N_9493,N_6419,N_5083);
nor U9494 (N_9494,N_6194,N_5312);
and U9495 (N_9495,N_6719,N_6842);
nor U9496 (N_9496,N_6609,N_7481);
xnor U9497 (N_9497,N_7457,N_6951);
or U9498 (N_9498,N_6892,N_6889);
or U9499 (N_9499,N_5777,N_5273);
nand U9500 (N_9500,N_5416,N_6118);
nand U9501 (N_9501,N_5422,N_5854);
nand U9502 (N_9502,N_5222,N_5468);
nand U9503 (N_9503,N_7194,N_7313);
and U9504 (N_9504,N_5955,N_6796);
or U9505 (N_9505,N_6204,N_5623);
and U9506 (N_9506,N_6169,N_6881);
or U9507 (N_9507,N_6408,N_5366);
or U9508 (N_9508,N_5839,N_7292);
nand U9509 (N_9509,N_6173,N_5866);
or U9510 (N_9510,N_5337,N_5906);
nor U9511 (N_9511,N_5367,N_5468);
or U9512 (N_9512,N_5857,N_6510);
or U9513 (N_9513,N_5810,N_7007);
or U9514 (N_9514,N_5274,N_6142);
nand U9515 (N_9515,N_6004,N_6360);
and U9516 (N_9516,N_5962,N_5929);
and U9517 (N_9517,N_5858,N_6212);
or U9518 (N_9518,N_7488,N_7385);
nor U9519 (N_9519,N_5312,N_6315);
and U9520 (N_9520,N_6639,N_6482);
or U9521 (N_9521,N_6269,N_6037);
nand U9522 (N_9522,N_6620,N_6984);
and U9523 (N_9523,N_5296,N_5531);
nor U9524 (N_9524,N_5254,N_6499);
nand U9525 (N_9525,N_6201,N_7483);
nand U9526 (N_9526,N_5996,N_5747);
nor U9527 (N_9527,N_5809,N_5479);
nor U9528 (N_9528,N_5267,N_5166);
xor U9529 (N_9529,N_6567,N_7105);
nor U9530 (N_9530,N_6787,N_7232);
and U9531 (N_9531,N_6964,N_7293);
nor U9532 (N_9532,N_6534,N_6557);
xnor U9533 (N_9533,N_5123,N_6472);
nand U9534 (N_9534,N_6123,N_6949);
and U9535 (N_9535,N_5283,N_7063);
nand U9536 (N_9536,N_6064,N_6886);
or U9537 (N_9537,N_7004,N_6847);
or U9538 (N_9538,N_6070,N_5906);
or U9539 (N_9539,N_5507,N_5680);
nor U9540 (N_9540,N_6179,N_7391);
or U9541 (N_9541,N_5754,N_7056);
nor U9542 (N_9542,N_6987,N_7339);
and U9543 (N_9543,N_7083,N_6616);
nand U9544 (N_9544,N_5812,N_6420);
and U9545 (N_9545,N_7126,N_5036);
or U9546 (N_9546,N_5494,N_7315);
xor U9547 (N_9547,N_6165,N_5572);
nor U9548 (N_9548,N_5238,N_7397);
and U9549 (N_9549,N_5843,N_6851);
xor U9550 (N_9550,N_6053,N_6825);
and U9551 (N_9551,N_6380,N_6732);
xnor U9552 (N_9552,N_6806,N_5037);
nand U9553 (N_9553,N_5149,N_6577);
nor U9554 (N_9554,N_6220,N_5163);
nand U9555 (N_9555,N_6473,N_6173);
xor U9556 (N_9556,N_6085,N_5988);
and U9557 (N_9557,N_7136,N_5143);
nor U9558 (N_9558,N_5042,N_6695);
nor U9559 (N_9559,N_6058,N_5968);
nor U9560 (N_9560,N_6020,N_7042);
and U9561 (N_9561,N_5973,N_7101);
or U9562 (N_9562,N_7086,N_6642);
nand U9563 (N_9563,N_5370,N_6624);
or U9564 (N_9564,N_6244,N_5260);
xor U9565 (N_9565,N_6162,N_6650);
and U9566 (N_9566,N_6687,N_6597);
nor U9567 (N_9567,N_5082,N_7363);
nand U9568 (N_9568,N_6284,N_5430);
or U9569 (N_9569,N_5424,N_6348);
or U9570 (N_9570,N_5216,N_6017);
nand U9571 (N_9571,N_7291,N_6243);
nand U9572 (N_9572,N_5189,N_5541);
or U9573 (N_9573,N_6399,N_6513);
nor U9574 (N_9574,N_7316,N_6023);
and U9575 (N_9575,N_7339,N_6434);
and U9576 (N_9576,N_6787,N_6249);
nand U9577 (N_9577,N_6007,N_6864);
or U9578 (N_9578,N_6048,N_6150);
and U9579 (N_9579,N_5457,N_6477);
xnor U9580 (N_9580,N_7292,N_6667);
nor U9581 (N_9581,N_6863,N_5476);
or U9582 (N_9582,N_7489,N_7153);
nand U9583 (N_9583,N_5694,N_6360);
nor U9584 (N_9584,N_6197,N_6889);
nand U9585 (N_9585,N_5567,N_5081);
or U9586 (N_9586,N_7206,N_6425);
xor U9587 (N_9587,N_5894,N_5250);
and U9588 (N_9588,N_6998,N_7127);
nand U9589 (N_9589,N_6983,N_6434);
and U9590 (N_9590,N_5364,N_5583);
nor U9591 (N_9591,N_5162,N_6843);
nand U9592 (N_9592,N_7106,N_6262);
nor U9593 (N_9593,N_6919,N_6459);
or U9594 (N_9594,N_5362,N_5147);
nor U9595 (N_9595,N_6318,N_5835);
nor U9596 (N_9596,N_5999,N_5404);
nand U9597 (N_9597,N_6135,N_5253);
nor U9598 (N_9598,N_6618,N_5075);
nand U9599 (N_9599,N_5832,N_6127);
nand U9600 (N_9600,N_7345,N_5932);
and U9601 (N_9601,N_6792,N_5498);
nand U9602 (N_9602,N_6847,N_7055);
and U9603 (N_9603,N_5558,N_7002);
nand U9604 (N_9604,N_7189,N_6440);
and U9605 (N_9605,N_7146,N_6732);
or U9606 (N_9606,N_7044,N_5048);
nor U9607 (N_9607,N_5267,N_6536);
and U9608 (N_9608,N_5407,N_6408);
xor U9609 (N_9609,N_7319,N_6202);
or U9610 (N_9610,N_5167,N_6360);
or U9611 (N_9611,N_5630,N_6956);
nor U9612 (N_9612,N_6041,N_5275);
nor U9613 (N_9613,N_6583,N_7226);
or U9614 (N_9614,N_5629,N_5786);
xnor U9615 (N_9615,N_5603,N_6827);
nand U9616 (N_9616,N_7408,N_6529);
nor U9617 (N_9617,N_6287,N_7123);
and U9618 (N_9618,N_7405,N_5895);
or U9619 (N_9619,N_5013,N_5080);
or U9620 (N_9620,N_5668,N_5585);
nor U9621 (N_9621,N_7446,N_5918);
nand U9622 (N_9622,N_6455,N_5574);
nor U9623 (N_9623,N_6396,N_6789);
or U9624 (N_9624,N_6368,N_7131);
nor U9625 (N_9625,N_7156,N_5611);
and U9626 (N_9626,N_6360,N_5068);
nor U9627 (N_9627,N_6418,N_5349);
and U9628 (N_9628,N_7389,N_7287);
nor U9629 (N_9629,N_7265,N_6355);
or U9630 (N_9630,N_7258,N_7085);
nand U9631 (N_9631,N_6260,N_5306);
nor U9632 (N_9632,N_6579,N_5287);
nor U9633 (N_9633,N_6961,N_6600);
or U9634 (N_9634,N_6239,N_7311);
nand U9635 (N_9635,N_6014,N_7428);
or U9636 (N_9636,N_6122,N_5454);
nand U9637 (N_9637,N_6058,N_6043);
or U9638 (N_9638,N_7218,N_6657);
nor U9639 (N_9639,N_5531,N_6394);
or U9640 (N_9640,N_7190,N_7096);
nand U9641 (N_9641,N_5809,N_5898);
and U9642 (N_9642,N_5375,N_6906);
xor U9643 (N_9643,N_7352,N_5562);
nor U9644 (N_9644,N_5504,N_7137);
nand U9645 (N_9645,N_5014,N_6702);
or U9646 (N_9646,N_6303,N_5561);
or U9647 (N_9647,N_6342,N_7239);
or U9648 (N_9648,N_6237,N_6108);
and U9649 (N_9649,N_6111,N_5022);
nand U9650 (N_9650,N_6693,N_5043);
nor U9651 (N_9651,N_6723,N_5576);
nor U9652 (N_9652,N_7185,N_6043);
nor U9653 (N_9653,N_5122,N_6901);
xnor U9654 (N_9654,N_6846,N_6275);
xor U9655 (N_9655,N_5025,N_6596);
xnor U9656 (N_9656,N_6821,N_5092);
nor U9657 (N_9657,N_7025,N_6353);
or U9658 (N_9658,N_5835,N_6691);
nor U9659 (N_9659,N_7293,N_5878);
nand U9660 (N_9660,N_5416,N_5065);
nand U9661 (N_9661,N_5399,N_6913);
and U9662 (N_9662,N_6072,N_5782);
nand U9663 (N_9663,N_6042,N_7023);
nand U9664 (N_9664,N_5060,N_7443);
nor U9665 (N_9665,N_7460,N_6911);
and U9666 (N_9666,N_6581,N_5473);
nand U9667 (N_9667,N_6130,N_7109);
and U9668 (N_9668,N_6107,N_5925);
nand U9669 (N_9669,N_6022,N_5505);
nand U9670 (N_9670,N_5282,N_7481);
nor U9671 (N_9671,N_7185,N_6569);
nand U9672 (N_9672,N_5584,N_7311);
nor U9673 (N_9673,N_5344,N_7395);
or U9674 (N_9674,N_6246,N_5479);
nand U9675 (N_9675,N_6216,N_6800);
or U9676 (N_9676,N_6268,N_5087);
xor U9677 (N_9677,N_7370,N_6177);
xnor U9678 (N_9678,N_6686,N_5815);
nor U9679 (N_9679,N_5132,N_5486);
xor U9680 (N_9680,N_5707,N_7420);
nand U9681 (N_9681,N_5951,N_6371);
or U9682 (N_9682,N_7274,N_5369);
and U9683 (N_9683,N_6443,N_5064);
or U9684 (N_9684,N_7418,N_6147);
nor U9685 (N_9685,N_6131,N_6157);
and U9686 (N_9686,N_6886,N_5083);
nand U9687 (N_9687,N_6028,N_5791);
nand U9688 (N_9688,N_5199,N_6915);
nand U9689 (N_9689,N_6614,N_6752);
nor U9690 (N_9690,N_7139,N_5924);
nand U9691 (N_9691,N_6252,N_5974);
nand U9692 (N_9692,N_6595,N_5175);
or U9693 (N_9693,N_5938,N_7124);
xnor U9694 (N_9694,N_6641,N_6715);
nor U9695 (N_9695,N_5782,N_5237);
and U9696 (N_9696,N_5552,N_7011);
nand U9697 (N_9697,N_6823,N_5871);
and U9698 (N_9698,N_7385,N_6606);
nand U9699 (N_9699,N_5213,N_5530);
nand U9700 (N_9700,N_6387,N_6121);
and U9701 (N_9701,N_5943,N_5435);
or U9702 (N_9702,N_5202,N_5702);
xnor U9703 (N_9703,N_5804,N_6121);
and U9704 (N_9704,N_5233,N_5199);
xor U9705 (N_9705,N_5990,N_6475);
nand U9706 (N_9706,N_7076,N_7355);
nand U9707 (N_9707,N_5528,N_5588);
nor U9708 (N_9708,N_6483,N_6356);
or U9709 (N_9709,N_6432,N_7287);
or U9710 (N_9710,N_7342,N_7179);
and U9711 (N_9711,N_5688,N_5702);
or U9712 (N_9712,N_7257,N_5475);
nor U9713 (N_9713,N_5173,N_5664);
nor U9714 (N_9714,N_7467,N_6226);
nand U9715 (N_9715,N_6703,N_6978);
and U9716 (N_9716,N_6213,N_6110);
nor U9717 (N_9717,N_6313,N_6049);
nor U9718 (N_9718,N_7239,N_5703);
and U9719 (N_9719,N_5355,N_5991);
nor U9720 (N_9720,N_5250,N_6485);
nor U9721 (N_9721,N_6752,N_6481);
xnor U9722 (N_9722,N_6627,N_7316);
nand U9723 (N_9723,N_5628,N_7199);
nor U9724 (N_9724,N_5597,N_7308);
nor U9725 (N_9725,N_6923,N_5517);
nor U9726 (N_9726,N_5667,N_5994);
nand U9727 (N_9727,N_6469,N_6853);
or U9728 (N_9728,N_6089,N_6406);
nand U9729 (N_9729,N_5617,N_5625);
or U9730 (N_9730,N_6510,N_7218);
nand U9731 (N_9731,N_5371,N_6980);
nand U9732 (N_9732,N_7102,N_5608);
nor U9733 (N_9733,N_6036,N_6483);
and U9734 (N_9734,N_7080,N_7483);
or U9735 (N_9735,N_5421,N_7225);
xnor U9736 (N_9736,N_5022,N_6095);
xnor U9737 (N_9737,N_5130,N_5460);
or U9738 (N_9738,N_5059,N_6183);
xor U9739 (N_9739,N_7241,N_6532);
nand U9740 (N_9740,N_5632,N_6510);
or U9741 (N_9741,N_5773,N_5961);
nand U9742 (N_9742,N_6999,N_6335);
xor U9743 (N_9743,N_7420,N_7317);
nand U9744 (N_9744,N_6464,N_5415);
or U9745 (N_9745,N_6754,N_7036);
and U9746 (N_9746,N_5699,N_5613);
nand U9747 (N_9747,N_6188,N_6412);
or U9748 (N_9748,N_5903,N_5734);
or U9749 (N_9749,N_5190,N_6283);
nand U9750 (N_9750,N_6873,N_6876);
or U9751 (N_9751,N_5355,N_6359);
or U9752 (N_9752,N_6137,N_7086);
and U9753 (N_9753,N_7340,N_5050);
and U9754 (N_9754,N_5059,N_5192);
or U9755 (N_9755,N_6330,N_6264);
nor U9756 (N_9756,N_5324,N_6719);
and U9757 (N_9757,N_6947,N_5082);
or U9758 (N_9758,N_5741,N_6872);
and U9759 (N_9759,N_6070,N_5073);
or U9760 (N_9760,N_7284,N_7269);
xor U9761 (N_9761,N_5835,N_6698);
or U9762 (N_9762,N_7314,N_6790);
and U9763 (N_9763,N_5015,N_5560);
and U9764 (N_9764,N_5565,N_6688);
and U9765 (N_9765,N_5095,N_5334);
xnor U9766 (N_9766,N_6358,N_5249);
or U9767 (N_9767,N_6029,N_7463);
nor U9768 (N_9768,N_5281,N_5617);
xor U9769 (N_9769,N_5222,N_6546);
nand U9770 (N_9770,N_6925,N_6722);
nor U9771 (N_9771,N_6519,N_6697);
nand U9772 (N_9772,N_6606,N_6674);
nor U9773 (N_9773,N_5397,N_5541);
nand U9774 (N_9774,N_7048,N_5873);
nand U9775 (N_9775,N_7461,N_6849);
nand U9776 (N_9776,N_6996,N_5621);
nand U9777 (N_9777,N_5712,N_5591);
or U9778 (N_9778,N_6948,N_6418);
nor U9779 (N_9779,N_6818,N_7206);
and U9780 (N_9780,N_5055,N_5165);
nor U9781 (N_9781,N_6999,N_7387);
or U9782 (N_9782,N_5589,N_5525);
or U9783 (N_9783,N_7147,N_6630);
nor U9784 (N_9784,N_5595,N_6719);
nor U9785 (N_9785,N_5282,N_5822);
and U9786 (N_9786,N_6596,N_7425);
or U9787 (N_9787,N_6820,N_6443);
and U9788 (N_9788,N_6101,N_5487);
nor U9789 (N_9789,N_6252,N_6244);
nor U9790 (N_9790,N_6274,N_7439);
and U9791 (N_9791,N_6406,N_5579);
or U9792 (N_9792,N_6612,N_6327);
or U9793 (N_9793,N_5126,N_6756);
and U9794 (N_9794,N_5379,N_6114);
or U9795 (N_9795,N_5558,N_6483);
or U9796 (N_9796,N_6471,N_6347);
or U9797 (N_9797,N_6596,N_6765);
and U9798 (N_9798,N_5177,N_5406);
or U9799 (N_9799,N_5323,N_5306);
nand U9800 (N_9800,N_6183,N_7151);
nor U9801 (N_9801,N_7343,N_5672);
nand U9802 (N_9802,N_6547,N_6266);
nor U9803 (N_9803,N_6255,N_5192);
or U9804 (N_9804,N_5680,N_5408);
and U9805 (N_9805,N_5270,N_7267);
and U9806 (N_9806,N_7132,N_5582);
nand U9807 (N_9807,N_5014,N_7376);
nor U9808 (N_9808,N_5891,N_5074);
xnor U9809 (N_9809,N_7438,N_7325);
nor U9810 (N_9810,N_6369,N_5792);
or U9811 (N_9811,N_7423,N_5699);
and U9812 (N_9812,N_6845,N_6543);
nand U9813 (N_9813,N_6140,N_6161);
nand U9814 (N_9814,N_5779,N_5457);
nand U9815 (N_9815,N_7323,N_7476);
and U9816 (N_9816,N_5896,N_6673);
xnor U9817 (N_9817,N_6147,N_7429);
nor U9818 (N_9818,N_7132,N_6292);
nor U9819 (N_9819,N_5790,N_5314);
nand U9820 (N_9820,N_7069,N_6540);
nand U9821 (N_9821,N_7155,N_5621);
nand U9822 (N_9822,N_5594,N_5782);
or U9823 (N_9823,N_7172,N_5311);
nand U9824 (N_9824,N_6421,N_6645);
nor U9825 (N_9825,N_6432,N_5466);
nor U9826 (N_9826,N_5880,N_5370);
xnor U9827 (N_9827,N_6851,N_6620);
or U9828 (N_9828,N_5390,N_6916);
nor U9829 (N_9829,N_5141,N_6553);
and U9830 (N_9830,N_5722,N_5317);
or U9831 (N_9831,N_5671,N_7423);
and U9832 (N_9832,N_5353,N_6267);
xor U9833 (N_9833,N_5015,N_5332);
nand U9834 (N_9834,N_7428,N_6016);
nor U9835 (N_9835,N_6236,N_5759);
nor U9836 (N_9836,N_5355,N_7341);
xor U9837 (N_9837,N_6783,N_6221);
nand U9838 (N_9838,N_7208,N_5609);
or U9839 (N_9839,N_7483,N_5843);
or U9840 (N_9840,N_5666,N_5146);
nor U9841 (N_9841,N_6423,N_7077);
nor U9842 (N_9842,N_5991,N_6338);
or U9843 (N_9843,N_5474,N_6410);
and U9844 (N_9844,N_6344,N_6626);
xnor U9845 (N_9845,N_6101,N_7103);
and U9846 (N_9846,N_5433,N_6710);
or U9847 (N_9847,N_5429,N_7166);
nand U9848 (N_9848,N_7498,N_5563);
and U9849 (N_9849,N_6689,N_7050);
or U9850 (N_9850,N_6995,N_5109);
and U9851 (N_9851,N_6550,N_5592);
xnor U9852 (N_9852,N_5001,N_6210);
and U9853 (N_9853,N_5372,N_6644);
or U9854 (N_9854,N_5387,N_6936);
and U9855 (N_9855,N_5063,N_5761);
nor U9856 (N_9856,N_6388,N_7011);
xnor U9857 (N_9857,N_7276,N_7225);
nor U9858 (N_9858,N_5494,N_7213);
and U9859 (N_9859,N_6779,N_6846);
or U9860 (N_9860,N_7359,N_6071);
or U9861 (N_9861,N_6311,N_6735);
nor U9862 (N_9862,N_5169,N_5831);
or U9863 (N_9863,N_5112,N_6205);
or U9864 (N_9864,N_7475,N_5486);
nor U9865 (N_9865,N_5564,N_7064);
nand U9866 (N_9866,N_6554,N_5945);
or U9867 (N_9867,N_5865,N_5538);
nand U9868 (N_9868,N_7036,N_5582);
or U9869 (N_9869,N_5716,N_6387);
nand U9870 (N_9870,N_6198,N_5560);
nor U9871 (N_9871,N_6047,N_5239);
nor U9872 (N_9872,N_5345,N_7341);
nand U9873 (N_9873,N_5734,N_7327);
nor U9874 (N_9874,N_6865,N_5932);
xor U9875 (N_9875,N_6883,N_7020);
nor U9876 (N_9876,N_6971,N_5893);
or U9877 (N_9877,N_5934,N_6045);
nand U9878 (N_9878,N_5361,N_6831);
nand U9879 (N_9879,N_5399,N_7155);
nand U9880 (N_9880,N_7061,N_6441);
nor U9881 (N_9881,N_5576,N_5305);
and U9882 (N_9882,N_6522,N_6304);
nand U9883 (N_9883,N_6632,N_6698);
and U9884 (N_9884,N_5339,N_5087);
nor U9885 (N_9885,N_5593,N_5411);
and U9886 (N_9886,N_7352,N_7431);
nand U9887 (N_9887,N_5602,N_6669);
and U9888 (N_9888,N_6762,N_6507);
nor U9889 (N_9889,N_6789,N_6298);
or U9890 (N_9890,N_7477,N_6738);
nand U9891 (N_9891,N_5490,N_5860);
and U9892 (N_9892,N_5495,N_5253);
or U9893 (N_9893,N_7065,N_6696);
nor U9894 (N_9894,N_5752,N_6647);
xnor U9895 (N_9895,N_7099,N_6609);
or U9896 (N_9896,N_6066,N_5940);
or U9897 (N_9897,N_7233,N_6901);
nor U9898 (N_9898,N_6820,N_7227);
nand U9899 (N_9899,N_5669,N_6803);
nand U9900 (N_9900,N_6979,N_5193);
nor U9901 (N_9901,N_7258,N_6365);
or U9902 (N_9902,N_6703,N_6006);
nand U9903 (N_9903,N_5435,N_6585);
and U9904 (N_9904,N_6839,N_6117);
and U9905 (N_9905,N_6942,N_7020);
xor U9906 (N_9906,N_5803,N_7185);
nor U9907 (N_9907,N_6877,N_7356);
and U9908 (N_9908,N_5184,N_5103);
and U9909 (N_9909,N_6374,N_7310);
or U9910 (N_9910,N_5452,N_5979);
nor U9911 (N_9911,N_6432,N_7035);
xnor U9912 (N_9912,N_6137,N_5844);
and U9913 (N_9913,N_6427,N_7117);
nor U9914 (N_9914,N_6354,N_6585);
nand U9915 (N_9915,N_5394,N_6126);
nor U9916 (N_9916,N_5780,N_6831);
nor U9917 (N_9917,N_5024,N_7108);
nor U9918 (N_9918,N_7107,N_7228);
and U9919 (N_9919,N_6529,N_6519);
or U9920 (N_9920,N_7046,N_7306);
nand U9921 (N_9921,N_6345,N_5211);
nand U9922 (N_9922,N_5613,N_7496);
xor U9923 (N_9923,N_5642,N_5460);
or U9924 (N_9924,N_6627,N_7171);
nor U9925 (N_9925,N_7252,N_5722);
or U9926 (N_9926,N_5439,N_6863);
or U9927 (N_9927,N_7108,N_5856);
or U9928 (N_9928,N_6096,N_7070);
nor U9929 (N_9929,N_7244,N_6312);
xnor U9930 (N_9930,N_6478,N_5244);
nand U9931 (N_9931,N_5887,N_5857);
nand U9932 (N_9932,N_5935,N_5182);
and U9933 (N_9933,N_6311,N_6714);
xor U9934 (N_9934,N_7235,N_6034);
nand U9935 (N_9935,N_5137,N_6708);
or U9936 (N_9936,N_6039,N_6520);
nor U9937 (N_9937,N_6383,N_6732);
xnor U9938 (N_9938,N_6265,N_6140);
and U9939 (N_9939,N_7286,N_6527);
or U9940 (N_9940,N_6097,N_5269);
nand U9941 (N_9941,N_7177,N_7067);
nand U9942 (N_9942,N_5679,N_7338);
nand U9943 (N_9943,N_6606,N_6072);
nor U9944 (N_9944,N_5933,N_5203);
xor U9945 (N_9945,N_6244,N_5084);
and U9946 (N_9946,N_5039,N_7121);
and U9947 (N_9947,N_6078,N_5952);
or U9948 (N_9948,N_7036,N_6090);
nand U9949 (N_9949,N_7281,N_5511);
nand U9950 (N_9950,N_7359,N_7469);
and U9951 (N_9951,N_6095,N_5640);
and U9952 (N_9952,N_7340,N_6945);
nand U9953 (N_9953,N_5289,N_6386);
and U9954 (N_9954,N_5855,N_6149);
nand U9955 (N_9955,N_5242,N_5957);
and U9956 (N_9956,N_5381,N_6994);
xor U9957 (N_9957,N_6971,N_6105);
nor U9958 (N_9958,N_6769,N_5754);
nand U9959 (N_9959,N_6863,N_7318);
nand U9960 (N_9960,N_6842,N_7322);
or U9961 (N_9961,N_7451,N_7268);
nor U9962 (N_9962,N_7049,N_7457);
and U9963 (N_9963,N_7411,N_5280);
nor U9964 (N_9964,N_7282,N_6104);
nor U9965 (N_9965,N_6841,N_5565);
xnor U9966 (N_9966,N_5413,N_7209);
nor U9967 (N_9967,N_6474,N_6591);
nand U9968 (N_9968,N_5435,N_5827);
or U9969 (N_9969,N_5613,N_5346);
or U9970 (N_9970,N_6143,N_6399);
nand U9971 (N_9971,N_6866,N_6924);
or U9972 (N_9972,N_5310,N_5157);
or U9973 (N_9973,N_6809,N_6186);
and U9974 (N_9974,N_7277,N_6480);
or U9975 (N_9975,N_6058,N_7072);
or U9976 (N_9976,N_6681,N_6359);
nand U9977 (N_9977,N_5190,N_6212);
xor U9978 (N_9978,N_5255,N_6120);
nor U9979 (N_9979,N_5091,N_7096);
nor U9980 (N_9980,N_5818,N_7031);
and U9981 (N_9981,N_7077,N_6311);
nand U9982 (N_9982,N_5904,N_5394);
and U9983 (N_9983,N_7070,N_6578);
nand U9984 (N_9984,N_6205,N_6111);
and U9985 (N_9985,N_6592,N_6194);
or U9986 (N_9986,N_6952,N_5065);
nand U9987 (N_9987,N_6433,N_6083);
nand U9988 (N_9988,N_6578,N_5784);
nand U9989 (N_9989,N_5911,N_5299);
nor U9990 (N_9990,N_5783,N_6197);
nand U9991 (N_9991,N_7064,N_6059);
or U9992 (N_9992,N_7286,N_6484);
or U9993 (N_9993,N_6644,N_6024);
nand U9994 (N_9994,N_6117,N_5728);
and U9995 (N_9995,N_5147,N_5602);
and U9996 (N_9996,N_5748,N_7480);
nand U9997 (N_9997,N_7198,N_5230);
nor U9998 (N_9998,N_6732,N_5725);
nand U9999 (N_9999,N_6275,N_6502);
xnor U10000 (N_10000,N_7857,N_9442);
nand U10001 (N_10001,N_8505,N_9729);
and U10002 (N_10002,N_9225,N_9224);
and U10003 (N_10003,N_7694,N_9458);
and U10004 (N_10004,N_8489,N_9912);
and U10005 (N_10005,N_8777,N_7940);
nand U10006 (N_10006,N_8724,N_8613);
and U10007 (N_10007,N_9069,N_9304);
and U10008 (N_10008,N_8024,N_8929);
or U10009 (N_10009,N_9311,N_9048);
and U10010 (N_10010,N_7731,N_9277);
or U10011 (N_10011,N_8753,N_8962);
nand U10012 (N_10012,N_8490,N_7678);
or U10013 (N_10013,N_8144,N_9668);
or U10014 (N_10014,N_7516,N_8185);
or U10015 (N_10015,N_9743,N_9056);
nand U10016 (N_10016,N_7789,N_9350);
or U10017 (N_10017,N_7621,N_8441);
nor U10018 (N_10018,N_8106,N_9986);
or U10019 (N_10019,N_7910,N_8416);
nand U10020 (N_10020,N_8282,N_9024);
or U10021 (N_10021,N_8181,N_8331);
and U10022 (N_10022,N_9866,N_9779);
xnor U10023 (N_10023,N_7672,N_9349);
nor U10024 (N_10024,N_8367,N_8050);
nand U10025 (N_10025,N_8027,N_9868);
xor U10026 (N_10026,N_8619,N_9127);
nor U10027 (N_10027,N_9393,N_9070);
nand U10028 (N_10028,N_8801,N_9303);
nor U10029 (N_10029,N_7812,N_8726);
nor U10030 (N_10030,N_9239,N_9187);
or U10031 (N_10031,N_9775,N_8544);
and U10032 (N_10032,N_9852,N_8161);
nor U10033 (N_10033,N_8974,N_9008);
and U10034 (N_10034,N_9074,N_8952);
and U10035 (N_10035,N_9190,N_8340);
and U10036 (N_10036,N_9020,N_9039);
nand U10037 (N_10037,N_8557,N_7778);
or U10038 (N_10038,N_8856,N_7598);
nor U10039 (N_10039,N_8029,N_9135);
nor U10040 (N_10040,N_9686,N_7639);
nor U10041 (N_10041,N_9254,N_8214);
xnor U10042 (N_10042,N_8858,N_9313);
and U10043 (N_10043,N_9540,N_9728);
nor U10044 (N_10044,N_9967,N_9267);
or U10045 (N_10045,N_9933,N_9805);
nand U10046 (N_10046,N_7928,N_8848);
xor U10047 (N_10047,N_9772,N_9642);
xor U10048 (N_10048,N_7870,N_8316);
and U10049 (N_10049,N_8804,N_7546);
and U10050 (N_10050,N_9700,N_8793);
nor U10051 (N_10051,N_9291,N_9250);
xor U10052 (N_10052,N_9312,N_7617);
or U10053 (N_10053,N_8243,N_9960);
and U10054 (N_10054,N_9719,N_7770);
xor U10055 (N_10055,N_9103,N_9042);
xor U10056 (N_10056,N_7898,N_7864);
xnor U10057 (N_10057,N_7693,N_8834);
or U10058 (N_10058,N_9257,N_9053);
nand U10059 (N_10059,N_8676,N_7967);
nor U10060 (N_10060,N_9812,N_8813);
and U10061 (N_10061,N_8370,N_9106);
nor U10062 (N_10062,N_9129,N_8889);
nor U10063 (N_10063,N_9154,N_8318);
xor U10064 (N_10064,N_8615,N_8465);
and U10065 (N_10065,N_9867,N_9598);
or U10066 (N_10066,N_9740,N_9915);
or U10067 (N_10067,N_7569,N_9976);
or U10068 (N_10068,N_8796,N_8873);
nor U10069 (N_10069,N_9518,N_7905);
nand U10070 (N_10070,N_7856,N_9230);
or U10071 (N_10071,N_9176,N_8948);
nor U10072 (N_10072,N_7725,N_7763);
xnor U10073 (N_10073,N_9721,N_8495);
xnor U10074 (N_10074,N_8004,N_9076);
xnor U10075 (N_10075,N_9876,N_8506);
or U10076 (N_10076,N_9457,N_8807);
nor U10077 (N_10077,N_9374,N_7842);
xnor U10078 (N_10078,N_9621,N_9751);
or U10079 (N_10079,N_9531,N_8642);
or U10080 (N_10080,N_9270,N_8978);
nor U10081 (N_10081,N_8084,N_9548);
or U10082 (N_10082,N_9123,N_7634);
or U10083 (N_10083,N_9242,N_8934);
nand U10084 (N_10084,N_7850,N_8440);
and U10085 (N_10085,N_8204,N_7846);
or U10086 (N_10086,N_8223,N_8965);
nor U10087 (N_10087,N_9498,N_7821);
nand U10088 (N_10088,N_8055,N_9731);
or U10089 (N_10089,N_7761,N_8943);
nor U10090 (N_10090,N_9208,N_9653);
nand U10091 (N_10091,N_8739,N_8134);
nor U10092 (N_10092,N_8819,N_8314);
and U10093 (N_10093,N_9541,N_8516);
and U10094 (N_10094,N_9379,N_8597);
or U10095 (N_10095,N_7990,N_7767);
xnor U10096 (N_10096,N_8372,N_8482);
or U10097 (N_10097,N_8009,N_7682);
and U10098 (N_10098,N_7995,N_9521);
nor U10099 (N_10099,N_9659,N_9031);
nand U10100 (N_10100,N_9551,N_9762);
nor U10101 (N_10101,N_9606,N_8632);
nor U10102 (N_10102,N_9758,N_9614);
or U10103 (N_10103,N_8829,N_8714);
nor U10104 (N_10104,N_8179,N_9692);
and U10105 (N_10105,N_8066,N_7899);
nand U10106 (N_10106,N_9191,N_8135);
nor U10107 (N_10107,N_8006,N_8885);
nor U10108 (N_10108,N_8337,N_7664);
or U10109 (N_10109,N_9633,N_7513);
nand U10110 (N_10110,N_7628,N_9683);
and U10111 (N_10111,N_9675,N_7648);
or U10112 (N_10112,N_7608,N_8564);
nand U10113 (N_10113,N_7640,N_9603);
nor U10114 (N_10114,N_9016,N_7661);
and U10115 (N_10115,N_9564,N_8045);
nor U10116 (N_10116,N_7970,N_7635);
xnor U10117 (N_10117,N_8594,N_8743);
nor U10118 (N_10118,N_8342,N_7573);
nand U10119 (N_10119,N_9180,N_9770);
nor U10120 (N_10120,N_8507,N_8323);
nor U10121 (N_10121,N_7885,N_8790);
nand U10122 (N_10122,N_8652,N_9273);
or U10123 (N_10123,N_7562,N_9328);
nor U10124 (N_10124,N_8076,N_8221);
nand U10125 (N_10125,N_7599,N_9107);
nand U10126 (N_10126,N_8396,N_8931);
xor U10127 (N_10127,N_8049,N_7755);
nand U10128 (N_10128,N_8643,N_9822);
xor U10129 (N_10129,N_8748,N_8442);
nand U10130 (N_10130,N_8320,N_7706);
nor U10131 (N_10131,N_8246,N_9950);
or U10132 (N_10132,N_8013,N_9892);
or U10133 (N_10133,N_8265,N_9321);
or U10134 (N_10134,N_8138,N_9409);
nand U10135 (N_10135,N_9138,N_8166);
or U10136 (N_10136,N_8114,N_8721);
nand U10137 (N_10137,N_7520,N_8556);
or U10138 (N_10138,N_8252,N_7897);
xnor U10139 (N_10139,N_9214,N_9280);
xnor U10140 (N_10140,N_9294,N_7587);
xor U10141 (N_10141,N_7802,N_9591);
and U10142 (N_10142,N_8865,N_9641);
or U10143 (N_10143,N_9987,N_7583);
or U10144 (N_10144,N_8887,N_9813);
and U10145 (N_10145,N_9702,N_9501);
nor U10146 (N_10146,N_8783,N_9279);
nand U10147 (N_10147,N_9783,N_9796);
or U10148 (N_10148,N_9872,N_8281);
and U10149 (N_10149,N_8317,N_9162);
and U10150 (N_10150,N_7539,N_8893);
and U10151 (N_10151,N_7961,N_8696);
nand U10152 (N_10152,N_7966,N_9099);
nand U10153 (N_10153,N_7948,N_8451);
nand U10154 (N_10154,N_9786,N_8357);
nand U10155 (N_10155,N_7515,N_7859);
or U10156 (N_10156,N_8010,N_8620);
nand U10157 (N_10157,N_8860,N_9677);
or U10158 (N_10158,N_9245,N_8047);
nor U10159 (N_10159,N_8108,N_7774);
or U10160 (N_10160,N_8382,N_9488);
nor U10161 (N_10161,N_9382,N_8303);
nor U10162 (N_10162,N_9814,N_9716);
nand U10163 (N_10163,N_8043,N_7919);
nand U10164 (N_10164,N_7510,N_8837);
and U10165 (N_10165,N_8062,N_9661);
nand U10166 (N_10166,N_9730,N_8278);
and U10167 (N_10167,N_8231,N_7909);
or U10168 (N_10168,N_8659,N_8525);
nand U10169 (N_10169,N_7975,N_7819);
nand U10170 (N_10170,N_9090,N_7519);
xnor U10171 (N_10171,N_8614,N_8876);
nor U10172 (N_10172,N_9901,N_9063);
or U10173 (N_10173,N_8773,N_8930);
nor U10174 (N_10174,N_9632,N_7645);
or U10175 (N_10175,N_9860,N_9412);
or U10176 (N_10176,N_8852,N_9497);
nor U10177 (N_10177,N_9147,N_9777);
and U10178 (N_10178,N_9274,N_8309);
and U10179 (N_10179,N_9195,N_9478);
nand U10180 (N_10180,N_8638,N_8792);
xor U10181 (N_10181,N_8483,N_8651);
or U10182 (N_10182,N_8000,N_8609);
nor U10183 (N_10183,N_8971,N_8037);
and U10184 (N_10184,N_9506,N_9526);
nor U10185 (N_10185,N_8170,N_9694);
nand U10186 (N_10186,N_9645,N_8582);
xor U10187 (N_10187,N_9970,N_7564);
and U10188 (N_10188,N_9470,N_8348);
nand U10189 (N_10189,N_7791,N_9262);
xnor U10190 (N_10190,N_9894,N_9984);
nor U10191 (N_10191,N_8032,N_8537);
nor U10192 (N_10192,N_9196,N_7551);
and U10193 (N_10193,N_8110,N_9482);
xor U10194 (N_10194,N_7709,N_8545);
and U10195 (N_10195,N_7922,N_8275);
nor U10196 (N_10196,N_8722,N_9619);
nand U10197 (N_10197,N_8436,N_8497);
nand U10198 (N_10198,N_9268,N_8761);
or U10199 (N_10199,N_7824,N_8859);
and U10200 (N_10200,N_8477,N_7743);
and U10201 (N_10201,N_7676,N_9825);
nor U10202 (N_10202,N_9080,N_9906);
nand U10203 (N_10203,N_8184,N_9649);
and U10204 (N_10204,N_8104,N_9736);
nand U10205 (N_10205,N_8890,N_9887);
or U10206 (N_10206,N_8881,N_7983);
nor U10207 (N_10207,N_9465,N_9781);
xor U10208 (N_10208,N_9459,N_9152);
or U10209 (N_10209,N_8028,N_7855);
xnor U10210 (N_10210,N_8260,N_8174);
or U10211 (N_10211,N_9395,N_8989);
or U10212 (N_10212,N_7652,N_8069);
or U10213 (N_10213,N_9856,N_9726);
nor U10214 (N_10214,N_9308,N_9732);
or U10215 (N_10215,N_8680,N_9168);
or U10216 (N_10216,N_7772,N_9553);
nand U10217 (N_10217,N_9701,N_9373);
nor U10218 (N_10218,N_7886,N_8664);
nand U10219 (N_10219,N_8142,N_9820);
xor U10220 (N_10220,N_8175,N_8498);
or U10221 (N_10221,N_8822,N_8227);
xnor U10222 (N_10222,N_8752,N_8727);
nor U10223 (N_10223,N_7536,N_9452);
xnor U10224 (N_10224,N_9390,N_8571);
xor U10225 (N_10225,N_8261,N_8186);
xnor U10226 (N_10226,N_9408,N_8584);
nor U10227 (N_10227,N_9169,N_9693);
or U10228 (N_10228,N_7826,N_8581);
xnor U10229 (N_10229,N_8888,N_8390);
xnor U10230 (N_10230,N_8800,N_8328);
or U10231 (N_10231,N_9480,N_7861);
nor U10232 (N_10232,N_8397,N_9445);
nand U10233 (N_10233,N_9744,N_9605);
nor U10234 (N_10234,N_9791,N_9681);
or U10235 (N_10235,N_7747,N_9865);
nor U10236 (N_10236,N_9845,N_8353);
or U10237 (N_10237,N_9184,N_9626);
nand U10238 (N_10238,N_8673,N_9010);
nand U10239 (N_10239,N_8250,N_9334);
nor U10240 (N_10240,N_9699,N_9229);
xnor U10241 (N_10241,N_9928,N_8710);
or U10242 (N_10242,N_8526,N_7646);
or U10243 (N_10243,N_7688,N_7765);
nor U10244 (N_10244,N_8457,N_7777);
or U10245 (N_10245,N_9908,N_8253);
nor U10246 (N_10246,N_9492,N_8349);
or U10247 (N_10247,N_7528,N_8277);
and U10248 (N_10248,N_9787,N_9114);
and U10249 (N_10249,N_8120,N_7538);
nor U10250 (N_10250,N_8668,N_8511);
xnor U10251 (N_10251,N_9949,N_8669);
and U10252 (N_10252,N_8162,N_7914);
or U10253 (N_10253,N_8606,N_8139);
nor U10254 (N_10254,N_9994,N_7845);
and U10255 (N_10255,N_9003,N_8901);
and U10256 (N_10256,N_9368,N_8406);
and U10257 (N_10257,N_9634,N_8681);
and U10258 (N_10258,N_8666,N_9358);
xnor U10259 (N_10259,N_9504,N_9171);
or U10260 (N_10260,N_8476,N_7653);
nor U10261 (N_10261,N_9620,N_8137);
nor U10262 (N_10262,N_9910,N_8258);
or U10263 (N_10263,N_8313,N_8570);
nor U10264 (N_10264,N_7533,N_8052);
or U10265 (N_10265,N_8445,N_8289);
nor U10266 (N_10266,N_8682,N_7982);
nor U10267 (N_10267,N_8823,N_9767);
nor U10268 (N_10268,N_9835,N_7744);
nor U10269 (N_10269,N_7759,N_9499);
or U10270 (N_10270,N_7997,N_9363);
nor U10271 (N_10271,N_9182,N_7602);
or U10272 (N_10272,N_9516,N_9883);
nor U10273 (N_10273,N_9370,N_9101);
nor U10274 (N_10274,N_9647,N_8663);
nor U10275 (N_10275,N_9665,N_8623);
or U10276 (N_10276,N_8454,N_9296);
xnor U10277 (N_10277,N_9007,N_8096);
and U10278 (N_10278,N_9017,N_9420);
nand U10279 (N_10279,N_8361,N_8466);
or U10280 (N_10280,N_7851,N_9596);
nand U10281 (N_10281,N_9177,N_8167);
and U10282 (N_10282,N_8533,N_8008);
nand U10283 (N_10283,N_9679,N_7702);
nor U10284 (N_10284,N_9018,N_8379);
nand U10285 (N_10285,N_7888,N_9573);
nor U10286 (N_10286,N_8405,N_9916);
nand U10287 (N_10287,N_8503,N_9194);
nor U10288 (N_10288,N_7553,N_9561);
or U10289 (N_10289,N_9232,N_8604);
and U10290 (N_10290,N_8884,N_8662);
nand U10291 (N_10291,N_8399,N_8216);
nand U10292 (N_10292,N_9778,N_8569);
or U10293 (N_10293,N_9151,N_8065);
nand U10294 (N_10294,N_8307,N_8305);
nand U10295 (N_10295,N_8156,N_9961);
nor U10296 (N_10296,N_9174,N_9853);
or U10297 (N_10297,N_9980,N_8732);
nor U10298 (N_10298,N_7929,N_9060);
nor U10299 (N_10299,N_9489,N_8070);
nor U10300 (N_10300,N_9510,N_8195);
and U10301 (N_10301,N_7558,N_9329);
xor U10302 (N_10302,N_8863,N_7580);
or U10303 (N_10303,N_9167,N_8061);
or U10304 (N_10304,N_8844,N_9335);
nand U10305 (N_10305,N_7853,N_7756);
or U10306 (N_10306,N_7656,N_9354);
nor U10307 (N_10307,N_7798,N_9907);
and U10308 (N_10308,N_9983,N_9713);
or U10309 (N_10309,N_8904,N_9185);
or U10310 (N_10310,N_7732,N_9446);
nor U10311 (N_10311,N_9166,N_9502);
or U10312 (N_10312,N_9939,N_7739);
xnor U10313 (N_10313,N_9071,N_9417);
or U10314 (N_10314,N_8658,N_9663);
or U10315 (N_10315,N_7511,N_8315);
nor U10316 (N_10316,N_8842,N_9473);
xnor U10317 (N_10317,N_7891,N_9365);
nand U10318 (N_10318,N_8546,N_9571);
nor U10319 (N_10319,N_7996,N_7878);
nand U10320 (N_10320,N_8444,N_7633);
and U10321 (N_10321,N_8363,N_7769);
and U10322 (N_10322,N_7504,N_9923);
or U10323 (N_10323,N_8407,N_7508);
nand U10324 (N_10324,N_9846,N_7659);
nor U10325 (N_10325,N_9925,N_8508);
nor U10326 (N_10326,N_8140,N_8979);
nor U10327 (N_10327,N_7957,N_8499);
nand U10328 (N_10328,N_9087,N_8479);
and U10329 (N_10329,N_7805,N_8287);
nor U10330 (N_10330,N_9742,N_9249);
nand U10331 (N_10331,N_9757,N_9124);
nor U10332 (N_10332,N_9266,N_7545);
nor U10333 (N_10333,N_7920,N_8913);
or U10334 (N_10334,N_8383,N_8095);
nand U10335 (N_10335,N_7781,N_8079);
or U10336 (N_10336,N_8755,N_8625);
nor U10337 (N_10337,N_8791,N_8836);
nand U10338 (N_10338,N_8808,N_8786);
xor U10339 (N_10339,N_7614,N_8951);
nor U10340 (N_10340,N_8500,N_8891);
or U10341 (N_10341,N_9589,N_9829);
and U10342 (N_10342,N_9133,N_9075);
nor U10343 (N_10343,N_8646,N_8236);
xor U10344 (N_10344,N_9464,N_8933);
xnor U10345 (N_10345,N_7740,N_8412);
nand U10346 (N_10346,N_7958,N_8271);
or U10347 (N_10347,N_9372,N_7729);
and U10348 (N_10348,N_8016,N_7749);
and U10349 (N_10349,N_7822,N_9049);
or U10350 (N_10350,N_8909,N_8158);
nand U10351 (N_10351,N_9914,N_9119);
and U10352 (N_10352,N_9064,N_9323);
nand U10353 (N_10353,N_9749,N_8715);
nor U10354 (N_10354,N_9886,N_9735);
nor U10355 (N_10355,N_8064,N_7655);
nand U10356 (N_10356,N_7594,N_7629);
or U10357 (N_10357,N_9431,N_8088);
nor U10358 (N_10358,N_9330,N_7716);
and U10359 (N_10359,N_8459,N_8924);
or U10360 (N_10360,N_7815,N_9227);
or U10361 (N_10361,N_9574,N_9893);
and U10362 (N_10362,N_8515,N_8333);
nand U10363 (N_10363,N_8048,N_7788);
nand U10364 (N_10364,N_8919,N_8912);
and U10365 (N_10365,N_9352,N_8756);
nor U10366 (N_10366,N_7529,N_8254);
nand U10367 (N_10367,N_8322,N_9202);
or U10368 (N_10368,N_7623,N_9585);
nand U10369 (N_10369,N_7620,N_7609);
nand U10370 (N_10370,N_8918,N_7890);
and U10371 (N_10371,N_9198,N_8846);
or U10372 (N_10372,N_8017,N_7872);
and U10373 (N_10373,N_8558,N_9996);
nor U10374 (N_10374,N_9423,N_9025);
nand U10375 (N_10375,N_7792,N_9284);
or U10376 (N_10376,N_8746,N_7913);
or U10377 (N_10377,N_8311,N_9121);
nor U10378 (N_10378,N_8081,N_9715);
or U10379 (N_10379,N_8877,N_9947);
and U10380 (N_10380,N_9292,N_8598);
nor U10381 (N_10381,N_9973,N_9377);
and U10382 (N_10382,N_9479,N_7968);
xor U10383 (N_10383,N_8700,N_9319);
nand U10384 (N_10384,N_9258,N_7657);
or U10385 (N_10385,N_7951,N_9369);
and U10386 (N_10386,N_8365,N_8798);
nor U10387 (N_10387,N_8220,N_9929);
or U10388 (N_10388,N_9922,N_9112);
or U10389 (N_10389,N_9529,N_8723);
nand U10390 (N_10390,N_9555,N_9275);
or U10391 (N_10391,N_8734,N_9919);
nand U10392 (N_10392,N_8622,N_9801);
and U10393 (N_10393,N_8704,N_7708);
nand U10394 (N_10394,N_8180,N_7862);
nand U10395 (N_10395,N_7523,N_8431);
and U10396 (N_10396,N_8075,N_7719);
or U10397 (N_10397,N_9221,N_9722);
and U10398 (N_10398,N_9942,N_7847);
and U10399 (N_10399,N_9386,N_9233);
and U10400 (N_10400,N_7939,N_8400);
xor U10401 (N_10401,N_7795,N_9997);
nor U10402 (N_10402,N_8915,N_7581);
nand U10403 (N_10403,N_8122,N_7838);
nor U10404 (N_10404,N_8802,N_8554);
xor U10405 (N_10405,N_7935,N_8855);
nor U10406 (N_10406,N_8218,N_7760);
and U10407 (N_10407,N_8882,N_8749);
or U10408 (N_10408,N_8085,N_8470);
or U10409 (N_10409,N_9451,N_9885);
or U10410 (N_10410,N_8942,N_8932);
nand U10411 (N_10411,N_9944,N_7860);
nand U10412 (N_10412,N_8414,N_8892);
and U10413 (N_10413,N_8063,N_7977);
and U10414 (N_10414,N_9857,N_8121);
or U10415 (N_10415,N_7949,N_8713);
xnor U10416 (N_10416,N_9660,N_9727);
or U10417 (N_10417,N_8742,N_9367);
xnor U10418 (N_10418,N_9341,N_8820);
nand U10419 (N_10419,N_9082,N_8034);
or U10420 (N_10420,N_9560,N_9200);
nor U10421 (N_10421,N_8921,N_8423);
and U10422 (N_10422,N_8267,N_8538);
or U10423 (N_10423,N_8857,N_8398);
xor U10424 (N_10424,N_8949,N_9037);
or U10425 (N_10425,N_9612,N_9132);
xor U10426 (N_10426,N_8778,N_8373);
nand U10427 (N_10427,N_8982,N_9988);
xor U10428 (N_10428,N_9131,N_9259);
nor U10429 (N_10429,N_8384,N_8968);
nor U10430 (N_10430,N_8381,N_9635);
nand U10431 (N_10431,N_9828,N_8270);
and U10432 (N_10432,N_8939,N_8201);
or U10433 (N_10433,N_7662,N_8716);
nand U10434 (N_10434,N_9746,N_8452);
or U10435 (N_10435,N_9794,N_8428);
or U10436 (N_10436,N_8975,N_9029);
and U10437 (N_10437,N_7517,N_8559);
or U10438 (N_10438,N_7556,N_9183);
nand U10439 (N_10439,N_8014,N_8364);
nor U10440 (N_10440,N_9240,N_7803);
xor U10441 (N_10441,N_9342,N_7809);
nor U10442 (N_10442,N_9302,N_7559);
nand U10443 (N_10443,N_7810,N_8954);
and U10444 (N_10444,N_8839,N_9260);
and U10445 (N_10445,N_8649,N_8657);
nor U10446 (N_10446,N_8502,N_7624);
or U10447 (N_10447,N_7547,N_8895);
nand U10448 (N_10448,N_9505,N_9955);
or U10449 (N_10449,N_9093,N_9116);
nand U10450 (N_10450,N_8393,N_9343);
or U10451 (N_10451,N_9345,N_8925);
nand U10452 (N_10452,N_9231,N_8344);
nor U10453 (N_10453,N_9036,N_8988);
and U10454 (N_10454,N_7535,N_9766);
and U10455 (N_10455,N_9572,N_7673);
nand U10456 (N_10456,N_7566,N_9785);
nor U10457 (N_10457,N_9696,N_9637);
or U10458 (N_10458,N_7830,N_8439);
nand U10459 (N_10459,N_9397,N_8816);
nand U10460 (N_10460,N_8072,N_8443);
and U10461 (N_10461,N_7554,N_8731);
nor U10462 (N_10462,N_8774,N_9780);
or U10463 (N_10463,N_8450,N_7690);
and U10464 (N_10464,N_8686,N_8080);
nand U10465 (N_10465,N_7991,N_8878);
or U10466 (N_10466,N_7783,N_9690);
or U10467 (N_10467,N_9963,N_7695);
nand U10468 (N_10468,N_9760,N_9269);
nand U10469 (N_10469,N_9437,N_8102);
and U10470 (N_10470,N_8553,N_9979);
and U10471 (N_10471,N_8678,N_8529);
xor U10472 (N_10472,N_9128,N_7685);
nand U10473 (N_10473,N_9869,N_9088);
or U10474 (N_10474,N_7900,N_9543);
nand U10475 (N_10475,N_8868,N_9160);
or U10476 (N_10476,N_8645,N_7960);
or U10477 (N_10477,N_9290,N_8896);
and U10478 (N_10478,N_9041,N_9765);
nor U10479 (N_10479,N_8226,N_9554);
nor U10480 (N_10480,N_9113,N_9559);
or U10481 (N_10481,N_7563,N_9440);
nand U10482 (N_10482,N_7895,N_9278);
or U10483 (N_10483,N_9537,N_8324);
or U10484 (N_10484,N_8205,N_7689);
or U10485 (N_10485,N_8264,N_9595);
nor U10486 (N_10486,N_9153,N_7941);
or U10487 (N_10487,N_7712,N_9858);
and U10488 (N_10488,N_7540,N_8765);
nor U10489 (N_10489,N_8321,N_8733);
or U10490 (N_10490,N_8005,N_9376);
nor U10491 (N_10491,N_8561,N_7978);
and U10492 (N_10492,N_8435,N_8972);
nand U10493 (N_10493,N_9579,N_7683);
or U10494 (N_10494,N_8200,N_7684);
nand U10495 (N_10495,N_8665,N_7985);
nor U10496 (N_10496,N_8094,N_8699);
nor U10497 (N_10497,N_9079,N_8605);
and U10498 (N_10498,N_9490,N_9806);
nand U10499 (N_10499,N_8990,N_9424);
nor U10500 (N_10500,N_9340,N_8776);
xor U10501 (N_10501,N_8136,N_9375);
nand U10502 (N_10502,N_8985,N_9466);
and U10503 (N_10503,N_7619,N_7671);
and U10504 (N_10504,N_9889,N_9021);
nand U10505 (N_10505,N_7813,N_9827);
or U10506 (N_10506,N_9247,N_8639);
nor U10507 (N_10507,N_9447,N_9832);
nor U10508 (N_10508,N_8667,N_9618);
and U10509 (N_10509,N_9314,N_9285);
nor U10510 (N_10510,N_7544,N_9899);
nor U10511 (N_10511,N_7721,N_7931);
nand U10512 (N_10512,N_8789,N_9484);
or U10513 (N_10513,N_8377,N_8833);
and U10514 (N_10514,N_7615,N_7816);
or U10515 (N_10515,N_8832,N_8284);
or U10516 (N_10516,N_9419,N_8617);
and U10517 (N_10517,N_8573,N_8164);
xnor U10518 (N_10518,N_8484,N_8946);
and U10519 (N_10519,N_8283,N_7787);
nor U10520 (N_10520,N_9590,N_8199);
or U10521 (N_10521,N_8251,N_8125);
or U10522 (N_10522,N_8212,N_9616);
and U10523 (N_10523,N_8916,N_7576);
nor U10524 (N_10524,N_9804,N_9186);
nor U10525 (N_10525,N_9246,N_9847);
nand U10526 (N_10526,N_8828,N_8105);
and U10527 (N_10527,N_7514,N_7925);
or U10528 (N_10528,N_7527,N_7954);
and U10529 (N_10529,N_8660,N_8935);
or U10530 (N_10530,N_8944,N_8419);
or U10531 (N_10531,N_9680,N_9125);
nand U10532 (N_10532,N_7613,N_8927);
nor U10533 (N_10533,N_8769,N_8923);
nor U10534 (N_10534,N_8228,N_9092);
nand U10535 (N_10535,N_9158,N_7503);
nor U10536 (N_10536,N_9644,N_7668);
nand U10537 (N_10537,N_8127,N_9159);
nand U10538 (N_10538,N_9669,N_8585);
or U10539 (N_10539,N_8718,N_7699);
and U10540 (N_10540,N_9584,N_9034);
nand U10541 (N_10541,N_8961,N_8831);
nand U10542 (N_10542,N_7943,N_8685);
nand U10543 (N_10543,N_9809,N_9831);
nor U10544 (N_10544,N_8413,N_7532);
or U10545 (N_10545,N_8474,N_8825);
nand U10546 (N_10546,N_9689,N_8523);
nand U10547 (N_10547,N_9648,N_9207);
nor U10548 (N_10548,N_7593,N_9172);
xnor U10549 (N_10549,N_9546,N_7686);
nor U10550 (N_10550,N_7717,N_8171);
or U10551 (N_10551,N_9297,N_8647);
or U10552 (N_10552,N_7701,N_8446);
xnor U10553 (N_10553,N_8119,N_9754);
and U10554 (N_10554,N_9491,N_7750);
or U10555 (N_10555,N_8957,N_8712);
and U10556 (N_10556,N_7549,N_9384);
or U10557 (N_10557,N_9611,N_9461);
nand U10558 (N_10558,N_7567,N_9309);
nand U10559 (N_10559,N_9674,N_9938);
nor U10560 (N_10560,N_8815,N_7703);
or U10561 (N_10561,N_7666,N_7754);
or U10562 (N_10562,N_7560,N_7938);
and U10563 (N_10563,N_9098,N_9035);
xnor U10564 (N_10564,N_8562,N_9052);
nand U10565 (N_10565,N_9199,N_7800);
and U10566 (N_10566,N_9897,N_9219);
nor U10567 (N_10567,N_9438,N_8151);
and U10568 (N_10568,N_8803,N_8725);
or U10569 (N_10569,N_9462,N_8698);
and U10570 (N_10570,N_8580,N_7650);
and U10571 (N_10571,N_7811,N_9870);
nor U10572 (N_10572,N_9205,N_9061);
xor U10573 (N_10573,N_8350,N_8964);
nand U10574 (N_10574,N_8346,N_8187);
and U10575 (N_10575,N_8402,N_8422);
nand U10576 (N_10576,N_7521,N_8023);
nor U10577 (N_10577,N_8233,N_8330);
nand U10578 (N_10578,N_9348,N_8310);
nand U10579 (N_10579,N_8551,N_9667);
or U10580 (N_10580,N_9398,N_8327);
nor U10581 (N_10581,N_8123,N_9065);
nor U10582 (N_10582,N_8298,N_9047);
or U10583 (N_10583,N_7727,N_8654);
nand U10584 (N_10584,N_8702,N_8552);
or U10585 (N_10585,N_9477,N_8602);
nor U10586 (N_10586,N_8782,N_9094);
nand U10587 (N_10587,N_9263,N_9353);
nor U10588 (N_10588,N_8449,N_9433);
nor U10589 (N_10589,N_8154,N_8438);
xor U10590 (N_10590,N_7921,N_8492);
nand U10591 (N_10591,N_8073,N_7715);
or U10592 (N_10592,N_8631,N_8897);
nand U10593 (N_10593,N_8098,N_8955);
and U10594 (N_10594,N_7987,N_8621);
and U10595 (N_10595,N_8589,N_8341);
nor U10596 (N_10596,N_7762,N_9797);
nand U10597 (N_10597,N_7570,N_8059);
nor U10598 (N_10598,N_8130,N_9613);
and U10599 (N_10599,N_8514,N_8359);
and U10600 (N_10600,N_7937,N_7873);
nand U10601 (N_10601,N_9811,N_9926);
or U10602 (N_10602,N_7992,N_9600);
xnor U10603 (N_10603,N_9295,N_8705);
nand U10604 (N_10604,N_9905,N_8297);
nor U10605 (N_10605,N_9911,N_7757);
nand U10606 (N_10606,N_8586,N_9389);
and U10607 (N_10607,N_8291,N_9753);
nor U10608 (N_10608,N_9117,N_9496);
nor U10609 (N_10609,N_7705,N_7625);
nor U10610 (N_10610,N_7828,N_8376);
and U10611 (N_10611,N_8003,N_8784);
nand U10612 (N_10612,N_8155,N_9575);
or U10613 (N_10613,N_9577,N_8177);
or U10614 (N_10614,N_7976,N_9509);
nor U10615 (N_10615,N_8209,N_8242);
nand U10616 (N_10616,N_8480,N_8021);
nor U10617 (N_10617,N_9104,N_9666);
nor U10618 (N_10618,N_7723,N_8071);
nor U10619 (N_10619,N_9238,N_8213);
nand U10620 (N_10620,N_9444,N_8688);
nand U10621 (N_10621,N_9366,N_8494);
nor U10622 (N_10622,N_7865,N_9519);
nor U10623 (N_10623,N_7577,N_9823);
xor U10624 (N_10624,N_7820,N_8118);
nor U10625 (N_10625,N_7808,N_8630);
nand U10626 (N_10626,N_9854,N_7748);
or U10627 (N_10627,N_9102,N_7785);
and U10628 (N_10628,N_8244,N_9532);
or U10629 (N_10629,N_7790,N_9627);
nand U10630 (N_10630,N_9821,N_7651);
or U10631 (N_10631,N_7934,N_8695);
nand U10632 (N_10632,N_9027,N_7746);
and U10633 (N_10633,N_9038,N_7726);
nand U10634 (N_10634,N_8936,N_9536);
and U10635 (N_10635,N_9415,N_7933);
or U10636 (N_10636,N_9977,N_7530);
nand U10637 (N_10637,N_9028,N_8997);
xor U10638 (N_10638,N_8078,N_9073);
and U10639 (N_10639,N_8741,N_9256);
and U10640 (N_10640,N_9771,N_9316);
and U10641 (N_10641,N_9752,N_9305);
and U10642 (N_10642,N_8408,N_7780);
nor U10643 (N_10643,N_9265,N_7641);
and U10644 (N_10644,N_9058,N_7814);
or U10645 (N_10645,N_9046,N_8684);
xor U10646 (N_10646,N_8111,N_9793);
nor U10647 (N_10647,N_9015,N_8115);
or U10648 (N_10648,N_8757,N_8953);
or U10649 (N_10649,N_8871,N_8217);
or U10650 (N_10650,N_9629,N_9120);
nor U10651 (N_10651,N_9547,N_7882);
xnor U10652 (N_10652,N_9628,N_9512);
or U10653 (N_10653,N_9400,N_7879);
nor U10654 (N_10654,N_8109,N_8387);
or U10655 (N_10655,N_9631,N_9346);
and U10656 (N_10656,N_7713,N_8239);
nand U10657 (N_10657,N_8430,N_8566);
nor U10658 (N_10658,N_8293,N_9687);
and U10659 (N_10659,N_7561,N_9909);
and U10660 (N_10660,N_9898,N_9001);
and U10661 (N_10661,N_8172,N_7710);
and U10662 (N_10662,N_9759,N_9819);
and U10663 (N_10663,N_9784,N_9456);
nand U10664 (N_10664,N_7591,N_8650);
nand U10665 (N_10665,N_9664,N_7603);
or U10666 (N_10666,N_9432,N_7947);
and U10667 (N_10667,N_7840,N_8814);
nand U10668 (N_10668,N_8485,N_8276);
xnor U10669 (N_10669,N_9951,N_8535);
or U10670 (N_10670,N_9359,N_8165);
and U10671 (N_10671,N_8543,N_9149);
or U10672 (N_10672,N_7852,N_8051);
or U10673 (N_10673,N_8304,N_7506);
xor U10674 (N_10674,N_9646,N_9426);
or U10675 (N_10675,N_7955,N_8129);
and U10676 (N_10676,N_9552,N_8610);
or U10677 (N_10677,N_9900,N_7832);
nand U10678 (N_10678,N_9818,N_8811);
nand U10679 (N_10679,N_8577,N_8089);
or U10680 (N_10680,N_9109,N_8854);
and U10681 (N_10681,N_8707,N_9576);
and U10682 (N_10682,N_8527,N_8751);
nand U10683 (N_10683,N_9213,N_8160);
and U10684 (N_10684,N_9173,N_8977);
or U10685 (N_10685,N_7730,N_8588);
nand U10686 (N_10686,N_9210,N_8203);
xnor U10687 (N_10687,N_9067,N_9720);
or U10688 (N_10688,N_8116,N_9429);
and U10689 (N_10689,N_8574,N_9043);
nand U10690 (N_10690,N_9150,N_7945);
and U10691 (N_10691,N_9272,N_9126);
and U10692 (N_10692,N_9836,N_8295);
or U10693 (N_10693,N_9493,N_8020);
nand U10694 (N_10694,N_7946,N_8240);
and U10695 (N_10695,N_9685,N_8022);
or U10696 (N_10696,N_8730,N_7902);
and U10697 (N_10697,N_9795,N_9896);
and U10698 (N_10698,N_9118,N_7758);
nor U10699 (N_10699,N_8640,N_9843);
or U10700 (N_10700,N_8074,N_7574);
nand U10701 (N_10701,N_9873,N_9019);
or U10702 (N_10702,N_8259,N_9243);
or U10703 (N_10703,N_8339,N_8425);
xnor U10704 (N_10704,N_7989,N_8809);
nor U10705 (N_10705,N_8945,N_8332);
or U10706 (N_10706,N_8183,N_9741);
nand U10707 (N_10707,N_8437,N_9441);
or U10708 (N_10708,N_9755,N_9850);
or U10709 (N_10709,N_9223,N_8867);
or U10710 (N_10710,N_8607,N_9724);
and U10711 (N_10711,N_7518,N_9235);
nand U10712 (N_10712,N_9189,N_9972);
xnor U10713 (N_10713,N_9990,N_8101);
nor U10714 (N_10714,N_9212,N_7680);
and U10715 (N_10715,N_8159,N_8455);
or U10716 (N_10716,N_8572,N_8128);
and U10717 (N_10717,N_7722,N_7881);
and U10718 (N_10718,N_8099,N_8448);
or U10719 (N_10719,N_9817,N_9022);
or U10720 (N_10720,N_7793,N_9436);
nor U10721 (N_10721,N_9884,N_8417);
or U10722 (N_10722,N_9032,N_8041);
and U10723 (N_10723,N_7696,N_7799);
nand U10724 (N_10724,N_9276,N_9298);
and U10725 (N_10725,N_8025,N_9364);
nor U10726 (N_10726,N_7796,N_9826);
and U10727 (N_10727,N_9640,N_7665);
or U10728 (N_10728,N_8720,N_7541);
nand U10729 (N_10729,N_9371,N_8157);
and U10730 (N_10730,N_8542,N_7883);
or U10731 (N_10731,N_8736,N_9077);
nand U10732 (N_10732,N_9450,N_9953);
or U10733 (N_10733,N_9201,N_9824);
nand U10734 (N_10734,N_9578,N_9084);
nand U10735 (N_10735,N_9958,N_9192);
xor U10736 (N_10736,N_7707,N_9544);
nor U10737 (N_10737,N_8996,N_8595);
xor U10738 (N_10738,N_8903,N_9218);
nand U10739 (N_10739,N_9882,N_8509);
nor U10740 (N_10740,N_9081,N_9322);
or U10741 (N_10741,N_9705,N_9924);
or U10742 (N_10742,N_7507,N_8056);
nor U10743 (N_10743,N_8152,N_8993);
nor U10744 (N_10744,N_7588,N_8843);
xnor U10745 (N_10745,N_9315,N_9562);
xnor U10746 (N_10746,N_8827,N_8475);
or U10747 (N_10747,N_9320,N_9964);
nand U10748 (N_10748,N_7752,N_9557);
or U10749 (N_10749,N_8775,N_9293);
and U10750 (N_10750,N_8468,N_9834);
and U10751 (N_10751,N_8229,N_7917);
and U10752 (N_10752,N_8378,N_7737);
nand U10753 (N_10753,N_8133,N_9237);
and U10754 (N_10754,N_9567,N_7637);
or U10755 (N_10755,N_8879,N_7971);
nand U10756 (N_10756,N_8970,N_7950);
nand U10757 (N_10757,N_7930,N_7901);
xnor U10758 (N_10758,N_8464,N_9799);
or U10759 (N_10759,N_7892,N_9652);
or U10760 (N_10760,N_8266,N_9156);
and U10761 (N_10761,N_8692,N_8401);
and U10762 (N_10762,N_8987,N_9638);
xnor U10763 (N_10763,N_9130,N_7936);
or U10764 (N_10764,N_9839,N_8268);
and U10765 (N_10765,N_9952,N_9416);
and U10766 (N_10766,N_7848,N_7512);
or U10767 (N_10767,N_9255,N_9830);
xnor U10768 (N_10768,N_8433,N_7896);
or U10769 (N_10769,N_7611,N_8866);
nand U10770 (N_10770,N_7876,N_7578);
nand U10771 (N_10771,N_9968,N_9682);
or U10772 (N_10772,N_8463,N_8883);
and U10773 (N_10773,N_9959,N_7691);
or U10774 (N_10774,N_9105,N_7817);
nor U10775 (N_10775,N_8611,N_8237);
nor U10776 (N_10776,N_9197,N_9930);
and U10777 (N_10777,N_9657,N_9511);
nand U10778 (N_10778,N_9601,N_7736);
or U10779 (N_10779,N_8030,N_7984);
xor U10780 (N_10780,N_8222,N_7550);
nand U10781 (N_10781,N_8616,N_8241);
and U10782 (N_10782,N_8198,N_8628);
nand U10783 (N_10783,N_8176,N_8596);
nor U10784 (N_10784,N_8518,N_8629);
nor U10785 (N_10785,N_8806,N_8694);
and U10786 (N_10786,N_8835,N_8576);
or U10787 (N_10787,N_7972,N_9507);
or U10788 (N_10788,N_8764,N_7866);
nor U10789 (N_10789,N_8750,N_9453);
or U10790 (N_10790,N_8103,N_9002);
nand U10791 (N_10791,N_9999,N_8656);
nand U10792 (N_10792,N_9401,N_9588);
and U10793 (N_10793,N_9337,N_9467);
nand U10794 (N_10794,N_8821,N_9317);
nand U10795 (N_10795,N_8547,N_9688);
xor U10796 (N_10796,N_9803,N_9671);
and U10797 (N_10797,N_8481,N_8215);
and U10798 (N_10798,N_8169,N_9747);
nor U10799 (N_10799,N_9097,N_9425);
xnor U10800 (N_10800,N_9085,N_9599);
or U10801 (N_10801,N_9975,N_9066);
nand U10802 (N_10802,N_9508,N_9528);
xor U10803 (N_10803,N_9932,N_7887);
and U10804 (N_10804,N_9844,N_9054);
nor U10805 (N_10805,N_8513,N_8235);
nor U10806 (N_10806,N_7753,N_9739);
or U10807 (N_10807,N_8097,N_8335);
nor U10808 (N_10808,N_9837,N_8190);
nor U10809 (N_10809,N_8817,N_8469);
nor U10810 (N_10810,N_9717,N_7916);
nor U10811 (N_10811,N_9863,N_9734);
nand U10812 (N_10812,N_8354,N_9157);
nand U10813 (N_10813,N_8626,N_9142);
xor U10814 (N_10814,N_8148,N_7642);
nor U10815 (N_10815,N_9422,N_8633);
nor U10816 (N_10816,N_8937,N_9656);
nor U10817 (N_10817,N_9602,N_9802);
xnor U10818 (N_10818,N_7907,N_8356);
nand U10819 (N_10819,N_7903,N_8427);
or U10820 (N_10820,N_8870,N_7973);
and U10821 (N_10821,N_9523,N_9222);
nor U10822 (N_10822,N_8288,N_9072);
and U10823 (N_10823,N_9875,N_8969);
nor U10824 (N_10824,N_9188,N_9798);
nand U10825 (N_10825,N_9630,N_8910);
nand U10826 (N_10826,N_7831,N_8539);
nand U10827 (N_10827,N_7596,N_8693);
nand U10828 (N_10828,N_8083,N_7745);
nor U10829 (N_10829,N_7616,N_7959);
nor U10830 (N_10830,N_8279,N_9851);
nor U10831 (N_10831,N_8426,N_7597);
or U10832 (N_10832,N_9495,N_8093);
or U10833 (N_10833,N_7626,N_9816);
nor U10834 (N_10834,N_7786,N_8966);
nand U10835 (N_10835,N_7500,N_9655);
and U10836 (N_10836,N_9193,N_8269);
nand U10837 (N_10837,N_7911,N_9111);
nor U10838 (N_10838,N_9710,N_8635);
nor U10839 (N_10839,N_8703,N_9244);
nor U10840 (N_10840,N_8182,N_9206);
and U10841 (N_10841,N_9472,N_8090);
xor U10842 (N_10842,N_9481,N_9623);
nand U10843 (N_10843,N_7779,N_8583);
xor U10844 (N_10844,N_8763,N_8082);
and U10845 (N_10845,N_8565,N_7841);
nand U10846 (N_10846,N_7868,N_8100);
and U10847 (N_10847,N_7565,N_9326);
or U10848 (N_10848,N_8368,N_9874);
or U10849 (N_10849,N_7969,N_7654);
nor U10850 (N_10850,N_9332,N_9520);
nand U10851 (N_10851,N_8294,N_8210);
nand U10852 (N_10852,N_7700,N_7880);
nor U10853 (N_10853,N_8744,N_7584);
and U10854 (N_10854,N_9234,N_7923);
and U10855 (N_10855,N_8528,N_8460);
nand U10856 (N_10856,N_8980,N_7579);
and U10857 (N_10857,N_9658,N_7734);
and U10858 (N_10858,N_8637,N_9385);
nand U10859 (N_10859,N_8675,N_9563);
nand U10860 (N_10860,N_9597,N_9723);
or U10861 (N_10861,N_8697,N_8163);
nand U10862 (N_10862,N_9362,N_8950);
nand U10863 (N_10863,N_9062,N_8760);
nor U10864 (N_10864,N_9421,N_9089);
and U10865 (N_10865,N_8329,N_9570);
nand U10866 (N_10866,N_9449,N_8296);
nor U10867 (N_10867,N_9299,N_8168);
or U10868 (N_10868,N_8410,N_9769);
nor U10869 (N_10869,N_9095,N_8255);
and U10870 (N_10870,N_9339,N_8976);
and U10871 (N_10871,N_8015,N_8512);
nor U10872 (N_10872,N_7827,N_9387);
and U10873 (N_10873,N_8234,N_9569);
and U10874 (N_10874,N_9026,N_8491);
nor U10875 (N_10875,N_8687,N_8928);
xnor U10876 (N_10876,N_9625,N_8599);
xor U10877 (N_10877,N_7844,N_8380);
and U10878 (N_10878,N_9051,N_9252);
nand U10879 (N_10879,N_8531,N_9643);
and U10880 (N_10880,N_7942,N_9418);
nand U10881 (N_10881,N_8728,N_8447);
nor U10882 (N_10882,N_9891,N_7877);
nand U10883 (N_10883,N_8197,N_8864);
nand U10884 (N_10884,N_8851,N_8301);
nand U10885 (N_10885,N_9888,N_8411);
and U10886 (N_10886,N_9969,N_8719);
nand U10887 (N_10887,N_8567,N_7612);
and U10888 (N_10888,N_8124,N_8958);
or U10889 (N_10889,N_8207,N_8126);
or U10890 (N_10890,N_7889,N_9714);
nand U10891 (N_10891,N_9522,N_8046);
or U10892 (N_10892,N_8420,N_9476);
and U10893 (N_10893,N_9513,N_8385);
nor U10894 (N_10894,N_9776,N_9514);
and U10895 (N_10895,N_8738,N_8555);
nand U10896 (N_10896,N_9006,N_8648);
nand U10897 (N_10897,N_7586,N_9995);
or U10898 (N_10898,N_9347,N_9404);
and U10899 (N_10899,N_8057,N_8563);
xor U10900 (N_10900,N_9695,N_8766);
xnor U10901 (N_10901,N_9750,N_9355);
xor U10902 (N_10902,N_8603,N_9411);
nor U10903 (N_10903,N_9178,N_9040);
nor U10904 (N_10904,N_8388,N_9164);
and U10905 (N_10905,N_9704,N_8040);
or U10906 (N_10906,N_8044,N_8369);
nand U10907 (N_10907,N_9864,N_8998);
xnor U10908 (N_10908,N_9678,N_8415);
nand U10909 (N_10909,N_8578,N_7681);
nand U10910 (N_10910,N_9108,N_7964);
and U10911 (N_10911,N_7807,N_9711);
nand U10912 (N_10912,N_7649,N_7893);
xor U10913 (N_10913,N_8467,N_7764);
nor U10914 (N_10914,N_9903,N_8493);
or U10915 (N_10915,N_8521,N_8956);
nor U10916 (N_10916,N_9985,N_7915);
nor U10917 (N_10917,N_7986,N_8849);
nand U10918 (N_10918,N_8007,N_8389);
nor U10919 (N_10919,N_9009,N_9044);
nand U10920 (N_10920,N_9300,N_8973);
and U10921 (N_10921,N_9204,N_8797);
nor U10922 (N_10922,N_8060,N_8188);
nand U10923 (N_10923,N_8326,N_8112);
nor U10924 (N_10924,N_9083,N_9962);
or U10925 (N_10925,N_8196,N_8900);
nand U10926 (N_10926,N_8143,N_9306);
or U10927 (N_10927,N_8053,N_9581);
or U10928 (N_10928,N_7998,N_9545);
nor U10929 (N_10929,N_7543,N_9978);
or U10930 (N_10930,N_9706,N_7738);
or U10931 (N_10931,N_9475,N_9937);
nor U10932 (N_10932,N_9289,N_8193);
xor U10933 (N_10933,N_7953,N_9881);
or U10934 (N_10934,N_7993,N_7784);
nor U10935 (N_10935,N_9146,N_9989);
nand U10936 (N_10936,N_9170,N_8230);
nor U10937 (N_10937,N_8208,N_8302);
and U10938 (N_10938,N_9862,N_8779);
nor U10939 (N_10939,N_7502,N_8366);
or U10940 (N_10940,N_7768,N_8374);
or U10941 (N_10941,N_8351,N_9761);
and U10942 (N_10942,N_8147,N_9998);
xnor U10943 (N_10943,N_9533,N_8362);
nand U10944 (N_10944,N_9356,N_7501);
or U10945 (N_10945,N_9861,N_9217);
nor U10946 (N_10946,N_9333,N_9954);
or U10947 (N_10947,N_8132,N_9413);
and U10948 (N_10948,N_8670,N_7806);
xnor U10949 (N_10949,N_8280,N_9005);
xor U10950 (N_10950,N_7924,N_9550);
nand U10951 (N_10951,N_9091,N_7610);
nor U10952 (N_10952,N_8395,N_9388);
xor U10953 (N_10953,N_9698,N_7604);
and U10954 (N_10954,N_9030,N_8249);
and U10955 (N_10955,N_8967,N_8840);
or U10956 (N_10956,N_7589,N_9485);
and U10957 (N_10957,N_8206,N_9271);
xnor U10958 (N_10958,N_9712,N_9800);
or U10959 (N_10959,N_8299,N_8473);
nor U10960 (N_10960,N_7963,N_7670);
and U10961 (N_10961,N_9610,N_7956);
and U10962 (N_10962,N_7509,N_8272);
nand U10963 (N_10963,N_7627,N_9718);
nor U10964 (N_10964,N_9023,N_9439);
nor U10965 (N_10965,N_8117,N_8285);
nor U10966 (N_10966,N_8787,N_7839);
or U10967 (N_10967,N_7849,N_7675);
or U10968 (N_10968,N_8661,N_8641);
and U10969 (N_10969,N_8907,N_8812);
nor U10970 (N_10970,N_8709,N_8312);
nand U10971 (N_10971,N_8434,N_8672);
nand U10972 (N_10972,N_8290,N_9764);
nand U10973 (N_10973,N_9524,N_9855);
xnor U10974 (N_10974,N_9463,N_8991);
nor U10975 (N_10975,N_8274,N_9494);
or U10976 (N_10976,N_7698,N_9013);
and U10977 (N_10977,N_7607,N_8612);
or U10978 (N_10978,N_9840,N_8677);
or U10979 (N_10979,N_8690,N_8386);
and U10980 (N_10980,N_9086,N_9228);
nor U10981 (N_10981,N_9921,N_9455);
or U10982 (N_10982,N_8624,N_9974);
xnor U10983 (N_10983,N_9636,N_9807);
nor U10984 (N_10984,N_8914,N_8587);
nor U10985 (N_10985,N_8471,N_8033);
and U10986 (N_10986,N_9141,N_7825);
nor U10987 (N_10987,N_8938,N_8805);
nor U10988 (N_10988,N_8941,N_7537);
xor U10989 (N_10989,N_8146,N_8194);
xor U10990 (N_10990,N_8847,N_9004);
or U10991 (N_10991,N_7733,N_7823);
xor U10992 (N_10992,N_8872,N_9261);
nor U10993 (N_10993,N_8894,N_9179);
or U10994 (N_10994,N_7782,N_7714);
and U10995 (N_10995,N_7692,N_7526);
nor U10996 (N_10996,N_9756,N_9788);
nand U10997 (N_10997,N_8926,N_9956);
nand U10998 (N_10998,N_9773,N_7548);
xnor U10999 (N_10999,N_8899,N_8421);
and U11000 (N_11000,N_9327,N_7618);
nor U11001 (N_11001,N_8319,N_8113);
and U11002 (N_11002,N_7647,N_9556);
nor U11003 (N_11003,N_9890,N_9407);
nand U11004 (N_11004,N_8042,N_8853);
xor U11005 (N_11005,N_9946,N_8355);
nor U11006 (N_11006,N_8826,N_8247);
nand U11007 (N_11007,N_8618,N_9991);
nor U11008 (N_11008,N_7801,N_9549);
nor U11009 (N_11009,N_7836,N_9920);
and U11010 (N_11010,N_8568,N_9487);
xnor U11011 (N_11011,N_8192,N_8038);
and U11012 (N_11012,N_8347,N_8905);
nand U11013 (N_11013,N_8701,N_9283);
nor U11014 (N_11014,N_8432,N_8758);
and U11015 (N_11015,N_8472,N_9639);
and U11016 (N_11016,N_9815,N_9163);
and U11017 (N_11017,N_7522,N_9360);
nand U11018 (N_11018,N_7874,N_9264);
nand U11019 (N_11019,N_8880,N_9586);
nor U11020 (N_11020,N_9654,N_7525);
and U11021 (N_11021,N_9934,N_8995);
nor U11022 (N_11022,N_9774,N_8519);
and U11023 (N_11023,N_7843,N_8532);
nor U11024 (N_11024,N_7658,N_7643);
and U11025 (N_11025,N_8145,N_9525);
nand U11026 (N_11026,N_9226,N_8908);
and U11027 (N_11027,N_9405,N_8653);
and U11028 (N_11028,N_9209,N_8772);
nand U11029 (N_11029,N_7974,N_8922);
nand U11030 (N_11030,N_8875,N_9448);
or U11031 (N_11031,N_7605,N_7724);
or U11032 (N_11032,N_7552,N_8039);
and U11033 (N_11033,N_9381,N_9287);
xnor U11034 (N_11034,N_7908,N_7638);
and U11035 (N_11035,N_9745,N_9877);
or U11036 (N_11036,N_8747,N_9175);
nand U11037 (N_11037,N_9336,N_8986);
nand U11038 (N_11038,N_8391,N_8343);
or U11039 (N_11039,N_9301,N_8706);
xor U11040 (N_11040,N_8092,N_8456);
and U11041 (N_11041,N_9136,N_9763);
or U11042 (N_11042,N_9331,N_9748);
nor U11043 (N_11043,N_7797,N_7775);
or U11044 (N_11044,N_9500,N_8634);
nand U11045 (N_11045,N_7697,N_8920);
or U11046 (N_11046,N_9622,N_9538);
xor U11047 (N_11047,N_8940,N_9012);
and U11048 (N_11048,N_8068,N_8504);
and U11049 (N_11049,N_9565,N_9527);
nor U11050 (N_11050,N_8981,N_9137);
or U11051 (N_11051,N_9651,N_8708);
nor U11052 (N_11052,N_7980,N_8360);
and U11053 (N_11053,N_7962,N_8418);
nor U11054 (N_11054,N_9936,N_8691);
nand U11055 (N_11055,N_8560,N_9357);
nor U11056 (N_11056,N_8845,N_9790);
and U11057 (N_11057,N_8150,N_9134);
and U11058 (N_11058,N_9378,N_7636);
and U11059 (N_11059,N_9838,N_7601);
xnor U11060 (N_11060,N_9414,N_9288);
or U11061 (N_11061,N_9241,N_9676);
nor U11062 (N_11062,N_8358,N_8352);
or U11063 (N_11063,N_8273,N_9148);
or U11064 (N_11064,N_8788,N_9215);
and U11065 (N_11065,N_8263,N_7834);
or U11066 (N_11066,N_9592,N_8189);
nand U11067 (N_11067,N_8262,N_9917);
or U11068 (N_11068,N_9181,N_9738);
and U11069 (N_11069,N_9059,N_8534);
and U11070 (N_11070,N_7884,N_7952);
or U11071 (N_11071,N_9486,N_9966);
xor U11072 (N_11072,N_9248,N_7742);
nor U11073 (N_11073,N_7505,N_8999);
and U11074 (N_11074,N_8087,N_7981);
nor U11075 (N_11075,N_7711,N_8338);
nand U11076 (N_11076,N_9725,N_9703);
nand U11077 (N_11077,N_8202,N_8478);
and U11078 (N_11078,N_7728,N_8149);
nand U11079 (N_11079,N_9430,N_9055);
or U11080 (N_11080,N_9737,N_9833);
nor U11081 (N_11081,N_9468,N_9943);
nand U11082 (N_11082,N_8627,N_8781);
or U11083 (N_11083,N_9361,N_7660);
or U11084 (N_11084,N_8232,N_7555);
or U11085 (N_11085,N_9434,N_7557);
and U11086 (N_11086,N_8371,N_7776);
xor U11087 (N_11087,N_9841,N_8683);
nor U11088 (N_11088,N_9325,N_8424);
or U11089 (N_11089,N_9391,N_8224);
or U11090 (N_11090,N_9708,N_9568);
or U11091 (N_11091,N_8501,N_7751);
and U11092 (N_11092,N_7965,N_7674);
nand U11093 (N_11093,N_9318,N_8256);
nor U11094 (N_11094,N_8754,N_9617);
and U11095 (N_11095,N_8067,N_7904);
or U11096 (N_11096,N_9483,N_8579);
nand U11097 (N_11097,N_8002,N_9650);
and U11098 (N_11098,N_7918,N_8404);
or U11099 (N_11099,N_7524,N_9515);
nor U11100 (N_11100,N_9402,N_7575);
nand U11101 (N_11101,N_7829,N_8759);
nor U11102 (N_11102,N_8409,N_8768);
nor U11103 (N_11103,N_9165,N_8077);
nand U11104 (N_11104,N_8711,N_9941);
and U11105 (N_11105,N_8593,N_8403);
and U11106 (N_11106,N_9879,N_8487);
or U11107 (N_11107,N_8917,N_7592);
nor U11108 (N_11108,N_8219,N_9871);
or U11109 (N_11109,N_9380,N_9454);
or U11110 (N_11110,N_8510,N_8153);
or U11111 (N_11111,N_8012,N_9842);
or U11112 (N_11112,N_8031,N_9607);
nand U11113 (N_11113,N_9709,N_7858);
nand U11114 (N_11114,N_8874,N_8141);
nor U11115 (N_11115,N_9144,N_9406);
or U11116 (N_11116,N_9033,N_9344);
nor U11117 (N_11117,N_9927,N_7630);
and U11118 (N_11118,N_7906,N_9460);
or U11119 (N_11119,N_8963,N_7871);
xor U11120 (N_11120,N_9057,N_9782);
or U11121 (N_11121,N_9707,N_9792);
and U11122 (N_11122,N_8838,N_8590);
nand U11123 (N_11123,N_9211,N_7572);
nor U11124 (N_11124,N_9410,N_8458);
or U11125 (N_11125,N_9068,N_8536);
nor U11126 (N_11126,N_7835,N_9399);
or U11127 (N_11127,N_9045,N_9155);
and U11128 (N_11128,N_9594,N_9392);
and U11129 (N_11129,N_8600,N_8785);
and U11130 (N_11130,N_8245,N_7804);
nor U11131 (N_11131,N_7669,N_9517);
and U11132 (N_11132,N_8992,N_8771);
xnor U11133 (N_11133,N_8035,N_9542);
and U11134 (N_11134,N_8862,N_7585);
xnor U11135 (N_11135,N_7867,N_7568);
nor U11136 (N_11136,N_7622,N_7994);
nor U11137 (N_11137,N_7534,N_9427);
nand U11138 (N_11138,N_9993,N_8591);
nor U11139 (N_11139,N_9582,N_9310);
and U11140 (N_11140,N_9535,N_8841);
or U11141 (N_11141,N_8869,N_7854);
or U11142 (N_11142,N_8173,N_9145);
or U11143 (N_11143,N_7663,N_9000);
nand U11144 (N_11144,N_9971,N_8575);
nand U11145 (N_11145,N_9945,N_9697);
nand U11146 (N_11146,N_8054,N_9615);
and U11147 (N_11147,N_8780,N_9931);
and U11148 (N_11148,N_8394,N_7869);
nor U11149 (N_11149,N_8850,N_8745);
xor U11150 (N_11150,N_9014,N_9324);
nand U11151 (N_11151,N_9580,N_9624);
nand U11152 (N_11152,N_8608,N_7582);
nor U11153 (N_11153,N_8091,N_9583);
nor U11154 (N_11154,N_8679,N_8740);
xnor U11155 (N_11155,N_7741,N_7988);
nor U11156 (N_11156,N_7571,N_7542);
or U11157 (N_11157,N_7531,N_9100);
and U11158 (N_11158,N_8959,N_8830);
and U11159 (N_11159,N_9122,N_7944);
nand U11160 (N_11160,N_8462,N_9115);
xnor U11161 (N_11161,N_9220,N_9282);
or U11162 (N_11162,N_7631,N_7999);
nor U11163 (N_11163,N_8257,N_7735);
nor U11164 (N_11164,N_8644,N_9534);
xnor U11165 (N_11165,N_8984,N_9428);
nor U11166 (N_11166,N_7600,N_8107);
and U11167 (N_11167,N_9351,N_8334);
nor U11168 (N_11168,N_8306,N_8524);
or U11169 (N_11169,N_8375,N_9808);
nor U11170 (N_11170,N_7837,N_9078);
or U11171 (N_11171,N_7766,N_8019);
and U11172 (N_11172,N_8636,N_8898);
nor U11173 (N_11173,N_9469,N_8238);
nor U11174 (N_11174,N_7773,N_8799);
or U11175 (N_11175,N_8001,N_7833);
nor U11176 (N_11176,N_7979,N_8906);
nor U11177 (N_11177,N_9251,N_8325);
or U11178 (N_11178,N_9880,N_9236);
nand U11179 (N_11179,N_9948,N_9918);
or U11180 (N_11180,N_9604,N_9940);
or U11181 (N_11181,N_8592,N_9672);
and U11182 (N_11182,N_9609,N_9558);
or U11183 (N_11183,N_9608,N_7912);
nand U11184 (N_11184,N_9904,N_8861);
nor U11185 (N_11185,N_8886,N_8550);
nor U11186 (N_11186,N_8540,N_9474);
nand U11187 (N_11187,N_9673,N_9396);
and U11188 (N_11188,N_8461,N_8336);
nor U11189 (N_11189,N_8548,N_9810);
and U11190 (N_11190,N_7875,N_8488);
or U11191 (N_11191,N_9307,N_8601);
xor U11192 (N_11192,N_9662,N_8292);
and U11193 (N_11193,N_9216,N_8011);
nor U11194 (N_11194,N_9895,N_9394);
and U11195 (N_11195,N_8810,N_9593);
nand U11196 (N_11196,N_7606,N_8794);
or U11197 (N_11197,N_8818,N_8737);
nand U11198 (N_11198,N_8541,N_8729);
and U11199 (N_11199,N_9503,N_9768);
or U11200 (N_11200,N_8671,N_8549);
or U11201 (N_11201,N_9143,N_9981);
nand U11202 (N_11202,N_8225,N_9471);
and U11203 (N_11203,N_8345,N_9539);
nor U11204 (N_11204,N_7644,N_8026);
nand U11205 (N_11205,N_7590,N_7667);
xnor U11206 (N_11206,N_8517,N_8392);
nand U11207 (N_11207,N_8286,N_8520);
nor U11208 (N_11208,N_9670,N_7794);
nand U11209 (N_11209,N_8178,N_8795);
nand U11210 (N_11210,N_9691,N_9096);
nand U11211 (N_11211,N_9733,N_9011);
or U11212 (N_11212,N_9203,N_9848);
xnor U11213 (N_11213,N_7932,N_8735);
nor U11214 (N_11214,N_8902,N_8770);
xnor U11215 (N_11215,N_7687,N_8486);
nor U11216 (N_11216,N_7720,N_9849);
nand U11217 (N_11217,N_9110,N_7926);
or U11218 (N_11218,N_9286,N_7927);
nor U11219 (N_11219,N_8767,N_8058);
or U11220 (N_11220,N_9435,N_8717);
nand U11221 (N_11221,N_9281,N_9913);
or U11222 (N_11222,N_9253,N_8429);
and U11223 (N_11223,N_8655,N_7771);
nor U11224 (N_11224,N_8018,N_8131);
nor U11225 (N_11225,N_9139,N_9338);
or U11226 (N_11226,N_9935,N_8762);
xor U11227 (N_11227,N_9902,N_9859);
nor U11228 (N_11228,N_8960,N_8086);
and U11229 (N_11229,N_9789,N_7704);
nor U11230 (N_11230,N_9140,N_7679);
nor U11231 (N_11231,N_9965,N_9957);
nor U11232 (N_11232,N_9982,N_8994);
and U11233 (N_11233,N_8522,N_7677);
or U11234 (N_11234,N_8191,N_8983);
or U11235 (N_11235,N_8300,N_8453);
nor U11236 (N_11236,N_8674,N_7718);
nand U11237 (N_11237,N_7863,N_9403);
or U11238 (N_11238,N_8689,N_8496);
nor U11239 (N_11239,N_9992,N_9878);
nor U11240 (N_11240,N_8308,N_9684);
and U11241 (N_11241,N_9587,N_9566);
and U11242 (N_11242,N_7595,N_7894);
nand U11243 (N_11243,N_8911,N_9530);
nand U11244 (N_11244,N_8530,N_8211);
nand U11245 (N_11245,N_8824,N_8248);
nor U11246 (N_11246,N_8036,N_9443);
or U11247 (N_11247,N_9383,N_7818);
or U11248 (N_11248,N_7632,N_9161);
or U11249 (N_11249,N_8947,N_9050);
nor U11250 (N_11250,N_8824,N_7714);
nand U11251 (N_11251,N_7665,N_9047);
nand U11252 (N_11252,N_7589,N_9480);
xnor U11253 (N_11253,N_7626,N_8004);
nor U11254 (N_11254,N_9296,N_9381);
nand U11255 (N_11255,N_7900,N_8240);
and U11256 (N_11256,N_7598,N_8152);
nand U11257 (N_11257,N_7658,N_8420);
or U11258 (N_11258,N_7612,N_8260);
nand U11259 (N_11259,N_7916,N_7729);
or U11260 (N_11260,N_8848,N_8591);
xnor U11261 (N_11261,N_9027,N_9826);
nor U11262 (N_11262,N_7635,N_9041);
nor U11263 (N_11263,N_9495,N_9014);
nand U11264 (N_11264,N_9345,N_8855);
and U11265 (N_11265,N_8935,N_9193);
nor U11266 (N_11266,N_7653,N_7724);
nor U11267 (N_11267,N_9328,N_8794);
and U11268 (N_11268,N_8363,N_9025);
or U11269 (N_11269,N_7604,N_9992);
nand U11270 (N_11270,N_9447,N_9351);
and U11271 (N_11271,N_7789,N_8412);
xnor U11272 (N_11272,N_9104,N_8232);
and U11273 (N_11273,N_9959,N_8632);
and U11274 (N_11274,N_8474,N_9272);
xnor U11275 (N_11275,N_8928,N_9933);
xnor U11276 (N_11276,N_9213,N_8357);
and U11277 (N_11277,N_7898,N_8624);
nand U11278 (N_11278,N_7589,N_9816);
nand U11279 (N_11279,N_8801,N_8286);
and U11280 (N_11280,N_7860,N_8843);
nand U11281 (N_11281,N_9371,N_8266);
and U11282 (N_11282,N_9065,N_7816);
nor U11283 (N_11283,N_9337,N_7948);
nor U11284 (N_11284,N_8774,N_8706);
nor U11285 (N_11285,N_8447,N_8232);
and U11286 (N_11286,N_8076,N_9032);
nand U11287 (N_11287,N_8786,N_7715);
xnor U11288 (N_11288,N_8707,N_9109);
and U11289 (N_11289,N_7670,N_8387);
xnor U11290 (N_11290,N_9834,N_9650);
or U11291 (N_11291,N_8070,N_9930);
or U11292 (N_11292,N_7657,N_8056);
and U11293 (N_11293,N_9839,N_9383);
or U11294 (N_11294,N_8270,N_9515);
or U11295 (N_11295,N_8643,N_7699);
nor U11296 (N_11296,N_7983,N_7644);
nor U11297 (N_11297,N_9165,N_7672);
and U11298 (N_11298,N_9099,N_7734);
nor U11299 (N_11299,N_8399,N_7845);
nand U11300 (N_11300,N_9712,N_8577);
nand U11301 (N_11301,N_9943,N_8718);
and U11302 (N_11302,N_7636,N_7626);
or U11303 (N_11303,N_8137,N_9497);
and U11304 (N_11304,N_7906,N_8974);
nand U11305 (N_11305,N_9770,N_8743);
and U11306 (N_11306,N_9910,N_7955);
xor U11307 (N_11307,N_9767,N_9405);
nand U11308 (N_11308,N_9121,N_8250);
and U11309 (N_11309,N_7650,N_8072);
nand U11310 (N_11310,N_8770,N_9614);
and U11311 (N_11311,N_8595,N_9196);
or U11312 (N_11312,N_9306,N_8065);
nand U11313 (N_11313,N_8380,N_8217);
and U11314 (N_11314,N_8049,N_8410);
nand U11315 (N_11315,N_8350,N_8016);
and U11316 (N_11316,N_7794,N_8957);
and U11317 (N_11317,N_9464,N_8257);
and U11318 (N_11318,N_8548,N_8618);
or U11319 (N_11319,N_8783,N_9307);
or U11320 (N_11320,N_9030,N_7876);
xnor U11321 (N_11321,N_7875,N_7899);
nor U11322 (N_11322,N_8665,N_9212);
nor U11323 (N_11323,N_8092,N_8622);
xnor U11324 (N_11324,N_8378,N_9081);
or U11325 (N_11325,N_8096,N_9748);
or U11326 (N_11326,N_9630,N_7987);
nand U11327 (N_11327,N_9294,N_9158);
nor U11328 (N_11328,N_8084,N_9868);
and U11329 (N_11329,N_9760,N_9213);
or U11330 (N_11330,N_7506,N_9480);
nor U11331 (N_11331,N_8297,N_8303);
and U11332 (N_11332,N_8531,N_9074);
nor U11333 (N_11333,N_8736,N_7824);
and U11334 (N_11334,N_8495,N_9670);
and U11335 (N_11335,N_7633,N_8861);
and U11336 (N_11336,N_8007,N_7680);
nor U11337 (N_11337,N_9743,N_7861);
nand U11338 (N_11338,N_8369,N_9324);
nor U11339 (N_11339,N_9206,N_9696);
or U11340 (N_11340,N_7554,N_7960);
and U11341 (N_11341,N_7516,N_8260);
nor U11342 (N_11342,N_7519,N_9020);
or U11343 (N_11343,N_8130,N_8588);
or U11344 (N_11344,N_8903,N_8810);
nor U11345 (N_11345,N_9290,N_8986);
nand U11346 (N_11346,N_9737,N_9822);
or U11347 (N_11347,N_8817,N_9203);
and U11348 (N_11348,N_9160,N_7984);
and U11349 (N_11349,N_8056,N_8826);
nand U11350 (N_11350,N_7799,N_8417);
xnor U11351 (N_11351,N_8475,N_9929);
nand U11352 (N_11352,N_7865,N_8088);
nand U11353 (N_11353,N_8843,N_8036);
and U11354 (N_11354,N_9292,N_8529);
nand U11355 (N_11355,N_8545,N_7721);
xor U11356 (N_11356,N_7865,N_7970);
nor U11357 (N_11357,N_9208,N_8269);
or U11358 (N_11358,N_7776,N_9605);
nor U11359 (N_11359,N_8829,N_7810);
nand U11360 (N_11360,N_7978,N_8241);
and U11361 (N_11361,N_8931,N_9611);
nor U11362 (N_11362,N_9007,N_7620);
nand U11363 (N_11363,N_8430,N_8580);
or U11364 (N_11364,N_9310,N_8568);
nand U11365 (N_11365,N_7800,N_8012);
nor U11366 (N_11366,N_9501,N_8251);
nor U11367 (N_11367,N_7781,N_8747);
nor U11368 (N_11368,N_7806,N_8084);
nor U11369 (N_11369,N_8234,N_7829);
nand U11370 (N_11370,N_9418,N_8173);
nor U11371 (N_11371,N_8704,N_9130);
nand U11372 (N_11372,N_9889,N_8333);
nor U11373 (N_11373,N_8228,N_7558);
nand U11374 (N_11374,N_7744,N_9393);
and U11375 (N_11375,N_9618,N_9798);
xnor U11376 (N_11376,N_9846,N_9573);
nor U11377 (N_11377,N_9631,N_8949);
nor U11378 (N_11378,N_9268,N_9570);
nand U11379 (N_11379,N_8243,N_8594);
or U11380 (N_11380,N_8720,N_7947);
nand U11381 (N_11381,N_7531,N_7889);
nand U11382 (N_11382,N_8377,N_8648);
nand U11383 (N_11383,N_8758,N_8974);
nand U11384 (N_11384,N_8539,N_9100);
or U11385 (N_11385,N_7513,N_9916);
or U11386 (N_11386,N_8183,N_9370);
or U11387 (N_11387,N_9026,N_9139);
and U11388 (N_11388,N_7976,N_8582);
and U11389 (N_11389,N_7837,N_8417);
nor U11390 (N_11390,N_9554,N_9426);
nor U11391 (N_11391,N_9288,N_8276);
xor U11392 (N_11392,N_8305,N_9570);
nand U11393 (N_11393,N_8326,N_8813);
nor U11394 (N_11394,N_8056,N_8734);
and U11395 (N_11395,N_9258,N_9913);
and U11396 (N_11396,N_8983,N_9895);
nand U11397 (N_11397,N_9448,N_7539);
xor U11398 (N_11398,N_7733,N_8846);
and U11399 (N_11399,N_8238,N_7894);
nor U11400 (N_11400,N_9224,N_8279);
nand U11401 (N_11401,N_8955,N_7952);
or U11402 (N_11402,N_8247,N_7970);
nor U11403 (N_11403,N_8331,N_8553);
or U11404 (N_11404,N_8163,N_9513);
or U11405 (N_11405,N_9731,N_9000);
xnor U11406 (N_11406,N_9843,N_8370);
nand U11407 (N_11407,N_9837,N_9805);
nor U11408 (N_11408,N_8477,N_8867);
nand U11409 (N_11409,N_8429,N_7984);
nand U11410 (N_11410,N_9492,N_9791);
and U11411 (N_11411,N_9824,N_9516);
nor U11412 (N_11412,N_9731,N_8617);
nand U11413 (N_11413,N_7530,N_9316);
nand U11414 (N_11414,N_8257,N_9405);
nand U11415 (N_11415,N_9283,N_7835);
nand U11416 (N_11416,N_8765,N_8402);
nor U11417 (N_11417,N_8926,N_8630);
and U11418 (N_11418,N_9125,N_9707);
or U11419 (N_11419,N_7614,N_9168);
and U11420 (N_11420,N_7616,N_7694);
nand U11421 (N_11421,N_8660,N_8190);
nor U11422 (N_11422,N_9412,N_9429);
and U11423 (N_11423,N_8599,N_9507);
xor U11424 (N_11424,N_8735,N_9089);
or U11425 (N_11425,N_8131,N_8903);
and U11426 (N_11426,N_7695,N_8427);
and U11427 (N_11427,N_9043,N_8709);
xor U11428 (N_11428,N_7867,N_9860);
xnor U11429 (N_11429,N_9249,N_9695);
and U11430 (N_11430,N_9203,N_9024);
nand U11431 (N_11431,N_8267,N_9101);
or U11432 (N_11432,N_8598,N_8694);
or U11433 (N_11433,N_9811,N_7660);
or U11434 (N_11434,N_7770,N_8907);
nand U11435 (N_11435,N_7797,N_9711);
and U11436 (N_11436,N_8114,N_9821);
nand U11437 (N_11437,N_9079,N_8148);
nor U11438 (N_11438,N_9353,N_9251);
and U11439 (N_11439,N_8219,N_9665);
nand U11440 (N_11440,N_8290,N_8364);
nor U11441 (N_11441,N_7824,N_8738);
and U11442 (N_11442,N_9530,N_7628);
nor U11443 (N_11443,N_9277,N_8064);
nand U11444 (N_11444,N_9210,N_7825);
and U11445 (N_11445,N_8228,N_8066);
and U11446 (N_11446,N_7734,N_8734);
xnor U11447 (N_11447,N_8358,N_9514);
xnor U11448 (N_11448,N_8327,N_8854);
or U11449 (N_11449,N_9644,N_8953);
or U11450 (N_11450,N_9144,N_7867);
nor U11451 (N_11451,N_7743,N_8186);
xnor U11452 (N_11452,N_9864,N_9575);
nor U11453 (N_11453,N_8188,N_8847);
nand U11454 (N_11454,N_8995,N_7816);
nand U11455 (N_11455,N_8389,N_9179);
xnor U11456 (N_11456,N_8491,N_9028);
nor U11457 (N_11457,N_8948,N_9712);
nor U11458 (N_11458,N_9170,N_9432);
nor U11459 (N_11459,N_9181,N_7623);
xnor U11460 (N_11460,N_8139,N_7752);
nand U11461 (N_11461,N_9090,N_9193);
nor U11462 (N_11462,N_9088,N_9628);
nand U11463 (N_11463,N_9596,N_9725);
or U11464 (N_11464,N_8720,N_8249);
and U11465 (N_11465,N_9819,N_9294);
xnor U11466 (N_11466,N_9274,N_9544);
xnor U11467 (N_11467,N_8818,N_7636);
and U11468 (N_11468,N_9996,N_9858);
nand U11469 (N_11469,N_8593,N_7561);
and U11470 (N_11470,N_8447,N_9617);
nand U11471 (N_11471,N_9619,N_8956);
and U11472 (N_11472,N_7620,N_9024);
or U11473 (N_11473,N_9971,N_8290);
or U11474 (N_11474,N_8591,N_8056);
nand U11475 (N_11475,N_7652,N_9232);
nand U11476 (N_11476,N_9882,N_8006);
nor U11477 (N_11477,N_7826,N_9384);
or U11478 (N_11478,N_9708,N_7684);
nand U11479 (N_11479,N_7560,N_8116);
and U11480 (N_11480,N_9841,N_9448);
nor U11481 (N_11481,N_9648,N_8095);
or U11482 (N_11482,N_9367,N_9079);
nand U11483 (N_11483,N_8203,N_9219);
nand U11484 (N_11484,N_9058,N_9183);
nand U11485 (N_11485,N_8852,N_8896);
or U11486 (N_11486,N_7749,N_7987);
nor U11487 (N_11487,N_9108,N_9008);
xor U11488 (N_11488,N_7875,N_8556);
or U11489 (N_11489,N_9052,N_8808);
or U11490 (N_11490,N_8299,N_8862);
and U11491 (N_11491,N_7500,N_9880);
nand U11492 (N_11492,N_9898,N_8785);
nand U11493 (N_11493,N_9377,N_9986);
and U11494 (N_11494,N_7956,N_9776);
nand U11495 (N_11495,N_9702,N_7952);
and U11496 (N_11496,N_8555,N_8185);
or U11497 (N_11497,N_9795,N_7950);
nor U11498 (N_11498,N_8134,N_9861);
xnor U11499 (N_11499,N_7804,N_8511);
and U11500 (N_11500,N_7505,N_8191);
nand U11501 (N_11501,N_9978,N_7814);
nand U11502 (N_11502,N_8808,N_8778);
or U11503 (N_11503,N_7742,N_7507);
and U11504 (N_11504,N_9407,N_9172);
and U11505 (N_11505,N_7599,N_8000);
nand U11506 (N_11506,N_8207,N_7989);
or U11507 (N_11507,N_8592,N_8021);
nor U11508 (N_11508,N_8423,N_7852);
nand U11509 (N_11509,N_9944,N_9239);
nand U11510 (N_11510,N_7621,N_7707);
nor U11511 (N_11511,N_9455,N_9700);
or U11512 (N_11512,N_7653,N_9146);
nor U11513 (N_11513,N_8221,N_7607);
or U11514 (N_11514,N_8999,N_8939);
and U11515 (N_11515,N_8376,N_9810);
and U11516 (N_11516,N_9839,N_9374);
or U11517 (N_11517,N_7921,N_8707);
and U11518 (N_11518,N_9115,N_7818);
nor U11519 (N_11519,N_8564,N_8841);
xnor U11520 (N_11520,N_8877,N_9089);
nor U11521 (N_11521,N_8537,N_9644);
nor U11522 (N_11522,N_7957,N_7582);
and U11523 (N_11523,N_7731,N_9310);
nand U11524 (N_11524,N_8277,N_8404);
nor U11525 (N_11525,N_8893,N_8875);
nor U11526 (N_11526,N_8844,N_7583);
nand U11527 (N_11527,N_9930,N_9779);
nor U11528 (N_11528,N_8664,N_7829);
and U11529 (N_11529,N_9805,N_8814);
or U11530 (N_11530,N_9416,N_7681);
and U11531 (N_11531,N_9304,N_7517);
and U11532 (N_11532,N_7803,N_9044);
nor U11533 (N_11533,N_9814,N_9909);
nand U11534 (N_11534,N_9287,N_7769);
and U11535 (N_11535,N_7954,N_8528);
nor U11536 (N_11536,N_9228,N_8396);
and U11537 (N_11537,N_8651,N_7776);
and U11538 (N_11538,N_8550,N_8870);
nand U11539 (N_11539,N_9094,N_8001);
nor U11540 (N_11540,N_9784,N_7738);
or U11541 (N_11541,N_9762,N_7821);
nor U11542 (N_11542,N_7742,N_8366);
nand U11543 (N_11543,N_8050,N_9892);
and U11544 (N_11544,N_8189,N_9688);
or U11545 (N_11545,N_7656,N_8705);
and U11546 (N_11546,N_7584,N_8439);
nand U11547 (N_11547,N_9425,N_7939);
and U11548 (N_11548,N_9342,N_8855);
nand U11549 (N_11549,N_8357,N_9473);
or U11550 (N_11550,N_8094,N_7903);
nor U11551 (N_11551,N_8572,N_9299);
and U11552 (N_11552,N_7936,N_7720);
and U11553 (N_11553,N_7702,N_9841);
or U11554 (N_11554,N_7644,N_8712);
or U11555 (N_11555,N_8870,N_9311);
nor U11556 (N_11556,N_9454,N_8292);
nor U11557 (N_11557,N_8261,N_8421);
and U11558 (N_11558,N_9349,N_7951);
xor U11559 (N_11559,N_7756,N_8583);
or U11560 (N_11560,N_9398,N_7703);
nand U11561 (N_11561,N_9390,N_8653);
nand U11562 (N_11562,N_9415,N_9053);
nor U11563 (N_11563,N_9792,N_9091);
nor U11564 (N_11564,N_8694,N_8211);
nand U11565 (N_11565,N_7529,N_8298);
nor U11566 (N_11566,N_9382,N_9255);
nor U11567 (N_11567,N_9040,N_7571);
and U11568 (N_11568,N_8043,N_7894);
or U11569 (N_11569,N_7775,N_9484);
nand U11570 (N_11570,N_7774,N_8111);
nor U11571 (N_11571,N_8648,N_8408);
nor U11572 (N_11572,N_9012,N_8018);
nand U11573 (N_11573,N_7705,N_9985);
nand U11574 (N_11574,N_8118,N_7736);
nand U11575 (N_11575,N_9944,N_8281);
xnor U11576 (N_11576,N_8180,N_7857);
nand U11577 (N_11577,N_8394,N_9419);
or U11578 (N_11578,N_9021,N_8643);
nor U11579 (N_11579,N_9618,N_8585);
nand U11580 (N_11580,N_9897,N_9042);
nand U11581 (N_11581,N_9154,N_7997);
nor U11582 (N_11582,N_8235,N_9655);
and U11583 (N_11583,N_7715,N_9575);
and U11584 (N_11584,N_8017,N_9663);
or U11585 (N_11585,N_9281,N_8886);
or U11586 (N_11586,N_9903,N_9127);
nand U11587 (N_11587,N_8380,N_8226);
nor U11588 (N_11588,N_9898,N_9350);
and U11589 (N_11589,N_9107,N_9334);
xor U11590 (N_11590,N_7961,N_8931);
or U11591 (N_11591,N_9347,N_8208);
and U11592 (N_11592,N_8580,N_7881);
xor U11593 (N_11593,N_8093,N_8554);
and U11594 (N_11594,N_7511,N_8312);
xnor U11595 (N_11595,N_8870,N_9323);
nand U11596 (N_11596,N_8885,N_9888);
and U11597 (N_11597,N_9795,N_7989);
nand U11598 (N_11598,N_7590,N_9539);
and U11599 (N_11599,N_8110,N_8847);
nand U11600 (N_11600,N_9235,N_8583);
and U11601 (N_11601,N_7797,N_9775);
nor U11602 (N_11602,N_8730,N_9390);
and U11603 (N_11603,N_8552,N_9618);
nor U11604 (N_11604,N_8961,N_8331);
and U11605 (N_11605,N_9678,N_8875);
or U11606 (N_11606,N_8647,N_8583);
nand U11607 (N_11607,N_8624,N_8042);
and U11608 (N_11608,N_7789,N_8279);
nand U11609 (N_11609,N_9381,N_9852);
nand U11610 (N_11610,N_8673,N_9535);
xor U11611 (N_11611,N_8730,N_9982);
nor U11612 (N_11612,N_9640,N_8323);
nor U11613 (N_11613,N_9367,N_8291);
and U11614 (N_11614,N_8010,N_9786);
and U11615 (N_11615,N_8916,N_7786);
and U11616 (N_11616,N_8481,N_7540);
nand U11617 (N_11617,N_9136,N_8166);
nand U11618 (N_11618,N_8985,N_7695);
and U11619 (N_11619,N_8679,N_8750);
and U11620 (N_11620,N_8527,N_8706);
nand U11621 (N_11621,N_8427,N_9745);
nand U11622 (N_11622,N_8277,N_9851);
nor U11623 (N_11623,N_8206,N_9733);
nor U11624 (N_11624,N_9933,N_8029);
nand U11625 (N_11625,N_9738,N_8916);
nor U11626 (N_11626,N_7545,N_8187);
xnor U11627 (N_11627,N_8933,N_7690);
nor U11628 (N_11628,N_8316,N_9864);
nor U11629 (N_11629,N_9818,N_8781);
nor U11630 (N_11630,N_9726,N_7602);
or U11631 (N_11631,N_9444,N_8947);
and U11632 (N_11632,N_7576,N_8719);
or U11633 (N_11633,N_8103,N_7969);
and U11634 (N_11634,N_7879,N_8746);
nand U11635 (N_11635,N_7513,N_8031);
or U11636 (N_11636,N_9972,N_8713);
or U11637 (N_11637,N_9745,N_8203);
nand U11638 (N_11638,N_9659,N_7755);
or U11639 (N_11639,N_9339,N_7516);
and U11640 (N_11640,N_8475,N_7985);
xnor U11641 (N_11641,N_9389,N_9333);
nand U11642 (N_11642,N_8634,N_8230);
nand U11643 (N_11643,N_9454,N_9819);
and U11644 (N_11644,N_9784,N_9543);
nor U11645 (N_11645,N_8979,N_8368);
or U11646 (N_11646,N_7787,N_9949);
nand U11647 (N_11647,N_8459,N_8270);
nor U11648 (N_11648,N_8727,N_9661);
nor U11649 (N_11649,N_8060,N_7749);
and U11650 (N_11650,N_9238,N_9329);
nor U11651 (N_11651,N_9335,N_7612);
nand U11652 (N_11652,N_8817,N_8543);
xor U11653 (N_11653,N_7683,N_7938);
or U11654 (N_11654,N_8873,N_8318);
or U11655 (N_11655,N_7625,N_8768);
nand U11656 (N_11656,N_8880,N_9927);
and U11657 (N_11657,N_8401,N_7856);
and U11658 (N_11658,N_8938,N_9210);
or U11659 (N_11659,N_8289,N_7509);
nand U11660 (N_11660,N_9777,N_7786);
nor U11661 (N_11661,N_9521,N_7923);
xnor U11662 (N_11662,N_9589,N_8844);
and U11663 (N_11663,N_9905,N_9128);
nand U11664 (N_11664,N_8000,N_9826);
nand U11665 (N_11665,N_9623,N_9901);
nand U11666 (N_11666,N_7700,N_8334);
nor U11667 (N_11667,N_8210,N_9951);
nor U11668 (N_11668,N_7663,N_8821);
nand U11669 (N_11669,N_9342,N_9382);
nor U11670 (N_11670,N_7905,N_7637);
and U11671 (N_11671,N_8205,N_8826);
or U11672 (N_11672,N_8576,N_7887);
xor U11673 (N_11673,N_9758,N_8993);
and U11674 (N_11674,N_9731,N_9761);
or U11675 (N_11675,N_8341,N_8479);
nand U11676 (N_11676,N_8572,N_8577);
nor U11677 (N_11677,N_7831,N_8376);
nand U11678 (N_11678,N_7672,N_8792);
and U11679 (N_11679,N_8012,N_7833);
or U11680 (N_11680,N_9207,N_7546);
nor U11681 (N_11681,N_7541,N_9847);
xnor U11682 (N_11682,N_8758,N_8025);
or U11683 (N_11683,N_7923,N_8580);
nand U11684 (N_11684,N_7699,N_7633);
xor U11685 (N_11685,N_8219,N_7812);
or U11686 (N_11686,N_8158,N_7938);
and U11687 (N_11687,N_9185,N_9325);
nor U11688 (N_11688,N_9321,N_7531);
or U11689 (N_11689,N_8667,N_7760);
or U11690 (N_11690,N_9045,N_8290);
nand U11691 (N_11691,N_9809,N_7697);
nand U11692 (N_11692,N_8797,N_9373);
or U11693 (N_11693,N_7619,N_8630);
nand U11694 (N_11694,N_8750,N_8259);
xor U11695 (N_11695,N_7677,N_8729);
or U11696 (N_11696,N_8405,N_7872);
nor U11697 (N_11697,N_8868,N_8083);
nand U11698 (N_11698,N_9146,N_7627);
and U11699 (N_11699,N_9585,N_7505);
xnor U11700 (N_11700,N_8013,N_9905);
nor U11701 (N_11701,N_9197,N_8775);
and U11702 (N_11702,N_9476,N_9594);
nand U11703 (N_11703,N_8028,N_9638);
nor U11704 (N_11704,N_9033,N_9452);
nand U11705 (N_11705,N_9827,N_7663);
nor U11706 (N_11706,N_8361,N_8903);
nor U11707 (N_11707,N_9116,N_8660);
or U11708 (N_11708,N_8308,N_8158);
xor U11709 (N_11709,N_9078,N_8063);
and U11710 (N_11710,N_9671,N_9699);
xnor U11711 (N_11711,N_9903,N_9880);
nor U11712 (N_11712,N_9505,N_8317);
nand U11713 (N_11713,N_8243,N_9662);
and U11714 (N_11714,N_8847,N_8551);
xnor U11715 (N_11715,N_7752,N_8997);
or U11716 (N_11716,N_7683,N_9186);
xnor U11717 (N_11717,N_8630,N_9228);
nor U11718 (N_11718,N_9976,N_9866);
and U11719 (N_11719,N_9772,N_7863);
and U11720 (N_11720,N_8506,N_7603);
and U11721 (N_11721,N_8689,N_8198);
or U11722 (N_11722,N_8396,N_7715);
or U11723 (N_11723,N_9610,N_9558);
xnor U11724 (N_11724,N_8817,N_8155);
nand U11725 (N_11725,N_9759,N_8203);
or U11726 (N_11726,N_9637,N_8437);
xnor U11727 (N_11727,N_8857,N_9448);
or U11728 (N_11728,N_7750,N_9567);
nand U11729 (N_11729,N_9394,N_8089);
and U11730 (N_11730,N_9456,N_7537);
nor U11731 (N_11731,N_8157,N_9113);
and U11732 (N_11732,N_8667,N_9561);
or U11733 (N_11733,N_8708,N_7731);
and U11734 (N_11734,N_7560,N_9756);
or U11735 (N_11735,N_9699,N_7785);
and U11736 (N_11736,N_9131,N_9827);
nand U11737 (N_11737,N_8176,N_9428);
or U11738 (N_11738,N_8041,N_8145);
xor U11739 (N_11739,N_7920,N_8474);
nand U11740 (N_11740,N_9385,N_8065);
or U11741 (N_11741,N_7734,N_9273);
nand U11742 (N_11742,N_9539,N_7914);
nor U11743 (N_11743,N_9898,N_8727);
or U11744 (N_11744,N_8585,N_8521);
nand U11745 (N_11745,N_9506,N_8190);
and U11746 (N_11746,N_9099,N_8237);
nor U11747 (N_11747,N_9288,N_7730);
or U11748 (N_11748,N_8212,N_8167);
or U11749 (N_11749,N_8725,N_9327);
or U11750 (N_11750,N_9458,N_8479);
and U11751 (N_11751,N_8365,N_8754);
and U11752 (N_11752,N_9425,N_8160);
nand U11753 (N_11753,N_7722,N_7742);
or U11754 (N_11754,N_9203,N_9454);
and U11755 (N_11755,N_9437,N_9929);
xnor U11756 (N_11756,N_7526,N_8811);
and U11757 (N_11757,N_8287,N_8036);
and U11758 (N_11758,N_8359,N_8322);
and U11759 (N_11759,N_9022,N_8756);
nor U11760 (N_11760,N_9605,N_8279);
nand U11761 (N_11761,N_9109,N_8121);
and U11762 (N_11762,N_8075,N_8519);
nor U11763 (N_11763,N_7627,N_9031);
nor U11764 (N_11764,N_7601,N_8328);
nand U11765 (N_11765,N_8947,N_7899);
nand U11766 (N_11766,N_8086,N_7858);
or U11767 (N_11767,N_9110,N_9626);
or U11768 (N_11768,N_7527,N_7594);
or U11769 (N_11769,N_9817,N_8649);
xnor U11770 (N_11770,N_9478,N_7721);
nor U11771 (N_11771,N_9992,N_9441);
or U11772 (N_11772,N_8776,N_9630);
or U11773 (N_11773,N_9840,N_7767);
nand U11774 (N_11774,N_7717,N_7858);
and U11775 (N_11775,N_9235,N_9607);
nor U11776 (N_11776,N_7880,N_8051);
or U11777 (N_11777,N_7645,N_7837);
and U11778 (N_11778,N_9066,N_7798);
or U11779 (N_11779,N_7797,N_8718);
nor U11780 (N_11780,N_8034,N_9170);
and U11781 (N_11781,N_9261,N_9094);
nor U11782 (N_11782,N_8249,N_8957);
nand U11783 (N_11783,N_9661,N_8717);
nand U11784 (N_11784,N_8831,N_9272);
and U11785 (N_11785,N_7723,N_9674);
or U11786 (N_11786,N_8597,N_9907);
and U11787 (N_11787,N_9322,N_8067);
nand U11788 (N_11788,N_8757,N_7974);
nand U11789 (N_11789,N_9995,N_7761);
and U11790 (N_11790,N_7838,N_9821);
nor U11791 (N_11791,N_7778,N_9975);
nand U11792 (N_11792,N_8666,N_7729);
nand U11793 (N_11793,N_9639,N_8760);
nor U11794 (N_11794,N_8749,N_9557);
xnor U11795 (N_11795,N_8374,N_8399);
or U11796 (N_11796,N_8344,N_9144);
or U11797 (N_11797,N_9721,N_8458);
nand U11798 (N_11798,N_9314,N_9352);
or U11799 (N_11799,N_8653,N_7583);
nand U11800 (N_11800,N_9255,N_7895);
nor U11801 (N_11801,N_8802,N_9041);
nand U11802 (N_11802,N_8076,N_9178);
nand U11803 (N_11803,N_8301,N_9249);
nor U11804 (N_11804,N_9227,N_9893);
nor U11805 (N_11805,N_7712,N_8056);
and U11806 (N_11806,N_9662,N_9775);
nor U11807 (N_11807,N_8385,N_9743);
and U11808 (N_11808,N_9558,N_9102);
nor U11809 (N_11809,N_8783,N_9407);
nor U11810 (N_11810,N_9543,N_9063);
nor U11811 (N_11811,N_9234,N_7538);
nor U11812 (N_11812,N_9410,N_7697);
nand U11813 (N_11813,N_8902,N_8251);
nand U11814 (N_11814,N_9387,N_7523);
nand U11815 (N_11815,N_7618,N_9585);
xnor U11816 (N_11816,N_9741,N_8900);
or U11817 (N_11817,N_9096,N_9574);
or U11818 (N_11818,N_7723,N_8742);
and U11819 (N_11819,N_8856,N_8266);
nor U11820 (N_11820,N_8175,N_8833);
xnor U11821 (N_11821,N_9811,N_8231);
xor U11822 (N_11822,N_7752,N_8231);
xnor U11823 (N_11823,N_8330,N_8029);
and U11824 (N_11824,N_7958,N_8556);
nor U11825 (N_11825,N_9235,N_8669);
or U11826 (N_11826,N_8631,N_9348);
nand U11827 (N_11827,N_8411,N_8341);
nand U11828 (N_11828,N_8645,N_9778);
and U11829 (N_11829,N_8856,N_7711);
nand U11830 (N_11830,N_8502,N_9545);
or U11831 (N_11831,N_7709,N_8511);
and U11832 (N_11832,N_9742,N_8443);
or U11833 (N_11833,N_9272,N_9536);
nand U11834 (N_11834,N_9537,N_8140);
and U11835 (N_11835,N_7920,N_8017);
nand U11836 (N_11836,N_8408,N_9245);
nand U11837 (N_11837,N_9744,N_7953);
and U11838 (N_11838,N_8787,N_8687);
nor U11839 (N_11839,N_7748,N_8036);
nand U11840 (N_11840,N_7964,N_9343);
and U11841 (N_11841,N_8117,N_9112);
nand U11842 (N_11842,N_7659,N_9680);
nor U11843 (N_11843,N_8420,N_8068);
and U11844 (N_11844,N_9221,N_8666);
nand U11845 (N_11845,N_7564,N_7806);
nand U11846 (N_11846,N_9880,N_8930);
nand U11847 (N_11847,N_9548,N_9386);
nor U11848 (N_11848,N_8228,N_8203);
nand U11849 (N_11849,N_8320,N_8291);
nand U11850 (N_11850,N_9045,N_9204);
nor U11851 (N_11851,N_8356,N_8090);
and U11852 (N_11852,N_8081,N_9807);
nand U11853 (N_11853,N_7759,N_8058);
and U11854 (N_11854,N_8550,N_7733);
nor U11855 (N_11855,N_9038,N_9087);
xnor U11856 (N_11856,N_7842,N_8009);
nor U11857 (N_11857,N_9293,N_8121);
nor U11858 (N_11858,N_9982,N_8482);
nor U11859 (N_11859,N_9447,N_7778);
nor U11860 (N_11860,N_9167,N_7723);
nand U11861 (N_11861,N_9013,N_7530);
or U11862 (N_11862,N_9061,N_9126);
nand U11863 (N_11863,N_8549,N_9221);
or U11864 (N_11864,N_9871,N_9325);
nor U11865 (N_11865,N_7546,N_8936);
or U11866 (N_11866,N_9508,N_8478);
and U11867 (N_11867,N_8503,N_9548);
xnor U11868 (N_11868,N_8444,N_8344);
nand U11869 (N_11869,N_9644,N_8452);
or U11870 (N_11870,N_8575,N_7877);
nand U11871 (N_11871,N_9364,N_8787);
and U11872 (N_11872,N_8694,N_8830);
nor U11873 (N_11873,N_7653,N_8892);
or U11874 (N_11874,N_9165,N_9402);
xnor U11875 (N_11875,N_9733,N_9664);
and U11876 (N_11876,N_8245,N_8828);
nor U11877 (N_11877,N_9100,N_9892);
nor U11878 (N_11878,N_8756,N_9219);
or U11879 (N_11879,N_9847,N_8581);
nor U11880 (N_11880,N_9921,N_8292);
nor U11881 (N_11881,N_9276,N_9170);
nand U11882 (N_11882,N_9098,N_8986);
and U11883 (N_11883,N_8515,N_7587);
or U11884 (N_11884,N_8870,N_8064);
or U11885 (N_11885,N_8839,N_8340);
nor U11886 (N_11886,N_8683,N_7721);
nor U11887 (N_11887,N_9049,N_8684);
nand U11888 (N_11888,N_7975,N_7621);
nor U11889 (N_11889,N_9821,N_8196);
nand U11890 (N_11890,N_7759,N_8596);
and U11891 (N_11891,N_8486,N_9848);
nor U11892 (N_11892,N_8442,N_9389);
or U11893 (N_11893,N_9381,N_9588);
nor U11894 (N_11894,N_9261,N_9116);
nand U11895 (N_11895,N_9638,N_9913);
or U11896 (N_11896,N_7867,N_8522);
xor U11897 (N_11897,N_8828,N_9126);
or U11898 (N_11898,N_9330,N_9614);
and U11899 (N_11899,N_7951,N_8557);
nor U11900 (N_11900,N_8274,N_8101);
or U11901 (N_11901,N_8278,N_9084);
xor U11902 (N_11902,N_9341,N_8432);
and U11903 (N_11903,N_8945,N_8126);
xor U11904 (N_11904,N_9364,N_8736);
and U11905 (N_11905,N_9718,N_9882);
or U11906 (N_11906,N_9088,N_8548);
and U11907 (N_11907,N_9688,N_9586);
nor U11908 (N_11908,N_8994,N_9497);
or U11909 (N_11909,N_8394,N_8839);
xnor U11910 (N_11910,N_9180,N_8658);
and U11911 (N_11911,N_8150,N_7682);
or U11912 (N_11912,N_8107,N_9049);
xor U11913 (N_11913,N_9292,N_9130);
nand U11914 (N_11914,N_8775,N_9560);
nand U11915 (N_11915,N_7519,N_9238);
nand U11916 (N_11916,N_9655,N_9191);
nand U11917 (N_11917,N_9133,N_8347);
and U11918 (N_11918,N_9903,N_9756);
nand U11919 (N_11919,N_8285,N_9435);
or U11920 (N_11920,N_7590,N_9454);
xor U11921 (N_11921,N_9340,N_9437);
nor U11922 (N_11922,N_8576,N_9825);
nand U11923 (N_11923,N_8206,N_7770);
nand U11924 (N_11924,N_8168,N_8852);
or U11925 (N_11925,N_9310,N_8536);
nor U11926 (N_11926,N_9751,N_9821);
nor U11927 (N_11927,N_9503,N_7744);
nor U11928 (N_11928,N_9693,N_9442);
and U11929 (N_11929,N_9558,N_9881);
nor U11930 (N_11930,N_7623,N_8839);
nand U11931 (N_11931,N_8083,N_7574);
nand U11932 (N_11932,N_8803,N_8777);
nor U11933 (N_11933,N_9210,N_9314);
nand U11934 (N_11934,N_8984,N_9548);
nand U11935 (N_11935,N_7752,N_8765);
xnor U11936 (N_11936,N_9330,N_9528);
and U11937 (N_11937,N_9275,N_8614);
or U11938 (N_11938,N_7875,N_8003);
nor U11939 (N_11939,N_9606,N_8551);
or U11940 (N_11940,N_8866,N_9037);
xnor U11941 (N_11941,N_8468,N_7804);
or U11942 (N_11942,N_9887,N_8974);
nand U11943 (N_11943,N_9146,N_7756);
or U11944 (N_11944,N_9233,N_8097);
nor U11945 (N_11945,N_9234,N_8705);
and U11946 (N_11946,N_8596,N_9271);
or U11947 (N_11947,N_8926,N_9868);
or U11948 (N_11948,N_7729,N_8028);
nor U11949 (N_11949,N_8776,N_8023);
nor U11950 (N_11950,N_8933,N_9113);
and U11951 (N_11951,N_8764,N_9394);
and U11952 (N_11952,N_7651,N_8371);
or U11953 (N_11953,N_8040,N_8220);
and U11954 (N_11954,N_8830,N_9442);
and U11955 (N_11955,N_7854,N_8865);
nand U11956 (N_11956,N_8245,N_8646);
nor U11957 (N_11957,N_8913,N_8880);
and U11958 (N_11958,N_8618,N_8499);
or U11959 (N_11959,N_8743,N_9475);
xnor U11960 (N_11960,N_9636,N_8253);
nor U11961 (N_11961,N_8820,N_9599);
nor U11962 (N_11962,N_9841,N_9289);
and U11963 (N_11963,N_9920,N_8918);
and U11964 (N_11964,N_8177,N_8067);
nand U11965 (N_11965,N_8107,N_8058);
nand U11966 (N_11966,N_8364,N_9055);
nor U11967 (N_11967,N_8179,N_9347);
or U11968 (N_11968,N_8063,N_7909);
nand U11969 (N_11969,N_8904,N_7729);
nor U11970 (N_11970,N_9643,N_8437);
and U11971 (N_11971,N_9587,N_8868);
nor U11972 (N_11972,N_8406,N_8765);
and U11973 (N_11973,N_9587,N_7651);
or U11974 (N_11974,N_9769,N_8011);
or U11975 (N_11975,N_9990,N_7813);
nor U11976 (N_11976,N_9625,N_9991);
nor U11977 (N_11977,N_7673,N_8681);
nand U11978 (N_11978,N_9969,N_9270);
and U11979 (N_11979,N_9397,N_9644);
nand U11980 (N_11980,N_8042,N_8459);
or U11981 (N_11981,N_9577,N_9328);
or U11982 (N_11982,N_8641,N_9756);
nor U11983 (N_11983,N_8332,N_8935);
and U11984 (N_11984,N_7609,N_9095);
nand U11985 (N_11985,N_9022,N_8730);
and U11986 (N_11986,N_8592,N_9504);
xor U11987 (N_11987,N_9270,N_8454);
and U11988 (N_11988,N_8822,N_9767);
nor U11989 (N_11989,N_8885,N_8486);
and U11990 (N_11990,N_9290,N_8583);
or U11991 (N_11991,N_8691,N_9208);
or U11992 (N_11992,N_8704,N_7540);
or U11993 (N_11993,N_9775,N_9168);
or U11994 (N_11994,N_7652,N_8568);
or U11995 (N_11995,N_9612,N_7816);
nand U11996 (N_11996,N_8812,N_9899);
and U11997 (N_11997,N_7519,N_8816);
nand U11998 (N_11998,N_8078,N_8779);
nor U11999 (N_11999,N_9492,N_9223);
nor U12000 (N_12000,N_7790,N_7606);
nor U12001 (N_12001,N_7553,N_8395);
or U12002 (N_12002,N_9154,N_8138);
xnor U12003 (N_12003,N_9708,N_8518);
nand U12004 (N_12004,N_8150,N_8791);
nand U12005 (N_12005,N_9117,N_7977);
and U12006 (N_12006,N_9888,N_9243);
nand U12007 (N_12007,N_8343,N_8104);
nor U12008 (N_12008,N_8857,N_9201);
or U12009 (N_12009,N_9612,N_9663);
nor U12010 (N_12010,N_8221,N_9684);
and U12011 (N_12011,N_8860,N_7902);
nand U12012 (N_12012,N_7913,N_8569);
or U12013 (N_12013,N_9733,N_8145);
nor U12014 (N_12014,N_8579,N_7990);
or U12015 (N_12015,N_9999,N_9321);
and U12016 (N_12016,N_8170,N_7838);
nor U12017 (N_12017,N_9821,N_9461);
and U12018 (N_12018,N_9133,N_9894);
xnor U12019 (N_12019,N_8824,N_7870);
or U12020 (N_12020,N_8377,N_9437);
nand U12021 (N_12021,N_9565,N_9603);
nor U12022 (N_12022,N_8242,N_8878);
nand U12023 (N_12023,N_9138,N_9401);
nand U12024 (N_12024,N_8184,N_8115);
xor U12025 (N_12025,N_7705,N_7691);
and U12026 (N_12026,N_8956,N_9575);
nor U12027 (N_12027,N_7783,N_7973);
nor U12028 (N_12028,N_8256,N_9512);
or U12029 (N_12029,N_9073,N_8035);
nand U12030 (N_12030,N_7939,N_9408);
nor U12031 (N_12031,N_8728,N_9588);
or U12032 (N_12032,N_8916,N_9700);
and U12033 (N_12033,N_8634,N_8242);
or U12034 (N_12034,N_9065,N_7828);
xor U12035 (N_12035,N_9639,N_7548);
nor U12036 (N_12036,N_9613,N_9800);
and U12037 (N_12037,N_7965,N_8044);
nor U12038 (N_12038,N_9886,N_8013);
nor U12039 (N_12039,N_9665,N_8756);
nand U12040 (N_12040,N_9679,N_8186);
nor U12041 (N_12041,N_8906,N_7588);
xor U12042 (N_12042,N_8638,N_8533);
nand U12043 (N_12043,N_8367,N_7922);
and U12044 (N_12044,N_9435,N_7570);
and U12045 (N_12045,N_8695,N_9976);
and U12046 (N_12046,N_8960,N_9173);
nand U12047 (N_12047,N_9255,N_7925);
nor U12048 (N_12048,N_9067,N_7913);
nand U12049 (N_12049,N_8195,N_7538);
nor U12050 (N_12050,N_8358,N_8167);
nand U12051 (N_12051,N_9375,N_8343);
and U12052 (N_12052,N_8175,N_7741);
and U12053 (N_12053,N_8275,N_9844);
or U12054 (N_12054,N_9737,N_8051);
nor U12055 (N_12055,N_9692,N_8866);
or U12056 (N_12056,N_8353,N_9709);
and U12057 (N_12057,N_9239,N_9268);
nand U12058 (N_12058,N_7723,N_7516);
and U12059 (N_12059,N_8664,N_8966);
nand U12060 (N_12060,N_7863,N_9608);
nand U12061 (N_12061,N_8956,N_9115);
nor U12062 (N_12062,N_7720,N_8088);
and U12063 (N_12063,N_8961,N_9763);
nor U12064 (N_12064,N_8611,N_7757);
nand U12065 (N_12065,N_9813,N_9084);
nand U12066 (N_12066,N_8708,N_7609);
nor U12067 (N_12067,N_8277,N_9026);
nand U12068 (N_12068,N_9512,N_8709);
and U12069 (N_12069,N_8502,N_9112);
and U12070 (N_12070,N_8300,N_9114);
nand U12071 (N_12071,N_8930,N_9201);
nor U12072 (N_12072,N_9760,N_8960);
or U12073 (N_12073,N_7796,N_8722);
nor U12074 (N_12074,N_8032,N_9133);
or U12075 (N_12075,N_8441,N_8074);
and U12076 (N_12076,N_7868,N_8618);
xnor U12077 (N_12077,N_9529,N_8707);
and U12078 (N_12078,N_9190,N_9482);
nand U12079 (N_12079,N_8961,N_7586);
nand U12080 (N_12080,N_9676,N_9644);
or U12081 (N_12081,N_9478,N_9583);
nand U12082 (N_12082,N_9886,N_7574);
nor U12083 (N_12083,N_9101,N_8694);
and U12084 (N_12084,N_8386,N_9261);
nand U12085 (N_12085,N_9455,N_8138);
nor U12086 (N_12086,N_9884,N_9356);
or U12087 (N_12087,N_7976,N_7622);
and U12088 (N_12088,N_9181,N_8231);
nor U12089 (N_12089,N_8257,N_9028);
nor U12090 (N_12090,N_8996,N_7728);
nor U12091 (N_12091,N_9541,N_7817);
and U12092 (N_12092,N_9827,N_9301);
or U12093 (N_12093,N_8418,N_9877);
and U12094 (N_12094,N_7611,N_8104);
nor U12095 (N_12095,N_9378,N_7690);
and U12096 (N_12096,N_9896,N_8941);
nor U12097 (N_12097,N_7733,N_8249);
or U12098 (N_12098,N_7714,N_8968);
nand U12099 (N_12099,N_7858,N_9410);
nor U12100 (N_12100,N_9926,N_8866);
nand U12101 (N_12101,N_7546,N_8054);
and U12102 (N_12102,N_9837,N_9638);
and U12103 (N_12103,N_8642,N_8937);
nor U12104 (N_12104,N_9653,N_7555);
or U12105 (N_12105,N_9676,N_9966);
xor U12106 (N_12106,N_9515,N_9276);
nor U12107 (N_12107,N_8774,N_8646);
nand U12108 (N_12108,N_7797,N_9406);
and U12109 (N_12109,N_8649,N_8442);
nand U12110 (N_12110,N_9060,N_8075);
nor U12111 (N_12111,N_7862,N_8189);
or U12112 (N_12112,N_8988,N_7772);
nor U12113 (N_12113,N_7981,N_7565);
or U12114 (N_12114,N_7841,N_7809);
or U12115 (N_12115,N_8637,N_7868);
nor U12116 (N_12116,N_9506,N_8143);
and U12117 (N_12117,N_9960,N_9873);
nor U12118 (N_12118,N_8284,N_8134);
or U12119 (N_12119,N_8982,N_9020);
or U12120 (N_12120,N_8775,N_8599);
nand U12121 (N_12121,N_8253,N_7624);
nor U12122 (N_12122,N_8044,N_9715);
nor U12123 (N_12123,N_7795,N_9872);
nor U12124 (N_12124,N_8488,N_9854);
xnor U12125 (N_12125,N_8632,N_8378);
nand U12126 (N_12126,N_9387,N_9778);
or U12127 (N_12127,N_7658,N_8978);
or U12128 (N_12128,N_7707,N_8347);
xor U12129 (N_12129,N_7504,N_9786);
nand U12130 (N_12130,N_7682,N_7826);
and U12131 (N_12131,N_8842,N_8241);
nor U12132 (N_12132,N_9705,N_8374);
nor U12133 (N_12133,N_8834,N_9074);
nor U12134 (N_12134,N_7781,N_8463);
nor U12135 (N_12135,N_9407,N_7777);
and U12136 (N_12136,N_9194,N_8942);
or U12137 (N_12137,N_9079,N_9779);
nor U12138 (N_12138,N_8149,N_8430);
and U12139 (N_12139,N_9142,N_8716);
nand U12140 (N_12140,N_8361,N_8136);
or U12141 (N_12141,N_9154,N_9671);
or U12142 (N_12142,N_9827,N_8805);
nand U12143 (N_12143,N_9980,N_9027);
xor U12144 (N_12144,N_7898,N_7723);
nand U12145 (N_12145,N_8546,N_7985);
nand U12146 (N_12146,N_9987,N_9918);
and U12147 (N_12147,N_7903,N_7739);
nor U12148 (N_12148,N_7946,N_8183);
nor U12149 (N_12149,N_9952,N_8403);
nor U12150 (N_12150,N_8508,N_7740);
or U12151 (N_12151,N_9330,N_8222);
xnor U12152 (N_12152,N_8234,N_9120);
and U12153 (N_12153,N_9906,N_9264);
and U12154 (N_12154,N_9578,N_8958);
and U12155 (N_12155,N_8004,N_8232);
and U12156 (N_12156,N_8079,N_7963);
and U12157 (N_12157,N_9313,N_7983);
nor U12158 (N_12158,N_8656,N_9071);
nand U12159 (N_12159,N_7983,N_9006);
nor U12160 (N_12160,N_9130,N_7503);
and U12161 (N_12161,N_8122,N_8594);
nor U12162 (N_12162,N_7793,N_8198);
nand U12163 (N_12163,N_8128,N_8472);
xor U12164 (N_12164,N_9380,N_8991);
xor U12165 (N_12165,N_9124,N_7541);
nor U12166 (N_12166,N_7975,N_9835);
nor U12167 (N_12167,N_8481,N_9793);
xor U12168 (N_12168,N_7651,N_9226);
and U12169 (N_12169,N_9074,N_9199);
nor U12170 (N_12170,N_7536,N_8980);
nor U12171 (N_12171,N_7559,N_7922);
or U12172 (N_12172,N_8337,N_8577);
or U12173 (N_12173,N_9718,N_9654);
nor U12174 (N_12174,N_8733,N_8096);
or U12175 (N_12175,N_7545,N_8839);
and U12176 (N_12176,N_9088,N_9490);
nor U12177 (N_12177,N_7679,N_9205);
xnor U12178 (N_12178,N_7681,N_8908);
nor U12179 (N_12179,N_7742,N_7815);
nor U12180 (N_12180,N_7983,N_9490);
nand U12181 (N_12181,N_8607,N_8593);
nor U12182 (N_12182,N_9941,N_7796);
or U12183 (N_12183,N_9437,N_8783);
or U12184 (N_12184,N_9999,N_9804);
nor U12185 (N_12185,N_8738,N_9743);
and U12186 (N_12186,N_9949,N_9434);
nand U12187 (N_12187,N_8778,N_8032);
nor U12188 (N_12188,N_7644,N_9087);
or U12189 (N_12189,N_9863,N_9699);
or U12190 (N_12190,N_9872,N_9129);
or U12191 (N_12191,N_9052,N_8923);
nor U12192 (N_12192,N_9620,N_7771);
xor U12193 (N_12193,N_7839,N_9579);
nand U12194 (N_12194,N_9360,N_8120);
nor U12195 (N_12195,N_8444,N_8111);
or U12196 (N_12196,N_9367,N_7569);
and U12197 (N_12197,N_9132,N_7714);
xor U12198 (N_12198,N_7660,N_7685);
nand U12199 (N_12199,N_9815,N_9381);
nor U12200 (N_12200,N_7902,N_8546);
nor U12201 (N_12201,N_9514,N_8655);
or U12202 (N_12202,N_7771,N_8140);
nor U12203 (N_12203,N_8910,N_8810);
and U12204 (N_12204,N_7544,N_8131);
nand U12205 (N_12205,N_7693,N_7728);
and U12206 (N_12206,N_9028,N_7897);
nor U12207 (N_12207,N_9213,N_9621);
or U12208 (N_12208,N_8914,N_8792);
or U12209 (N_12209,N_7826,N_9955);
and U12210 (N_12210,N_8435,N_7589);
nand U12211 (N_12211,N_8200,N_7901);
xnor U12212 (N_12212,N_9918,N_8529);
or U12213 (N_12213,N_9339,N_7979);
nand U12214 (N_12214,N_8230,N_9896);
xor U12215 (N_12215,N_9056,N_9292);
nor U12216 (N_12216,N_9748,N_8621);
or U12217 (N_12217,N_8003,N_8804);
or U12218 (N_12218,N_9853,N_9418);
or U12219 (N_12219,N_9761,N_9952);
nor U12220 (N_12220,N_7820,N_7962);
or U12221 (N_12221,N_7718,N_8249);
nor U12222 (N_12222,N_7761,N_9778);
and U12223 (N_12223,N_8641,N_9521);
nand U12224 (N_12224,N_8795,N_8540);
nand U12225 (N_12225,N_9872,N_9825);
and U12226 (N_12226,N_9351,N_7522);
xnor U12227 (N_12227,N_8257,N_9331);
nor U12228 (N_12228,N_9197,N_9717);
and U12229 (N_12229,N_8373,N_9106);
xor U12230 (N_12230,N_7585,N_9736);
nor U12231 (N_12231,N_9887,N_8284);
xnor U12232 (N_12232,N_9915,N_8212);
and U12233 (N_12233,N_9727,N_7956);
or U12234 (N_12234,N_9511,N_7651);
and U12235 (N_12235,N_8387,N_9353);
or U12236 (N_12236,N_9077,N_8064);
nor U12237 (N_12237,N_9743,N_8344);
nor U12238 (N_12238,N_9061,N_9720);
or U12239 (N_12239,N_8529,N_8763);
nand U12240 (N_12240,N_8577,N_9093);
and U12241 (N_12241,N_9203,N_7883);
nor U12242 (N_12242,N_9193,N_9119);
nor U12243 (N_12243,N_7880,N_7711);
and U12244 (N_12244,N_9985,N_7731);
and U12245 (N_12245,N_9099,N_7661);
and U12246 (N_12246,N_7579,N_9341);
or U12247 (N_12247,N_8544,N_8146);
and U12248 (N_12248,N_8963,N_8225);
nand U12249 (N_12249,N_9680,N_9449);
and U12250 (N_12250,N_9500,N_7613);
and U12251 (N_12251,N_9007,N_9603);
or U12252 (N_12252,N_9376,N_8377);
and U12253 (N_12253,N_9102,N_9074);
nor U12254 (N_12254,N_9581,N_8522);
nand U12255 (N_12255,N_8659,N_8838);
nand U12256 (N_12256,N_8445,N_9102);
nand U12257 (N_12257,N_8795,N_7562);
nand U12258 (N_12258,N_8818,N_8261);
nand U12259 (N_12259,N_8003,N_8393);
and U12260 (N_12260,N_9172,N_8770);
and U12261 (N_12261,N_9722,N_8861);
nand U12262 (N_12262,N_9679,N_9601);
or U12263 (N_12263,N_9798,N_8730);
nor U12264 (N_12264,N_9144,N_7724);
and U12265 (N_12265,N_8242,N_8554);
nand U12266 (N_12266,N_9317,N_8723);
nand U12267 (N_12267,N_8465,N_8973);
and U12268 (N_12268,N_9769,N_8855);
nor U12269 (N_12269,N_8909,N_9574);
and U12270 (N_12270,N_9750,N_9012);
and U12271 (N_12271,N_9406,N_7509);
or U12272 (N_12272,N_8014,N_7930);
and U12273 (N_12273,N_8661,N_7541);
or U12274 (N_12274,N_8329,N_9409);
nor U12275 (N_12275,N_9995,N_9481);
nor U12276 (N_12276,N_8552,N_9368);
or U12277 (N_12277,N_7637,N_8016);
or U12278 (N_12278,N_8815,N_8388);
nand U12279 (N_12279,N_7513,N_9150);
or U12280 (N_12280,N_9273,N_8210);
xnor U12281 (N_12281,N_9790,N_7949);
and U12282 (N_12282,N_8528,N_8971);
nand U12283 (N_12283,N_9715,N_9325);
nand U12284 (N_12284,N_8670,N_8453);
and U12285 (N_12285,N_9997,N_9836);
xor U12286 (N_12286,N_7766,N_9700);
or U12287 (N_12287,N_9762,N_7551);
nand U12288 (N_12288,N_8224,N_9288);
or U12289 (N_12289,N_8986,N_7813);
nand U12290 (N_12290,N_7591,N_7754);
nand U12291 (N_12291,N_9036,N_9641);
and U12292 (N_12292,N_7941,N_9211);
nor U12293 (N_12293,N_9443,N_8306);
xor U12294 (N_12294,N_7534,N_9119);
or U12295 (N_12295,N_8636,N_9272);
nand U12296 (N_12296,N_7719,N_9643);
nor U12297 (N_12297,N_9485,N_7616);
nand U12298 (N_12298,N_9820,N_9282);
and U12299 (N_12299,N_8088,N_9645);
nor U12300 (N_12300,N_9803,N_8285);
or U12301 (N_12301,N_7895,N_9891);
xnor U12302 (N_12302,N_7906,N_9867);
nor U12303 (N_12303,N_8326,N_7889);
nand U12304 (N_12304,N_8179,N_8205);
nor U12305 (N_12305,N_8346,N_9992);
nor U12306 (N_12306,N_8131,N_8013);
xor U12307 (N_12307,N_7670,N_9634);
xor U12308 (N_12308,N_9824,N_8115);
nor U12309 (N_12309,N_9359,N_8621);
nand U12310 (N_12310,N_7728,N_9238);
and U12311 (N_12311,N_7811,N_7654);
nand U12312 (N_12312,N_9865,N_7804);
nand U12313 (N_12313,N_9737,N_8029);
or U12314 (N_12314,N_9627,N_7725);
and U12315 (N_12315,N_9544,N_8501);
nand U12316 (N_12316,N_7674,N_9656);
and U12317 (N_12317,N_9571,N_7674);
nor U12318 (N_12318,N_7858,N_8656);
or U12319 (N_12319,N_7604,N_8329);
or U12320 (N_12320,N_9322,N_7830);
and U12321 (N_12321,N_9719,N_9567);
or U12322 (N_12322,N_8567,N_9031);
or U12323 (N_12323,N_8103,N_7906);
nand U12324 (N_12324,N_7761,N_9574);
nand U12325 (N_12325,N_7728,N_8185);
nand U12326 (N_12326,N_9997,N_8234);
and U12327 (N_12327,N_7878,N_8586);
and U12328 (N_12328,N_7660,N_8389);
xor U12329 (N_12329,N_8020,N_8939);
nand U12330 (N_12330,N_9737,N_9872);
nor U12331 (N_12331,N_9868,N_9481);
nor U12332 (N_12332,N_8120,N_9819);
or U12333 (N_12333,N_8349,N_9367);
xnor U12334 (N_12334,N_8280,N_9829);
and U12335 (N_12335,N_9328,N_7685);
and U12336 (N_12336,N_7627,N_8219);
nand U12337 (N_12337,N_9629,N_8561);
nand U12338 (N_12338,N_7871,N_9541);
nand U12339 (N_12339,N_7567,N_9336);
or U12340 (N_12340,N_9175,N_9876);
nand U12341 (N_12341,N_9064,N_9192);
or U12342 (N_12342,N_9014,N_9973);
nor U12343 (N_12343,N_8839,N_8955);
nand U12344 (N_12344,N_9174,N_9514);
or U12345 (N_12345,N_9558,N_8596);
or U12346 (N_12346,N_9905,N_8121);
nor U12347 (N_12347,N_7778,N_7857);
xnor U12348 (N_12348,N_8753,N_9400);
xor U12349 (N_12349,N_7669,N_9782);
nor U12350 (N_12350,N_9930,N_9902);
nor U12351 (N_12351,N_7520,N_7913);
or U12352 (N_12352,N_7787,N_9024);
and U12353 (N_12353,N_7683,N_7764);
and U12354 (N_12354,N_9197,N_9863);
nand U12355 (N_12355,N_9359,N_8464);
and U12356 (N_12356,N_8444,N_9161);
or U12357 (N_12357,N_8975,N_8501);
or U12358 (N_12358,N_8760,N_9731);
nor U12359 (N_12359,N_9845,N_7567);
nor U12360 (N_12360,N_9800,N_7728);
nand U12361 (N_12361,N_9997,N_9512);
or U12362 (N_12362,N_7531,N_8534);
xnor U12363 (N_12363,N_9875,N_8007);
and U12364 (N_12364,N_8321,N_9661);
xor U12365 (N_12365,N_8535,N_8037);
and U12366 (N_12366,N_8936,N_8217);
nor U12367 (N_12367,N_8963,N_7847);
nand U12368 (N_12368,N_9730,N_9164);
xnor U12369 (N_12369,N_9924,N_7796);
or U12370 (N_12370,N_8507,N_8487);
and U12371 (N_12371,N_7552,N_8813);
and U12372 (N_12372,N_9256,N_9014);
xor U12373 (N_12373,N_9784,N_8523);
nor U12374 (N_12374,N_7997,N_9283);
xor U12375 (N_12375,N_7745,N_9153);
and U12376 (N_12376,N_9040,N_9574);
or U12377 (N_12377,N_9406,N_9686);
or U12378 (N_12378,N_7928,N_9071);
xnor U12379 (N_12379,N_8757,N_8689);
xnor U12380 (N_12380,N_7980,N_9237);
nand U12381 (N_12381,N_8151,N_7672);
or U12382 (N_12382,N_7735,N_8605);
nor U12383 (N_12383,N_7503,N_9310);
or U12384 (N_12384,N_8468,N_9094);
and U12385 (N_12385,N_9329,N_9775);
xor U12386 (N_12386,N_8005,N_9450);
nand U12387 (N_12387,N_8643,N_8414);
or U12388 (N_12388,N_7626,N_9783);
and U12389 (N_12389,N_9586,N_9034);
and U12390 (N_12390,N_8078,N_8365);
nand U12391 (N_12391,N_8424,N_9655);
and U12392 (N_12392,N_9107,N_9242);
and U12393 (N_12393,N_9870,N_9938);
nor U12394 (N_12394,N_9612,N_8013);
nand U12395 (N_12395,N_8449,N_9735);
and U12396 (N_12396,N_8781,N_9749);
and U12397 (N_12397,N_9294,N_8543);
nand U12398 (N_12398,N_9121,N_9594);
or U12399 (N_12399,N_8597,N_8073);
or U12400 (N_12400,N_8871,N_9341);
or U12401 (N_12401,N_7938,N_8161);
nand U12402 (N_12402,N_9187,N_7771);
or U12403 (N_12403,N_9395,N_7913);
nand U12404 (N_12404,N_8798,N_9805);
or U12405 (N_12405,N_8067,N_7669);
or U12406 (N_12406,N_9711,N_7968);
nand U12407 (N_12407,N_7840,N_8411);
and U12408 (N_12408,N_8648,N_8498);
nor U12409 (N_12409,N_9609,N_9439);
or U12410 (N_12410,N_8699,N_9680);
nand U12411 (N_12411,N_9537,N_8009);
nand U12412 (N_12412,N_7918,N_9667);
nor U12413 (N_12413,N_9482,N_7940);
xnor U12414 (N_12414,N_9558,N_9442);
nor U12415 (N_12415,N_8788,N_9641);
or U12416 (N_12416,N_9101,N_9457);
or U12417 (N_12417,N_8115,N_8226);
nand U12418 (N_12418,N_9236,N_8140);
or U12419 (N_12419,N_9172,N_8573);
or U12420 (N_12420,N_7618,N_9671);
nand U12421 (N_12421,N_7550,N_8657);
and U12422 (N_12422,N_8489,N_7698);
nor U12423 (N_12423,N_8305,N_9992);
nor U12424 (N_12424,N_8332,N_8997);
or U12425 (N_12425,N_9794,N_8982);
or U12426 (N_12426,N_8886,N_7557);
nand U12427 (N_12427,N_9144,N_9036);
or U12428 (N_12428,N_9548,N_9219);
nand U12429 (N_12429,N_7962,N_7796);
and U12430 (N_12430,N_9755,N_8838);
nand U12431 (N_12431,N_9492,N_9692);
xnor U12432 (N_12432,N_7661,N_9264);
or U12433 (N_12433,N_9031,N_9616);
nand U12434 (N_12434,N_9204,N_7994);
and U12435 (N_12435,N_9325,N_9191);
xnor U12436 (N_12436,N_7971,N_8450);
nor U12437 (N_12437,N_9275,N_7860);
and U12438 (N_12438,N_9673,N_9079);
or U12439 (N_12439,N_8263,N_9183);
nand U12440 (N_12440,N_9988,N_9990);
or U12441 (N_12441,N_8349,N_8127);
and U12442 (N_12442,N_8653,N_8834);
xnor U12443 (N_12443,N_7921,N_7872);
or U12444 (N_12444,N_9804,N_8479);
nor U12445 (N_12445,N_9596,N_8475);
and U12446 (N_12446,N_9342,N_7532);
xnor U12447 (N_12447,N_8620,N_8256);
or U12448 (N_12448,N_8026,N_8209);
xnor U12449 (N_12449,N_9049,N_8697);
or U12450 (N_12450,N_9229,N_9746);
or U12451 (N_12451,N_8581,N_9397);
nor U12452 (N_12452,N_8739,N_8743);
nor U12453 (N_12453,N_9777,N_9020);
or U12454 (N_12454,N_9408,N_8945);
and U12455 (N_12455,N_9661,N_9155);
nand U12456 (N_12456,N_9528,N_9649);
or U12457 (N_12457,N_8715,N_8924);
nand U12458 (N_12458,N_8915,N_8572);
and U12459 (N_12459,N_9802,N_9820);
nand U12460 (N_12460,N_7897,N_8548);
nor U12461 (N_12461,N_7887,N_7553);
xnor U12462 (N_12462,N_7846,N_8596);
nand U12463 (N_12463,N_9294,N_9185);
nand U12464 (N_12464,N_8079,N_9264);
or U12465 (N_12465,N_8574,N_8279);
and U12466 (N_12466,N_8651,N_9187);
or U12467 (N_12467,N_7737,N_9733);
or U12468 (N_12468,N_8794,N_7878);
and U12469 (N_12469,N_8560,N_9867);
or U12470 (N_12470,N_9488,N_8655);
and U12471 (N_12471,N_8682,N_8958);
nor U12472 (N_12472,N_9271,N_9718);
or U12473 (N_12473,N_9371,N_9476);
nor U12474 (N_12474,N_8926,N_8565);
or U12475 (N_12475,N_8676,N_8517);
nor U12476 (N_12476,N_8840,N_8657);
nor U12477 (N_12477,N_9697,N_9155);
nand U12478 (N_12478,N_9235,N_8500);
nand U12479 (N_12479,N_7897,N_8519);
and U12480 (N_12480,N_9460,N_7948);
and U12481 (N_12481,N_9627,N_8780);
and U12482 (N_12482,N_8210,N_9595);
or U12483 (N_12483,N_9927,N_7707);
nor U12484 (N_12484,N_9728,N_9508);
xor U12485 (N_12485,N_9283,N_9282);
nor U12486 (N_12486,N_7624,N_7975);
and U12487 (N_12487,N_7646,N_7613);
and U12488 (N_12488,N_9484,N_9349);
nor U12489 (N_12489,N_9884,N_8935);
or U12490 (N_12490,N_8034,N_9605);
nor U12491 (N_12491,N_8750,N_8622);
xor U12492 (N_12492,N_8195,N_9941);
nand U12493 (N_12493,N_8545,N_7651);
nor U12494 (N_12494,N_7997,N_7624);
xor U12495 (N_12495,N_9470,N_7957);
nor U12496 (N_12496,N_9440,N_7944);
nor U12497 (N_12497,N_8085,N_8141);
nor U12498 (N_12498,N_9896,N_7572);
nand U12499 (N_12499,N_8453,N_8970);
or U12500 (N_12500,N_10879,N_11431);
nand U12501 (N_12501,N_11512,N_11907);
nand U12502 (N_12502,N_10079,N_10954);
nor U12503 (N_12503,N_10063,N_10558);
or U12504 (N_12504,N_10003,N_11786);
nand U12505 (N_12505,N_10297,N_10163);
and U12506 (N_12506,N_10648,N_10687);
and U12507 (N_12507,N_12301,N_12028);
nand U12508 (N_12508,N_11259,N_11815);
nand U12509 (N_12509,N_10179,N_11166);
nand U12510 (N_12510,N_11377,N_10674);
or U12511 (N_12511,N_11586,N_11578);
nand U12512 (N_12512,N_11539,N_12458);
and U12513 (N_12513,N_10897,N_12061);
xnor U12514 (N_12514,N_12260,N_10190);
and U12515 (N_12515,N_10430,N_11873);
and U12516 (N_12516,N_10012,N_11067);
or U12517 (N_12517,N_10632,N_10437);
nor U12518 (N_12518,N_11519,N_10072);
nor U12519 (N_12519,N_11318,N_11210);
and U12520 (N_12520,N_12396,N_11986);
nor U12521 (N_12521,N_10336,N_10733);
nand U12522 (N_12522,N_10928,N_10852);
nor U12523 (N_12523,N_11725,N_12094);
and U12524 (N_12524,N_10896,N_12346);
nand U12525 (N_12525,N_10989,N_12071);
or U12526 (N_12526,N_12119,N_10022);
nand U12527 (N_12527,N_11972,N_10882);
or U12528 (N_12528,N_12242,N_10419);
nand U12529 (N_12529,N_12059,N_11711);
and U12530 (N_12530,N_11205,N_10763);
nand U12531 (N_12531,N_10185,N_12058);
nor U12532 (N_12532,N_10106,N_10358);
nor U12533 (N_12533,N_12116,N_11253);
and U12534 (N_12534,N_12415,N_11899);
and U12535 (N_12535,N_12103,N_12039);
nand U12536 (N_12536,N_10409,N_10211);
nor U12537 (N_12537,N_11783,N_10694);
and U12538 (N_12538,N_11079,N_11187);
or U12539 (N_12539,N_10475,N_10976);
and U12540 (N_12540,N_11626,N_10286);
and U12541 (N_12541,N_10771,N_10904);
and U12542 (N_12542,N_10870,N_11323);
nor U12543 (N_12543,N_11439,N_10304);
or U12544 (N_12544,N_11189,N_10946);
nor U12545 (N_12545,N_11167,N_11928);
nor U12546 (N_12546,N_11707,N_10044);
nor U12547 (N_12547,N_12113,N_12120);
and U12548 (N_12548,N_10337,N_12251);
nand U12549 (N_12549,N_10488,N_11092);
or U12550 (N_12550,N_10355,N_10050);
and U12551 (N_12551,N_11973,N_10149);
xnor U12552 (N_12552,N_10945,N_11840);
nor U12553 (N_12553,N_12304,N_10381);
xnor U12554 (N_12554,N_11123,N_11833);
nand U12555 (N_12555,N_11788,N_10210);
and U12556 (N_12556,N_10467,N_10743);
nand U12557 (N_12557,N_10939,N_11097);
nand U12558 (N_12558,N_11593,N_10835);
nand U12559 (N_12559,N_11970,N_11800);
or U12560 (N_12560,N_12008,N_10324);
and U12561 (N_12561,N_12055,N_11152);
nor U12562 (N_12562,N_11057,N_11639);
xnor U12563 (N_12563,N_12087,N_11037);
xor U12564 (N_12564,N_11630,N_10957);
and U12565 (N_12565,N_10914,N_10237);
or U12566 (N_12566,N_11179,N_11546);
or U12567 (N_12567,N_10706,N_10585);
nor U12568 (N_12568,N_11749,N_11031);
nand U12569 (N_12569,N_11341,N_11008);
or U12570 (N_12570,N_11902,N_10907);
and U12571 (N_12571,N_12015,N_11803);
and U12572 (N_12572,N_12264,N_11299);
and U12573 (N_12573,N_10636,N_11016);
or U12574 (N_12574,N_12033,N_12351);
nor U12575 (N_12575,N_11868,N_10098);
xnor U12576 (N_12576,N_10645,N_10744);
nor U12577 (N_12577,N_10829,N_11818);
nor U12578 (N_12578,N_10507,N_11679);
nand U12579 (N_12579,N_11369,N_12140);
nand U12580 (N_12580,N_10735,N_10096);
nand U12581 (N_12581,N_10600,N_10081);
or U12582 (N_12582,N_11908,N_11676);
and U12583 (N_12583,N_10794,N_11081);
and U12584 (N_12584,N_11114,N_10684);
nand U12585 (N_12585,N_12338,N_10095);
nand U12586 (N_12586,N_11589,N_12115);
nor U12587 (N_12587,N_11584,N_12474);
and U12588 (N_12588,N_11681,N_10953);
nor U12589 (N_12589,N_10580,N_10532);
or U12590 (N_12590,N_10257,N_12130);
nand U12591 (N_12591,N_11610,N_12286);
nor U12592 (N_12592,N_11478,N_11825);
nor U12593 (N_12593,N_11145,N_11202);
and U12594 (N_12594,N_12089,N_12259);
or U12595 (N_12595,N_10695,N_10545);
and U12596 (N_12596,N_12313,N_11476);
and U12597 (N_12597,N_11754,N_10749);
nand U12598 (N_12598,N_11646,N_11449);
nor U12599 (N_12599,N_11820,N_12318);
nor U12600 (N_12600,N_11623,N_10084);
or U12601 (N_12601,N_12299,N_12029);
nor U12602 (N_12602,N_11311,N_11883);
and U12603 (N_12603,N_10254,N_10622);
and U12604 (N_12604,N_12454,N_10469);
and U12605 (N_12605,N_11433,N_11074);
or U12606 (N_12606,N_10589,N_11521);
nor U12607 (N_12607,N_10170,N_10745);
nand U12608 (N_12608,N_12037,N_11291);
or U12609 (N_12609,N_11385,N_10762);
or U12610 (N_12610,N_10736,N_11629);
or U12611 (N_12611,N_12020,N_12312);
nor U12612 (N_12612,N_11154,N_10028);
nor U12613 (N_12613,N_11680,N_10032);
nor U12614 (N_12614,N_10171,N_12300);
or U12615 (N_12615,N_10110,N_11772);
nor U12616 (N_12616,N_10857,N_10252);
and U12617 (N_12617,N_11326,N_10797);
nor U12618 (N_12618,N_10851,N_10992);
nand U12619 (N_12619,N_11743,N_11258);
and U12620 (N_12620,N_11251,N_11391);
or U12621 (N_12621,N_11019,N_12409);
nor U12622 (N_12622,N_10780,N_10544);
and U12623 (N_12623,N_10222,N_12155);
xor U12624 (N_12624,N_10754,N_11134);
and U12625 (N_12625,N_11319,N_11988);
or U12626 (N_12626,N_12297,N_11475);
xnor U12627 (N_12627,N_10868,N_10202);
and U12628 (N_12628,N_11766,N_11828);
nor U12629 (N_12629,N_10055,N_10356);
or U12630 (N_12630,N_10932,N_11028);
or U12631 (N_12631,N_10476,N_11588);
or U12632 (N_12632,N_11550,N_11601);
xnor U12633 (N_12633,N_11487,N_10231);
nand U12634 (N_12634,N_12105,N_11556);
nand U12635 (N_12635,N_11914,N_10923);
nand U12636 (N_12636,N_10327,N_11091);
nor U12637 (N_12637,N_10959,N_11795);
xor U12638 (N_12638,N_11327,N_12434);
or U12639 (N_12639,N_11156,N_11760);
or U12640 (N_12640,N_10727,N_10630);
and U12641 (N_12641,N_11477,N_10264);
and U12642 (N_12642,N_10315,N_12147);
nand U12643 (N_12643,N_10140,N_11456);
or U12644 (N_12644,N_11903,N_10302);
or U12645 (N_12645,N_10740,N_12226);
xnor U12646 (N_12646,N_12056,N_10993);
nor U12647 (N_12647,N_12319,N_10987);
xor U12648 (N_12648,N_11894,N_10118);
nand U12649 (N_12649,N_11242,N_10586);
or U12650 (N_12650,N_11075,N_11922);
nand U12651 (N_12651,N_11523,N_10485);
nor U12652 (N_12652,N_12229,N_10145);
and U12653 (N_12653,N_11400,N_12298);
and U12654 (N_12654,N_11463,N_11612);
and U12655 (N_12655,N_10714,N_12065);
xnor U12656 (N_12656,N_11822,N_10689);
or U12657 (N_12657,N_11437,N_10962);
and U12658 (N_12658,N_12218,N_12412);
and U12659 (N_12659,N_10561,N_11222);
or U12660 (N_12660,N_10093,N_11194);
or U12661 (N_12661,N_11513,N_11984);
and U12662 (N_12662,N_12287,N_10972);
nor U12663 (N_12663,N_10114,N_10538);
or U12664 (N_12664,N_12280,N_12159);
nand U12665 (N_12665,N_10970,N_12010);
and U12666 (N_12666,N_10439,N_10217);
nand U12667 (N_12667,N_10030,N_10018);
nor U12668 (N_12668,N_12151,N_11144);
nor U12669 (N_12669,N_11090,N_10508);
and U12670 (N_12670,N_12288,N_12278);
or U12671 (N_12671,N_11280,N_10865);
and U12672 (N_12672,N_12011,N_11193);
or U12673 (N_12673,N_10153,N_10563);
nand U12674 (N_12674,N_11733,N_10269);
or U12675 (N_12675,N_12202,N_11034);
or U12676 (N_12676,N_10380,N_11816);
nand U12677 (N_12677,N_11536,N_11959);
nand U12678 (N_12678,N_11673,N_11246);
nor U12679 (N_12679,N_10180,N_10633);
or U12680 (N_12680,N_12333,N_10479);
nand U12681 (N_12681,N_11324,N_11943);
nand U12682 (N_12682,N_10504,N_11622);
and U12683 (N_12683,N_12186,N_10646);
or U12684 (N_12684,N_10655,N_11579);
nand U12685 (N_12685,N_10524,N_11320);
and U12686 (N_12686,N_10331,N_11875);
and U12687 (N_12687,N_11184,N_11102);
or U12688 (N_12688,N_12201,N_10542);
or U12689 (N_12689,N_10301,N_12084);
nand U12690 (N_12690,N_11684,N_12073);
and U12691 (N_12691,N_11633,N_11613);
or U12692 (N_12692,N_11649,N_10390);
nor U12693 (N_12693,N_11412,N_11200);
or U12694 (N_12694,N_12368,N_10427);
nor U12695 (N_12695,N_12342,N_12187);
or U12696 (N_12696,N_11399,N_10201);
nand U12697 (N_12697,N_11503,N_10457);
or U12698 (N_12698,N_11462,N_10560);
and U12699 (N_12699,N_12230,N_10176);
and U12700 (N_12700,N_11926,N_12244);
xor U12701 (N_12701,N_11784,N_12355);
and U12702 (N_12702,N_10873,N_12265);
and U12703 (N_12703,N_11813,N_10635);
xor U12704 (N_12704,N_11804,N_10746);
nand U12705 (N_12705,N_10661,N_10604);
xnor U12706 (N_12706,N_10772,N_12173);
and U12707 (N_12707,N_10268,N_11862);
nor U12708 (N_12708,N_12361,N_10965);
nor U12709 (N_12709,N_12437,N_11013);
or U12710 (N_12710,N_12169,N_11295);
nor U12711 (N_12711,N_11070,N_10844);
and U12712 (N_12712,N_12335,N_11064);
xor U12713 (N_12713,N_11609,N_10000);
nor U12714 (N_12714,N_11349,N_11871);
nand U12715 (N_12715,N_10826,N_12377);
nor U12716 (N_12716,N_12408,N_10319);
and U12717 (N_12717,N_10291,N_10830);
and U12718 (N_12718,N_11055,N_10191);
nand U12719 (N_12719,N_10553,N_12375);
or U12720 (N_12720,N_10624,N_11290);
or U12721 (N_12721,N_10117,N_10434);
nor U12722 (N_12722,N_11287,N_12380);
nand U12723 (N_12723,N_10433,N_10471);
xnor U12724 (N_12724,N_11805,N_10186);
nor U12725 (N_12725,N_11559,N_10901);
and U12726 (N_12726,N_12072,N_12357);
xor U12727 (N_12727,N_12213,N_10383);
and U12728 (N_12728,N_11450,N_11562);
nor U12729 (N_12729,N_12464,N_12165);
nand U12730 (N_12730,N_11826,N_12080);
and U12731 (N_12731,N_12145,N_10934);
nand U12732 (N_12732,N_10782,N_10663);
nor U12733 (N_12733,N_10531,N_11552);
nand U12734 (N_12734,N_11504,N_10866);
or U12735 (N_12735,N_12382,N_11133);
and U12736 (N_12736,N_11351,N_11595);
and U12737 (N_12737,N_10199,N_12488);
and U12738 (N_12738,N_11239,N_11590);
xor U12739 (N_12739,N_12180,N_11175);
or U12740 (N_12740,N_12423,N_11611);
or U12741 (N_12741,N_10869,N_11047);
and U12742 (N_12742,N_11597,N_10951);
xor U12743 (N_12743,N_11505,N_11538);
and U12744 (N_12744,N_11480,N_11457);
or U12745 (N_12745,N_10513,N_10097);
and U12746 (N_12746,N_12499,N_12107);
nand U12747 (N_12747,N_11348,N_11614);
nor U12748 (N_12748,N_10623,N_11365);
xnor U12749 (N_12749,N_10379,N_10481);
and U12750 (N_12750,N_12303,N_12066);
nand U12751 (N_12751,N_10892,N_11464);
nor U12752 (N_12752,N_10265,N_10718);
nor U12753 (N_12753,N_11853,N_11455);
nor U12754 (N_12754,N_10020,N_12344);
nand U12755 (N_12755,N_11855,N_11471);
and U12756 (N_12756,N_11050,N_12076);
xnor U12757 (N_12757,N_11930,N_10207);
nand U12758 (N_12758,N_10647,N_11838);
or U12759 (N_12759,N_10119,N_11953);
nor U12760 (N_12760,N_10124,N_10443);
nand U12761 (N_12761,N_11426,N_10966);
nand U12762 (N_12762,N_12021,N_11044);
or U12763 (N_12763,N_10444,N_10602);
nor U12764 (N_12764,N_10593,N_12403);
nand U12765 (N_12765,N_10594,N_10064);
nand U12766 (N_12766,N_11007,N_10209);
nand U12767 (N_12767,N_10960,N_11151);
nor U12768 (N_12768,N_10339,N_10378);
and U12769 (N_12769,N_11137,N_10537);
or U12770 (N_12770,N_11583,N_11916);
or U12771 (N_12771,N_10157,N_11359);
and U12772 (N_12772,N_12188,N_11925);
nor U12773 (N_12773,N_11999,N_10223);
nand U12774 (N_12774,N_10637,N_10823);
nor U12775 (N_12775,N_10332,N_12389);
or U12776 (N_12776,N_10426,N_10458);
or U12777 (N_12777,N_11744,N_11077);
nor U12778 (N_12778,N_10348,N_10748);
or U12779 (N_12779,N_10193,N_10592);
nand U12780 (N_12780,N_11454,N_10468);
and U12781 (N_12781,N_10683,N_10528);
or U12782 (N_12782,N_12426,N_10385);
or U12783 (N_12783,N_10420,N_11960);
nor U12784 (N_12784,N_12197,N_11276);
nand U12785 (N_12785,N_11951,N_11110);
or U12786 (N_12786,N_11900,N_10307);
or U12787 (N_12787,N_10539,N_10878);
nor U12788 (N_12788,N_11421,N_11876);
or U12789 (N_12789,N_10569,N_10527);
or U12790 (N_12790,N_11850,N_10952);
and U12791 (N_12791,N_12152,N_11052);
and U12792 (N_12792,N_10295,N_12024);
or U12793 (N_12793,N_10854,N_11344);
nand U12794 (N_12794,N_11765,N_11432);
and U12795 (N_12795,N_11024,N_10352);
and U12796 (N_12796,N_11026,N_10747);
and U12797 (N_12797,N_11640,N_11366);
nor U12798 (N_12798,N_10243,N_11168);
xor U12799 (N_12799,N_11461,N_12217);
xor U12800 (N_12800,N_12134,N_10078);
or U12801 (N_12801,N_11025,N_11058);
xnor U12802 (N_12802,N_10455,N_11987);
nand U12803 (N_12803,N_11897,N_12214);
xor U12804 (N_12804,N_12290,N_10449);
and U12805 (N_12805,N_12253,N_12471);
and U12806 (N_12806,N_10376,N_11491);
or U12807 (N_12807,N_10833,N_10737);
or U12808 (N_12808,N_10858,N_10465);
and U12809 (N_12809,N_11098,N_11216);
or U12810 (N_12810,N_10871,N_10926);
and U12811 (N_12811,N_10521,N_10918);
or U12812 (N_12812,N_11206,N_10891);
nand U12813 (N_12813,N_11962,N_10599);
nand U12814 (N_12814,N_10460,N_12305);
or U12815 (N_12815,N_12281,N_11674);
nand U12816 (N_12816,N_12388,N_11762);
nor U12817 (N_12817,N_12402,N_11218);
nand U12818 (N_12818,N_11572,N_12164);
xnor U12819 (N_12819,N_11036,N_10391);
nand U12820 (N_12820,N_12171,N_10396);
and U12821 (N_12821,N_11895,N_10054);
nor U12822 (N_12822,N_11657,N_11186);
nor U12823 (N_12823,N_11856,N_12157);
nand U12824 (N_12824,N_12367,N_12466);
and U12825 (N_12825,N_10898,N_12496);
nor U12826 (N_12826,N_12406,N_11996);
and U12827 (N_12827,N_10716,N_10318);
and U12828 (N_12828,N_10877,N_10860);
xnor U12829 (N_12829,N_12199,N_10841);
or U12830 (N_12830,N_11923,N_12381);
nand U12831 (N_12831,N_12407,N_10935);
xor U12832 (N_12832,N_12181,N_10496);
xor U12833 (N_12833,N_12459,N_10101);
and U12834 (N_12834,N_10998,N_11516);
nor U12835 (N_12835,N_10653,N_11938);
nor U12836 (N_12836,N_12472,N_12341);
or U12837 (N_12837,N_11022,N_11231);
nor U12838 (N_12838,N_10678,N_11790);
nor U12839 (N_12839,N_11402,N_11874);
nand U12840 (N_12840,N_12441,N_10685);
or U12841 (N_12841,N_11220,N_11105);
nand U12842 (N_12842,N_12349,N_11274);
nor U12843 (N_12843,N_12436,N_11940);
and U12844 (N_12844,N_11185,N_12206);
or U12845 (N_12845,N_11732,N_10876);
nand U12846 (N_12846,N_10523,N_11130);
xor U12847 (N_12847,N_11333,N_10472);
nand U12848 (N_12848,N_12234,N_10533);
nand U12849 (N_12849,N_10205,N_11709);
and U12850 (N_12850,N_11362,N_11226);
or U12851 (N_12851,N_12476,N_11136);
nand U12852 (N_12852,N_11283,N_11672);
and U12853 (N_12853,N_11298,N_10731);
or U12854 (N_12854,N_11997,N_12284);
and U12855 (N_12855,N_12438,N_11252);
nor U12856 (N_12856,N_10247,N_10280);
or U12857 (N_12857,N_12467,N_12495);
xor U12858 (N_12858,N_10491,N_11380);
nor U12859 (N_12859,N_10256,N_11779);
nor U12860 (N_12860,N_10839,N_11106);
and U12861 (N_12861,N_11886,N_11697);
xor U12862 (N_12862,N_11071,N_11702);
or U12863 (N_12863,N_10421,N_11135);
nor U12864 (N_12864,N_11677,N_11864);
xnor U12865 (N_12865,N_10795,N_11357);
xor U12866 (N_12866,N_10392,N_10130);
nand U12867 (N_12867,N_10616,N_11924);
nor U12868 (N_12868,N_10314,N_12205);
and U12869 (N_12869,N_11419,N_11778);
and U12870 (N_12870,N_12099,N_12210);
and U12871 (N_12871,N_10224,N_10942);
nand U12872 (N_12872,N_11496,N_10813);
and U12873 (N_12873,N_10729,N_11666);
nand U12874 (N_12874,N_11889,N_10732);
nor U12875 (N_12875,N_12399,N_12490);
or U12876 (N_12876,N_12121,N_10956);
nand U12877 (N_12877,N_11140,N_11248);
xnor U12878 (N_12878,N_11670,N_12168);
nand U12879 (N_12879,N_11934,N_11761);
xnor U12880 (N_12880,N_12445,N_12394);
nor U12881 (N_12881,N_11753,N_10131);
and U12882 (N_12882,N_11568,N_10828);
nor U12883 (N_12883,N_11269,N_10981);
or U12884 (N_12884,N_11228,N_10525);
nand U12885 (N_12885,N_10397,N_10936);
nor U12886 (N_12886,N_10399,N_12296);
or U12887 (N_12887,N_10151,N_10010);
nand U12888 (N_12888,N_10758,N_12443);
and U12889 (N_12889,N_10424,N_10824);
or U12890 (N_12890,N_11303,N_10053);
nand U12891 (N_12891,N_12209,N_10719);
or U12892 (N_12892,N_10529,N_12497);
or U12893 (N_12893,N_11484,N_10750);
nor U12894 (N_12894,N_11992,N_11401);
and U12895 (N_12895,N_11101,N_11386);
nand U12896 (N_12896,N_10173,N_10900);
and U12897 (N_12897,N_10177,N_12207);
and U12898 (N_12898,N_10009,N_10775);
nand U12899 (N_12899,N_11501,N_11499);
or U12900 (N_12900,N_12292,N_11961);
nand U12901 (N_12901,N_11625,N_11606);
and U12902 (N_12902,N_11658,N_11627);
or U12903 (N_12903,N_11466,N_10517);
nor U12904 (N_12904,N_10061,N_12391);
or U12905 (N_12905,N_11937,N_10410);
nor U12906 (N_12906,N_10920,N_11650);
nand U12907 (N_12907,N_12309,N_10345);
xor U12908 (N_12908,N_10321,N_11139);
or U12909 (N_12909,N_12270,N_11155);
nand U12910 (N_12910,N_12468,N_11302);
xnor U12911 (N_12911,N_10271,N_12200);
or U12912 (N_12912,N_12254,N_10997);
or U12913 (N_12913,N_12078,N_11279);
nand U12914 (N_12914,N_10334,N_11289);
nand U12915 (N_12915,N_11416,N_11498);
and U12916 (N_12916,N_11817,N_10627);
or U12917 (N_12917,N_11963,N_10006);
xnor U12918 (N_12918,N_11909,N_11409);
nor U12919 (N_12919,N_12189,N_10040);
and U12920 (N_12920,N_11423,N_12422);
or U12921 (N_12921,N_10608,N_11214);
nor U12922 (N_12922,N_11018,N_12461);
or U12923 (N_12923,N_11919,N_12215);
nand U12924 (N_12924,N_12135,N_12345);
and U12925 (N_12925,N_10484,N_12117);
and U12926 (N_12926,N_11729,N_11901);
nand U12927 (N_12927,N_11624,N_12032);
nor U12928 (N_12928,N_11527,N_11212);
xor U12929 (N_12929,N_11159,N_12354);
nand U12930 (N_12930,N_11892,N_11882);
and U12931 (N_12931,N_11844,N_10776);
nand U12932 (N_12932,N_10221,N_10559);
or U12933 (N_12933,N_10711,N_11254);
xnor U12934 (N_12934,N_11541,N_10790);
nand U12935 (N_12935,N_11076,N_10577);
nor U12936 (N_12936,N_11950,N_10875);
xor U12937 (N_12937,N_10122,N_12240);
xor U12938 (N_12938,N_11334,N_12228);
nor U12939 (N_12939,N_10365,N_10510);
nand U12940 (N_12940,N_10405,N_12393);
nor U12941 (N_12941,N_10628,N_10004);
and U12942 (N_12942,N_10575,N_12469);
or U12943 (N_12943,N_11387,N_11294);
nand U12944 (N_12944,N_10849,N_10492);
nor U12945 (N_12945,N_10233,N_12285);
nand U12946 (N_12946,N_10283,N_11330);
nor U12947 (N_12947,N_10300,N_12343);
nand U12948 (N_12948,N_11814,N_10698);
nand U12949 (N_12949,N_11734,N_11296);
and U12950 (N_12950,N_11967,N_10487);
nor U12951 (N_12951,N_10086,N_10169);
or U12952 (N_12952,N_10500,N_10774);
nor U12953 (N_12953,N_11285,N_12035);
nand U12954 (N_12954,N_10969,N_12125);
and U12955 (N_12955,N_12144,N_11748);
nand U12956 (N_12956,N_11667,N_11858);
and U12957 (N_12957,N_10768,N_11379);
xor U12958 (N_12958,N_10943,N_10245);
xnor U12959 (N_12959,N_11099,N_11860);
xor U12960 (N_12960,N_11635,N_10219);
xor U12961 (N_12961,N_11575,N_10329);
and U12962 (N_12962,N_10335,N_10846);
and U12963 (N_12963,N_11605,N_10933);
or U12964 (N_12964,N_11941,N_11196);
or U12965 (N_12965,N_12175,N_11724);
nand U12966 (N_12966,N_10979,N_12167);
nor U12967 (N_12967,N_11810,N_12446);
or U12968 (N_12968,N_11708,N_11616);
nor U12969 (N_12969,N_10292,N_11413);
nor U12970 (N_12970,N_11979,N_12162);
or U12971 (N_12971,N_11001,N_11109);
or U12972 (N_12972,N_12249,N_12353);
nand U12973 (N_12973,N_10546,N_11878);
nor U12974 (N_12974,N_10549,N_11440);
nor U12975 (N_12975,N_10349,N_11971);
or U12976 (N_12976,N_12455,N_10584);
nand U12977 (N_12977,N_11404,N_10804);
nor U12978 (N_12978,N_10669,N_10212);
xor U12979 (N_12979,N_11411,N_10890);
nand U12980 (N_12980,N_11170,N_11338);
and U12981 (N_12981,N_11763,N_11585);
nor U12982 (N_12982,N_11715,N_10051);
and U12983 (N_12983,N_11321,N_10917);
and U12984 (N_12984,N_11208,N_11794);
xor U12985 (N_12985,N_11192,N_12031);
and U12986 (N_12986,N_10042,N_12386);
or U12987 (N_12987,N_10371,N_12090);
or U12988 (N_12988,N_11558,N_11243);
xor U12989 (N_12989,N_10742,N_11481);
nand U12990 (N_12990,N_10834,N_11436);
nor U12991 (N_12991,N_12384,N_11373);
nor U12992 (N_12992,N_11881,N_10428);
nor U12993 (N_12993,N_11162,N_12314);
xnor U12994 (N_12994,N_12272,N_12231);
nor U12995 (N_12995,N_12350,N_11495);
nand U12996 (N_12996,N_12000,N_10293);
or U12997 (N_12997,N_10692,N_12060);
xnor U12998 (N_12998,N_11087,N_11195);
nand U12999 (N_12999,N_11719,N_11773);
and U13000 (N_13000,N_11500,N_10103);
nand U13001 (N_13001,N_11257,N_11172);
or U13002 (N_13002,N_10195,N_12079);
nor U13003 (N_13003,N_10251,N_10069);
or U13004 (N_13004,N_10657,N_11122);
nand U13005 (N_13005,N_10127,N_11775);
nor U13006 (N_13006,N_10978,N_12129);
and U13007 (N_13007,N_10842,N_12005);
nand U13008 (N_13008,N_10340,N_10715);
and U13009 (N_13009,N_10760,N_10367);
or U13010 (N_13010,N_10576,N_11347);
or U13011 (N_13011,N_11352,N_11782);
nand U13012 (N_13012,N_10654,N_10609);
or U13013 (N_13013,N_10074,N_10995);
nor U13014 (N_13014,N_10950,N_11010);
nand U13015 (N_13015,N_11266,N_10407);
and U13016 (N_13016,N_11554,N_10175);
and U13017 (N_13017,N_12481,N_10634);
xnor U13018 (N_13018,N_12102,N_11180);
or U13019 (N_13019,N_11913,N_11354);
or U13020 (N_13020,N_11278,N_10466);
nand U13021 (N_13021,N_12273,N_12179);
nand U13022 (N_13022,N_12414,N_11685);
or U13023 (N_13023,N_10905,N_10425);
nand U13024 (N_13024,N_11931,N_10066);
nand U13025 (N_13025,N_12081,N_11126);
or U13026 (N_13026,N_11418,N_10764);
nor U13027 (N_13027,N_10658,N_10696);
or U13028 (N_13028,N_12095,N_11486);
nand U13029 (N_13029,N_11918,N_10982);
nand U13030 (N_13030,N_10429,N_10279);
nor U13031 (N_13031,N_11631,N_11129);
nand U13032 (N_13032,N_11582,N_10342);
or U13033 (N_13033,N_11372,N_10029);
or U13034 (N_13034,N_10226,N_11002);
nor U13035 (N_13035,N_11660,N_10373);
xor U13036 (N_13036,N_10255,N_11683);
and U13037 (N_13037,N_10990,N_11331);
nor U13038 (N_13038,N_12366,N_11759);
nand U13039 (N_13039,N_12294,N_10230);
and U13040 (N_13040,N_12022,N_12379);
nor U13041 (N_13041,N_11509,N_10075);
nand U13042 (N_13042,N_11005,N_12027);
or U13043 (N_13043,N_10354,N_11093);
nor U13044 (N_13044,N_10143,N_10708);
xor U13045 (N_13045,N_10232,N_11511);
or U13046 (N_13046,N_10713,N_10741);
nand U13047 (N_13047,N_11698,N_12092);
nand U13048 (N_13048,N_12158,N_12348);
or U13049 (N_13049,N_12250,N_10693);
nor U13050 (N_13050,N_11406,N_12203);
xnor U13051 (N_13051,N_12276,N_10887);
nor U13052 (N_13052,N_11103,N_11383);
nand U13053 (N_13053,N_10362,N_10902);
or U13054 (N_13054,N_10401,N_12337);
nand U13055 (N_13055,N_11229,N_10406);
and U13056 (N_13056,N_11799,N_11469);
and U13057 (N_13057,N_11488,N_11265);
xor U13058 (N_13058,N_10578,N_10007);
nand U13059 (N_13059,N_11273,N_12246);
or U13060 (N_13060,N_10903,N_10435);
xor U13061 (N_13061,N_12450,N_12126);
xnor U13062 (N_13062,N_11211,N_10515);
nand U13063 (N_13063,N_12470,N_11035);
and U13064 (N_13064,N_11394,N_11730);
and U13065 (N_13065,N_12263,N_12405);
nor U13066 (N_13066,N_10152,N_10991);
nand U13067 (N_13067,N_10611,N_12012);
and U13068 (N_13068,N_12216,N_10817);
xor U13069 (N_13069,N_10543,N_12332);
nand U13070 (N_13070,N_12325,N_12269);
nor U13071 (N_13071,N_11821,N_10767);
or U13072 (N_13072,N_11332,N_10784);
and U13073 (N_13073,N_10587,N_10431);
nor U13074 (N_13074,N_12385,N_12457);
nand U13075 (N_13075,N_11435,N_11000);
nand U13076 (N_13076,N_10412,N_12427);
or U13077 (N_13077,N_11525,N_11848);
and U13078 (N_13078,N_11978,N_11577);
nor U13079 (N_13079,N_12177,N_12052);
or U13080 (N_13080,N_10619,N_10659);
nor U13081 (N_13081,N_10512,N_11793);
nor U13082 (N_13082,N_11549,N_10192);
or U13083 (N_13083,N_11617,N_11304);
xor U13084 (N_13084,N_11806,N_12484);
or U13085 (N_13085,N_11742,N_10388);
nor U13086 (N_13086,N_10244,N_10710);
nand U13087 (N_13087,N_11990,N_11407);
xnor U13088 (N_13088,N_12241,N_11735);
nor U13089 (N_13089,N_11542,N_11221);
nor U13090 (N_13090,N_10441,N_11427);
nor U13091 (N_13091,N_11510,N_11392);
or U13092 (N_13092,N_10206,N_11599);
or U13093 (N_13093,N_11116,N_10005);
or U13094 (N_13094,N_12100,N_12362);
nand U13095 (N_13095,N_11428,N_11989);
xnor U13096 (N_13096,N_11796,N_11085);
and U13097 (N_13097,N_10246,N_10141);
or U13098 (N_13098,N_11004,N_11173);
nand U13099 (N_13099,N_10023,N_10912);
or U13100 (N_13100,N_11410,N_11768);
nor U13101 (N_13101,N_11866,N_12046);
nor U13102 (N_13102,N_11183,N_10451);
nand U13103 (N_13103,N_11169,N_12452);
and U13104 (N_13104,N_12424,N_11644);
nand U13105 (N_13105,N_11048,N_12358);
nor U13106 (N_13106,N_10105,N_10888);
xnor U13107 (N_13107,N_12238,N_11514);
nand U13108 (N_13108,N_10453,N_10160);
or U13109 (N_13109,N_12232,N_10639);
nor U13110 (N_13110,N_11722,N_11381);
xnor U13111 (N_13111,N_11458,N_10071);
nand U13112 (N_13112,N_11236,N_10721);
nand U13113 (N_13113,N_12091,N_11203);
xor U13114 (N_13114,N_10322,N_11506);
or U13115 (N_13115,N_10121,N_10422);
or U13116 (N_13116,N_12146,N_11147);
nor U13117 (N_13117,N_10369,N_11929);
and U13118 (N_13118,N_10432,N_10166);
nand U13119 (N_13119,N_11376,N_12404);
or U13120 (N_13120,N_10704,N_11755);
nand U13121 (N_13121,N_12463,N_11260);
and U13122 (N_13122,N_11078,N_10884);
or U13123 (N_13123,N_10603,N_11567);
nand U13124 (N_13124,N_10941,N_11238);
and U13125 (N_13125,N_10783,N_11198);
or U13126 (N_13126,N_10922,N_12044);
or U13127 (N_13127,N_10514,N_12172);
nor U13128 (N_13128,N_11665,N_12373);
nor U13129 (N_13129,N_12248,N_12137);
or U13130 (N_13130,N_10757,N_10499);
nor U13131 (N_13131,N_10415,N_11204);
nand U13132 (N_13132,N_10060,N_10436);
and U13133 (N_13133,N_11465,N_12063);
nand U13134 (N_13134,N_10203,N_11507);
xnor U13135 (N_13135,N_11638,N_10135);
nor U13136 (N_13136,N_11792,N_11745);
or U13137 (N_13137,N_10493,N_12143);
or U13138 (N_13138,N_11712,N_11936);
and U13139 (N_13139,N_10234,N_12139);
and U13140 (N_13140,N_11824,N_11378);
and U13141 (N_13141,N_10534,N_11060);
and U13142 (N_13142,N_10359,N_10077);
nor U13143 (N_13143,N_12034,N_11396);
or U13144 (N_13144,N_12323,N_11301);
xnor U13145 (N_13145,N_10100,N_12266);
and U13146 (N_13146,N_11857,N_10214);
nor U13147 (N_13147,N_11393,N_10720);
nand U13148 (N_13148,N_11920,N_10015);
or U13149 (N_13149,N_11017,N_11153);
nand U13150 (N_13150,N_12395,N_12227);
and U13151 (N_13151,N_10281,N_12485);
nor U13152 (N_13152,N_10501,N_10102);
nand U13153 (N_13153,N_10184,N_11890);
or U13154 (N_13154,N_10643,N_11245);
nand U13155 (N_13155,N_11851,N_10555);
and U13156 (N_13156,N_10261,N_11096);
or U13157 (N_13157,N_10800,N_10303);
and U13158 (N_13158,N_10773,N_12363);
or U13159 (N_13159,N_10109,N_11655);
nor U13160 (N_13160,N_10403,N_12018);
nand U13161 (N_13161,N_12174,N_10473);
and U13162 (N_13162,N_11801,N_10417);
and U13163 (N_13163,N_12184,N_11863);
or U13164 (N_13164,N_12036,N_10438);
nand U13165 (N_13165,N_11374,N_10574);
nor U13166 (N_13166,N_11165,N_10266);
nand U13167 (N_13167,N_10700,N_11069);
nor U13168 (N_13168,N_12096,N_11811);
or U13169 (N_13169,N_10021,N_10881);
or U13170 (N_13170,N_12327,N_11781);
nor U13171 (N_13171,N_10518,N_11921);
nor U13172 (N_13172,N_11250,N_10346);
xor U13173 (N_13173,N_11056,N_12085);
nand U13174 (N_13174,N_11600,N_10111);
nor U13175 (N_13175,N_10208,N_10867);
and U13176 (N_13176,N_11741,N_11408);
or U13177 (N_13177,N_11607,N_11335);
and U13178 (N_13178,N_11974,N_10477);
or U13179 (N_13179,N_11240,N_11720);
nand U13180 (N_13180,N_10855,N_10344);
nand U13181 (N_13181,N_11422,N_10240);
nor U13182 (N_13182,N_12493,N_12315);
nor U13183 (N_13183,N_10320,N_11532);
or U13184 (N_13184,N_10387,N_10506);
xnor U13185 (N_13185,N_10091,N_10285);
nor U13186 (N_13186,N_12465,N_10831);
nand U13187 (N_13187,N_11854,N_10906);
nor U13188 (N_13188,N_12161,N_12256);
and U13189 (N_13189,N_12068,N_12326);
nor U13190 (N_13190,N_12019,N_10400);
or U13191 (N_13191,N_11181,N_10258);
nor U13192 (N_13192,N_12009,N_10822);
nor U13193 (N_13193,N_11714,N_12237);
xnor U13194 (N_13194,N_10672,N_10447);
nor U13195 (N_13195,N_11580,N_11746);
and U13196 (N_13196,N_10819,N_11117);
nor U13197 (N_13197,N_10310,N_11176);
and U13198 (N_13198,N_10155,N_12328);
nor U13199 (N_13199,N_10921,N_10489);
nand U13200 (N_13200,N_10677,N_10238);
nand U13201 (N_13201,N_11118,N_12223);
nor U13202 (N_13202,N_11264,N_11954);
nor U13203 (N_13203,N_11446,N_10058);
nor U13204 (N_13204,N_10011,N_11736);
nand U13205 (N_13205,N_12433,N_11594);
or U13206 (N_13206,N_11777,N_12336);
xnor U13207 (N_13207,N_12483,N_12245);
xnor U13208 (N_13208,N_11642,N_11027);
or U13209 (N_13209,N_10927,N_11769);
nand U13210 (N_13210,N_12420,N_10540);
nand U13211 (N_13211,N_11415,N_12132);
nor U13212 (N_13212,N_10810,N_10495);
nand U13213 (N_13213,N_10899,N_10550);
or U13214 (N_13214,N_10364,N_10394);
or U13215 (N_13215,N_11910,N_11812);
nand U13216 (N_13216,N_10699,N_11015);
or U13217 (N_13217,N_12045,N_10734);
nor U13218 (N_13218,N_10838,N_10343);
nor U13219 (N_13219,N_11620,N_11217);
and U13220 (N_13220,N_10347,N_10606);
or U13221 (N_13221,N_10625,N_10673);
nor U13222 (N_13222,N_10404,N_11830);
nor U13223 (N_13223,N_10666,N_11718);
nand U13224 (N_13224,N_11089,N_10984);
nor U13225 (N_13225,N_10445,N_11682);
xnor U13226 (N_13226,N_12002,N_11199);
or U13227 (N_13227,N_10803,N_11694);
nand U13228 (N_13228,N_11149,N_11837);
and U13229 (N_13229,N_10931,N_10601);
nand U13230 (N_13230,N_10765,N_12293);
xor U13231 (N_13231,N_10919,N_11063);
nand U13232 (N_13232,N_12017,N_10617);
xnor U13233 (N_13233,N_10861,N_12439);
or U13234 (N_13234,N_12093,N_11489);
nor U13235 (N_13235,N_10668,N_10181);
or U13236 (N_13236,N_10641,N_11038);
nor U13237 (N_13237,N_12317,N_11329);
nand U13238 (N_13238,N_10325,N_11643);
nor U13239 (N_13239,N_11148,N_12182);
nor U13240 (N_13240,N_12320,N_10129);
or U13241 (N_13241,N_10788,N_10218);
nor U13242 (N_13242,N_11494,N_11687);
and U13243 (N_13243,N_12311,N_10798);
nor U13244 (N_13244,N_11297,N_11654);
xor U13245 (N_13245,N_11981,N_11121);
and U13246 (N_13246,N_11947,N_11482);
nand U13247 (N_13247,N_11945,N_10705);
or U13248 (N_13248,N_10681,N_10853);
nor U13249 (N_13249,N_10650,N_10198);
or U13250 (N_13250,N_10288,N_10112);
nand U13251 (N_13251,N_11739,N_11747);
and U13252 (N_13252,N_11982,N_11006);
and U13253 (N_13253,N_11780,N_10967);
and U13254 (N_13254,N_12101,N_12435);
nand U13255 (N_13255,N_11524,N_10290);
nor U13256 (N_13256,N_10787,N_12419);
or U13257 (N_13257,N_10260,N_10649);
and U13258 (N_13258,N_10662,N_10278);
xor U13259 (N_13259,N_11662,N_10660);
nand U13260 (N_13260,N_10893,N_10618);
and U13261 (N_13261,N_12070,N_10880);
nand U13262 (N_13262,N_10996,N_10094);
nor U13263 (N_13263,N_12243,N_11345);
or U13264 (N_13264,N_10194,N_11809);
nor U13265 (N_13265,N_11598,N_12097);
or U13266 (N_13266,N_11424,N_10450);
or U13267 (N_13267,N_11158,N_10631);
nor U13268 (N_13268,N_11030,N_11219);
xnor U13269 (N_13269,N_10910,N_10411);
nor U13270 (N_13270,N_12447,N_10626);
or U13271 (N_13271,N_10026,N_10859);
and U13272 (N_13272,N_12030,N_11459);
and U13273 (N_13273,N_10948,N_10464);
nor U13274 (N_13274,N_11115,N_10068);
nor U13275 (N_13275,N_10305,N_12440);
or U13276 (N_13276,N_11764,N_10323);
and U13277 (N_13277,N_12051,N_10595);
and U13278 (N_13278,N_12478,N_11807);
nand U13279 (N_13279,N_11360,N_12411);
nor U13280 (N_13280,N_10675,N_10667);
or U13281 (N_13281,N_11234,N_12392);
nand U13282 (N_13282,N_10452,N_11281);
xor U13283 (N_13283,N_11138,N_11268);
or U13284 (N_13284,N_10272,N_10478);
or U13285 (N_13285,N_12486,N_10818);
nor U13286 (N_13286,N_11716,N_12212);
and U13287 (N_13287,N_10955,N_10498);
xor U13288 (N_13288,N_12178,N_11430);
and U13289 (N_13289,N_10656,N_10299);
nand U13290 (N_13290,N_11995,N_10812);
xnor U13291 (N_13291,N_10591,N_10115);
or U13292 (N_13292,N_11776,N_11686);
xor U13293 (N_13293,N_11086,N_10353);
nand U13294 (N_13294,N_11073,N_10686);
and U13295 (N_13295,N_10133,N_10123);
nor U13296 (N_13296,N_10583,N_10070);
nand U13297 (N_13297,N_10259,N_10267);
nor U13298 (N_13298,N_10092,N_10188);
nor U13299 (N_13299,N_11322,N_11191);
nor U13300 (N_13300,N_11740,N_11977);
nand U13301 (N_13301,N_11717,N_10605);
or U13302 (N_13302,N_11839,N_10582);
and U13303 (N_13303,N_12106,N_11425);
nor U13304 (N_13304,N_12082,N_12131);
or U13305 (N_13305,N_12487,N_10423);
nand U13306 (N_13306,N_11441,N_11602);
and U13307 (N_13307,N_10530,N_10548);
or U13308 (N_13308,N_10691,N_10330);
and U13309 (N_13309,N_10554,N_11468);
nor U13310 (N_13310,N_12307,N_11307);
nor U13311 (N_13311,N_11157,N_11653);
and U13312 (N_13312,N_11367,N_10132);
nand U13313 (N_13313,N_10014,N_11171);
nor U13314 (N_13314,N_10973,N_10845);
or U13315 (N_13315,N_10013,N_12050);
xor U13316 (N_13316,N_10802,N_12431);
and U13317 (N_13317,N_10816,N_11353);
xnor U13318 (N_13318,N_11976,N_12138);
nor U13319 (N_13319,N_10250,N_11045);
and U13320 (N_13320,N_10035,N_10316);
nor U13321 (N_13321,N_12222,N_12111);
xnor U13322 (N_13322,N_10724,N_12416);
or U13323 (N_13323,N_12421,N_11869);
nor U13324 (N_13324,N_11703,N_11272);
nand U13325 (N_13325,N_12160,N_10309);
nor U13326 (N_13326,N_10895,N_11980);
nor U13327 (N_13327,N_10338,N_10726);
or U13328 (N_13328,N_10370,N_10139);
and U13329 (N_13329,N_11692,N_11223);
nand U13330 (N_13330,N_10215,N_10147);
nor U13331 (N_13331,N_10885,N_11497);
xor U13332 (N_13332,N_11618,N_10516);
and U13333 (N_13333,N_10270,N_11738);
nand U13334 (N_13334,N_10375,N_11062);
xnor U13335 (N_13335,N_12224,N_11576);
nand U13336 (N_13336,N_10413,N_10886);
nor U13337 (N_13337,N_11548,N_10057);
xnor U13338 (N_13338,N_12114,N_10083);
and U13339 (N_13339,N_11100,N_10395);
nand U13340 (N_13340,N_11355,N_11284);
and U13341 (N_13341,N_12014,N_10805);
and U13342 (N_13342,N_11188,N_11949);
xnor U13343 (N_13343,N_11596,N_10463);
and U13344 (N_13344,N_12400,N_11808);
or U13345 (N_13345,N_10916,N_10864);
nor U13346 (N_13346,N_12306,N_10642);
or U13347 (N_13347,N_11958,N_10062);
or U13348 (N_13348,N_10676,N_12352);
nand U13349 (N_13349,N_11068,N_11721);
nor U13350 (N_13350,N_12262,N_11420);
nor U13351 (N_13351,N_10236,N_10679);
and U13352 (N_13352,N_10806,N_12053);
or U13353 (N_13353,N_11647,N_10761);
nand U13354 (N_13354,N_11445,N_12108);
xor U13355 (N_13355,N_10228,N_11787);
or U13356 (N_13356,N_11518,N_12359);
and U13357 (N_13357,N_11942,N_10474);
nand U13358 (N_13358,N_10402,N_10766);
or U13359 (N_13359,N_10248,N_11132);
nor U13360 (N_13360,N_10613,N_12124);
nand U13361 (N_13361,N_12149,N_12442);
or U13362 (N_13362,N_10128,N_11182);
or U13363 (N_13363,N_10386,N_11011);
and U13364 (N_13364,N_10059,N_10811);
and U13365 (N_13365,N_11964,N_11414);
and U13366 (N_13366,N_11143,N_12239);
and U13367 (N_13367,N_12310,N_10126);
nand U13368 (N_13368,N_11150,N_12233);
or U13369 (N_13369,N_11308,N_11131);
and U13370 (N_13370,N_11905,N_12267);
or U13371 (N_13371,N_11261,N_11314);
nor U13372 (N_13372,N_11213,N_10308);
or U13373 (N_13373,N_12475,N_11933);
xnor U13374 (N_13374,N_10863,N_11994);
and U13375 (N_13375,N_11040,N_10730);
and U13376 (N_13376,N_11340,N_10227);
xnor U13377 (N_13377,N_10480,N_11564);
nand U13378 (N_13378,N_11443,N_11288);
nor U13379 (N_13379,N_12195,N_10930);
and U13380 (N_13380,N_10688,N_10273);
or U13381 (N_13381,N_10187,N_11975);
or U13382 (N_13382,N_10041,N_11767);
or U13383 (N_13383,N_12185,N_11472);
nor U13384 (N_13384,N_10148,N_11847);
and U13385 (N_13385,N_10189,N_12211);
nor U13386 (N_13386,N_12040,N_11845);
xor U13387 (N_13387,N_12261,N_11530);
xnor U13388 (N_13388,N_12252,N_10317);
or U13389 (N_13389,N_11473,N_11361);
nand U13390 (N_13390,N_11621,N_10883);
and U13391 (N_13391,N_11834,N_11267);
nor U13392 (N_13392,N_11517,N_11880);
and U13393 (N_13393,N_10294,N_10547);
or U13394 (N_13394,N_12154,N_12378);
nand U13395 (N_13395,N_11628,N_10827);
xor U13396 (N_13396,N_10980,N_12192);
nor U13397 (N_13397,N_11831,N_12016);
nand U13398 (N_13398,N_10638,N_12498);
nand U13399 (N_13399,N_11033,N_12316);
and U13400 (N_13400,N_11244,N_10043);
nor U13401 (N_13401,N_11823,N_12271);
and U13402 (N_13402,N_11520,N_10680);
or U13403 (N_13403,N_11270,N_10461);
nand U13404 (N_13404,N_11574,N_11688);
nand U13405 (N_13405,N_10572,N_11533);
nor U13406 (N_13406,N_10738,N_12410);
xnor U13407 (N_13407,N_11209,N_11342);
or U13408 (N_13408,N_10146,N_11515);
and U13409 (N_13409,N_11750,N_10486);
and U13410 (N_13410,N_12128,N_11112);
xor U13411 (N_13411,N_10526,N_12295);
xor U13412 (N_13412,N_10938,N_10416);
nor U13413 (N_13413,N_11142,N_11846);
nand U13414 (N_13414,N_11946,N_10312);
or U13415 (N_13415,N_11003,N_10505);
nor U13416 (N_13416,N_10253,N_10949);
nand U13417 (N_13417,N_11948,N_10777);
nor U13418 (N_13418,N_10671,N_10620);
or U13419 (N_13419,N_11865,N_12006);
nor U13420 (N_13420,N_10848,N_11225);
nor U13421 (N_13421,N_11615,N_10511);
and U13422 (N_13422,N_11395,N_11177);
and U13423 (N_13423,N_12123,N_11966);
and U13424 (N_13424,N_11119,N_10456);
nor U13425 (N_13425,N_12148,N_12074);
nand U13426 (N_13426,N_12141,N_10847);
and U13427 (N_13427,N_10363,N_11434);
and U13428 (N_13428,N_10144,N_10756);
nor U13429 (N_13429,N_11233,N_11912);
nor U13430 (N_13430,N_12324,N_10937);
and U13431 (N_13431,N_10366,N_11867);
or U13432 (N_13432,N_11346,N_11088);
nand U13433 (N_13433,N_10929,N_11032);
and U13434 (N_13434,N_11356,N_12127);
or U13435 (N_13435,N_12494,N_11619);
or U13436 (N_13436,N_11020,N_10759);
nand U13437 (N_13437,N_11453,N_12104);
and U13438 (N_13438,N_10911,N_11128);
xor U13439 (N_13439,N_11141,N_12489);
or U13440 (N_13440,N_11669,N_10807);
or U13441 (N_13441,N_10821,N_12339);
nand U13442 (N_13442,N_10614,N_11728);
or U13443 (N_13443,N_12356,N_11502);
and U13444 (N_13444,N_12477,N_11689);
and U13445 (N_13445,N_11569,N_10104);
or U13446 (N_13446,N_10197,N_11178);
nor U13447 (N_13447,N_11652,N_11054);
nand U13448 (N_13448,N_10697,N_11991);
or U13449 (N_13449,N_10262,N_11887);
and U13450 (N_13450,N_10690,N_12112);
and U13451 (N_13451,N_11791,N_10048);
nand U13452 (N_13452,N_11965,N_12166);
or U13453 (N_13453,N_12003,N_11785);
and U13454 (N_13454,N_11592,N_10045);
nor U13455 (N_13455,N_12370,N_11553);
or U13456 (N_13456,N_12057,N_10755);
and U13457 (N_13457,N_12142,N_12444);
nor U13458 (N_13458,N_11277,N_11160);
xor U13459 (N_13459,N_12150,N_12221);
and U13460 (N_13460,N_10999,N_11164);
and U13461 (N_13461,N_11343,N_11849);
or U13462 (N_13462,N_10204,N_12401);
and U13463 (N_13463,N_10161,N_10065);
xnor U13464 (N_13464,N_10158,N_10494);
nor U13465 (N_13465,N_11888,N_12163);
nand U13466 (N_13466,N_10961,N_10167);
nand U13467 (N_13467,N_11690,N_12364);
or U13468 (N_13468,N_10276,N_10770);
xor U13469 (N_13469,N_12330,N_12041);
and U13470 (N_13470,N_11207,N_11029);
or U13471 (N_13471,N_11829,N_10398);
or U13472 (N_13472,N_10038,N_12086);
nand U13473 (N_13473,N_11636,N_12122);
or U13474 (N_13474,N_11042,N_11710);
nor U13475 (N_13475,N_11798,N_11350);
nor U13476 (N_13476,N_10520,N_11852);
and U13477 (N_13477,N_12049,N_11939);
or U13478 (N_13478,N_11551,N_11835);
or U13479 (N_13479,N_12110,N_10116);
nor U13480 (N_13480,N_12220,N_12235);
nand U13481 (N_13481,N_11911,N_11249);
and U13482 (N_13482,N_11896,N_11389);
or U13483 (N_13483,N_11444,N_10113);
xnor U13484 (N_13484,N_10579,N_10596);
nand U13485 (N_13485,N_12170,N_10994);
nor U13486 (N_13486,N_10008,N_10808);
or U13487 (N_13487,N_12255,N_12383);
nor U13488 (N_13488,N_11370,N_11656);
or U13489 (N_13489,N_12329,N_11363);
nor U13490 (N_13490,N_10986,N_10174);
nor U13491 (N_13491,N_11906,N_12067);
nand U13492 (N_13492,N_10306,N_10368);
and U13493 (N_13493,N_10311,N_10769);
and U13494 (N_13494,N_10408,N_10047);
and U13495 (N_13495,N_10052,N_10016);
nor U13496 (N_13496,N_11111,N_10136);
nand U13497 (N_13497,N_10017,N_12176);
xor U13498 (N_13498,N_10535,N_11313);
xor U13499 (N_13499,N_12283,N_12417);
and U13500 (N_13500,N_11447,N_10182);
xnor U13501 (N_13501,N_10225,N_11061);
or U13502 (N_13502,N_10497,N_11384);
and U13503 (N_13503,N_10778,N_10753);
or U13504 (N_13504,N_10287,N_11043);
nor U13505 (N_13505,N_10551,N_11756);
and U13506 (N_13506,N_10974,N_10099);
xnor U13507 (N_13507,N_11695,N_10815);
or U13508 (N_13508,N_11634,N_11241);
nand U13509 (N_13509,N_11292,N_10220);
or U13510 (N_13510,N_12038,N_10351);
or U13511 (N_13511,N_10971,N_11460);
nand U13512 (N_13512,N_11161,N_10350);
or U13513 (N_13513,N_11023,N_12369);
nor U13514 (N_13514,N_11842,N_10709);
xor U13515 (N_13515,N_12236,N_11232);
or U13516 (N_13516,N_10564,N_10717);
xnor U13517 (N_13517,N_12451,N_11581);
and U13518 (N_13518,N_11547,N_10360);
nor U13519 (N_13519,N_10249,N_10107);
and U13520 (N_13520,N_11337,N_11713);
nor U13521 (N_13521,N_10090,N_10786);
nor U13522 (N_13522,N_10154,N_10019);
or U13523 (N_13523,N_10739,N_10216);
nor U13524 (N_13524,N_11879,N_10509);
nor U13525 (N_13525,N_11479,N_10089);
nand U13526 (N_13526,N_11452,N_12390);
and U13527 (N_13527,N_11014,N_12347);
and U13528 (N_13528,N_11604,N_12004);
xor U13529 (N_13529,N_12425,N_11836);
and U13530 (N_13530,N_12449,N_11247);
and U13531 (N_13531,N_11645,N_10850);
nand U13532 (N_13532,N_10874,N_10454);
nor U13533 (N_13533,N_11066,N_12204);
and U13534 (N_13534,N_11146,N_10814);
and U13535 (N_13535,N_10651,N_12453);
nand U13536 (N_13536,N_11565,N_10183);
xnor U13537 (N_13537,N_10284,N_12013);
and U13538 (N_13538,N_12322,N_10702);
nor U13539 (N_13539,N_10977,N_12277);
xnor U13540 (N_13540,N_12048,N_12418);
or U13541 (N_13541,N_10440,N_10567);
nand U13542 (N_13542,N_11570,N_10562);
and U13543 (N_13543,N_10644,N_11364);
nand U13544 (N_13544,N_11540,N_12183);
nand U13545 (N_13545,N_10947,N_11557);
or U13546 (N_13546,N_12462,N_10840);
or U13547 (N_13547,N_12153,N_10082);
nand U13548 (N_13548,N_12282,N_12268);
nor U13549 (N_13549,N_11317,N_11235);
and U13550 (N_13550,N_11508,N_12054);
and U13551 (N_13551,N_12007,N_11663);
nand U13552 (N_13552,N_10377,N_11637);
or U13553 (N_13553,N_10789,N_11771);
and U13554 (N_13554,N_11293,N_11107);
nand U13555 (N_13555,N_12397,N_10610);
or U13556 (N_13556,N_10541,N_11819);
and U13557 (N_13557,N_10615,N_10703);
nand U13558 (N_13558,N_10178,N_10964);
and U13559 (N_13559,N_10988,N_10080);
or U13560 (N_13560,N_10665,N_12001);
nand U13561 (N_13561,N_11859,N_10590);
or U13562 (N_13562,N_10522,N_10393);
xor U13563 (N_13563,N_12075,N_11608);
nand U13564 (N_13564,N_10566,N_10792);
or U13565 (N_13565,N_11083,N_12482);
or U13566 (N_13566,N_11012,N_12083);
nor U13567 (N_13567,N_11429,N_11082);
and U13568 (N_13568,N_12429,N_10581);
or U13569 (N_13569,N_11328,N_10820);
or U13570 (N_13570,N_10168,N_10357);
or U13571 (N_13571,N_12047,N_10384);
nor U13572 (N_13572,N_10924,N_12374);
or U13573 (N_13573,N_11691,N_10134);
nand U13574 (N_13574,N_11944,N_10985);
or U13575 (N_13575,N_11041,N_11275);
or U13576 (N_13576,N_11770,N_11021);
or U13577 (N_13577,N_10915,N_10791);
and U13578 (N_13578,N_11723,N_10296);
nor U13579 (N_13579,N_12136,N_11442);
xor U13580 (N_13580,N_10607,N_11358);
xnor U13581 (N_13581,N_11286,N_10725);
nor U13582 (N_13582,N_10263,N_11651);
nor U13583 (N_13583,N_11113,N_12365);
nand U13584 (N_13584,N_11375,N_10894);
nor U13585 (N_13585,N_11336,N_11125);
or U13586 (N_13586,N_11065,N_11648);
xor U13587 (N_13587,N_11659,N_10277);
or U13588 (N_13588,N_11310,N_11049);
xnor U13589 (N_13589,N_10836,N_11870);
and U13590 (N_13590,N_11306,N_10707);
nand U13591 (N_13591,N_10229,N_10172);
nor U13592 (N_13592,N_10120,N_11543);
nand U13593 (N_13593,N_11727,N_12042);
nor U13594 (N_13594,N_12275,N_11544);
and U13595 (N_13595,N_10570,N_12190);
nor U13596 (N_13596,N_10940,N_10025);
xor U13597 (N_13597,N_11388,N_11325);
nor U13598 (N_13598,N_12334,N_10612);
nor U13599 (N_13599,N_10372,N_12274);
nand U13600 (N_13600,N_11534,N_10571);
or U13601 (N_13601,N_11789,N_10557);
xor U13602 (N_13602,N_10242,N_10361);
nand U13603 (N_13603,N_12291,N_11603);
nor U13604 (N_13604,N_11693,N_11467);
and U13605 (N_13605,N_11752,N_12428);
or U13606 (N_13606,N_10067,N_11832);
nand U13607 (N_13607,N_11315,N_11262);
or U13608 (N_13608,N_12340,N_10701);
or U13609 (N_13609,N_11535,N_11877);
and U13610 (N_13610,N_10165,N_12371);
and U13611 (N_13611,N_11124,N_10125);
and U13612 (N_13612,N_12480,N_12257);
xnor U13613 (N_13613,N_11127,N_11668);
or U13614 (N_13614,N_10033,N_11282);
nor U13615 (N_13615,N_12025,N_10751);
or U13616 (N_13616,N_10200,N_10446);
nand U13617 (N_13617,N_11935,N_10793);
nor U13618 (N_13618,N_11300,N_10442);
or U13619 (N_13619,N_12118,N_11368);
or U13620 (N_13620,N_10682,N_10552);
nand U13621 (N_13621,N_12258,N_12225);
nor U13622 (N_13622,N_10908,N_11104);
or U13623 (N_13623,N_12064,N_11403);
or U13624 (N_13624,N_10049,N_10925);
nand U13625 (N_13625,N_11405,N_11046);
nand U13626 (N_13626,N_11985,N_12308);
xor U13627 (N_13627,N_10087,N_10137);
xnor U13628 (N_13628,N_11522,N_11957);
or U13629 (N_13629,N_10983,N_11545);
or U13630 (N_13630,N_11726,N_10856);
or U13631 (N_13631,N_11587,N_11256);
xnor U13632 (N_13632,N_11661,N_11898);
xor U13633 (N_13633,N_10809,N_11316);
nand U13634 (N_13634,N_10239,N_10326);
and U13635 (N_13635,N_10801,N_12069);
or U13636 (N_13636,N_11737,N_11678);
nand U13637 (N_13637,N_10502,N_11998);
and U13638 (N_13638,N_12247,N_11891);
nor U13639 (N_13639,N_10024,N_11952);
or U13640 (N_13640,N_11915,N_11094);
or U13641 (N_13641,N_10598,N_12321);
nand U13642 (N_13642,N_12479,N_11560);
nand U13643 (N_13643,N_11051,N_11490);
and U13644 (N_13644,N_10164,N_10621);
xnor U13645 (N_13645,N_11493,N_12023);
nand U13646 (N_13646,N_12448,N_11704);
or U13647 (N_13647,N_12491,N_11009);
nand U13648 (N_13648,N_10799,N_11758);
nand U13649 (N_13649,N_10862,N_10150);
and U13650 (N_13650,N_10039,N_12088);
nor U13651 (N_13651,N_10958,N_10490);
xnor U13652 (N_13652,N_12043,N_10909);
or U13653 (N_13653,N_12456,N_11309);
and U13654 (N_13654,N_11371,N_11774);
nor U13655 (N_13655,N_10374,N_10837);
or U13656 (N_13656,N_11053,N_11802);
nor U13657 (N_13657,N_11827,N_11224);
and U13658 (N_13658,N_12098,N_11632);
or U13659 (N_13659,N_10470,N_12191);
nor U13660 (N_13660,N_11571,N_12198);
nor U13661 (N_13661,N_10073,N_10565);
and U13662 (N_13662,N_10142,N_10723);
and U13663 (N_13663,N_10503,N_10138);
xor U13664 (N_13664,N_10282,N_10274);
and U13665 (N_13665,N_12413,N_10712);
xnor U13666 (N_13666,N_11932,N_10843);
nand U13667 (N_13667,N_10597,N_10556);
nor U13668 (N_13668,N_11163,N_11339);
or U13669 (N_13669,N_10213,N_10519);
xor U13670 (N_13670,N_12133,N_12196);
and U13671 (N_13671,N_11573,N_11174);
and U13672 (N_13672,N_10796,N_10313);
and U13673 (N_13673,N_11537,N_11237);
nor U13674 (N_13674,N_11893,N_11927);
nand U13675 (N_13675,N_11120,N_11529);
and U13676 (N_13676,N_10002,N_10568);
or U13677 (N_13677,N_10046,N_10832);
nand U13678 (N_13678,N_12376,N_10963);
xor U13679 (N_13679,N_12372,N_10462);
xor U13680 (N_13680,N_12279,N_10483);
nand U13681 (N_13681,N_12026,N_10298);
nor U13682 (N_13682,N_10156,N_11566);
nand U13683 (N_13683,N_11555,N_11757);
or U13684 (N_13684,N_11448,N_10027);
and U13685 (N_13685,N_10414,N_10482);
nor U13686 (N_13686,N_11095,N_11797);
and U13687 (N_13687,N_11227,N_10159);
nor U13688 (N_13688,N_10056,N_11485);
nand U13689 (N_13689,N_12492,N_10573);
and U13690 (N_13690,N_10289,N_11706);
or U13691 (N_13691,N_12398,N_11470);
and U13692 (N_13692,N_11969,N_11483);
nand U13693 (N_13693,N_10034,N_10001);
nand U13694 (N_13694,N_10728,N_11563);
or U13695 (N_13695,N_11696,N_10108);
and U13696 (N_13696,N_11190,N_12193);
and U13697 (N_13697,N_10459,N_10722);
nor U13698 (N_13698,N_10588,N_11474);
nand U13699 (N_13699,N_10085,N_11664);
nor U13700 (N_13700,N_11397,N_10088);
nand U13701 (N_13701,N_11438,N_11591);
nand U13702 (N_13702,N_11968,N_10889);
xor U13703 (N_13703,N_12302,N_10036);
xnor U13704 (N_13704,N_10640,N_10872);
nor U13705 (N_13705,N_10913,N_11917);
nor U13706 (N_13706,N_11699,N_12387);
or U13707 (N_13707,N_10275,N_10536);
and U13708 (N_13708,N_12430,N_11417);
or U13709 (N_13709,N_11526,N_11872);
and U13710 (N_13710,N_11993,N_11398);
nand U13711 (N_13711,N_11080,N_11201);
and U13712 (N_13712,N_12473,N_11641);
and U13713 (N_13713,N_11751,N_12077);
nor U13714 (N_13714,N_12156,N_10418);
or U13715 (N_13715,N_11382,N_11263);
nor U13716 (N_13716,N_10629,N_11305);
or U13717 (N_13717,N_11255,N_10944);
nand U13718 (N_13718,N_12109,N_11197);
and U13719 (N_13719,N_11528,N_12219);
and U13720 (N_13720,N_11561,N_12208);
and U13721 (N_13721,N_11884,N_10162);
nand U13722 (N_13722,N_11956,N_11885);
nand U13723 (N_13723,N_12289,N_12331);
xnor U13724 (N_13724,N_11108,N_10664);
nor U13725 (N_13725,N_11705,N_10241);
nand U13726 (N_13726,N_11451,N_12194);
or U13727 (N_13727,N_10752,N_12460);
or U13728 (N_13728,N_11039,N_12360);
nand U13729 (N_13729,N_10781,N_10031);
nand U13730 (N_13730,N_11700,N_11983);
or U13731 (N_13731,N_11215,N_11841);
and U13732 (N_13732,N_11955,N_10968);
nand U13733 (N_13733,N_10975,N_11701);
nor U13734 (N_13734,N_10333,N_10235);
nand U13735 (N_13735,N_11675,N_10037);
or U13736 (N_13736,N_10382,N_11072);
nand U13737 (N_13737,N_10076,N_10785);
nor U13738 (N_13738,N_10196,N_10779);
or U13739 (N_13739,N_11084,N_11861);
nand U13740 (N_13740,N_12432,N_11492);
or U13741 (N_13741,N_10341,N_11230);
nor U13742 (N_13742,N_10670,N_12062);
nand U13743 (N_13743,N_11671,N_10652);
or U13744 (N_13744,N_10825,N_11731);
and U13745 (N_13745,N_10328,N_11059);
or U13746 (N_13746,N_10389,N_11390);
nand U13747 (N_13747,N_11312,N_11531);
xnor U13748 (N_13748,N_11904,N_11843);
nand U13749 (N_13749,N_11271,N_10448);
nor U13750 (N_13750,N_11946,N_10332);
and U13751 (N_13751,N_11431,N_11343);
nand U13752 (N_13752,N_12179,N_11769);
and U13753 (N_13753,N_11790,N_12293);
and U13754 (N_13754,N_11088,N_10445);
xnor U13755 (N_13755,N_10130,N_10062);
nand U13756 (N_13756,N_12256,N_10246);
or U13757 (N_13757,N_12428,N_12416);
and U13758 (N_13758,N_10674,N_11663);
and U13759 (N_13759,N_10011,N_12228);
and U13760 (N_13760,N_10531,N_12428);
nand U13761 (N_13761,N_11960,N_11418);
and U13762 (N_13762,N_12132,N_11000);
or U13763 (N_13763,N_12328,N_11074);
or U13764 (N_13764,N_11582,N_11998);
xnor U13765 (N_13765,N_12133,N_12342);
or U13766 (N_13766,N_12420,N_11533);
or U13767 (N_13767,N_10674,N_12363);
nor U13768 (N_13768,N_11426,N_11635);
nor U13769 (N_13769,N_12478,N_10835);
and U13770 (N_13770,N_11079,N_11289);
nor U13771 (N_13771,N_11503,N_10415);
and U13772 (N_13772,N_10158,N_10478);
and U13773 (N_13773,N_11616,N_12011);
nand U13774 (N_13774,N_10937,N_11675);
nand U13775 (N_13775,N_11259,N_11488);
nor U13776 (N_13776,N_10519,N_10379);
nor U13777 (N_13777,N_10090,N_11928);
nand U13778 (N_13778,N_11232,N_10117);
and U13779 (N_13779,N_12377,N_11499);
and U13780 (N_13780,N_11960,N_10909);
and U13781 (N_13781,N_10811,N_10522);
or U13782 (N_13782,N_10364,N_12299);
and U13783 (N_13783,N_11100,N_11774);
nor U13784 (N_13784,N_10760,N_11594);
and U13785 (N_13785,N_12238,N_10456);
nor U13786 (N_13786,N_11326,N_11653);
and U13787 (N_13787,N_12188,N_10774);
and U13788 (N_13788,N_10135,N_10452);
xnor U13789 (N_13789,N_11250,N_10322);
and U13790 (N_13790,N_11528,N_11134);
nand U13791 (N_13791,N_12135,N_12071);
and U13792 (N_13792,N_10609,N_11458);
nand U13793 (N_13793,N_11385,N_11849);
and U13794 (N_13794,N_12157,N_10752);
nand U13795 (N_13795,N_10090,N_11785);
or U13796 (N_13796,N_10714,N_12189);
or U13797 (N_13797,N_10790,N_10684);
or U13798 (N_13798,N_12386,N_10131);
or U13799 (N_13799,N_12279,N_11040);
or U13800 (N_13800,N_10830,N_12313);
and U13801 (N_13801,N_11670,N_10162);
and U13802 (N_13802,N_11298,N_11908);
and U13803 (N_13803,N_10322,N_10567);
nand U13804 (N_13804,N_10267,N_10806);
and U13805 (N_13805,N_10660,N_11786);
nor U13806 (N_13806,N_10295,N_10436);
nand U13807 (N_13807,N_12473,N_11883);
or U13808 (N_13808,N_11543,N_11667);
and U13809 (N_13809,N_11146,N_10607);
and U13810 (N_13810,N_11548,N_12030);
nor U13811 (N_13811,N_12423,N_11041);
and U13812 (N_13812,N_12161,N_11507);
or U13813 (N_13813,N_10840,N_10784);
nor U13814 (N_13814,N_11405,N_10347);
and U13815 (N_13815,N_10514,N_12402);
nor U13816 (N_13816,N_10866,N_11245);
and U13817 (N_13817,N_11369,N_12336);
and U13818 (N_13818,N_12449,N_11843);
nand U13819 (N_13819,N_10710,N_11037);
or U13820 (N_13820,N_10565,N_12169);
xnor U13821 (N_13821,N_11973,N_10634);
nor U13822 (N_13822,N_11833,N_11274);
or U13823 (N_13823,N_10866,N_11863);
nand U13824 (N_13824,N_10947,N_11943);
nor U13825 (N_13825,N_11224,N_10879);
and U13826 (N_13826,N_10096,N_11886);
or U13827 (N_13827,N_10402,N_10502);
or U13828 (N_13828,N_11954,N_10270);
nand U13829 (N_13829,N_10994,N_11357);
and U13830 (N_13830,N_11759,N_12105);
and U13831 (N_13831,N_11116,N_11248);
nor U13832 (N_13832,N_11819,N_11139);
xnor U13833 (N_13833,N_10579,N_10175);
nor U13834 (N_13834,N_12308,N_10951);
and U13835 (N_13835,N_12477,N_11763);
nor U13836 (N_13836,N_10205,N_11020);
and U13837 (N_13837,N_11790,N_10625);
nand U13838 (N_13838,N_10266,N_11087);
nand U13839 (N_13839,N_10909,N_10161);
nand U13840 (N_13840,N_11367,N_11688);
nor U13841 (N_13841,N_10182,N_10634);
nor U13842 (N_13842,N_11803,N_11445);
nor U13843 (N_13843,N_10711,N_10084);
and U13844 (N_13844,N_10466,N_12168);
and U13845 (N_13845,N_11707,N_12333);
or U13846 (N_13846,N_10379,N_10032);
or U13847 (N_13847,N_12230,N_10336);
nand U13848 (N_13848,N_10020,N_11211);
and U13849 (N_13849,N_10919,N_10187);
and U13850 (N_13850,N_10012,N_10634);
nand U13851 (N_13851,N_11883,N_10532);
nand U13852 (N_13852,N_11277,N_10573);
or U13853 (N_13853,N_10719,N_10912);
xnor U13854 (N_13854,N_11479,N_12252);
nand U13855 (N_13855,N_11713,N_10140);
nor U13856 (N_13856,N_11331,N_12328);
nor U13857 (N_13857,N_10022,N_10609);
or U13858 (N_13858,N_12467,N_12286);
or U13859 (N_13859,N_11938,N_12322);
nor U13860 (N_13860,N_10379,N_10435);
and U13861 (N_13861,N_10685,N_10979);
nand U13862 (N_13862,N_10593,N_10951);
or U13863 (N_13863,N_10352,N_11998);
and U13864 (N_13864,N_11401,N_10588);
nand U13865 (N_13865,N_10501,N_12244);
xnor U13866 (N_13866,N_11923,N_11735);
and U13867 (N_13867,N_11576,N_10671);
nor U13868 (N_13868,N_10390,N_11265);
nand U13869 (N_13869,N_12075,N_12415);
nand U13870 (N_13870,N_10427,N_10068);
nor U13871 (N_13871,N_11518,N_10087);
or U13872 (N_13872,N_12152,N_12089);
nor U13873 (N_13873,N_10444,N_10319);
nor U13874 (N_13874,N_12020,N_11015);
nor U13875 (N_13875,N_10631,N_11081);
nand U13876 (N_13876,N_10429,N_11755);
and U13877 (N_13877,N_12009,N_11171);
nor U13878 (N_13878,N_11071,N_11441);
and U13879 (N_13879,N_10859,N_12453);
nand U13880 (N_13880,N_12114,N_10555);
nand U13881 (N_13881,N_11242,N_10192);
nor U13882 (N_13882,N_10439,N_12084);
nand U13883 (N_13883,N_10275,N_10099);
and U13884 (N_13884,N_12290,N_11002);
nor U13885 (N_13885,N_10703,N_11083);
or U13886 (N_13886,N_10752,N_11369);
nor U13887 (N_13887,N_12064,N_12469);
and U13888 (N_13888,N_10725,N_11208);
nor U13889 (N_13889,N_10803,N_10617);
nand U13890 (N_13890,N_11106,N_12046);
or U13891 (N_13891,N_12099,N_11357);
nand U13892 (N_13892,N_12296,N_10193);
or U13893 (N_13893,N_10744,N_10218);
nand U13894 (N_13894,N_11559,N_10817);
nor U13895 (N_13895,N_12438,N_11855);
nor U13896 (N_13896,N_10246,N_11679);
and U13897 (N_13897,N_11874,N_11890);
nand U13898 (N_13898,N_11597,N_10432);
nor U13899 (N_13899,N_10083,N_11044);
nor U13900 (N_13900,N_11335,N_10376);
or U13901 (N_13901,N_10481,N_11016);
or U13902 (N_13902,N_10639,N_10221);
nand U13903 (N_13903,N_10361,N_11001);
nor U13904 (N_13904,N_12254,N_10434);
or U13905 (N_13905,N_11611,N_11606);
or U13906 (N_13906,N_11250,N_10891);
nor U13907 (N_13907,N_12209,N_10167);
nor U13908 (N_13908,N_11916,N_10908);
nand U13909 (N_13909,N_11941,N_10532);
and U13910 (N_13910,N_10170,N_11929);
nand U13911 (N_13911,N_11188,N_11059);
and U13912 (N_13912,N_12315,N_10124);
nor U13913 (N_13913,N_10139,N_10384);
or U13914 (N_13914,N_12416,N_10104);
xnor U13915 (N_13915,N_11488,N_11377);
nand U13916 (N_13916,N_10819,N_12434);
and U13917 (N_13917,N_10793,N_11790);
nand U13918 (N_13918,N_10049,N_10654);
nand U13919 (N_13919,N_10598,N_10896);
nand U13920 (N_13920,N_12033,N_11685);
nand U13921 (N_13921,N_10553,N_10824);
nor U13922 (N_13922,N_10581,N_12138);
xnor U13923 (N_13923,N_10376,N_10078);
or U13924 (N_13924,N_12442,N_10909);
and U13925 (N_13925,N_11275,N_10094);
and U13926 (N_13926,N_12173,N_12370);
and U13927 (N_13927,N_10911,N_12366);
or U13928 (N_13928,N_11388,N_10157);
nand U13929 (N_13929,N_11814,N_11600);
and U13930 (N_13930,N_10409,N_10088);
nor U13931 (N_13931,N_10837,N_11298);
and U13932 (N_13932,N_11174,N_10876);
or U13933 (N_13933,N_10099,N_11159);
nor U13934 (N_13934,N_11584,N_11064);
nand U13935 (N_13935,N_11089,N_11333);
nand U13936 (N_13936,N_12238,N_11747);
nor U13937 (N_13937,N_12434,N_11445);
or U13938 (N_13938,N_11932,N_11852);
nand U13939 (N_13939,N_11028,N_10584);
xor U13940 (N_13940,N_10915,N_11888);
or U13941 (N_13941,N_11151,N_10531);
nand U13942 (N_13942,N_11578,N_11522);
nor U13943 (N_13943,N_10634,N_11301);
xnor U13944 (N_13944,N_12134,N_11531);
nor U13945 (N_13945,N_10571,N_11337);
and U13946 (N_13946,N_10080,N_10105);
or U13947 (N_13947,N_12367,N_11933);
and U13948 (N_13948,N_11064,N_10354);
nor U13949 (N_13949,N_10439,N_12211);
nand U13950 (N_13950,N_12003,N_11776);
nand U13951 (N_13951,N_11542,N_11868);
nor U13952 (N_13952,N_11756,N_11443);
nor U13953 (N_13953,N_12340,N_10889);
nand U13954 (N_13954,N_11578,N_10473);
xnor U13955 (N_13955,N_10042,N_10725);
xor U13956 (N_13956,N_11040,N_12275);
or U13957 (N_13957,N_12006,N_11506);
nand U13958 (N_13958,N_11215,N_11994);
and U13959 (N_13959,N_11440,N_10380);
nor U13960 (N_13960,N_11682,N_10382);
and U13961 (N_13961,N_10583,N_11867);
or U13962 (N_13962,N_12126,N_10701);
and U13963 (N_13963,N_11022,N_11841);
and U13964 (N_13964,N_12133,N_11100);
xnor U13965 (N_13965,N_12263,N_10271);
or U13966 (N_13966,N_12289,N_10791);
nand U13967 (N_13967,N_11029,N_10318);
nand U13968 (N_13968,N_11920,N_11344);
and U13969 (N_13969,N_11004,N_12083);
or U13970 (N_13970,N_11409,N_11970);
nand U13971 (N_13971,N_12354,N_11141);
nand U13972 (N_13972,N_11900,N_10370);
nor U13973 (N_13973,N_10142,N_12161);
or U13974 (N_13974,N_12172,N_10719);
and U13975 (N_13975,N_11491,N_11317);
and U13976 (N_13976,N_11068,N_12298);
xor U13977 (N_13977,N_10187,N_10544);
xor U13978 (N_13978,N_10695,N_12051);
nor U13979 (N_13979,N_12433,N_10301);
or U13980 (N_13980,N_10265,N_12118);
nor U13981 (N_13981,N_10965,N_12307);
or U13982 (N_13982,N_11658,N_10022);
or U13983 (N_13983,N_12178,N_11695);
or U13984 (N_13984,N_12390,N_11576);
and U13985 (N_13985,N_11102,N_11899);
or U13986 (N_13986,N_11219,N_10447);
or U13987 (N_13987,N_10244,N_12325);
or U13988 (N_13988,N_10109,N_10185);
or U13989 (N_13989,N_12293,N_11922);
nand U13990 (N_13990,N_10501,N_11425);
nand U13991 (N_13991,N_11795,N_10794);
nand U13992 (N_13992,N_10571,N_10187);
nand U13993 (N_13993,N_11489,N_10378);
or U13994 (N_13994,N_12350,N_12077);
and U13995 (N_13995,N_11714,N_11613);
or U13996 (N_13996,N_11579,N_12058);
nor U13997 (N_13997,N_11486,N_11123);
nor U13998 (N_13998,N_12487,N_11503);
and U13999 (N_13999,N_11855,N_11081);
nor U14000 (N_14000,N_10942,N_12207);
and U14001 (N_14001,N_10313,N_11846);
nor U14002 (N_14002,N_11740,N_11339);
nand U14003 (N_14003,N_12166,N_12182);
nand U14004 (N_14004,N_10615,N_11629);
nor U14005 (N_14005,N_11748,N_10764);
nand U14006 (N_14006,N_11539,N_10957);
nand U14007 (N_14007,N_11276,N_11086);
xor U14008 (N_14008,N_10352,N_10223);
or U14009 (N_14009,N_10656,N_10435);
and U14010 (N_14010,N_11664,N_10087);
nand U14011 (N_14011,N_10661,N_12126);
nor U14012 (N_14012,N_10738,N_10552);
and U14013 (N_14013,N_10538,N_12328);
and U14014 (N_14014,N_11732,N_10967);
nand U14015 (N_14015,N_11851,N_10808);
xnor U14016 (N_14016,N_10645,N_12467);
or U14017 (N_14017,N_11329,N_10636);
and U14018 (N_14018,N_10020,N_11067);
and U14019 (N_14019,N_11123,N_11485);
nor U14020 (N_14020,N_10176,N_11076);
xnor U14021 (N_14021,N_11481,N_10931);
and U14022 (N_14022,N_11529,N_11761);
or U14023 (N_14023,N_11801,N_12411);
xnor U14024 (N_14024,N_11038,N_11172);
nand U14025 (N_14025,N_11759,N_11130);
or U14026 (N_14026,N_12291,N_11059);
and U14027 (N_14027,N_11641,N_10588);
or U14028 (N_14028,N_10290,N_11245);
nand U14029 (N_14029,N_10175,N_12112);
and U14030 (N_14030,N_10304,N_12316);
nand U14031 (N_14031,N_11439,N_10180);
nor U14032 (N_14032,N_12472,N_11756);
nor U14033 (N_14033,N_11624,N_10137);
nand U14034 (N_14034,N_11024,N_10165);
or U14035 (N_14035,N_11780,N_12442);
nand U14036 (N_14036,N_10606,N_10416);
xnor U14037 (N_14037,N_11447,N_11771);
nand U14038 (N_14038,N_10799,N_11302);
or U14039 (N_14039,N_11485,N_10490);
nand U14040 (N_14040,N_10984,N_12365);
or U14041 (N_14041,N_12142,N_10941);
nor U14042 (N_14042,N_10956,N_10810);
and U14043 (N_14043,N_11777,N_10996);
nand U14044 (N_14044,N_10871,N_10395);
xor U14045 (N_14045,N_11812,N_10107);
nor U14046 (N_14046,N_12490,N_11177);
nand U14047 (N_14047,N_11532,N_10894);
or U14048 (N_14048,N_11320,N_12106);
or U14049 (N_14049,N_11808,N_11707);
or U14050 (N_14050,N_12004,N_12140);
xnor U14051 (N_14051,N_11928,N_11414);
and U14052 (N_14052,N_12270,N_11593);
xor U14053 (N_14053,N_10984,N_10659);
nand U14054 (N_14054,N_11459,N_11965);
nor U14055 (N_14055,N_11471,N_11650);
nand U14056 (N_14056,N_12362,N_11780);
nand U14057 (N_14057,N_10115,N_11699);
xor U14058 (N_14058,N_11121,N_11777);
nand U14059 (N_14059,N_11344,N_11761);
or U14060 (N_14060,N_11845,N_10061);
nor U14061 (N_14061,N_12389,N_11308);
or U14062 (N_14062,N_11910,N_12126);
and U14063 (N_14063,N_12205,N_12114);
nand U14064 (N_14064,N_10328,N_11554);
and U14065 (N_14065,N_10354,N_11631);
and U14066 (N_14066,N_11093,N_11443);
nand U14067 (N_14067,N_11053,N_10941);
xnor U14068 (N_14068,N_10753,N_11755);
and U14069 (N_14069,N_12435,N_11681);
and U14070 (N_14070,N_10664,N_11549);
or U14071 (N_14071,N_10840,N_11626);
and U14072 (N_14072,N_11750,N_11979);
nand U14073 (N_14073,N_11533,N_12237);
or U14074 (N_14074,N_10957,N_10008);
and U14075 (N_14075,N_10075,N_11655);
and U14076 (N_14076,N_11233,N_10777);
nand U14077 (N_14077,N_11646,N_11279);
nand U14078 (N_14078,N_11048,N_10135);
nor U14079 (N_14079,N_11044,N_12075);
nor U14080 (N_14080,N_10454,N_10811);
and U14081 (N_14081,N_12231,N_11143);
and U14082 (N_14082,N_12152,N_11193);
nor U14083 (N_14083,N_11785,N_10065);
and U14084 (N_14084,N_10910,N_10077);
or U14085 (N_14085,N_10916,N_11267);
nor U14086 (N_14086,N_10759,N_10637);
or U14087 (N_14087,N_10310,N_11840);
nor U14088 (N_14088,N_10582,N_12129);
nand U14089 (N_14089,N_11958,N_10071);
or U14090 (N_14090,N_12184,N_11026);
nor U14091 (N_14091,N_12073,N_10416);
or U14092 (N_14092,N_12130,N_10281);
xor U14093 (N_14093,N_12073,N_11745);
or U14094 (N_14094,N_11394,N_12443);
nor U14095 (N_14095,N_10874,N_11044);
or U14096 (N_14096,N_10909,N_10930);
xor U14097 (N_14097,N_11033,N_10742);
nor U14098 (N_14098,N_10775,N_12201);
nor U14099 (N_14099,N_10503,N_11754);
and U14100 (N_14100,N_12004,N_12169);
or U14101 (N_14101,N_10691,N_10867);
and U14102 (N_14102,N_11076,N_11263);
and U14103 (N_14103,N_10526,N_10576);
nand U14104 (N_14104,N_10495,N_11594);
xnor U14105 (N_14105,N_10857,N_11931);
and U14106 (N_14106,N_10886,N_11292);
or U14107 (N_14107,N_10090,N_11211);
nand U14108 (N_14108,N_10870,N_11833);
and U14109 (N_14109,N_12304,N_11741);
or U14110 (N_14110,N_11313,N_12479);
or U14111 (N_14111,N_11135,N_11968);
nand U14112 (N_14112,N_10801,N_10019);
or U14113 (N_14113,N_12450,N_11174);
or U14114 (N_14114,N_11706,N_12121);
or U14115 (N_14115,N_10405,N_10331);
or U14116 (N_14116,N_11412,N_10376);
nand U14117 (N_14117,N_11959,N_11086);
nand U14118 (N_14118,N_12375,N_12205);
nor U14119 (N_14119,N_10075,N_11542);
xnor U14120 (N_14120,N_10300,N_10578);
or U14121 (N_14121,N_10318,N_10233);
xnor U14122 (N_14122,N_11249,N_10854);
xor U14123 (N_14123,N_10052,N_12000);
or U14124 (N_14124,N_11066,N_10319);
xnor U14125 (N_14125,N_10292,N_10707);
nor U14126 (N_14126,N_10947,N_11628);
nor U14127 (N_14127,N_11356,N_10945);
or U14128 (N_14128,N_11440,N_11836);
nor U14129 (N_14129,N_10307,N_11381);
xnor U14130 (N_14130,N_10331,N_11828);
or U14131 (N_14131,N_10533,N_11440);
xnor U14132 (N_14132,N_10071,N_12341);
or U14133 (N_14133,N_11514,N_11772);
xor U14134 (N_14134,N_11755,N_12252);
or U14135 (N_14135,N_11091,N_11779);
nand U14136 (N_14136,N_11865,N_12489);
or U14137 (N_14137,N_12071,N_11477);
nand U14138 (N_14138,N_12236,N_11201);
or U14139 (N_14139,N_10426,N_11819);
and U14140 (N_14140,N_10023,N_11105);
nand U14141 (N_14141,N_10863,N_11415);
nand U14142 (N_14142,N_10216,N_11282);
and U14143 (N_14143,N_11908,N_11956);
or U14144 (N_14144,N_11270,N_10766);
and U14145 (N_14145,N_11555,N_10142);
and U14146 (N_14146,N_11867,N_10351);
and U14147 (N_14147,N_11837,N_11198);
nand U14148 (N_14148,N_10440,N_12319);
or U14149 (N_14149,N_11870,N_12160);
nor U14150 (N_14150,N_11783,N_10995);
nand U14151 (N_14151,N_11434,N_10387);
xor U14152 (N_14152,N_10373,N_10056);
or U14153 (N_14153,N_10327,N_10143);
nor U14154 (N_14154,N_10040,N_11802);
xnor U14155 (N_14155,N_11396,N_10134);
nand U14156 (N_14156,N_11825,N_12376);
and U14157 (N_14157,N_11385,N_11522);
or U14158 (N_14158,N_10638,N_11838);
or U14159 (N_14159,N_11348,N_10014);
nor U14160 (N_14160,N_11837,N_11303);
nand U14161 (N_14161,N_11641,N_12148);
and U14162 (N_14162,N_10100,N_10345);
nand U14163 (N_14163,N_10957,N_12212);
or U14164 (N_14164,N_12067,N_11346);
xnor U14165 (N_14165,N_11255,N_11888);
nor U14166 (N_14166,N_12067,N_10085);
or U14167 (N_14167,N_11092,N_12417);
or U14168 (N_14168,N_12346,N_10143);
nor U14169 (N_14169,N_10756,N_12431);
and U14170 (N_14170,N_11224,N_11261);
nand U14171 (N_14171,N_11620,N_10678);
nor U14172 (N_14172,N_12249,N_10058);
or U14173 (N_14173,N_10764,N_11747);
and U14174 (N_14174,N_11794,N_12074);
nor U14175 (N_14175,N_10030,N_11400);
nor U14176 (N_14176,N_12325,N_12109);
nor U14177 (N_14177,N_10257,N_11270);
nor U14178 (N_14178,N_11962,N_10420);
or U14179 (N_14179,N_10410,N_10304);
and U14180 (N_14180,N_11056,N_10527);
or U14181 (N_14181,N_12478,N_10729);
or U14182 (N_14182,N_12141,N_12466);
nand U14183 (N_14183,N_10586,N_11447);
nor U14184 (N_14184,N_11967,N_10227);
nand U14185 (N_14185,N_11003,N_12441);
and U14186 (N_14186,N_11621,N_10611);
nor U14187 (N_14187,N_12093,N_10680);
xnor U14188 (N_14188,N_11926,N_11810);
nor U14189 (N_14189,N_12192,N_12466);
nor U14190 (N_14190,N_11955,N_10608);
nor U14191 (N_14191,N_11709,N_12023);
and U14192 (N_14192,N_10957,N_11148);
nand U14193 (N_14193,N_12099,N_11591);
nor U14194 (N_14194,N_11879,N_12178);
nand U14195 (N_14195,N_11531,N_10181);
and U14196 (N_14196,N_12159,N_11442);
or U14197 (N_14197,N_11154,N_12014);
and U14198 (N_14198,N_10138,N_12269);
and U14199 (N_14199,N_12114,N_10093);
nand U14200 (N_14200,N_11230,N_12356);
nand U14201 (N_14201,N_10383,N_11219);
nor U14202 (N_14202,N_11844,N_11016);
xor U14203 (N_14203,N_11284,N_10108);
or U14204 (N_14204,N_12280,N_11558);
and U14205 (N_14205,N_11181,N_10735);
nor U14206 (N_14206,N_11732,N_10955);
nor U14207 (N_14207,N_11958,N_11720);
nand U14208 (N_14208,N_11805,N_12004);
nor U14209 (N_14209,N_11247,N_10128);
or U14210 (N_14210,N_12134,N_10757);
or U14211 (N_14211,N_11955,N_11527);
and U14212 (N_14212,N_12465,N_11530);
xnor U14213 (N_14213,N_10941,N_12491);
or U14214 (N_14214,N_11764,N_12094);
xor U14215 (N_14215,N_12071,N_10620);
xor U14216 (N_14216,N_12232,N_10789);
nor U14217 (N_14217,N_12281,N_11530);
and U14218 (N_14218,N_11196,N_11928);
nand U14219 (N_14219,N_10832,N_11838);
and U14220 (N_14220,N_10981,N_11648);
or U14221 (N_14221,N_10954,N_12069);
nor U14222 (N_14222,N_11975,N_10198);
nand U14223 (N_14223,N_10013,N_10873);
nand U14224 (N_14224,N_11133,N_10857);
nor U14225 (N_14225,N_10354,N_10153);
nor U14226 (N_14226,N_10337,N_11211);
nor U14227 (N_14227,N_12185,N_11724);
nor U14228 (N_14228,N_12144,N_10394);
or U14229 (N_14229,N_12440,N_10212);
and U14230 (N_14230,N_11344,N_11553);
or U14231 (N_14231,N_11103,N_12155);
or U14232 (N_14232,N_10496,N_10517);
or U14233 (N_14233,N_10786,N_11469);
nor U14234 (N_14234,N_10776,N_10119);
xnor U14235 (N_14235,N_10836,N_12274);
and U14236 (N_14236,N_11741,N_10729);
and U14237 (N_14237,N_12414,N_10379);
and U14238 (N_14238,N_11151,N_12413);
and U14239 (N_14239,N_11845,N_10462);
and U14240 (N_14240,N_11540,N_10063);
nand U14241 (N_14241,N_12154,N_12112);
and U14242 (N_14242,N_11606,N_10767);
and U14243 (N_14243,N_10870,N_12233);
xnor U14244 (N_14244,N_10076,N_11814);
or U14245 (N_14245,N_11968,N_10995);
and U14246 (N_14246,N_11808,N_11116);
nand U14247 (N_14247,N_10598,N_11226);
xnor U14248 (N_14248,N_10397,N_11610);
nor U14249 (N_14249,N_12035,N_10337);
nor U14250 (N_14250,N_11412,N_11129);
nand U14251 (N_14251,N_12377,N_10972);
nor U14252 (N_14252,N_10999,N_11567);
or U14253 (N_14253,N_11429,N_11011);
and U14254 (N_14254,N_11717,N_10379);
or U14255 (N_14255,N_11632,N_12110);
and U14256 (N_14256,N_11106,N_12257);
nor U14257 (N_14257,N_11507,N_11996);
nor U14258 (N_14258,N_10712,N_10816);
and U14259 (N_14259,N_10040,N_12310);
nand U14260 (N_14260,N_10021,N_11042);
nor U14261 (N_14261,N_10727,N_11192);
or U14262 (N_14262,N_11908,N_11703);
xor U14263 (N_14263,N_10352,N_11299);
and U14264 (N_14264,N_10339,N_11525);
nand U14265 (N_14265,N_12389,N_10737);
nor U14266 (N_14266,N_11384,N_11916);
nor U14267 (N_14267,N_10903,N_10221);
or U14268 (N_14268,N_10676,N_10819);
nand U14269 (N_14269,N_10514,N_11886);
or U14270 (N_14270,N_10279,N_11613);
xnor U14271 (N_14271,N_12499,N_11253);
and U14272 (N_14272,N_10468,N_10651);
nor U14273 (N_14273,N_11650,N_10978);
nor U14274 (N_14274,N_10583,N_11409);
xnor U14275 (N_14275,N_11327,N_11747);
or U14276 (N_14276,N_12112,N_11839);
or U14277 (N_14277,N_11741,N_11825);
nor U14278 (N_14278,N_10899,N_10785);
xnor U14279 (N_14279,N_10476,N_10686);
or U14280 (N_14280,N_10109,N_12425);
and U14281 (N_14281,N_11655,N_12411);
xnor U14282 (N_14282,N_10775,N_11957);
nand U14283 (N_14283,N_12035,N_12047);
nand U14284 (N_14284,N_10868,N_11782);
or U14285 (N_14285,N_10773,N_11453);
nand U14286 (N_14286,N_11019,N_10795);
or U14287 (N_14287,N_12464,N_10071);
xnor U14288 (N_14288,N_10774,N_11647);
nand U14289 (N_14289,N_12441,N_11584);
and U14290 (N_14290,N_10388,N_10321);
and U14291 (N_14291,N_11126,N_12054);
nor U14292 (N_14292,N_10139,N_11684);
nand U14293 (N_14293,N_10342,N_11067);
or U14294 (N_14294,N_10414,N_12350);
and U14295 (N_14295,N_12301,N_10481);
or U14296 (N_14296,N_11738,N_10378);
or U14297 (N_14297,N_11796,N_11934);
nor U14298 (N_14298,N_10791,N_11854);
or U14299 (N_14299,N_12044,N_10633);
nand U14300 (N_14300,N_10632,N_10882);
nor U14301 (N_14301,N_12351,N_11113);
and U14302 (N_14302,N_12495,N_10397);
xor U14303 (N_14303,N_11524,N_12175);
and U14304 (N_14304,N_11147,N_11000);
nor U14305 (N_14305,N_11803,N_11604);
or U14306 (N_14306,N_11381,N_10114);
xnor U14307 (N_14307,N_10509,N_12067);
nor U14308 (N_14308,N_12193,N_10686);
or U14309 (N_14309,N_12238,N_11268);
nor U14310 (N_14310,N_10248,N_10973);
or U14311 (N_14311,N_11469,N_10443);
nand U14312 (N_14312,N_11851,N_12004);
or U14313 (N_14313,N_10364,N_10296);
nor U14314 (N_14314,N_10797,N_11064);
and U14315 (N_14315,N_11558,N_10462);
nor U14316 (N_14316,N_12452,N_11753);
and U14317 (N_14317,N_10055,N_10374);
and U14318 (N_14318,N_11150,N_10417);
nand U14319 (N_14319,N_10301,N_11843);
nand U14320 (N_14320,N_12426,N_11485);
or U14321 (N_14321,N_10504,N_12108);
nand U14322 (N_14322,N_12292,N_11123);
and U14323 (N_14323,N_11195,N_10629);
or U14324 (N_14324,N_10030,N_10875);
and U14325 (N_14325,N_12196,N_10177);
xor U14326 (N_14326,N_11321,N_12140);
and U14327 (N_14327,N_10058,N_12216);
nor U14328 (N_14328,N_11188,N_11413);
xor U14329 (N_14329,N_10974,N_12098);
or U14330 (N_14330,N_11404,N_10177);
nor U14331 (N_14331,N_10730,N_10754);
nor U14332 (N_14332,N_11300,N_10250);
and U14333 (N_14333,N_10440,N_12216);
xor U14334 (N_14334,N_10491,N_12236);
nand U14335 (N_14335,N_10363,N_12492);
nor U14336 (N_14336,N_11227,N_11362);
or U14337 (N_14337,N_11983,N_10193);
or U14338 (N_14338,N_10783,N_10454);
xor U14339 (N_14339,N_11072,N_10068);
and U14340 (N_14340,N_10311,N_11170);
and U14341 (N_14341,N_11948,N_10782);
nor U14342 (N_14342,N_11228,N_10608);
nor U14343 (N_14343,N_10782,N_11765);
and U14344 (N_14344,N_12274,N_10056);
and U14345 (N_14345,N_12393,N_10598);
nand U14346 (N_14346,N_11725,N_10657);
and U14347 (N_14347,N_12230,N_10506);
nor U14348 (N_14348,N_10248,N_11309);
and U14349 (N_14349,N_11434,N_10286);
nor U14350 (N_14350,N_11709,N_11020);
nor U14351 (N_14351,N_11717,N_10169);
and U14352 (N_14352,N_10031,N_11098);
or U14353 (N_14353,N_10529,N_12170);
xor U14354 (N_14354,N_12270,N_11339);
or U14355 (N_14355,N_11671,N_12206);
and U14356 (N_14356,N_12212,N_12443);
nor U14357 (N_14357,N_10641,N_12453);
xor U14358 (N_14358,N_10839,N_10388);
nand U14359 (N_14359,N_12242,N_10118);
and U14360 (N_14360,N_11900,N_12304);
nand U14361 (N_14361,N_10149,N_11686);
nor U14362 (N_14362,N_11430,N_11224);
and U14363 (N_14363,N_12322,N_10079);
xnor U14364 (N_14364,N_12091,N_11053);
nand U14365 (N_14365,N_10114,N_10197);
and U14366 (N_14366,N_10212,N_12396);
or U14367 (N_14367,N_11791,N_10464);
nor U14368 (N_14368,N_11228,N_10926);
nand U14369 (N_14369,N_10163,N_11633);
and U14370 (N_14370,N_10150,N_12430);
nor U14371 (N_14371,N_10558,N_12164);
nor U14372 (N_14372,N_11024,N_10366);
nand U14373 (N_14373,N_10190,N_10159);
or U14374 (N_14374,N_11852,N_11103);
nand U14375 (N_14375,N_11818,N_11730);
nand U14376 (N_14376,N_11794,N_10381);
and U14377 (N_14377,N_10470,N_10492);
nor U14378 (N_14378,N_10748,N_10741);
or U14379 (N_14379,N_12371,N_10672);
and U14380 (N_14380,N_12490,N_10060);
nor U14381 (N_14381,N_10693,N_12155);
nor U14382 (N_14382,N_12466,N_11100);
nor U14383 (N_14383,N_10639,N_11596);
and U14384 (N_14384,N_10749,N_12394);
and U14385 (N_14385,N_11886,N_10470);
nand U14386 (N_14386,N_11237,N_12452);
or U14387 (N_14387,N_11271,N_11672);
or U14388 (N_14388,N_11871,N_10815);
nor U14389 (N_14389,N_10388,N_10561);
xor U14390 (N_14390,N_10923,N_11837);
or U14391 (N_14391,N_11111,N_10002);
nand U14392 (N_14392,N_10074,N_10540);
nor U14393 (N_14393,N_12189,N_10843);
nor U14394 (N_14394,N_12465,N_10078);
or U14395 (N_14395,N_10265,N_12112);
nor U14396 (N_14396,N_11392,N_10078);
and U14397 (N_14397,N_12082,N_10207);
or U14398 (N_14398,N_10622,N_12137);
or U14399 (N_14399,N_10852,N_10698);
and U14400 (N_14400,N_11939,N_10293);
nor U14401 (N_14401,N_10364,N_11424);
or U14402 (N_14402,N_10733,N_10307);
or U14403 (N_14403,N_12377,N_12216);
or U14404 (N_14404,N_10446,N_12021);
nand U14405 (N_14405,N_11639,N_10052);
and U14406 (N_14406,N_10945,N_11545);
nor U14407 (N_14407,N_11354,N_12063);
or U14408 (N_14408,N_11971,N_12131);
or U14409 (N_14409,N_12051,N_11217);
nor U14410 (N_14410,N_12436,N_10074);
nor U14411 (N_14411,N_10533,N_10071);
nor U14412 (N_14412,N_11979,N_11705);
nand U14413 (N_14413,N_10621,N_10447);
and U14414 (N_14414,N_10797,N_11032);
nor U14415 (N_14415,N_10173,N_11856);
nor U14416 (N_14416,N_11194,N_10066);
nand U14417 (N_14417,N_12060,N_11265);
nand U14418 (N_14418,N_11627,N_10666);
nand U14419 (N_14419,N_10251,N_10848);
and U14420 (N_14420,N_10134,N_12132);
or U14421 (N_14421,N_10459,N_12123);
and U14422 (N_14422,N_10205,N_11279);
and U14423 (N_14423,N_10328,N_10929);
nor U14424 (N_14424,N_10205,N_11503);
nand U14425 (N_14425,N_10533,N_10164);
or U14426 (N_14426,N_11118,N_12383);
or U14427 (N_14427,N_11715,N_11693);
nor U14428 (N_14428,N_10371,N_11854);
and U14429 (N_14429,N_12006,N_10954);
nand U14430 (N_14430,N_11622,N_12152);
or U14431 (N_14431,N_10917,N_11618);
nor U14432 (N_14432,N_12149,N_11586);
or U14433 (N_14433,N_12453,N_10781);
nor U14434 (N_14434,N_10329,N_10898);
xor U14435 (N_14435,N_10559,N_11568);
nor U14436 (N_14436,N_10262,N_11529);
nand U14437 (N_14437,N_11417,N_10749);
nor U14438 (N_14438,N_10526,N_10088);
or U14439 (N_14439,N_12047,N_11632);
nor U14440 (N_14440,N_12069,N_12225);
nor U14441 (N_14441,N_12385,N_12078);
nor U14442 (N_14442,N_11979,N_11869);
nor U14443 (N_14443,N_11076,N_10399);
nand U14444 (N_14444,N_10831,N_10757);
or U14445 (N_14445,N_11592,N_10799);
or U14446 (N_14446,N_12408,N_10752);
nand U14447 (N_14447,N_10017,N_10518);
and U14448 (N_14448,N_11254,N_12011);
and U14449 (N_14449,N_11726,N_10492);
or U14450 (N_14450,N_10985,N_11886);
nand U14451 (N_14451,N_11539,N_10813);
or U14452 (N_14452,N_10036,N_12070);
and U14453 (N_14453,N_11450,N_11881);
nor U14454 (N_14454,N_11738,N_10617);
nor U14455 (N_14455,N_12264,N_10431);
or U14456 (N_14456,N_11816,N_11310);
nor U14457 (N_14457,N_10950,N_10132);
or U14458 (N_14458,N_11317,N_11250);
or U14459 (N_14459,N_11086,N_12140);
or U14460 (N_14460,N_10548,N_11654);
nand U14461 (N_14461,N_11714,N_12099);
or U14462 (N_14462,N_10454,N_10527);
nand U14463 (N_14463,N_10543,N_11885);
nand U14464 (N_14464,N_10460,N_10124);
and U14465 (N_14465,N_10984,N_10824);
xor U14466 (N_14466,N_10102,N_10422);
nor U14467 (N_14467,N_10155,N_10100);
nor U14468 (N_14468,N_11129,N_11750);
or U14469 (N_14469,N_11746,N_10304);
and U14470 (N_14470,N_12008,N_12305);
and U14471 (N_14471,N_10461,N_11878);
nand U14472 (N_14472,N_11270,N_11918);
or U14473 (N_14473,N_11917,N_10643);
or U14474 (N_14474,N_11496,N_11001);
nand U14475 (N_14475,N_10923,N_11112);
nor U14476 (N_14476,N_11541,N_11306);
and U14477 (N_14477,N_11282,N_10655);
xnor U14478 (N_14478,N_11092,N_10239);
xor U14479 (N_14479,N_12127,N_10699);
nor U14480 (N_14480,N_11308,N_10769);
nor U14481 (N_14481,N_12458,N_12207);
nand U14482 (N_14482,N_11689,N_10431);
nor U14483 (N_14483,N_10115,N_11710);
nand U14484 (N_14484,N_10456,N_10062);
nor U14485 (N_14485,N_11970,N_11615);
nor U14486 (N_14486,N_11190,N_11958);
xor U14487 (N_14487,N_10168,N_11027);
and U14488 (N_14488,N_11514,N_11862);
or U14489 (N_14489,N_11721,N_11944);
nor U14490 (N_14490,N_12311,N_10856);
and U14491 (N_14491,N_11729,N_11063);
or U14492 (N_14492,N_12448,N_12183);
or U14493 (N_14493,N_11669,N_12147);
nor U14494 (N_14494,N_10453,N_10536);
nand U14495 (N_14495,N_10754,N_12461);
or U14496 (N_14496,N_10874,N_11842);
nand U14497 (N_14497,N_11947,N_10211);
nand U14498 (N_14498,N_12089,N_10515);
or U14499 (N_14499,N_10871,N_10442);
and U14500 (N_14500,N_11292,N_10879);
nand U14501 (N_14501,N_11115,N_11338);
nor U14502 (N_14502,N_11380,N_10157);
nor U14503 (N_14503,N_10280,N_12473);
and U14504 (N_14504,N_11001,N_11651);
and U14505 (N_14505,N_12434,N_12449);
nor U14506 (N_14506,N_11449,N_12198);
or U14507 (N_14507,N_11989,N_10616);
and U14508 (N_14508,N_12138,N_10350);
nor U14509 (N_14509,N_10033,N_11962);
nand U14510 (N_14510,N_10233,N_10309);
nand U14511 (N_14511,N_11898,N_11894);
nor U14512 (N_14512,N_11084,N_12263);
or U14513 (N_14513,N_10613,N_10760);
or U14514 (N_14514,N_10578,N_10983);
and U14515 (N_14515,N_11561,N_10844);
or U14516 (N_14516,N_11850,N_11408);
nor U14517 (N_14517,N_11401,N_11249);
and U14518 (N_14518,N_11716,N_11407);
xor U14519 (N_14519,N_10787,N_10259);
and U14520 (N_14520,N_10776,N_11784);
nor U14521 (N_14521,N_10847,N_10910);
xor U14522 (N_14522,N_11648,N_12296);
nor U14523 (N_14523,N_10698,N_10364);
nor U14524 (N_14524,N_12360,N_12489);
and U14525 (N_14525,N_10947,N_10577);
and U14526 (N_14526,N_12354,N_12292);
nand U14527 (N_14527,N_11569,N_10513);
xnor U14528 (N_14528,N_10930,N_12221);
or U14529 (N_14529,N_12087,N_10351);
xnor U14530 (N_14530,N_11342,N_10452);
nor U14531 (N_14531,N_11365,N_11769);
nand U14532 (N_14532,N_11906,N_10831);
or U14533 (N_14533,N_10932,N_10213);
and U14534 (N_14534,N_12488,N_11126);
or U14535 (N_14535,N_12168,N_12455);
nand U14536 (N_14536,N_11964,N_12242);
or U14537 (N_14537,N_11512,N_10923);
and U14538 (N_14538,N_10425,N_11171);
or U14539 (N_14539,N_12082,N_11317);
nor U14540 (N_14540,N_11445,N_11650);
or U14541 (N_14541,N_11089,N_10335);
nand U14542 (N_14542,N_10421,N_11288);
or U14543 (N_14543,N_12005,N_12103);
nor U14544 (N_14544,N_11643,N_11236);
nand U14545 (N_14545,N_10513,N_11492);
nor U14546 (N_14546,N_10969,N_10924);
and U14547 (N_14547,N_12239,N_10930);
xor U14548 (N_14548,N_11159,N_11967);
nand U14549 (N_14549,N_12458,N_12253);
nand U14550 (N_14550,N_11203,N_12002);
or U14551 (N_14551,N_10389,N_11642);
nor U14552 (N_14552,N_10550,N_10301);
nand U14553 (N_14553,N_12357,N_10836);
or U14554 (N_14554,N_11640,N_11212);
and U14555 (N_14555,N_10256,N_12144);
nor U14556 (N_14556,N_11745,N_10996);
or U14557 (N_14557,N_12119,N_11017);
nor U14558 (N_14558,N_11369,N_11086);
nor U14559 (N_14559,N_11198,N_10318);
nor U14560 (N_14560,N_10208,N_10352);
xor U14561 (N_14561,N_10801,N_12163);
nor U14562 (N_14562,N_11415,N_10468);
nor U14563 (N_14563,N_11201,N_10954);
and U14564 (N_14564,N_10816,N_10119);
nand U14565 (N_14565,N_11367,N_12137);
nand U14566 (N_14566,N_11826,N_11573);
nand U14567 (N_14567,N_11302,N_10210);
nor U14568 (N_14568,N_11821,N_12192);
and U14569 (N_14569,N_12320,N_11060);
or U14570 (N_14570,N_10453,N_11731);
nor U14571 (N_14571,N_12100,N_10538);
nor U14572 (N_14572,N_11913,N_10266);
and U14573 (N_14573,N_10537,N_10293);
or U14574 (N_14574,N_10836,N_10994);
nor U14575 (N_14575,N_11548,N_10971);
nor U14576 (N_14576,N_11657,N_11282);
and U14577 (N_14577,N_10102,N_11171);
or U14578 (N_14578,N_10334,N_11911);
nor U14579 (N_14579,N_12466,N_10533);
or U14580 (N_14580,N_10622,N_10996);
nor U14581 (N_14581,N_10146,N_10734);
nand U14582 (N_14582,N_10068,N_12366);
nand U14583 (N_14583,N_12304,N_12247);
nand U14584 (N_14584,N_11718,N_10943);
and U14585 (N_14585,N_12300,N_11069);
or U14586 (N_14586,N_12458,N_11118);
and U14587 (N_14587,N_11943,N_10257);
or U14588 (N_14588,N_12098,N_10479);
nor U14589 (N_14589,N_12316,N_11159);
or U14590 (N_14590,N_11389,N_10559);
and U14591 (N_14591,N_11589,N_10192);
nor U14592 (N_14592,N_10339,N_12087);
xor U14593 (N_14593,N_10669,N_10237);
xor U14594 (N_14594,N_10552,N_11880);
nor U14595 (N_14595,N_12276,N_11806);
xnor U14596 (N_14596,N_10798,N_11605);
or U14597 (N_14597,N_11402,N_10419);
or U14598 (N_14598,N_11715,N_10447);
nor U14599 (N_14599,N_12346,N_12264);
nand U14600 (N_14600,N_10631,N_10506);
nand U14601 (N_14601,N_11386,N_11078);
xor U14602 (N_14602,N_12279,N_10732);
nand U14603 (N_14603,N_12304,N_11367);
or U14604 (N_14604,N_11103,N_10182);
and U14605 (N_14605,N_10055,N_10187);
or U14606 (N_14606,N_11554,N_11782);
nor U14607 (N_14607,N_11614,N_10555);
or U14608 (N_14608,N_12364,N_11105);
or U14609 (N_14609,N_10594,N_10482);
nor U14610 (N_14610,N_10776,N_11365);
nand U14611 (N_14611,N_11889,N_11044);
nor U14612 (N_14612,N_10442,N_10853);
and U14613 (N_14613,N_10560,N_12126);
nor U14614 (N_14614,N_10366,N_12261);
xor U14615 (N_14615,N_11104,N_12228);
or U14616 (N_14616,N_12245,N_12212);
nor U14617 (N_14617,N_11667,N_11746);
nand U14618 (N_14618,N_10395,N_10437);
nand U14619 (N_14619,N_11072,N_11276);
nor U14620 (N_14620,N_10811,N_10729);
nand U14621 (N_14621,N_10743,N_10025);
or U14622 (N_14622,N_11036,N_10958);
and U14623 (N_14623,N_12499,N_12036);
and U14624 (N_14624,N_11260,N_10239);
nand U14625 (N_14625,N_10170,N_10095);
and U14626 (N_14626,N_11273,N_11787);
xnor U14627 (N_14627,N_12097,N_10278);
nor U14628 (N_14628,N_10818,N_10955);
and U14629 (N_14629,N_12333,N_10946);
or U14630 (N_14630,N_11486,N_11570);
nor U14631 (N_14631,N_12114,N_10142);
xor U14632 (N_14632,N_11141,N_12323);
or U14633 (N_14633,N_11616,N_10502);
xnor U14634 (N_14634,N_11804,N_12080);
nor U14635 (N_14635,N_11634,N_11391);
nand U14636 (N_14636,N_11902,N_11448);
or U14637 (N_14637,N_11006,N_11865);
and U14638 (N_14638,N_11787,N_11877);
or U14639 (N_14639,N_10912,N_11461);
nand U14640 (N_14640,N_10038,N_12216);
nand U14641 (N_14641,N_11549,N_12306);
xor U14642 (N_14642,N_12117,N_10094);
or U14643 (N_14643,N_11928,N_11748);
nand U14644 (N_14644,N_10195,N_11599);
nor U14645 (N_14645,N_11220,N_11307);
nor U14646 (N_14646,N_11827,N_11371);
or U14647 (N_14647,N_10637,N_11863);
nor U14648 (N_14648,N_11643,N_12237);
nand U14649 (N_14649,N_12453,N_10212);
or U14650 (N_14650,N_11928,N_10606);
or U14651 (N_14651,N_12092,N_11757);
or U14652 (N_14652,N_12116,N_11420);
and U14653 (N_14653,N_12481,N_11534);
nand U14654 (N_14654,N_11416,N_11984);
xor U14655 (N_14655,N_10855,N_10427);
nand U14656 (N_14656,N_12022,N_10530);
or U14657 (N_14657,N_10297,N_11285);
nor U14658 (N_14658,N_12068,N_12226);
nor U14659 (N_14659,N_10964,N_11377);
nor U14660 (N_14660,N_11865,N_12075);
nand U14661 (N_14661,N_11966,N_12248);
or U14662 (N_14662,N_10803,N_11778);
and U14663 (N_14663,N_11214,N_12106);
and U14664 (N_14664,N_10519,N_11099);
or U14665 (N_14665,N_10622,N_10461);
nor U14666 (N_14666,N_12386,N_11056);
nand U14667 (N_14667,N_11707,N_10723);
nor U14668 (N_14668,N_10152,N_12104);
nand U14669 (N_14669,N_11722,N_10515);
or U14670 (N_14670,N_11952,N_12355);
or U14671 (N_14671,N_10144,N_10626);
xnor U14672 (N_14672,N_10720,N_10189);
and U14673 (N_14673,N_11002,N_11801);
xor U14674 (N_14674,N_12373,N_10875);
and U14675 (N_14675,N_12267,N_10067);
xor U14676 (N_14676,N_10620,N_11877);
or U14677 (N_14677,N_12400,N_11302);
nor U14678 (N_14678,N_12050,N_10563);
and U14679 (N_14679,N_12047,N_10421);
nand U14680 (N_14680,N_11655,N_12105);
xnor U14681 (N_14681,N_10566,N_10558);
and U14682 (N_14682,N_11026,N_11076);
xnor U14683 (N_14683,N_11565,N_10474);
or U14684 (N_14684,N_11811,N_11531);
xnor U14685 (N_14685,N_10158,N_11963);
or U14686 (N_14686,N_11075,N_11970);
nand U14687 (N_14687,N_12129,N_10857);
xor U14688 (N_14688,N_10589,N_12144);
nand U14689 (N_14689,N_12216,N_11531);
or U14690 (N_14690,N_11609,N_10455);
and U14691 (N_14691,N_11759,N_10281);
and U14692 (N_14692,N_11618,N_11558);
xor U14693 (N_14693,N_10124,N_10164);
nand U14694 (N_14694,N_11244,N_11112);
nand U14695 (N_14695,N_10556,N_10346);
xor U14696 (N_14696,N_11060,N_10631);
and U14697 (N_14697,N_12093,N_12194);
or U14698 (N_14698,N_10029,N_10147);
and U14699 (N_14699,N_10238,N_11118);
or U14700 (N_14700,N_12474,N_10552);
nor U14701 (N_14701,N_10208,N_11098);
nor U14702 (N_14702,N_11239,N_11631);
nand U14703 (N_14703,N_10761,N_10149);
nand U14704 (N_14704,N_10769,N_11410);
or U14705 (N_14705,N_11274,N_10429);
nor U14706 (N_14706,N_10224,N_12272);
and U14707 (N_14707,N_10319,N_10156);
and U14708 (N_14708,N_12193,N_10242);
xnor U14709 (N_14709,N_11440,N_11140);
nand U14710 (N_14710,N_10037,N_10227);
xnor U14711 (N_14711,N_12472,N_11980);
and U14712 (N_14712,N_11733,N_11771);
and U14713 (N_14713,N_10476,N_10513);
or U14714 (N_14714,N_11973,N_10019);
and U14715 (N_14715,N_10023,N_10943);
nor U14716 (N_14716,N_11548,N_11073);
nand U14717 (N_14717,N_10685,N_11394);
nand U14718 (N_14718,N_11880,N_11528);
nor U14719 (N_14719,N_11435,N_10131);
and U14720 (N_14720,N_11448,N_10740);
nor U14721 (N_14721,N_10168,N_10106);
nor U14722 (N_14722,N_11035,N_10582);
nor U14723 (N_14723,N_11666,N_12446);
nor U14724 (N_14724,N_10722,N_10865);
nand U14725 (N_14725,N_10610,N_11883);
nand U14726 (N_14726,N_10631,N_10960);
xor U14727 (N_14727,N_10963,N_10279);
or U14728 (N_14728,N_10977,N_11393);
and U14729 (N_14729,N_10275,N_12071);
and U14730 (N_14730,N_10899,N_10510);
nor U14731 (N_14731,N_11383,N_10224);
or U14732 (N_14732,N_10874,N_10462);
and U14733 (N_14733,N_10017,N_10204);
or U14734 (N_14734,N_11000,N_10420);
nand U14735 (N_14735,N_11061,N_12432);
or U14736 (N_14736,N_11206,N_10228);
and U14737 (N_14737,N_12260,N_12041);
or U14738 (N_14738,N_12262,N_10259);
and U14739 (N_14739,N_11366,N_12477);
nand U14740 (N_14740,N_11984,N_12489);
or U14741 (N_14741,N_10235,N_11290);
nor U14742 (N_14742,N_11209,N_11235);
and U14743 (N_14743,N_10335,N_11150);
and U14744 (N_14744,N_11529,N_10942);
and U14745 (N_14745,N_12110,N_12038);
or U14746 (N_14746,N_10693,N_10238);
nor U14747 (N_14747,N_10301,N_10423);
nand U14748 (N_14748,N_10386,N_10496);
nor U14749 (N_14749,N_10010,N_10910);
or U14750 (N_14750,N_11874,N_10659);
or U14751 (N_14751,N_12359,N_11129);
nand U14752 (N_14752,N_10046,N_11884);
nand U14753 (N_14753,N_12348,N_10252);
or U14754 (N_14754,N_10897,N_11460);
nor U14755 (N_14755,N_12446,N_12427);
nor U14756 (N_14756,N_12437,N_12351);
nor U14757 (N_14757,N_12090,N_12402);
or U14758 (N_14758,N_11040,N_11597);
nand U14759 (N_14759,N_11155,N_12138);
nand U14760 (N_14760,N_10351,N_12310);
or U14761 (N_14761,N_11737,N_10883);
nand U14762 (N_14762,N_11694,N_10197);
xnor U14763 (N_14763,N_10260,N_12482);
nor U14764 (N_14764,N_12381,N_10699);
nand U14765 (N_14765,N_10671,N_12322);
nand U14766 (N_14766,N_11830,N_11044);
or U14767 (N_14767,N_11093,N_10239);
or U14768 (N_14768,N_11256,N_10214);
and U14769 (N_14769,N_12487,N_11351);
and U14770 (N_14770,N_11398,N_10022);
or U14771 (N_14771,N_12246,N_11184);
or U14772 (N_14772,N_12457,N_11644);
nor U14773 (N_14773,N_11985,N_11127);
nand U14774 (N_14774,N_11283,N_12389);
xor U14775 (N_14775,N_10197,N_10444);
nor U14776 (N_14776,N_10203,N_10127);
nor U14777 (N_14777,N_10966,N_10419);
and U14778 (N_14778,N_10460,N_11208);
nor U14779 (N_14779,N_10718,N_10103);
xnor U14780 (N_14780,N_11673,N_10810);
nand U14781 (N_14781,N_11747,N_10771);
nor U14782 (N_14782,N_10732,N_11171);
and U14783 (N_14783,N_11450,N_10758);
nor U14784 (N_14784,N_10272,N_12312);
nor U14785 (N_14785,N_11798,N_11163);
xnor U14786 (N_14786,N_10211,N_12265);
and U14787 (N_14787,N_11612,N_11731);
nor U14788 (N_14788,N_10514,N_10603);
nor U14789 (N_14789,N_10664,N_10439);
or U14790 (N_14790,N_12172,N_12029);
and U14791 (N_14791,N_10052,N_10291);
nand U14792 (N_14792,N_11267,N_12206);
nand U14793 (N_14793,N_10503,N_12191);
and U14794 (N_14794,N_11426,N_10830);
and U14795 (N_14795,N_11785,N_10133);
and U14796 (N_14796,N_10105,N_11227);
or U14797 (N_14797,N_10753,N_11616);
nor U14798 (N_14798,N_10728,N_12031);
nor U14799 (N_14799,N_11147,N_10037);
nand U14800 (N_14800,N_10646,N_12250);
nor U14801 (N_14801,N_11204,N_11037);
nor U14802 (N_14802,N_11882,N_11137);
or U14803 (N_14803,N_11993,N_11387);
or U14804 (N_14804,N_11404,N_10437);
or U14805 (N_14805,N_11883,N_10004);
nand U14806 (N_14806,N_10033,N_10718);
nand U14807 (N_14807,N_11707,N_12395);
and U14808 (N_14808,N_11037,N_10301);
nand U14809 (N_14809,N_11908,N_11046);
nor U14810 (N_14810,N_10742,N_10028);
nor U14811 (N_14811,N_10042,N_11958);
and U14812 (N_14812,N_10700,N_10256);
or U14813 (N_14813,N_11766,N_10219);
nor U14814 (N_14814,N_10279,N_12417);
or U14815 (N_14815,N_10969,N_11543);
nor U14816 (N_14816,N_10917,N_11608);
nor U14817 (N_14817,N_12427,N_10289);
nor U14818 (N_14818,N_10366,N_10102);
or U14819 (N_14819,N_12165,N_10133);
and U14820 (N_14820,N_10697,N_11959);
nand U14821 (N_14821,N_10183,N_11351);
and U14822 (N_14822,N_11155,N_11063);
and U14823 (N_14823,N_12197,N_10736);
or U14824 (N_14824,N_12493,N_10031);
and U14825 (N_14825,N_10619,N_10401);
nor U14826 (N_14826,N_12283,N_10443);
nor U14827 (N_14827,N_10015,N_11168);
nand U14828 (N_14828,N_10270,N_10589);
xnor U14829 (N_14829,N_11251,N_10948);
xnor U14830 (N_14830,N_10838,N_11248);
nand U14831 (N_14831,N_10755,N_11129);
nand U14832 (N_14832,N_10442,N_11646);
or U14833 (N_14833,N_11962,N_10006);
and U14834 (N_14834,N_11475,N_10835);
and U14835 (N_14835,N_11393,N_10744);
xnor U14836 (N_14836,N_10717,N_10273);
and U14837 (N_14837,N_10674,N_10095);
nand U14838 (N_14838,N_11330,N_11165);
or U14839 (N_14839,N_10024,N_10609);
nor U14840 (N_14840,N_12429,N_10843);
nand U14841 (N_14841,N_10527,N_11671);
nand U14842 (N_14842,N_11867,N_12154);
nor U14843 (N_14843,N_11301,N_11405);
xor U14844 (N_14844,N_11684,N_10552);
and U14845 (N_14845,N_12347,N_11686);
or U14846 (N_14846,N_10973,N_10385);
or U14847 (N_14847,N_10750,N_12187);
or U14848 (N_14848,N_10691,N_10914);
and U14849 (N_14849,N_11126,N_10604);
and U14850 (N_14850,N_10335,N_11158);
nor U14851 (N_14851,N_12430,N_10876);
and U14852 (N_14852,N_12137,N_10552);
nor U14853 (N_14853,N_10489,N_12368);
or U14854 (N_14854,N_11134,N_10342);
and U14855 (N_14855,N_11098,N_10572);
nand U14856 (N_14856,N_10800,N_10798);
nand U14857 (N_14857,N_11926,N_12011);
xor U14858 (N_14858,N_11232,N_12353);
or U14859 (N_14859,N_10484,N_12457);
nand U14860 (N_14860,N_12301,N_12117);
nor U14861 (N_14861,N_11934,N_10490);
or U14862 (N_14862,N_10227,N_12113);
nor U14863 (N_14863,N_12432,N_10409);
nor U14864 (N_14864,N_10787,N_10470);
or U14865 (N_14865,N_12035,N_10678);
or U14866 (N_14866,N_12482,N_11280);
nor U14867 (N_14867,N_12412,N_10398);
and U14868 (N_14868,N_11331,N_11336);
nor U14869 (N_14869,N_11039,N_11858);
nand U14870 (N_14870,N_11272,N_11955);
and U14871 (N_14871,N_10336,N_10498);
or U14872 (N_14872,N_10315,N_12159);
or U14873 (N_14873,N_10981,N_11055);
and U14874 (N_14874,N_10719,N_12279);
nand U14875 (N_14875,N_11947,N_10351);
or U14876 (N_14876,N_11441,N_11479);
nor U14877 (N_14877,N_12045,N_12429);
and U14878 (N_14878,N_10505,N_11623);
or U14879 (N_14879,N_10121,N_12077);
nand U14880 (N_14880,N_12323,N_11172);
or U14881 (N_14881,N_10526,N_11497);
nand U14882 (N_14882,N_10028,N_11046);
and U14883 (N_14883,N_12021,N_12456);
and U14884 (N_14884,N_11393,N_12133);
nand U14885 (N_14885,N_11267,N_11713);
and U14886 (N_14886,N_10145,N_10053);
nor U14887 (N_14887,N_12477,N_11598);
or U14888 (N_14888,N_12433,N_10478);
xnor U14889 (N_14889,N_11516,N_11648);
nand U14890 (N_14890,N_11329,N_11655);
or U14891 (N_14891,N_10664,N_12397);
nand U14892 (N_14892,N_10264,N_11546);
and U14893 (N_14893,N_11956,N_10749);
xnor U14894 (N_14894,N_11717,N_12354);
and U14895 (N_14895,N_10996,N_10962);
nand U14896 (N_14896,N_10710,N_11015);
or U14897 (N_14897,N_12237,N_11311);
or U14898 (N_14898,N_11485,N_10387);
nor U14899 (N_14899,N_11340,N_10514);
nor U14900 (N_14900,N_10093,N_10538);
nor U14901 (N_14901,N_12396,N_11791);
or U14902 (N_14902,N_10329,N_10546);
nor U14903 (N_14903,N_11429,N_10861);
nand U14904 (N_14904,N_11346,N_10756);
nor U14905 (N_14905,N_11985,N_12496);
nand U14906 (N_14906,N_10484,N_12244);
xor U14907 (N_14907,N_11319,N_10039);
or U14908 (N_14908,N_11302,N_12201);
and U14909 (N_14909,N_11099,N_10368);
and U14910 (N_14910,N_11575,N_11707);
xor U14911 (N_14911,N_10569,N_11327);
nor U14912 (N_14912,N_10088,N_12239);
nor U14913 (N_14913,N_11045,N_11606);
nor U14914 (N_14914,N_10435,N_10334);
or U14915 (N_14915,N_12261,N_11544);
and U14916 (N_14916,N_11978,N_11362);
nand U14917 (N_14917,N_11567,N_11371);
nor U14918 (N_14918,N_11713,N_11159);
nand U14919 (N_14919,N_10502,N_12439);
or U14920 (N_14920,N_10589,N_12358);
or U14921 (N_14921,N_10380,N_10015);
nand U14922 (N_14922,N_11220,N_12326);
or U14923 (N_14923,N_10931,N_11194);
nand U14924 (N_14924,N_10083,N_11137);
or U14925 (N_14925,N_11303,N_10224);
nor U14926 (N_14926,N_12240,N_10457);
and U14927 (N_14927,N_10030,N_10791);
and U14928 (N_14928,N_10841,N_12193);
nor U14929 (N_14929,N_12065,N_11943);
or U14930 (N_14930,N_12443,N_11141);
and U14931 (N_14931,N_10130,N_10655);
xnor U14932 (N_14932,N_10142,N_11704);
or U14933 (N_14933,N_12470,N_10120);
nor U14934 (N_14934,N_10832,N_11551);
nor U14935 (N_14935,N_12149,N_12159);
or U14936 (N_14936,N_10625,N_10495);
or U14937 (N_14937,N_11028,N_10540);
xor U14938 (N_14938,N_10452,N_11119);
nand U14939 (N_14939,N_11703,N_11343);
and U14940 (N_14940,N_11962,N_11058);
nand U14941 (N_14941,N_11800,N_10302);
and U14942 (N_14942,N_11181,N_11212);
nand U14943 (N_14943,N_10220,N_11199);
xor U14944 (N_14944,N_11292,N_10030);
and U14945 (N_14945,N_11204,N_10719);
nand U14946 (N_14946,N_11712,N_10371);
or U14947 (N_14947,N_11327,N_10324);
nand U14948 (N_14948,N_11179,N_11994);
xnor U14949 (N_14949,N_11489,N_11938);
nand U14950 (N_14950,N_11635,N_11203);
xnor U14951 (N_14951,N_11055,N_10820);
nor U14952 (N_14952,N_11550,N_10204);
nand U14953 (N_14953,N_11220,N_10980);
and U14954 (N_14954,N_10479,N_12386);
or U14955 (N_14955,N_10649,N_11445);
nor U14956 (N_14956,N_10475,N_10171);
nor U14957 (N_14957,N_11802,N_10606);
and U14958 (N_14958,N_11673,N_10235);
xor U14959 (N_14959,N_11728,N_11838);
nand U14960 (N_14960,N_10396,N_11679);
and U14961 (N_14961,N_11939,N_11712);
nand U14962 (N_14962,N_12482,N_10846);
nor U14963 (N_14963,N_12435,N_10346);
nor U14964 (N_14964,N_10679,N_12221);
nand U14965 (N_14965,N_10817,N_11090);
xnor U14966 (N_14966,N_11861,N_12244);
and U14967 (N_14967,N_11696,N_11909);
or U14968 (N_14968,N_11923,N_11640);
nand U14969 (N_14969,N_10737,N_11108);
xnor U14970 (N_14970,N_10329,N_10503);
or U14971 (N_14971,N_12238,N_10688);
nand U14972 (N_14972,N_10706,N_12351);
nand U14973 (N_14973,N_10184,N_11756);
or U14974 (N_14974,N_10574,N_12464);
nand U14975 (N_14975,N_11859,N_10372);
nor U14976 (N_14976,N_11923,N_11535);
or U14977 (N_14977,N_11799,N_11608);
or U14978 (N_14978,N_11729,N_11908);
or U14979 (N_14979,N_10795,N_10734);
xor U14980 (N_14980,N_10745,N_10427);
or U14981 (N_14981,N_11542,N_11528);
nor U14982 (N_14982,N_11152,N_12431);
or U14983 (N_14983,N_11802,N_12112);
nor U14984 (N_14984,N_11119,N_10028);
nand U14985 (N_14985,N_11084,N_10501);
or U14986 (N_14986,N_10477,N_10655);
nand U14987 (N_14987,N_10483,N_11183);
nand U14988 (N_14988,N_11821,N_11863);
and U14989 (N_14989,N_10703,N_11796);
and U14990 (N_14990,N_10334,N_11538);
and U14991 (N_14991,N_11575,N_10366);
or U14992 (N_14992,N_12281,N_11159);
nor U14993 (N_14993,N_11962,N_12102);
nor U14994 (N_14994,N_10569,N_12413);
nand U14995 (N_14995,N_11508,N_10891);
xnor U14996 (N_14996,N_10466,N_12267);
and U14997 (N_14997,N_11350,N_10771);
or U14998 (N_14998,N_10372,N_10483);
nand U14999 (N_14999,N_10225,N_11204);
nand U15000 (N_15000,N_12967,N_12709);
or U15001 (N_15001,N_13981,N_12540);
nor U15002 (N_15002,N_13148,N_13832);
and U15003 (N_15003,N_14674,N_13635);
nor U15004 (N_15004,N_13095,N_14154);
nor U15005 (N_15005,N_14123,N_13028);
or U15006 (N_15006,N_14333,N_13762);
nand U15007 (N_15007,N_13657,N_12924);
and U15008 (N_15008,N_12985,N_14953);
nor U15009 (N_15009,N_12989,N_13269);
or U15010 (N_15010,N_13172,N_13447);
nor U15011 (N_15011,N_14245,N_12689);
nor U15012 (N_15012,N_14105,N_13619);
nand U15013 (N_15013,N_14803,N_14931);
nor U15014 (N_15014,N_13106,N_12559);
or U15015 (N_15015,N_12671,N_13519);
nand U15016 (N_15016,N_13501,N_12839);
nand U15017 (N_15017,N_13822,N_14808);
nand U15018 (N_15018,N_14992,N_13354);
or U15019 (N_15019,N_13339,N_14051);
or U15020 (N_15020,N_14131,N_14463);
xor U15021 (N_15021,N_12759,N_13488);
or U15022 (N_15022,N_12968,N_14113);
or U15023 (N_15023,N_14689,N_13013);
nor U15024 (N_15024,N_13340,N_14912);
nor U15025 (N_15025,N_14576,N_14714);
nor U15026 (N_15026,N_12717,N_13472);
and U15027 (N_15027,N_12631,N_13192);
or U15028 (N_15028,N_14868,N_14987);
nor U15029 (N_15029,N_13764,N_14967);
xor U15030 (N_15030,N_14523,N_14046);
or U15031 (N_15031,N_14181,N_13716);
and U15032 (N_15032,N_14276,N_14966);
nand U15033 (N_15033,N_13734,N_14741);
nand U15034 (N_15034,N_12529,N_13471);
nor U15035 (N_15035,N_14422,N_14448);
nor U15036 (N_15036,N_14325,N_12750);
nor U15037 (N_15037,N_14455,N_14350);
nor U15038 (N_15038,N_13211,N_12683);
and U15039 (N_15039,N_13161,N_12783);
nand U15040 (N_15040,N_14215,N_14032);
nor U15041 (N_15041,N_14942,N_12686);
and U15042 (N_15042,N_14745,N_14853);
xor U15043 (N_15043,N_13539,N_14048);
nand U15044 (N_15044,N_13986,N_12518);
nor U15045 (N_15045,N_12713,N_14227);
or U15046 (N_15046,N_14795,N_13553);
and U15047 (N_15047,N_12746,N_14343);
nand U15048 (N_15048,N_13837,N_12542);
xnor U15049 (N_15049,N_12579,N_14749);
nand U15050 (N_15050,N_14704,N_13032);
and U15051 (N_15051,N_13755,N_13493);
nor U15052 (N_15052,N_14581,N_13191);
xor U15053 (N_15053,N_12807,N_14974);
and U15054 (N_15054,N_14817,N_13468);
xnor U15055 (N_15055,N_13546,N_13079);
xor U15056 (N_15056,N_13378,N_12606);
or U15057 (N_15057,N_14417,N_13248);
or U15058 (N_15058,N_14374,N_13630);
xor U15059 (N_15059,N_13512,N_14190);
nor U15060 (N_15060,N_13311,N_13479);
xnor U15061 (N_15061,N_14057,N_13955);
nor U15062 (N_15062,N_13111,N_13499);
and U15063 (N_15063,N_13157,N_14321);
and U15064 (N_15064,N_12587,N_12840);
xnor U15065 (N_15065,N_14027,N_13025);
nand U15066 (N_15066,N_13902,N_13906);
nor U15067 (N_15067,N_14490,N_14693);
or U15068 (N_15068,N_13633,N_13490);
nand U15069 (N_15069,N_13541,N_13850);
and U15070 (N_15070,N_12639,N_14452);
nand U15071 (N_15071,N_13708,N_13104);
xnor U15072 (N_15072,N_12948,N_13187);
or U15073 (N_15073,N_14952,N_14641);
and U15074 (N_15074,N_13632,N_12655);
nor U15075 (N_15075,N_14198,N_13403);
or U15076 (N_15076,N_12550,N_13272);
nor U15077 (N_15077,N_12771,N_13126);
or U15078 (N_15078,N_13420,N_12660);
nand U15079 (N_15079,N_14908,N_13418);
and U15080 (N_15080,N_14110,N_13421);
or U15081 (N_15081,N_13386,N_14259);
nand U15082 (N_15082,N_14766,N_14064);
nand U15083 (N_15083,N_14429,N_12982);
and U15084 (N_15084,N_12860,N_13010);
and U15085 (N_15085,N_12932,N_12563);
xor U15086 (N_15086,N_14059,N_13449);
and U15087 (N_15087,N_12941,N_12621);
nand U15088 (N_15088,N_13536,N_13326);
nand U15089 (N_15089,N_12749,N_14486);
or U15090 (N_15090,N_13655,N_12926);
xor U15091 (N_15091,N_14171,N_13586);
nor U15092 (N_15092,N_12635,N_14017);
and U15093 (N_15093,N_14661,N_14193);
nand U15094 (N_15094,N_13377,N_13394);
nand U15095 (N_15095,N_13252,N_12755);
nand U15096 (N_15096,N_12641,N_14118);
or U15097 (N_15097,N_14183,N_13243);
nand U15098 (N_15098,N_14068,N_14652);
or U15099 (N_15099,N_14530,N_14251);
xnor U15100 (N_15100,N_13469,N_13615);
nor U15101 (N_15101,N_12902,N_12761);
nand U15102 (N_15102,N_13116,N_13786);
or U15103 (N_15103,N_12500,N_12907);
nand U15104 (N_15104,N_14407,N_14135);
or U15105 (N_15105,N_13690,N_12585);
nand U15106 (N_15106,N_12520,N_14638);
or U15107 (N_15107,N_14443,N_14380);
or U15108 (N_15108,N_14869,N_13180);
nor U15109 (N_15109,N_12690,N_14377);
and U15110 (N_15110,N_12541,N_12573);
or U15111 (N_15111,N_13034,N_13925);
xor U15112 (N_15112,N_13941,N_12675);
nand U15113 (N_15113,N_13276,N_13895);
or U15114 (N_15114,N_12789,N_12917);
and U15115 (N_15115,N_13004,N_14695);
nand U15116 (N_15116,N_13531,N_13054);
nor U15117 (N_15117,N_12990,N_13369);
nor U15118 (N_15118,N_13450,N_13090);
nand U15119 (N_15119,N_14209,N_12528);
and U15120 (N_15120,N_13149,N_13933);
nor U15121 (N_15121,N_14628,N_13367);
nand U15122 (N_15122,N_13576,N_14594);
and U15123 (N_15123,N_14454,N_13617);
nor U15124 (N_15124,N_12741,N_14290);
nor U15125 (N_15125,N_13330,N_13346);
and U15126 (N_15126,N_13799,N_14717);
or U15127 (N_15127,N_13834,N_13560);
nor U15128 (N_15128,N_14986,N_13274);
nor U15129 (N_15129,N_14881,N_12855);
xor U15130 (N_15130,N_14849,N_13058);
or U15131 (N_15131,N_14143,N_12915);
or U15132 (N_15132,N_12583,N_12963);
nor U15133 (N_15133,N_14816,N_13807);
and U15134 (N_15134,N_14438,N_13757);
xor U15135 (N_15135,N_14832,N_14201);
nand U15136 (N_15136,N_13975,N_13598);
nand U15137 (N_15137,N_13721,N_12938);
or U15138 (N_15138,N_13171,N_13007);
and U15139 (N_15139,N_13724,N_14911);
or U15140 (N_15140,N_14132,N_13894);
or U15141 (N_15141,N_14929,N_14610);
or U15142 (N_15142,N_14780,N_14405);
or U15143 (N_15143,N_14657,N_13684);
and U15144 (N_15144,N_14859,N_13069);
nand U15145 (N_15145,N_14999,N_14239);
and U15146 (N_15146,N_14044,N_14677);
nand U15147 (N_15147,N_14169,N_13525);
and U15148 (N_15148,N_13517,N_12527);
nand U15149 (N_15149,N_12797,N_13736);
or U15150 (N_15150,N_13431,N_12548);
nor U15151 (N_15151,N_14735,N_14563);
nand U15152 (N_15152,N_13543,N_14034);
nor U15153 (N_15153,N_12972,N_13821);
nor U15154 (N_15154,N_12584,N_12833);
and U15155 (N_15155,N_14274,N_12906);
nor U15156 (N_15156,N_14412,N_13137);
xnor U15157 (N_15157,N_12707,N_13545);
nor U15158 (N_15158,N_13751,N_12533);
and U15159 (N_15159,N_12880,N_13990);
nor U15160 (N_15160,N_12590,N_13068);
or U15161 (N_15161,N_12796,N_13454);
and U15162 (N_15162,N_13489,N_14872);
nor U15163 (N_15163,N_12653,N_13145);
and U15164 (N_15164,N_12888,N_12558);
or U15165 (N_15165,N_14702,N_13198);
nand U15166 (N_15166,N_14371,N_13816);
nand U15167 (N_15167,N_13230,N_14852);
and U15168 (N_15168,N_12599,N_12719);
nand U15169 (N_15169,N_13527,N_13959);
nor U15170 (N_15170,N_12571,N_14208);
or U15171 (N_15171,N_13524,N_12992);
nand U15172 (N_15172,N_12658,N_12512);
nor U15173 (N_15173,N_14372,N_12838);
and U15174 (N_15174,N_13582,N_14993);
and U15175 (N_15175,N_13830,N_14386);
xor U15176 (N_15176,N_13446,N_13001);
nand U15177 (N_15177,N_13364,N_14360);
nand U15178 (N_15178,N_12504,N_14867);
nor U15179 (N_15179,N_13485,N_13915);
and U15180 (N_15180,N_12645,N_13491);
and U15181 (N_15181,N_14841,N_12617);
and U15182 (N_15182,N_13967,N_14344);
and U15183 (N_15183,N_14876,N_12923);
nor U15184 (N_15184,N_13650,N_13701);
nor U15185 (N_15185,N_14682,N_13119);
and U15186 (N_15186,N_12501,N_13996);
and U15187 (N_15187,N_14409,N_13196);
nor U15188 (N_15188,N_13885,N_13162);
nand U15189 (N_15189,N_13238,N_14379);
or U15190 (N_15190,N_13995,N_14444);
nand U15191 (N_15191,N_14678,N_14725);
or U15192 (N_15192,N_13671,N_12710);
and U15193 (N_15193,N_12775,N_14591);
nor U15194 (N_15194,N_14025,N_14280);
nor U15195 (N_15195,N_14896,N_14546);
or U15196 (N_15196,N_12800,N_13642);
or U15197 (N_15197,N_14261,N_12736);
nor U15198 (N_15198,N_14042,N_12505);
or U15199 (N_15199,N_14436,N_14771);
nand U15200 (N_15200,N_14363,N_14187);
nand U15201 (N_15201,N_14398,N_14618);
nor U15202 (N_15202,N_12572,N_13629);
and U15203 (N_15203,N_12899,N_13011);
nor U15204 (N_15204,N_13968,N_13964);
and U15205 (N_15205,N_13298,N_13924);
nor U15206 (N_15206,N_12859,N_14865);
or U15207 (N_15207,N_14621,N_13224);
and U15208 (N_15208,N_13960,N_13511);
or U15209 (N_15209,N_13686,N_14310);
nand U15210 (N_15210,N_14010,N_14100);
xnor U15211 (N_15211,N_14770,N_14514);
nand U15212 (N_15212,N_13206,N_14778);
nand U15213 (N_15213,N_13002,N_14570);
and U15214 (N_15214,N_14294,N_14312);
nand U15215 (N_15215,N_12918,N_12753);
nand U15216 (N_15216,N_12703,N_13522);
nor U15217 (N_15217,N_13153,N_13048);
nor U15218 (N_15218,N_12715,N_13273);
xor U15219 (N_15219,N_12580,N_12969);
nor U15220 (N_15220,N_12594,N_14843);
and U15221 (N_15221,N_13950,N_13646);
nand U15222 (N_15222,N_14728,N_14602);
nand U15223 (N_15223,N_12619,N_14699);
or U15224 (N_15224,N_14821,N_14271);
or U15225 (N_15225,N_13218,N_14041);
nand U15226 (N_15226,N_12945,N_12662);
and U15227 (N_15227,N_14352,N_13801);
nand U15228 (N_15228,N_12592,N_12965);
and U15229 (N_15229,N_13666,N_14128);
nand U15230 (N_15230,N_14499,N_14058);
nand U15231 (N_15231,N_13572,N_14680);
or U15232 (N_15232,N_14178,N_13453);
nor U15233 (N_15233,N_14098,N_12966);
and U15234 (N_15234,N_13208,N_13936);
nor U15235 (N_15235,N_14762,N_13678);
nor U15236 (N_15236,N_14604,N_13637);
nand U15237 (N_15237,N_14767,N_14583);
and U15238 (N_15238,N_12596,N_14093);
and U15239 (N_15239,N_14909,N_12947);
xnor U15240 (N_15240,N_13215,N_14777);
and U15241 (N_15241,N_14804,N_12851);
nor U15242 (N_15242,N_13306,N_14985);
or U15243 (N_15243,N_13983,N_14529);
or U15244 (N_15244,N_14081,N_14461);
nor U15245 (N_15245,N_12776,N_13518);
or U15246 (N_15246,N_14316,N_14283);
xnor U15247 (N_15247,N_13791,N_14229);
or U15248 (N_15248,N_14266,N_12987);
and U15249 (N_15249,N_13513,N_13426);
or U15250 (N_15250,N_14785,N_14216);
xor U15251 (N_15251,N_14149,N_13739);
or U15252 (N_15252,N_13315,N_14014);
and U15253 (N_15253,N_13288,N_14424);
or U15254 (N_15254,N_14792,N_13839);
nor U15255 (N_15255,N_14401,N_13336);
nand U15256 (N_15256,N_13201,N_13703);
nand U15257 (N_15257,N_14439,N_14561);
nand U15258 (N_15258,N_13737,N_12806);
nand U15259 (N_15259,N_13840,N_12552);
and U15260 (N_15260,N_12757,N_13029);
or U15261 (N_15261,N_12943,N_14532);
xnor U15262 (N_15262,N_13889,N_12661);
nor U15263 (N_15263,N_14200,N_14440);
nor U15264 (N_15264,N_13664,N_12513);
nand U15265 (N_15265,N_13929,N_12685);
nand U15266 (N_15266,N_13796,N_14511);
and U15267 (N_15267,N_14844,N_13831);
nand U15268 (N_15268,N_12980,N_12524);
nand U15269 (N_15269,N_12567,N_13689);
xor U15270 (N_15270,N_14148,N_13170);
or U15271 (N_15271,N_13815,N_14115);
and U15272 (N_15272,N_12701,N_14164);
or U15273 (N_15273,N_14559,N_12700);
and U15274 (N_15274,N_14427,N_14395);
xnor U15275 (N_15275,N_13535,N_14207);
nand U15276 (N_15276,N_14501,N_13754);
nand U15277 (N_15277,N_13085,N_12756);
and U15278 (N_15278,N_12691,N_12673);
nor U15279 (N_15279,N_14815,N_13140);
nand U15280 (N_15280,N_14731,N_12808);
nor U15281 (N_15281,N_12962,N_12852);
xnor U15282 (N_15282,N_12821,N_14159);
or U15283 (N_15283,N_13563,N_14775);
and U15284 (N_15284,N_14472,N_14716);
and U15285 (N_15285,N_13712,N_14217);
nand U15286 (N_15286,N_13970,N_12971);
nor U15287 (N_15287,N_14161,N_12976);
nand U15288 (N_15288,N_12679,N_13455);
and U15289 (N_15289,N_14644,N_13595);
or U15290 (N_15290,N_12726,N_14267);
nand U15291 (N_15291,N_13898,N_14568);
and U15292 (N_15292,N_13030,N_12799);
or U15293 (N_15293,N_12603,N_14060);
nand U15294 (N_15294,N_12654,N_13350);
nand U15295 (N_15295,N_12648,N_14936);
nor U15296 (N_15296,N_13564,N_12886);
or U15297 (N_15297,N_14323,N_14700);
or U15298 (N_15298,N_14203,N_14988);
and U15299 (N_15299,N_13949,N_14155);
nand U15300 (N_15300,N_13761,N_14813);
nor U15301 (N_15301,N_12916,N_14650);
or U15302 (N_15302,N_14550,N_13718);
nand U15303 (N_15303,N_13413,N_14074);
and U15304 (N_15304,N_12725,N_14662);
nor U15305 (N_15305,N_13858,N_14957);
xor U15306 (N_15306,N_14219,N_14194);
and U15307 (N_15307,N_13132,N_14537);
nor U15308 (N_15308,N_12729,N_13334);
nor U15309 (N_15309,N_12826,N_13317);
nor U15310 (N_15310,N_14491,N_13884);
or U15311 (N_15311,N_14531,N_12752);
or U15312 (N_15312,N_13798,N_14166);
and U15313 (N_15313,N_13168,N_13649);
nor U15314 (N_15314,N_13193,N_14527);
nor U15315 (N_15315,N_13320,N_13961);
nor U15316 (N_15316,N_13258,N_13121);
xor U15317 (N_15317,N_14697,N_14920);
nor U15318 (N_15318,N_14337,N_12844);
nand U15319 (N_15319,N_13870,N_13297);
or U15320 (N_15320,N_14619,N_13973);
or U15321 (N_15321,N_13720,N_12870);
xor U15322 (N_15322,N_13901,N_13596);
xor U15323 (N_15323,N_12837,N_13345);
and U15324 (N_15324,N_14431,N_13711);
or U15325 (N_15325,N_12530,N_13337);
and U15326 (N_15326,N_13352,N_13189);
xor U15327 (N_15327,N_14989,N_14705);
and U15328 (N_15328,N_12861,N_14718);
and U15329 (N_15329,N_13185,N_14710);
or U15330 (N_15330,N_13747,N_13966);
nor U15331 (N_15331,N_13370,N_14249);
nor U15332 (N_15332,N_12910,N_13963);
xnor U15333 (N_15333,N_14631,N_13730);
and U15334 (N_15334,N_12908,N_13999);
or U15335 (N_15335,N_13125,N_13144);
nor U15336 (N_15336,N_13097,N_12677);
xnor U15337 (N_15337,N_13480,N_14268);
nand U15338 (N_15338,N_12921,N_13780);
and U15339 (N_15339,N_14740,N_13289);
nor U15340 (N_15340,N_12885,N_13406);
xnor U15341 (N_15341,N_14306,N_14946);
nor U15342 (N_15342,N_13587,N_14636);
or U15343 (N_15343,N_13552,N_13989);
or U15344 (N_15344,N_13382,N_13433);
xor U15345 (N_15345,N_14456,N_12986);
nor U15346 (N_15346,N_13246,N_14943);
xor U15347 (N_15347,N_14420,N_13448);
nor U15348 (N_15348,N_13284,N_14457);
nand U15349 (N_15349,N_14663,N_12818);
and U15350 (N_15350,N_13062,N_13991);
or U15351 (N_15351,N_14473,N_14856);
or U15352 (N_15352,N_14752,N_13935);
or U15353 (N_15353,N_13205,N_13329);
and U15354 (N_15354,N_14493,N_14759);
nor U15355 (N_15355,N_14298,N_12944);
nand U15356 (N_15356,N_13749,N_13390);
xnor U15357 (N_15357,N_13893,N_13738);
or U15358 (N_15358,N_14122,N_13475);
nand U15359 (N_15359,N_14314,N_13235);
nand U15360 (N_15360,N_13903,N_14389);
nand U15361 (N_15361,N_12984,N_13237);
xnor U15362 (N_15362,N_13809,N_14842);
nor U15363 (N_15363,N_13139,N_13881);
nand U15364 (N_15364,N_12723,N_14688);
xor U15365 (N_15365,N_14968,N_13729);
nand U15366 (N_15366,N_13200,N_12640);
nand U15367 (N_15367,N_14787,N_13926);
nor U15368 (N_15368,N_14554,N_12638);
nand U15369 (N_15369,N_13270,N_13653);
xnor U15370 (N_15370,N_14675,N_14180);
xor U15371 (N_15371,N_13003,N_14270);
and U15372 (N_15372,N_14134,N_13212);
and U15373 (N_15373,N_13251,N_13688);
nor U15374 (N_15374,N_14022,N_13395);
nand U15375 (N_15375,N_14263,N_13639);
nand U15376 (N_15376,N_13302,N_14676);
nand U15377 (N_15377,N_13725,N_14139);
or U15378 (N_15378,N_13958,N_14860);
nor U15379 (N_15379,N_14418,N_14525);
and U15380 (N_15380,N_14684,N_14300);
nor U15381 (N_15381,N_13027,N_12845);
xnor U15382 (N_15382,N_14996,N_12743);
or U15383 (N_15383,N_14781,N_13052);
or U15384 (N_15384,N_14757,N_12722);
or U15385 (N_15385,N_13474,N_13759);
nand U15386 (N_15386,N_12942,N_14696);
nor U15387 (N_15387,N_13808,N_14713);
and U15388 (N_15388,N_14130,N_13457);
nor U15389 (N_15389,N_14519,N_12934);
or U15390 (N_15390,N_14789,N_14221);
xor U15391 (N_15391,N_13865,N_13462);
and U15392 (N_15392,N_13673,N_12734);
and U15393 (N_15393,N_14308,N_13951);
nor U15394 (N_15394,N_14145,N_13940);
nand U15395 (N_15395,N_14620,N_14228);
nor U15396 (N_15396,N_14031,N_14573);
and U15397 (N_15397,N_13089,N_14367);
nand U15398 (N_15398,N_13624,N_12663);
nor U15399 (N_15399,N_14562,N_14277);
and U15400 (N_15400,N_12622,N_13366);
xnor U15401 (N_15401,N_13669,N_13213);
xor U15402 (N_15402,N_12656,N_14390);
nor U15403 (N_15403,N_13435,N_14857);
nand U15404 (N_15404,N_14050,N_13687);
and U15405 (N_15405,N_13473,N_14253);
nor U15406 (N_15406,N_14886,N_12554);
nand U15407 (N_15407,N_14230,N_13477);
nor U15408 (N_15408,N_13784,N_14827);
or U15409 (N_15409,N_13900,N_14430);
and U15410 (N_15410,N_13110,N_13355);
nand U15411 (N_15411,N_13652,N_12531);
or U15412 (N_15412,N_12697,N_13920);
and U15413 (N_15413,N_13937,N_13323);
or U15414 (N_15414,N_12576,N_13872);
xor U15415 (N_15415,N_13239,N_14520);
or U15416 (N_15416,N_14858,N_14796);
xnor U15417 (N_15417,N_12875,N_14466);
and U15418 (N_15418,N_14078,N_13574);
and U15419 (N_15419,N_12718,N_13072);
xor U15420 (N_15420,N_12801,N_13266);
nor U15421 (N_15421,N_14667,N_12695);
nor U15422 (N_15422,N_13074,N_14304);
nor U15423 (N_15423,N_13672,N_13609);
nand U15424 (N_15424,N_13108,N_14913);
nand U15425 (N_15425,N_13897,N_13380);
nor U15426 (N_15426,N_12716,N_14241);
nor U15427 (N_15427,N_14038,N_14692);
and U15428 (N_15428,N_12857,N_13668);
and U15429 (N_15429,N_13826,N_13226);
or U15430 (N_15430,N_14421,N_12925);
nand U15431 (N_15431,N_13282,N_13067);
nor U15432 (N_15432,N_12620,N_13216);
xor U15433 (N_15433,N_13982,N_14391);
and U15434 (N_15434,N_14930,N_14236);
nor U15435 (N_15435,N_13084,N_14978);
or U15436 (N_15436,N_13422,N_13165);
nor U15437 (N_15437,N_14332,N_13877);
or U15438 (N_15438,N_12618,N_13250);
nor U15439 (N_15439,N_13023,N_13614);
nand U15440 (N_15440,N_13777,N_14601);
nor U15441 (N_15441,N_14744,N_13828);
or U15442 (N_15442,N_14726,N_14838);
nand U15443 (N_15443,N_12706,N_14806);
or U15444 (N_15444,N_13594,N_13663);
and U15445 (N_15445,N_14192,N_14877);
nor U15446 (N_15446,N_14874,N_14863);
or U15447 (N_15447,N_12682,N_14924);
nor U15448 (N_15448,N_13411,N_14036);
nor U15449 (N_15449,N_14335,N_14346);
nand U15450 (N_15450,N_12961,N_12739);
and U15451 (N_15451,N_13083,N_14005);
nand U15452 (N_15452,N_12795,N_14470);
nand U15453 (N_15453,N_14719,N_13997);
xnor U15454 (N_15454,N_14585,N_13379);
nor U15455 (N_15455,N_12785,N_13965);
nand U15456 (N_15456,N_12568,N_14625);
xor U15457 (N_15457,N_14224,N_13580);
and U15458 (N_15458,N_14776,N_13221);
nor U15459 (N_15459,N_13878,N_13158);
or U15460 (N_15460,N_13167,N_13107);
nor U15461 (N_15461,N_13363,N_13064);
nand U15462 (N_15462,N_13114,N_12794);
nand U15463 (N_15463,N_13939,N_13980);
nor U15464 (N_15464,N_14013,N_12869);
nor U15465 (N_15465,N_14588,N_13727);
and U15466 (N_15466,N_14980,N_13497);
xnor U15467 (N_15467,N_12588,N_13636);
nand U15468 (N_15468,N_14605,N_12871);
xor U15469 (N_15469,N_12774,N_14954);
or U15470 (N_15470,N_14818,N_13886);
nand U15471 (N_15471,N_13694,N_14516);
and U15472 (N_15472,N_13508,N_12704);
nor U15473 (N_15473,N_14536,N_14094);
nand U15474 (N_15474,N_14907,N_13682);
or U15475 (N_15475,N_14165,N_14845);
nor U15476 (N_15476,N_14934,N_12991);
xor U15477 (N_15477,N_13548,N_14369);
and U15478 (N_15478,N_13043,N_12853);
xnor U15479 (N_15479,N_14299,N_13923);
xnor U15480 (N_15480,N_14708,N_13410);
nand U15481 (N_15481,N_14173,N_13102);
nand U15482 (N_15482,N_14982,N_12681);
or U15483 (N_15483,N_14542,N_13271);
and U15484 (N_15484,N_12762,N_13500);
or U15485 (N_15485,N_13645,N_14285);
and U15486 (N_15486,N_14730,N_14077);
or U15487 (N_15487,N_14750,N_13476);
nor U15488 (N_15488,N_14703,N_13229);
and U15489 (N_15489,N_12633,N_14979);
and U15490 (N_15490,N_13843,N_13098);
nand U15491 (N_15491,N_13581,N_14729);
nor U15492 (N_15492,N_14096,N_13583);
and U15493 (N_15493,N_13484,N_13735);
nand U15494 (N_15494,N_14072,N_14235);
and U15495 (N_15495,N_14141,N_13746);
nor U15496 (N_15496,N_13763,N_14348);
nand U15497 (N_15497,N_13376,N_14834);
and U15498 (N_15498,N_14969,N_13348);
or U15499 (N_15499,N_13338,N_12672);
or U15500 (N_15500,N_14887,N_13498);
or U15501 (N_15501,N_13082,N_14076);
or U15502 (N_15502,N_12767,N_14671);
nor U15503 (N_15503,N_14960,N_13452);
and U15504 (N_15504,N_13245,N_14011);
nor U15505 (N_15505,N_12896,N_14382);
xor U15506 (N_15506,N_12960,N_14172);
nand U15507 (N_15507,N_12608,N_12744);
and U15508 (N_15508,N_14737,N_14672);
nor U15509 (N_15509,N_14024,N_13827);
or U15510 (N_15510,N_13998,N_14721);
xnor U15511 (N_15511,N_13841,N_13254);
nor U15512 (N_15512,N_14883,N_14928);
xnor U15513 (N_15513,N_13740,N_14106);
nand U15514 (N_15514,N_14875,N_13823);
or U15515 (N_15515,N_14480,N_14471);
and U15516 (N_15516,N_14513,N_12667);
xor U15517 (N_15517,N_12507,N_14275);
and U15518 (N_15518,N_13241,N_12868);
nand U15519 (N_15519,N_14528,N_14426);
and U15520 (N_15520,N_14445,N_14289);
and U15521 (N_15521,N_13874,N_14204);
and U15522 (N_15522,N_14071,N_14903);
or U15523 (N_15523,N_13859,N_13533);
or U15524 (N_15524,N_14317,N_14615);
or U15525 (N_15525,N_14645,N_13232);
nor U15526 (N_15526,N_12534,N_12825);
xor U15527 (N_15527,N_12610,N_13295);
or U15528 (N_15528,N_13781,N_13863);
nand U15529 (N_15529,N_13717,N_12792);
or U15530 (N_15530,N_14467,N_14174);
nand U15531 (N_15531,N_13019,N_13327);
nor U15532 (N_15532,N_14892,N_13341);
or U15533 (N_15533,N_14938,N_13423);
or U15534 (N_15534,N_14400,N_13434);
nand U15535 (N_15535,N_13464,N_14428);
nand U15536 (N_15536,N_13209,N_14948);
and U15537 (N_15537,N_13060,N_12630);
nand U15538 (N_15538,N_14670,N_14889);
nor U15539 (N_15539,N_14167,N_13875);
or U15540 (N_15540,N_14080,N_13482);
or U15541 (N_15541,N_14894,N_14634);
nor U15542 (N_15542,N_14237,N_13318);
nand U15543 (N_15543,N_14595,N_13660);
xnor U15544 (N_15544,N_12809,N_14555);
and U15545 (N_15545,N_12854,N_13974);
and U15546 (N_15546,N_13549,N_14213);
or U15547 (N_15547,N_14811,N_12836);
and U15548 (N_15548,N_13620,N_14756);
and U15549 (N_15549,N_14373,N_13589);
nand U15550 (N_15550,N_13597,N_14265);
or U15551 (N_15551,N_14142,N_13388);
nand U15552 (N_15552,N_13538,N_13039);
nand U15553 (N_15553,N_13432,N_14399);
nor U15554 (N_15554,N_14496,N_13120);
and U15555 (N_15555,N_12889,N_14878);
xor U15556 (N_15556,N_14927,N_13222);
and U15557 (N_15557,N_13918,N_14376);
nand U15558 (N_15558,N_14260,N_13478);
nor U15559 (N_15559,N_13743,N_14281);
or U15560 (N_15560,N_13506,N_13676);
or U15561 (N_15561,N_14751,N_12856);
nand U15562 (N_15562,N_14854,N_13299);
and U15563 (N_15563,N_13806,N_13709);
nor U15564 (N_15564,N_14691,N_13921);
nor U15565 (N_15565,N_14545,N_13756);
xnor U15566 (N_15566,N_14250,N_14584);
nand U15567 (N_15567,N_14066,N_12903);
or U15568 (N_15568,N_12543,N_13662);
and U15569 (N_15569,N_14385,N_13020);
and U15570 (N_15570,N_13515,N_14956);
nand U15571 (N_15571,N_12830,N_12842);
nor U15572 (N_15572,N_13627,N_12577);
nor U15573 (N_15573,N_14774,N_13199);
or U15574 (N_15574,N_13123,N_14334);
or U15575 (N_15575,N_13804,N_12549);
xor U15576 (N_15576,N_14724,N_14160);
nor U15577 (N_15577,N_14917,N_13705);
and U15578 (N_15578,N_13142,N_12626);
nand U15579 (N_15579,N_12502,N_12632);
nand U15580 (N_15580,N_13324,N_13136);
nor U15581 (N_15581,N_12914,N_12705);
nand U15582 (N_15582,N_14088,N_13319);
nand U15583 (N_15583,N_13316,N_14309);
nor U15584 (N_15584,N_14891,N_13634);
and U15585 (N_15585,N_13914,N_14611);
and U15586 (N_15586,N_14353,N_13036);
nand U15587 (N_15587,N_14837,N_13887);
or U15588 (N_15588,N_13049,N_14836);
or U15589 (N_15589,N_14626,N_12953);
nor U15590 (N_15590,N_12887,N_12522);
nand U15591 (N_15591,N_14823,N_12930);
nand U15592 (N_15592,N_13631,N_13159);
and U15593 (N_15593,N_14474,N_13385);
and U15594 (N_15594,N_14915,N_14880);
nor U15595 (N_15595,N_13231,N_12575);
nor U15596 (N_15596,N_13602,N_14286);
and U15597 (N_15597,N_13190,N_14587);
nor U15598 (N_15598,N_14524,N_14177);
nor U15599 (N_15599,N_14895,N_14152);
and U15600 (N_15600,N_14240,N_12952);
xor U15601 (N_15601,N_12538,N_14720);
or U15602 (N_15602,N_13812,N_13803);
nand U15603 (N_15603,N_12738,N_14359);
nor U15604 (N_15604,N_13401,N_13891);
and U15605 (N_15605,N_13405,N_13467);
nand U15606 (N_15606,N_13101,N_13381);
or U15607 (N_15607,N_14754,N_12866);
nand U15608 (N_15608,N_13606,N_13992);
or U15609 (N_15609,N_13012,N_13117);
nor U15610 (N_15610,N_12816,N_13957);
or U15611 (N_15611,N_12773,N_14962);
nand U15612 (N_15612,N_14303,N_14690);
or U15613 (N_15613,N_14822,N_14184);
and U15614 (N_15614,N_13436,N_13134);
xor U15615 (N_15615,N_14861,N_14330);
nor U15616 (N_15616,N_14478,N_13706);
and U15617 (N_15617,N_12511,N_14451);
nand U15618 (N_15618,N_14922,N_13700);
and U15619 (N_15619,N_14313,N_14487);
and U15620 (N_15620,N_13625,N_13197);
and U15621 (N_15621,N_14539,N_12834);
xnor U15622 (N_15622,N_12546,N_12509);
or U15623 (N_15623,N_14949,N_12803);
nor U15624 (N_15624,N_12748,N_13943);
or U15625 (N_15625,N_14170,N_14392);
and U15626 (N_15626,N_12946,N_13817);
nor U15627 (N_15627,N_14415,N_14340);
nand U15628 (N_15628,N_14238,N_13045);
nor U15629 (N_15629,N_12936,N_12780);
or U15630 (N_15630,N_13994,N_13188);
and U15631 (N_15631,N_13829,N_12847);
and U15632 (N_15632,N_14509,N_13439);
xnor U15633 (N_15633,N_13483,N_13260);
nor U15634 (N_15634,N_14341,N_13772);
nor U15635 (N_15635,N_13138,N_13281);
or U15636 (N_15636,N_13607,N_13307);
nor U15637 (N_15637,N_14706,N_13322);
or U15638 (N_15638,N_12999,N_13932);
nand U15639 (N_15639,N_13156,N_13835);
or U15640 (N_15640,N_14168,N_13063);
nand U15641 (N_15641,N_12778,N_14965);
or U15642 (N_15642,N_14345,N_13509);
and U15643 (N_15643,N_14109,N_14772);
nand U15644 (N_15644,N_12883,N_13623);
xnor U15645 (N_15645,N_12850,N_13766);
nor U15646 (N_15646,N_13692,N_14681);
or U15647 (N_15647,N_13456,N_14319);
nand U15648 (N_15648,N_13309,N_14768);
nor U15649 (N_15649,N_13510,N_13584);
and U15650 (N_15650,N_14035,N_14764);
nand U15651 (N_15651,N_14632,N_13392);
and U15652 (N_15652,N_13600,N_14599);
or U15653 (N_15653,N_13301,N_12913);
nand U15654 (N_15654,N_12565,N_13728);
or U15655 (N_15655,N_14598,N_13523);
nand U15656 (N_15656,N_13031,N_13819);
and U15657 (N_15657,N_13601,N_13776);
and U15658 (N_15658,N_13516,N_12714);
nor U15659 (N_15659,N_14328,N_13585);
or U15660 (N_15660,N_14484,N_14107);
nor U15661 (N_15661,N_12574,N_14596);
xor U15662 (N_15662,N_12607,N_13041);
xor U15663 (N_15663,N_13788,N_14001);
nor U15664 (N_15664,N_14906,N_13278);
and U15665 (N_15665,N_12754,N_13035);
nand U15666 (N_15666,N_14893,N_14571);
nand U15667 (N_15667,N_12813,N_13109);
or U15668 (N_15668,N_12802,N_12788);
nand U15669 (N_15669,N_14256,N_12612);
nand U15670 (N_15670,N_13407,N_12911);
nand U15671 (N_15671,N_14809,N_12772);
and U15672 (N_15672,N_13308,N_13987);
or U15673 (N_15673,N_13103,N_13792);
or U15674 (N_15674,N_14202,N_14623);
nor U15675 (N_15675,N_13782,N_12634);
or U15676 (N_15676,N_13704,N_14257);
xor U15677 (N_15677,N_14507,N_13554);
xnor U15678 (N_15678,N_14541,N_12779);
or U15679 (N_15679,N_12874,N_12589);
or U15680 (N_15680,N_14084,N_12996);
or U15681 (N_15681,N_14665,N_12532);
xnor U15682 (N_15682,N_13820,N_14709);
nand U15683 (N_15683,N_14701,N_13285);
and U15684 (N_15684,N_12508,N_14904);
xor U15685 (N_15685,N_14322,N_13504);
and U15686 (N_15686,N_12553,N_12740);
nand U15687 (N_15687,N_13919,N_14820);
nand U15688 (N_15688,N_12994,N_14069);
xnor U15689 (N_15689,N_12760,N_14799);
and U15690 (N_15690,N_13015,N_13146);
and U15691 (N_15691,N_14939,N_14383);
nor U15692 (N_15692,N_14637,N_14921);
nand U15693 (N_15693,N_13922,N_14534);
or U15694 (N_15694,N_13534,N_14950);
or U15695 (N_15695,N_14797,N_13021);
nand U15696 (N_15696,N_14885,N_13628);
nor U15697 (N_15697,N_13356,N_12666);
nand U15698 (N_15698,N_14305,N_14103);
nor U15699 (N_15699,N_13143,N_13047);
and U15700 (N_15700,N_14790,N_13293);
and U15701 (N_15701,N_12694,N_13862);
xnor U15702 (N_15702,N_13971,N_14941);
and U15703 (N_15703,N_12712,N_14944);
and U15704 (N_15704,N_14423,N_13945);
nor U15705 (N_15705,N_14961,N_14589);
xnor U15706 (N_15706,N_13359,N_12882);
or U15707 (N_15707,N_13825,N_14847);
nor U15708 (N_15708,N_14075,N_14282);
or U15709 (N_15709,N_13693,N_13075);
and U15710 (N_15710,N_12831,N_14453);
nand U15711 (N_15711,N_14358,N_14413);
and U15712 (N_15712,N_13953,N_13934);
nor U15713 (N_15713,N_14375,N_13313);
or U15714 (N_15714,N_14108,N_12609);
or U15715 (N_15715,N_13240,N_14447);
nor U15716 (N_15716,N_14018,N_14825);
and U15717 (N_15717,N_14711,N_14600);
or U15718 (N_15718,N_14416,N_14381);
nand U15719 (N_15719,N_12770,N_13166);
nand U15720 (N_15720,N_14083,N_12858);
or U15721 (N_15721,N_14234,N_13417);
nor U15722 (N_15722,N_13268,N_14579);
xor U15723 (N_15723,N_13445,N_13438);
nor U15724 (N_15724,N_13351,N_12676);
or U15725 (N_15725,N_14362,N_14826);
and U15726 (N_15726,N_13679,N_13860);
nor U15727 (N_15727,N_13537,N_14252);
and U15728 (N_15728,N_14608,N_14535);
nor U15729 (N_15729,N_13066,N_14043);
and U15730 (N_15730,N_13430,N_12822);
or U15731 (N_15731,N_13869,N_13969);
and U15732 (N_15732,N_13264,N_14477);
nand U15733 (N_15733,N_13093,N_14864);
or U15734 (N_15734,N_14793,N_14408);
or U15735 (N_15735,N_13026,N_13133);
xor U15736 (N_15736,N_14425,N_14030);
nand U15737 (N_15737,N_14970,N_13593);
or U15738 (N_15738,N_12824,N_14357);
nand U15739 (N_15739,N_12892,N_13864);
and U15740 (N_15740,N_12790,N_13612);
nand U15741 (N_15741,N_12636,N_13459);
nor U15742 (N_15742,N_13466,N_12669);
nand U15743 (N_15743,N_14176,N_14147);
nand U15744 (N_15744,N_14747,N_14481);
and U15745 (N_15745,N_12922,N_14791);
nand U15746 (N_15746,N_14521,N_12555);
and U15747 (N_15747,N_14722,N_13750);
xnor U15748 (N_15748,N_14761,N_14121);
xor U15749 (N_15749,N_13851,N_12909);
and U15750 (N_15750,N_14156,N_13389);
and U15751 (N_15751,N_14897,N_14016);
nand U15752 (N_15752,N_14150,N_14153);
nand U15753 (N_15753,N_12781,N_14318);
or U15754 (N_15754,N_14432,N_13427);
and U15755 (N_15755,N_12595,N_14522);
and U15756 (N_15756,N_13626,N_12733);
and U15757 (N_15757,N_12651,N_13115);
nor U15758 (N_15758,N_13722,N_13547);
and U15759 (N_15759,N_13540,N_14510);
xnor U15760 (N_15760,N_12937,N_13696);
nand U15761 (N_15761,N_14666,N_14779);
nand U15762 (N_15762,N_14862,N_14067);
nor U15763 (N_15763,N_13038,N_14070);
xor U15764 (N_15764,N_12848,N_14404);
nand U15765 (N_15765,N_13494,N_14937);
xnor U15766 (N_15766,N_14021,N_14218);
nor U15767 (N_15767,N_14575,N_13393);
xor U15768 (N_15768,N_13460,N_14963);
or U15769 (N_15769,N_14464,N_12623);
nor U15770 (N_15770,N_13908,N_13988);
or U15771 (N_15771,N_14087,N_13733);
and U15772 (N_15772,N_14648,N_14533);
or U15773 (N_15773,N_13770,N_14654);
and U15774 (N_15774,N_14095,N_14125);
and U15775 (N_15775,N_13578,N_13715);
nor U15776 (N_15776,N_13181,N_13972);
xor U15777 (N_15777,N_13360,N_12805);
nor U15778 (N_15778,N_12535,N_14882);
nand U15779 (N_15779,N_14609,N_14073);
nand U15780 (N_15780,N_13178,N_12556);
and U15781 (N_15781,N_13904,N_14460);
or U15782 (N_15782,N_14951,N_12698);
nand U15783 (N_15783,N_14998,N_12642);
nand U15784 (N_15784,N_13573,N_13558);
and U15785 (N_15785,N_13892,N_13530);
nand U15786 (N_15786,N_14396,N_12904);
and U15787 (N_15787,N_14397,N_12890);
nor U15788 (N_15788,N_14248,N_14111);
nand U15789 (N_15789,N_13654,N_14450);
nor U15790 (N_15790,N_12864,N_14955);
and U15791 (N_15791,N_14848,N_14214);
and U15792 (N_15792,N_14144,N_12692);
nor U15793 (N_15793,N_14800,N_13118);
nand U15794 (N_15794,N_14743,N_13046);
nor U15795 (N_15795,N_14712,N_14124);
and U15796 (N_15796,N_14053,N_14590);
and U15797 (N_15797,N_14622,N_13677);
nor U15798 (N_15798,N_13217,N_14824);
xor U15799 (N_15799,N_12862,N_14851);
or U15800 (N_15800,N_12919,N_12643);
nor U15801 (N_15801,N_13014,N_14007);
nor U15802 (N_15802,N_12523,N_13849);
and U15803 (N_15803,N_14288,N_14244);
nor U15804 (N_15804,N_14393,N_13458);
nor U15805 (N_15805,N_13263,N_13916);
xor U15806 (N_15806,N_13024,N_13911);
and U15807 (N_15807,N_12849,N_14324);
and U15808 (N_15808,N_13183,N_14403);
and U15809 (N_15809,N_13437,N_13310);
nand U15810 (N_15810,N_13797,N_12949);
xor U15811 (N_15811,N_14065,N_13526);
nor U15812 (N_15812,N_12927,N_12578);
nand U15813 (N_15813,N_12637,N_14212);
or U15814 (N_15814,N_12898,N_14758);
nor U15815 (N_15815,N_14659,N_12973);
nor U15816 (N_15816,N_12829,N_14916);
nand U15817 (N_15817,N_14786,N_14086);
nand U15818 (N_15818,N_12525,N_14411);
nand U15819 (N_15819,N_12817,N_14765);
and U15820 (N_15820,N_12503,N_12758);
nor U15821 (N_15821,N_14196,N_14140);
nor U15822 (N_15822,N_13033,N_14354);
nand U15823 (N_15823,N_12601,N_14551);
and U15824 (N_15824,N_13481,N_14734);
and U15825 (N_15825,N_13557,N_13055);
nor U15826 (N_15826,N_14040,N_14222);
nand U15827 (N_15827,N_13429,N_14592);
or U15828 (N_15828,N_12863,N_14612);
and U15829 (N_15829,N_14899,N_13910);
xnor U15830 (N_15830,N_13880,N_13053);
nand U15831 (N_15831,N_14707,N_14114);
and U15832 (N_15832,N_14888,N_13163);
nor U15833 (N_15833,N_13616,N_12879);
or U15834 (N_15834,N_13265,N_12920);
nand U15835 (N_15835,N_14435,N_13387);
or U15836 (N_15836,N_14660,N_14560);
and U15837 (N_15837,N_14538,N_14388);
or U15838 (N_15838,N_13207,N_12564);
or U15839 (N_15839,N_14578,N_14365);
nand U15840 (N_15840,N_13977,N_14515);
nand U15841 (N_15841,N_14468,N_13503);
nor U15842 (N_15842,N_13719,N_13505);
nor U15843 (N_15843,N_12602,N_14901);
nand U15844 (N_15844,N_13174,N_14338);
and U15845 (N_15845,N_14462,N_13312);
nor U15846 (N_15846,N_13135,N_12625);
nand U15847 (N_15847,N_13368,N_14378);
or U15848 (N_15848,N_13374,N_13332);
nand U15849 (N_15849,N_12557,N_13846);
and U15850 (N_15850,N_13016,N_13328);
or U15851 (N_15851,N_13247,N_12647);
nor U15852 (N_15852,N_12819,N_13592);
or U15853 (N_15853,N_13077,N_13568);
nand U15854 (N_15854,N_14349,N_13065);
and U15855 (N_15855,N_14127,N_14246);
nand U15856 (N_15856,N_13732,N_14910);
and U15857 (N_15857,N_12912,N_13888);
nor U15858 (N_15858,N_12628,N_14629);
nor U15859 (N_15859,N_13599,N_14655);
nor U15860 (N_15860,N_14686,N_14326);
and U15861 (N_15861,N_14199,N_13373);
or U15862 (N_15862,N_13707,N_13362);
nor U15863 (N_15863,N_14687,N_13164);
nand U15864 (N_15864,N_13249,N_12804);
and U15865 (N_15865,N_13760,N_13882);
and U15866 (N_15866,N_13202,N_13847);
nand U15867 (N_15867,N_12519,N_14195);
nor U15868 (N_15868,N_14158,N_14651);
nor U15869 (N_15869,N_12988,N_13868);
and U15870 (N_15870,N_13561,N_14635);
nor U15871 (N_15871,N_12566,N_13731);
or U15872 (N_15872,N_12768,N_12605);
nand U15873 (N_15873,N_13234,N_14090);
and U15874 (N_15874,N_13502,N_13186);
nor U15875 (N_15875,N_13461,N_14933);
nand U15876 (N_15876,N_14855,N_13131);
nand U15877 (N_15877,N_13402,N_13160);
and U15878 (N_15878,N_14301,N_12843);
nor U15879 (N_15879,N_12721,N_13818);
and U15880 (N_15880,N_13775,N_14441);
or U15881 (N_15881,N_14553,N_13428);
nor U15882 (N_15882,N_13985,N_14351);
nor U15883 (N_15883,N_14871,N_14446);
and U15884 (N_15884,N_14753,N_13399);
or U15885 (N_15885,N_14459,N_12537);
or U15886 (N_15886,N_14220,N_13242);
or U15887 (N_15887,N_14805,N_14492);
nand U15888 (N_15888,N_12591,N_12702);
and U15889 (N_15889,N_13397,N_14669);
nor U15890 (N_15890,N_13141,N_12950);
nor U15891 (N_15891,N_14293,N_14763);
nor U15892 (N_15892,N_14476,N_12597);
nand U15893 (N_15893,N_14442,N_13487);
or U15894 (N_15894,N_12878,N_14873);
nor U15895 (N_15895,N_14162,N_13441);
or U15896 (N_15896,N_12516,N_13314);
nor U15897 (N_15897,N_14231,N_12928);
or U15898 (N_15898,N_12674,N_13177);
nor U15899 (N_15899,N_13056,N_14356);
nand U15900 (N_15900,N_14475,N_12586);
nor U15901 (N_15901,N_14003,N_12820);
nor U15902 (N_15902,N_13383,N_14054);
nand U15903 (N_15903,N_12593,N_13286);
nand U15904 (N_15904,N_14658,N_14574);
and U15905 (N_15905,N_13371,N_13567);
and U15906 (N_15906,N_14732,N_13442);
or U15907 (N_15907,N_12545,N_14727);
nor U15908 (N_15908,N_14656,N_13419);
or U15909 (N_15909,N_14269,N_13050);
and U15910 (N_15910,N_13769,N_13976);
and U15911 (N_15911,N_13765,N_12570);
or U15912 (N_15912,N_13094,N_14079);
xor U15913 (N_15913,N_14146,N_13542);
nand U15914 (N_15914,N_14919,N_12782);
and U15915 (N_15915,N_14976,N_14627);
or U15916 (N_15916,N_13555,N_14833);
xor U15917 (N_15917,N_13022,N_13225);
nor U15918 (N_15918,N_13070,N_13353);
and U15919 (N_15919,N_14835,N_14572);
nand U15920 (N_15920,N_14009,N_12786);
nand U15921 (N_15921,N_13656,N_14284);
and U15922 (N_15922,N_14940,N_14495);
or U15923 (N_15923,N_14788,N_12514);
and U15924 (N_15924,N_14157,N_12664);
xnor U15925 (N_15925,N_13325,N_12668);
or U15926 (N_15926,N_13179,N_14810);
and U15927 (N_15927,N_14566,N_12977);
nor U15928 (N_15928,N_14959,N_12665);
and U15929 (N_15929,N_14097,N_13907);
nand U15930 (N_15930,N_14698,N_13292);
and U15931 (N_15931,N_14469,N_12611);
nand U15932 (N_15932,N_14739,N_14091);
nand U15933 (N_15933,N_14580,N_13277);
and U15934 (N_15934,N_13848,N_12615);
or U15935 (N_15935,N_14273,N_13529);
and U15936 (N_15936,N_13122,N_14742);
nor U15937 (N_15937,N_13795,N_13037);
nor U15938 (N_15938,N_12764,N_14630);
nor U15939 (N_15939,N_12727,N_12867);
nor U15940 (N_15940,N_13194,N_14019);
nand U15941 (N_15941,N_14846,N_14994);
or U15942 (N_15942,N_13375,N_13384);
xor U15943 (N_15943,N_14736,N_14991);
or U15944 (N_15944,N_14479,N_14331);
nand U15945 (N_15945,N_13774,N_13040);
nor U15946 (N_15946,N_12763,N_14485);
nand U15947 (N_15947,N_14182,N_12895);
nor U15948 (N_15948,N_13802,N_13984);
and U15949 (N_15949,N_13905,N_14292);
and U15950 (N_15950,N_13790,N_13946);
and U15951 (N_15951,N_12766,N_13603);
and U15952 (N_15952,N_13571,N_13883);
and U15953 (N_15953,N_13566,N_14755);
nor U15954 (N_15954,N_14517,N_13667);
nand U15955 (N_15955,N_12933,N_14006);
or U15956 (N_15956,N_12846,N_14565);
or U15957 (N_15957,N_13873,N_13372);
or U15958 (N_15958,N_13096,N_14633);
xnor U15959 (N_15959,N_13279,N_14926);
and U15960 (N_15960,N_14782,N_12649);
or U15961 (N_15961,N_13771,N_13866);
or U15962 (N_15962,N_13228,N_12958);
nand U15963 (N_15963,N_13440,N_12970);
nand U15964 (N_15964,N_14564,N_13173);
or U15965 (N_15965,N_14850,N_12891);
and U15966 (N_15966,N_12688,N_13570);
and U15967 (N_15967,N_13008,N_14037);
xnor U15968 (N_15968,N_14465,N_12957);
or U15969 (N_15969,N_13233,N_12569);
nor U15970 (N_15970,N_14567,N_14232);
and U15971 (N_15971,N_14983,N_12929);
nand U15972 (N_15972,N_14586,N_13854);
and U15973 (N_15973,N_12693,N_12765);
or U15974 (N_15974,N_12983,N_14026);
or U15975 (N_15975,N_12959,N_12745);
nor U15976 (N_15976,N_13357,N_14419);
nand U15977 (N_15977,N_13006,N_13305);
nand U15978 (N_15978,N_14258,N_14089);
xor U15979 (N_15979,N_13793,N_14830);
nor U15980 (N_15980,N_14624,N_14975);
and U15981 (N_15981,N_13280,N_13244);
or U15982 (N_15982,N_14020,N_14569);
and U15983 (N_15983,N_14336,N_12974);
and U15984 (N_15984,N_13059,N_12732);
and U15985 (N_15985,N_13073,N_13425);
or U15986 (N_15986,N_13528,N_13203);
xor U15987 (N_15987,N_14997,N_13748);
nor U15988 (N_15988,N_14543,N_13824);
nand U15989 (N_15989,N_13569,N_14327);
or U15990 (N_15990,N_14434,N_13391);
xnor U15991 (N_15991,N_14023,N_14092);
nor U15992 (N_15992,N_12521,N_14890);
nor U15993 (N_15993,N_12613,N_14045);
or U15994 (N_15994,N_14540,N_13726);
xor U15995 (N_15995,N_13577,N_13551);
xor U15996 (N_15996,N_13683,N_13219);
nor U15997 (N_15997,N_13605,N_12751);
xnor U15998 (N_15998,N_13051,N_12561);
and U15999 (N_15999,N_14649,N_13253);
and U16000 (N_16000,N_14126,N_14898);
xnor U16001 (N_16001,N_13414,N_14502);
xor U16002 (N_16002,N_13514,N_13088);
xnor U16003 (N_16003,N_13532,N_13470);
and U16004 (N_16004,N_13702,N_12614);
nand U16005 (N_16005,N_12769,N_13805);
nor U16006 (N_16006,N_13758,N_14639);
and U16007 (N_16007,N_12884,N_13155);
nand U16008 (N_16008,N_13659,N_13257);
or U16009 (N_16009,N_12678,N_14506);
and U16010 (N_16010,N_13852,N_13647);
nand U16011 (N_16011,N_14047,N_13018);
nor U16012 (N_16012,N_14482,N_12810);
and U16013 (N_16013,N_13182,N_14829);
or U16014 (N_16014,N_14402,N_14646);
or U16015 (N_16015,N_13794,N_13408);
and U16016 (N_16016,N_13283,N_14320);
or U16017 (N_16017,N_14368,N_14012);
or U16018 (N_16018,N_14039,N_13262);
or U16019 (N_16019,N_14494,N_13942);
nand U16020 (N_16020,N_14387,N_13291);
or U16021 (N_16021,N_13741,N_14802);
and U16022 (N_16022,N_14394,N_13349);
nand U16023 (N_16023,N_13938,N_12841);
and U16024 (N_16024,N_14243,N_14784);
and U16025 (N_16025,N_13303,N_13343);
nor U16026 (N_16026,N_12551,N_14879);
nor U16027 (N_16027,N_14255,N_13061);
xor U16028 (N_16028,N_14254,N_12997);
or U16029 (N_16029,N_14603,N_13810);
and U16030 (N_16030,N_13768,N_13896);
nand U16031 (N_16031,N_14414,N_13544);
and U16032 (N_16032,N_13124,N_14370);
nor U16033 (N_16033,N_13800,N_12798);
and U16034 (N_16034,N_13608,N_12547);
or U16035 (N_16035,N_13618,N_12893);
or U16036 (N_16036,N_14870,N_12995);
nor U16037 (N_16037,N_14508,N_14297);
xnor U16038 (N_16038,N_13778,N_12724);
nand U16039 (N_16039,N_13644,N_14518);
or U16040 (N_16040,N_13150,N_13665);
and U16041 (N_16041,N_12978,N_14947);
xor U16042 (N_16042,N_14307,N_14973);
and U16043 (N_16043,N_13565,N_14458);
or U16044 (N_16044,N_14188,N_14062);
or U16045 (N_16045,N_13685,N_13917);
nand U16046 (N_16046,N_12901,N_13853);
nand U16047 (N_16047,N_13931,N_13147);
xnor U16048 (N_16048,N_14812,N_12791);
and U16049 (N_16049,N_13091,N_14679);
nor U16050 (N_16050,N_13913,N_14489);
nand U16051 (N_16051,N_14279,N_13210);
or U16052 (N_16052,N_14773,N_12873);
and U16053 (N_16053,N_14971,N_13744);
and U16054 (N_16054,N_13267,N_13643);
nand U16055 (N_16055,N_14647,N_14840);
nor U16056 (N_16056,N_14738,N_13294);
or U16057 (N_16057,N_13753,N_12812);
xor U16058 (N_16058,N_13681,N_14694);
xnor U16059 (N_16059,N_14668,N_13833);
and U16060 (N_16060,N_13227,N_14801);
or U16061 (N_16061,N_13333,N_14189);
or U16062 (N_16062,N_13661,N_13767);
nand U16063 (N_16063,N_13152,N_12581);
nor U16064 (N_16064,N_13928,N_12616);
or U16065 (N_16065,N_13811,N_14205);
nand U16066 (N_16066,N_13899,N_14673);
and U16067 (N_16067,N_14433,N_12680);
nor U16068 (N_16068,N_12629,N_14008);
nor U16069 (N_16069,N_12940,N_12835);
or U16070 (N_16070,N_12720,N_14769);
and U16071 (N_16071,N_13076,N_14210);
nand U16072 (N_16072,N_13424,N_14120);
nand U16073 (N_16073,N_13590,N_13952);
and U16074 (N_16074,N_13347,N_13255);
nor U16075 (N_16075,N_14798,N_13195);
nand U16076 (N_16076,N_14925,N_13261);
nand U16077 (N_16077,N_14339,N_13979);
xnor U16078 (N_16078,N_13492,N_13713);
or U16079 (N_16079,N_14311,N_13745);
nand U16080 (N_16080,N_13300,N_14117);
nor U16081 (N_16081,N_14175,N_14839);
nand U16082 (N_16082,N_13358,N_12784);
or U16083 (N_16083,N_14242,N_14342);
nand U16084 (N_16084,N_13057,N_12877);
and U16085 (N_16085,N_13092,N_13861);
nor U16086 (N_16086,N_14505,N_14287);
nand U16087 (N_16087,N_13236,N_13151);
and U16088 (N_16088,N_12598,N_13610);
and U16089 (N_16089,N_13714,N_14990);
xor U16090 (N_16090,N_13009,N_13912);
nor U16091 (N_16091,N_12998,N_13658);
and U16092 (N_16092,N_13876,N_14923);
or U16093 (N_16093,N_14406,N_13842);
xor U16094 (N_16094,N_13651,N_12931);
nor U16095 (N_16095,N_14794,N_14556);
or U16096 (N_16096,N_13562,N_14138);
or U16097 (N_16097,N_13005,N_13400);
nor U16098 (N_16098,N_12905,N_14900);
nor U16099 (N_16099,N_13042,N_14197);
nand U16100 (N_16100,N_12562,N_12708);
xor U16101 (N_16101,N_14449,N_13100);
nand U16102 (N_16102,N_13398,N_13559);
nand U16103 (N_16103,N_14029,N_13081);
nor U16104 (N_16104,N_14361,N_14945);
and U16105 (N_16105,N_12659,N_14552);
and U16106 (N_16106,N_12684,N_14614);
nor U16107 (N_16107,N_13495,N_14082);
nor U16108 (N_16108,N_14315,N_13890);
and U16109 (N_16109,N_14364,N_13836);
and U16110 (N_16110,N_13783,N_12536);
nor U16111 (N_16111,N_14512,N_14366);
nor U16112 (N_16112,N_13845,N_14914);
or U16113 (N_16113,N_14577,N_14498);
nor U16114 (N_16114,N_14116,N_13978);
nor U16115 (N_16115,N_14206,N_13128);
xor U16116 (N_16116,N_13496,N_14137);
nand U16117 (N_16117,N_13579,N_14814);
nor U16118 (N_16118,N_13344,N_13078);
and U16119 (N_16119,N_14984,N_13993);
nand U16120 (N_16120,N_12539,N_13879);
and U16121 (N_16121,N_12600,N_14606);
or U16122 (N_16122,N_14642,N_14163);
or U16123 (N_16123,N_13071,N_14557);
nor U16124 (N_16124,N_14247,N_13695);
nand U16125 (N_16125,N_13622,N_14055);
and U16126 (N_16126,N_14526,N_14497);
and U16127 (N_16127,N_12964,N_13550);
nor U16128 (N_16128,N_14828,N_12979);
nor U16129 (N_16129,N_13927,N_14932);
nand U16130 (N_16130,N_12900,N_12730);
nor U16131 (N_16131,N_14102,N_12981);
nor U16132 (N_16132,N_13697,N_13404);
nand U16133 (N_16133,N_14549,N_12737);
nor U16134 (N_16134,N_14483,N_13112);
xnor U16135 (N_16135,N_14384,N_14866);
xnor U16136 (N_16136,N_14643,N_14902);
nor U16137 (N_16137,N_13752,N_14616);
nand U16138 (N_16138,N_12652,N_13956);
nor U16139 (N_16139,N_14104,N_13304);
and U16140 (N_16140,N_14329,N_12699);
nor U16141 (N_16141,N_13670,N_13130);
or U16142 (N_16142,N_14653,N_13909);
or U16143 (N_16143,N_14504,N_12515);
nand U16144 (N_16144,N_12828,N_14296);
nor U16145 (N_16145,N_12894,N_12876);
nand U16146 (N_16146,N_14918,N_12955);
or U16147 (N_16147,N_13867,N_13699);
and U16148 (N_16148,N_14831,N_13099);
nor U16149 (N_16149,N_13641,N_12711);
nand U16150 (N_16150,N_14291,N_13275);
and U16151 (N_16151,N_13575,N_14099);
or U16152 (N_16152,N_13176,N_13444);
nand U16153 (N_16153,N_12735,N_13710);
nand U16154 (N_16154,N_14302,N_14437);
and U16155 (N_16155,N_13296,N_12939);
nand U16156 (N_16156,N_13184,N_13604);
or U16157 (N_16157,N_14225,N_14063);
nor U16158 (N_16158,N_14995,N_13220);
nor U16159 (N_16159,N_13621,N_14548);
or U16160 (N_16160,N_14819,N_13814);
nor U16161 (N_16161,N_12728,N_14226);
nand U16162 (N_16162,N_14597,N_12742);
xor U16163 (N_16163,N_12897,N_12935);
and U16164 (N_16164,N_12951,N_14347);
or U16165 (N_16165,N_12993,N_13675);
and U16166 (N_16166,N_14905,N_12560);
nand U16167 (N_16167,N_12881,N_13813);
and U16168 (N_16168,N_13000,N_13087);
nand U16169 (N_16169,N_14101,N_13948);
or U16170 (N_16170,N_14211,N_12956);
xor U16171 (N_16171,N_12823,N_13930);
or U16172 (N_16172,N_13680,N_14004);
or U16173 (N_16173,N_14607,N_13465);
nand U16174 (N_16174,N_12815,N_13204);
or U16175 (N_16175,N_14733,N_12827);
and U16176 (N_16176,N_12787,N_14613);
or U16177 (N_16177,N_12644,N_14715);
nor U16178 (N_16178,N_14233,N_14783);
or U16179 (N_16179,N_13086,N_13638);
nor U16180 (N_16180,N_12506,N_12517);
nand U16181 (N_16181,N_13856,N_13591);
and U16182 (N_16182,N_13416,N_14056);
nor U16183 (N_16183,N_14617,N_13451);
and U16184 (N_16184,N_13954,N_12510);
nand U16185 (N_16185,N_13409,N_14544);
nor U16186 (N_16186,N_12975,N_13613);
and U16187 (N_16187,N_14760,N_14151);
or U16188 (N_16188,N_14136,N_13611);
and U16189 (N_16189,N_14807,N_13785);
nor U16190 (N_16190,N_12646,N_14191);
nor U16191 (N_16191,N_14748,N_13342);
nand U16192 (N_16192,N_14272,N_14179);
nor U16193 (N_16193,N_13415,N_13773);
xor U16194 (N_16194,N_14186,N_14981);
xnor U16195 (N_16195,N_12696,N_12650);
nor U16196 (N_16196,N_14223,N_13443);
xnor U16197 (N_16197,N_13256,N_13290);
nand U16198 (N_16198,N_13779,N_13396);
nor U16199 (N_16199,N_13857,N_13855);
nor U16200 (N_16200,N_13789,N_12687);
or U16201 (N_16201,N_13044,N_12832);
and U16202 (N_16202,N_13154,N_14547);
xnor U16203 (N_16203,N_13556,N_12627);
and U16204 (N_16204,N_14558,N_14410);
nor U16205 (N_16205,N_14683,N_12544);
and U16206 (N_16206,N_14085,N_14723);
nand U16207 (N_16207,N_12865,N_14503);
nor U16208 (N_16208,N_13321,N_14049);
or U16209 (N_16209,N_14264,N_13287);
and U16210 (N_16210,N_13871,N_14185);
and U16211 (N_16211,N_13335,N_13844);
or U16212 (N_16212,N_14488,N_13113);
or U16213 (N_16213,N_14129,N_13463);
or U16214 (N_16214,N_13331,N_14355);
and U16215 (N_16215,N_14278,N_14972);
or U16216 (N_16216,N_13486,N_14935);
nand U16217 (N_16217,N_12670,N_13169);
nand U16218 (N_16218,N_13723,N_14262);
or U16219 (N_16219,N_13640,N_14582);
and U16220 (N_16220,N_13947,N_14061);
nand U16221 (N_16221,N_14500,N_14958);
nand U16222 (N_16222,N_12814,N_14015);
nand U16223 (N_16223,N_13838,N_12731);
nor U16224 (N_16224,N_13698,N_12526);
or U16225 (N_16225,N_13962,N_13674);
and U16226 (N_16226,N_13507,N_13223);
nor U16227 (N_16227,N_14964,N_13080);
nor U16228 (N_16228,N_13361,N_13214);
nand U16229 (N_16229,N_14685,N_13017);
or U16230 (N_16230,N_12604,N_13127);
or U16231 (N_16231,N_14295,N_13520);
nor U16232 (N_16232,N_12582,N_12811);
and U16233 (N_16233,N_13175,N_12954);
and U16234 (N_16234,N_14977,N_14052);
and U16235 (N_16235,N_13259,N_13742);
nor U16236 (N_16236,N_13521,N_14640);
xnor U16237 (N_16237,N_14664,N_12872);
and U16238 (N_16238,N_14746,N_14000);
or U16239 (N_16239,N_14133,N_14884);
nand U16240 (N_16240,N_14112,N_12657);
and U16241 (N_16241,N_13365,N_12793);
nand U16242 (N_16242,N_12624,N_12777);
or U16243 (N_16243,N_13648,N_13412);
nor U16244 (N_16244,N_14119,N_13691);
nand U16245 (N_16245,N_14593,N_12747);
and U16246 (N_16246,N_13944,N_13129);
xnor U16247 (N_16247,N_13787,N_13588);
and U16248 (N_16248,N_14002,N_14028);
nor U16249 (N_16249,N_14033,N_13105);
or U16250 (N_16250,N_13328,N_13500);
or U16251 (N_16251,N_12598,N_14569);
and U16252 (N_16252,N_14327,N_13460);
and U16253 (N_16253,N_13949,N_14193);
xnor U16254 (N_16254,N_14451,N_12672);
and U16255 (N_16255,N_12634,N_14050);
and U16256 (N_16256,N_14044,N_14066);
nor U16257 (N_16257,N_13506,N_13653);
nor U16258 (N_16258,N_13721,N_13487);
xor U16259 (N_16259,N_14699,N_13154);
and U16260 (N_16260,N_13409,N_12649);
nand U16261 (N_16261,N_14130,N_13781);
nor U16262 (N_16262,N_12503,N_12900);
nor U16263 (N_16263,N_13379,N_14765);
nand U16264 (N_16264,N_13338,N_14784);
or U16265 (N_16265,N_14247,N_13571);
xnor U16266 (N_16266,N_12782,N_13765);
xor U16267 (N_16267,N_12677,N_13744);
nand U16268 (N_16268,N_14935,N_14590);
xnor U16269 (N_16269,N_14771,N_13323);
nand U16270 (N_16270,N_12685,N_14393);
nand U16271 (N_16271,N_14110,N_12646);
or U16272 (N_16272,N_13463,N_14001);
nor U16273 (N_16273,N_14471,N_13255);
and U16274 (N_16274,N_13169,N_14919);
xor U16275 (N_16275,N_14332,N_12739);
nand U16276 (N_16276,N_14818,N_12737);
nor U16277 (N_16277,N_13925,N_13802);
or U16278 (N_16278,N_12607,N_12876);
nand U16279 (N_16279,N_12905,N_13578);
and U16280 (N_16280,N_13495,N_14465);
and U16281 (N_16281,N_13883,N_12677);
nand U16282 (N_16282,N_12645,N_14900);
or U16283 (N_16283,N_13063,N_13622);
nor U16284 (N_16284,N_12925,N_13154);
or U16285 (N_16285,N_14976,N_14130);
or U16286 (N_16286,N_14690,N_12699);
or U16287 (N_16287,N_12797,N_14293);
nor U16288 (N_16288,N_13119,N_14646);
xor U16289 (N_16289,N_14391,N_13459);
nand U16290 (N_16290,N_12977,N_14016);
nand U16291 (N_16291,N_13980,N_14413);
or U16292 (N_16292,N_13259,N_14491);
or U16293 (N_16293,N_14102,N_14179);
nor U16294 (N_16294,N_13526,N_14361);
and U16295 (N_16295,N_13396,N_13599);
and U16296 (N_16296,N_13579,N_14568);
xor U16297 (N_16297,N_13397,N_13555);
nand U16298 (N_16298,N_14783,N_13274);
nand U16299 (N_16299,N_13957,N_14676);
nor U16300 (N_16300,N_14884,N_13792);
and U16301 (N_16301,N_12921,N_14266);
nand U16302 (N_16302,N_13721,N_13312);
nand U16303 (N_16303,N_12556,N_12955);
nand U16304 (N_16304,N_13561,N_14049);
nand U16305 (N_16305,N_14253,N_14114);
nand U16306 (N_16306,N_14956,N_14357);
nand U16307 (N_16307,N_14175,N_13361);
or U16308 (N_16308,N_13065,N_13331);
nor U16309 (N_16309,N_13031,N_13734);
nor U16310 (N_16310,N_12836,N_14859);
nand U16311 (N_16311,N_12846,N_13192);
nand U16312 (N_16312,N_13700,N_14526);
or U16313 (N_16313,N_14785,N_14779);
nor U16314 (N_16314,N_12938,N_12728);
or U16315 (N_16315,N_14106,N_13362);
nand U16316 (N_16316,N_14091,N_14930);
and U16317 (N_16317,N_13780,N_12687);
and U16318 (N_16318,N_14869,N_13698);
xnor U16319 (N_16319,N_14977,N_13671);
xor U16320 (N_16320,N_13924,N_12919);
and U16321 (N_16321,N_12578,N_13288);
xnor U16322 (N_16322,N_13709,N_13974);
or U16323 (N_16323,N_12592,N_14614);
nor U16324 (N_16324,N_14804,N_14386);
or U16325 (N_16325,N_14070,N_14334);
nor U16326 (N_16326,N_12643,N_12997);
nand U16327 (N_16327,N_14959,N_12614);
or U16328 (N_16328,N_13014,N_14401);
and U16329 (N_16329,N_14771,N_13202);
and U16330 (N_16330,N_13746,N_13179);
nand U16331 (N_16331,N_14286,N_13481);
xor U16332 (N_16332,N_12873,N_14605);
nor U16333 (N_16333,N_13095,N_14395);
nor U16334 (N_16334,N_14407,N_14168);
and U16335 (N_16335,N_13944,N_14451);
or U16336 (N_16336,N_12607,N_13137);
nand U16337 (N_16337,N_14582,N_13109);
or U16338 (N_16338,N_12708,N_12922);
and U16339 (N_16339,N_13489,N_14263);
nor U16340 (N_16340,N_14378,N_13662);
nand U16341 (N_16341,N_14540,N_12758);
nor U16342 (N_16342,N_13113,N_13516);
xor U16343 (N_16343,N_13673,N_13867);
or U16344 (N_16344,N_12682,N_14183);
or U16345 (N_16345,N_12593,N_14321);
or U16346 (N_16346,N_14053,N_13130);
or U16347 (N_16347,N_14484,N_13071);
nor U16348 (N_16348,N_12682,N_13505);
nor U16349 (N_16349,N_13348,N_13226);
and U16350 (N_16350,N_13136,N_13695);
nor U16351 (N_16351,N_14526,N_14082);
and U16352 (N_16352,N_14859,N_13655);
xor U16353 (N_16353,N_14627,N_12906);
nand U16354 (N_16354,N_13078,N_13340);
nor U16355 (N_16355,N_14785,N_12975);
or U16356 (N_16356,N_13572,N_13695);
or U16357 (N_16357,N_14721,N_14881);
and U16358 (N_16358,N_14177,N_14831);
or U16359 (N_16359,N_13619,N_14651);
or U16360 (N_16360,N_14993,N_14673);
and U16361 (N_16361,N_13128,N_13809);
and U16362 (N_16362,N_13839,N_12838);
and U16363 (N_16363,N_12674,N_12508);
and U16364 (N_16364,N_13698,N_12848);
xnor U16365 (N_16365,N_14857,N_12519);
and U16366 (N_16366,N_14150,N_13723);
nor U16367 (N_16367,N_13342,N_14507);
xor U16368 (N_16368,N_13929,N_14865);
or U16369 (N_16369,N_13928,N_14100);
or U16370 (N_16370,N_14372,N_12683);
or U16371 (N_16371,N_13293,N_14020);
and U16372 (N_16372,N_14260,N_14571);
and U16373 (N_16373,N_12654,N_14460);
and U16374 (N_16374,N_13846,N_14978);
nor U16375 (N_16375,N_14971,N_12582);
nand U16376 (N_16376,N_13396,N_14379);
and U16377 (N_16377,N_12843,N_13320);
nand U16378 (N_16378,N_13141,N_14325);
and U16379 (N_16379,N_14075,N_12901);
or U16380 (N_16380,N_14439,N_13179);
nor U16381 (N_16381,N_14986,N_12597);
nor U16382 (N_16382,N_13715,N_13933);
nand U16383 (N_16383,N_13874,N_13106);
and U16384 (N_16384,N_14253,N_14325);
or U16385 (N_16385,N_14318,N_13453);
or U16386 (N_16386,N_13267,N_14746);
or U16387 (N_16387,N_13864,N_14384);
nor U16388 (N_16388,N_13602,N_13712);
nor U16389 (N_16389,N_13700,N_12805);
and U16390 (N_16390,N_13756,N_13790);
and U16391 (N_16391,N_13712,N_13446);
or U16392 (N_16392,N_14694,N_13219);
nand U16393 (N_16393,N_12994,N_13312);
nor U16394 (N_16394,N_14611,N_13499);
or U16395 (N_16395,N_14659,N_14114);
and U16396 (N_16396,N_13825,N_13299);
and U16397 (N_16397,N_12598,N_13082);
xor U16398 (N_16398,N_14780,N_13746);
xor U16399 (N_16399,N_13672,N_13002);
or U16400 (N_16400,N_13398,N_13309);
nor U16401 (N_16401,N_12863,N_13323);
nand U16402 (N_16402,N_14148,N_12718);
and U16403 (N_16403,N_13773,N_14589);
xnor U16404 (N_16404,N_12837,N_12555);
xor U16405 (N_16405,N_14520,N_14304);
nand U16406 (N_16406,N_14537,N_14660);
or U16407 (N_16407,N_13374,N_13888);
and U16408 (N_16408,N_13842,N_13321);
or U16409 (N_16409,N_13157,N_13260);
nor U16410 (N_16410,N_14459,N_13871);
nor U16411 (N_16411,N_13510,N_13173);
xor U16412 (N_16412,N_14387,N_13917);
or U16413 (N_16413,N_12779,N_12627);
and U16414 (N_16414,N_14673,N_14444);
xnor U16415 (N_16415,N_12608,N_13672);
xnor U16416 (N_16416,N_13332,N_14877);
nor U16417 (N_16417,N_14052,N_14289);
and U16418 (N_16418,N_13221,N_14566);
nand U16419 (N_16419,N_14027,N_14164);
or U16420 (N_16420,N_13421,N_12504);
nand U16421 (N_16421,N_13964,N_14899);
nor U16422 (N_16422,N_14542,N_12752);
or U16423 (N_16423,N_12549,N_12924);
nor U16424 (N_16424,N_13130,N_14349);
xnor U16425 (N_16425,N_13818,N_14773);
xor U16426 (N_16426,N_13773,N_13395);
xnor U16427 (N_16427,N_14355,N_13932);
nand U16428 (N_16428,N_14937,N_13257);
nor U16429 (N_16429,N_13962,N_14502);
and U16430 (N_16430,N_14887,N_13992);
nor U16431 (N_16431,N_13351,N_12862);
and U16432 (N_16432,N_12999,N_12610);
and U16433 (N_16433,N_13683,N_12955);
nand U16434 (N_16434,N_12831,N_14735);
or U16435 (N_16435,N_14923,N_13202);
and U16436 (N_16436,N_14862,N_14485);
nor U16437 (N_16437,N_13841,N_12591);
or U16438 (N_16438,N_14279,N_13873);
or U16439 (N_16439,N_14302,N_14743);
and U16440 (N_16440,N_12974,N_13920);
and U16441 (N_16441,N_13468,N_14589);
and U16442 (N_16442,N_13244,N_13085);
nand U16443 (N_16443,N_14818,N_12548);
and U16444 (N_16444,N_14731,N_14196);
xnor U16445 (N_16445,N_12812,N_12724);
xnor U16446 (N_16446,N_13031,N_13105);
nor U16447 (N_16447,N_13715,N_14473);
xnor U16448 (N_16448,N_13131,N_14490);
nand U16449 (N_16449,N_13322,N_14466);
nand U16450 (N_16450,N_13551,N_13909);
and U16451 (N_16451,N_13755,N_13988);
or U16452 (N_16452,N_13718,N_14430);
nand U16453 (N_16453,N_14924,N_13673);
xor U16454 (N_16454,N_14906,N_13009);
nand U16455 (N_16455,N_13914,N_12942);
and U16456 (N_16456,N_12576,N_12904);
nand U16457 (N_16457,N_14176,N_13321);
xor U16458 (N_16458,N_12510,N_13890);
and U16459 (N_16459,N_14076,N_13824);
nand U16460 (N_16460,N_13972,N_14489);
xor U16461 (N_16461,N_14012,N_13478);
nand U16462 (N_16462,N_12925,N_13947);
or U16463 (N_16463,N_13429,N_12977);
and U16464 (N_16464,N_13832,N_13595);
and U16465 (N_16465,N_13789,N_13800);
nor U16466 (N_16466,N_14422,N_14609);
and U16467 (N_16467,N_13506,N_14932);
or U16468 (N_16468,N_13667,N_14117);
or U16469 (N_16469,N_12799,N_12588);
or U16470 (N_16470,N_14003,N_13845);
or U16471 (N_16471,N_13815,N_14057);
nor U16472 (N_16472,N_14313,N_13711);
nor U16473 (N_16473,N_13112,N_14425);
nand U16474 (N_16474,N_14240,N_13419);
or U16475 (N_16475,N_13695,N_12753);
nor U16476 (N_16476,N_13425,N_13135);
nand U16477 (N_16477,N_12551,N_14830);
or U16478 (N_16478,N_13364,N_12677);
nand U16479 (N_16479,N_13767,N_13225);
and U16480 (N_16480,N_13263,N_13702);
or U16481 (N_16481,N_12802,N_13766);
and U16482 (N_16482,N_13465,N_13856);
xor U16483 (N_16483,N_14802,N_14442);
nor U16484 (N_16484,N_13801,N_13496);
nand U16485 (N_16485,N_13161,N_14965);
nand U16486 (N_16486,N_13630,N_14116);
nor U16487 (N_16487,N_14540,N_14625);
nand U16488 (N_16488,N_14023,N_12596);
xnor U16489 (N_16489,N_13758,N_13280);
nor U16490 (N_16490,N_14316,N_13294);
nor U16491 (N_16491,N_13446,N_13594);
nor U16492 (N_16492,N_14835,N_14180);
nand U16493 (N_16493,N_12722,N_12544);
or U16494 (N_16494,N_14157,N_13152);
xnor U16495 (N_16495,N_13636,N_13710);
nor U16496 (N_16496,N_14852,N_13973);
or U16497 (N_16497,N_14335,N_13933);
xor U16498 (N_16498,N_13529,N_13286);
and U16499 (N_16499,N_14435,N_13847);
nor U16500 (N_16500,N_12725,N_13055);
or U16501 (N_16501,N_14532,N_13909);
nand U16502 (N_16502,N_13119,N_14687);
and U16503 (N_16503,N_13297,N_12756);
nor U16504 (N_16504,N_13926,N_13261);
or U16505 (N_16505,N_13094,N_14710);
nand U16506 (N_16506,N_12519,N_14172);
nor U16507 (N_16507,N_13905,N_14640);
nor U16508 (N_16508,N_14334,N_12618);
nand U16509 (N_16509,N_13605,N_13141);
nor U16510 (N_16510,N_14836,N_12508);
or U16511 (N_16511,N_13187,N_12877);
nor U16512 (N_16512,N_13711,N_12765);
nand U16513 (N_16513,N_13040,N_12559);
and U16514 (N_16514,N_14379,N_12914);
nand U16515 (N_16515,N_14564,N_13498);
nor U16516 (N_16516,N_13325,N_14959);
nor U16517 (N_16517,N_14713,N_13723);
nand U16518 (N_16518,N_13636,N_14603);
nor U16519 (N_16519,N_14802,N_12826);
or U16520 (N_16520,N_13746,N_12979);
nor U16521 (N_16521,N_12644,N_14696);
and U16522 (N_16522,N_13658,N_13417);
nor U16523 (N_16523,N_12998,N_14926);
nor U16524 (N_16524,N_14569,N_13930);
nor U16525 (N_16525,N_14899,N_14379);
or U16526 (N_16526,N_13653,N_14734);
nand U16527 (N_16527,N_14675,N_13079);
and U16528 (N_16528,N_13218,N_12724);
or U16529 (N_16529,N_13820,N_13340);
nand U16530 (N_16530,N_13730,N_12502);
or U16531 (N_16531,N_14126,N_13041);
nand U16532 (N_16532,N_13002,N_12728);
or U16533 (N_16533,N_13488,N_13922);
nor U16534 (N_16534,N_12727,N_14317);
nor U16535 (N_16535,N_14082,N_13005);
nand U16536 (N_16536,N_12687,N_14388);
or U16537 (N_16537,N_13455,N_14365);
nor U16538 (N_16538,N_14676,N_13098);
nand U16539 (N_16539,N_14464,N_13250);
nand U16540 (N_16540,N_14856,N_13236);
xnor U16541 (N_16541,N_14739,N_14727);
nor U16542 (N_16542,N_14363,N_13367);
nand U16543 (N_16543,N_12972,N_14831);
nor U16544 (N_16544,N_13521,N_12509);
and U16545 (N_16545,N_13979,N_12739);
nor U16546 (N_16546,N_12875,N_14500);
nor U16547 (N_16547,N_13819,N_14262);
or U16548 (N_16548,N_13260,N_12603);
or U16549 (N_16549,N_12941,N_14299);
and U16550 (N_16550,N_13967,N_13633);
nand U16551 (N_16551,N_12989,N_13974);
xnor U16552 (N_16552,N_12902,N_12658);
nor U16553 (N_16553,N_13067,N_14634);
nand U16554 (N_16554,N_12545,N_14913);
and U16555 (N_16555,N_13206,N_13204);
xnor U16556 (N_16556,N_14391,N_13869);
and U16557 (N_16557,N_13284,N_14633);
nor U16558 (N_16558,N_14227,N_13552);
nand U16559 (N_16559,N_12787,N_12821);
nor U16560 (N_16560,N_13986,N_12880);
and U16561 (N_16561,N_13393,N_14477);
nor U16562 (N_16562,N_14021,N_14188);
and U16563 (N_16563,N_13176,N_13644);
or U16564 (N_16564,N_13653,N_14961);
or U16565 (N_16565,N_12922,N_14267);
nor U16566 (N_16566,N_12959,N_12887);
nor U16567 (N_16567,N_13534,N_13034);
and U16568 (N_16568,N_13513,N_14491);
nand U16569 (N_16569,N_14604,N_13841);
or U16570 (N_16570,N_13602,N_14764);
or U16571 (N_16571,N_13879,N_14841);
nand U16572 (N_16572,N_13841,N_14067);
and U16573 (N_16573,N_14195,N_12818);
or U16574 (N_16574,N_13933,N_14731);
and U16575 (N_16575,N_13210,N_12881);
xor U16576 (N_16576,N_12999,N_13716);
nor U16577 (N_16577,N_14897,N_13170);
and U16578 (N_16578,N_14421,N_12888);
and U16579 (N_16579,N_12639,N_12942);
or U16580 (N_16580,N_13258,N_13927);
nor U16581 (N_16581,N_13394,N_13885);
and U16582 (N_16582,N_14213,N_14840);
and U16583 (N_16583,N_13964,N_13361);
xnor U16584 (N_16584,N_13035,N_14315);
and U16585 (N_16585,N_14583,N_14322);
nand U16586 (N_16586,N_12808,N_14762);
nor U16587 (N_16587,N_13437,N_12685);
and U16588 (N_16588,N_14408,N_13094);
and U16589 (N_16589,N_14360,N_13838);
xor U16590 (N_16590,N_12654,N_13197);
or U16591 (N_16591,N_12740,N_14062);
or U16592 (N_16592,N_13658,N_13804);
nor U16593 (N_16593,N_12756,N_14253);
or U16594 (N_16594,N_13709,N_12584);
xnor U16595 (N_16595,N_13221,N_12998);
nand U16596 (N_16596,N_13700,N_13675);
or U16597 (N_16597,N_12924,N_13239);
and U16598 (N_16598,N_13099,N_14508);
xnor U16599 (N_16599,N_12930,N_14173);
or U16600 (N_16600,N_14013,N_12922);
or U16601 (N_16601,N_14834,N_13224);
nor U16602 (N_16602,N_14967,N_12548);
nand U16603 (N_16603,N_12567,N_12972);
nor U16604 (N_16604,N_12932,N_12626);
or U16605 (N_16605,N_12761,N_13840);
and U16606 (N_16606,N_14656,N_14183);
nand U16607 (N_16607,N_12672,N_12529);
nand U16608 (N_16608,N_14592,N_14428);
or U16609 (N_16609,N_14367,N_13027);
nand U16610 (N_16610,N_13815,N_13321);
xnor U16611 (N_16611,N_14384,N_14209);
nor U16612 (N_16612,N_13839,N_13900);
or U16613 (N_16613,N_13160,N_14340);
nor U16614 (N_16614,N_13844,N_14136);
and U16615 (N_16615,N_13371,N_13635);
xnor U16616 (N_16616,N_13605,N_13566);
nand U16617 (N_16617,N_14247,N_14409);
and U16618 (N_16618,N_13660,N_13608);
xor U16619 (N_16619,N_12551,N_13512);
or U16620 (N_16620,N_12773,N_14740);
nor U16621 (N_16621,N_14612,N_12588);
xor U16622 (N_16622,N_13193,N_13718);
nor U16623 (N_16623,N_12684,N_12716);
xor U16624 (N_16624,N_12661,N_13618);
nand U16625 (N_16625,N_14120,N_13350);
or U16626 (N_16626,N_13424,N_12962);
nand U16627 (N_16627,N_14029,N_14165);
nor U16628 (N_16628,N_13731,N_14867);
nand U16629 (N_16629,N_12735,N_12915);
nand U16630 (N_16630,N_13443,N_14984);
and U16631 (N_16631,N_14272,N_13737);
and U16632 (N_16632,N_14828,N_14646);
xnor U16633 (N_16633,N_13635,N_14366);
nor U16634 (N_16634,N_12635,N_13862);
and U16635 (N_16635,N_13890,N_13929);
and U16636 (N_16636,N_12810,N_14836);
nand U16637 (N_16637,N_13343,N_14426);
nor U16638 (N_16638,N_13632,N_14959);
or U16639 (N_16639,N_14233,N_13086);
xnor U16640 (N_16640,N_14929,N_14783);
nand U16641 (N_16641,N_14522,N_14219);
or U16642 (N_16642,N_13021,N_14125);
xnor U16643 (N_16643,N_13993,N_12693);
nor U16644 (N_16644,N_13260,N_14385);
or U16645 (N_16645,N_14504,N_12948);
nand U16646 (N_16646,N_13352,N_13476);
or U16647 (N_16647,N_13328,N_13672);
and U16648 (N_16648,N_13076,N_14322);
and U16649 (N_16649,N_12977,N_12656);
nand U16650 (N_16650,N_14447,N_14966);
and U16651 (N_16651,N_13486,N_13174);
nor U16652 (N_16652,N_12915,N_13483);
and U16653 (N_16653,N_12584,N_14657);
nand U16654 (N_16654,N_12903,N_13540);
nand U16655 (N_16655,N_12980,N_13408);
or U16656 (N_16656,N_13418,N_14901);
nor U16657 (N_16657,N_13393,N_13473);
and U16658 (N_16658,N_12661,N_12982);
nor U16659 (N_16659,N_13733,N_13534);
and U16660 (N_16660,N_13621,N_14758);
and U16661 (N_16661,N_13785,N_13128);
or U16662 (N_16662,N_14045,N_14182);
nand U16663 (N_16663,N_14411,N_13769);
and U16664 (N_16664,N_13906,N_14124);
and U16665 (N_16665,N_12734,N_14194);
or U16666 (N_16666,N_13360,N_13963);
nor U16667 (N_16667,N_13708,N_12688);
or U16668 (N_16668,N_13962,N_12816);
and U16669 (N_16669,N_14867,N_14317);
xnor U16670 (N_16670,N_12931,N_13814);
nor U16671 (N_16671,N_14410,N_14275);
nor U16672 (N_16672,N_14096,N_14521);
or U16673 (N_16673,N_14354,N_13261);
nor U16674 (N_16674,N_14857,N_14738);
xor U16675 (N_16675,N_14962,N_14839);
nand U16676 (N_16676,N_14992,N_13908);
nor U16677 (N_16677,N_13384,N_13368);
and U16678 (N_16678,N_13828,N_13756);
nor U16679 (N_16679,N_14840,N_12557);
nor U16680 (N_16680,N_12790,N_13474);
nor U16681 (N_16681,N_14325,N_13013);
nand U16682 (N_16682,N_14249,N_14377);
xor U16683 (N_16683,N_14267,N_14309);
nor U16684 (N_16684,N_13719,N_14011);
and U16685 (N_16685,N_13376,N_12800);
and U16686 (N_16686,N_13975,N_12777);
nand U16687 (N_16687,N_14091,N_12944);
nor U16688 (N_16688,N_14615,N_12731);
nand U16689 (N_16689,N_13285,N_13660);
or U16690 (N_16690,N_14846,N_14762);
nand U16691 (N_16691,N_13416,N_12627);
nand U16692 (N_16692,N_13730,N_14089);
nand U16693 (N_16693,N_14949,N_14538);
nand U16694 (N_16694,N_13727,N_14667);
nor U16695 (N_16695,N_14020,N_14719);
nor U16696 (N_16696,N_14808,N_12738);
or U16697 (N_16697,N_14347,N_14821);
nand U16698 (N_16698,N_14712,N_14874);
nor U16699 (N_16699,N_13763,N_12822);
xnor U16700 (N_16700,N_13232,N_13623);
nand U16701 (N_16701,N_12903,N_13761);
nand U16702 (N_16702,N_12873,N_13937);
or U16703 (N_16703,N_14246,N_13930);
or U16704 (N_16704,N_13586,N_14833);
or U16705 (N_16705,N_14149,N_13821);
or U16706 (N_16706,N_12799,N_12686);
and U16707 (N_16707,N_13607,N_12561);
or U16708 (N_16708,N_12689,N_13732);
or U16709 (N_16709,N_12889,N_12800);
nand U16710 (N_16710,N_14578,N_12802);
nand U16711 (N_16711,N_14876,N_14312);
and U16712 (N_16712,N_13755,N_14562);
nand U16713 (N_16713,N_13303,N_14716);
or U16714 (N_16714,N_13430,N_12979);
xnor U16715 (N_16715,N_13084,N_14722);
nor U16716 (N_16716,N_14755,N_14743);
nor U16717 (N_16717,N_13335,N_13828);
nand U16718 (N_16718,N_14934,N_12642);
nor U16719 (N_16719,N_12591,N_12795);
nor U16720 (N_16720,N_13757,N_12878);
nor U16721 (N_16721,N_14586,N_14555);
nor U16722 (N_16722,N_13488,N_14418);
and U16723 (N_16723,N_13344,N_14933);
nand U16724 (N_16724,N_13623,N_13626);
and U16725 (N_16725,N_12584,N_13293);
and U16726 (N_16726,N_13785,N_14329);
or U16727 (N_16727,N_14152,N_13335);
xor U16728 (N_16728,N_14142,N_12987);
or U16729 (N_16729,N_13853,N_14026);
or U16730 (N_16730,N_13187,N_14793);
xnor U16731 (N_16731,N_13324,N_14882);
nand U16732 (N_16732,N_14963,N_14642);
or U16733 (N_16733,N_13510,N_13727);
nand U16734 (N_16734,N_12554,N_13861);
or U16735 (N_16735,N_14215,N_14768);
xnor U16736 (N_16736,N_13959,N_14672);
nand U16737 (N_16737,N_14224,N_14192);
and U16738 (N_16738,N_14497,N_14441);
and U16739 (N_16739,N_13128,N_12651);
or U16740 (N_16740,N_13675,N_14606);
nand U16741 (N_16741,N_13342,N_14160);
xor U16742 (N_16742,N_14137,N_13662);
nand U16743 (N_16743,N_14044,N_14865);
or U16744 (N_16744,N_13524,N_12557);
nand U16745 (N_16745,N_14541,N_13895);
and U16746 (N_16746,N_14454,N_12586);
nand U16747 (N_16747,N_13832,N_14245);
nand U16748 (N_16748,N_13736,N_13927);
nor U16749 (N_16749,N_14802,N_13433);
nor U16750 (N_16750,N_14544,N_13481);
and U16751 (N_16751,N_13877,N_13443);
or U16752 (N_16752,N_14986,N_13664);
nand U16753 (N_16753,N_13325,N_13984);
or U16754 (N_16754,N_14465,N_13499);
xor U16755 (N_16755,N_14341,N_13177);
nor U16756 (N_16756,N_12962,N_14035);
nand U16757 (N_16757,N_13033,N_14451);
xnor U16758 (N_16758,N_13551,N_14102);
or U16759 (N_16759,N_12953,N_13820);
xor U16760 (N_16760,N_13327,N_13883);
nor U16761 (N_16761,N_14013,N_14315);
nand U16762 (N_16762,N_14963,N_14928);
and U16763 (N_16763,N_12963,N_14840);
xor U16764 (N_16764,N_14925,N_13236);
and U16765 (N_16765,N_12529,N_14628);
nor U16766 (N_16766,N_13539,N_13856);
nor U16767 (N_16767,N_12994,N_13296);
and U16768 (N_16768,N_13283,N_14792);
or U16769 (N_16769,N_13363,N_14239);
nand U16770 (N_16770,N_13098,N_14465);
nand U16771 (N_16771,N_14638,N_14340);
xor U16772 (N_16772,N_14644,N_12819);
nand U16773 (N_16773,N_14303,N_13366);
and U16774 (N_16774,N_13914,N_13454);
and U16775 (N_16775,N_12553,N_14285);
and U16776 (N_16776,N_13637,N_13275);
and U16777 (N_16777,N_14333,N_13845);
xnor U16778 (N_16778,N_13295,N_13887);
nor U16779 (N_16779,N_12651,N_14249);
nor U16780 (N_16780,N_14857,N_13360);
nor U16781 (N_16781,N_12953,N_14432);
nor U16782 (N_16782,N_14931,N_12868);
nand U16783 (N_16783,N_14316,N_12523);
or U16784 (N_16784,N_14108,N_13718);
and U16785 (N_16785,N_12853,N_14679);
or U16786 (N_16786,N_13151,N_14727);
and U16787 (N_16787,N_13109,N_14518);
nand U16788 (N_16788,N_14235,N_13920);
nand U16789 (N_16789,N_14945,N_13792);
nand U16790 (N_16790,N_13970,N_14238);
nor U16791 (N_16791,N_14613,N_14887);
and U16792 (N_16792,N_13909,N_14677);
nand U16793 (N_16793,N_14264,N_14437);
nor U16794 (N_16794,N_14643,N_13488);
and U16795 (N_16795,N_14830,N_12722);
nor U16796 (N_16796,N_12738,N_12610);
nand U16797 (N_16797,N_12609,N_14525);
and U16798 (N_16798,N_13322,N_14283);
nand U16799 (N_16799,N_14650,N_14142);
and U16800 (N_16800,N_14743,N_13312);
nand U16801 (N_16801,N_14398,N_14925);
nor U16802 (N_16802,N_13011,N_13736);
or U16803 (N_16803,N_14561,N_12907);
or U16804 (N_16804,N_13389,N_13633);
nor U16805 (N_16805,N_12704,N_14428);
xnor U16806 (N_16806,N_12883,N_14962);
or U16807 (N_16807,N_13577,N_13379);
or U16808 (N_16808,N_14995,N_13811);
or U16809 (N_16809,N_12523,N_14639);
nor U16810 (N_16810,N_14674,N_12704);
nand U16811 (N_16811,N_13733,N_12509);
or U16812 (N_16812,N_12940,N_14886);
xor U16813 (N_16813,N_12611,N_13732);
xnor U16814 (N_16814,N_12896,N_12624);
or U16815 (N_16815,N_13846,N_13734);
and U16816 (N_16816,N_13892,N_13968);
nor U16817 (N_16817,N_12596,N_14314);
nor U16818 (N_16818,N_14105,N_13009);
xnor U16819 (N_16819,N_13965,N_14738);
and U16820 (N_16820,N_13003,N_14956);
nor U16821 (N_16821,N_14319,N_14569);
or U16822 (N_16822,N_14201,N_14199);
nand U16823 (N_16823,N_13844,N_14632);
or U16824 (N_16824,N_14072,N_14618);
nand U16825 (N_16825,N_14615,N_12638);
or U16826 (N_16826,N_14759,N_13905);
and U16827 (N_16827,N_14880,N_13589);
xor U16828 (N_16828,N_13540,N_14083);
nor U16829 (N_16829,N_13792,N_14664);
or U16830 (N_16830,N_14896,N_12943);
nor U16831 (N_16831,N_13127,N_12695);
nor U16832 (N_16832,N_13432,N_14367);
or U16833 (N_16833,N_14121,N_14670);
or U16834 (N_16834,N_14330,N_13141);
xor U16835 (N_16835,N_14441,N_13872);
nand U16836 (N_16836,N_12985,N_13603);
or U16837 (N_16837,N_14916,N_14633);
and U16838 (N_16838,N_12924,N_13217);
nor U16839 (N_16839,N_14010,N_14142);
xor U16840 (N_16840,N_13798,N_14910);
and U16841 (N_16841,N_13004,N_13523);
or U16842 (N_16842,N_13188,N_14100);
and U16843 (N_16843,N_14274,N_14316);
and U16844 (N_16844,N_14424,N_14313);
nand U16845 (N_16845,N_13754,N_13312);
nand U16846 (N_16846,N_14086,N_13819);
nand U16847 (N_16847,N_12528,N_12865);
nand U16848 (N_16848,N_14690,N_12682);
nand U16849 (N_16849,N_12554,N_14645);
or U16850 (N_16850,N_13447,N_13314);
or U16851 (N_16851,N_13783,N_14999);
nor U16852 (N_16852,N_12615,N_14736);
nor U16853 (N_16853,N_12565,N_12518);
nor U16854 (N_16854,N_12652,N_14124);
or U16855 (N_16855,N_14216,N_14455);
xnor U16856 (N_16856,N_14251,N_12581);
or U16857 (N_16857,N_14870,N_13359);
and U16858 (N_16858,N_12648,N_14857);
and U16859 (N_16859,N_12631,N_12860);
or U16860 (N_16860,N_14416,N_13374);
and U16861 (N_16861,N_14784,N_14404);
and U16862 (N_16862,N_14481,N_13051);
and U16863 (N_16863,N_13669,N_13967);
and U16864 (N_16864,N_14784,N_14631);
nand U16865 (N_16865,N_12605,N_13174);
or U16866 (N_16866,N_14744,N_13940);
nor U16867 (N_16867,N_14666,N_13160);
xnor U16868 (N_16868,N_14167,N_12543);
nor U16869 (N_16869,N_13059,N_13072);
or U16870 (N_16870,N_14373,N_12574);
or U16871 (N_16871,N_13233,N_12640);
and U16872 (N_16872,N_14478,N_13345);
or U16873 (N_16873,N_13467,N_13201);
and U16874 (N_16874,N_14849,N_13948);
nor U16875 (N_16875,N_14795,N_12863);
nand U16876 (N_16876,N_14360,N_13329);
or U16877 (N_16877,N_14339,N_13307);
and U16878 (N_16878,N_12954,N_14454);
nand U16879 (N_16879,N_14840,N_14764);
and U16880 (N_16880,N_13193,N_14352);
or U16881 (N_16881,N_13733,N_13421);
nand U16882 (N_16882,N_14703,N_13893);
or U16883 (N_16883,N_14946,N_13138);
and U16884 (N_16884,N_12947,N_13980);
and U16885 (N_16885,N_12680,N_13889);
and U16886 (N_16886,N_13423,N_12964);
nand U16887 (N_16887,N_14341,N_13911);
nand U16888 (N_16888,N_13168,N_14728);
and U16889 (N_16889,N_13202,N_13398);
nand U16890 (N_16890,N_14092,N_12635);
nand U16891 (N_16891,N_12793,N_13667);
and U16892 (N_16892,N_14306,N_14628);
or U16893 (N_16893,N_13074,N_14778);
or U16894 (N_16894,N_13039,N_13353);
nor U16895 (N_16895,N_13306,N_13266);
nor U16896 (N_16896,N_14951,N_13996);
xnor U16897 (N_16897,N_13236,N_13970);
nand U16898 (N_16898,N_14544,N_14871);
and U16899 (N_16899,N_14801,N_13836);
xnor U16900 (N_16900,N_13564,N_14319);
or U16901 (N_16901,N_14349,N_14772);
nor U16902 (N_16902,N_13518,N_13494);
and U16903 (N_16903,N_14920,N_14176);
and U16904 (N_16904,N_13880,N_12556);
nand U16905 (N_16905,N_13676,N_14032);
nor U16906 (N_16906,N_12856,N_14245);
or U16907 (N_16907,N_14567,N_14570);
nand U16908 (N_16908,N_13079,N_14085);
nand U16909 (N_16909,N_14411,N_13787);
and U16910 (N_16910,N_13784,N_13674);
nor U16911 (N_16911,N_13606,N_13646);
or U16912 (N_16912,N_13952,N_13728);
nand U16913 (N_16913,N_14427,N_12813);
nor U16914 (N_16914,N_12627,N_14030);
nor U16915 (N_16915,N_14339,N_13015);
xnor U16916 (N_16916,N_13084,N_12816);
or U16917 (N_16917,N_13930,N_12994);
nor U16918 (N_16918,N_13098,N_12985);
xor U16919 (N_16919,N_14999,N_13897);
or U16920 (N_16920,N_14337,N_14703);
or U16921 (N_16921,N_13584,N_12945);
nor U16922 (N_16922,N_14229,N_14891);
nand U16923 (N_16923,N_14831,N_14002);
or U16924 (N_16924,N_12940,N_13129);
or U16925 (N_16925,N_14920,N_13917);
and U16926 (N_16926,N_14755,N_12653);
nor U16927 (N_16927,N_14581,N_14157);
nand U16928 (N_16928,N_13193,N_12872);
or U16929 (N_16929,N_13987,N_13650);
nor U16930 (N_16930,N_14286,N_14641);
and U16931 (N_16931,N_14866,N_14560);
nor U16932 (N_16932,N_14700,N_14718);
nand U16933 (N_16933,N_14946,N_12864);
and U16934 (N_16934,N_13382,N_13004);
xor U16935 (N_16935,N_12549,N_13995);
and U16936 (N_16936,N_12544,N_13398);
and U16937 (N_16937,N_13895,N_12592);
nand U16938 (N_16938,N_13193,N_14776);
nor U16939 (N_16939,N_14059,N_14725);
and U16940 (N_16940,N_13986,N_13427);
nand U16941 (N_16941,N_14768,N_14581);
nor U16942 (N_16942,N_13511,N_13036);
xor U16943 (N_16943,N_12793,N_14133);
nand U16944 (N_16944,N_14753,N_13045);
xnor U16945 (N_16945,N_13156,N_14183);
nor U16946 (N_16946,N_14331,N_12870);
and U16947 (N_16947,N_12559,N_14521);
or U16948 (N_16948,N_12550,N_14369);
nand U16949 (N_16949,N_14046,N_13202);
nand U16950 (N_16950,N_14592,N_14412);
nor U16951 (N_16951,N_12619,N_13670);
xor U16952 (N_16952,N_13320,N_13177);
or U16953 (N_16953,N_13452,N_13940);
or U16954 (N_16954,N_13138,N_13003);
nand U16955 (N_16955,N_13357,N_13969);
nand U16956 (N_16956,N_14096,N_13172);
nand U16957 (N_16957,N_13392,N_13295);
nor U16958 (N_16958,N_14027,N_14190);
and U16959 (N_16959,N_14756,N_13755);
nand U16960 (N_16960,N_14985,N_12544);
and U16961 (N_16961,N_14452,N_13218);
nand U16962 (N_16962,N_13036,N_13801);
nand U16963 (N_16963,N_14331,N_13785);
or U16964 (N_16964,N_14522,N_14932);
nor U16965 (N_16965,N_13347,N_12928);
and U16966 (N_16966,N_14305,N_13144);
nand U16967 (N_16967,N_14919,N_13692);
xnor U16968 (N_16968,N_13507,N_14668);
and U16969 (N_16969,N_14075,N_13277);
and U16970 (N_16970,N_13650,N_14020);
nand U16971 (N_16971,N_13618,N_12877);
nand U16972 (N_16972,N_12969,N_13886);
nand U16973 (N_16973,N_14250,N_14844);
nor U16974 (N_16974,N_13941,N_13013);
nand U16975 (N_16975,N_12794,N_14048);
nand U16976 (N_16976,N_13684,N_12876);
or U16977 (N_16977,N_12540,N_13273);
nor U16978 (N_16978,N_12675,N_13707);
or U16979 (N_16979,N_13396,N_13406);
xor U16980 (N_16980,N_13772,N_13320);
nand U16981 (N_16981,N_14072,N_14445);
or U16982 (N_16982,N_12768,N_12601);
or U16983 (N_16983,N_14295,N_14838);
nor U16984 (N_16984,N_14613,N_13753);
or U16985 (N_16985,N_14579,N_13647);
or U16986 (N_16986,N_14117,N_14669);
nand U16987 (N_16987,N_12561,N_14716);
and U16988 (N_16988,N_13815,N_13780);
and U16989 (N_16989,N_13870,N_14394);
and U16990 (N_16990,N_14552,N_12867);
or U16991 (N_16991,N_13333,N_13882);
and U16992 (N_16992,N_12505,N_13861);
or U16993 (N_16993,N_13602,N_13999);
nand U16994 (N_16994,N_14159,N_13228);
nand U16995 (N_16995,N_13240,N_13635);
xor U16996 (N_16996,N_12817,N_13601);
nand U16997 (N_16997,N_14327,N_14714);
and U16998 (N_16998,N_12853,N_13010);
nor U16999 (N_16999,N_13473,N_14742);
or U17000 (N_17000,N_14806,N_13614);
nor U17001 (N_17001,N_12740,N_12793);
or U17002 (N_17002,N_13340,N_13869);
xnor U17003 (N_17003,N_12898,N_12950);
nor U17004 (N_17004,N_12913,N_14899);
nand U17005 (N_17005,N_14230,N_14362);
nand U17006 (N_17006,N_13516,N_13453);
nor U17007 (N_17007,N_13524,N_12984);
and U17008 (N_17008,N_13948,N_14720);
nand U17009 (N_17009,N_14502,N_14765);
and U17010 (N_17010,N_14823,N_14889);
nor U17011 (N_17011,N_14503,N_12886);
or U17012 (N_17012,N_14154,N_13671);
xnor U17013 (N_17013,N_13745,N_12676);
or U17014 (N_17014,N_14897,N_13201);
nor U17015 (N_17015,N_12743,N_14336);
and U17016 (N_17016,N_12769,N_13941);
and U17017 (N_17017,N_13483,N_13869);
and U17018 (N_17018,N_14728,N_12965);
and U17019 (N_17019,N_12847,N_12549);
and U17020 (N_17020,N_14726,N_13742);
nor U17021 (N_17021,N_14294,N_13031);
or U17022 (N_17022,N_12546,N_14539);
nand U17023 (N_17023,N_13722,N_12599);
and U17024 (N_17024,N_14426,N_12948);
nor U17025 (N_17025,N_14639,N_14196);
nand U17026 (N_17026,N_13634,N_13675);
or U17027 (N_17027,N_14432,N_12949);
nor U17028 (N_17028,N_14548,N_13907);
and U17029 (N_17029,N_13516,N_13398);
nand U17030 (N_17030,N_13415,N_14294);
and U17031 (N_17031,N_13504,N_13165);
or U17032 (N_17032,N_14710,N_14482);
nand U17033 (N_17033,N_14094,N_14731);
nor U17034 (N_17034,N_12869,N_13519);
or U17035 (N_17035,N_13275,N_14789);
nand U17036 (N_17036,N_14273,N_12763);
and U17037 (N_17037,N_13133,N_14080);
nor U17038 (N_17038,N_12722,N_14090);
or U17039 (N_17039,N_13638,N_14373);
xnor U17040 (N_17040,N_12563,N_13592);
nor U17041 (N_17041,N_14857,N_13265);
nor U17042 (N_17042,N_12894,N_13929);
and U17043 (N_17043,N_14174,N_12750);
or U17044 (N_17044,N_12682,N_13783);
or U17045 (N_17045,N_13188,N_12530);
nor U17046 (N_17046,N_13288,N_14606);
or U17047 (N_17047,N_14961,N_14916);
nor U17048 (N_17048,N_13548,N_14568);
and U17049 (N_17049,N_12961,N_13855);
and U17050 (N_17050,N_13094,N_14193);
nor U17051 (N_17051,N_14065,N_14048);
or U17052 (N_17052,N_13522,N_13725);
nor U17053 (N_17053,N_13355,N_14415);
and U17054 (N_17054,N_12853,N_14327);
nor U17055 (N_17055,N_14668,N_14868);
and U17056 (N_17056,N_14985,N_13210);
nand U17057 (N_17057,N_14860,N_12892);
or U17058 (N_17058,N_13789,N_13302);
and U17059 (N_17059,N_13079,N_13395);
nor U17060 (N_17060,N_12668,N_14004);
nor U17061 (N_17061,N_14932,N_12897);
nand U17062 (N_17062,N_14407,N_14632);
or U17063 (N_17063,N_13912,N_13900);
nand U17064 (N_17064,N_13246,N_14359);
or U17065 (N_17065,N_13505,N_14329);
or U17066 (N_17066,N_13620,N_13242);
nor U17067 (N_17067,N_14830,N_12513);
nor U17068 (N_17068,N_12617,N_13158);
nand U17069 (N_17069,N_14995,N_14468);
and U17070 (N_17070,N_13932,N_13671);
nor U17071 (N_17071,N_14005,N_14674);
nor U17072 (N_17072,N_12725,N_13236);
and U17073 (N_17073,N_14055,N_13295);
xor U17074 (N_17074,N_14738,N_13305);
nand U17075 (N_17075,N_13682,N_12982);
nor U17076 (N_17076,N_12820,N_13445);
nor U17077 (N_17077,N_13018,N_14223);
nor U17078 (N_17078,N_13266,N_13719);
and U17079 (N_17079,N_13352,N_13713);
or U17080 (N_17080,N_13174,N_13914);
nand U17081 (N_17081,N_14500,N_13517);
nor U17082 (N_17082,N_13371,N_14492);
nand U17083 (N_17083,N_14412,N_14642);
and U17084 (N_17084,N_13244,N_14279);
and U17085 (N_17085,N_14749,N_13872);
and U17086 (N_17086,N_12824,N_13160);
and U17087 (N_17087,N_12950,N_14287);
or U17088 (N_17088,N_14568,N_14272);
or U17089 (N_17089,N_13175,N_14843);
or U17090 (N_17090,N_14172,N_14782);
nor U17091 (N_17091,N_14460,N_14389);
nor U17092 (N_17092,N_13433,N_14559);
or U17093 (N_17093,N_13841,N_14330);
and U17094 (N_17094,N_14021,N_14907);
nor U17095 (N_17095,N_13781,N_12796);
and U17096 (N_17096,N_12561,N_14901);
and U17097 (N_17097,N_14906,N_13907);
nand U17098 (N_17098,N_12509,N_14177);
nor U17099 (N_17099,N_13514,N_13803);
nand U17100 (N_17100,N_13383,N_14715);
or U17101 (N_17101,N_14162,N_13915);
nand U17102 (N_17102,N_14967,N_14563);
or U17103 (N_17103,N_14097,N_14159);
nor U17104 (N_17104,N_13327,N_13561);
and U17105 (N_17105,N_13216,N_13680);
or U17106 (N_17106,N_14198,N_14664);
nand U17107 (N_17107,N_14594,N_14944);
nand U17108 (N_17108,N_12902,N_14069);
and U17109 (N_17109,N_12863,N_14585);
and U17110 (N_17110,N_14021,N_14633);
and U17111 (N_17111,N_12652,N_14430);
nor U17112 (N_17112,N_13021,N_14212);
or U17113 (N_17113,N_14635,N_13230);
and U17114 (N_17114,N_12697,N_12579);
and U17115 (N_17115,N_12707,N_12731);
and U17116 (N_17116,N_14839,N_12815);
xnor U17117 (N_17117,N_12927,N_13708);
nand U17118 (N_17118,N_13583,N_14559);
nand U17119 (N_17119,N_14878,N_13307);
or U17120 (N_17120,N_14671,N_14203);
or U17121 (N_17121,N_14265,N_13826);
or U17122 (N_17122,N_13148,N_14513);
or U17123 (N_17123,N_13714,N_13718);
nand U17124 (N_17124,N_14489,N_14492);
and U17125 (N_17125,N_13607,N_13936);
nor U17126 (N_17126,N_14447,N_14928);
nor U17127 (N_17127,N_13531,N_14687);
and U17128 (N_17128,N_13896,N_13989);
nor U17129 (N_17129,N_12646,N_14079);
nand U17130 (N_17130,N_13859,N_14552);
and U17131 (N_17131,N_14644,N_14902);
and U17132 (N_17132,N_12762,N_14064);
and U17133 (N_17133,N_14130,N_14572);
nor U17134 (N_17134,N_12935,N_12991);
nor U17135 (N_17135,N_14552,N_13569);
and U17136 (N_17136,N_14432,N_13061);
and U17137 (N_17137,N_14419,N_13418);
or U17138 (N_17138,N_13268,N_13542);
or U17139 (N_17139,N_13261,N_14643);
nor U17140 (N_17140,N_13426,N_12871);
and U17141 (N_17141,N_12830,N_14581);
or U17142 (N_17142,N_12666,N_13856);
or U17143 (N_17143,N_13036,N_12750);
nor U17144 (N_17144,N_14033,N_14254);
and U17145 (N_17145,N_13448,N_14633);
xor U17146 (N_17146,N_13258,N_12789);
nor U17147 (N_17147,N_12828,N_13837);
nand U17148 (N_17148,N_13594,N_14376);
nand U17149 (N_17149,N_13313,N_14954);
nor U17150 (N_17150,N_14025,N_14515);
nor U17151 (N_17151,N_14875,N_14213);
nor U17152 (N_17152,N_13072,N_12774);
and U17153 (N_17153,N_14482,N_14601);
nand U17154 (N_17154,N_13192,N_14641);
and U17155 (N_17155,N_12590,N_14296);
or U17156 (N_17156,N_12575,N_14300);
nand U17157 (N_17157,N_14911,N_14741);
or U17158 (N_17158,N_12929,N_14721);
nor U17159 (N_17159,N_14988,N_14721);
nor U17160 (N_17160,N_13302,N_13165);
and U17161 (N_17161,N_13205,N_12906);
nor U17162 (N_17162,N_13153,N_13248);
or U17163 (N_17163,N_14644,N_13990);
nand U17164 (N_17164,N_14955,N_13048);
nand U17165 (N_17165,N_14407,N_12610);
nand U17166 (N_17166,N_14300,N_13722);
nor U17167 (N_17167,N_12781,N_13372);
and U17168 (N_17168,N_13837,N_14200);
xor U17169 (N_17169,N_13616,N_14678);
nor U17170 (N_17170,N_13113,N_12869);
nand U17171 (N_17171,N_12848,N_14183);
and U17172 (N_17172,N_12568,N_13123);
nor U17173 (N_17173,N_14298,N_12740);
xor U17174 (N_17174,N_12600,N_13108);
nand U17175 (N_17175,N_14357,N_13640);
and U17176 (N_17176,N_14392,N_14300);
nand U17177 (N_17177,N_14017,N_12596);
nand U17178 (N_17178,N_14108,N_14419);
or U17179 (N_17179,N_13384,N_13495);
and U17180 (N_17180,N_14032,N_12985);
nand U17181 (N_17181,N_14065,N_13854);
nand U17182 (N_17182,N_14847,N_12752);
and U17183 (N_17183,N_13107,N_12685);
or U17184 (N_17184,N_14177,N_13437);
and U17185 (N_17185,N_13431,N_14197);
and U17186 (N_17186,N_14547,N_14305);
or U17187 (N_17187,N_14066,N_13238);
nand U17188 (N_17188,N_14878,N_12933);
or U17189 (N_17189,N_12935,N_13972);
xnor U17190 (N_17190,N_13431,N_14385);
and U17191 (N_17191,N_13014,N_12831);
nor U17192 (N_17192,N_14091,N_14839);
or U17193 (N_17193,N_13336,N_14874);
xnor U17194 (N_17194,N_13411,N_14291);
nor U17195 (N_17195,N_13466,N_14888);
nor U17196 (N_17196,N_13208,N_14920);
nor U17197 (N_17197,N_14448,N_14523);
nor U17198 (N_17198,N_14038,N_14377);
or U17199 (N_17199,N_14748,N_13343);
or U17200 (N_17200,N_14470,N_12890);
nand U17201 (N_17201,N_14877,N_13322);
or U17202 (N_17202,N_13037,N_12794);
nand U17203 (N_17203,N_12805,N_14386);
xor U17204 (N_17204,N_14173,N_14825);
nor U17205 (N_17205,N_14060,N_14251);
nor U17206 (N_17206,N_13202,N_12796);
nor U17207 (N_17207,N_14021,N_14128);
and U17208 (N_17208,N_14822,N_13936);
nand U17209 (N_17209,N_13148,N_13677);
nor U17210 (N_17210,N_14107,N_13359);
nor U17211 (N_17211,N_14689,N_13117);
nor U17212 (N_17212,N_12909,N_14274);
or U17213 (N_17213,N_14656,N_14464);
nand U17214 (N_17214,N_13780,N_14978);
or U17215 (N_17215,N_12598,N_14098);
nand U17216 (N_17216,N_14725,N_13479);
nor U17217 (N_17217,N_13226,N_13051);
or U17218 (N_17218,N_13328,N_14933);
or U17219 (N_17219,N_14016,N_14110);
xor U17220 (N_17220,N_12859,N_12614);
xnor U17221 (N_17221,N_13361,N_14706);
and U17222 (N_17222,N_12732,N_13406);
or U17223 (N_17223,N_14853,N_12659);
nand U17224 (N_17224,N_12643,N_14018);
and U17225 (N_17225,N_13434,N_12775);
or U17226 (N_17226,N_14919,N_14503);
nor U17227 (N_17227,N_13270,N_12607);
nor U17228 (N_17228,N_14057,N_13958);
nor U17229 (N_17229,N_14863,N_13931);
or U17230 (N_17230,N_13906,N_13839);
nand U17231 (N_17231,N_13431,N_12751);
nor U17232 (N_17232,N_14035,N_13544);
or U17233 (N_17233,N_12940,N_12756);
or U17234 (N_17234,N_12953,N_14589);
nand U17235 (N_17235,N_13284,N_13112);
nand U17236 (N_17236,N_13020,N_14763);
xor U17237 (N_17237,N_12611,N_13785);
or U17238 (N_17238,N_12519,N_13331);
or U17239 (N_17239,N_14276,N_14253);
nand U17240 (N_17240,N_12833,N_13826);
nor U17241 (N_17241,N_13197,N_12686);
and U17242 (N_17242,N_12516,N_14819);
nand U17243 (N_17243,N_14394,N_13666);
nor U17244 (N_17244,N_14290,N_13413);
nor U17245 (N_17245,N_12701,N_14805);
xnor U17246 (N_17246,N_14881,N_13916);
xor U17247 (N_17247,N_14994,N_13513);
xnor U17248 (N_17248,N_13729,N_14179);
and U17249 (N_17249,N_12804,N_14626);
or U17250 (N_17250,N_12607,N_14866);
and U17251 (N_17251,N_14851,N_14314);
nand U17252 (N_17252,N_12637,N_13409);
and U17253 (N_17253,N_13595,N_14735);
and U17254 (N_17254,N_13310,N_14713);
nor U17255 (N_17255,N_13629,N_12747);
or U17256 (N_17256,N_14398,N_14910);
xor U17257 (N_17257,N_13400,N_13040);
nand U17258 (N_17258,N_12688,N_13503);
nor U17259 (N_17259,N_14839,N_12961);
nor U17260 (N_17260,N_14114,N_13849);
and U17261 (N_17261,N_14465,N_14919);
nand U17262 (N_17262,N_14783,N_14947);
nor U17263 (N_17263,N_13192,N_14098);
and U17264 (N_17264,N_13519,N_14153);
nand U17265 (N_17265,N_14259,N_14673);
nand U17266 (N_17266,N_12793,N_14021);
nand U17267 (N_17267,N_13541,N_14197);
and U17268 (N_17268,N_12758,N_13589);
nand U17269 (N_17269,N_14161,N_13734);
or U17270 (N_17270,N_14014,N_12677);
nand U17271 (N_17271,N_12609,N_14617);
nand U17272 (N_17272,N_13938,N_13812);
nand U17273 (N_17273,N_14388,N_12573);
or U17274 (N_17274,N_13961,N_14313);
and U17275 (N_17275,N_13294,N_14751);
nor U17276 (N_17276,N_13144,N_12875);
xor U17277 (N_17277,N_13966,N_13835);
nand U17278 (N_17278,N_13599,N_12785);
or U17279 (N_17279,N_13144,N_13073);
nand U17280 (N_17280,N_13082,N_14445);
and U17281 (N_17281,N_13676,N_13566);
nand U17282 (N_17282,N_14584,N_14526);
and U17283 (N_17283,N_12889,N_12731);
xor U17284 (N_17284,N_13362,N_12717);
or U17285 (N_17285,N_12770,N_12824);
nor U17286 (N_17286,N_14365,N_14944);
nor U17287 (N_17287,N_13822,N_14358);
or U17288 (N_17288,N_14378,N_14895);
or U17289 (N_17289,N_12580,N_14906);
or U17290 (N_17290,N_12703,N_13419);
nand U17291 (N_17291,N_14820,N_12851);
and U17292 (N_17292,N_12595,N_14868);
nand U17293 (N_17293,N_13317,N_14941);
nor U17294 (N_17294,N_12524,N_13480);
nand U17295 (N_17295,N_13220,N_14488);
or U17296 (N_17296,N_12873,N_12508);
nand U17297 (N_17297,N_14671,N_12982);
or U17298 (N_17298,N_13485,N_14966);
nand U17299 (N_17299,N_13068,N_13763);
xor U17300 (N_17300,N_12641,N_13540);
or U17301 (N_17301,N_13790,N_13878);
nand U17302 (N_17302,N_14500,N_14529);
nand U17303 (N_17303,N_12558,N_13699);
and U17304 (N_17304,N_13347,N_13594);
nand U17305 (N_17305,N_14475,N_14577);
xor U17306 (N_17306,N_12956,N_14362);
and U17307 (N_17307,N_13156,N_14081);
nand U17308 (N_17308,N_13911,N_13502);
nor U17309 (N_17309,N_12765,N_13405);
or U17310 (N_17310,N_13721,N_14202);
nor U17311 (N_17311,N_14961,N_13569);
nor U17312 (N_17312,N_14088,N_13035);
nand U17313 (N_17313,N_13195,N_14729);
or U17314 (N_17314,N_12696,N_13422);
and U17315 (N_17315,N_12638,N_14746);
and U17316 (N_17316,N_12766,N_12654);
and U17317 (N_17317,N_13499,N_13171);
nor U17318 (N_17318,N_14620,N_12642);
nand U17319 (N_17319,N_14168,N_13074);
and U17320 (N_17320,N_13670,N_13091);
or U17321 (N_17321,N_13830,N_13378);
nand U17322 (N_17322,N_12742,N_13549);
or U17323 (N_17323,N_13825,N_12688);
or U17324 (N_17324,N_13281,N_14169);
and U17325 (N_17325,N_14129,N_12834);
and U17326 (N_17326,N_14436,N_13632);
or U17327 (N_17327,N_13782,N_14165);
or U17328 (N_17328,N_13904,N_13672);
nor U17329 (N_17329,N_13176,N_14904);
or U17330 (N_17330,N_14474,N_14389);
and U17331 (N_17331,N_12678,N_13148);
or U17332 (N_17332,N_14044,N_12773);
nand U17333 (N_17333,N_13800,N_14461);
nand U17334 (N_17334,N_14978,N_13271);
and U17335 (N_17335,N_14464,N_12935);
nand U17336 (N_17336,N_14748,N_14030);
nand U17337 (N_17337,N_13602,N_13726);
and U17338 (N_17338,N_13584,N_13127);
nor U17339 (N_17339,N_14812,N_14537);
nor U17340 (N_17340,N_13689,N_14079);
or U17341 (N_17341,N_12986,N_14283);
or U17342 (N_17342,N_13571,N_14250);
or U17343 (N_17343,N_14449,N_13660);
and U17344 (N_17344,N_14837,N_14145);
nand U17345 (N_17345,N_14729,N_13303);
nor U17346 (N_17346,N_13304,N_14657);
nand U17347 (N_17347,N_13472,N_13912);
nor U17348 (N_17348,N_12921,N_14515);
nor U17349 (N_17349,N_14962,N_14286);
or U17350 (N_17350,N_12748,N_13914);
nand U17351 (N_17351,N_13765,N_14625);
nand U17352 (N_17352,N_14128,N_12882);
or U17353 (N_17353,N_14044,N_14803);
nor U17354 (N_17354,N_13772,N_14585);
nor U17355 (N_17355,N_14610,N_14666);
xnor U17356 (N_17356,N_13002,N_12503);
nand U17357 (N_17357,N_14526,N_13699);
nand U17358 (N_17358,N_13070,N_13728);
and U17359 (N_17359,N_13383,N_14611);
nor U17360 (N_17360,N_14340,N_12795);
nand U17361 (N_17361,N_14046,N_13909);
or U17362 (N_17362,N_12622,N_12844);
and U17363 (N_17363,N_13804,N_13642);
or U17364 (N_17364,N_14433,N_14140);
or U17365 (N_17365,N_13656,N_13615);
nor U17366 (N_17366,N_14714,N_13515);
nand U17367 (N_17367,N_14437,N_13849);
nand U17368 (N_17368,N_13597,N_14260);
or U17369 (N_17369,N_13887,N_14390);
nand U17370 (N_17370,N_13678,N_13002);
nor U17371 (N_17371,N_14405,N_12682);
nand U17372 (N_17372,N_13199,N_14224);
or U17373 (N_17373,N_12691,N_13759);
nand U17374 (N_17374,N_14196,N_13106);
or U17375 (N_17375,N_14312,N_13262);
or U17376 (N_17376,N_13236,N_13825);
or U17377 (N_17377,N_14741,N_13739);
or U17378 (N_17378,N_14572,N_13733);
and U17379 (N_17379,N_13248,N_13839);
and U17380 (N_17380,N_13167,N_12714);
and U17381 (N_17381,N_13042,N_13864);
and U17382 (N_17382,N_14196,N_14505);
xnor U17383 (N_17383,N_13650,N_12942);
or U17384 (N_17384,N_13135,N_14994);
nor U17385 (N_17385,N_14404,N_13407);
nand U17386 (N_17386,N_14574,N_12523);
or U17387 (N_17387,N_12657,N_13682);
or U17388 (N_17388,N_14705,N_14832);
or U17389 (N_17389,N_14978,N_14073);
and U17390 (N_17390,N_14697,N_14628);
and U17391 (N_17391,N_13857,N_14615);
or U17392 (N_17392,N_13732,N_13351);
or U17393 (N_17393,N_13601,N_14113);
xor U17394 (N_17394,N_12872,N_12674);
nand U17395 (N_17395,N_12764,N_14443);
xnor U17396 (N_17396,N_12708,N_13073);
and U17397 (N_17397,N_13978,N_13615);
nor U17398 (N_17398,N_14312,N_13328);
nand U17399 (N_17399,N_13502,N_14689);
nor U17400 (N_17400,N_14207,N_12969);
and U17401 (N_17401,N_14116,N_13126);
and U17402 (N_17402,N_14339,N_14481);
and U17403 (N_17403,N_13187,N_13329);
nand U17404 (N_17404,N_12764,N_13374);
and U17405 (N_17405,N_12706,N_12951);
nand U17406 (N_17406,N_12636,N_14056);
nand U17407 (N_17407,N_13048,N_14520);
nand U17408 (N_17408,N_14828,N_13806);
nor U17409 (N_17409,N_13237,N_13769);
nand U17410 (N_17410,N_13249,N_12829);
or U17411 (N_17411,N_13850,N_13853);
or U17412 (N_17412,N_14476,N_14624);
and U17413 (N_17413,N_14363,N_12573);
and U17414 (N_17414,N_13549,N_14676);
and U17415 (N_17415,N_13202,N_14649);
nor U17416 (N_17416,N_14365,N_14818);
nand U17417 (N_17417,N_14849,N_14039);
nor U17418 (N_17418,N_14538,N_13013);
nand U17419 (N_17419,N_12860,N_12787);
xnor U17420 (N_17420,N_14548,N_13826);
and U17421 (N_17421,N_13463,N_13488);
xnor U17422 (N_17422,N_12840,N_13537);
nand U17423 (N_17423,N_14309,N_12550);
xnor U17424 (N_17424,N_13450,N_12574);
or U17425 (N_17425,N_14983,N_12705);
and U17426 (N_17426,N_13245,N_13176);
or U17427 (N_17427,N_12856,N_12775);
or U17428 (N_17428,N_13933,N_13584);
nand U17429 (N_17429,N_13288,N_13033);
nand U17430 (N_17430,N_13001,N_12953);
or U17431 (N_17431,N_13481,N_12676);
or U17432 (N_17432,N_12888,N_13733);
or U17433 (N_17433,N_12525,N_13077);
xor U17434 (N_17434,N_14486,N_14762);
and U17435 (N_17435,N_13509,N_14212);
and U17436 (N_17436,N_14120,N_13187);
nand U17437 (N_17437,N_13971,N_13036);
and U17438 (N_17438,N_13360,N_13336);
xor U17439 (N_17439,N_14446,N_13712);
nand U17440 (N_17440,N_14007,N_13811);
nand U17441 (N_17441,N_13846,N_14698);
nor U17442 (N_17442,N_14197,N_13922);
nand U17443 (N_17443,N_13151,N_12823);
nand U17444 (N_17444,N_13938,N_13901);
or U17445 (N_17445,N_14391,N_13837);
nor U17446 (N_17446,N_14483,N_12954);
nor U17447 (N_17447,N_14721,N_14747);
xor U17448 (N_17448,N_13531,N_14408);
nand U17449 (N_17449,N_13644,N_13841);
xor U17450 (N_17450,N_13537,N_14381);
or U17451 (N_17451,N_14161,N_13866);
nor U17452 (N_17452,N_13215,N_14421);
nand U17453 (N_17453,N_13233,N_13903);
xnor U17454 (N_17454,N_12663,N_13309);
or U17455 (N_17455,N_14336,N_14665);
or U17456 (N_17456,N_14484,N_13811);
xnor U17457 (N_17457,N_12832,N_13267);
nand U17458 (N_17458,N_13485,N_13436);
nor U17459 (N_17459,N_14493,N_14277);
nand U17460 (N_17460,N_12958,N_13047);
or U17461 (N_17461,N_13873,N_13799);
nand U17462 (N_17462,N_13681,N_13288);
nand U17463 (N_17463,N_13016,N_14426);
nor U17464 (N_17464,N_12740,N_13373);
and U17465 (N_17465,N_14587,N_14535);
nor U17466 (N_17466,N_13711,N_12866);
nor U17467 (N_17467,N_13786,N_13678);
or U17468 (N_17468,N_12550,N_13993);
or U17469 (N_17469,N_14104,N_14727);
or U17470 (N_17470,N_13824,N_14405);
nor U17471 (N_17471,N_13776,N_13933);
and U17472 (N_17472,N_14108,N_14770);
nor U17473 (N_17473,N_12788,N_12932);
or U17474 (N_17474,N_13589,N_13327);
nand U17475 (N_17475,N_14904,N_14581);
nand U17476 (N_17476,N_14550,N_14299);
nor U17477 (N_17477,N_14672,N_13446);
nor U17478 (N_17478,N_14412,N_14409);
and U17479 (N_17479,N_12566,N_12851);
or U17480 (N_17480,N_14984,N_14284);
nor U17481 (N_17481,N_13637,N_13076);
nor U17482 (N_17482,N_14559,N_13158);
and U17483 (N_17483,N_14751,N_12878);
or U17484 (N_17484,N_13391,N_14690);
nor U17485 (N_17485,N_14957,N_13107);
or U17486 (N_17486,N_13121,N_13565);
and U17487 (N_17487,N_13481,N_14753);
xnor U17488 (N_17488,N_13681,N_14781);
or U17489 (N_17489,N_14682,N_13991);
nor U17490 (N_17490,N_14247,N_14114);
nor U17491 (N_17491,N_13412,N_14298);
and U17492 (N_17492,N_12586,N_14239);
xnor U17493 (N_17493,N_13733,N_13767);
nor U17494 (N_17494,N_14641,N_14156);
nand U17495 (N_17495,N_13070,N_12531);
nand U17496 (N_17496,N_13288,N_12741);
nor U17497 (N_17497,N_13358,N_12896);
xnor U17498 (N_17498,N_12713,N_12930);
or U17499 (N_17499,N_14213,N_13771);
nor U17500 (N_17500,N_16872,N_16441);
and U17501 (N_17501,N_16213,N_16518);
and U17502 (N_17502,N_16774,N_16795);
nand U17503 (N_17503,N_15869,N_16664);
nor U17504 (N_17504,N_17254,N_15318);
and U17505 (N_17505,N_17132,N_15621);
or U17506 (N_17506,N_16968,N_16477);
or U17507 (N_17507,N_16417,N_17090);
and U17508 (N_17508,N_17215,N_17048);
or U17509 (N_17509,N_17034,N_15913);
nor U17510 (N_17510,N_15376,N_15779);
xor U17511 (N_17511,N_17310,N_15684);
nor U17512 (N_17512,N_16648,N_16360);
nand U17513 (N_17513,N_16473,N_15940);
or U17514 (N_17514,N_15328,N_16025);
or U17515 (N_17515,N_15240,N_17062);
nor U17516 (N_17516,N_15487,N_17042);
nand U17517 (N_17517,N_15829,N_17299);
and U17518 (N_17518,N_17138,N_17358);
or U17519 (N_17519,N_16099,N_17346);
or U17520 (N_17520,N_16359,N_16547);
nor U17521 (N_17521,N_16143,N_15601);
and U17522 (N_17522,N_17009,N_17490);
and U17523 (N_17523,N_16301,N_16969);
and U17524 (N_17524,N_16005,N_17499);
and U17525 (N_17525,N_15321,N_16493);
nor U17526 (N_17526,N_15781,N_15868);
nand U17527 (N_17527,N_16031,N_16341);
nand U17528 (N_17528,N_15517,N_15374);
or U17529 (N_17529,N_15973,N_16408);
or U17530 (N_17530,N_15138,N_16410);
and U17531 (N_17531,N_15160,N_17244);
nor U17532 (N_17532,N_16890,N_15100);
nand U17533 (N_17533,N_15447,N_16576);
and U17534 (N_17534,N_15945,N_16788);
nor U17535 (N_17535,N_15439,N_15468);
xnor U17536 (N_17536,N_17051,N_16353);
xnor U17537 (N_17537,N_17201,N_16762);
xor U17538 (N_17538,N_15928,N_15052);
xnor U17539 (N_17539,N_17454,N_16511);
nand U17540 (N_17540,N_16034,N_16431);
or U17541 (N_17541,N_15588,N_15354);
or U17542 (N_17542,N_15101,N_17091);
nor U17543 (N_17543,N_17283,N_15802);
or U17544 (N_17544,N_16864,N_16930);
or U17545 (N_17545,N_17344,N_17230);
nor U17546 (N_17546,N_15436,N_16804);
and U17547 (N_17547,N_16538,N_16685);
or U17548 (N_17548,N_15429,N_16910);
nor U17549 (N_17549,N_16394,N_15576);
nor U17550 (N_17550,N_16237,N_15417);
or U17551 (N_17551,N_16815,N_17243);
and U17552 (N_17552,N_16085,N_17417);
xnor U17553 (N_17553,N_16616,N_16227);
nor U17554 (N_17554,N_17455,N_16054);
nor U17555 (N_17555,N_17181,N_16636);
nor U17556 (N_17556,N_15622,N_17222);
and U17557 (N_17557,N_15933,N_15078);
or U17558 (N_17558,N_16841,N_16110);
nor U17559 (N_17559,N_16332,N_16934);
nand U17560 (N_17560,N_15999,N_15244);
nand U17561 (N_17561,N_16634,N_16751);
or U17562 (N_17562,N_16033,N_15366);
nand U17563 (N_17563,N_16418,N_16255);
nor U17564 (N_17564,N_15809,N_17288);
or U17565 (N_17565,N_16909,N_16081);
or U17566 (N_17566,N_15590,N_15368);
nand U17567 (N_17567,N_16138,N_16334);
and U17568 (N_17568,N_16597,N_15414);
nand U17569 (N_17569,N_17427,N_16991);
or U17570 (N_17570,N_16502,N_17405);
or U17571 (N_17571,N_17095,N_16853);
nand U17572 (N_17572,N_16615,N_15213);
and U17573 (N_17573,N_15125,N_17452);
and U17574 (N_17574,N_17493,N_16783);
and U17575 (N_17575,N_17311,N_15126);
nand U17576 (N_17576,N_15864,N_16567);
nand U17577 (N_17577,N_15330,N_16194);
nor U17578 (N_17578,N_15128,N_15316);
nor U17579 (N_17579,N_16624,N_16595);
nor U17580 (N_17580,N_15730,N_17206);
nor U17581 (N_17581,N_17149,N_16283);
nand U17582 (N_17582,N_16737,N_16637);
nand U17583 (N_17583,N_15412,N_15259);
or U17584 (N_17584,N_16541,N_16537);
and U17585 (N_17585,N_16376,N_16197);
or U17586 (N_17586,N_17073,N_16221);
and U17587 (N_17587,N_16328,N_15946);
and U17588 (N_17588,N_15390,N_17225);
nor U17589 (N_17589,N_15109,N_17497);
or U17590 (N_17590,N_16368,N_15494);
and U17591 (N_17591,N_16661,N_17218);
or U17592 (N_17592,N_16736,N_16520);
nor U17593 (N_17593,N_17361,N_15168);
or U17594 (N_17594,N_15117,N_16643);
and U17595 (N_17595,N_15932,N_15996);
or U17596 (N_17596,N_15431,N_15993);
nor U17597 (N_17597,N_16561,N_17207);
nor U17598 (N_17598,N_15580,N_15790);
and U17599 (N_17599,N_15971,N_16438);
nand U17600 (N_17600,N_15575,N_17433);
nor U17601 (N_17601,N_15907,N_16193);
nand U17602 (N_17602,N_17019,N_15824);
or U17603 (N_17603,N_15253,N_15617);
and U17604 (N_17604,N_15740,N_16100);
nor U17605 (N_17605,N_15513,N_16126);
nand U17606 (N_17606,N_15013,N_16101);
nor U17607 (N_17607,N_17468,N_16210);
and U17608 (N_17608,N_17307,N_16793);
or U17609 (N_17609,N_17135,N_15484);
nand U17610 (N_17610,N_16173,N_15036);
or U17611 (N_17611,N_16524,N_15333);
nand U17612 (N_17612,N_17457,N_15844);
nand U17613 (N_17613,N_17354,N_16055);
nor U17614 (N_17614,N_17316,N_15323);
xnor U17615 (N_17615,N_15975,N_16988);
nor U17616 (N_17616,N_17128,N_16510);
xor U17617 (N_17617,N_16144,N_15122);
or U17618 (N_17618,N_16844,N_15169);
or U17619 (N_17619,N_15678,N_16282);
xnor U17620 (N_17620,N_15827,N_15055);
and U17621 (N_17621,N_17148,N_16906);
nor U17622 (N_17622,N_15093,N_16926);
nor U17623 (N_17623,N_16933,N_16794);
xnor U17624 (N_17624,N_16164,N_16504);
or U17625 (N_17625,N_15605,N_16366);
and U17626 (N_17626,N_15363,N_16010);
xor U17627 (N_17627,N_16722,N_15107);
nor U17628 (N_17628,N_15948,N_15839);
and U17629 (N_17629,N_16008,N_16580);
or U17630 (N_17630,N_15015,N_15005);
nor U17631 (N_17631,N_17485,N_16363);
nor U17632 (N_17632,N_17265,N_16843);
nand U17633 (N_17633,N_16551,N_15609);
and U17634 (N_17634,N_16225,N_15927);
or U17635 (N_17635,N_16188,N_16084);
nor U17636 (N_17636,N_17349,N_16784);
nand U17637 (N_17637,N_15378,N_16350);
nor U17638 (N_17638,N_16591,N_15749);
nand U17639 (N_17639,N_15774,N_16396);
or U17640 (N_17640,N_17018,N_15269);
and U17641 (N_17641,N_16730,N_15962);
and U17642 (N_17642,N_16923,N_16782);
or U17643 (N_17643,N_15862,N_16501);
or U17644 (N_17644,N_15921,N_16187);
and U17645 (N_17645,N_15179,N_16049);
nor U17646 (N_17646,N_17247,N_15771);
and U17647 (N_17647,N_16155,N_16542);
or U17648 (N_17648,N_15021,N_17453);
nand U17649 (N_17649,N_15966,N_15937);
nand U17650 (N_17650,N_15514,N_15049);
or U17651 (N_17651,N_15947,N_15950);
nand U17652 (N_17652,N_17210,N_15400);
nor U17653 (N_17653,N_17328,N_16007);
nand U17654 (N_17654,N_17326,N_16831);
nor U17655 (N_17655,N_15235,N_17136);
nor U17656 (N_17656,N_17327,N_17082);
or U17657 (N_17657,N_15581,N_16190);
and U17658 (N_17658,N_16594,N_17476);
or U17659 (N_17659,N_16308,N_15832);
nand U17660 (N_17660,N_15067,N_16092);
and U17661 (N_17661,N_16397,N_15938);
or U17662 (N_17662,N_15242,N_15681);
or U17663 (N_17663,N_17382,N_15196);
nand U17664 (N_17664,N_17366,N_15880);
nor U17665 (N_17665,N_16826,N_17268);
and U17666 (N_17666,N_17140,N_15442);
nor U17667 (N_17667,N_15770,N_15645);
xnor U17668 (N_17668,N_16306,N_15184);
or U17669 (N_17669,N_16663,N_15619);
and U17670 (N_17670,N_16873,N_15964);
nor U17671 (N_17671,N_15625,N_17087);
nand U17672 (N_17672,N_16427,N_16768);
or U17673 (N_17673,N_15134,N_15452);
or U17674 (N_17674,N_15450,N_16797);
nor U17675 (N_17675,N_15828,N_15025);
and U17676 (N_17676,N_15696,N_16810);
nand U17677 (N_17677,N_15387,N_16822);
xnor U17678 (N_17678,N_16146,N_17432);
nand U17679 (N_17679,N_16902,N_15592);
nand U17680 (N_17680,N_17280,N_16086);
nand U17681 (N_17681,N_17383,N_15340);
and U17682 (N_17682,N_16461,N_15761);
nand U17683 (N_17683,N_15531,N_15367);
nand U17684 (N_17684,N_16691,N_16936);
nand U17685 (N_17685,N_15427,N_15438);
and U17686 (N_17686,N_17246,N_17281);
nor U17687 (N_17687,N_15399,N_17159);
nor U17688 (N_17688,N_15075,N_16728);
nor U17689 (N_17689,N_17269,N_15532);
and U17690 (N_17690,N_16167,N_17055);
or U17691 (N_17691,N_16488,N_15448);
nor U17692 (N_17692,N_17237,N_16045);
or U17693 (N_17693,N_16199,N_15509);
or U17694 (N_17694,N_16435,N_15744);
nand U17695 (N_17695,N_16956,N_15370);
nand U17696 (N_17696,N_15922,N_16851);
xor U17697 (N_17697,N_16162,N_17263);
or U17698 (N_17698,N_16627,N_16953);
or U17699 (N_17699,N_15338,N_15606);
xnor U17700 (N_17700,N_15108,N_16203);
nand U17701 (N_17701,N_16927,N_16932);
nand U17702 (N_17702,N_15292,N_15879);
and U17703 (N_17703,N_15251,N_16985);
and U17704 (N_17704,N_17040,N_17340);
and U17705 (N_17705,N_15456,N_16620);
xor U17706 (N_17706,N_15845,N_16997);
and U17707 (N_17707,N_17496,N_15663);
nor U17708 (N_17708,N_17459,N_15132);
nor U17709 (N_17709,N_16121,N_15463);
xor U17710 (N_17710,N_16258,N_15857);
nor U17711 (N_17711,N_15270,N_16151);
and U17712 (N_17712,N_17267,N_16606);
nor U17713 (N_17713,N_15926,N_16354);
or U17714 (N_17714,N_17076,N_16867);
or U17715 (N_17715,N_17302,N_15389);
and U17716 (N_17716,N_17146,N_15265);
nor U17717 (N_17717,N_17155,N_15916);
or U17718 (N_17718,N_15293,N_16669);
nor U17719 (N_17719,N_16564,N_15028);
and U17720 (N_17720,N_15904,N_15079);
nand U17721 (N_17721,N_15657,N_17294);
nor U17722 (N_17722,N_17185,N_15643);
nor U17723 (N_17723,N_16814,N_16087);
and U17724 (N_17724,N_17190,N_15212);
nand U17725 (N_17725,N_15104,N_15523);
or U17726 (N_17726,N_17421,N_17020);
and U17727 (N_17727,N_16449,N_16463);
or U17728 (N_17728,N_15551,N_17204);
nor U17729 (N_17729,N_16130,N_16954);
nor U17730 (N_17730,N_16068,N_15068);
and U17731 (N_17731,N_16484,N_16280);
nand U17732 (N_17732,N_16714,N_15310);
nor U17733 (N_17733,N_16242,N_16471);
nand U17734 (N_17734,N_16119,N_17111);
nand U17735 (N_17735,N_17022,N_17184);
and U17736 (N_17736,N_15788,N_15812);
nor U17737 (N_17737,N_17122,N_16051);
nor U17738 (N_17738,N_16073,N_16671);
and U17739 (N_17739,N_15754,N_16016);
and U17740 (N_17740,N_16917,N_16738);
nand U17741 (N_17741,N_16950,N_15566);
nor U17742 (N_17742,N_15713,N_16267);
nor U17743 (N_17743,N_15291,N_15026);
xnor U17744 (N_17744,N_15508,N_15209);
or U17745 (N_17745,N_15140,N_17012);
nor U17746 (N_17746,N_17050,N_15193);
or U17747 (N_17747,N_15453,N_17304);
or U17748 (N_17748,N_15748,N_15525);
nor U17749 (N_17749,N_16293,N_15519);
nor U17750 (N_17750,N_16743,N_15976);
and U17751 (N_17751,N_15673,N_15407);
and U17752 (N_17752,N_17063,N_15180);
or U17753 (N_17753,N_16223,N_16381);
and U17754 (N_17754,N_15563,N_15538);
nand U17755 (N_17755,N_16881,N_16569);
nand U17756 (N_17756,N_16063,N_16649);
and U17757 (N_17757,N_17115,N_16772);
xnor U17758 (N_17758,N_17420,N_16106);
and U17759 (N_17759,N_16982,N_15102);
nor U17760 (N_17760,N_16529,N_15614);
or U17761 (N_17761,N_15556,N_16082);
or U17762 (N_17762,N_16224,N_16204);
nor U17763 (N_17763,N_15382,N_16820);
and U17764 (N_17764,N_15313,N_16388);
nand U17765 (N_17765,N_15098,N_17364);
xnor U17766 (N_17766,N_15432,N_15320);
or U17767 (N_17767,N_16114,N_16995);
xnor U17768 (N_17768,N_17345,N_15472);
nor U17769 (N_17769,N_15446,N_15041);
xnor U17770 (N_17770,N_17378,N_15986);
and U17771 (N_17771,N_16840,N_15396);
or U17772 (N_17772,N_16407,N_16905);
nor U17773 (N_17773,N_15097,N_17440);
xor U17774 (N_17774,N_15796,N_16159);
and U17775 (N_17775,N_17166,N_16787);
or U17776 (N_17776,N_15115,N_16708);
or U17777 (N_17777,N_15943,N_16064);
nand U17778 (N_17778,N_16048,N_15949);
nand U17779 (N_17779,N_15148,N_17449);
or U17780 (N_17780,N_15324,N_16458);
nor U17781 (N_17781,N_16827,N_15279);
or U17782 (N_17782,N_15658,N_17229);
nand U17783 (N_17783,N_15358,N_15655);
nand U17784 (N_17784,N_15383,N_15243);
or U17785 (N_17785,N_15751,N_16614);
nor U17786 (N_17786,N_17429,N_16182);
nor U17787 (N_17787,N_16260,N_16653);
and U17788 (N_17788,N_17387,N_17072);
nand U17789 (N_17789,N_16076,N_16185);
and U17790 (N_17790,N_17100,N_15155);
nand U17791 (N_17791,N_16414,N_15939);
nor U17792 (N_17792,N_16939,N_16123);
and U17793 (N_17793,N_15651,N_15159);
and U17794 (N_17794,N_17235,N_16248);
and U17795 (N_17795,N_15351,N_17406);
and U17796 (N_17796,N_16043,N_17093);
xnor U17797 (N_17797,N_17415,N_15511);
or U17798 (N_17798,N_15489,N_15598);
and U17799 (N_17799,N_15664,N_15051);
or U17800 (N_17800,N_16865,N_17151);
and U17801 (N_17801,N_15612,N_15860);
nand U17802 (N_17802,N_15290,N_17197);
nand U17803 (N_17803,N_15995,N_16657);
nand U17804 (N_17804,N_15226,N_16713);
and U17805 (N_17805,N_15967,N_15162);
or U17806 (N_17806,N_16131,N_16503);
nor U17807 (N_17807,N_15755,N_15863);
or U17808 (N_17808,N_15236,N_17052);
or U17809 (N_17809,N_15706,N_16771);
and U17810 (N_17810,N_17092,N_17029);
or U17811 (N_17811,N_16442,N_16701);
and U17812 (N_17812,N_15165,N_16240);
and U17813 (N_17813,N_17451,N_16948);
or U17814 (N_17814,N_16535,N_15170);
nor U17815 (N_17815,N_16451,N_16333);
or U17816 (N_17816,N_15894,N_15053);
nand U17817 (N_17817,N_16599,N_17306);
and U17818 (N_17818,N_16120,N_16852);
xnor U17819 (N_17819,N_17450,N_15114);
and U17820 (N_17820,N_16113,N_16269);
or U17821 (N_17821,N_16666,N_15349);
xnor U17822 (N_17822,N_17372,N_17202);
nor U17823 (N_17823,N_15952,N_15561);
or U17824 (N_17824,N_16147,N_17279);
nor U17825 (N_17825,N_17318,N_15500);
or U17826 (N_17826,N_15173,N_16554);
or U17827 (N_17827,N_15018,N_16566);
and U17828 (N_17828,N_16891,N_16592);
nand U17829 (N_17829,N_16758,N_17370);
or U17830 (N_17830,N_16300,N_17213);
nand U17831 (N_17831,N_15183,N_16989);
or U17832 (N_17832,N_15840,N_15794);
nand U17833 (N_17833,N_17043,N_17084);
nand U17834 (N_17834,N_15559,N_15283);
nor U17835 (N_17835,N_15589,N_15359);
or U17836 (N_17836,N_16655,N_17110);
nor U17837 (N_17837,N_16393,N_15615);
and U17838 (N_17838,N_17038,N_17160);
nor U17839 (N_17839,N_15958,N_15301);
nor U17840 (N_17840,N_16205,N_16125);
and U17841 (N_17841,N_15604,N_15662);
nand U17842 (N_17842,N_17396,N_15174);
or U17843 (N_17843,N_16707,N_15888);
or U17844 (N_17844,N_15882,N_17097);
or U17845 (N_17845,N_15300,N_16790);
or U17846 (N_17846,N_15111,N_17030);
nand U17847 (N_17847,N_16103,N_16543);
nor U17848 (N_17848,N_15153,N_16999);
and U17849 (N_17849,N_15762,N_17338);
or U17850 (N_17850,N_16078,N_16605);
nor U17851 (N_17851,N_16344,N_16466);
nor U17852 (N_17852,N_17231,N_16975);
nand U17853 (N_17853,N_16860,N_17272);
nor U17854 (N_17854,N_15195,N_15764);
nand U17855 (N_17855,N_16578,N_16295);
xnor U17856 (N_17856,N_15070,N_16009);
nand U17857 (N_17857,N_16839,N_15640);
nor U17858 (N_17858,N_15203,N_16492);
or U17859 (N_17859,N_15821,N_16035);
nand U17860 (N_17860,N_15488,N_17023);
or U17861 (N_17861,N_16482,N_16108);
or U17862 (N_17862,N_16745,N_15144);
nand U17863 (N_17863,N_15022,N_15903);
nor U17864 (N_17864,N_16791,N_15527);
nor U17865 (N_17865,N_16302,N_15066);
or U17866 (N_17866,N_17033,N_15006);
or U17867 (N_17867,N_17350,N_16095);
and U17868 (N_17868,N_16725,N_16265);
nand U17869 (N_17869,N_17170,N_15677);
nand U17870 (N_17870,N_15746,N_15000);
and U17871 (N_17871,N_16483,N_16059);
and U17872 (N_17872,N_17035,N_15482);
or U17873 (N_17873,N_16253,N_15951);
and U17874 (N_17874,N_16195,N_16135);
nand U17875 (N_17875,N_15676,N_16370);
nor U17876 (N_17876,N_16490,N_15276);
xnor U17877 (N_17877,N_17445,N_16623);
or U17878 (N_17878,N_16311,N_17203);
nor U17879 (N_17879,N_17362,N_15397);
nor U17880 (N_17880,N_16673,N_16986);
or U17881 (N_17881,N_15573,N_15200);
nand U17882 (N_17882,N_17343,N_17162);
and U17883 (N_17883,N_16047,N_15024);
nor U17884 (N_17884,N_16962,N_16878);
nor U17885 (N_17885,N_17465,N_16142);
nor U17886 (N_17886,N_15116,N_15987);
nand U17887 (N_17887,N_15685,N_16153);
nor U17888 (N_17888,N_15766,N_17386);
nand U17889 (N_17889,N_15145,N_15364);
or U17890 (N_17890,N_16924,N_16337);
nor U17891 (N_17891,N_16343,N_15080);
or U17892 (N_17892,N_16717,N_16403);
and U17893 (N_17893,N_15418,N_16735);
nor U17894 (N_17894,N_15475,N_16645);
and U17895 (N_17895,N_15957,N_17105);
nand U17896 (N_17896,N_15668,N_15027);
and U17897 (N_17897,N_15247,N_16012);
nand U17898 (N_17898,N_16964,N_16882);
nand U17899 (N_17899,N_16491,N_15653);
nor U17900 (N_17900,N_16992,N_16709);
or U17901 (N_17901,N_16452,N_16298);
xor U17902 (N_17902,N_15884,N_17291);
and U17903 (N_17903,N_15011,N_17355);
or U17904 (N_17904,N_15734,N_17320);
nor U17905 (N_17905,N_17284,N_15600);
and U17906 (N_17906,N_16895,N_16896);
xor U17907 (N_17907,N_16176,N_16780);
xnor U17908 (N_17908,N_17003,N_15808);
xnor U17909 (N_17909,N_15239,N_15050);
nor U17910 (N_17910,N_15570,N_16854);
xnor U17911 (N_17911,N_16915,N_15188);
and U17912 (N_17912,N_15325,N_15158);
nor U17913 (N_17913,N_17456,N_16998);
xor U17914 (N_17914,N_16877,N_15620);
nor U17915 (N_17915,N_15039,N_16026);
nand U17916 (N_17916,N_15076,N_16601);
or U17917 (N_17917,N_15002,N_16373);
nor U17918 (N_17918,N_16675,N_16575);
nor U17919 (N_17919,N_16274,N_17436);
nand U17920 (N_17920,N_15392,N_16152);
nor U17921 (N_17921,N_16404,N_15786);
nor U17922 (N_17922,N_16979,N_16446);
and U17923 (N_17923,N_16022,N_16468);
or U17924 (N_17924,N_17224,N_15874);
xor U17925 (N_17925,N_17194,N_15991);
nand U17926 (N_17926,N_16695,N_15222);
nand U17927 (N_17927,N_15035,N_16355);
and U17928 (N_17928,N_15268,N_17489);
nor U17929 (N_17929,N_16519,N_15234);
xnor U17930 (N_17930,N_16356,N_16874);
xnor U17931 (N_17931,N_16846,N_15020);
xnor U17932 (N_17932,N_15833,N_15595);
or U17933 (N_17933,N_15982,N_16455);
nand U17934 (N_17934,N_17464,N_16568);
and U17935 (N_17935,N_16208,N_15727);
nor U17936 (N_17936,N_15955,N_15217);
or U17937 (N_17937,N_16678,N_15742);
nand U17938 (N_17938,N_17017,N_17319);
nand U17939 (N_17939,N_16244,N_15697);
nand U17940 (N_17940,N_16763,N_15223);
nand U17941 (N_17941,N_17195,N_16424);
or U17942 (N_17942,N_15229,N_16799);
nand U17943 (N_17943,N_15683,N_16157);
nand U17944 (N_17944,N_15872,N_16044);
and U17945 (N_17945,N_15065,N_16074);
and U17946 (N_17946,N_17120,N_16305);
nor U17947 (N_17947,N_15810,N_15799);
xor U17948 (N_17948,N_17067,N_16565);
nor U17949 (N_17949,N_16764,N_15785);
or U17950 (N_17950,N_15717,N_16241);
nand U17951 (N_17951,N_15670,N_17333);
nand U17952 (N_17952,N_15186,N_15635);
nand U17953 (N_17953,N_15486,N_15284);
nand U17954 (N_17954,N_15665,N_16129);
nor U17955 (N_17955,N_16245,N_15281);
nand U17956 (N_17956,N_17479,N_16154);
nand U17957 (N_17957,N_15142,N_16422);
nand U17958 (N_17958,N_16207,N_16700);
xor U17959 (N_17959,N_15637,N_16724);
and U17960 (N_17960,N_17000,N_15403);
xor U17961 (N_17961,N_17086,N_17175);
or U17962 (N_17962,N_16377,N_16230);
nor U17963 (N_17963,N_15225,N_15758);
or U17964 (N_17964,N_17205,N_17080);
nor U17965 (N_17965,N_15547,N_15492);
nand U17966 (N_17966,N_16361,N_15900);
or U17967 (N_17967,N_15731,N_15516);
nand U17968 (N_17968,N_15972,N_17053);
nor U17969 (N_17969,N_15047,N_16105);
or U17970 (N_17970,N_15064,N_16586);
nand U17971 (N_17971,N_17488,N_15315);
and U17972 (N_17972,N_17466,N_16670);
and U17973 (N_17973,N_15485,N_15189);
xor U17974 (N_17974,N_15215,N_15759);
nor U17975 (N_17975,N_16018,N_16749);
nor U17976 (N_17976,N_16444,N_16433);
or U17977 (N_17977,N_16139,N_16065);
or U17978 (N_17978,N_16824,N_15411);
and U17979 (N_17979,N_16229,N_16046);
nand U17980 (N_17980,N_15695,N_17253);
xor U17981 (N_17981,N_15515,N_15019);
or U17982 (N_17982,N_17167,N_17379);
nor U17983 (N_17983,N_15666,N_16517);
nor U17984 (N_17984,N_15769,N_15750);
nor U17985 (N_17985,N_16413,N_17130);
nand U17986 (N_17986,N_16960,N_15917);
and U17987 (N_17987,N_17388,N_17483);
nor U17988 (N_17988,N_17047,N_15433);
xor U17989 (N_17989,N_16888,N_17198);
and U17990 (N_17990,N_16457,N_17257);
or U17991 (N_17991,N_17068,N_15257);
and U17992 (N_17992,N_17347,N_16801);
and U17993 (N_17993,N_16478,N_17404);
or U17994 (N_17994,N_16498,N_16702);
nor U17995 (N_17995,N_15783,N_16385);
or U17996 (N_17996,N_15819,N_15745);
nor U17997 (N_17997,N_15194,N_16371);
xnor U17998 (N_17998,N_16235,N_16056);
nor U17999 (N_17999,N_16037,N_16961);
xor U18000 (N_18000,N_16165,N_17348);
and U18001 (N_18001,N_16515,N_15633);
nand U18002 (N_18002,N_15878,N_16596);
nor U18003 (N_18003,N_16312,N_16994);
or U18004 (N_18004,N_15136,N_16384);
nor U18005 (N_18005,N_16416,N_16289);
nor U18006 (N_18006,N_17081,N_17236);
xnor U18007 (N_18007,N_16178,N_17251);
nor U18008 (N_18008,N_16651,N_15757);
or U18009 (N_18009,N_17153,N_17187);
nand U18010 (N_18010,N_16262,N_17303);
and U18011 (N_18011,N_16970,N_15627);
nor U18012 (N_18012,N_16398,N_15813);
xnor U18013 (N_18013,N_15385,N_17238);
xor U18014 (N_18014,N_16734,N_16352);
or U18015 (N_18015,N_15478,N_15347);
and U18016 (N_18016,N_16522,N_17252);
or U18017 (N_18017,N_17492,N_17367);
and U18018 (N_18018,N_17178,N_17389);
and U18019 (N_18019,N_16617,N_15061);
nand U18020 (N_18020,N_15660,N_16557);
nand U18021 (N_18021,N_16598,N_16689);
xor U18022 (N_18022,N_16358,N_15371);
or U18023 (N_18023,N_16401,N_15255);
or U18024 (N_18024,N_17004,N_17077);
and U18025 (N_18025,N_15739,N_16102);
and U18026 (N_18026,N_17056,N_16476);
and U18027 (N_18027,N_15638,N_15069);
nand U18028 (N_18028,N_17079,N_15649);
or U18029 (N_18029,N_17463,N_17352);
or U18030 (N_18030,N_15038,N_17470);
nor U18031 (N_18031,N_16472,N_15565);
nand U18032 (N_18032,N_15702,N_16607);
or U18033 (N_18033,N_15549,N_16303);
nor U18034 (N_18034,N_15521,N_15369);
and U18035 (N_18035,N_16641,N_15906);
and U18036 (N_18036,N_17308,N_17227);
or U18037 (N_18037,N_16186,N_15554);
or U18038 (N_18038,N_16180,N_17223);
nand U18039 (N_18039,N_16057,N_16856);
or U18040 (N_18040,N_16549,N_15607);
or U18041 (N_18041,N_16629,N_17117);
nor U18042 (N_18042,N_15540,N_15143);
or U18043 (N_18043,N_16279,N_16214);
or U18044 (N_18044,N_15352,N_15406);
or U18045 (N_18045,N_15546,N_15274);
xor U18046 (N_18046,N_15130,N_16117);
and U18047 (N_18047,N_15629,N_15185);
and U18048 (N_18048,N_17498,N_17199);
and U18049 (N_18049,N_16166,N_15709);
or U18050 (N_18050,N_15801,N_16757);
xor U18051 (N_18051,N_15543,N_16818);
or U18052 (N_18052,N_17085,N_17031);
xor U18053 (N_18053,N_17005,N_15218);
nor U18054 (N_18054,N_16775,N_15451);
nand U18055 (N_18055,N_16609,N_15510);
or U18056 (N_18056,N_15208,N_17474);
and U18057 (N_18057,N_15384,N_17221);
and U18058 (N_18058,N_16340,N_17103);
nand U18059 (N_18059,N_16263,N_16247);
nor U18060 (N_18060,N_16278,N_17270);
or U18061 (N_18061,N_15007,N_15254);
nand U18062 (N_18062,N_16965,N_16239);
and U18063 (N_18063,N_15797,N_16281);
xor U18064 (N_18064,N_16218,N_16516);
nor U18065 (N_18065,N_15963,N_17065);
xor U18066 (N_18066,N_17480,N_17032);
and U18067 (N_18067,N_16573,N_16475);
nor U18068 (N_18068,N_16633,N_17484);
nor U18069 (N_18069,N_16487,N_15469);
or U18070 (N_18070,N_17232,N_16816);
nand U18071 (N_18071,N_16765,N_16859);
nor U18072 (N_18072,N_16369,N_16972);
nor U18073 (N_18073,N_16993,N_17002);
nand U18074 (N_18074,N_16200,N_16944);
and U18075 (N_18075,N_16217,N_15777);
nand U18076 (N_18076,N_15644,N_16539);
nand U18077 (N_18077,N_16550,N_16505);
nor U18078 (N_18078,N_15309,N_16329);
and U18079 (N_18079,N_15329,N_17107);
or U18080 (N_18080,N_17475,N_15924);
nor U18081 (N_18081,N_15388,N_16094);
or U18082 (N_18082,N_15715,N_16323);
and U18083 (N_18083,N_15923,N_17013);
or U18084 (N_18084,N_17192,N_15842);
nor U18085 (N_18085,N_17189,N_15176);
and U18086 (N_18086,N_16583,N_16789);
xor U18087 (N_18087,N_15736,N_17098);
or U18088 (N_18088,N_16072,N_15033);
nor U18089 (N_18089,N_15008,N_16706);
or U18090 (N_18090,N_15772,N_15379);
and U18091 (N_18091,N_15214,N_16618);
nand U18092 (N_18092,N_15567,N_15445);
and U18093 (N_18093,N_15425,N_17321);
xor U18094 (N_18094,N_16090,N_15336);
and U18095 (N_18095,N_16336,N_15161);
or U18096 (N_18096,N_16704,N_16644);
or U18097 (N_18097,N_15732,N_17139);
and U18098 (N_18098,N_15703,N_15669);
xor U18099 (N_18099,N_16869,N_16177);
xor U18100 (N_18100,N_15373,N_17133);
and U18101 (N_18101,N_15584,N_16058);
nand U18102 (N_18102,N_16863,N_15848);
or U18103 (N_18103,N_15800,N_15377);
and U18104 (N_18104,N_17447,N_16069);
and U18105 (N_18105,N_16088,N_16286);
or U18106 (N_18106,N_16423,N_15853);
or U18107 (N_18107,N_16409,N_17460);
nor U18108 (N_18108,N_17339,N_16083);
nand U18109 (N_18109,N_15342,N_17437);
or U18110 (N_18110,N_15099,N_17390);
nor U18111 (N_18111,N_16705,N_15082);
nor U18112 (N_18112,N_17300,N_15404);
or U18113 (N_18113,N_15843,N_16897);
and U18114 (N_18114,N_16331,N_17060);
nor U18115 (N_18115,N_16912,N_15671);
or U18116 (N_18116,N_16171,N_17039);
nor U18117 (N_18117,N_15464,N_17430);
nor U18118 (N_18118,N_15712,N_16019);
nand U18119 (N_18119,N_16006,N_16039);
nand U18120 (N_18120,N_16588,N_16243);
xor U18121 (N_18121,N_15231,N_15569);
nand U18122 (N_18122,N_16823,N_17228);
xnor U18123 (N_18123,N_15564,N_16715);
or U18124 (N_18124,N_16145,N_16805);
or U18125 (N_18125,N_17169,N_15199);
nand U18126 (N_18126,N_15124,N_16957);
and U18127 (N_18127,N_15711,N_17255);
or U18128 (N_18128,N_15341,N_15959);
or U18129 (N_18129,N_16903,N_15056);
nor U18130 (N_18130,N_15238,N_16779);
or U18131 (N_18131,N_17070,N_15555);
or U18132 (N_18132,N_16067,N_17371);
or U18133 (N_18133,N_16556,N_15820);
xor U18134 (N_18134,N_16526,N_15123);
and U18135 (N_18135,N_17341,N_15030);
nand U18136 (N_18136,N_16681,N_15046);
nor U18137 (N_18137,N_16904,N_15348);
nor U18138 (N_18138,N_15562,N_15823);
nor U18139 (N_18139,N_16506,N_16434);
and U18140 (N_18140,N_17127,N_17487);
nor U18141 (N_18141,N_17314,N_15550);
nand U18142 (N_18142,N_15944,N_16421);
or U18143 (N_18143,N_15803,N_15545);
nand U18144 (N_18144,N_16955,N_16838);
nand U18145 (N_18145,N_15694,N_16546);
nor U18146 (N_18146,N_16158,N_17274);
and U18147 (N_18147,N_15306,N_15072);
xor U18148 (N_18148,N_17481,N_17219);
or U18149 (N_18149,N_17315,N_15434);
and U18150 (N_18150,N_16315,N_16677);
nor U18151 (N_18151,N_16639,N_16104);
nand U18152 (N_18152,N_15294,N_17006);
xnor U18153 (N_18153,N_15322,N_17446);
and U18154 (N_18154,N_17337,N_16602);
or U18155 (N_18155,N_16600,N_15499);
xnor U18156 (N_18156,N_17241,N_15163);
or U18157 (N_18157,N_17239,N_15577);
and U18158 (N_18158,N_15981,N_16480);
or U18159 (N_18159,N_17412,N_15441);
xor U18160 (N_18160,N_17143,N_16212);
nand U18161 (N_18161,N_15867,N_15381);
and U18162 (N_18162,N_15308,N_15258);
and U18163 (N_18163,N_15205,N_16628);
or U18164 (N_18164,N_16777,N_15262);
and U18165 (N_18165,N_15127,N_15430);
and U18166 (N_18166,N_17164,N_16430);
nand U18167 (N_18167,N_15910,N_16321);
nor U18168 (N_18168,N_15830,N_15260);
nand U18169 (N_18169,N_16942,N_16378);
nand U18170 (N_18170,N_16454,N_15707);
nand U18171 (N_18171,N_16536,N_16949);
nor U18172 (N_18172,N_15652,N_16003);
and U18173 (N_18173,N_15063,N_15299);
or U18174 (N_18174,N_15582,N_17161);
and U18175 (N_18175,N_15303,N_16291);
nor U18176 (N_18176,N_16866,N_16273);
or U18177 (N_18177,N_17240,N_15335);
nand U18178 (N_18178,N_15421,N_15267);
or U18179 (N_18179,N_16211,N_16870);
nand U18180 (N_18180,N_15861,N_15151);
nand U18181 (N_18181,N_15929,N_17419);
and U18182 (N_18182,N_15305,N_17114);
or U18183 (N_18183,N_15768,N_15723);
or U18184 (N_18184,N_16978,N_16662);
or U18185 (N_18185,N_16761,N_15084);
and U18186 (N_18186,N_15150,N_16109);
nand U18187 (N_18187,N_15542,N_16766);
nand U18188 (N_18188,N_15728,N_16920);
and U18189 (N_18189,N_16880,N_16813);
or U18190 (N_18190,N_16357,N_16495);
and U18191 (N_18191,N_16727,N_15426);
nand U18192 (N_18192,N_17322,N_16299);
and U18193 (N_18193,N_15071,N_15206);
or U18194 (N_18194,N_15202,N_15956);
nand U18195 (N_18195,N_17398,N_15719);
nor U18196 (N_18196,N_15775,N_16889);
nor U18197 (N_18197,N_15327,N_16387);
xor U18198 (N_18198,N_15881,N_16935);
or U18199 (N_18199,N_16236,N_17220);
nor U18200 (N_18200,N_15798,N_17037);
nand U18201 (N_18201,N_16445,N_16015);
nor U18202 (N_18202,N_15192,N_15187);
and U18203 (N_18203,N_15031,N_16729);
nor U18204 (N_18204,N_15302,N_16603);
nand U18205 (N_18205,N_16107,N_15455);
nand U18206 (N_18206,N_16496,N_15818);
nand U18207 (N_18207,N_15286,N_16811);
or U18208 (N_18208,N_16938,N_16364);
and U18209 (N_18209,N_15642,N_17234);
or U18210 (N_18210,N_15228,N_16553);
and U18211 (N_18211,N_17331,N_15250);
or U18212 (N_18212,N_15282,N_17407);
nand U18213 (N_18213,N_15297,N_16532);
nor U18214 (N_18214,N_15154,N_15477);
xnor U18215 (N_18215,N_17026,N_15571);
nand U18216 (N_18216,N_17041,N_16079);
or U18217 (N_18217,N_15095,N_16579);
nor U18218 (N_18218,N_15522,N_15659);
or U18219 (N_18219,N_16676,N_16703);
nand U18220 (N_18220,N_17426,N_16029);
and U18221 (N_18221,N_15850,N_15978);
or U18222 (N_18222,N_16389,N_15585);
or U18223 (N_18223,N_16711,N_16175);
and U18224 (N_18224,N_16558,N_17400);
nand U18225 (N_18225,N_17125,N_15763);
or U18226 (N_18226,N_15277,N_16412);
nor U18227 (N_18227,N_17486,N_17101);
or U18228 (N_18228,N_15724,N_17262);
nand U18229 (N_18229,N_15059,N_15897);
nand U18230 (N_18230,N_17045,N_16133);
or U18231 (N_18231,N_16161,N_16342);
and U18232 (N_18232,N_15834,N_16324);
xnor U18233 (N_18233,N_16124,N_16367);
xor U18234 (N_18234,N_15618,N_16460);
and U18235 (N_18235,N_15859,N_16497);
nand U18236 (N_18236,N_17008,N_15435);
or U18237 (N_18237,N_15023,N_15083);
xor U18238 (N_18238,N_15990,N_17357);
nor U18239 (N_18239,N_16066,N_16001);
or U18240 (N_18240,N_17360,N_16581);
nand U18241 (N_18241,N_17021,N_16170);
nor U18242 (N_18242,N_17177,N_15825);
nor U18243 (N_18243,N_16313,N_17168);
or U18244 (N_18244,N_16885,N_16612);
and U18245 (N_18245,N_15139,N_16608);
or U18246 (N_18246,N_17109,N_15647);
or U18247 (N_18247,N_16544,N_16070);
nor U18248 (N_18248,N_16365,N_15146);
or U18249 (N_18249,N_16169,N_17011);
nand U18250 (N_18250,N_16326,N_17373);
and U18251 (N_18251,N_15413,N_16391);
and U18252 (N_18252,N_16876,N_16249);
nor U18253 (N_18253,N_17402,N_16901);
or U18254 (N_18254,N_15743,N_15210);
xnor U18255 (N_18255,N_15483,N_16275);
and U18256 (N_18256,N_15895,N_16692);
nor U18257 (N_18257,N_17188,N_15557);
nand U18258 (N_18258,N_16834,N_16322);
or U18259 (N_18259,N_16201,N_16345);
or U18260 (N_18260,N_16577,N_16115);
nor U18261 (N_18261,N_17152,N_15191);
xnor U18262 (N_18262,N_16660,N_15345);
nand U18263 (N_18263,N_15776,N_15885);
nand U18264 (N_18264,N_17472,N_17027);
and U18265 (N_18265,N_16559,N_15476);
or U18266 (N_18266,N_16786,N_15423);
or U18267 (N_18267,N_15930,N_16020);
nor U18268 (N_18268,N_16481,N_15044);
nand U18269 (N_18269,N_16319,N_16191);
and U18270 (N_18270,N_17410,N_16908);
nand U18271 (N_18271,N_17448,N_15893);
and U18272 (N_18272,N_16428,N_17106);
nand U18273 (N_18273,N_16952,N_15220);
and U18274 (N_18274,N_17108,N_17064);
nand U18275 (N_18275,N_16741,N_16990);
or U18276 (N_18276,N_15503,N_16832);
nand U18277 (N_18277,N_15314,N_15062);
or U18278 (N_18278,N_16694,N_15171);
nor U18279 (N_18279,N_16499,N_16122);
and U18280 (N_18280,N_17173,N_15437);
nand U18281 (N_18281,N_17129,N_17066);
nor U18282 (N_18282,N_15524,N_16089);
nor U18283 (N_18283,N_16971,N_15232);
and U18284 (N_18284,N_15471,N_15273);
nand U18285 (N_18285,N_16233,N_17495);
or U18286 (N_18286,N_16593,N_15714);
nand U18287 (N_18287,N_17259,N_17381);
or U18288 (N_18288,N_17428,N_17121);
nand U18289 (N_18289,N_15536,N_15735);
nand U18290 (N_18290,N_16552,N_16587);
nand U18291 (N_18291,N_17332,N_15221);
nand U18292 (N_18292,N_16590,N_15835);
nor U18293 (N_18293,N_16626,N_17317);
nand U18294 (N_18294,N_17282,N_15890);
nor U18295 (N_18295,N_16527,N_16149);
or U18296 (N_18296,N_16759,N_15700);
or U18297 (N_18297,N_15636,N_16437);
nor U18298 (N_18298,N_15245,N_15493);
nor U18299 (N_18299,N_15156,N_15674);
or U18300 (N_18300,N_15831,N_16755);
xor U18301 (N_18301,N_16687,N_16830);
nor U18302 (N_18302,N_15586,N_16307);
or U18303 (N_18303,N_16000,N_17423);
or U18304 (N_18304,N_15460,N_15989);
and U18305 (N_18305,N_17124,N_16156);
or U18306 (N_18306,N_15402,N_16395);
and U18307 (N_18307,N_15918,N_16682);
nand U18308 (N_18308,N_17182,N_16183);
or U18309 (N_18309,N_15889,N_16440);
and U18310 (N_18310,N_16746,N_16405);
or U18311 (N_18311,N_15911,N_15841);
xor U18312 (N_18312,N_16718,N_17059);
or U18313 (N_18313,N_15462,N_15656);
or U18314 (N_18314,N_15805,N_15086);
or U18315 (N_18315,N_15866,N_16148);
nor U18316 (N_18316,N_17256,N_16686);
xor U18317 (N_18317,N_16582,N_17329);
or U18318 (N_18318,N_16925,N_16574);
and U18319 (N_18319,N_16272,N_17094);
xor U18320 (N_18320,N_16011,N_15773);
nor U18321 (N_18321,N_15149,N_16380);
nand U18322 (N_18322,N_16062,N_17351);
and U18323 (N_18323,N_17323,N_16479);
nand U18324 (N_18324,N_16459,N_16375);
nand U18325 (N_18325,N_15587,N_16320);
or U18326 (N_18326,N_16947,N_17297);
xor U18327 (N_18327,N_15256,N_17296);
nand U18328 (N_18328,N_15846,N_17165);
or U18329 (N_18329,N_15870,N_15871);
nand U18330 (N_18330,N_15876,N_16747);
xnor U18331 (N_18331,N_15942,N_16292);
xnor U18332 (N_18332,N_15395,N_16168);
or U18333 (N_18333,N_16919,N_15908);
or U18334 (N_18334,N_16621,N_16837);
or U18335 (N_18335,N_15454,N_16362);
and U18336 (N_18336,N_16238,N_15988);
and U18337 (N_18337,N_15641,N_17112);
nor U18338 (N_18338,N_15498,N_17075);
or U18339 (N_18339,N_15806,N_15909);
and U18340 (N_18340,N_15248,N_17145);
and U18341 (N_18341,N_16346,N_17147);
xor U18342 (N_18342,N_17438,N_15856);
nor U18343 (N_18343,N_15854,N_15380);
and U18344 (N_18344,N_16310,N_16928);
or U18345 (N_18345,N_15602,N_16946);
or U18346 (N_18346,N_15470,N_15747);
and U18347 (N_18347,N_15361,N_15077);
nand U18348 (N_18348,N_16509,N_16382);
nand U18349 (N_18349,N_17007,N_16189);
nor U18350 (N_18350,N_16339,N_16821);
nor U18351 (N_18351,N_15443,N_15705);
or U18352 (N_18352,N_15689,N_15899);
or U18353 (N_18353,N_17482,N_16785);
or U18354 (N_18354,N_16937,N_16271);
nor U18355 (N_18355,N_15416,N_17356);
and U18356 (N_18356,N_15365,N_17458);
nor U18357 (N_18357,N_15449,N_17377);
nand U18358 (N_18358,N_16770,N_16351);
nand U18359 (N_18359,N_15865,N_17209);
nand U18360 (N_18360,N_17200,N_16533);
or U18361 (N_18361,N_17275,N_16017);
or U18362 (N_18362,N_16439,N_17261);
nand U18363 (N_18363,N_16647,N_15716);
nand U18364 (N_18364,N_17416,N_17353);
and U18365 (N_18365,N_15334,N_17399);
or U18366 (N_18366,N_15631,N_15060);
and U18367 (N_18367,N_15693,N_16512);
nand U18368 (N_18368,N_15935,N_15765);
nor U18369 (N_18369,N_15237,N_15816);
or U18370 (N_18370,N_16489,N_17174);
nor U18371 (N_18371,N_15722,N_16053);
or U18372 (N_18372,N_17154,N_16884);
nor U18373 (N_18373,N_15968,N_15954);
and U18374 (N_18374,N_15690,N_15375);
xor U18375 (N_18375,N_15181,N_15394);
or U18376 (N_18376,N_15997,N_15386);
or U18377 (N_18377,N_17271,N_15778);
or U18378 (N_18378,N_16684,N_15211);
nor U18379 (N_18379,N_16809,N_16585);
nor U18380 (N_18380,N_15591,N_16096);
or U18381 (N_18381,N_16383,N_16215);
xor U18382 (N_18382,N_17088,N_15054);
nor U18383 (N_18383,N_15198,N_16467);
and U18384 (N_18384,N_16297,N_15409);
nand U18385 (N_18385,N_15037,N_15961);
nor U18386 (N_18386,N_16918,N_16050);
nor U18387 (N_18387,N_17444,N_15648);
xnor U18388 (N_18388,N_16800,N_16419);
or U18389 (N_18389,N_16773,N_16940);
xnor U18390 (N_18390,N_15898,N_15467);
and U18391 (N_18391,N_16256,N_15410);
or U18392 (N_18392,N_15105,N_16625);
xor U18393 (N_18393,N_16679,N_16808);
nand U18394 (N_18394,N_15568,N_15272);
and U18395 (N_18395,N_15855,N_17313);
nor U18396 (N_18396,N_17494,N_16325);
and U18397 (N_18397,N_17431,N_17290);
xnor U18398 (N_18398,N_15440,N_16374);
nand U18399 (N_18399,N_16447,N_15458);
nand U18400 (N_18400,N_15634,N_15393);
and U18401 (N_18401,N_16807,N_16513);
and U18402 (N_18402,N_17156,N_15172);
or U18403 (N_18403,N_17462,N_16667);
nand U18404 (N_18404,N_15419,N_15616);
nor U18405 (N_18405,N_16665,N_15495);
nand U18406 (N_18406,N_16137,N_16028);
or U18407 (N_18407,N_16753,N_16432);
nor U18408 (N_18408,N_16443,N_17301);
or U18409 (N_18409,N_15147,N_16112);
and U18410 (N_18410,N_16893,N_17425);
nor U18411 (N_18411,N_15398,N_15197);
and U18412 (N_18412,N_15275,N_17216);
nand U18413 (N_18413,N_17123,N_15480);
nor U18414 (N_18414,N_16696,N_15886);
and U18415 (N_18415,N_16967,N_16631);
and U18416 (N_18416,N_16849,N_15701);
nand U18417 (N_18417,N_16042,N_16220);
or U18418 (N_18418,N_17439,N_17158);
and U18419 (N_18419,N_15583,N_15473);
and U18420 (N_18420,N_16128,N_16030);
nor U18421 (N_18421,N_15915,N_15001);
nor U18422 (N_18422,N_17211,N_17309);
xnor U18423 (N_18423,N_15137,N_15630);
nand U18424 (N_18424,N_15356,N_16710);
xor U18425 (N_18425,N_15767,N_15353);
nor U18426 (N_18426,N_16338,N_15307);
and U18427 (N_18427,N_16179,N_16562);
and U18428 (N_18428,N_16638,N_15698);
nand U18429 (N_18429,N_15496,N_15331);
or U18430 (N_18430,N_15103,N_16690);
or U18431 (N_18431,N_15849,N_17054);
or U18432 (N_18432,N_15249,N_15029);
nor U18433 (N_18433,N_17150,N_17025);
nand U18434 (N_18434,N_16032,N_16219);
and U18435 (N_18435,N_16683,N_17172);
nor U18436 (N_18436,N_16828,N_17071);
and U18437 (N_18437,N_16425,N_15623);
nor U18438 (N_18438,N_16469,N_15691);
nand U18439 (N_18439,N_15682,N_16958);
or U18440 (N_18440,N_16060,N_15597);
nor U18441 (N_18441,N_16514,N_16379);
nor U18442 (N_18442,N_16977,N_16726);
xnor U18443 (N_18443,N_15057,N_16270);
nor U18444 (N_18444,N_15167,N_15672);
nand U18445 (N_18445,N_17141,N_16610);
or U18446 (N_18446,N_17001,N_16571);
xor U18447 (N_18447,N_16091,N_15710);
xnor U18448 (N_18448,N_15970,N_15479);
and U18449 (N_18449,N_15012,N_17435);
nor U18450 (N_18450,N_16754,N_16732);
xnor U18451 (N_18451,N_15296,N_15408);
or U18452 (N_18452,N_15501,N_15073);
nand U18453 (N_18453,N_16659,N_15733);
nand U18454 (N_18454,N_16750,N_15780);
nand U18455 (N_18455,N_15687,N_15548);
and U18456 (N_18456,N_15692,N_16222);
xnor U18457 (N_18457,N_16817,N_15009);
nand U18458 (N_18458,N_17413,N_15541);
xnor U18459 (N_18459,N_17245,N_15977);
and U18460 (N_18460,N_17342,N_15852);
or U18461 (N_18461,N_15466,N_15784);
nor U18462 (N_18462,N_17046,N_15680);
nand U18463 (N_18463,N_17144,N_16525);
nand U18464 (N_18464,N_17096,N_16951);
xnor U18465 (N_18465,N_15626,N_15791);
nor U18466 (N_18466,N_16531,N_16879);
nor U18467 (N_18467,N_16132,N_16931);
nand U18468 (N_18468,N_15405,N_16760);
nor U18469 (N_18469,N_15085,N_15266);
and U18470 (N_18470,N_15157,N_15688);
or U18471 (N_18471,N_16226,N_16150);
xor U18472 (N_18472,N_15795,N_15216);
or U18473 (N_18473,N_15241,N_16974);
nand U18474 (N_18474,N_16309,N_15883);
nand U18475 (N_18475,N_16752,N_16654);
and U18476 (N_18476,N_16984,N_16652);
or U18477 (N_18477,N_15121,N_15133);
and U18478 (N_18478,N_15782,N_16996);
and U18479 (N_18479,N_17391,N_15088);
nor U18480 (N_18480,N_15985,N_16792);
xnor U18481 (N_18481,N_15994,N_17242);
and U18482 (N_18482,N_16916,N_16680);
nand U18483 (N_18483,N_16184,N_15014);
nand U18484 (N_18484,N_16098,N_16871);
nor U18485 (N_18485,N_17191,N_16898);
nand U18486 (N_18486,N_15807,N_17285);
nand U18487 (N_18487,N_16259,N_17273);
and U18488 (N_18488,N_15787,N_16436);
nand U18489 (N_18489,N_15974,N_15135);
and U18490 (N_18490,N_15016,N_16160);
nor U18491 (N_18491,N_15873,N_15444);
nand U18492 (N_18492,N_16004,N_15112);
or U18493 (N_18493,N_15639,N_16400);
and U18494 (N_18494,N_16163,N_15089);
or U18495 (N_18495,N_15304,N_16181);
nor U18496 (N_18496,N_17365,N_16252);
and U18497 (N_18497,N_16500,N_16257);
or U18498 (N_18498,N_15401,N_15343);
xnor U18499 (N_18499,N_16327,N_17374);
or U18500 (N_18500,N_16894,N_17324);
and U18501 (N_18501,N_17286,N_17264);
nand U18502 (N_18502,N_15457,N_15901);
and U18503 (N_18503,N_15465,N_16448);
nand U18504 (N_18504,N_15896,N_15288);
and U18505 (N_18505,N_15624,N_15979);
nand U18506 (N_18506,N_17102,N_16494);
and U18507 (N_18507,N_15391,N_15737);
nand U18508 (N_18508,N_17214,N_15611);
nand U18509 (N_18509,N_15686,N_17044);
or U18510 (N_18510,N_15699,N_17137);
xnor U18511 (N_18511,N_15350,N_16118);
nand U18512 (N_18512,N_15357,N_15289);
nand U18513 (N_18513,N_17477,N_16330);
nand U18514 (N_18514,N_15969,N_16555);
and U18515 (N_18515,N_15608,N_16530);
or U18516 (N_18516,N_15596,N_15537);
or U18517 (N_18517,N_15118,N_16075);
xor U18518 (N_18518,N_16875,N_17393);
nand U18519 (N_18519,N_17157,N_17295);
nor U18520 (N_18520,N_16296,N_16318);
nor U18521 (N_18521,N_17089,N_15992);
and U18522 (N_18522,N_17193,N_15919);
nand U18523 (N_18523,N_16402,N_17186);
nand U18524 (N_18524,N_15497,N_17078);
nor U18525 (N_18525,N_17057,N_17024);
and U18526 (N_18526,N_17183,N_17401);
xor U18527 (N_18527,N_16731,N_16802);
or U18528 (N_18528,N_16172,N_15428);
or U18529 (N_18529,N_15998,N_16040);
and U18530 (N_18530,N_15836,N_16929);
nor U18531 (N_18531,N_16077,N_16563);
xor U18532 (N_18532,N_17116,N_15902);
and U18533 (N_18533,N_15838,N_15518);
and U18534 (N_18534,N_16027,N_15752);
and U18535 (N_18535,N_16134,N_16116);
and U18536 (N_18536,N_15074,N_16712);
nand U18537 (N_18537,N_16136,N_15560);
or U18538 (N_18538,N_17375,N_17016);
nand U18539 (N_18539,N_16907,N_17104);
nor U18540 (N_18540,N_15043,N_15599);
or U18541 (N_18541,N_16023,N_15720);
nor U18542 (N_18542,N_16348,N_15129);
and U18543 (N_18543,N_15891,N_17380);
or U18544 (N_18544,N_16796,N_16900);
and U18545 (N_18545,N_17083,N_16453);
or U18546 (N_18546,N_16921,N_15920);
or U18547 (N_18547,N_15081,N_16868);
and U18548 (N_18548,N_15230,N_16987);
and U18549 (N_18549,N_15905,N_15360);
and U18550 (N_18550,N_16198,N_17233);
or U18551 (N_18551,N_15983,N_16833);
xnor U18552 (N_18552,N_15708,N_15520);
nor U18553 (N_18553,N_15017,N_17409);
nand U18554 (N_18554,N_16913,N_16973);
or U18555 (N_18555,N_16836,N_16052);
nand U18556 (N_18556,N_17305,N_16983);
nand U18557 (N_18557,N_16981,N_15789);
nand U18558 (N_18558,N_15572,N_16507);
and U18559 (N_18559,N_16630,N_16390);
or U18560 (N_18560,N_15756,N_15980);
or U18561 (N_18561,N_17292,N_16485);
nor U18562 (N_18562,N_15814,N_15152);
nand U18563 (N_18563,N_16426,N_16668);
xor U18564 (N_18564,N_16911,N_16038);
xnor U18565 (N_18565,N_17248,N_16922);
or U18566 (N_18566,N_17325,N_16697);
nand U18567 (N_18567,N_16462,N_16486);
or U18568 (N_18568,N_16250,N_17258);
or U18569 (N_18569,N_17163,N_17414);
and U18570 (N_18570,N_17397,N_17179);
xor U18571 (N_18571,N_17442,N_16589);
and U18572 (N_18572,N_16723,N_16740);
nand U18573 (N_18573,N_16349,N_15553);
or U18574 (N_18574,N_17369,N_15337);
or U18575 (N_18575,N_16698,N_16386);
nor U18576 (N_18576,N_16656,N_15533);
and U18577 (N_18577,N_17471,N_15346);
and U18578 (N_18578,N_17473,N_15579);
nand U18579 (N_18579,N_16528,N_17478);
or U18580 (N_18580,N_15332,N_15953);
nand U18581 (N_18581,N_16658,N_15178);
or U18582 (N_18582,N_15887,N_16963);
or U18583 (N_18583,N_15792,N_17249);
nor U18584 (N_18584,N_17394,N_16406);
and U18585 (N_18585,N_15362,N_16842);
or U18586 (N_18586,N_15578,N_16862);
xor U18587 (N_18587,N_15042,N_16024);
and U18588 (N_18588,N_16111,N_16264);
nand U18589 (N_18589,N_17126,N_15204);
or U18590 (N_18590,N_15941,N_17298);
nand U18591 (N_18591,N_17196,N_15628);
and U18592 (N_18592,N_15164,N_16861);
nand U18593 (N_18593,N_16097,N_16650);
or U18594 (N_18594,N_15120,N_17359);
and U18595 (N_18595,N_16781,N_16847);
nor U18596 (N_18596,N_15502,N_15826);
nand U18597 (N_18597,N_15593,N_17208);
or U18598 (N_18598,N_17014,N_16246);
xnor U18599 (N_18599,N_15227,N_15326);
or U18600 (N_18600,N_15461,N_15032);
and U18601 (N_18601,N_16192,N_16429);
or U18602 (N_18602,N_17408,N_17293);
or U18603 (N_18603,N_16456,N_15246);
nor U18604 (N_18604,N_16002,N_15096);
xor U18605 (N_18605,N_15804,N_16521);
nand U18606 (N_18606,N_16399,N_15741);
and U18607 (N_18607,N_15175,N_16721);
nand U18608 (N_18608,N_16845,N_16733);
and U18609 (N_18609,N_15094,N_15912);
nand U18610 (N_18610,N_15298,N_15512);
or U18611 (N_18611,N_16914,N_17469);
and U18612 (N_18612,N_15474,N_15718);
nand U18613 (N_18613,N_16672,N_15675);
nor U18614 (N_18614,N_17061,N_17491);
or U18615 (N_18615,N_17113,N_15287);
xnor U18616 (N_18616,N_17217,N_16959);
nor U18617 (N_18617,N_15729,N_15264);
nand U18618 (N_18618,N_16812,N_17074);
or U18619 (N_18619,N_15295,N_16347);
xor U18620 (N_18620,N_15875,N_17226);
or U18621 (N_18621,N_15420,N_17376);
nor U18622 (N_18622,N_15271,N_16613);
nor U18623 (N_18623,N_16209,N_16857);
nand U18624 (N_18624,N_17171,N_16642);
nor U18625 (N_18625,N_15190,N_17142);
and U18626 (N_18626,N_15507,N_17363);
nand U18627 (N_18627,N_16474,N_15317);
or U18628 (N_18628,N_16268,N_16855);
nand U18629 (N_18629,N_17134,N_15793);
nand U18630 (N_18630,N_16013,N_17411);
nand U18631 (N_18631,N_16470,N_15311);
nand U18632 (N_18632,N_15113,N_16622);
or U18633 (N_18633,N_15851,N_15280);
xnor U18634 (N_18634,N_16560,N_16251);
and U18635 (N_18635,N_16548,N_15339);
nand U18636 (N_18636,N_15934,N_15040);
or U18637 (N_18637,N_16835,N_16254);
nand U18638 (N_18638,N_15877,N_15594);
and U18639 (N_18639,N_17036,N_15558);
and U18640 (N_18640,N_16767,N_15965);
and U18641 (N_18641,N_15738,N_15285);
nand U18642 (N_18642,N_15087,N_17212);
nand U18643 (N_18643,N_17467,N_16335);
nand U18644 (N_18644,N_16945,N_16604);
xor U18645 (N_18645,N_15535,N_15481);
nor U18646 (N_18646,N_16196,N_17176);
and U18647 (N_18647,N_15422,N_15045);
nand U18648 (N_18648,N_15372,N_15177);
nor U18649 (N_18649,N_16699,N_17180);
or U18650 (N_18650,N_16798,N_15822);
nor U18651 (N_18651,N_16411,N_17385);
nor U18652 (N_18652,N_15526,N_16776);
nor U18653 (N_18653,N_16277,N_15319);
and U18654 (N_18654,N_16261,N_17330);
nand U18655 (N_18655,N_15090,N_17287);
xnor U18656 (N_18656,N_16314,N_16234);
nor U18657 (N_18657,N_16858,N_16720);
and U18658 (N_18658,N_17395,N_16883);
or U18659 (N_18659,N_17443,N_15490);
or U18660 (N_18660,N_15491,N_17336);
nor U18661 (N_18661,N_16829,N_15632);
nor U18662 (N_18662,N_15646,N_16508);
nor U18663 (N_18663,N_17334,N_16744);
or U18664 (N_18664,N_15892,N_16231);
or U18665 (N_18665,N_16141,N_16071);
or U18666 (N_18666,N_15110,N_16688);
and U18667 (N_18667,N_16523,N_15858);
and U18668 (N_18668,N_16976,N_17424);
nor U18669 (N_18669,N_16206,N_15034);
and U18670 (N_18670,N_15936,N_16850);
nand U18671 (N_18671,N_15837,N_15505);
or U18672 (N_18672,N_17028,N_16886);
nor U18673 (N_18673,N_17099,N_17058);
and U18674 (N_18674,N_17461,N_15003);
and U18675 (N_18675,N_17384,N_17434);
nand U18676 (N_18676,N_16372,N_16756);
and U18677 (N_18677,N_16041,N_15650);
nor U18678 (N_18678,N_16232,N_16803);
or U18679 (N_18679,N_16769,N_15092);
and U18680 (N_18680,N_16825,N_17119);
or U18681 (N_18681,N_15753,N_15811);
or U18682 (N_18682,N_16742,N_15931);
or U18683 (N_18683,N_15534,N_15704);
xor U18684 (N_18684,N_15263,N_16887);
xnor U18685 (N_18685,N_15613,N_17266);
or U18686 (N_18686,N_16061,N_15219);
nand U18687 (N_18687,N_15984,N_16415);
or U18688 (N_18688,N_16719,N_17118);
nor U18689 (N_18689,N_15914,N_15182);
nand U18690 (N_18690,N_16748,N_15817);
nor U18691 (N_18691,N_15010,N_17289);
or U18692 (N_18692,N_15528,N_15233);
or U18693 (N_18693,N_15721,N_15610);
and U18694 (N_18694,N_15278,N_16465);
nand U18695 (N_18695,N_16545,N_16674);
or U18696 (N_18696,N_17335,N_16202);
nand U18697 (N_18697,N_16941,N_16464);
nand U18698 (N_18698,N_16540,N_15925);
nand U18699 (N_18699,N_16127,N_17403);
nand U18700 (N_18700,N_16014,N_15207);
nor U18701 (N_18701,N_15960,N_15530);
and U18702 (N_18702,N_15252,N_15726);
and U18703 (N_18703,N_15847,N_15459);
or U18704 (N_18704,N_16450,N_16980);
nor U18705 (N_18705,N_16266,N_15119);
or U18706 (N_18706,N_16174,N_17131);
nand U18707 (N_18707,N_15725,N_16392);
nand U18708 (N_18708,N_15058,N_16635);
or U18709 (N_18709,N_17418,N_17276);
xnor U18710 (N_18710,N_17392,N_17260);
nor U18711 (N_18711,N_16284,N_15261);
or U18712 (N_18712,N_15552,N_16080);
nor U18713 (N_18713,N_16899,N_16294);
or U18714 (N_18714,N_15544,N_17441);
nor U18715 (N_18715,N_15815,N_15424);
and U18716 (N_18716,N_16778,N_17010);
nand U18717 (N_18717,N_16848,N_16216);
and U18718 (N_18718,N_16693,N_16534);
xor U18719 (N_18719,N_15539,N_15661);
and U18720 (N_18720,N_15504,N_15091);
nor U18721 (N_18721,N_16287,N_15141);
or U18722 (N_18722,N_15106,N_16276);
and U18723 (N_18723,N_16228,N_16966);
xnor U18724 (N_18724,N_15048,N_17049);
nor U18725 (N_18725,N_15312,N_17069);
and U18726 (N_18726,N_16611,N_16140);
nor U18727 (N_18727,N_16093,N_15224);
and U18728 (N_18728,N_16570,N_15603);
and U18729 (N_18729,N_16892,N_15667);
nand U18730 (N_18730,N_16304,N_16806);
and U18731 (N_18731,N_16317,N_15760);
and U18732 (N_18732,N_15415,N_15344);
and U18733 (N_18733,N_16716,N_15004);
nor U18734 (N_18734,N_16572,N_15654);
nand U18735 (N_18735,N_17278,N_15529);
and U18736 (N_18736,N_16943,N_17015);
xor U18737 (N_18737,N_17368,N_15574);
and U18738 (N_18738,N_17250,N_15131);
xor U18739 (N_18739,N_16036,N_16646);
and U18740 (N_18740,N_16420,N_16739);
xor U18741 (N_18741,N_15506,N_16285);
nand U18742 (N_18742,N_16632,N_15201);
or U18743 (N_18743,N_17422,N_15355);
and U18744 (N_18744,N_16021,N_16316);
xor U18745 (N_18745,N_17277,N_16819);
nand U18746 (N_18746,N_16290,N_15166);
nand U18747 (N_18747,N_16619,N_16584);
nor U18748 (N_18748,N_17312,N_16288);
and U18749 (N_18749,N_15679,N_16640);
nor U18750 (N_18750,N_15206,N_16806);
and U18751 (N_18751,N_16202,N_15309);
or U18752 (N_18752,N_15409,N_15285);
or U18753 (N_18753,N_15962,N_16321);
and U18754 (N_18754,N_15722,N_17467);
and U18755 (N_18755,N_16938,N_15727);
or U18756 (N_18756,N_16978,N_16419);
nor U18757 (N_18757,N_16691,N_17401);
nor U18758 (N_18758,N_15790,N_17456);
nor U18759 (N_18759,N_15100,N_16357);
nand U18760 (N_18760,N_15101,N_16366);
nor U18761 (N_18761,N_16436,N_15182);
and U18762 (N_18762,N_16125,N_16766);
xnor U18763 (N_18763,N_15871,N_16903);
nand U18764 (N_18764,N_16508,N_16706);
nor U18765 (N_18765,N_16681,N_17230);
nor U18766 (N_18766,N_16699,N_16090);
or U18767 (N_18767,N_16086,N_16630);
and U18768 (N_18768,N_16221,N_15829);
xor U18769 (N_18769,N_15383,N_16517);
nor U18770 (N_18770,N_15725,N_15250);
or U18771 (N_18771,N_16391,N_17318);
nor U18772 (N_18772,N_15341,N_15206);
nand U18773 (N_18773,N_16998,N_17326);
and U18774 (N_18774,N_16864,N_15155);
nor U18775 (N_18775,N_17460,N_17270);
or U18776 (N_18776,N_16492,N_16030);
nand U18777 (N_18777,N_15265,N_17189);
nand U18778 (N_18778,N_15141,N_16380);
or U18779 (N_18779,N_15399,N_17108);
xor U18780 (N_18780,N_16573,N_15653);
xnor U18781 (N_18781,N_16560,N_15828);
and U18782 (N_18782,N_17022,N_16000);
nand U18783 (N_18783,N_15678,N_15663);
xor U18784 (N_18784,N_17447,N_15036);
nand U18785 (N_18785,N_15785,N_17119);
nand U18786 (N_18786,N_15303,N_17117);
or U18787 (N_18787,N_17146,N_16998);
nand U18788 (N_18788,N_16855,N_16454);
nand U18789 (N_18789,N_17104,N_15836);
nand U18790 (N_18790,N_15117,N_16218);
nor U18791 (N_18791,N_15420,N_15472);
or U18792 (N_18792,N_16784,N_15561);
or U18793 (N_18793,N_17138,N_16513);
nand U18794 (N_18794,N_16874,N_16751);
or U18795 (N_18795,N_17445,N_16789);
or U18796 (N_18796,N_16271,N_17310);
xnor U18797 (N_18797,N_17238,N_15904);
and U18798 (N_18798,N_15879,N_17194);
nand U18799 (N_18799,N_16945,N_16441);
and U18800 (N_18800,N_15794,N_15963);
nor U18801 (N_18801,N_17493,N_15724);
or U18802 (N_18802,N_15337,N_17155);
nor U18803 (N_18803,N_16885,N_17139);
and U18804 (N_18804,N_15632,N_17165);
xnor U18805 (N_18805,N_15980,N_15500);
xnor U18806 (N_18806,N_15313,N_16247);
nor U18807 (N_18807,N_15774,N_15962);
nand U18808 (N_18808,N_15857,N_17065);
or U18809 (N_18809,N_15929,N_16023);
or U18810 (N_18810,N_17036,N_16570);
and U18811 (N_18811,N_15068,N_16996);
or U18812 (N_18812,N_15412,N_16577);
nand U18813 (N_18813,N_15129,N_17043);
nand U18814 (N_18814,N_16311,N_16157);
xor U18815 (N_18815,N_16542,N_16642);
nand U18816 (N_18816,N_16122,N_17449);
xor U18817 (N_18817,N_16154,N_16433);
nor U18818 (N_18818,N_15061,N_16291);
and U18819 (N_18819,N_16681,N_16358);
nand U18820 (N_18820,N_15084,N_15543);
nor U18821 (N_18821,N_17495,N_17012);
nand U18822 (N_18822,N_16571,N_15444);
nand U18823 (N_18823,N_16335,N_17286);
and U18824 (N_18824,N_16190,N_15426);
nor U18825 (N_18825,N_15828,N_17301);
and U18826 (N_18826,N_17375,N_16439);
or U18827 (N_18827,N_17076,N_16540);
and U18828 (N_18828,N_17290,N_15340);
or U18829 (N_18829,N_16071,N_17104);
and U18830 (N_18830,N_16908,N_15904);
nand U18831 (N_18831,N_17293,N_16947);
and U18832 (N_18832,N_16409,N_16344);
nand U18833 (N_18833,N_16598,N_16334);
nand U18834 (N_18834,N_16487,N_16403);
nand U18835 (N_18835,N_15584,N_16336);
and U18836 (N_18836,N_15467,N_15221);
nor U18837 (N_18837,N_16656,N_16972);
nor U18838 (N_18838,N_15344,N_16465);
xor U18839 (N_18839,N_17141,N_17259);
nor U18840 (N_18840,N_16170,N_17194);
nor U18841 (N_18841,N_17483,N_16992);
or U18842 (N_18842,N_15444,N_16142);
nand U18843 (N_18843,N_17499,N_15211);
nor U18844 (N_18844,N_17321,N_16402);
xnor U18845 (N_18845,N_17327,N_15802);
nor U18846 (N_18846,N_17461,N_16106);
nor U18847 (N_18847,N_15063,N_15940);
nor U18848 (N_18848,N_16937,N_17256);
nand U18849 (N_18849,N_15158,N_16624);
nand U18850 (N_18850,N_15354,N_15727);
nand U18851 (N_18851,N_15275,N_16421);
and U18852 (N_18852,N_16831,N_16374);
nand U18853 (N_18853,N_16966,N_15452);
nand U18854 (N_18854,N_17117,N_17347);
or U18855 (N_18855,N_17271,N_16583);
nand U18856 (N_18856,N_17341,N_17022);
and U18857 (N_18857,N_16513,N_16267);
or U18858 (N_18858,N_15038,N_15267);
or U18859 (N_18859,N_17431,N_16598);
nand U18860 (N_18860,N_16852,N_16790);
nor U18861 (N_18861,N_15988,N_16374);
nand U18862 (N_18862,N_16160,N_15730);
nor U18863 (N_18863,N_17128,N_15468);
nand U18864 (N_18864,N_15268,N_16293);
nand U18865 (N_18865,N_15861,N_15567);
and U18866 (N_18866,N_15642,N_15119);
and U18867 (N_18867,N_15985,N_15491);
and U18868 (N_18868,N_16837,N_15100);
nor U18869 (N_18869,N_15596,N_16685);
and U18870 (N_18870,N_17019,N_15549);
nor U18871 (N_18871,N_15177,N_17196);
or U18872 (N_18872,N_17425,N_16995);
and U18873 (N_18873,N_16530,N_15816);
nor U18874 (N_18874,N_15209,N_15561);
nor U18875 (N_18875,N_17270,N_15841);
and U18876 (N_18876,N_15681,N_15486);
xnor U18877 (N_18877,N_17308,N_16456);
nor U18878 (N_18878,N_15016,N_16695);
or U18879 (N_18879,N_16320,N_15509);
nor U18880 (N_18880,N_15959,N_15305);
and U18881 (N_18881,N_15340,N_16610);
and U18882 (N_18882,N_16116,N_15831);
nor U18883 (N_18883,N_16440,N_17416);
nand U18884 (N_18884,N_15626,N_15764);
or U18885 (N_18885,N_16750,N_16094);
nor U18886 (N_18886,N_15750,N_15605);
or U18887 (N_18887,N_16699,N_15891);
nor U18888 (N_18888,N_16872,N_15783);
nor U18889 (N_18889,N_16960,N_17326);
or U18890 (N_18890,N_17493,N_16395);
nor U18891 (N_18891,N_17137,N_17160);
xnor U18892 (N_18892,N_15882,N_16860);
nand U18893 (N_18893,N_15280,N_15861);
nor U18894 (N_18894,N_16252,N_16391);
or U18895 (N_18895,N_16860,N_16833);
or U18896 (N_18896,N_17305,N_17420);
nor U18897 (N_18897,N_16068,N_17460);
and U18898 (N_18898,N_15638,N_16961);
and U18899 (N_18899,N_15426,N_15947);
and U18900 (N_18900,N_17005,N_17047);
nand U18901 (N_18901,N_15099,N_15969);
nor U18902 (N_18902,N_16251,N_16019);
or U18903 (N_18903,N_15657,N_17186);
or U18904 (N_18904,N_17383,N_16851);
nor U18905 (N_18905,N_16264,N_15502);
nand U18906 (N_18906,N_16487,N_17292);
nand U18907 (N_18907,N_17321,N_16831);
nor U18908 (N_18908,N_17002,N_16887);
and U18909 (N_18909,N_17207,N_15027);
nor U18910 (N_18910,N_15324,N_16859);
nor U18911 (N_18911,N_16861,N_16780);
nand U18912 (N_18912,N_17308,N_17021);
nand U18913 (N_18913,N_17186,N_15096);
nand U18914 (N_18914,N_16306,N_16012);
nand U18915 (N_18915,N_16453,N_15917);
or U18916 (N_18916,N_16307,N_15922);
nor U18917 (N_18917,N_15063,N_17037);
xnor U18918 (N_18918,N_15421,N_15337);
xor U18919 (N_18919,N_17412,N_16674);
nand U18920 (N_18920,N_15693,N_15390);
or U18921 (N_18921,N_16799,N_16062);
or U18922 (N_18922,N_16447,N_16232);
nor U18923 (N_18923,N_17185,N_16655);
and U18924 (N_18924,N_15994,N_15189);
or U18925 (N_18925,N_16637,N_17261);
nand U18926 (N_18926,N_15456,N_15555);
nand U18927 (N_18927,N_16884,N_15363);
and U18928 (N_18928,N_16493,N_17406);
nor U18929 (N_18929,N_16049,N_15316);
or U18930 (N_18930,N_16652,N_16842);
nor U18931 (N_18931,N_16762,N_16025);
or U18932 (N_18932,N_15828,N_17157);
nand U18933 (N_18933,N_16656,N_16416);
nor U18934 (N_18934,N_15587,N_16541);
and U18935 (N_18935,N_15932,N_15501);
or U18936 (N_18936,N_15107,N_17479);
nand U18937 (N_18937,N_15780,N_15303);
and U18938 (N_18938,N_16293,N_16679);
or U18939 (N_18939,N_15684,N_17360);
and U18940 (N_18940,N_17383,N_16371);
and U18941 (N_18941,N_17166,N_15717);
and U18942 (N_18942,N_17055,N_17023);
nor U18943 (N_18943,N_15722,N_16686);
nand U18944 (N_18944,N_16704,N_15533);
and U18945 (N_18945,N_15956,N_15662);
xnor U18946 (N_18946,N_16063,N_15890);
nor U18947 (N_18947,N_15296,N_15948);
and U18948 (N_18948,N_15230,N_17019);
and U18949 (N_18949,N_16500,N_17478);
nor U18950 (N_18950,N_15459,N_15635);
and U18951 (N_18951,N_16469,N_17274);
and U18952 (N_18952,N_16983,N_17382);
nand U18953 (N_18953,N_16411,N_16982);
nand U18954 (N_18954,N_16706,N_15071);
nand U18955 (N_18955,N_16723,N_17387);
and U18956 (N_18956,N_17339,N_15819);
or U18957 (N_18957,N_16736,N_15028);
or U18958 (N_18958,N_16821,N_17239);
and U18959 (N_18959,N_16085,N_17086);
xnor U18960 (N_18960,N_15050,N_17445);
or U18961 (N_18961,N_16701,N_15799);
or U18962 (N_18962,N_16112,N_15933);
nand U18963 (N_18963,N_16296,N_15673);
nand U18964 (N_18964,N_16907,N_15055);
and U18965 (N_18965,N_15380,N_16028);
nor U18966 (N_18966,N_17184,N_16738);
or U18967 (N_18967,N_17414,N_15075);
nor U18968 (N_18968,N_17002,N_17249);
nand U18969 (N_18969,N_15552,N_17105);
nand U18970 (N_18970,N_16153,N_17109);
nor U18971 (N_18971,N_15496,N_16779);
nand U18972 (N_18972,N_15198,N_16941);
nor U18973 (N_18973,N_16910,N_15381);
nor U18974 (N_18974,N_15859,N_16124);
nor U18975 (N_18975,N_15306,N_17298);
xnor U18976 (N_18976,N_15585,N_15237);
xor U18977 (N_18977,N_15721,N_16654);
nand U18978 (N_18978,N_15698,N_16247);
xnor U18979 (N_18979,N_15848,N_15122);
nor U18980 (N_18980,N_15480,N_16960);
and U18981 (N_18981,N_15497,N_17387);
and U18982 (N_18982,N_15827,N_15590);
or U18983 (N_18983,N_15260,N_16533);
nand U18984 (N_18984,N_16419,N_16272);
nor U18985 (N_18985,N_17287,N_15216);
nand U18986 (N_18986,N_15765,N_15621);
nand U18987 (N_18987,N_16010,N_16081);
nor U18988 (N_18988,N_16462,N_17069);
nand U18989 (N_18989,N_17490,N_15584);
and U18990 (N_18990,N_15511,N_15986);
nor U18991 (N_18991,N_15774,N_16208);
nand U18992 (N_18992,N_15620,N_16081);
nand U18993 (N_18993,N_16441,N_17462);
or U18994 (N_18994,N_16919,N_17154);
and U18995 (N_18995,N_15961,N_15361);
or U18996 (N_18996,N_17002,N_15034);
or U18997 (N_18997,N_15067,N_16764);
nand U18998 (N_18998,N_15084,N_16637);
or U18999 (N_18999,N_15558,N_17352);
and U19000 (N_19000,N_15477,N_15758);
and U19001 (N_19001,N_16515,N_15588);
and U19002 (N_19002,N_16646,N_15796);
and U19003 (N_19003,N_17026,N_16485);
xnor U19004 (N_19004,N_17186,N_15357);
nand U19005 (N_19005,N_16744,N_16617);
nand U19006 (N_19006,N_17009,N_15773);
and U19007 (N_19007,N_16760,N_16491);
nand U19008 (N_19008,N_15770,N_17428);
xnor U19009 (N_19009,N_17070,N_15121);
or U19010 (N_19010,N_17386,N_16130);
nor U19011 (N_19011,N_16153,N_15025);
or U19012 (N_19012,N_16627,N_16003);
and U19013 (N_19013,N_16696,N_15066);
or U19014 (N_19014,N_16409,N_15826);
xor U19015 (N_19015,N_16790,N_17143);
or U19016 (N_19016,N_15531,N_17469);
and U19017 (N_19017,N_16014,N_15359);
and U19018 (N_19018,N_15309,N_15868);
nor U19019 (N_19019,N_16509,N_16695);
and U19020 (N_19020,N_15912,N_15613);
and U19021 (N_19021,N_15004,N_16127);
and U19022 (N_19022,N_16699,N_16353);
or U19023 (N_19023,N_15510,N_16502);
and U19024 (N_19024,N_16464,N_16340);
and U19025 (N_19025,N_16767,N_17355);
and U19026 (N_19026,N_15350,N_15195);
or U19027 (N_19027,N_16011,N_15340);
nand U19028 (N_19028,N_15726,N_15663);
nand U19029 (N_19029,N_17057,N_16801);
and U19030 (N_19030,N_15618,N_15204);
nor U19031 (N_19031,N_16005,N_16168);
nand U19032 (N_19032,N_17255,N_15088);
nand U19033 (N_19033,N_16553,N_15532);
nand U19034 (N_19034,N_17388,N_15214);
nand U19035 (N_19035,N_16816,N_16614);
or U19036 (N_19036,N_15693,N_16459);
nor U19037 (N_19037,N_16124,N_16802);
and U19038 (N_19038,N_15014,N_17060);
nand U19039 (N_19039,N_16104,N_16115);
nand U19040 (N_19040,N_16270,N_16548);
nor U19041 (N_19041,N_17178,N_17168);
nand U19042 (N_19042,N_15333,N_16843);
and U19043 (N_19043,N_15612,N_15954);
nor U19044 (N_19044,N_16731,N_15811);
or U19045 (N_19045,N_15626,N_16367);
or U19046 (N_19046,N_16326,N_17137);
or U19047 (N_19047,N_17200,N_16926);
and U19048 (N_19048,N_16528,N_17043);
xnor U19049 (N_19049,N_17095,N_16458);
and U19050 (N_19050,N_16976,N_15256);
nand U19051 (N_19051,N_17498,N_16988);
and U19052 (N_19052,N_15615,N_17283);
xnor U19053 (N_19053,N_16751,N_16667);
nand U19054 (N_19054,N_15124,N_17194);
nor U19055 (N_19055,N_17413,N_16107);
nand U19056 (N_19056,N_17132,N_16411);
nand U19057 (N_19057,N_16202,N_17017);
nand U19058 (N_19058,N_17257,N_16351);
or U19059 (N_19059,N_17449,N_16834);
and U19060 (N_19060,N_17096,N_15300);
and U19061 (N_19061,N_15830,N_16775);
or U19062 (N_19062,N_15887,N_16720);
nor U19063 (N_19063,N_15823,N_17320);
nand U19064 (N_19064,N_15645,N_16965);
or U19065 (N_19065,N_17328,N_15201);
and U19066 (N_19066,N_15482,N_16975);
nand U19067 (N_19067,N_15998,N_17285);
xnor U19068 (N_19068,N_15111,N_15516);
and U19069 (N_19069,N_15027,N_15411);
nor U19070 (N_19070,N_15935,N_15882);
nor U19071 (N_19071,N_15246,N_15879);
and U19072 (N_19072,N_17197,N_15767);
and U19073 (N_19073,N_16467,N_15468);
nor U19074 (N_19074,N_17253,N_15850);
nand U19075 (N_19075,N_17401,N_15145);
nand U19076 (N_19076,N_17027,N_17486);
nand U19077 (N_19077,N_15365,N_15913);
nor U19078 (N_19078,N_17249,N_16967);
and U19079 (N_19079,N_16273,N_15242);
and U19080 (N_19080,N_15363,N_15541);
and U19081 (N_19081,N_15060,N_16397);
or U19082 (N_19082,N_17358,N_17146);
nand U19083 (N_19083,N_16837,N_15266);
or U19084 (N_19084,N_15030,N_16049);
or U19085 (N_19085,N_15732,N_15945);
xnor U19086 (N_19086,N_16754,N_16552);
and U19087 (N_19087,N_15287,N_15898);
nand U19088 (N_19088,N_15633,N_16062);
nor U19089 (N_19089,N_16409,N_15165);
and U19090 (N_19090,N_16308,N_17253);
and U19091 (N_19091,N_17189,N_16876);
or U19092 (N_19092,N_16441,N_15413);
nor U19093 (N_19093,N_16694,N_16811);
nand U19094 (N_19094,N_16868,N_15136);
xor U19095 (N_19095,N_15737,N_15814);
nand U19096 (N_19096,N_16417,N_17332);
nand U19097 (N_19097,N_15465,N_17228);
nor U19098 (N_19098,N_15589,N_16009);
nand U19099 (N_19099,N_15745,N_16273);
or U19100 (N_19100,N_15356,N_15144);
and U19101 (N_19101,N_16217,N_17149);
nor U19102 (N_19102,N_16872,N_16462);
xnor U19103 (N_19103,N_17022,N_16944);
nand U19104 (N_19104,N_16112,N_15246);
nor U19105 (N_19105,N_15287,N_16719);
nand U19106 (N_19106,N_16122,N_16006);
and U19107 (N_19107,N_15042,N_15278);
or U19108 (N_19108,N_15223,N_16351);
nor U19109 (N_19109,N_16688,N_16654);
or U19110 (N_19110,N_17493,N_16672);
nand U19111 (N_19111,N_15086,N_17339);
or U19112 (N_19112,N_17157,N_15564);
nand U19113 (N_19113,N_15098,N_15427);
or U19114 (N_19114,N_16774,N_15064);
nand U19115 (N_19115,N_15843,N_15666);
and U19116 (N_19116,N_17300,N_17443);
nand U19117 (N_19117,N_17067,N_16216);
and U19118 (N_19118,N_15647,N_16055);
nand U19119 (N_19119,N_17367,N_16494);
or U19120 (N_19120,N_16664,N_16455);
and U19121 (N_19121,N_15068,N_17214);
or U19122 (N_19122,N_15747,N_16449);
nor U19123 (N_19123,N_15744,N_15694);
or U19124 (N_19124,N_17311,N_16735);
or U19125 (N_19125,N_15490,N_17374);
or U19126 (N_19126,N_15015,N_15768);
nor U19127 (N_19127,N_17398,N_15098);
nor U19128 (N_19128,N_16695,N_15707);
xor U19129 (N_19129,N_16722,N_16038);
and U19130 (N_19130,N_15279,N_17242);
nand U19131 (N_19131,N_15244,N_15096);
nor U19132 (N_19132,N_17383,N_15656);
nand U19133 (N_19133,N_17170,N_16094);
nor U19134 (N_19134,N_15413,N_16649);
nor U19135 (N_19135,N_15628,N_16410);
xnor U19136 (N_19136,N_16244,N_16847);
or U19137 (N_19137,N_15419,N_17055);
xor U19138 (N_19138,N_15891,N_15547);
or U19139 (N_19139,N_17481,N_16546);
nor U19140 (N_19140,N_16952,N_15649);
and U19141 (N_19141,N_17125,N_15563);
and U19142 (N_19142,N_16980,N_17438);
or U19143 (N_19143,N_15871,N_15977);
and U19144 (N_19144,N_15503,N_16181);
nand U19145 (N_19145,N_16988,N_17160);
nand U19146 (N_19146,N_15484,N_16072);
nand U19147 (N_19147,N_15374,N_17108);
nand U19148 (N_19148,N_16472,N_16888);
and U19149 (N_19149,N_16539,N_15440);
nand U19150 (N_19150,N_16545,N_16763);
nand U19151 (N_19151,N_16596,N_16175);
or U19152 (N_19152,N_16503,N_17042);
nand U19153 (N_19153,N_15191,N_17277);
or U19154 (N_19154,N_16757,N_17156);
nor U19155 (N_19155,N_17287,N_15256);
and U19156 (N_19156,N_15448,N_15750);
nor U19157 (N_19157,N_15806,N_16953);
and U19158 (N_19158,N_15605,N_17237);
nand U19159 (N_19159,N_15248,N_15235);
nand U19160 (N_19160,N_15202,N_15980);
nor U19161 (N_19161,N_15818,N_16774);
nor U19162 (N_19162,N_17498,N_15426);
xor U19163 (N_19163,N_15988,N_16049);
xor U19164 (N_19164,N_16297,N_16216);
nand U19165 (N_19165,N_17256,N_15617);
xor U19166 (N_19166,N_17391,N_16232);
nand U19167 (N_19167,N_16538,N_16475);
or U19168 (N_19168,N_16801,N_16850);
nand U19169 (N_19169,N_17049,N_16167);
and U19170 (N_19170,N_16043,N_15665);
and U19171 (N_19171,N_16769,N_15363);
nand U19172 (N_19172,N_15524,N_15621);
nand U19173 (N_19173,N_15812,N_15480);
nor U19174 (N_19174,N_17204,N_17487);
nand U19175 (N_19175,N_17223,N_15914);
and U19176 (N_19176,N_16780,N_17269);
nor U19177 (N_19177,N_15548,N_17236);
nand U19178 (N_19178,N_16716,N_16766);
or U19179 (N_19179,N_17371,N_15357);
or U19180 (N_19180,N_16293,N_16288);
and U19181 (N_19181,N_15708,N_16863);
and U19182 (N_19182,N_17017,N_16237);
nand U19183 (N_19183,N_16009,N_15015);
and U19184 (N_19184,N_17460,N_17132);
nor U19185 (N_19185,N_15840,N_17210);
and U19186 (N_19186,N_15625,N_15189);
or U19187 (N_19187,N_15865,N_16556);
nand U19188 (N_19188,N_15154,N_17139);
and U19189 (N_19189,N_16000,N_16424);
nand U19190 (N_19190,N_15370,N_17297);
or U19191 (N_19191,N_15581,N_17061);
nand U19192 (N_19192,N_16225,N_16809);
nor U19193 (N_19193,N_15072,N_15854);
nor U19194 (N_19194,N_16325,N_16560);
nor U19195 (N_19195,N_16289,N_15029);
nand U19196 (N_19196,N_15358,N_16794);
nor U19197 (N_19197,N_17165,N_15736);
and U19198 (N_19198,N_17259,N_16201);
or U19199 (N_19199,N_16255,N_16461);
nor U19200 (N_19200,N_17346,N_15889);
nor U19201 (N_19201,N_17370,N_16925);
or U19202 (N_19202,N_16411,N_17383);
and U19203 (N_19203,N_15076,N_17238);
or U19204 (N_19204,N_15300,N_16176);
and U19205 (N_19205,N_15157,N_16575);
nand U19206 (N_19206,N_15071,N_15632);
or U19207 (N_19207,N_16444,N_17112);
and U19208 (N_19208,N_15543,N_17205);
or U19209 (N_19209,N_17016,N_16855);
nor U19210 (N_19210,N_17231,N_15492);
and U19211 (N_19211,N_16757,N_15135);
and U19212 (N_19212,N_15459,N_16410);
xnor U19213 (N_19213,N_15906,N_16947);
and U19214 (N_19214,N_15201,N_16790);
nor U19215 (N_19215,N_17236,N_17218);
or U19216 (N_19216,N_15395,N_15763);
nand U19217 (N_19217,N_15902,N_17438);
and U19218 (N_19218,N_17026,N_15076);
or U19219 (N_19219,N_15623,N_15575);
nor U19220 (N_19220,N_15472,N_15374);
nand U19221 (N_19221,N_15372,N_16028);
and U19222 (N_19222,N_17258,N_17217);
and U19223 (N_19223,N_16225,N_16748);
or U19224 (N_19224,N_15735,N_17174);
nand U19225 (N_19225,N_15827,N_15011);
nand U19226 (N_19226,N_15401,N_15879);
xnor U19227 (N_19227,N_17108,N_15755);
and U19228 (N_19228,N_15040,N_15736);
nand U19229 (N_19229,N_16865,N_17317);
nand U19230 (N_19230,N_17247,N_17462);
nor U19231 (N_19231,N_16818,N_16723);
or U19232 (N_19232,N_16050,N_17045);
nor U19233 (N_19233,N_15357,N_17375);
nand U19234 (N_19234,N_17180,N_16837);
xnor U19235 (N_19235,N_16245,N_17149);
or U19236 (N_19236,N_16194,N_16113);
nand U19237 (N_19237,N_15945,N_16937);
or U19238 (N_19238,N_16516,N_15019);
or U19239 (N_19239,N_15176,N_16959);
or U19240 (N_19240,N_17416,N_15083);
nor U19241 (N_19241,N_16224,N_17313);
and U19242 (N_19242,N_16544,N_16902);
nand U19243 (N_19243,N_16214,N_17428);
and U19244 (N_19244,N_17160,N_16948);
nor U19245 (N_19245,N_17313,N_15835);
or U19246 (N_19246,N_16552,N_15829);
nand U19247 (N_19247,N_17262,N_15543);
or U19248 (N_19248,N_15547,N_16697);
and U19249 (N_19249,N_16287,N_16746);
nor U19250 (N_19250,N_15877,N_16857);
and U19251 (N_19251,N_15628,N_16121);
nand U19252 (N_19252,N_16341,N_16131);
or U19253 (N_19253,N_16979,N_15426);
and U19254 (N_19254,N_16680,N_17026);
nand U19255 (N_19255,N_16941,N_16363);
nand U19256 (N_19256,N_16905,N_16238);
nand U19257 (N_19257,N_15965,N_16393);
and U19258 (N_19258,N_16089,N_17289);
nand U19259 (N_19259,N_15049,N_16421);
xor U19260 (N_19260,N_17144,N_16729);
nor U19261 (N_19261,N_15167,N_17190);
nor U19262 (N_19262,N_16635,N_16456);
or U19263 (N_19263,N_17478,N_15230);
nor U19264 (N_19264,N_16938,N_16229);
nor U19265 (N_19265,N_16095,N_15459);
nand U19266 (N_19266,N_15990,N_16746);
nand U19267 (N_19267,N_16782,N_15407);
nor U19268 (N_19268,N_15385,N_15313);
or U19269 (N_19269,N_15832,N_15524);
xnor U19270 (N_19270,N_17203,N_16777);
nor U19271 (N_19271,N_16134,N_15107);
nand U19272 (N_19272,N_16715,N_15369);
and U19273 (N_19273,N_17034,N_17452);
nand U19274 (N_19274,N_16977,N_15201);
or U19275 (N_19275,N_17389,N_16173);
nor U19276 (N_19276,N_15688,N_17079);
or U19277 (N_19277,N_16016,N_17012);
or U19278 (N_19278,N_16967,N_16722);
and U19279 (N_19279,N_16530,N_16434);
nand U19280 (N_19280,N_16335,N_15144);
nor U19281 (N_19281,N_15980,N_17287);
xor U19282 (N_19282,N_15714,N_15063);
nand U19283 (N_19283,N_16609,N_15060);
nor U19284 (N_19284,N_15996,N_17218);
nand U19285 (N_19285,N_16124,N_16912);
and U19286 (N_19286,N_15326,N_15098);
nor U19287 (N_19287,N_15431,N_16148);
or U19288 (N_19288,N_17269,N_17398);
and U19289 (N_19289,N_16600,N_17484);
nor U19290 (N_19290,N_15070,N_16165);
nand U19291 (N_19291,N_15248,N_16249);
nor U19292 (N_19292,N_15447,N_16585);
or U19293 (N_19293,N_16443,N_16796);
and U19294 (N_19294,N_17094,N_15147);
and U19295 (N_19295,N_15218,N_15415);
nor U19296 (N_19296,N_15439,N_17251);
nand U19297 (N_19297,N_16814,N_15913);
nand U19298 (N_19298,N_16702,N_16850);
xor U19299 (N_19299,N_16440,N_15044);
and U19300 (N_19300,N_16687,N_17460);
nor U19301 (N_19301,N_16007,N_17237);
nor U19302 (N_19302,N_17441,N_16344);
nor U19303 (N_19303,N_15908,N_16549);
xor U19304 (N_19304,N_17139,N_15300);
and U19305 (N_19305,N_15694,N_17056);
or U19306 (N_19306,N_15237,N_16784);
and U19307 (N_19307,N_15328,N_16609);
and U19308 (N_19308,N_15796,N_15409);
nand U19309 (N_19309,N_15910,N_16776);
nor U19310 (N_19310,N_17359,N_16199);
nor U19311 (N_19311,N_16262,N_15332);
or U19312 (N_19312,N_17166,N_17170);
and U19313 (N_19313,N_16183,N_16711);
or U19314 (N_19314,N_15659,N_16140);
or U19315 (N_19315,N_17183,N_17223);
nor U19316 (N_19316,N_16787,N_16109);
and U19317 (N_19317,N_16650,N_15813);
or U19318 (N_19318,N_17493,N_16729);
or U19319 (N_19319,N_16784,N_15304);
nand U19320 (N_19320,N_16686,N_15184);
nand U19321 (N_19321,N_16567,N_17154);
xnor U19322 (N_19322,N_15649,N_15202);
and U19323 (N_19323,N_15015,N_16239);
nor U19324 (N_19324,N_16696,N_16399);
and U19325 (N_19325,N_16515,N_17025);
nand U19326 (N_19326,N_17373,N_17072);
nand U19327 (N_19327,N_17481,N_16164);
and U19328 (N_19328,N_17157,N_16228);
nor U19329 (N_19329,N_15745,N_15515);
or U19330 (N_19330,N_16249,N_15729);
and U19331 (N_19331,N_17330,N_16727);
nor U19332 (N_19332,N_15054,N_15218);
and U19333 (N_19333,N_15064,N_16648);
nor U19334 (N_19334,N_16956,N_15871);
or U19335 (N_19335,N_15357,N_15124);
and U19336 (N_19336,N_15510,N_16586);
or U19337 (N_19337,N_15456,N_16479);
and U19338 (N_19338,N_17093,N_16628);
nor U19339 (N_19339,N_17315,N_15507);
nand U19340 (N_19340,N_16007,N_15629);
nor U19341 (N_19341,N_16869,N_16390);
and U19342 (N_19342,N_16568,N_17169);
and U19343 (N_19343,N_17295,N_15384);
nand U19344 (N_19344,N_15080,N_17389);
and U19345 (N_19345,N_16200,N_15922);
or U19346 (N_19346,N_17103,N_15120);
or U19347 (N_19347,N_16084,N_15552);
nor U19348 (N_19348,N_15912,N_17435);
xor U19349 (N_19349,N_16126,N_15036);
and U19350 (N_19350,N_17402,N_17290);
nor U19351 (N_19351,N_17398,N_15380);
nor U19352 (N_19352,N_15181,N_17213);
and U19353 (N_19353,N_16138,N_17125);
and U19354 (N_19354,N_15921,N_16276);
xnor U19355 (N_19355,N_16090,N_15357);
and U19356 (N_19356,N_16333,N_16426);
nor U19357 (N_19357,N_16433,N_17168);
xor U19358 (N_19358,N_16512,N_15660);
nand U19359 (N_19359,N_15502,N_16243);
nor U19360 (N_19360,N_15584,N_15604);
and U19361 (N_19361,N_15990,N_16919);
nand U19362 (N_19362,N_15116,N_15862);
nor U19363 (N_19363,N_17486,N_17478);
or U19364 (N_19364,N_16661,N_16711);
and U19365 (N_19365,N_17371,N_15289);
and U19366 (N_19366,N_17144,N_16962);
nor U19367 (N_19367,N_15331,N_15925);
xor U19368 (N_19368,N_16460,N_17429);
and U19369 (N_19369,N_17397,N_15309);
or U19370 (N_19370,N_16716,N_17391);
and U19371 (N_19371,N_15287,N_16267);
and U19372 (N_19372,N_17298,N_15799);
or U19373 (N_19373,N_16832,N_16595);
or U19374 (N_19374,N_16177,N_15902);
nand U19375 (N_19375,N_17292,N_16415);
and U19376 (N_19376,N_16022,N_15229);
nand U19377 (N_19377,N_17301,N_17107);
or U19378 (N_19378,N_16486,N_17329);
or U19379 (N_19379,N_16128,N_15073);
or U19380 (N_19380,N_15007,N_16103);
and U19381 (N_19381,N_16751,N_16127);
nor U19382 (N_19382,N_17267,N_15196);
nand U19383 (N_19383,N_15857,N_17475);
or U19384 (N_19384,N_16144,N_16341);
nor U19385 (N_19385,N_16715,N_15302);
or U19386 (N_19386,N_15223,N_16961);
xnor U19387 (N_19387,N_15357,N_16158);
nor U19388 (N_19388,N_15133,N_15976);
or U19389 (N_19389,N_16815,N_16584);
nand U19390 (N_19390,N_15297,N_15394);
nor U19391 (N_19391,N_17361,N_15768);
nor U19392 (N_19392,N_16835,N_16963);
and U19393 (N_19393,N_16378,N_15810);
xnor U19394 (N_19394,N_15012,N_16323);
nor U19395 (N_19395,N_15010,N_15995);
xnor U19396 (N_19396,N_15495,N_16479);
nand U19397 (N_19397,N_16105,N_15170);
nor U19398 (N_19398,N_15445,N_15366);
xnor U19399 (N_19399,N_17387,N_16462);
nor U19400 (N_19400,N_16005,N_15347);
and U19401 (N_19401,N_16021,N_16244);
nor U19402 (N_19402,N_15872,N_17268);
nand U19403 (N_19403,N_17125,N_15177);
xor U19404 (N_19404,N_16221,N_17467);
and U19405 (N_19405,N_17312,N_16646);
xor U19406 (N_19406,N_15135,N_17176);
and U19407 (N_19407,N_16354,N_16103);
nor U19408 (N_19408,N_15758,N_17055);
nor U19409 (N_19409,N_16188,N_17032);
nand U19410 (N_19410,N_17323,N_15117);
nor U19411 (N_19411,N_16005,N_15022);
or U19412 (N_19412,N_16953,N_16647);
xnor U19413 (N_19413,N_15645,N_15377);
nor U19414 (N_19414,N_16618,N_16801);
and U19415 (N_19415,N_17053,N_17396);
nand U19416 (N_19416,N_17336,N_15708);
xnor U19417 (N_19417,N_16414,N_17173);
and U19418 (N_19418,N_16416,N_16515);
and U19419 (N_19419,N_16275,N_16288);
nor U19420 (N_19420,N_15412,N_15343);
nor U19421 (N_19421,N_16609,N_15545);
nor U19422 (N_19422,N_15523,N_15171);
or U19423 (N_19423,N_16640,N_16382);
xnor U19424 (N_19424,N_16072,N_17112);
or U19425 (N_19425,N_16264,N_16339);
and U19426 (N_19426,N_17105,N_16000);
nand U19427 (N_19427,N_15992,N_17320);
nand U19428 (N_19428,N_15508,N_16014);
xnor U19429 (N_19429,N_15301,N_16420);
nand U19430 (N_19430,N_15561,N_16889);
nand U19431 (N_19431,N_17052,N_17391);
and U19432 (N_19432,N_16608,N_15379);
nor U19433 (N_19433,N_15830,N_15510);
nor U19434 (N_19434,N_16183,N_17227);
or U19435 (N_19435,N_15048,N_16459);
nand U19436 (N_19436,N_15054,N_16570);
nand U19437 (N_19437,N_15113,N_15048);
nand U19438 (N_19438,N_16922,N_17085);
or U19439 (N_19439,N_16788,N_17232);
nand U19440 (N_19440,N_17124,N_15043);
or U19441 (N_19441,N_15756,N_15056);
and U19442 (N_19442,N_16848,N_16659);
or U19443 (N_19443,N_16432,N_17078);
nand U19444 (N_19444,N_15026,N_15906);
and U19445 (N_19445,N_15556,N_15925);
xnor U19446 (N_19446,N_16018,N_17409);
xor U19447 (N_19447,N_17176,N_15173);
nand U19448 (N_19448,N_15281,N_15793);
or U19449 (N_19449,N_15955,N_17234);
or U19450 (N_19450,N_15797,N_15977);
nor U19451 (N_19451,N_16567,N_17428);
xor U19452 (N_19452,N_16563,N_15093);
or U19453 (N_19453,N_15760,N_16765);
or U19454 (N_19454,N_17373,N_15634);
or U19455 (N_19455,N_15522,N_15665);
nand U19456 (N_19456,N_16543,N_15486);
and U19457 (N_19457,N_15754,N_16587);
xnor U19458 (N_19458,N_15464,N_15509);
and U19459 (N_19459,N_17203,N_15059);
nor U19460 (N_19460,N_16175,N_16248);
nor U19461 (N_19461,N_15251,N_16696);
and U19462 (N_19462,N_15448,N_16141);
or U19463 (N_19463,N_15519,N_16163);
nand U19464 (N_19464,N_16827,N_17488);
nor U19465 (N_19465,N_16048,N_15478);
nor U19466 (N_19466,N_15024,N_15563);
xnor U19467 (N_19467,N_15009,N_15791);
xnor U19468 (N_19468,N_17416,N_16815);
xnor U19469 (N_19469,N_15233,N_15761);
nand U19470 (N_19470,N_15589,N_16696);
nand U19471 (N_19471,N_16147,N_16160);
and U19472 (N_19472,N_16971,N_15259);
or U19473 (N_19473,N_17337,N_15837);
or U19474 (N_19474,N_16338,N_15659);
and U19475 (N_19475,N_16168,N_16630);
or U19476 (N_19476,N_15145,N_15870);
nor U19477 (N_19477,N_17132,N_16305);
nor U19478 (N_19478,N_16778,N_16544);
and U19479 (N_19479,N_17223,N_15309);
nand U19480 (N_19480,N_16890,N_15875);
or U19481 (N_19481,N_15174,N_15883);
nand U19482 (N_19482,N_17078,N_16088);
nor U19483 (N_19483,N_16067,N_17420);
nor U19484 (N_19484,N_16311,N_16228);
nor U19485 (N_19485,N_16082,N_16100);
or U19486 (N_19486,N_15571,N_15367);
or U19487 (N_19487,N_16651,N_17005);
nor U19488 (N_19488,N_16820,N_16636);
and U19489 (N_19489,N_15094,N_17058);
nor U19490 (N_19490,N_15203,N_15304);
and U19491 (N_19491,N_15345,N_16480);
nand U19492 (N_19492,N_15071,N_17047);
nand U19493 (N_19493,N_15220,N_15241);
nand U19494 (N_19494,N_16903,N_17383);
xor U19495 (N_19495,N_16626,N_16084);
nor U19496 (N_19496,N_17338,N_16935);
nor U19497 (N_19497,N_16539,N_16281);
nor U19498 (N_19498,N_15826,N_16059);
xnor U19499 (N_19499,N_17010,N_15920);
nand U19500 (N_19500,N_16746,N_17225);
nor U19501 (N_19501,N_15698,N_16403);
nand U19502 (N_19502,N_15103,N_15991);
nor U19503 (N_19503,N_15853,N_16988);
and U19504 (N_19504,N_16430,N_16378);
nor U19505 (N_19505,N_16072,N_15111);
nor U19506 (N_19506,N_16713,N_17229);
nor U19507 (N_19507,N_15246,N_15171);
or U19508 (N_19508,N_17401,N_16777);
xnor U19509 (N_19509,N_16844,N_16176);
and U19510 (N_19510,N_16884,N_17418);
nand U19511 (N_19511,N_16208,N_17081);
or U19512 (N_19512,N_16980,N_17015);
nand U19513 (N_19513,N_15576,N_15505);
and U19514 (N_19514,N_17239,N_16579);
nand U19515 (N_19515,N_15917,N_15810);
and U19516 (N_19516,N_17269,N_15971);
nand U19517 (N_19517,N_17193,N_16575);
nand U19518 (N_19518,N_17140,N_15493);
nand U19519 (N_19519,N_16343,N_15756);
or U19520 (N_19520,N_16559,N_16101);
nand U19521 (N_19521,N_15692,N_16856);
and U19522 (N_19522,N_15677,N_16627);
and U19523 (N_19523,N_15574,N_16166);
nand U19524 (N_19524,N_16033,N_16429);
and U19525 (N_19525,N_15485,N_16069);
xnor U19526 (N_19526,N_15329,N_17018);
nor U19527 (N_19527,N_17146,N_15245);
nor U19528 (N_19528,N_17051,N_15283);
xnor U19529 (N_19529,N_16478,N_16068);
or U19530 (N_19530,N_16191,N_15490);
and U19531 (N_19531,N_16007,N_16894);
and U19532 (N_19532,N_17249,N_15232);
nand U19533 (N_19533,N_16961,N_16658);
and U19534 (N_19534,N_15403,N_15691);
and U19535 (N_19535,N_15466,N_15948);
and U19536 (N_19536,N_16592,N_16875);
nand U19537 (N_19537,N_17046,N_16010);
nor U19538 (N_19538,N_16099,N_17471);
or U19539 (N_19539,N_15229,N_15497);
and U19540 (N_19540,N_16336,N_15827);
or U19541 (N_19541,N_15154,N_17392);
xor U19542 (N_19542,N_15459,N_17104);
and U19543 (N_19543,N_17358,N_16021);
or U19544 (N_19544,N_17200,N_17110);
and U19545 (N_19545,N_16422,N_16636);
and U19546 (N_19546,N_15174,N_17162);
and U19547 (N_19547,N_16539,N_16782);
nor U19548 (N_19548,N_16930,N_17149);
and U19549 (N_19549,N_15015,N_16021);
or U19550 (N_19550,N_15047,N_16078);
nor U19551 (N_19551,N_16483,N_15825);
nor U19552 (N_19552,N_16674,N_16392);
nand U19553 (N_19553,N_16912,N_15365);
nand U19554 (N_19554,N_17037,N_17047);
nor U19555 (N_19555,N_15338,N_16868);
and U19556 (N_19556,N_15774,N_15513);
nor U19557 (N_19557,N_15802,N_15887);
nor U19558 (N_19558,N_15178,N_16756);
xnor U19559 (N_19559,N_16677,N_15935);
nor U19560 (N_19560,N_17422,N_17385);
or U19561 (N_19561,N_17477,N_15427);
or U19562 (N_19562,N_17409,N_15742);
and U19563 (N_19563,N_15827,N_15147);
xnor U19564 (N_19564,N_17098,N_15338);
nand U19565 (N_19565,N_16043,N_16947);
and U19566 (N_19566,N_16855,N_15448);
xor U19567 (N_19567,N_16412,N_17496);
nand U19568 (N_19568,N_16957,N_17369);
nand U19569 (N_19569,N_16730,N_15528);
nand U19570 (N_19570,N_15811,N_17166);
or U19571 (N_19571,N_15397,N_16942);
or U19572 (N_19572,N_16729,N_16752);
xor U19573 (N_19573,N_15048,N_16803);
nor U19574 (N_19574,N_16223,N_16893);
or U19575 (N_19575,N_17459,N_16386);
or U19576 (N_19576,N_17267,N_17492);
nand U19577 (N_19577,N_15096,N_17416);
and U19578 (N_19578,N_15920,N_16161);
and U19579 (N_19579,N_16622,N_15281);
or U19580 (N_19580,N_15266,N_15291);
and U19581 (N_19581,N_16803,N_16677);
and U19582 (N_19582,N_15792,N_15624);
and U19583 (N_19583,N_15753,N_15953);
nor U19584 (N_19584,N_17243,N_16158);
or U19585 (N_19585,N_17006,N_15672);
or U19586 (N_19586,N_16483,N_16082);
or U19587 (N_19587,N_17212,N_17389);
or U19588 (N_19588,N_15499,N_15342);
nor U19589 (N_19589,N_16526,N_16437);
nand U19590 (N_19590,N_16933,N_16793);
and U19591 (N_19591,N_15702,N_16055);
or U19592 (N_19592,N_15892,N_17232);
or U19593 (N_19593,N_15838,N_16012);
and U19594 (N_19594,N_16640,N_16495);
nor U19595 (N_19595,N_16468,N_17070);
nor U19596 (N_19596,N_16105,N_17421);
nand U19597 (N_19597,N_16256,N_16809);
nor U19598 (N_19598,N_16005,N_16109);
xnor U19599 (N_19599,N_15987,N_15825);
nand U19600 (N_19600,N_16013,N_16184);
or U19601 (N_19601,N_15733,N_15314);
nor U19602 (N_19602,N_16795,N_15107);
nand U19603 (N_19603,N_16951,N_15992);
and U19604 (N_19604,N_15903,N_15369);
nand U19605 (N_19605,N_16196,N_16028);
and U19606 (N_19606,N_17316,N_15131);
nand U19607 (N_19607,N_15551,N_15991);
or U19608 (N_19608,N_15396,N_17355);
or U19609 (N_19609,N_17197,N_17147);
or U19610 (N_19610,N_16818,N_15618);
or U19611 (N_19611,N_15051,N_16255);
and U19612 (N_19612,N_15272,N_16639);
or U19613 (N_19613,N_16274,N_16189);
or U19614 (N_19614,N_15868,N_16867);
nand U19615 (N_19615,N_16076,N_17400);
nand U19616 (N_19616,N_15421,N_17363);
or U19617 (N_19617,N_15456,N_17151);
nand U19618 (N_19618,N_15203,N_15920);
nor U19619 (N_19619,N_17148,N_15497);
nor U19620 (N_19620,N_16149,N_16510);
nand U19621 (N_19621,N_16336,N_16060);
xnor U19622 (N_19622,N_16660,N_15710);
nand U19623 (N_19623,N_16601,N_15538);
xor U19624 (N_19624,N_17018,N_16074);
and U19625 (N_19625,N_15501,N_15588);
nand U19626 (N_19626,N_17428,N_16770);
or U19627 (N_19627,N_15162,N_16706);
or U19628 (N_19628,N_16158,N_15539);
and U19629 (N_19629,N_17358,N_16226);
nand U19630 (N_19630,N_17283,N_16098);
nand U19631 (N_19631,N_15577,N_17443);
and U19632 (N_19632,N_17284,N_15759);
nand U19633 (N_19633,N_17244,N_16772);
nor U19634 (N_19634,N_15555,N_16780);
nor U19635 (N_19635,N_16518,N_16436);
nor U19636 (N_19636,N_16345,N_16110);
nand U19637 (N_19637,N_16234,N_16138);
xor U19638 (N_19638,N_15182,N_16218);
or U19639 (N_19639,N_17493,N_16517);
nand U19640 (N_19640,N_16435,N_16229);
or U19641 (N_19641,N_15926,N_15042);
or U19642 (N_19642,N_15617,N_16266);
or U19643 (N_19643,N_15915,N_15067);
nand U19644 (N_19644,N_15685,N_15416);
nand U19645 (N_19645,N_15437,N_16252);
xor U19646 (N_19646,N_15061,N_16521);
nor U19647 (N_19647,N_16480,N_15724);
nor U19648 (N_19648,N_17497,N_16087);
nand U19649 (N_19649,N_17168,N_16121);
nor U19650 (N_19650,N_15274,N_16685);
nor U19651 (N_19651,N_17174,N_16455);
and U19652 (N_19652,N_16894,N_16600);
nor U19653 (N_19653,N_16928,N_16923);
and U19654 (N_19654,N_15497,N_15203);
nor U19655 (N_19655,N_15074,N_16145);
and U19656 (N_19656,N_15246,N_16860);
nor U19657 (N_19657,N_16645,N_15129);
or U19658 (N_19658,N_15617,N_17094);
or U19659 (N_19659,N_16123,N_16259);
or U19660 (N_19660,N_15789,N_16794);
or U19661 (N_19661,N_16848,N_16825);
and U19662 (N_19662,N_15817,N_16745);
xnor U19663 (N_19663,N_15737,N_16704);
nor U19664 (N_19664,N_17225,N_16316);
nor U19665 (N_19665,N_15697,N_16802);
or U19666 (N_19666,N_17376,N_16270);
and U19667 (N_19667,N_15521,N_17141);
nand U19668 (N_19668,N_16571,N_17320);
and U19669 (N_19669,N_15677,N_17203);
and U19670 (N_19670,N_15648,N_15883);
nor U19671 (N_19671,N_16653,N_15280);
xnor U19672 (N_19672,N_15974,N_16802);
nor U19673 (N_19673,N_17060,N_16913);
or U19674 (N_19674,N_15391,N_16930);
nor U19675 (N_19675,N_15734,N_16465);
nand U19676 (N_19676,N_15700,N_16451);
and U19677 (N_19677,N_15160,N_15314);
nor U19678 (N_19678,N_15107,N_16974);
or U19679 (N_19679,N_16519,N_16372);
and U19680 (N_19680,N_17236,N_16548);
nor U19681 (N_19681,N_15494,N_17302);
or U19682 (N_19682,N_16657,N_15712);
nor U19683 (N_19683,N_16452,N_15896);
nand U19684 (N_19684,N_15834,N_15881);
or U19685 (N_19685,N_17151,N_16888);
or U19686 (N_19686,N_16617,N_15270);
and U19687 (N_19687,N_15067,N_15432);
nand U19688 (N_19688,N_15153,N_16235);
xnor U19689 (N_19689,N_16622,N_16459);
nor U19690 (N_19690,N_16626,N_16119);
nand U19691 (N_19691,N_16699,N_16285);
nor U19692 (N_19692,N_15100,N_17191);
nand U19693 (N_19693,N_16136,N_16821);
or U19694 (N_19694,N_15065,N_15918);
and U19695 (N_19695,N_15046,N_15233);
or U19696 (N_19696,N_17160,N_16827);
nor U19697 (N_19697,N_15105,N_16567);
and U19698 (N_19698,N_15284,N_16614);
xnor U19699 (N_19699,N_16930,N_15906);
nor U19700 (N_19700,N_15660,N_15693);
and U19701 (N_19701,N_15624,N_16440);
nand U19702 (N_19702,N_16385,N_16625);
nor U19703 (N_19703,N_16129,N_16831);
and U19704 (N_19704,N_17381,N_16629);
and U19705 (N_19705,N_15771,N_16054);
nor U19706 (N_19706,N_16916,N_15517);
nand U19707 (N_19707,N_17471,N_17201);
and U19708 (N_19708,N_16360,N_16344);
nand U19709 (N_19709,N_15535,N_15436);
and U19710 (N_19710,N_17093,N_16230);
and U19711 (N_19711,N_15017,N_17130);
nor U19712 (N_19712,N_16028,N_16031);
xor U19713 (N_19713,N_15576,N_16715);
and U19714 (N_19714,N_15826,N_15186);
xor U19715 (N_19715,N_17486,N_15791);
nor U19716 (N_19716,N_17461,N_16456);
nor U19717 (N_19717,N_15101,N_15514);
nand U19718 (N_19718,N_16019,N_17466);
nand U19719 (N_19719,N_15766,N_15670);
or U19720 (N_19720,N_17157,N_15948);
and U19721 (N_19721,N_15934,N_17382);
nor U19722 (N_19722,N_15663,N_15027);
or U19723 (N_19723,N_15728,N_17487);
or U19724 (N_19724,N_17493,N_16717);
or U19725 (N_19725,N_17134,N_17397);
nor U19726 (N_19726,N_16579,N_15741);
nor U19727 (N_19727,N_15989,N_16494);
nor U19728 (N_19728,N_15807,N_16520);
or U19729 (N_19729,N_15161,N_16489);
or U19730 (N_19730,N_16177,N_16312);
and U19731 (N_19731,N_16414,N_16471);
nand U19732 (N_19732,N_15520,N_16870);
or U19733 (N_19733,N_16922,N_15206);
nor U19734 (N_19734,N_16985,N_15085);
xnor U19735 (N_19735,N_15769,N_15217);
nor U19736 (N_19736,N_15290,N_15553);
and U19737 (N_19737,N_15577,N_16492);
nor U19738 (N_19738,N_15622,N_17324);
nand U19739 (N_19739,N_16875,N_15719);
nand U19740 (N_19740,N_16131,N_17184);
nand U19741 (N_19741,N_16301,N_16499);
and U19742 (N_19742,N_15761,N_16565);
or U19743 (N_19743,N_16960,N_17115);
nand U19744 (N_19744,N_15746,N_17103);
nand U19745 (N_19745,N_16879,N_16639);
or U19746 (N_19746,N_15004,N_15773);
and U19747 (N_19747,N_15441,N_15526);
and U19748 (N_19748,N_15491,N_15803);
nand U19749 (N_19749,N_15719,N_17048);
nor U19750 (N_19750,N_15669,N_15784);
nor U19751 (N_19751,N_15702,N_15075);
nand U19752 (N_19752,N_16446,N_15261);
nor U19753 (N_19753,N_16635,N_15025);
nand U19754 (N_19754,N_15612,N_16622);
and U19755 (N_19755,N_17367,N_15402);
xor U19756 (N_19756,N_15018,N_16503);
nand U19757 (N_19757,N_15635,N_15701);
nor U19758 (N_19758,N_15196,N_15189);
and U19759 (N_19759,N_15523,N_17205);
nand U19760 (N_19760,N_16570,N_15942);
or U19761 (N_19761,N_17052,N_16340);
and U19762 (N_19762,N_15511,N_16023);
nand U19763 (N_19763,N_15773,N_16544);
nand U19764 (N_19764,N_16288,N_15731);
and U19765 (N_19765,N_16362,N_16297);
nand U19766 (N_19766,N_15431,N_17210);
nor U19767 (N_19767,N_15944,N_16292);
nand U19768 (N_19768,N_15417,N_16949);
and U19769 (N_19769,N_17133,N_17497);
xnor U19770 (N_19770,N_16307,N_16908);
or U19771 (N_19771,N_17329,N_15749);
xor U19772 (N_19772,N_16922,N_16531);
and U19773 (N_19773,N_16099,N_17048);
and U19774 (N_19774,N_16890,N_16996);
or U19775 (N_19775,N_15889,N_16171);
and U19776 (N_19776,N_17438,N_16090);
nor U19777 (N_19777,N_16612,N_17282);
nand U19778 (N_19778,N_16511,N_15984);
or U19779 (N_19779,N_16226,N_17321);
or U19780 (N_19780,N_15465,N_15085);
nand U19781 (N_19781,N_15421,N_15197);
or U19782 (N_19782,N_15934,N_15672);
nand U19783 (N_19783,N_15703,N_16298);
nand U19784 (N_19784,N_15818,N_17415);
or U19785 (N_19785,N_15151,N_15227);
or U19786 (N_19786,N_15146,N_16999);
or U19787 (N_19787,N_16892,N_17052);
xnor U19788 (N_19788,N_17319,N_15227);
and U19789 (N_19789,N_16440,N_17059);
and U19790 (N_19790,N_16611,N_15761);
nand U19791 (N_19791,N_15705,N_15697);
or U19792 (N_19792,N_15200,N_16934);
nand U19793 (N_19793,N_16904,N_15511);
nand U19794 (N_19794,N_16604,N_15140);
nor U19795 (N_19795,N_17491,N_17214);
or U19796 (N_19796,N_15180,N_15271);
and U19797 (N_19797,N_17439,N_17340);
nand U19798 (N_19798,N_15644,N_16869);
nor U19799 (N_19799,N_17191,N_16219);
or U19800 (N_19800,N_17399,N_15113);
nor U19801 (N_19801,N_16086,N_15585);
and U19802 (N_19802,N_15321,N_16190);
nand U19803 (N_19803,N_15866,N_16007);
or U19804 (N_19804,N_16371,N_15269);
nand U19805 (N_19805,N_17407,N_15960);
nand U19806 (N_19806,N_17365,N_15853);
nor U19807 (N_19807,N_16633,N_15413);
nor U19808 (N_19808,N_16853,N_16003);
nand U19809 (N_19809,N_17144,N_15653);
nand U19810 (N_19810,N_17437,N_15881);
nor U19811 (N_19811,N_15202,N_17185);
and U19812 (N_19812,N_15564,N_16295);
nor U19813 (N_19813,N_17278,N_17117);
xnor U19814 (N_19814,N_16621,N_15461);
and U19815 (N_19815,N_17319,N_15925);
or U19816 (N_19816,N_15432,N_17417);
and U19817 (N_19817,N_16336,N_15090);
and U19818 (N_19818,N_17331,N_16297);
and U19819 (N_19819,N_17412,N_17217);
nand U19820 (N_19820,N_17013,N_17360);
xor U19821 (N_19821,N_15438,N_17443);
nand U19822 (N_19822,N_15791,N_15541);
or U19823 (N_19823,N_16319,N_15886);
and U19824 (N_19824,N_16750,N_17475);
or U19825 (N_19825,N_16767,N_15025);
and U19826 (N_19826,N_16610,N_17432);
and U19827 (N_19827,N_17075,N_16129);
or U19828 (N_19828,N_15483,N_15371);
nor U19829 (N_19829,N_16017,N_15429);
nor U19830 (N_19830,N_16889,N_15920);
or U19831 (N_19831,N_17104,N_15956);
xnor U19832 (N_19832,N_17307,N_15057);
nand U19833 (N_19833,N_17192,N_16246);
or U19834 (N_19834,N_16542,N_17342);
and U19835 (N_19835,N_15933,N_15003);
nand U19836 (N_19836,N_17083,N_15820);
or U19837 (N_19837,N_16733,N_15030);
and U19838 (N_19838,N_17392,N_15882);
nor U19839 (N_19839,N_17050,N_15789);
nor U19840 (N_19840,N_15570,N_16042);
nand U19841 (N_19841,N_16745,N_16965);
or U19842 (N_19842,N_16368,N_16790);
nor U19843 (N_19843,N_17302,N_17275);
and U19844 (N_19844,N_16914,N_15885);
or U19845 (N_19845,N_15924,N_16878);
or U19846 (N_19846,N_16735,N_16010);
or U19847 (N_19847,N_16001,N_15937);
nor U19848 (N_19848,N_15509,N_15570);
and U19849 (N_19849,N_15534,N_15858);
nand U19850 (N_19850,N_15747,N_16436);
nand U19851 (N_19851,N_15961,N_16081);
and U19852 (N_19852,N_15764,N_16981);
nand U19853 (N_19853,N_16308,N_15211);
nand U19854 (N_19854,N_15851,N_16307);
nand U19855 (N_19855,N_15533,N_15222);
nand U19856 (N_19856,N_15623,N_17293);
and U19857 (N_19857,N_15235,N_16468);
nor U19858 (N_19858,N_17476,N_16465);
nand U19859 (N_19859,N_17116,N_16731);
and U19860 (N_19860,N_15397,N_17148);
nor U19861 (N_19861,N_17123,N_15790);
or U19862 (N_19862,N_16021,N_16421);
and U19863 (N_19863,N_17113,N_15956);
nand U19864 (N_19864,N_15651,N_16381);
or U19865 (N_19865,N_17018,N_15734);
and U19866 (N_19866,N_16324,N_16462);
nand U19867 (N_19867,N_17066,N_16192);
nand U19868 (N_19868,N_16354,N_17370);
or U19869 (N_19869,N_16475,N_17203);
xnor U19870 (N_19870,N_17201,N_17378);
nand U19871 (N_19871,N_16159,N_15995);
and U19872 (N_19872,N_15618,N_16353);
and U19873 (N_19873,N_15204,N_15489);
and U19874 (N_19874,N_15007,N_16238);
nand U19875 (N_19875,N_15517,N_17120);
nor U19876 (N_19876,N_16512,N_16632);
nor U19877 (N_19877,N_16970,N_16115);
nand U19878 (N_19878,N_15571,N_15065);
or U19879 (N_19879,N_15695,N_15796);
or U19880 (N_19880,N_15780,N_15147);
nand U19881 (N_19881,N_16899,N_15060);
and U19882 (N_19882,N_17481,N_15717);
nor U19883 (N_19883,N_16990,N_15870);
nor U19884 (N_19884,N_17366,N_15062);
or U19885 (N_19885,N_16069,N_16154);
xor U19886 (N_19886,N_15763,N_17143);
or U19887 (N_19887,N_16583,N_17428);
and U19888 (N_19888,N_15351,N_15374);
nor U19889 (N_19889,N_15899,N_17391);
or U19890 (N_19890,N_16373,N_16988);
and U19891 (N_19891,N_17039,N_17214);
nand U19892 (N_19892,N_15022,N_17055);
or U19893 (N_19893,N_16941,N_15260);
nor U19894 (N_19894,N_15555,N_15670);
and U19895 (N_19895,N_17233,N_15251);
nand U19896 (N_19896,N_15590,N_17279);
nor U19897 (N_19897,N_16727,N_16362);
xor U19898 (N_19898,N_15183,N_15357);
nand U19899 (N_19899,N_15918,N_15219);
and U19900 (N_19900,N_15819,N_16022);
nand U19901 (N_19901,N_16330,N_15783);
nor U19902 (N_19902,N_16968,N_16846);
nor U19903 (N_19903,N_17368,N_15104);
and U19904 (N_19904,N_15204,N_15037);
and U19905 (N_19905,N_17204,N_15756);
nor U19906 (N_19906,N_17174,N_15701);
and U19907 (N_19907,N_15841,N_16236);
xnor U19908 (N_19908,N_16944,N_15195);
and U19909 (N_19909,N_15630,N_17103);
nand U19910 (N_19910,N_16801,N_16299);
or U19911 (N_19911,N_15752,N_17082);
nand U19912 (N_19912,N_15141,N_15649);
and U19913 (N_19913,N_15189,N_15305);
nor U19914 (N_19914,N_17344,N_16101);
and U19915 (N_19915,N_16484,N_16361);
and U19916 (N_19916,N_16061,N_16224);
nand U19917 (N_19917,N_15389,N_15453);
xor U19918 (N_19918,N_15952,N_16520);
nor U19919 (N_19919,N_15542,N_16791);
nor U19920 (N_19920,N_16270,N_16615);
and U19921 (N_19921,N_15267,N_17020);
nand U19922 (N_19922,N_16827,N_16070);
nor U19923 (N_19923,N_17498,N_15456);
nor U19924 (N_19924,N_16262,N_16075);
nor U19925 (N_19925,N_15022,N_15345);
or U19926 (N_19926,N_16507,N_15795);
xnor U19927 (N_19927,N_15961,N_16308);
nand U19928 (N_19928,N_15821,N_17333);
and U19929 (N_19929,N_15752,N_17189);
nand U19930 (N_19930,N_15998,N_17487);
and U19931 (N_19931,N_16797,N_17024);
nand U19932 (N_19932,N_17344,N_17436);
or U19933 (N_19933,N_15843,N_17286);
xnor U19934 (N_19934,N_16278,N_16069);
nor U19935 (N_19935,N_17168,N_15633);
nor U19936 (N_19936,N_17249,N_17095);
and U19937 (N_19937,N_16799,N_17321);
xor U19938 (N_19938,N_16936,N_17450);
and U19939 (N_19939,N_15969,N_15240);
nand U19940 (N_19940,N_16509,N_16626);
nand U19941 (N_19941,N_15621,N_16410);
nor U19942 (N_19942,N_16617,N_16522);
nand U19943 (N_19943,N_15328,N_15759);
nand U19944 (N_19944,N_16536,N_17148);
or U19945 (N_19945,N_15699,N_15714);
and U19946 (N_19946,N_16173,N_15083);
or U19947 (N_19947,N_16585,N_15076);
nand U19948 (N_19948,N_16011,N_16429);
nand U19949 (N_19949,N_16545,N_16972);
nor U19950 (N_19950,N_17467,N_15850);
or U19951 (N_19951,N_17217,N_15655);
nand U19952 (N_19952,N_16154,N_15046);
nand U19953 (N_19953,N_15149,N_15378);
or U19954 (N_19954,N_15616,N_16563);
nand U19955 (N_19955,N_17101,N_17076);
xor U19956 (N_19956,N_17110,N_15714);
nand U19957 (N_19957,N_16326,N_16639);
nor U19958 (N_19958,N_17312,N_15180);
nand U19959 (N_19959,N_16749,N_16471);
or U19960 (N_19960,N_16699,N_17210);
and U19961 (N_19961,N_15538,N_15449);
nand U19962 (N_19962,N_16963,N_17269);
and U19963 (N_19963,N_15846,N_15917);
nand U19964 (N_19964,N_16869,N_15544);
and U19965 (N_19965,N_16814,N_16116);
nand U19966 (N_19966,N_16697,N_15942);
and U19967 (N_19967,N_16990,N_17291);
xor U19968 (N_19968,N_15981,N_15465);
or U19969 (N_19969,N_16220,N_16507);
or U19970 (N_19970,N_15678,N_17430);
nor U19971 (N_19971,N_16693,N_17222);
xnor U19972 (N_19972,N_17165,N_16625);
and U19973 (N_19973,N_15738,N_16753);
and U19974 (N_19974,N_15372,N_16004);
nand U19975 (N_19975,N_16813,N_16502);
nor U19976 (N_19976,N_15693,N_17292);
nand U19977 (N_19977,N_16424,N_17340);
nor U19978 (N_19978,N_16229,N_16998);
xor U19979 (N_19979,N_15868,N_15014);
and U19980 (N_19980,N_15955,N_15092);
nand U19981 (N_19981,N_15974,N_16687);
nand U19982 (N_19982,N_15918,N_15892);
or U19983 (N_19983,N_16801,N_15099);
nor U19984 (N_19984,N_17256,N_15765);
nor U19985 (N_19985,N_16607,N_16295);
nor U19986 (N_19986,N_17282,N_16894);
xor U19987 (N_19987,N_15765,N_15617);
nor U19988 (N_19988,N_17033,N_15815);
and U19989 (N_19989,N_15364,N_16312);
nand U19990 (N_19990,N_15668,N_15976);
nand U19991 (N_19991,N_16948,N_16120);
nand U19992 (N_19992,N_15342,N_16219);
nor U19993 (N_19993,N_16701,N_15565);
nor U19994 (N_19994,N_15423,N_17319);
nor U19995 (N_19995,N_15464,N_17418);
or U19996 (N_19996,N_17179,N_15280);
and U19997 (N_19997,N_15043,N_16943);
or U19998 (N_19998,N_15115,N_16673);
and U19999 (N_19999,N_15146,N_16819);
nor U20000 (N_20000,N_19097,N_19903);
nor U20001 (N_20001,N_19309,N_19955);
xnor U20002 (N_20002,N_19360,N_18536);
nand U20003 (N_20003,N_19859,N_17690);
nand U20004 (N_20004,N_18891,N_18965);
and U20005 (N_20005,N_17915,N_19749);
nor U20006 (N_20006,N_18340,N_19145);
nor U20007 (N_20007,N_18740,N_18657);
nand U20008 (N_20008,N_19174,N_19515);
nand U20009 (N_20009,N_19448,N_18303);
or U20010 (N_20010,N_19775,N_19176);
and U20011 (N_20011,N_17591,N_19742);
nand U20012 (N_20012,N_18755,N_19525);
or U20013 (N_20013,N_19285,N_17699);
or U20014 (N_20014,N_18379,N_19855);
nor U20015 (N_20015,N_18869,N_19409);
nand U20016 (N_20016,N_19825,N_19817);
or U20017 (N_20017,N_19968,N_18830);
nand U20018 (N_20018,N_18613,N_17773);
nand U20019 (N_20019,N_19573,N_17860);
or U20020 (N_20020,N_17501,N_17571);
and U20021 (N_20021,N_19348,N_18052);
or U20022 (N_20022,N_18136,N_17570);
or U20023 (N_20023,N_17522,N_19978);
or U20024 (N_20024,N_18614,N_17696);
nand U20025 (N_20025,N_19137,N_18405);
and U20026 (N_20026,N_18535,N_19080);
nor U20027 (N_20027,N_18245,N_18234);
nor U20028 (N_20028,N_19985,N_18729);
nand U20029 (N_20029,N_19592,N_19280);
or U20030 (N_20030,N_19513,N_18364);
and U20031 (N_20031,N_17956,N_18647);
nor U20032 (N_20032,N_17708,N_19984);
nand U20033 (N_20033,N_18971,N_18999);
nand U20034 (N_20034,N_18956,N_19722);
or U20035 (N_20035,N_18476,N_17531);
nand U20036 (N_20036,N_17697,N_18734);
or U20037 (N_20037,N_18759,N_18210);
nor U20038 (N_20038,N_17864,N_19276);
or U20039 (N_20039,N_18758,N_17700);
and U20040 (N_20040,N_19271,N_19512);
nand U20041 (N_20041,N_19247,N_19188);
nand U20042 (N_20042,N_18727,N_17528);
nand U20043 (N_20043,N_17950,N_18043);
or U20044 (N_20044,N_17841,N_19996);
nand U20045 (N_20045,N_17657,N_18412);
or U20046 (N_20046,N_19673,N_19833);
nor U20047 (N_20047,N_18519,N_18514);
and U20048 (N_20048,N_19433,N_18938);
or U20049 (N_20049,N_19956,N_18120);
nand U20050 (N_20050,N_18717,N_19300);
nand U20051 (N_20051,N_19056,N_17715);
or U20052 (N_20052,N_17741,N_17590);
or U20053 (N_20053,N_17502,N_17752);
and U20054 (N_20054,N_17881,N_18014);
xnor U20055 (N_20055,N_19637,N_17782);
nor U20056 (N_20056,N_18279,N_18857);
and U20057 (N_20057,N_19766,N_18192);
nor U20058 (N_20058,N_18266,N_19190);
nand U20059 (N_20059,N_17664,N_18592);
and U20060 (N_20060,N_19149,N_17695);
nor U20061 (N_20061,N_18829,N_18724);
or U20062 (N_20062,N_18222,N_18056);
nor U20063 (N_20063,N_19158,N_19493);
nand U20064 (N_20064,N_18552,N_19320);
or U20065 (N_20065,N_18749,N_19549);
nand U20066 (N_20066,N_18472,N_17595);
nor U20067 (N_20067,N_18308,N_17930);
and U20068 (N_20068,N_18431,N_19298);
xnor U20069 (N_20069,N_18010,N_19844);
and U20070 (N_20070,N_19782,N_18282);
or U20071 (N_20071,N_19571,N_19070);
or U20072 (N_20072,N_19245,N_17945);
or U20073 (N_20073,N_17527,N_18141);
or U20074 (N_20074,N_18400,N_18917);
or U20075 (N_20075,N_19543,N_19077);
nand U20076 (N_20076,N_19769,N_18861);
and U20077 (N_20077,N_19481,N_18445);
nand U20078 (N_20078,N_18934,N_17799);
nand U20079 (N_20079,N_19356,N_19652);
nand U20080 (N_20080,N_19861,N_18809);
and U20081 (N_20081,N_19330,N_18672);
nand U20082 (N_20082,N_17928,N_18155);
and U20083 (N_20083,N_18774,N_18042);
and U20084 (N_20084,N_18211,N_19230);
nand U20085 (N_20085,N_18252,N_19404);
and U20086 (N_20086,N_18277,N_17687);
xnor U20087 (N_20087,N_19819,N_17827);
and U20088 (N_20088,N_19868,N_19754);
xnor U20089 (N_20089,N_19881,N_19971);
nor U20090 (N_20090,N_18538,N_19175);
and U20091 (N_20091,N_19304,N_18660);
and U20092 (N_20092,N_18617,N_19691);
nor U20093 (N_20093,N_18990,N_18888);
nor U20094 (N_20094,N_17854,N_18641);
nor U20095 (N_20095,N_19429,N_18508);
xnor U20096 (N_20096,N_19197,N_19504);
nand U20097 (N_20097,N_17565,N_17744);
or U20098 (N_20098,N_18452,N_19347);
nand U20099 (N_20099,N_19902,N_19048);
nand U20100 (N_20100,N_19328,N_18294);
xnor U20101 (N_20101,N_19144,N_19069);
or U20102 (N_20102,N_19969,N_17671);
or U20103 (N_20103,N_19455,N_19622);
xor U20104 (N_20104,N_17897,N_17780);
or U20105 (N_20105,N_19849,N_19936);
or U20106 (N_20106,N_17896,N_19873);
nor U20107 (N_20107,N_19026,N_18163);
nand U20108 (N_20108,N_17851,N_19887);
or U20109 (N_20109,N_19514,N_18251);
nor U20110 (N_20110,N_18102,N_19604);
nand U20111 (N_20111,N_18616,N_18725);
xnor U20112 (N_20112,N_19628,N_18807);
or U20113 (N_20113,N_18644,N_18576);
and U20114 (N_20114,N_18417,N_18559);
nand U20115 (N_20115,N_18448,N_18035);
or U20116 (N_20116,N_17966,N_18439);
and U20117 (N_20117,N_19596,N_17635);
or U20118 (N_20118,N_18183,N_18233);
or U20119 (N_20119,N_19675,N_19747);
or U20120 (N_20120,N_19142,N_19806);
and U20121 (N_20121,N_18179,N_19728);
or U20122 (N_20122,N_18298,N_19863);
nor U20123 (N_20123,N_19828,N_19439);
or U20124 (N_20124,N_18390,N_18290);
or U20125 (N_20125,N_19415,N_18314);
and U20126 (N_20126,N_19061,N_18925);
or U20127 (N_20127,N_19576,N_18894);
nor U20128 (N_20128,N_19703,N_17818);
and U20129 (N_20129,N_19520,N_18152);
and U20130 (N_20130,N_18632,N_19641);
xor U20131 (N_20131,N_18106,N_19168);
and U20132 (N_20132,N_17674,N_19349);
and U20133 (N_20133,N_19339,N_18305);
nand U20134 (N_20134,N_18387,N_19627);
and U20135 (N_20135,N_19643,N_18811);
nand U20136 (N_20136,N_19226,N_17685);
and U20137 (N_20137,N_18873,N_19361);
or U20138 (N_20138,N_19314,N_19063);
xor U20139 (N_20139,N_19021,N_18059);
or U20140 (N_20140,N_18909,N_19617);
xnor U20141 (N_20141,N_19606,N_19460);
nor U20142 (N_20142,N_19476,N_18718);
or U20143 (N_20143,N_18404,N_18663);
nor U20144 (N_20144,N_19618,N_19709);
xor U20145 (N_20145,N_19005,N_18877);
nand U20146 (N_20146,N_18478,N_17556);
nand U20147 (N_20147,N_18515,N_19425);
or U20148 (N_20148,N_18310,N_18506);
and U20149 (N_20149,N_19727,N_19423);
and U20150 (N_20150,N_19710,N_19116);
nor U20151 (N_20151,N_17888,N_19187);
or U20152 (N_20152,N_18399,N_19052);
nand U20153 (N_20153,N_18003,N_19561);
or U20154 (N_20154,N_19718,N_17990);
nand U20155 (N_20155,N_18586,N_17969);
xor U20156 (N_20156,N_19741,N_17720);
or U20157 (N_20157,N_19967,N_18895);
or U20158 (N_20158,N_19699,N_19102);
and U20159 (N_20159,N_19386,N_18064);
and U20160 (N_20160,N_19022,N_18306);
nand U20161 (N_20161,N_19426,N_18425);
nand U20162 (N_20162,N_18567,N_19060);
nor U20163 (N_20163,N_17766,N_18093);
or U20164 (N_20164,N_18849,N_19359);
nand U20165 (N_20165,N_18459,N_19225);
xnor U20166 (N_20166,N_19951,N_17820);
or U20167 (N_20167,N_18673,N_18363);
and U20168 (N_20168,N_18646,N_18777);
nor U20169 (N_20169,N_18768,N_19153);
nand U20170 (N_20170,N_18549,N_19181);
nor U20171 (N_20171,N_17762,N_19720);
and U20172 (N_20172,N_18747,N_18598);
xor U20173 (N_20173,N_17750,N_19273);
nand U20174 (N_20174,N_18422,N_19394);
nand U20175 (N_20175,N_18621,N_18767);
or U20176 (N_20176,N_18021,N_18333);
xor U20177 (N_20177,N_19882,N_18490);
nor U20178 (N_20178,N_19745,N_19018);
nand U20179 (N_20179,N_19192,N_18868);
nor U20180 (N_20180,N_18815,N_18295);
or U20181 (N_20181,N_18151,N_17588);
nand U20182 (N_20182,N_18175,N_19418);
nand U20183 (N_20183,N_19905,N_18300);
nand U20184 (N_20184,N_17584,N_18786);
or U20185 (N_20185,N_18595,N_18882);
or U20186 (N_20186,N_19680,N_18181);
or U20187 (N_20187,N_18739,N_18193);
nand U20188 (N_20188,N_17821,N_19480);
and U20189 (N_20189,N_18612,N_18369);
nand U20190 (N_20190,N_17650,N_18943);
and U20191 (N_20191,N_19874,N_17927);
nor U20192 (N_20192,N_17692,N_18413);
nor U20193 (N_20193,N_19143,N_19935);
and U20194 (N_20194,N_17646,N_19150);
nand U20195 (N_20195,N_17684,N_18113);
and U20196 (N_20196,N_18212,N_19218);
nand U20197 (N_20197,N_18671,N_19194);
nor U20198 (N_20198,N_17508,N_18982);
xor U20199 (N_20199,N_18912,N_17934);
and U20200 (N_20200,N_18121,N_19335);
and U20201 (N_20201,N_19950,N_19536);
nand U20202 (N_20202,N_18962,N_19471);
or U20203 (N_20203,N_18752,N_19161);
and U20204 (N_20204,N_18092,N_18597);
nor U20205 (N_20205,N_19364,N_18159);
nand U20206 (N_20206,N_19698,N_19575);
nand U20207 (N_20207,N_19160,N_18770);
and U20208 (N_20208,N_19039,N_19909);
nand U20209 (N_20209,N_18027,N_18127);
nor U20210 (N_20210,N_18649,N_18221);
nor U20211 (N_20211,N_19672,N_19707);
and U20212 (N_20212,N_18793,N_18633);
or U20213 (N_20213,N_17525,N_19193);
nand U20214 (N_20214,N_18931,N_18676);
nor U20215 (N_20215,N_18855,N_19095);
xor U20216 (N_20216,N_18914,N_19616);
nor U20217 (N_20217,N_17914,N_18769);
nor U20218 (N_20218,N_17797,N_18693);
xnor U20219 (N_20219,N_18823,N_19156);
or U20220 (N_20220,N_19408,N_19577);
nand U20221 (N_20221,N_17628,N_19407);
or U20222 (N_20222,N_17844,N_18382);
nor U20223 (N_20223,N_17911,N_19338);
or U20224 (N_20224,N_17737,N_19171);
nor U20225 (N_20225,N_18426,N_19926);
and U20226 (N_20226,N_18964,N_18985);
nor U20227 (N_20227,N_19282,N_18356);
and U20228 (N_20228,N_18146,N_19997);
nor U20229 (N_20229,N_18087,N_18737);
nand U20230 (N_20230,N_17811,N_18902);
and U20231 (N_20231,N_18821,N_17879);
and U20232 (N_20232,N_19841,N_18575);
nor U20233 (N_20233,N_18007,N_18098);
nand U20234 (N_20234,N_17771,N_18083);
and U20235 (N_20235,N_17778,N_19387);
nand U20236 (N_20236,N_19500,N_19484);
and U20237 (N_20237,N_18446,N_19554);
nand U20238 (N_20238,N_17748,N_18194);
nor U20239 (N_20239,N_18715,N_17763);
and U20240 (N_20240,N_18041,N_18499);
nand U20241 (N_20241,N_17970,N_18907);
nor U20242 (N_20242,N_18296,N_19995);
and U20243 (N_20243,N_19453,N_18267);
nor U20244 (N_20244,N_18634,N_18189);
nand U20245 (N_20245,N_18989,N_17603);
and U20246 (N_20246,N_19733,N_18652);
nor U20247 (N_20247,N_18883,N_17564);
or U20248 (N_20248,N_17958,N_19959);
or U20249 (N_20249,N_19659,N_19100);
nand U20250 (N_20250,N_18780,N_18698);
nand U20251 (N_20251,N_19399,N_17803);
and U20252 (N_20252,N_18284,N_19494);
nand U20253 (N_20253,N_17596,N_19261);
nor U20254 (N_20254,N_18126,N_17722);
and U20255 (N_20255,N_19334,N_18032);
nor U20256 (N_20256,N_17648,N_19810);
xnor U20257 (N_20257,N_19847,N_18153);
or U20258 (N_20258,N_18455,N_19451);
nand U20259 (N_20259,N_18498,N_19837);
nand U20260 (N_20260,N_19921,N_18254);
nor U20261 (N_20261,N_18415,N_18860);
or U20262 (N_20262,N_19786,N_19293);
and U20263 (N_20263,N_17996,N_19840);
and U20264 (N_20264,N_18385,N_18462);
nor U20265 (N_20265,N_19925,N_19008);
and U20266 (N_20266,N_18033,N_19866);
nand U20267 (N_20267,N_18795,N_17714);
xnor U20268 (N_20268,N_18929,N_18218);
nand U20269 (N_20269,N_19507,N_18642);
nand U20270 (N_20270,N_18471,N_17840);
nor U20271 (N_20271,N_18378,N_17575);
nand U20272 (N_20272,N_18858,N_19495);
and U20273 (N_20273,N_17680,N_18975);
and U20274 (N_20274,N_19384,N_17688);
nand U20275 (N_20275,N_19016,N_17772);
xor U20276 (N_20276,N_18488,N_19565);
nor U20277 (N_20277,N_18878,N_19560);
nand U20278 (N_20278,N_19353,N_17542);
nor U20279 (N_20279,N_19803,N_18450);
or U20280 (N_20280,N_18605,N_19224);
and U20281 (N_20281,N_17561,N_19006);
and U20282 (N_20282,N_18000,N_19678);
xnor U20283 (N_20283,N_19558,N_17649);
nor U20284 (N_20284,N_19167,N_17526);
nor U20285 (N_20285,N_18044,N_17909);
or U20286 (N_20286,N_19367,N_18608);
nand U20287 (N_20287,N_17701,N_17889);
nand U20288 (N_20288,N_18474,N_19875);
nand U20289 (N_20289,N_17783,N_18825);
and U20290 (N_20290,N_18738,N_17913);
or U20291 (N_20291,N_18260,N_19712);
and U20292 (N_20292,N_18827,N_17882);
nor U20293 (N_20293,N_18143,N_18338);
and U20294 (N_20294,N_17832,N_17544);
nor U20295 (N_20295,N_19067,N_19275);
nand U20296 (N_20296,N_18456,N_19258);
nand U20297 (N_20297,N_19796,N_19283);
nor U20298 (N_20298,N_18002,N_19219);
xor U20299 (N_20299,N_17619,N_18689);
nor U20300 (N_20300,N_18246,N_18224);
and U20301 (N_20301,N_17833,N_19671);
or U20302 (N_20302,N_17511,N_18540);
nand U20303 (N_20303,N_19938,N_19203);
or U20304 (N_20304,N_18216,N_19634);
nor U20305 (N_20305,N_18564,N_19465);
nor U20306 (N_20306,N_19835,N_19750);
nand U20307 (N_20307,N_17775,N_18451);
and U20308 (N_20308,N_17919,N_17899);
and U20309 (N_20309,N_18012,N_18022);
nand U20310 (N_20310,N_17558,N_17823);
nand U20311 (N_20311,N_17517,N_17757);
nand U20312 (N_20312,N_18818,N_17637);
nor U20313 (N_20313,N_17920,N_18247);
or U20314 (N_20314,N_18703,N_19834);
or U20315 (N_20315,N_18708,N_19196);
nor U20316 (N_20316,N_17634,N_19157);
nor U20317 (N_20317,N_19055,N_19785);
nand U20318 (N_20318,N_19579,N_18105);
or U20319 (N_20319,N_18761,N_17548);
nor U20320 (N_20320,N_19474,N_19567);
and U20321 (N_20321,N_18437,N_17954);
nor U20322 (N_20322,N_19035,N_19856);
nor U20323 (N_20323,N_19928,N_19207);
or U20324 (N_20324,N_18094,N_18741);
or U20325 (N_20325,N_17798,N_19839);
or U20326 (N_20326,N_18635,N_17702);
or U20327 (N_20327,N_17764,N_18289);
and U20328 (N_20328,N_18876,N_18227);
or U20329 (N_20329,N_18916,N_19411);
nand U20330 (N_20330,N_19331,N_19546);
or U20331 (N_20331,N_18966,N_17887);
and U20332 (N_20332,N_19265,N_19631);
nand U20333 (N_20333,N_18560,N_17629);
and U20334 (N_20334,N_18150,N_19030);
or U20335 (N_20335,N_18276,N_19090);
nand U20336 (N_20336,N_19570,N_19379);
nand U20337 (N_20337,N_18493,N_19539);
nand U20338 (N_20338,N_18255,N_19180);
and U20339 (N_20339,N_18073,N_19913);
nor U20340 (N_20340,N_18682,N_18637);
and U20341 (N_20341,N_18697,N_18972);
nor U20342 (N_20342,N_18037,N_17639);
and U20343 (N_20343,N_17733,N_18664);
xor U20344 (N_20344,N_18836,N_19578);
or U20345 (N_20345,N_18961,N_18360);
nor U20346 (N_20346,N_18053,N_18440);
nand U20347 (N_20347,N_18668,N_19389);
or U20348 (N_20348,N_18636,N_17658);
and U20349 (N_20349,N_18579,N_18974);
nand U20350 (N_20350,N_18323,N_18623);
nor U20351 (N_20351,N_17786,N_18223);
nor U20352 (N_20352,N_17904,N_19082);
xor U20353 (N_20353,N_19146,N_18615);
nor U20354 (N_20354,N_18551,N_19681);
xnor U20355 (N_20355,N_18449,N_19371);
and U20356 (N_20356,N_18469,N_17886);
and U20357 (N_20357,N_18963,N_19896);
or U20358 (N_20358,N_17875,N_19485);
and U20359 (N_20359,N_17532,N_19735);
and U20360 (N_20360,N_19731,N_18475);
or U20361 (N_20361,N_19942,N_19799);
nor U20362 (N_20362,N_19108,N_19450);
nand U20363 (N_20363,N_19305,N_18401);
nor U20364 (N_20364,N_18104,N_19049);
nand U20365 (N_20365,N_19041,N_19763);
nand U20366 (N_20366,N_17843,N_19398);
nand U20367 (N_20367,N_19620,N_18775);
and U20368 (N_20368,N_19303,N_18100);
and U20369 (N_20369,N_18397,N_19899);
and U20370 (N_20370,N_18928,N_19322);
nor U20371 (N_20371,N_18319,N_19534);
nand U20372 (N_20372,N_19934,N_19636);
nand U20373 (N_20373,N_18367,N_18355);
nand U20374 (N_20374,N_18979,N_18651);
or U20375 (N_20375,N_19036,N_18969);
xor U20376 (N_20376,N_17938,N_17663);
or U20377 (N_20377,N_19326,N_18908);
or U20378 (N_20378,N_17632,N_19944);
and U20379 (N_20379,N_19011,N_18373);
nor U20380 (N_20380,N_18610,N_19777);
and U20381 (N_20381,N_19732,N_18539);
xor U20382 (N_20382,N_17998,N_18197);
or U20383 (N_20383,N_19173,N_17706);
or U20384 (N_20384,N_17640,N_18144);
or U20385 (N_20385,N_17847,N_17600);
nor U20386 (N_20386,N_19169,N_19498);
nor U20387 (N_20387,N_18903,N_18005);
or U20388 (N_20388,N_19290,N_19264);
nor U20389 (N_20389,N_18072,N_19092);
and U20390 (N_20390,N_19099,N_17933);
nor U20391 (N_20391,N_18470,N_18172);
nor U20392 (N_20392,N_17725,N_19164);
or U20393 (N_20393,N_18846,N_18661);
nor U20394 (N_20394,N_17880,N_18050);
nor U20395 (N_20395,N_17900,N_18123);
nor U20396 (N_20396,N_18833,N_18765);
and U20397 (N_20397,N_19430,N_19880);
nand U20398 (N_20398,N_18428,N_18352);
nand U20399 (N_20399,N_19831,N_17952);
nand U20400 (N_20400,N_18955,N_18942);
or U20401 (N_20401,N_18871,N_17689);
and U20402 (N_20402,N_19209,N_17845);
nor U20403 (N_20403,N_18901,N_18485);
nor U20404 (N_20404,N_17946,N_18288);
and U20405 (N_20405,N_17676,N_19003);
nand U20406 (N_20406,N_19540,N_18238);
nor U20407 (N_20407,N_19235,N_18243);
nand U20408 (N_20408,N_18486,N_19396);
nor U20409 (N_20409,N_19807,N_19961);
nor U20410 (N_20410,N_17867,N_18862);
and U20411 (N_20411,N_19487,N_18864);
and U20412 (N_20412,N_18336,N_18429);
and U20413 (N_20413,N_18346,N_18513);
nor U20414 (N_20414,N_19132,N_19015);
nand U20415 (N_20415,N_19668,N_18702);
nand U20416 (N_20416,N_18923,N_19007);
and U20417 (N_20417,N_19979,N_18722);
or U20418 (N_20418,N_17559,N_17810);
and U20419 (N_20419,N_17961,N_19179);
xor U20420 (N_20420,N_17795,N_18079);
and U20421 (N_20421,N_17529,N_18958);
nand U20422 (N_20422,N_19296,N_18867);
nand U20423 (N_20423,N_19524,N_18160);
nand U20424 (N_20424,N_17739,N_17807);
nor U20425 (N_20425,N_19310,N_18244);
and U20426 (N_20426,N_17838,N_19109);
nor U20427 (N_20427,N_18483,N_19748);
or U20428 (N_20428,N_18317,N_17709);
and U20429 (N_20429,N_18640,N_18341);
or U20430 (N_20430,N_18436,N_17812);
xor U20431 (N_20431,N_19890,N_19585);
nor U20432 (N_20432,N_19992,N_19151);
nand U20433 (N_20433,N_18984,N_18489);
and U20434 (N_20434,N_18297,N_17997);
xnor U20435 (N_20435,N_17551,N_19713);
or U20436 (N_20436,N_19079,N_19526);
and U20437 (N_20437,N_17948,N_18763);
nor U20438 (N_20438,N_17866,N_18024);
nand U20439 (N_20439,N_19813,N_17618);
nor U20440 (N_20440,N_17801,N_18593);
xor U20441 (N_20441,N_18492,N_17587);
nor U20442 (N_20442,N_17652,N_19832);
nand U20443 (N_20443,N_19352,N_18957);
or U20444 (N_20444,N_17781,N_17622);
nor U20445 (N_20445,N_19093,N_19688);
nand U20446 (N_20446,N_18937,N_18344);
nor U20447 (N_20447,N_17800,N_17574);
nor U20448 (N_20448,N_18270,N_18435);
or U20449 (N_20449,N_18922,N_19045);
nand U20450 (N_20450,N_18619,N_18139);
or U20451 (N_20451,N_19004,N_18906);
nor U20452 (N_20452,N_17607,N_18720);
nor U20453 (N_20453,N_17834,N_19449);
xor U20454 (N_20454,N_19345,N_17965);
and U20455 (N_20455,N_19853,N_19288);
and U20456 (N_20456,N_18392,N_19690);
nor U20457 (N_20457,N_18563,N_17955);
or U20458 (N_20458,N_18116,N_18960);
or U20459 (N_20459,N_17894,N_17981);
nor U20460 (N_20460,N_19040,N_18528);
or U20461 (N_20461,N_17734,N_18541);
or U20462 (N_20462,N_19594,N_18692);
nand U20463 (N_20463,N_18302,N_18748);
nor U20464 (N_20464,N_17509,N_19162);
or U20465 (N_20465,N_18186,N_18932);
or U20466 (N_20466,N_19580,N_19664);
nor U20467 (N_20467,N_17560,N_18026);
nand U20468 (N_20468,N_18550,N_17850);
or U20469 (N_20469,N_19406,N_18351);
nand U20470 (N_20470,N_18719,N_18603);
nor U20471 (N_20471,N_18347,N_18119);
or U20472 (N_20472,N_17906,N_19363);
or U20473 (N_20473,N_17724,N_18068);
or U20474 (N_20474,N_18601,N_19544);
and U20475 (N_20475,N_19836,N_18841);
nand U20476 (N_20476,N_19574,N_19670);
nand U20477 (N_20477,N_17510,N_19700);
and U20478 (N_20478,N_18607,N_19708);
nor U20479 (N_20479,N_18534,N_17636);
nand U20480 (N_20480,N_17694,N_18790);
nor U20481 (N_20481,N_18688,N_18842);
and U20482 (N_20482,N_18804,N_19202);
xor U20483 (N_20483,N_19736,N_19315);
or U20484 (N_20484,N_19216,N_19469);
nand U20485 (N_20485,N_19958,N_17539);
xnor U20486 (N_20486,N_17554,N_18587);
nor U20487 (N_20487,N_18434,N_18799);
nor U20488 (N_20488,N_19010,N_18580);
nand U20489 (N_20489,N_18555,N_17633);
or U20490 (N_20490,N_19869,N_18203);
xnor U20491 (N_20491,N_17994,N_18918);
or U20492 (N_20492,N_18546,N_19597);
nor U20493 (N_20493,N_17848,N_18318);
or U20494 (N_20494,N_19329,N_17562);
and U20495 (N_20495,N_18140,N_18154);
nor U20496 (N_20496,N_18060,N_18258);
or U20497 (N_20497,N_17836,N_19467);
nor U20498 (N_20498,N_18025,N_19970);
nand U20499 (N_20499,N_19506,N_18304);
nor U20500 (N_20500,N_19630,N_18988);
nor U20501 (N_20501,N_19584,N_19083);
and U20502 (N_20502,N_19268,N_19333);
nand U20503 (N_20503,N_18854,N_18156);
nor U20504 (N_20504,N_19768,N_19737);
nor U20505 (N_20505,N_19072,N_19538);
or U20506 (N_20506,N_19692,N_19598);
and U20507 (N_20507,N_19440,N_17580);
xor U20508 (N_20508,N_19227,N_19729);
nand U20509 (N_20509,N_18309,N_18132);
nand U20510 (N_20510,N_19686,N_17730);
and U20511 (N_20511,N_19445,N_19250);
and U20512 (N_20512,N_19136,N_17767);
nor U20513 (N_20513,N_18125,N_18886);
or U20514 (N_20514,N_18710,N_19456);
or U20515 (N_20515,N_19900,N_18843);
or U20516 (N_20516,N_19809,N_19734);
and U20517 (N_20517,N_19915,N_18744);
or U20518 (N_20518,N_19871,N_19657);
or U20519 (N_20519,N_18504,N_17686);
and U20520 (N_20520,N_19980,N_18185);
nand U20521 (N_20521,N_19117,N_18473);
nand U20522 (N_20522,N_17765,N_18174);
or U20523 (N_20523,N_19390,N_17751);
nor U20524 (N_20524,N_19139,N_18695);
and U20525 (N_20525,N_18684,N_19325);
nor U20526 (N_20526,N_19037,N_18705);
nand U20527 (N_20527,N_18835,N_19308);
xnor U20528 (N_20528,N_18018,N_19421);
nand U20529 (N_20529,N_18980,N_19547);
nor U20530 (N_20530,N_19846,N_17506);
nor U20531 (N_20531,N_17568,N_18507);
nand U20532 (N_20532,N_19753,N_18265);
nor U20533 (N_20533,N_19054,N_17758);
nand U20534 (N_20534,N_19564,N_17541);
or U20535 (N_20535,N_19464,N_18533);
and U20536 (N_20536,N_19518,N_19563);
and U20537 (N_20537,N_18525,N_19756);
or U20538 (N_20538,N_18997,N_17721);
nand U20539 (N_20539,N_18466,N_19212);
nor U20540 (N_20540,N_17895,N_18118);
or U20541 (N_20541,N_19393,N_19042);
and U20542 (N_20542,N_17578,N_19344);
xnor U20543 (N_20543,N_19417,N_18381);
or U20544 (N_20544,N_18596,N_19013);
or U20545 (N_20545,N_18678,N_18165);
xor U20546 (N_20546,N_17785,N_19447);
nand U20547 (N_20547,N_17536,N_17967);
and U20548 (N_20548,N_19388,N_19463);
and U20549 (N_20549,N_17835,N_18169);
nand U20550 (N_20550,N_17514,N_19351);
or U20551 (N_20551,N_17540,N_19633);
or U20552 (N_20552,N_19666,N_17784);
or U20553 (N_20553,N_19973,N_18249);
nor U20554 (N_20554,N_17825,N_18464);
xor U20555 (N_20555,N_17853,N_18209);
or U20556 (N_20556,N_18274,N_18269);
nor U20557 (N_20557,N_18884,N_18396);
or U20558 (N_20558,N_19537,N_19208);
nand U20559 (N_20559,N_18313,N_18076);
nor U20560 (N_20560,N_17666,N_18147);
or U20561 (N_20561,N_18177,N_19808);
and U20562 (N_20562,N_18581,N_17660);
nor U20563 (N_20563,N_18572,N_18728);
and U20564 (N_20564,N_17774,N_17760);
nand U20565 (N_20565,N_17520,N_19313);
and U20566 (N_20566,N_19318,N_19215);
nand U20567 (N_20567,N_17643,N_18751);
or U20568 (N_20568,N_19989,N_18582);
nand U20569 (N_20569,N_17589,N_19274);
and U20570 (N_20570,N_19199,N_19983);
or U20571 (N_20571,N_18038,N_18813);
and U20572 (N_20572,N_18950,N_18182);
or U20573 (N_20573,N_19918,N_19665);
or U20574 (N_20574,N_19557,N_19762);
or U20575 (N_20575,N_19302,N_18020);
or U20576 (N_20576,N_19380,N_18287);
nand U20577 (N_20577,N_19530,N_18733);
nand U20578 (N_20578,N_18531,N_17805);
nor U20579 (N_20579,N_19793,N_19679);
and U20580 (N_20580,N_19883,N_17655);
xor U20581 (N_20581,N_19663,N_19764);
nor U20582 (N_20582,N_19907,N_19497);
and U20583 (N_20583,N_18897,N_19615);
or U20584 (N_20584,N_19551,N_19438);
xnor U20585 (N_20585,N_17521,N_18712);
nor U20586 (N_20586,N_17719,N_17917);
and U20587 (N_20587,N_18700,N_18518);
xnor U20588 (N_20588,N_18001,N_17705);
xor U20589 (N_20589,N_19795,N_19138);
nor U20590 (N_20590,N_17581,N_17547);
or U20591 (N_20591,N_19569,N_19301);
nor U20592 (N_20592,N_18669,N_18838);
or U20593 (N_20593,N_19319,N_19029);
nor U20594 (N_20594,N_17957,N_17908);
nor U20595 (N_20595,N_19475,N_18129);
nand U20596 (N_20596,N_17638,N_18754);
or U20597 (N_20597,N_18981,N_17505);
or U20598 (N_20598,N_18686,N_17583);
nand U20599 (N_20599,N_17662,N_17918);
and U20600 (N_20600,N_19231,N_19204);
or U20601 (N_20601,N_18913,N_19694);
nand U20602 (N_20602,N_18383,N_17516);
nand U20603 (N_20603,N_19987,N_19505);
and U20604 (N_20604,N_19249,N_19267);
or U20605 (N_20605,N_18859,N_18949);
and U20606 (N_20606,N_19112,N_18034);
nor U20607 (N_20607,N_19922,N_17626);
and U20608 (N_20608,N_19755,N_19801);
or U20609 (N_20609,N_19701,N_19977);
or U20610 (N_20610,N_17837,N_17552);
and U20611 (N_20611,N_19454,N_18784);
nor U20612 (N_20612,N_17883,N_18013);
and U20613 (N_20613,N_17761,N_19255);
or U20614 (N_20614,N_18257,N_18164);
or U20615 (N_20615,N_19542,N_18259);
or U20616 (N_20616,N_19677,N_18548);
nand U20617 (N_20617,N_18898,N_19788);
nand U20618 (N_20618,N_18558,N_18114);
nand U20619 (N_20619,N_19009,N_19241);
xnor U20620 (N_20620,N_19901,N_17631);
and U20621 (N_20621,N_19391,N_18225);
nor U20622 (N_20622,N_17592,N_19818);
or U20623 (N_20623,N_18939,N_18526);
nand U20624 (N_20624,N_19858,N_18031);
and U20625 (N_20625,N_17586,N_18643);
and U20626 (N_20626,N_19130,N_18993);
nor U20627 (N_20627,N_17576,N_18783);
nor U20628 (N_20628,N_19726,N_19076);
or U20629 (N_20629,N_18028,N_18658);
and U20630 (N_20630,N_18879,N_19046);
and U20631 (N_20631,N_19613,N_18122);
nand U20632 (N_20632,N_18736,N_17891);
nor U20633 (N_20633,N_17791,N_17831);
xor U20634 (N_20634,N_19614,N_19532);
or U20635 (N_20635,N_19403,N_17858);
nor U20636 (N_20636,N_18968,N_19297);
or U20637 (N_20637,N_19278,N_17808);
and U20638 (N_20638,N_18810,N_19533);
nor U20639 (N_20639,N_17983,N_18509);
nor U20640 (N_20640,N_18794,N_17873);
nor U20641 (N_20641,N_18250,N_19541);
or U20642 (N_20642,N_19589,N_19891);
xnor U20643 (N_20643,N_19519,N_18566);
nor U20644 (N_20644,N_18411,N_18946);
or U20645 (N_20645,N_17623,N_17726);
nand U20646 (N_20646,N_19244,N_18653);
or U20647 (N_20647,N_17665,N_19317);
nor U20648 (N_20648,N_17874,N_18766);
nand U20649 (N_20649,N_17976,N_18110);
or U20650 (N_20650,N_19781,N_19452);
or U20651 (N_20651,N_19624,N_18510);
nor U20652 (N_20652,N_19738,N_19032);
and U20653 (N_20653,N_19719,N_19797);
nand U20654 (N_20654,N_18852,N_17901);
nor U20655 (N_20655,N_18826,N_19599);
nor U20656 (N_20656,N_19307,N_19894);
or U20657 (N_20657,N_19802,N_18561);
xor U20658 (N_20658,N_19377,N_18690);
nand U20659 (N_20659,N_17617,N_18131);
nor U20660 (N_20660,N_18229,N_18286);
nor U20661 (N_20661,N_17543,N_18199);
nor U20662 (N_20662,N_19252,N_17977);
and U20663 (N_20663,N_18188,N_19912);
nor U20664 (N_20664,N_18162,N_18611);
nor U20665 (N_20665,N_17842,N_18680);
nor U20666 (N_20666,N_19327,N_19044);
nor U20667 (N_20667,N_18389,N_17546);
nor U20668 (N_20668,N_17585,N_19413);
nor U20669 (N_20669,N_18930,N_19787);
nand U20670 (N_20670,N_19517,N_17944);
and U20671 (N_20671,N_19086,N_19744);
nand U20672 (N_20672,N_17828,N_19205);
nor U20673 (N_20673,N_19826,N_17746);
or U20674 (N_20674,N_17893,N_18402);
or U20675 (N_20675,N_17611,N_19658);
or U20676 (N_20676,N_19716,N_18995);
and U20677 (N_20677,N_19213,N_19660);
nor U20678 (N_20678,N_18433,N_19845);
and U20679 (N_20679,N_19583,N_19000);
xnor U20680 (N_20680,N_17959,N_18307);
xor U20681 (N_20681,N_19172,N_19929);
and U20682 (N_20682,N_18029,N_18421);
nand U20683 (N_20683,N_18782,N_18142);
or U20684 (N_20684,N_19906,N_17512);
or U20685 (N_20685,N_18242,N_19155);
and U20686 (N_20686,N_18215,N_19640);
and U20687 (N_20687,N_18248,N_18945);
nand U20688 (N_20688,N_17939,N_18792);
nor U20689 (N_20689,N_17723,N_18554);
xnor U20690 (N_20690,N_18423,N_19886);
or U20691 (N_20691,N_19655,N_18731);
or U20692 (N_20692,N_18594,N_19251);
and U20693 (N_20693,N_18316,N_19644);
and U20694 (N_20694,N_18206,N_18384);
nand U20695 (N_20695,N_19816,N_17538);
nand U20696 (N_20696,N_19759,N_18441);
and U20697 (N_20697,N_18571,N_18732);
nor U20698 (N_20698,N_18213,N_18874);
xor U20699 (N_20699,N_18565,N_18967);
and U20700 (N_20700,N_19346,N_19201);
xor U20701 (N_20701,N_18500,N_19765);
and U20702 (N_20702,N_17868,N_18796);
and U20703 (N_20703,N_18345,N_18845);
or U20704 (N_20704,N_18128,N_19508);
and U20705 (N_20705,N_19645,N_19186);
nor U20706 (N_20706,N_18557,N_18291);
and U20707 (N_20707,N_19354,N_19689);
and U20708 (N_20708,N_17878,N_17577);
and U20709 (N_20709,N_19647,N_19098);
or U20710 (N_20710,N_18927,N_19324);
or U20711 (N_20711,N_18124,N_18687);
or U20712 (N_20712,N_19123,N_18444);
or U20713 (N_20713,N_19610,N_18926);
nand U20714 (N_20714,N_17973,N_17572);
and U20715 (N_20715,N_19410,N_17630);
or U20716 (N_20716,N_18494,N_18482);
nand U20717 (N_20717,N_18870,N_18030);
nand U20718 (N_20718,N_18602,N_17624);
xnor U20719 (N_20719,N_19740,N_17553);
nor U20720 (N_20720,N_18416,N_18933);
or U20721 (N_20721,N_18350,N_18591);
and U20722 (N_20722,N_17537,N_18487);
nand U20723 (N_20723,N_19200,N_17608);
nor U20724 (N_20724,N_19521,N_18149);
xor U20725 (N_20725,N_19917,N_18406);
nor U20726 (N_20726,N_17569,N_19277);
or U20727 (N_20727,N_19034,N_19259);
and U20728 (N_20728,N_17602,N_18201);
nor U20729 (N_20729,N_17892,N_19914);
nor U20730 (N_20730,N_19316,N_18089);
and U20731 (N_20731,N_18023,N_18443);
xnor U20732 (N_20732,N_18407,N_19587);
nor U20733 (N_20733,N_18532,N_19653);
nand U20734 (N_20734,N_17683,N_19272);
or U20735 (N_20735,N_19930,N_19422);
nor U20736 (N_20736,N_17852,N_19375);
nand U20737 (N_20737,N_18568,N_19242);
nor U20738 (N_20738,N_19395,N_19704);
or U20739 (N_20739,N_19864,N_19170);
nor U20740 (N_20740,N_17727,N_18370);
and U20741 (N_20741,N_19243,N_19870);
and U20742 (N_20742,N_17610,N_18756);
nor U20743 (N_20743,N_18685,N_18312);
nand U20744 (N_20744,N_19473,N_18730);
nor U20745 (N_20745,N_19074,N_18271);
nor U20746 (N_20746,N_17653,N_17747);
nand U20747 (N_20747,N_19489,N_18187);
nor U20748 (N_20748,N_18656,N_18590);
and U20749 (N_20749,N_19115,N_17682);
nand U20750 (N_20750,N_19378,N_18099);
nor U20751 (N_20751,N_18896,N_18970);
nor U20752 (N_20752,N_19998,N_19625);
and U20753 (N_20753,N_18716,N_19023);
and U20754 (N_20754,N_17898,N_18418);
or U20755 (N_20755,N_18872,N_19949);
and U20756 (N_20756,N_18115,N_18019);
nand U20757 (N_20757,N_18393,N_18742);
xnor U20758 (N_20758,N_18588,N_19088);
and U20759 (N_20759,N_17871,N_19877);
nor U20760 (N_20760,N_18088,N_18890);
or U20761 (N_20761,N_18239,N_18465);
or U20762 (N_20762,N_19358,N_18674);
nor U20763 (N_20763,N_18359,N_17621);
and U20764 (N_20764,N_18349,N_19994);
or U20765 (N_20765,N_19412,N_19621);
nand U20766 (N_20766,N_17862,N_19342);
nor U20767 (N_20767,N_18496,N_18683);
and U20768 (N_20768,N_19829,N_18065);
and U20769 (N_20769,N_17625,N_19369);
or U20770 (N_20770,N_18987,N_17661);
xor U20771 (N_20771,N_19051,N_19383);
or U20772 (N_20772,N_19791,N_18824);
and U20773 (N_20773,N_17902,N_19025);
xor U20774 (N_20774,N_18817,N_19178);
nor U20775 (N_20775,N_17656,N_19428);
nor U20776 (N_20776,N_18556,N_17605);
nor U20777 (N_20777,N_19020,N_19295);
or U20778 (N_20778,N_19287,N_19595);
and U20779 (N_20779,N_17856,N_19770);
and U20780 (N_20780,N_19550,N_18178);
nand U20781 (N_20781,N_19746,N_17777);
nor U20782 (N_20782,N_19084,N_19695);
and U20783 (N_20783,N_19441,N_18335);
and U20784 (N_20784,N_18348,N_18503);
nand U20785 (N_20785,N_19884,N_18573);
nor U20786 (N_20786,N_17877,N_18628);
nand U20787 (N_20787,N_17731,N_18039);
xor U20788 (N_20788,N_19966,N_19028);
and U20789 (N_20789,N_19236,N_18529);
nor U20790 (N_20790,N_17979,N_18847);
nor U20791 (N_20791,N_17668,N_18327);
nor U20792 (N_20792,N_17794,N_18226);
and U20793 (N_20793,N_18109,N_18322);
nand U20794 (N_20794,N_18797,N_19685);
or U20795 (N_20795,N_17740,N_19924);
or U20796 (N_20796,N_17792,N_18848);
xor U20797 (N_20797,N_19229,N_17941);
nor U20798 (N_20798,N_19814,N_18569);
nor U20799 (N_20799,N_18398,N_17606);
and U20800 (N_20800,N_17995,N_18424);
nor U20801 (N_20801,N_19923,N_18137);
nand U20802 (N_20802,N_19066,N_19374);
nor U20803 (N_20803,N_19073,N_18948);
or U20804 (N_20804,N_17716,N_18654);
nand U20805 (N_20805,N_17507,N_17513);
nand U20806 (N_20806,N_18263,N_19693);
nor U20807 (N_20807,N_17609,N_18228);
or U20808 (N_20808,N_17675,N_18753);
and U20809 (N_20809,N_18745,N_18017);
and U20810 (N_20810,N_19605,N_17916);
or U20811 (N_20811,N_17742,N_17770);
or U20812 (N_20812,N_18630,N_18057);
and U20813 (N_20813,N_18280,N_19611);
and U20814 (N_20814,N_18394,N_18292);
nand U20815 (N_20815,N_18167,N_19405);
nor U20816 (N_20816,N_19381,N_18011);
nor U20817 (N_20817,N_18430,N_17962);
and U20818 (N_20818,N_18706,N_19752);
or U20819 (N_20819,N_18992,N_18330);
nor U20820 (N_20820,N_19824,N_18542);
nand U20821 (N_20821,N_19669,N_18976);
or U20822 (N_20822,N_17756,N_18495);
or U20823 (N_20823,N_18709,N_17802);
nand U20824 (N_20824,N_17987,N_18924);
nand U20825 (N_20825,N_19889,N_18820);
and U20826 (N_20826,N_19081,N_17787);
nand U20827 (N_20827,N_19113,N_18543);
or U20828 (N_20828,N_19545,N_18851);
nor U20829 (N_20829,N_18816,N_18983);
and U20830 (N_20830,N_17885,N_19492);
and U20831 (N_20831,N_17829,N_19548);
xnor U20832 (N_20832,N_19152,N_17601);
xor U20833 (N_20833,N_19850,N_18195);
or U20834 (N_20834,N_19458,N_18453);
xnor U20835 (N_20835,N_18788,N_19119);
nand U20836 (N_20836,N_19047,N_19974);
nand U20837 (N_20837,N_18638,N_19401);
nor U20838 (N_20838,N_19976,N_19773);
or U20839 (N_20839,N_18048,N_17903);
nor U20840 (N_20840,N_18253,N_19125);
or U20841 (N_20841,N_17597,N_18331);
nor U20842 (N_20842,N_17703,N_18420);
nand U20843 (N_20843,N_19999,N_18704);
nand U20844 (N_20844,N_18648,N_18108);
nand U20845 (N_20845,N_18618,N_17788);
nand U20846 (N_20846,N_17670,N_18545);
xnor U20847 (N_20847,N_19851,N_19270);
or U20848 (N_20848,N_19432,N_17745);
nor U20849 (N_20849,N_18977,N_17579);
or U20850 (N_20850,N_19607,N_17816);
nor U20851 (N_20851,N_19661,N_19436);
or U20852 (N_20852,N_17989,N_19312);
nand U20853 (N_20853,N_19602,N_18457);
and U20854 (N_20854,N_19101,N_18723);
nand U20855 (N_20855,N_17776,N_18885);
and U20856 (N_20856,N_17921,N_17857);
nor U20857 (N_20857,N_18148,N_18626);
nand U20858 (N_20858,N_18502,N_18231);
nor U20859 (N_20859,N_19129,N_19248);
or U20860 (N_20860,N_17870,N_18046);
nor U20861 (N_20861,N_19148,N_17755);
nand U20862 (N_20862,N_19772,N_18477);
and U20863 (N_20863,N_18391,N_18281);
xnor U20864 (N_20864,N_18940,N_17712);
nand U20865 (N_20865,N_19159,N_19075);
and U20866 (N_20866,N_18071,N_19717);
and U20867 (N_20867,N_17713,N_19166);
nand U20868 (N_20868,N_19916,N_18537);
nor U20869 (N_20869,N_19572,N_18427);
nor U20870 (N_20870,N_19350,N_19058);
xnor U20871 (N_20871,N_17993,N_18701);
nor U20872 (N_20872,N_19446,N_18324);
and U20873 (N_20873,N_19848,N_17693);
or U20874 (N_20874,N_19911,N_18241);
or U20875 (N_20875,N_18837,N_19778);
nand U20876 (N_20876,N_19937,N_19437);
xor U20877 (N_20877,N_18078,N_19114);
nor U20878 (N_20878,N_18840,N_19012);
or U20879 (N_20879,N_19362,N_17768);
or U20880 (N_20880,N_18952,N_18776);
or U20881 (N_20881,N_19651,N_19355);
xor U20882 (N_20882,N_17884,N_19581);
and U20883 (N_20883,N_17550,N_18321);
nand U20884 (N_20884,N_17645,N_18447);
or U20885 (N_20885,N_18278,N_17796);
nand U20886 (N_20886,N_19128,N_17524);
nand U20887 (N_20887,N_19368,N_19337);
xnor U20888 (N_20888,N_19472,N_19050);
and U20889 (N_20889,N_19878,N_18915);
and U20890 (N_20890,N_18419,N_17924);
or U20891 (N_20891,N_19562,N_19804);
or U20892 (N_20892,N_19635,N_19953);
nor U20893 (N_20893,N_17819,N_18585);
nor U20894 (N_20894,N_18320,N_19126);
nand U20895 (N_20895,N_19262,N_18577);
or U20896 (N_20896,N_18196,N_18171);
nor U20897 (N_20897,N_19591,N_18522);
and U20898 (N_20898,N_17735,N_19397);
and U20899 (N_20899,N_19110,N_19443);
or U20900 (N_20900,N_17953,N_19263);
nor U20901 (N_20901,N_18625,N_19294);
or U20902 (N_20902,N_19684,N_19743);
nor U20903 (N_20903,N_19147,N_17972);
nor U20904 (N_20904,N_19365,N_18208);
xor U20905 (N_20905,N_18395,N_19656);
nand U20906 (N_20906,N_19553,N_19991);
or U20907 (N_20907,N_19254,N_19529);
and U20908 (N_20908,N_19981,N_18819);
nand U20909 (N_20909,N_17582,N_19723);
nor U20910 (N_20910,N_18166,N_18750);
and U20911 (N_20911,N_18998,N_19931);
nand U20912 (N_20912,N_18045,N_19948);
and U20913 (N_20913,N_19779,N_17651);
nor U20914 (N_20914,N_18009,N_17503);
xor U20915 (N_20915,N_19424,N_18839);
or U20916 (N_20916,N_19952,N_18040);
or U20917 (N_20917,N_19087,N_19774);
and U20918 (N_20918,N_19842,N_19879);
and U20919 (N_20919,N_18726,N_18919);
nor U20920 (N_20920,N_18055,N_17642);
and U20921 (N_20921,N_18375,N_18696);
nor U20922 (N_20922,N_17616,N_19908);
nand U20923 (N_20923,N_18670,N_17974);
nor U20924 (N_20924,N_18299,N_18757);
nor U20925 (N_20925,N_19427,N_17518);
or U20926 (N_20926,N_19523,N_19094);
or U20927 (N_20927,N_17809,N_19648);
or U20928 (N_20928,N_19642,N_19027);
nand U20929 (N_20929,N_18054,N_17813);
nor U20930 (N_20930,N_18806,N_18342);
and U20931 (N_20931,N_19033,N_19590);
or U20932 (N_20932,N_19392,N_19867);
nor U20933 (N_20933,N_18589,N_19414);
and U20934 (N_20934,N_19586,N_18337);
xnor U20935 (N_20935,N_18236,N_19237);
or U20936 (N_20936,N_19556,N_17968);
xor U20937 (N_20937,N_18951,N_18074);
and U20938 (N_20938,N_19852,N_18666);
or U20939 (N_20939,N_18329,N_18530);
or U20940 (N_20940,N_18762,N_18480);
or U20941 (N_20941,N_18578,N_18230);
nor U20942 (N_20942,N_17641,N_18574);
and U20943 (N_20943,N_18772,N_19478);
and U20944 (N_20944,N_18235,N_19528);
nor U20945 (N_20945,N_19191,N_18662);
or U20946 (N_20946,N_18714,N_17985);
or U20947 (N_20947,N_18272,N_17963);
nor U20948 (N_20948,N_18361,N_18366);
nand U20949 (N_20949,N_17718,N_18374);
or U20950 (N_20950,N_19057,N_18834);
and U20951 (N_20951,N_19141,N_18432);
xnor U20952 (N_20952,N_19163,N_17949);
and U20953 (N_20953,N_19662,N_19739);
nor U20954 (N_20954,N_19758,N_17566);
nand U20955 (N_20955,N_17815,N_19821);
xor U20956 (N_20956,N_18198,N_18803);
nor U20957 (N_20957,N_18107,N_18112);
xor U20958 (N_20958,N_17717,N_19706);
and U20959 (N_20959,N_18831,N_18624);
nand U20960 (N_20960,N_18675,N_18491);
nor U20961 (N_20961,N_19014,N_18372);
and U20962 (N_20962,N_18328,N_18047);
xor U20963 (N_20963,N_18067,N_18629);
nor U20964 (N_20964,N_19096,N_18881);
and U20965 (N_20965,N_19131,N_17704);
nand U20966 (N_20966,N_18785,N_18639);
or U20967 (N_20967,N_17644,N_18944);
nand U20968 (N_20968,N_19711,N_18386);
nand U20969 (N_20969,N_17991,N_18764);
nor U20970 (N_20970,N_19214,N_19933);
nor U20971 (N_20971,N_19975,N_18544);
nand U20972 (N_20972,N_19111,N_18899);
nand U20973 (N_20973,N_18268,N_19206);
and U20974 (N_20974,N_19822,N_17573);
nand U20975 (N_20975,N_17988,N_18905);
and U20976 (N_20976,N_18315,N_18454);
or U20977 (N_20977,N_19400,N_18667);
or U20978 (N_20978,N_18133,N_19794);
nand U20979 (N_20979,N_19827,N_19402);
nand U20980 (N_20980,N_19457,N_18645);
and U20981 (N_20981,N_17754,N_19857);
and U20982 (N_20982,N_18161,N_18458);
nand U20983 (N_20983,N_18547,N_19127);
nand U20984 (N_20984,N_19140,N_17937);
or U20985 (N_20985,N_18015,N_18735);
nor U20986 (N_20986,N_19246,N_19820);
nor U20987 (N_20987,N_18058,N_17620);
and U20988 (N_20988,N_17743,N_19601);
and U20989 (N_20989,N_18081,N_18828);
nor U20990 (N_20990,N_18583,N_19089);
xor U20991 (N_20991,N_18665,N_18061);
nand U20992 (N_20992,N_19751,N_19284);
and U20993 (N_20993,N_18217,N_18679);
xor U20994 (N_20994,N_19919,N_19222);
or U20995 (N_20995,N_19893,N_17980);
nor U20996 (N_20996,N_19600,N_18214);
or U20997 (N_20997,N_19001,N_18911);
or U20998 (N_20998,N_18219,N_19470);
nand U20999 (N_20999,N_17971,N_19503);
nor U21000 (N_21000,N_18677,N_19420);
nor U21001 (N_21001,N_17711,N_18953);
or U21002 (N_21002,N_17677,N_18791);
or U21003 (N_21003,N_18517,N_17523);
nor U21004 (N_21004,N_19972,N_18787);
and U21005 (N_21005,N_19434,N_17984);
nor U21006 (N_21006,N_17861,N_18332);
nor U21007 (N_21007,N_19134,N_18371);
nor U21008 (N_21008,N_18262,N_19960);
nor U21009 (N_21009,N_19502,N_18004);
nand U21010 (N_21010,N_19466,N_18524);
and U21011 (N_21011,N_19963,N_18135);
nor U21012 (N_21012,N_19555,N_17549);
and U21013 (N_21013,N_18256,N_18184);
and U21014 (N_21014,N_18410,N_19531);
nand U21015 (N_21015,N_19725,N_17922);
nor U21016 (N_21016,N_18954,N_17667);
xnor U21017 (N_21017,N_17839,N_17931);
nor U21018 (N_21018,N_17698,N_19510);
xor U21019 (N_21019,N_18176,N_18293);
and U21020 (N_21020,N_18283,N_17849);
and U21021 (N_21021,N_18947,N_19609);
nand U21022 (N_21022,N_19183,N_18362);
nand U21023 (N_21023,N_17691,N_18880);
and U21024 (N_21024,N_19509,N_19062);
nor U21025 (N_21025,N_19291,N_19461);
nor U21026 (N_21026,N_18631,N_18063);
and U21027 (N_21027,N_17599,N_17830);
nand U21028 (N_21028,N_18168,N_19721);
nand U21029 (N_21029,N_17515,N_18959);
nand U21030 (N_21030,N_18365,N_19522);
or U21031 (N_21031,N_18138,N_18204);
nand U21032 (N_21032,N_19416,N_18357);
nor U21033 (N_21033,N_18994,N_17659);
or U21034 (N_21034,N_19639,N_18111);
nand U21035 (N_21035,N_17504,N_17647);
xor U21036 (N_21036,N_18802,N_19311);
nand U21037 (N_21037,N_19431,N_19185);
nor U21038 (N_21038,N_18805,N_18096);
nand U21039 (N_21039,N_19910,N_19286);
nand U21040 (N_21040,N_17779,N_19527);
xor U21041 (N_21041,N_17729,N_17563);
nand U21042 (N_21042,N_19442,N_17804);
nand U21043 (N_21043,N_17555,N_19357);
xnor U21044 (N_21044,N_19107,N_19988);
and U21045 (N_21045,N_18066,N_18822);
or U21046 (N_21046,N_17593,N_19823);
nand U21047 (N_21047,N_17846,N_18264);
nand U21048 (N_21048,N_17872,N_18200);
nand U21049 (N_21049,N_19468,N_17960);
nand U21050 (N_21050,N_17817,N_19376);
nand U21051 (N_21051,N_19696,N_19784);
or U21052 (N_21052,N_18986,N_18521);
and U21053 (N_21053,N_19702,N_17910);
or U21054 (N_21054,N_18844,N_19830);
or U21055 (N_21055,N_18694,N_19233);
nand U21056 (N_21056,N_19805,N_17942);
nor U21057 (N_21057,N_19940,N_18261);
nor U21058 (N_21058,N_18442,N_17964);
nand U21059 (N_21059,N_18460,N_18527);
nand U21060 (N_21060,N_18285,N_18889);
or U21061 (N_21061,N_19306,N_18438);
nor U21062 (N_21062,N_18097,N_19260);
xor U21063 (N_21063,N_19730,N_19120);
xnor U21064 (N_21064,N_18376,N_17926);
and U21065 (N_21065,N_19238,N_18377);
nand U21066 (N_21066,N_18921,N_18505);
and U21067 (N_21067,N_19954,N_17863);
xor U21068 (N_21068,N_19993,N_18865);
nand U21069 (N_21069,N_17793,N_19121);
or U21070 (N_21070,N_18086,N_19124);
nor U21071 (N_21071,N_19341,N_17594);
or U21072 (N_21072,N_17982,N_19511);
nor U21073 (N_21073,N_18380,N_18584);
nand U21074 (N_21074,N_18077,N_18358);
nand U21075 (N_21075,N_17999,N_18006);
or U21076 (N_21076,N_19444,N_19122);
or U21077 (N_21077,N_19945,N_18409);
xnor U21078 (N_21078,N_18622,N_17869);
nor U21079 (N_21079,N_19221,N_19626);
or U21080 (N_21080,N_19957,N_19568);
and U21081 (N_21081,N_18343,N_19279);
nand U21082 (N_21082,N_19177,N_17673);
xnor U21083 (N_21083,N_19812,N_19697);
and U21084 (N_21084,N_17947,N_19608);
xor U21085 (N_21085,N_19986,N_18892);
nor U21086 (N_21086,N_18085,N_19053);
xnor U21087 (N_21087,N_17936,N_19340);
nand U21088 (N_21088,N_18900,N_18743);
nand U21089 (N_21089,N_18339,N_18620);
and U21090 (N_21090,N_19516,N_19854);
nor U21091 (N_21091,N_17534,N_17912);
or U21092 (N_21092,N_18850,N_17669);
nor U21093 (N_21093,N_18778,N_19789);
nand U21094 (N_21094,N_17790,N_18501);
or U21095 (N_21095,N_19593,N_18084);
nand U21096 (N_21096,N_19705,N_18463);
and U21097 (N_21097,N_17932,N_17753);
or U21098 (N_21098,N_19490,N_18008);
or U21099 (N_21099,N_18650,N_18134);
nand U21100 (N_21100,N_19895,N_19281);
xnor U21101 (N_21101,N_18190,N_18101);
xnor U21102 (N_21102,N_18655,N_19002);
and U21103 (N_21103,N_18095,N_19862);
and U21104 (N_21104,N_17978,N_17749);
or U21105 (N_21105,N_19990,N_19483);
nor U21106 (N_21106,N_17925,N_19031);
or U21107 (N_21107,N_17992,N_18516);
or U21108 (N_21108,N_19619,N_19195);
or U21109 (N_21109,N_18205,N_19501);
nand U21110 (N_21110,N_18941,N_19582);
nor U21111 (N_21111,N_19435,N_17814);
nand U21112 (N_21112,N_19217,N_18553);
nand U21113 (N_21113,N_19920,N_19240);
xnor U21114 (N_21114,N_19078,N_19479);
and U21115 (N_21115,N_17935,N_19232);
and U21116 (N_21116,N_19059,N_18691);
nor U21117 (N_21117,N_19024,N_19650);
nand U21118 (N_21118,N_19373,N_17806);
nand U21119 (N_21119,N_17789,N_19800);
or U21120 (N_21120,N_19269,N_19043);
nor U21121 (N_21121,N_19499,N_19947);
xnor U21122 (N_21122,N_18808,N_19682);
nor U21123 (N_21123,N_18713,N_17865);
xor U21124 (N_21124,N_19962,N_18479);
nand U21125 (N_21125,N_19876,N_17533);
nand U21126 (N_21126,N_17557,N_19792);
and U21127 (N_21127,N_18388,N_18062);
xnor U21128 (N_21128,N_18798,N_19811);
nor U21129 (N_21129,N_18863,N_18887);
or U21130 (N_21130,N_18080,N_19676);
or U21131 (N_21131,N_17654,N_18158);
nand U21132 (N_21132,N_19496,N_18570);
nor U21133 (N_21133,N_18103,N_18275);
nor U21134 (N_21134,N_18232,N_19674);
nand U21135 (N_21135,N_18414,N_19488);
nor U21136 (N_21136,N_19336,N_18814);
or U21137 (N_21137,N_18202,N_18403);
nor U21138 (N_21138,N_17929,N_19106);
and U21139 (N_21139,N_19683,N_17822);
nand U21140 (N_21140,N_18523,N_18910);
xor U21141 (N_21141,N_18812,N_19228);
and U21142 (N_21142,N_18627,N_19790);
nor U21143 (N_21143,N_19623,N_19552);
or U21144 (N_21144,N_19761,N_18049);
or U21145 (N_21145,N_17876,N_19239);
nand U21146 (N_21146,N_18481,N_17615);
nor U21147 (N_21147,N_19182,N_19798);
and U21148 (N_21148,N_18604,N_19071);
nor U21149 (N_21149,N_19927,N_18353);
nor U21150 (N_21150,N_17598,N_18904);
nor U21151 (N_21151,N_19482,N_19189);
nand U21152 (N_21152,N_19964,N_18368);
nor U21153 (N_21153,N_18157,N_17707);
or U21154 (N_21154,N_19654,N_18760);
nor U21155 (N_21155,N_19198,N_18273);
nor U21156 (N_21156,N_19323,N_17826);
or U21157 (N_21157,N_19366,N_17769);
and U21158 (N_21158,N_19588,N_19982);
nor U21159 (N_21159,N_17951,N_19632);
nor U21160 (N_21160,N_19477,N_18781);
xor U21161 (N_21161,N_19815,N_19370);
nor U21162 (N_21162,N_19667,N_18773);
nand U21163 (N_21163,N_19133,N_17612);
nand U21164 (N_21164,N_19687,N_19118);
or U21165 (N_21165,N_19776,N_19838);
nand U21166 (N_21166,N_17567,N_18800);
nand U21167 (N_21167,N_17923,N_18497);
or U21168 (N_21168,N_18354,N_19105);
nor U21169 (N_21169,N_17535,N_17890);
xor U21170 (N_21170,N_19603,N_17728);
xor U21171 (N_21171,N_19382,N_18075);
nand U21172 (N_21172,N_17678,N_18600);
and U21173 (N_21173,N_19939,N_17986);
and U21174 (N_21174,N_18746,N_19885);
or U21175 (N_21175,N_17855,N_19566);
or U21176 (N_21176,N_18016,N_19289);
or U21177 (N_21177,N_18511,N_19299);
nor U21178 (N_21178,N_18082,N_18681);
nor U21179 (N_21179,N_19649,N_18920);
nor U21180 (N_21180,N_18220,N_19211);
nand U21181 (N_21181,N_19135,N_18484);
nor U21182 (N_21182,N_19019,N_19419);
nor U21183 (N_21183,N_19385,N_19860);
xnor U21184 (N_21184,N_18721,N_19559);
and U21185 (N_21185,N_18207,N_18117);
nor U21186 (N_21186,N_18978,N_18771);
nor U21187 (N_21187,N_18801,N_19064);
and U21188 (N_21188,N_19068,N_17681);
or U21189 (N_21189,N_18091,N_18520);
xor U21190 (N_21190,N_19904,N_17975);
nor U21191 (N_21191,N_19256,N_19462);
or U21192 (N_21192,N_18973,N_18145);
nor U21193 (N_21193,N_18935,N_19154);
xnor U21194 (N_21194,N_17613,N_18325);
and U21195 (N_21195,N_19757,N_19165);
xor U21196 (N_21196,N_19897,N_17824);
nor U21197 (N_21197,N_19943,N_19321);
or U21198 (N_21198,N_18853,N_18408);
nor U21199 (N_21199,N_19535,N_19760);
or U21200 (N_21200,N_17545,N_18996);
nand U21201 (N_21201,N_18609,N_19266);
and U21202 (N_21202,N_18237,N_17530);
nand U21203 (N_21203,N_19103,N_17627);
xor U21204 (N_21204,N_18240,N_19783);
or U21205 (N_21205,N_19085,N_17738);
or U21206 (N_21206,N_17679,N_18180);
and U21207 (N_21207,N_19932,N_18461);
and U21208 (N_21208,N_17710,N_18789);
or U21209 (N_21209,N_19459,N_19941);
nand U21210 (N_21210,N_19888,N_17500);
nand U21211 (N_21211,N_19332,N_19104);
nand U21212 (N_21212,N_19715,N_19843);
nand U21213 (N_21213,N_19065,N_18779);
and U21214 (N_21214,N_18173,N_17907);
nor U21215 (N_21215,N_17672,N_19486);
or U21216 (N_21216,N_18659,N_19038);
or U21217 (N_21217,N_18856,N_17759);
nand U21218 (N_21218,N_18301,N_18599);
or U21219 (N_21219,N_18090,N_18334);
or U21220 (N_21220,N_18467,N_18936);
xor U21221 (N_21221,N_19491,N_19184);
or U21222 (N_21222,N_18991,N_19646);
nand U21223 (N_21223,N_18893,N_19767);
xnor U21224 (N_21224,N_18875,N_19892);
nand U21225 (N_21225,N_19629,N_18170);
nand U21226 (N_21226,N_17732,N_17736);
nor U21227 (N_21227,N_18711,N_19017);
or U21228 (N_21228,N_17519,N_18070);
and U21229 (N_21229,N_18036,N_18051);
xnor U21230 (N_21230,N_18326,N_18512);
nor U21231 (N_21231,N_19946,N_18866);
nand U21232 (N_21232,N_17604,N_18311);
nand U21233 (N_21233,N_17905,N_18069);
and U21234 (N_21234,N_19223,N_19234);
or U21235 (N_21235,N_19965,N_19220);
nand U21236 (N_21236,N_19210,N_19780);
xnor U21237 (N_21237,N_19372,N_19612);
nand U21238 (N_21238,N_18699,N_19257);
or U21239 (N_21239,N_17943,N_18562);
nand U21240 (N_21240,N_17859,N_18707);
nor U21241 (N_21241,N_18130,N_18468);
nor U21242 (N_21242,N_17940,N_19771);
and U21243 (N_21243,N_19253,N_18832);
and U21244 (N_21244,N_17614,N_18191);
nand U21245 (N_21245,N_19638,N_18606);
and U21246 (N_21246,N_19292,N_19724);
and U21247 (N_21247,N_19865,N_19872);
or U21248 (N_21248,N_19898,N_19714);
and U21249 (N_21249,N_19091,N_19343);
nor U21250 (N_21250,N_19665,N_17640);
or U21251 (N_21251,N_18033,N_18973);
nor U21252 (N_21252,N_17977,N_19259);
nor U21253 (N_21253,N_17924,N_19453);
nand U21254 (N_21254,N_17795,N_17994);
nor U21255 (N_21255,N_17978,N_18238);
nand U21256 (N_21256,N_18237,N_19271);
xnor U21257 (N_21257,N_18600,N_18872);
or U21258 (N_21258,N_19346,N_18965);
and U21259 (N_21259,N_17509,N_19694);
xor U21260 (N_21260,N_19654,N_19732);
and U21261 (N_21261,N_19656,N_17883);
and U21262 (N_21262,N_17763,N_17917);
nand U21263 (N_21263,N_19639,N_18289);
and U21264 (N_21264,N_18934,N_17773);
or U21265 (N_21265,N_17908,N_19286);
xor U21266 (N_21266,N_17671,N_19009);
nand U21267 (N_21267,N_18046,N_18159);
nor U21268 (N_21268,N_18207,N_18555);
nand U21269 (N_21269,N_17914,N_18591);
nor U21270 (N_21270,N_19813,N_18554);
and U21271 (N_21271,N_18576,N_17853);
and U21272 (N_21272,N_18383,N_19999);
or U21273 (N_21273,N_18498,N_17922);
nand U21274 (N_21274,N_19647,N_19007);
and U21275 (N_21275,N_18499,N_19200);
nand U21276 (N_21276,N_19378,N_19905);
and U21277 (N_21277,N_19178,N_18415);
and U21278 (N_21278,N_17500,N_18556);
nand U21279 (N_21279,N_18559,N_19806);
or U21280 (N_21280,N_19820,N_18667);
or U21281 (N_21281,N_18993,N_19340);
nand U21282 (N_21282,N_19004,N_18837);
nor U21283 (N_21283,N_17501,N_19469);
nor U21284 (N_21284,N_17979,N_17693);
nor U21285 (N_21285,N_19736,N_17848);
nand U21286 (N_21286,N_18629,N_18078);
nor U21287 (N_21287,N_17744,N_19144);
or U21288 (N_21288,N_17995,N_17654);
and U21289 (N_21289,N_18506,N_18014);
and U21290 (N_21290,N_19799,N_19413);
nand U21291 (N_21291,N_19493,N_18619);
or U21292 (N_21292,N_18424,N_17700);
and U21293 (N_21293,N_18950,N_19822);
xor U21294 (N_21294,N_17885,N_19023);
and U21295 (N_21295,N_19335,N_17707);
and U21296 (N_21296,N_19759,N_19521);
and U21297 (N_21297,N_18054,N_18568);
and U21298 (N_21298,N_19519,N_18451);
and U21299 (N_21299,N_18417,N_18838);
or U21300 (N_21300,N_17747,N_19871);
nor U21301 (N_21301,N_18839,N_19201);
xnor U21302 (N_21302,N_18240,N_19795);
and U21303 (N_21303,N_19701,N_17935);
or U21304 (N_21304,N_18605,N_19532);
and U21305 (N_21305,N_19624,N_19952);
or U21306 (N_21306,N_18227,N_18825);
and U21307 (N_21307,N_19594,N_18162);
or U21308 (N_21308,N_18095,N_19057);
or U21309 (N_21309,N_19967,N_19396);
nor U21310 (N_21310,N_19765,N_18092);
or U21311 (N_21311,N_18328,N_18789);
nor U21312 (N_21312,N_18588,N_17984);
nor U21313 (N_21313,N_19200,N_18285);
nor U21314 (N_21314,N_19521,N_18230);
or U21315 (N_21315,N_19457,N_19589);
nand U21316 (N_21316,N_19052,N_18778);
or U21317 (N_21317,N_19164,N_18119);
nor U21318 (N_21318,N_18512,N_17607);
nor U21319 (N_21319,N_18849,N_17958);
nor U21320 (N_21320,N_19367,N_19504);
nor U21321 (N_21321,N_17668,N_19963);
and U21322 (N_21322,N_19436,N_17797);
xnor U21323 (N_21323,N_18110,N_18302);
nand U21324 (N_21324,N_19896,N_19267);
nor U21325 (N_21325,N_18436,N_19320);
or U21326 (N_21326,N_19271,N_19903);
nor U21327 (N_21327,N_19451,N_18022);
nor U21328 (N_21328,N_17959,N_17764);
xor U21329 (N_21329,N_18163,N_18369);
or U21330 (N_21330,N_19713,N_18651);
and U21331 (N_21331,N_19874,N_18275);
nor U21332 (N_21332,N_18949,N_19738);
nand U21333 (N_21333,N_17536,N_19245);
or U21334 (N_21334,N_19709,N_18328);
xor U21335 (N_21335,N_18087,N_17753);
nand U21336 (N_21336,N_17592,N_19647);
xnor U21337 (N_21337,N_18997,N_19467);
xor U21338 (N_21338,N_18211,N_18639);
nor U21339 (N_21339,N_19560,N_18070);
nor U21340 (N_21340,N_18726,N_18909);
or U21341 (N_21341,N_17832,N_18642);
nand U21342 (N_21342,N_18957,N_18936);
and U21343 (N_21343,N_17843,N_19381);
nand U21344 (N_21344,N_17893,N_19117);
nor U21345 (N_21345,N_19656,N_19559);
nor U21346 (N_21346,N_19376,N_19784);
nand U21347 (N_21347,N_17945,N_18529);
or U21348 (N_21348,N_18074,N_18369);
nor U21349 (N_21349,N_19813,N_18101);
nor U21350 (N_21350,N_18884,N_19756);
nor U21351 (N_21351,N_19719,N_19788);
nor U21352 (N_21352,N_18646,N_19343);
nand U21353 (N_21353,N_18690,N_19510);
nand U21354 (N_21354,N_18145,N_19091);
nor U21355 (N_21355,N_19884,N_19017);
nand U21356 (N_21356,N_18870,N_17616);
and U21357 (N_21357,N_18391,N_18462);
and U21358 (N_21358,N_19280,N_18633);
and U21359 (N_21359,N_17956,N_17580);
and U21360 (N_21360,N_18323,N_17888);
or U21361 (N_21361,N_19325,N_18904);
nand U21362 (N_21362,N_17627,N_19577);
nand U21363 (N_21363,N_19295,N_18158);
and U21364 (N_21364,N_19585,N_19857);
nor U21365 (N_21365,N_18069,N_18495);
xnor U21366 (N_21366,N_17738,N_19154);
or U21367 (N_21367,N_19739,N_18330);
nor U21368 (N_21368,N_17933,N_18094);
nor U21369 (N_21369,N_17622,N_19764);
or U21370 (N_21370,N_19693,N_19878);
or U21371 (N_21371,N_19560,N_19051);
and U21372 (N_21372,N_19005,N_17502);
and U21373 (N_21373,N_19236,N_17868);
nand U21374 (N_21374,N_18082,N_18378);
or U21375 (N_21375,N_19716,N_18526);
or U21376 (N_21376,N_19826,N_19677);
or U21377 (N_21377,N_19461,N_17785);
xor U21378 (N_21378,N_17950,N_19183);
or U21379 (N_21379,N_18662,N_19578);
and U21380 (N_21380,N_19831,N_19219);
or U21381 (N_21381,N_19043,N_17958);
nand U21382 (N_21382,N_18445,N_19052);
and U21383 (N_21383,N_19307,N_17707);
nor U21384 (N_21384,N_18873,N_19617);
nand U21385 (N_21385,N_19398,N_18782);
nor U21386 (N_21386,N_18503,N_18219);
nand U21387 (N_21387,N_18817,N_17675);
nor U21388 (N_21388,N_19347,N_18279);
nor U21389 (N_21389,N_19584,N_19964);
nand U21390 (N_21390,N_17717,N_18219);
xor U21391 (N_21391,N_19589,N_19557);
and U21392 (N_21392,N_19880,N_18048);
nand U21393 (N_21393,N_19967,N_18275);
nor U21394 (N_21394,N_18781,N_17651);
nor U21395 (N_21395,N_19302,N_19911);
nor U21396 (N_21396,N_17890,N_18019);
or U21397 (N_21397,N_18567,N_19792);
and U21398 (N_21398,N_19466,N_18237);
and U21399 (N_21399,N_18097,N_17952);
and U21400 (N_21400,N_19042,N_17797);
and U21401 (N_21401,N_18627,N_18854);
nand U21402 (N_21402,N_18493,N_19786);
nor U21403 (N_21403,N_19637,N_19392);
and U21404 (N_21404,N_18652,N_17962);
and U21405 (N_21405,N_17959,N_18860);
nand U21406 (N_21406,N_18170,N_19462);
and U21407 (N_21407,N_18546,N_18521);
nor U21408 (N_21408,N_18287,N_18058);
nor U21409 (N_21409,N_19273,N_19338);
and U21410 (N_21410,N_18831,N_19678);
or U21411 (N_21411,N_19811,N_18172);
or U21412 (N_21412,N_18547,N_18244);
nor U21413 (N_21413,N_18839,N_19598);
nor U21414 (N_21414,N_19487,N_17515);
xor U21415 (N_21415,N_19733,N_18073);
or U21416 (N_21416,N_19345,N_18443);
xnor U21417 (N_21417,N_18271,N_18884);
xnor U21418 (N_21418,N_19333,N_19042);
and U21419 (N_21419,N_18935,N_17844);
nand U21420 (N_21420,N_18690,N_19248);
xnor U21421 (N_21421,N_18146,N_18572);
nor U21422 (N_21422,N_19651,N_18907);
and U21423 (N_21423,N_17884,N_18151);
nor U21424 (N_21424,N_19575,N_18467);
and U21425 (N_21425,N_18213,N_18412);
and U21426 (N_21426,N_18981,N_18172);
and U21427 (N_21427,N_19000,N_19145);
or U21428 (N_21428,N_19034,N_18556);
and U21429 (N_21429,N_17777,N_19404);
nor U21430 (N_21430,N_19233,N_19802);
nor U21431 (N_21431,N_17501,N_18958);
nor U21432 (N_21432,N_19583,N_17966);
nand U21433 (N_21433,N_18530,N_18973);
nor U21434 (N_21434,N_17992,N_17516);
nand U21435 (N_21435,N_19545,N_19226);
or U21436 (N_21436,N_19930,N_17684);
and U21437 (N_21437,N_19457,N_18605);
and U21438 (N_21438,N_18734,N_18704);
or U21439 (N_21439,N_18630,N_17721);
and U21440 (N_21440,N_19366,N_18511);
nand U21441 (N_21441,N_17812,N_19288);
nor U21442 (N_21442,N_18622,N_17567);
nor U21443 (N_21443,N_19151,N_18937);
nand U21444 (N_21444,N_18758,N_19548);
and U21445 (N_21445,N_18360,N_19751);
nor U21446 (N_21446,N_18272,N_17961);
and U21447 (N_21447,N_18291,N_17758);
nand U21448 (N_21448,N_18482,N_19508);
or U21449 (N_21449,N_19336,N_18491);
nor U21450 (N_21450,N_19611,N_19303);
and U21451 (N_21451,N_19659,N_19750);
nor U21452 (N_21452,N_18922,N_17743);
nor U21453 (N_21453,N_19487,N_19137);
or U21454 (N_21454,N_19028,N_17518);
nand U21455 (N_21455,N_18268,N_18131);
nor U21456 (N_21456,N_18569,N_18334);
and U21457 (N_21457,N_19349,N_18018);
or U21458 (N_21458,N_19957,N_18293);
nor U21459 (N_21459,N_19670,N_18406);
nor U21460 (N_21460,N_18732,N_18873);
xor U21461 (N_21461,N_17506,N_17812);
nand U21462 (N_21462,N_19506,N_17966);
and U21463 (N_21463,N_19416,N_18619);
nand U21464 (N_21464,N_18490,N_19496);
nand U21465 (N_21465,N_18339,N_19957);
nor U21466 (N_21466,N_19183,N_19886);
nand U21467 (N_21467,N_19636,N_18837);
nand U21468 (N_21468,N_18836,N_19408);
nor U21469 (N_21469,N_19087,N_19572);
or U21470 (N_21470,N_18899,N_18669);
or U21471 (N_21471,N_19390,N_17986);
and U21472 (N_21472,N_17550,N_18023);
nand U21473 (N_21473,N_18184,N_18693);
xor U21474 (N_21474,N_17669,N_18579);
and U21475 (N_21475,N_18620,N_19279);
xor U21476 (N_21476,N_17651,N_18155);
xor U21477 (N_21477,N_18074,N_17594);
xnor U21478 (N_21478,N_18043,N_18810);
xnor U21479 (N_21479,N_18698,N_18973);
and U21480 (N_21480,N_19504,N_19289);
and U21481 (N_21481,N_18714,N_17695);
or U21482 (N_21482,N_18736,N_18181);
nand U21483 (N_21483,N_17983,N_19522);
and U21484 (N_21484,N_17840,N_17667);
nand U21485 (N_21485,N_17620,N_18836);
or U21486 (N_21486,N_19079,N_19532);
nor U21487 (N_21487,N_19752,N_18214);
and U21488 (N_21488,N_17858,N_17820);
or U21489 (N_21489,N_17975,N_18667);
nor U21490 (N_21490,N_19834,N_19838);
and U21491 (N_21491,N_18959,N_19379);
and U21492 (N_21492,N_18636,N_18072);
or U21493 (N_21493,N_18777,N_18347);
and U21494 (N_21494,N_17912,N_18622);
nor U21495 (N_21495,N_19367,N_17718);
nor U21496 (N_21496,N_19485,N_19769);
nor U21497 (N_21497,N_17739,N_19481);
nand U21498 (N_21498,N_19114,N_19942);
nand U21499 (N_21499,N_19032,N_18961);
or U21500 (N_21500,N_17693,N_17841);
nor U21501 (N_21501,N_18803,N_17588);
nand U21502 (N_21502,N_18649,N_17649);
and U21503 (N_21503,N_17691,N_17670);
nor U21504 (N_21504,N_19272,N_17979);
or U21505 (N_21505,N_19334,N_18312);
or U21506 (N_21506,N_18272,N_19742);
xnor U21507 (N_21507,N_17864,N_18147);
or U21508 (N_21508,N_17594,N_19834);
nor U21509 (N_21509,N_19707,N_19510);
and U21510 (N_21510,N_17807,N_19740);
nor U21511 (N_21511,N_19378,N_18108);
or U21512 (N_21512,N_18641,N_19323);
nand U21513 (N_21513,N_19535,N_18631);
or U21514 (N_21514,N_18510,N_19806);
nor U21515 (N_21515,N_17805,N_18640);
and U21516 (N_21516,N_17956,N_17784);
nor U21517 (N_21517,N_19211,N_18360);
nor U21518 (N_21518,N_18364,N_19546);
and U21519 (N_21519,N_19782,N_17731);
nand U21520 (N_21520,N_18060,N_18530);
and U21521 (N_21521,N_19817,N_18372);
or U21522 (N_21522,N_19469,N_18680);
and U21523 (N_21523,N_18552,N_18543);
or U21524 (N_21524,N_18389,N_19839);
nor U21525 (N_21525,N_18187,N_19877);
and U21526 (N_21526,N_18556,N_19156);
nand U21527 (N_21527,N_18946,N_19261);
nor U21528 (N_21528,N_18881,N_19783);
nand U21529 (N_21529,N_19706,N_18083);
nand U21530 (N_21530,N_19444,N_19891);
or U21531 (N_21531,N_19257,N_17938);
nor U21532 (N_21532,N_18028,N_19609);
and U21533 (N_21533,N_18914,N_18245);
xor U21534 (N_21534,N_17695,N_19644);
nand U21535 (N_21535,N_18487,N_19434);
nor U21536 (N_21536,N_17510,N_18037);
or U21537 (N_21537,N_19943,N_17695);
nand U21538 (N_21538,N_18210,N_19482);
nand U21539 (N_21539,N_19986,N_19565);
and U21540 (N_21540,N_18142,N_19466);
and U21541 (N_21541,N_18959,N_18101);
and U21542 (N_21542,N_18673,N_19614);
xor U21543 (N_21543,N_19456,N_17660);
nand U21544 (N_21544,N_18606,N_18711);
and U21545 (N_21545,N_18469,N_18655);
xnor U21546 (N_21546,N_19077,N_18909);
nand U21547 (N_21547,N_18470,N_17709);
nand U21548 (N_21548,N_19776,N_18677);
nand U21549 (N_21549,N_17661,N_19625);
and U21550 (N_21550,N_17668,N_18782);
nor U21551 (N_21551,N_18612,N_19711);
nand U21552 (N_21552,N_18142,N_19007);
or U21553 (N_21553,N_17897,N_19249);
and U21554 (N_21554,N_18629,N_18554);
or U21555 (N_21555,N_19959,N_18591);
nor U21556 (N_21556,N_18649,N_17683);
or U21557 (N_21557,N_19758,N_19398);
and U21558 (N_21558,N_17851,N_19810);
nand U21559 (N_21559,N_19887,N_18083);
or U21560 (N_21560,N_18423,N_17506);
nor U21561 (N_21561,N_18188,N_19880);
or U21562 (N_21562,N_19299,N_17657);
and U21563 (N_21563,N_18391,N_18852);
or U21564 (N_21564,N_19511,N_19812);
nand U21565 (N_21565,N_17971,N_19925);
and U21566 (N_21566,N_19195,N_18468);
nor U21567 (N_21567,N_19068,N_19434);
and U21568 (N_21568,N_17792,N_18277);
and U21569 (N_21569,N_18791,N_19893);
nor U21570 (N_21570,N_19673,N_18671);
nand U21571 (N_21571,N_18011,N_19531);
xnor U21572 (N_21572,N_19157,N_18925);
and U21573 (N_21573,N_18016,N_18117);
and U21574 (N_21574,N_18210,N_19845);
nor U21575 (N_21575,N_19821,N_18275);
or U21576 (N_21576,N_19286,N_19690);
nor U21577 (N_21577,N_18104,N_17926);
nor U21578 (N_21578,N_19799,N_18078);
or U21579 (N_21579,N_18194,N_19301);
or U21580 (N_21580,N_17806,N_17584);
nand U21581 (N_21581,N_18101,N_19150);
or U21582 (N_21582,N_18178,N_17927);
and U21583 (N_21583,N_19412,N_19077);
xnor U21584 (N_21584,N_18765,N_18705);
and U21585 (N_21585,N_19469,N_17819);
and U21586 (N_21586,N_19923,N_18467);
nor U21587 (N_21587,N_18357,N_17595);
and U21588 (N_21588,N_17969,N_18266);
or U21589 (N_21589,N_19501,N_17538);
and U21590 (N_21590,N_19493,N_17502);
nand U21591 (N_21591,N_19395,N_19415);
or U21592 (N_21592,N_19717,N_17742);
nor U21593 (N_21593,N_19282,N_18836);
or U21594 (N_21594,N_18735,N_18357);
and U21595 (N_21595,N_19171,N_18001);
xnor U21596 (N_21596,N_18525,N_18906);
xor U21597 (N_21597,N_18948,N_18900);
nand U21598 (N_21598,N_17522,N_18763);
and U21599 (N_21599,N_19736,N_18248);
nor U21600 (N_21600,N_18907,N_17932);
nand U21601 (N_21601,N_19337,N_18868);
and U21602 (N_21602,N_19999,N_18439);
and U21603 (N_21603,N_19679,N_19229);
and U21604 (N_21604,N_19738,N_18547);
nor U21605 (N_21605,N_19690,N_18853);
nor U21606 (N_21606,N_19197,N_18207);
nor U21607 (N_21607,N_19383,N_19756);
nand U21608 (N_21608,N_17966,N_19837);
and U21609 (N_21609,N_19082,N_19896);
and U21610 (N_21610,N_17647,N_19222);
nand U21611 (N_21611,N_19245,N_18490);
nor U21612 (N_21612,N_18734,N_19120);
or U21613 (N_21613,N_19184,N_17576);
or U21614 (N_21614,N_18660,N_18680);
xor U21615 (N_21615,N_18116,N_18223);
or U21616 (N_21616,N_19733,N_18099);
and U21617 (N_21617,N_17639,N_18090);
nand U21618 (N_21618,N_19033,N_18989);
xnor U21619 (N_21619,N_18166,N_18241);
nor U21620 (N_21620,N_19101,N_19813);
nand U21621 (N_21621,N_17899,N_17687);
and U21622 (N_21622,N_17751,N_18339);
nand U21623 (N_21623,N_17771,N_18168);
nand U21624 (N_21624,N_17881,N_19622);
or U21625 (N_21625,N_19378,N_18147);
nor U21626 (N_21626,N_17686,N_18029);
nor U21627 (N_21627,N_19893,N_18167);
and U21628 (N_21628,N_18448,N_17507);
nor U21629 (N_21629,N_19115,N_19621);
or U21630 (N_21630,N_17718,N_19244);
nand U21631 (N_21631,N_18859,N_18745);
or U21632 (N_21632,N_19433,N_18881);
nand U21633 (N_21633,N_17952,N_19275);
or U21634 (N_21634,N_19229,N_17895);
nor U21635 (N_21635,N_18058,N_19535);
or U21636 (N_21636,N_17585,N_19085);
and U21637 (N_21637,N_18984,N_19461);
xnor U21638 (N_21638,N_17862,N_18508);
and U21639 (N_21639,N_19104,N_18479);
nand U21640 (N_21640,N_17584,N_18467);
and U21641 (N_21641,N_18477,N_18336);
nand U21642 (N_21642,N_19617,N_18633);
nand U21643 (N_21643,N_19894,N_17646);
and U21644 (N_21644,N_18534,N_19334);
nor U21645 (N_21645,N_18852,N_19647);
xnor U21646 (N_21646,N_19561,N_17724);
and U21647 (N_21647,N_17944,N_19055);
or U21648 (N_21648,N_19585,N_19815);
nor U21649 (N_21649,N_19803,N_18290);
nand U21650 (N_21650,N_17805,N_19627);
and U21651 (N_21651,N_19586,N_18091);
nand U21652 (N_21652,N_17718,N_17806);
or U21653 (N_21653,N_17846,N_19446);
and U21654 (N_21654,N_18634,N_19854);
and U21655 (N_21655,N_18208,N_19618);
or U21656 (N_21656,N_18733,N_19203);
or U21657 (N_21657,N_19653,N_18751);
or U21658 (N_21658,N_19850,N_19337);
or U21659 (N_21659,N_18318,N_18380);
and U21660 (N_21660,N_19529,N_18333);
nand U21661 (N_21661,N_17627,N_18293);
nor U21662 (N_21662,N_17827,N_19856);
nand U21663 (N_21663,N_17653,N_17858);
nand U21664 (N_21664,N_19992,N_18684);
nor U21665 (N_21665,N_18944,N_18106);
or U21666 (N_21666,N_19061,N_18067);
nor U21667 (N_21667,N_19700,N_18974);
or U21668 (N_21668,N_17898,N_19398);
nand U21669 (N_21669,N_18369,N_19840);
nand U21670 (N_21670,N_18428,N_19896);
nand U21671 (N_21671,N_18060,N_17790);
and U21672 (N_21672,N_19448,N_17563);
and U21673 (N_21673,N_17561,N_19552);
nand U21674 (N_21674,N_19499,N_17938);
xnor U21675 (N_21675,N_19966,N_18494);
nand U21676 (N_21676,N_19226,N_18990);
nor U21677 (N_21677,N_19916,N_17870);
nand U21678 (N_21678,N_18507,N_19565);
and U21679 (N_21679,N_18660,N_18912);
nand U21680 (N_21680,N_17522,N_18417);
xor U21681 (N_21681,N_19149,N_18742);
and U21682 (N_21682,N_19298,N_19748);
nand U21683 (N_21683,N_17880,N_19453);
nand U21684 (N_21684,N_18604,N_19684);
nor U21685 (N_21685,N_19357,N_18591);
and U21686 (N_21686,N_18205,N_19690);
or U21687 (N_21687,N_18578,N_17635);
and U21688 (N_21688,N_18200,N_17888);
and U21689 (N_21689,N_19792,N_19946);
xor U21690 (N_21690,N_19646,N_17690);
or U21691 (N_21691,N_17647,N_18488);
nand U21692 (N_21692,N_19026,N_18920);
and U21693 (N_21693,N_19524,N_18912);
or U21694 (N_21694,N_18153,N_18311);
nand U21695 (N_21695,N_17728,N_19547);
xor U21696 (N_21696,N_19715,N_18989);
or U21697 (N_21697,N_18979,N_17633);
nor U21698 (N_21698,N_19821,N_18351);
or U21699 (N_21699,N_19125,N_19768);
nor U21700 (N_21700,N_19784,N_19344);
nand U21701 (N_21701,N_19117,N_17610);
xnor U21702 (N_21702,N_18206,N_19024);
nor U21703 (N_21703,N_18693,N_19497);
or U21704 (N_21704,N_18701,N_18886);
or U21705 (N_21705,N_19138,N_19970);
nor U21706 (N_21706,N_19138,N_18620);
nand U21707 (N_21707,N_18846,N_17654);
xnor U21708 (N_21708,N_18164,N_19793);
and U21709 (N_21709,N_18275,N_18299);
xor U21710 (N_21710,N_17576,N_18190);
nand U21711 (N_21711,N_17694,N_19263);
or U21712 (N_21712,N_18297,N_19218);
nand U21713 (N_21713,N_19910,N_19732);
or U21714 (N_21714,N_19397,N_18505);
nand U21715 (N_21715,N_17511,N_18163);
or U21716 (N_21716,N_18395,N_19940);
nor U21717 (N_21717,N_19578,N_18636);
nor U21718 (N_21718,N_19607,N_18752);
nor U21719 (N_21719,N_19604,N_18305);
nand U21720 (N_21720,N_17801,N_19168);
nand U21721 (N_21721,N_17793,N_19636);
xor U21722 (N_21722,N_18453,N_17984);
or U21723 (N_21723,N_18785,N_17688);
or U21724 (N_21724,N_19722,N_18128);
or U21725 (N_21725,N_19305,N_19744);
or U21726 (N_21726,N_18053,N_17878);
nand U21727 (N_21727,N_19986,N_18060);
and U21728 (N_21728,N_18492,N_18385);
or U21729 (N_21729,N_19528,N_19540);
and U21730 (N_21730,N_19648,N_19766);
xnor U21731 (N_21731,N_18538,N_19358);
nor U21732 (N_21732,N_18933,N_19438);
nand U21733 (N_21733,N_18946,N_17710);
and U21734 (N_21734,N_19979,N_18092);
nand U21735 (N_21735,N_19616,N_19545);
nor U21736 (N_21736,N_19985,N_18855);
nand U21737 (N_21737,N_17705,N_18330);
or U21738 (N_21738,N_19505,N_19461);
nand U21739 (N_21739,N_17942,N_18449);
nand U21740 (N_21740,N_17936,N_19064);
and U21741 (N_21741,N_17547,N_18896);
or U21742 (N_21742,N_19783,N_18855);
nor U21743 (N_21743,N_17532,N_19899);
nand U21744 (N_21744,N_18946,N_19210);
or U21745 (N_21745,N_17647,N_19287);
and U21746 (N_21746,N_19618,N_17940);
and U21747 (N_21747,N_19488,N_18145);
nor U21748 (N_21748,N_18109,N_18761);
nor U21749 (N_21749,N_18274,N_19513);
and U21750 (N_21750,N_19141,N_17951);
or U21751 (N_21751,N_17567,N_17879);
or U21752 (N_21752,N_18957,N_19905);
nand U21753 (N_21753,N_17844,N_17763);
or U21754 (N_21754,N_18588,N_19836);
and U21755 (N_21755,N_19430,N_18526);
and U21756 (N_21756,N_17730,N_17792);
nand U21757 (N_21757,N_19897,N_18111);
and U21758 (N_21758,N_19994,N_18437);
or U21759 (N_21759,N_19261,N_17999);
nor U21760 (N_21760,N_17855,N_19671);
or U21761 (N_21761,N_18342,N_18598);
nor U21762 (N_21762,N_19586,N_19954);
nor U21763 (N_21763,N_19486,N_17685);
nor U21764 (N_21764,N_17650,N_19609);
and U21765 (N_21765,N_19275,N_17507);
nand U21766 (N_21766,N_18061,N_19668);
nor U21767 (N_21767,N_18029,N_19619);
or U21768 (N_21768,N_18705,N_17913);
or U21769 (N_21769,N_19766,N_18088);
and U21770 (N_21770,N_17746,N_19916);
or U21771 (N_21771,N_17805,N_19565);
nand U21772 (N_21772,N_18019,N_19885);
nor U21773 (N_21773,N_17790,N_19174);
xnor U21774 (N_21774,N_17775,N_19224);
or U21775 (N_21775,N_19709,N_18186);
nor U21776 (N_21776,N_18029,N_18835);
and U21777 (N_21777,N_18145,N_19708);
nand U21778 (N_21778,N_18895,N_17604);
xor U21779 (N_21779,N_18970,N_17693);
and U21780 (N_21780,N_17707,N_17854);
nor U21781 (N_21781,N_19118,N_19699);
and U21782 (N_21782,N_19182,N_18669);
and U21783 (N_21783,N_19893,N_18058);
nand U21784 (N_21784,N_19220,N_19911);
and U21785 (N_21785,N_18628,N_19156);
or U21786 (N_21786,N_19014,N_18255);
nand U21787 (N_21787,N_19331,N_18681);
xor U21788 (N_21788,N_19800,N_19111);
or U21789 (N_21789,N_19173,N_19880);
and U21790 (N_21790,N_19963,N_17793);
or U21791 (N_21791,N_17820,N_19905);
or U21792 (N_21792,N_18011,N_17892);
or U21793 (N_21793,N_17589,N_19302);
and U21794 (N_21794,N_17648,N_17976);
nor U21795 (N_21795,N_19645,N_19620);
nor U21796 (N_21796,N_19235,N_19421);
or U21797 (N_21797,N_17622,N_19955);
or U21798 (N_21798,N_19358,N_18913);
nor U21799 (N_21799,N_18461,N_18441);
and U21800 (N_21800,N_18026,N_19510);
xnor U21801 (N_21801,N_18093,N_19830);
and U21802 (N_21802,N_18762,N_18833);
and U21803 (N_21803,N_19616,N_19770);
nor U21804 (N_21804,N_19237,N_18865);
nor U21805 (N_21805,N_19926,N_19081);
nand U21806 (N_21806,N_17718,N_19713);
nor U21807 (N_21807,N_19508,N_19101);
or U21808 (N_21808,N_19159,N_17699);
nor U21809 (N_21809,N_19461,N_19450);
xnor U21810 (N_21810,N_19223,N_17793);
or U21811 (N_21811,N_19492,N_17508);
or U21812 (N_21812,N_18732,N_18943);
nand U21813 (N_21813,N_19230,N_17691);
and U21814 (N_21814,N_19352,N_19987);
nor U21815 (N_21815,N_18261,N_17881);
and U21816 (N_21816,N_18139,N_18808);
or U21817 (N_21817,N_17595,N_19287);
nand U21818 (N_21818,N_19448,N_17733);
nand U21819 (N_21819,N_18947,N_18776);
nor U21820 (N_21820,N_19045,N_19575);
or U21821 (N_21821,N_19932,N_17645);
nand U21822 (N_21822,N_17795,N_18315);
nor U21823 (N_21823,N_19800,N_17679);
and U21824 (N_21824,N_18000,N_19943);
nor U21825 (N_21825,N_19633,N_18541);
nand U21826 (N_21826,N_17532,N_19967);
nor U21827 (N_21827,N_19938,N_18688);
and U21828 (N_21828,N_19352,N_19766);
and U21829 (N_21829,N_18181,N_19342);
xnor U21830 (N_21830,N_19518,N_18779);
nor U21831 (N_21831,N_19125,N_17628);
nor U21832 (N_21832,N_18525,N_17627);
or U21833 (N_21833,N_19280,N_18309);
nand U21834 (N_21834,N_19264,N_19292);
nand U21835 (N_21835,N_18994,N_19608);
nand U21836 (N_21836,N_17886,N_18042);
nor U21837 (N_21837,N_17691,N_19565);
or U21838 (N_21838,N_19805,N_17706);
and U21839 (N_21839,N_18270,N_19105);
nand U21840 (N_21840,N_19116,N_18659);
nand U21841 (N_21841,N_19382,N_17695);
or U21842 (N_21842,N_17603,N_18897);
or U21843 (N_21843,N_18404,N_18311);
nand U21844 (N_21844,N_17772,N_17991);
or U21845 (N_21845,N_17838,N_18449);
nand U21846 (N_21846,N_18211,N_18794);
or U21847 (N_21847,N_19844,N_18197);
nand U21848 (N_21848,N_17851,N_17715);
and U21849 (N_21849,N_19110,N_19735);
and U21850 (N_21850,N_17637,N_18205);
and U21851 (N_21851,N_19053,N_19608);
xor U21852 (N_21852,N_18198,N_19408);
nand U21853 (N_21853,N_17881,N_19284);
or U21854 (N_21854,N_18544,N_17621);
nand U21855 (N_21855,N_18597,N_19574);
xor U21856 (N_21856,N_19111,N_18539);
and U21857 (N_21857,N_17676,N_18426);
or U21858 (N_21858,N_19678,N_19865);
and U21859 (N_21859,N_18197,N_19578);
nor U21860 (N_21860,N_18566,N_17518);
or U21861 (N_21861,N_17748,N_18912);
or U21862 (N_21862,N_19364,N_18917);
and U21863 (N_21863,N_18089,N_18725);
nand U21864 (N_21864,N_18319,N_19046);
and U21865 (N_21865,N_18269,N_18166);
or U21866 (N_21866,N_19326,N_17514);
nor U21867 (N_21867,N_19322,N_19962);
or U21868 (N_21868,N_19338,N_18223);
and U21869 (N_21869,N_19104,N_18325);
or U21870 (N_21870,N_18513,N_18969);
or U21871 (N_21871,N_19366,N_18351);
or U21872 (N_21872,N_19187,N_18405);
and U21873 (N_21873,N_19032,N_19482);
or U21874 (N_21874,N_18978,N_18485);
nor U21875 (N_21875,N_19974,N_17786);
nor U21876 (N_21876,N_19524,N_18289);
and U21877 (N_21877,N_18677,N_19194);
nand U21878 (N_21878,N_17550,N_18802);
or U21879 (N_21879,N_17956,N_19338);
nand U21880 (N_21880,N_19264,N_17747);
or U21881 (N_21881,N_19472,N_17665);
or U21882 (N_21882,N_19044,N_18803);
nor U21883 (N_21883,N_19637,N_18137);
nor U21884 (N_21884,N_19007,N_18634);
nor U21885 (N_21885,N_19108,N_17718);
xnor U21886 (N_21886,N_18368,N_18896);
and U21887 (N_21887,N_19169,N_19170);
nor U21888 (N_21888,N_18493,N_17996);
nor U21889 (N_21889,N_19442,N_19490);
xnor U21890 (N_21890,N_18242,N_18284);
and U21891 (N_21891,N_19465,N_18598);
and U21892 (N_21892,N_18535,N_19156);
nor U21893 (N_21893,N_17565,N_19944);
or U21894 (N_21894,N_19735,N_17571);
and U21895 (N_21895,N_19324,N_19560);
nor U21896 (N_21896,N_19157,N_18734);
nand U21897 (N_21897,N_18577,N_19604);
nor U21898 (N_21898,N_19263,N_18294);
xor U21899 (N_21899,N_17858,N_17616);
nor U21900 (N_21900,N_19677,N_18591);
nand U21901 (N_21901,N_19159,N_17973);
nand U21902 (N_21902,N_18686,N_18288);
nor U21903 (N_21903,N_18929,N_18480);
and U21904 (N_21904,N_18226,N_18425);
or U21905 (N_21905,N_18256,N_17590);
and U21906 (N_21906,N_19554,N_19285);
nor U21907 (N_21907,N_19250,N_19491);
nor U21908 (N_21908,N_19198,N_17537);
nor U21909 (N_21909,N_18073,N_19621);
nand U21910 (N_21910,N_17857,N_18246);
nand U21911 (N_21911,N_17743,N_19421);
nor U21912 (N_21912,N_18244,N_19810);
nand U21913 (N_21913,N_18421,N_19989);
or U21914 (N_21914,N_18517,N_18563);
nand U21915 (N_21915,N_19125,N_18056);
nor U21916 (N_21916,N_19870,N_18748);
nor U21917 (N_21917,N_19364,N_18850);
or U21918 (N_21918,N_19233,N_18857);
and U21919 (N_21919,N_17582,N_19765);
nand U21920 (N_21920,N_19278,N_19336);
or U21921 (N_21921,N_18526,N_19471);
or U21922 (N_21922,N_18572,N_18831);
nor U21923 (N_21923,N_18567,N_18626);
nor U21924 (N_21924,N_19509,N_18272);
or U21925 (N_21925,N_19924,N_19259);
nand U21926 (N_21926,N_18833,N_18125);
nand U21927 (N_21927,N_17723,N_19498);
nor U21928 (N_21928,N_17724,N_17889);
xor U21929 (N_21929,N_19776,N_19034);
nand U21930 (N_21930,N_18107,N_19866);
nor U21931 (N_21931,N_17817,N_17543);
and U21932 (N_21932,N_18893,N_18097);
or U21933 (N_21933,N_18832,N_19431);
nand U21934 (N_21934,N_18124,N_19644);
xnor U21935 (N_21935,N_18117,N_18328);
nor U21936 (N_21936,N_18428,N_18133);
nor U21937 (N_21937,N_19977,N_19878);
nand U21938 (N_21938,N_18771,N_17708);
nor U21939 (N_21939,N_18230,N_19264);
or U21940 (N_21940,N_19367,N_17932);
or U21941 (N_21941,N_18025,N_18393);
nand U21942 (N_21942,N_18676,N_18437);
or U21943 (N_21943,N_19288,N_18520);
xor U21944 (N_21944,N_18984,N_18397);
and U21945 (N_21945,N_18070,N_19001);
nand U21946 (N_21946,N_19941,N_18262);
nor U21947 (N_21947,N_17789,N_18790);
nor U21948 (N_21948,N_19666,N_18378);
nand U21949 (N_21949,N_18105,N_18726);
or U21950 (N_21950,N_19264,N_17618);
nand U21951 (N_21951,N_18511,N_17801);
and U21952 (N_21952,N_17516,N_19266);
nand U21953 (N_21953,N_18496,N_18997);
and U21954 (N_21954,N_19931,N_19736);
and U21955 (N_21955,N_19324,N_18177);
xnor U21956 (N_21956,N_17754,N_18736);
or U21957 (N_21957,N_19172,N_19684);
nor U21958 (N_21958,N_18892,N_18442);
and U21959 (N_21959,N_19964,N_19082);
nand U21960 (N_21960,N_19089,N_19478);
xnor U21961 (N_21961,N_17656,N_19496);
nand U21962 (N_21962,N_19876,N_19991);
nor U21963 (N_21963,N_18052,N_17805);
nand U21964 (N_21964,N_18747,N_19430);
and U21965 (N_21965,N_17789,N_19617);
nor U21966 (N_21966,N_18785,N_18424);
and U21967 (N_21967,N_18228,N_18374);
and U21968 (N_21968,N_18748,N_18182);
or U21969 (N_21969,N_18603,N_18586);
nor U21970 (N_21970,N_17916,N_17745);
and U21971 (N_21971,N_17753,N_18600);
and U21972 (N_21972,N_18769,N_19800);
and U21973 (N_21973,N_18807,N_17714);
nand U21974 (N_21974,N_18953,N_19779);
or U21975 (N_21975,N_19110,N_18310);
nor U21976 (N_21976,N_18635,N_19978);
xor U21977 (N_21977,N_19791,N_18614);
nand U21978 (N_21978,N_18651,N_17856);
and U21979 (N_21979,N_19440,N_17824);
or U21980 (N_21980,N_19681,N_19604);
nor U21981 (N_21981,N_19593,N_18439);
or U21982 (N_21982,N_19349,N_18243);
and U21983 (N_21983,N_19992,N_19125);
nand U21984 (N_21984,N_18609,N_19174);
nor U21985 (N_21985,N_17509,N_18835);
and U21986 (N_21986,N_17864,N_18939);
nor U21987 (N_21987,N_18800,N_19613);
nor U21988 (N_21988,N_19275,N_19271);
and U21989 (N_21989,N_19072,N_19168);
nor U21990 (N_21990,N_19421,N_18958);
nand U21991 (N_21991,N_19816,N_19437);
nand U21992 (N_21992,N_19042,N_18012);
nor U21993 (N_21993,N_17503,N_19501);
and U21994 (N_21994,N_19796,N_18755);
nor U21995 (N_21995,N_19332,N_19660);
xnor U21996 (N_21996,N_19312,N_19358);
and U21997 (N_21997,N_18235,N_19697);
and U21998 (N_21998,N_17698,N_19783);
and U21999 (N_21999,N_18491,N_18394);
nor U22000 (N_22000,N_18224,N_18764);
or U22001 (N_22001,N_18554,N_17687);
nand U22002 (N_22002,N_19452,N_18565);
or U22003 (N_22003,N_19447,N_17650);
nor U22004 (N_22004,N_18657,N_19190);
and U22005 (N_22005,N_17735,N_17673);
or U22006 (N_22006,N_18015,N_18954);
nand U22007 (N_22007,N_19010,N_19487);
nor U22008 (N_22008,N_18182,N_19631);
nor U22009 (N_22009,N_19894,N_18961);
nor U22010 (N_22010,N_18605,N_19833);
nand U22011 (N_22011,N_17518,N_18144);
and U22012 (N_22012,N_19703,N_17827);
nor U22013 (N_22013,N_18369,N_18228);
or U22014 (N_22014,N_19161,N_19831);
nand U22015 (N_22015,N_18140,N_19200);
and U22016 (N_22016,N_19154,N_19123);
or U22017 (N_22017,N_18510,N_17950);
nor U22018 (N_22018,N_17913,N_19502);
and U22019 (N_22019,N_19718,N_19923);
nand U22020 (N_22020,N_18682,N_18161);
or U22021 (N_22021,N_18127,N_17780);
nand U22022 (N_22022,N_18590,N_18703);
nand U22023 (N_22023,N_19136,N_19601);
and U22024 (N_22024,N_18520,N_19857);
xor U22025 (N_22025,N_19369,N_18474);
or U22026 (N_22026,N_18878,N_17962);
nor U22027 (N_22027,N_19227,N_17995);
and U22028 (N_22028,N_19427,N_19136);
xor U22029 (N_22029,N_17924,N_19815);
nor U22030 (N_22030,N_19173,N_18616);
nand U22031 (N_22031,N_18339,N_19289);
and U22032 (N_22032,N_17586,N_19063);
nor U22033 (N_22033,N_19543,N_18713);
nand U22034 (N_22034,N_18018,N_18632);
nor U22035 (N_22035,N_19082,N_18226);
or U22036 (N_22036,N_17558,N_17822);
xor U22037 (N_22037,N_18292,N_19246);
and U22038 (N_22038,N_17834,N_18711);
xor U22039 (N_22039,N_19626,N_19590);
nor U22040 (N_22040,N_19067,N_17976);
nor U22041 (N_22041,N_17633,N_19705);
xnor U22042 (N_22042,N_17557,N_17985);
nor U22043 (N_22043,N_19856,N_19034);
nand U22044 (N_22044,N_17728,N_18648);
nor U22045 (N_22045,N_17575,N_19549);
or U22046 (N_22046,N_18675,N_18691);
and U22047 (N_22047,N_17619,N_19549);
nand U22048 (N_22048,N_19229,N_18170);
or U22049 (N_22049,N_18790,N_17896);
nand U22050 (N_22050,N_19179,N_19061);
nand U22051 (N_22051,N_19753,N_19110);
and U22052 (N_22052,N_17798,N_18008);
and U22053 (N_22053,N_19643,N_17954);
or U22054 (N_22054,N_19981,N_19053);
nand U22055 (N_22055,N_18668,N_17507);
or U22056 (N_22056,N_17553,N_18003);
nand U22057 (N_22057,N_17692,N_19936);
xnor U22058 (N_22058,N_19125,N_19180);
nor U22059 (N_22059,N_19806,N_18482);
nor U22060 (N_22060,N_18990,N_19151);
xnor U22061 (N_22061,N_19636,N_17982);
and U22062 (N_22062,N_18668,N_19063);
or U22063 (N_22063,N_18088,N_19235);
and U22064 (N_22064,N_18480,N_18630);
and U22065 (N_22065,N_19455,N_19297);
and U22066 (N_22066,N_18509,N_19301);
or U22067 (N_22067,N_19080,N_18653);
or U22068 (N_22068,N_17867,N_19533);
or U22069 (N_22069,N_19785,N_19044);
nor U22070 (N_22070,N_18644,N_18889);
or U22071 (N_22071,N_19379,N_17973);
and U22072 (N_22072,N_19557,N_19652);
and U22073 (N_22073,N_18428,N_19345);
or U22074 (N_22074,N_18266,N_19204);
and U22075 (N_22075,N_19650,N_17605);
nor U22076 (N_22076,N_19383,N_19580);
and U22077 (N_22077,N_17987,N_19869);
xor U22078 (N_22078,N_18009,N_19013);
nand U22079 (N_22079,N_17763,N_17818);
or U22080 (N_22080,N_17586,N_18365);
and U22081 (N_22081,N_17505,N_19224);
or U22082 (N_22082,N_18763,N_18964);
nor U22083 (N_22083,N_17606,N_18023);
or U22084 (N_22084,N_17939,N_19331);
nand U22085 (N_22085,N_17763,N_19016);
xor U22086 (N_22086,N_19405,N_17865);
nand U22087 (N_22087,N_19622,N_19818);
nor U22088 (N_22088,N_19753,N_19653);
nand U22089 (N_22089,N_19712,N_18227);
nor U22090 (N_22090,N_17812,N_18693);
and U22091 (N_22091,N_19044,N_18589);
nor U22092 (N_22092,N_18206,N_18557);
or U22093 (N_22093,N_19135,N_18385);
nand U22094 (N_22094,N_17719,N_19191);
nand U22095 (N_22095,N_18492,N_19178);
nor U22096 (N_22096,N_18483,N_18098);
nor U22097 (N_22097,N_19993,N_19490);
or U22098 (N_22098,N_19053,N_18843);
nand U22099 (N_22099,N_19262,N_18430);
xor U22100 (N_22100,N_17916,N_18562);
xor U22101 (N_22101,N_18117,N_19849);
nand U22102 (N_22102,N_18489,N_18488);
nand U22103 (N_22103,N_19924,N_18105);
and U22104 (N_22104,N_18726,N_17648);
nor U22105 (N_22105,N_19358,N_19880);
or U22106 (N_22106,N_19157,N_18854);
and U22107 (N_22107,N_18512,N_18842);
or U22108 (N_22108,N_19705,N_17719);
and U22109 (N_22109,N_19235,N_17666);
or U22110 (N_22110,N_17588,N_17502);
nor U22111 (N_22111,N_19104,N_17892);
nand U22112 (N_22112,N_18362,N_18243);
xnor U22113 (N_22113,N_19107,N_17700);
xor U22114 (N_22114,N_18620,N_18849);
or U22115 (N_22115,N_17885,N_19447);
xor U22116 (N_22116,N_17862,N_17593);
or U22117 (N_22117,N_18257,N_19707);
or U22118 (N_22118,N_19667,N_19769);
nor U22119 (N_22119,N_18633,N_19443);
and U22120 (N_22120,N_17862,N_18502);
and U22121 (N_22121,N_18579,N_18015);
nor U22122 (N_22122,N_17928,N_18102);
and U22123 (N_22123,N_19857,N_18912);
and U22124 (N_22124,N_19748,N_19033);
and U22125 (N_22125,N_17583,N_19104);
nand U22126 (N_22126,N_18732,N_19292);
and U22127 (N_22127,N_19785,N_17980);
nor U22128 (N_22128,N_18286,N_17858);
nand U22129 (N_22129,N_19457,N_18770);
nor U22130 (N_22130,N_19146,N_19454);
nor U22131 (N_22131,N_19154,N_19211);
xor U22132 (N_22132,N_17992,N_18507);
and U22133 (N_22133,N_17875,N_18407);
nand U22134 (N_22134,N_18449,N_18611);
nand U22135 (N_22135,N_19364,N_18884);
xor U22136 (N_22136,N_18761,N_19384);
nand U22137 (N_22137,N_19610,N_18428);
nor U22138 (N_22138,N_19506,N_18495);
or U22139 (N_22139,N_19022,N_19222);
nor U22140 (N_22140,N_19179,N_17507);
or U22141 (N_22141,N_18384,N_18273);
or U22142 (N_22142,N_18541,N_19934);
or U22143 (N_22143,N_17525,N_19494);
nor U22144 (N_22144,N_19854,N_19292);
nor U22145 (N_22145,N_18402,N_18576);
or U22146 (N_22146,N_18435,N_19813);
or U22147 (N_22147,N_18397,N_18861);
or U22148 (N_22148,N_19583,N_17837);
nand U22149 (N_22149,N_17549,N_18607);
and U22150 (N_22150,N_18664,N_18004);
or U22151 (N_22151,N_19828,N_19053);
nor U22152 (N_22152,N_19111,N_18646);
nand U22153 (N_22153,N_19606,N_17629);
or U22154 (N_22154,N_18907,N_19270);
or U22155 (N_22155,N_18955,N_19838);
nand U22156 (N_22156,N_17747,N_17516);
nand U22157 (N_22157,N_19337,N_17990);
or U22158 (N_22158,N_18546,N_19433);
nor U22159 (N_22159,N_18176,N_17642);
xor U22160 (N_22160,N_19311,N_18972);
or U22161 (N_22161,N_18770,N_18755);
nor U22162 (N_22162,N_19910,N_19657);
xor U22163 (N_22163,N_18310,N_17512);
nor U22164 (N_22164,N_18176,N_18949);
xnor U22165 (N_22165,N_19682,N_19905);
nor U22166 (N_22166,N_17561,N_18702);
xnor U22167 (N_22167,N_17743,N_17618);
nor U22168 (N_22168,N_19104,N_19896);
or U22169 (N_22169,N_19692,N_19651);
or U22170 (N_22170,N_18414,N_18905);
and U22171 (N_22171,N_17739,N_17742);
and U22172 (N_22172,N_19869,N_17569);
or U22173 (N_22173,N_18562,N_17758);
nand U22174 (N_22174,N_19357,N_18163);
nor U22175 (N_22175,N_19469,N_18623);
or U22176 (N_22176,N_19160,N_17788);
nor U22177 (N_22177,N_17762,N_18105);
or U22178 (N_22178,N_18871,N_17644);
nor U22179 (N_22179,N_18987,N_19404);
nand U22180 (N_22180,N_18704,N_18142);
nand U22181 (N_22181,N_17724,N_17990);
xor U22182 (N_22182,N_17970,N_18781);
and U22183 (N_22183,N_18052,N_17751);
nand U22184 (N_22184,N_17939,N_18696);
and U22185 (N_22185,N_19265,N_18066);
nor U22186 (N_22186,N_17567,N_19777);
nand U22187 (N_22187,N_17874,N_18889);
nand U22188 (N_22188,N_19973,N_17976);
and U22189 (N_22189,N_19207,N_18622);
or U22190 (N_22190,N_19563,N_17726);
or U22191 (N_22191,N_18638,N_17791);
xnor U22192 (N_22192,N_18528,N_18104);
nand U22193 (N_22193,N_18143,N_18534);
and U22194 (N_22194,N_19795,N_19220);
nand U22195 (N_22195,N_18228,N_18941);
nand U22196 (N_22196,N_19789,N_17500);
nor U22197 (N_22197,N_19641,N_18852);
and U22198 (N_22198,N_17646,N_18958);
or U22199 (N_22199,N_19966,N_17628);
nor U22200 (N_22200,N_17951,N_18093);
or U22201 (N_22201,N_19804,N_17623);
or U22202 (N_22202,N_19385,N_18846);
xor U22203 (N_22203,N_18592,N_17927);
nand U22204 (N_22204,N_19098,N_19534);
and U22205 (N_22205,N_17936,N_19800);
nor U22206 (N_22206,N_18366,N_19112);
and U22207 (N_22207,N_18761,N_17872);
nand U22208 (N_22208,N_17855,N_17990);
or U22209 (N_22209,N_17802,N_18041);
nor U22210 (N_22210,N_17902,N_17654);
nand U22211 (N_22211,N_19192,N_19212);
or U22212 (N_22212,N_18271,N_19788);
nor U22213 (N_22213,N_18280,N_19128);
or U22214 (N_22214,N_19721,N_18959);
nor U22215 (N_22215,N_19033,N_17554);
nand U22216 (N_22216,N_19441,N_18355);
nand U22217 (N_22217,N_18647,N_18298);
nor U22218 (N_22218,N_19614,N_17533);
and U22219 (N_22219,N_17762,N_18392);
or U22220 (N_22220,N_17907,N_19884);
nor U22221 (N_22221,N_18895,N_19867);
nand U22222 (N_22222,N_18864,N_17893);
nand U22223 (N_22223,N_18761,N_19232);
or U22224 (N_22224,N_18714,N_19629);
or U22225 (N_22225,N_19504,N_19624);
or U22226 (N_22226,N_19501,N_19974);
nand U22227 (N_22227,N_19268,N_18691);
or U22228 (N_22228,N_18211,N_18664);
nand U22229 (N_22229,N_17547,N_19309);
nand U22230 (N_22230,N_17946,N_18696);
nand U22231 (N_22231,N_19574,N_18591);
xor U22232 (N_22232,N_18010,N_17591);
nor U22233 (N_22233,N_19665,N_19097);
nor U22234 (N_22234,N_17803,N_17919);
or U22235 (N_22235,N_19041,N_19661);
nor U22236 (N_22236,N_17627,N_19817);
or U22237 (N_22237,N_18857,N_17834);
nand U22238 (N_22238,N_17863,N_17616);
or U22239 (N_22239,N_17866,N_17741);
nor U22240 (N_22240,N_19178,N_18611);
nor U22241 (N_22241,N_18866,N_19024);
and U22242 (N_22242,N_19368,N_19183);
nand U22243 (N_22243,N_18425,N_17623);
or U22244 (N_22244,N_17602,N_19842);
nor U22245 (N_22245,N_18354,N_19260);
nor U22246 (N_22246,N_19245,N_17854);
or U22247 (N_22247,N_18134,N_18146);
and U22248 (N_22248,N_18213,N_19253);
nor U22249 (N_22249,N_17580,N_18383);
or U22250 (N_22250,N_19791,N_18511);
or U22251 (N_22251,N_17544,N_17664);
or U22252 (N_22252,N_19897,N_19213);
nand U22253 (N_22253,N_19070,N_18959);
and U22254 (N_22254,N_18489,N_19731);
or U22255 (N_22255,N_18046,N_19608);
and U22256 (N_22256,N_19758,N_19526);
and U22257 (N_22257,N_17502,N_18233);
nor U22258 (N_22258,N_18258,N_19164);
and U22259 (N_22259,N_17940,N_17918);
nor U22260 (N_22260,N_18195,N_18969);
nor U22261 (N_22261,N_19625,N_18314);
or U22262 (N_22262,N_19695,N_19729);
and U22263 (N_22263,N_18544,N_19052);
xnor U22264 (N_22264,N_18306,N_18013);
xnor U22265 (N_22265,N_18271,N_19193);
and U22266 (N_22266,N_19428,N_18771);
nor U22267 (N_22267,N_18602,N_19021);
or U22268 (N_22268,N_19514,N_19905);
and U22269 (N_22269,N_19720,N_19400);
or U22270 (N_22270,N_19719,N_18455);
and U22271 (N_22271,N_18353,N_19504);
nand U22272 (N_22272,N_18927,N_18817);
and U22273 (N_22273,N_18719,N_17581);
nand U22274 (N_22274,N_18938,N_18741);
xnor U22275 (N_22275,N_18891,N_17880);
and U22276 (N_22276,N_19591,N_19746);
or U22277 (N_22277,N_17653,N_19889);
xor U22278 (N_22278,N_19330,N_19357);
nor U22279 (N_22279,N_18753,N_19721);
xnor U22280 (N_22280,N_17743,N_19584);
nor U22281 (N_22281,N_18959,N_19317);
nor U22282 (N_22282,N_19280,N_19951);
xnor U22283 (N_22283,N_19387,N_17809);
nand U22284 (N_22284,N_19029,N_17955);
nor U22285 (N_22285,N_19718,N_19621);
nor U22286 (N_22286,N_19544,N_18315);
and U22287 (N_22287,N_18937,N_17559);
or U22288 (N_22288,N_17911,N_17987);
xor U22289 (N_22289,N_19232,N_19137);
or U22290 (N_22290,N_18515,N_19936);
or U22291 (N_22291,N_17867,N_19925);
nor U22292 (N_22292,N_19476,N_19402);
xor U22293 (N_22293,N_18150,N_17757);
nand U22294 (N_22294,N_17653,N_19159);
and U22295 (N_22295,N_17957,N_19831);
and U22296 (N_22296,N_17820,N_17546);
nand U22297 (N_22297,N_18337,N_19925);
and U22298 (N_22298,N_19545,N_19632);
nor U22299 (N_22299,N_19868,N_19360);
nor U22300 (N_22300,N_19519,N_18549);
and U22301 (N_22301,N_18962,N_17991);
and U22302 (N_22302,N_18669,N_17664);
or U22303 (N_22303,N_17782,N_18648);
or U22304 (N_22304,N_18655,N_19313);
nand U22305 (N_22305,N_17793,N_17670);
nand U22306 (N_22306,N_19259,N_19775);
or U22307 (N_22307,N_18712,N_19237);
and U22308 (N_22308,N_19390,N_18854);
xnor U22309 (N_22309,N_19446,N_19797);
nor U22310 (N_22310,N_18148,N_18443);
and U22311 (N_22311,N_19374,N_18769);
or U22312 (N_22312,N_17742,N_18122);
or U22313 (N_22313,N_18401,N_19662);
nor U22314 (N_22314,N_19878,N_18333);
or U22315 (N_22315,N_17527,N_19515);
and U22316 (N_22316,N_17891,N_17815);
nor U22317 (N_22317,N_18380,N_18809);
nand U22318 (N_22318,N_19536,N_19736);
or U22319 (N_22319,N_19608,N_18196);
and U22320 (N_22320,N_19416,N_18798);
xor U22321 (N_22321,N_19921,N_18533);
nor U22322 (N_22322,N_19492,N_18944);
and U22323 (N_22323,N_19045,N_19706);
nor U22324 (N_22324,N_18288,N_19267);
and U22325 (N_22325,N_18780,N_17666);
nor U22326 (N_22326,N_17719,N_18593);
or U22327 (N_22327,N_19154,N_19019);
and U22328 (N_22328,N_19096,N_18943);
or U22329 (N_22329,N_18303,N_18955);
and U22330 (N_22330,N_19896,N_17551);
or U22331 (N_22331,N_17907,N_19003);
and U22332 (N_22332,N_19089,N_19127);
or U22333 (N_22333,N_17768,N_18558);
nor U22334 (N_22334,N_19740,N_19036);
nor U22335 (N_22335,N_17725,N_19370);
and U22336 (N_22336,N_19620,N_19300);
nor U22337 (N_22337,N_18730,N_18969);
nand U22338 (N_22338,N_18983,N_17905);
nand U22339 (N_22339,N_17935,N_19660);
xnor U22340 (N_22340,N_18281,N_19967);
and U22341 (N_22341,N_18484,N_19709);
nand U22342 (N_22342,N_18781,N_19280);
and U22343 (N_22343,N_18874,N_19190);
or U22344 (N_22344,N_19057,N_19117);
nand U22345 (N_22345,N_17771,N_19622);
nor U22346 (N_22346,N_19472,N_17661);
nand U22347 (N_22347,N_17662,N_17714);
xor U22348 (N_22348,N_17688,N_17708);
nand U22349 (N_22349,N_17942,N_19276);
and U22350 (N_22350,N_17668,N_17793);
or U22351 (N_22351,N_17560,N_19434);
xnor U22352 (N_22352,N_18404,N_17526);
xor U22353 (N_22353,N_19352,N_19166);
nor U22354 (N_22354,N_19603,N_18663);
and U22355 (N_22355,N_18459,N_18762);
or U22356 (N_22356,N_18102,N_18275);
and U22357 (N_22357,N_18878,N_19109);
nand U22358 (N_22358,N_17878,N_18985);
nand U22359 (N_22359,N_19916,N_19927);
xor U22360 (N_22360,N_17525,N_18281);
and U22361 (N_22361,N_18102,N_19846);
xor U22362 (N_22362,N_18971,N_19701);
nor U22363 (N_22363,N_18238,N_19139);
and U22364 (N_22364,N_18170,N_19597);
nand U22365 (N_22365,N_18542,N_19119);
xnor U22366 (N_22366,N_18946,N_19875);
nor U22367 (N_22367,N_19769,N_18733);
nand U22368 (N_22368,N_19735,N_19320);
or U22369 (N_22369,N_18491,N_17656);
nand U22370 (N_22370,N_18894,N_19106);
or U22371 (N_22371,N_19331,N_19173);
and U22372 (N_22372,N_17661,N_18103);
nand U22373 (N_22373,N_18165,N_19041);
or U22374 (N_22374,N_18980,N_19326);
and U22375 (N_22375,N_19077,N_18613);
nor U22376 (N_22376,N_18052,N_17794);
nor U22377 (N_22377,N_18668,N_17905);
nor U22378 (N_22378,N_17600,N_19190);
xor U22379 (N_22379,N_19764,N_18032);
nor U22380 (N_22380,N_19487,N_17792);
or U22381 (N_22381,N_19286,N_19605);
and U22382 (N_22382,N_18112,N_19959);
nor U22383 (N_22383,N_19491,N_19026);
and U22384 (N_22384,N_19522,N_19156);
nand U22385 (N_22385,N_19008,N_18967);
or U22386 (N_22386,N_19282,N_19940);
and U22387 (N_22387,N_19315,N_18671);
xor U22388 (N_22388,N_19211,N_18049);
or U22389 (N_22389,N_18052,N_19256);
nor U22390 (N_22390,N_17977,N_18900);
or U22391 (N_22391,N_19952,N_19130);
nor U22392 (N_22392,N_19127,N_19616);
xnor U22393 (N_22393,N_18703,N_19115);
nand U22394 (N_22394,N_18754,N_19351);
and U22395 (N_22395,N_18517,N_17978);
and U22396 (N_22396,N_18983,N_19625);
or U22397 (N_22397,N_18858,N_19965);
nand U22398 (N_22398,N_17870,N_17951);
nor U22399 (N_22399,N_18298,N_18878);
and U22400 (N_22400,N_19782,N_18818);
nand U22401 (N_22401,N_19868,N_17946);
nor U22402 (N_22402,N_18006,N_18989);
nand U22403 (N_22403,N_18439,N_19969);
nor U22404 (N_22404,N_17603,N_18855);
xor U22405 (N_22405,N_17627,N_18848);
and U22406 (N_22406,N_19918,N_18319);
or U22407 (N_22407,N_19261,N_19013);
and U22408 (N_22408,N_19946,N_17606);
nand U22409 (N_22409,N_18302,N_18922);
and U22410 (N_22410,N_18604,N_19114);
or U22411 (N_22411,N_17903,N_18520);
and U22412 (N_22412,N_19149,N_18959);
nand U22413 (N_22413,N_19695,N_18485);
and U22414 (N_22414,N_17604,N_17833);
nand U22415 (N_22415,N_19854,N_19773);
nor U22416 (N_22416,N_18966,N_19562);
nand U22417 (N_22417,N_17994,N_19639);
or U22418 (N_22418,N_18522,N_18962);
nand U22419 (N_22419,N_17739,N_18069);
nor U22420 (N_22420,N_19852,N_17553);
and U22421 (N_22421,N_18239,N_19227);
nor U22422 (N_22422,N_19725,N_19426);
xor U22423 (N_22423,N_18666,N_19041);
nand U22424 (N_22424,N_19590,N_18185);
and U22425 (N_22425,N_19915,N_19574);
nor U22426 (N_22426,N_17867,N_18014);
nor U22427 (N_22427,N_19245,N_17585);
and U22428 (N_22428,N_18960,N_17622);
or U22429 (N_22429,N_18172,N_19280);
or U22430 (N_22430,N_18284,N_19861);
or U22431 (N_22431,N_19011,N_17511);
or U22432 (N_22432,N_17964,N_18737);
or U22433 (N_22433,N_18946,N_18233);
nor U22434 (N_22434,N_19935,N_18116);
or U22435 (N_22435,N_19974,N_18861);
nand U22436 (N_22436,N_19212,N_19762);
and U22437 (N_22437,N_18542,N_19466);
nor U22438 (N_22438,N_19981,N_17923);
and U22439 (N_22439,N_18143,N_19890);
and U22440 (N_22440,N_17796,N_19282);
nor U22441 (N_22441,N_17831,N_19585);
nand U22442 (N_22442,N_18854,N_17699);
or U22443 (N_22443,N_18260,N_19059);
nor U22444 (N_22444,N_18124,N_19311);
nor U22445 (N_22445,N_18740,N_19925);
or U22446 (N_22446,N_18886,N_18141);
nand U22447 (N_22447,N_18921,N_17834);
nand U22448 (N_22448,N_18341,N_17859);
nor U22449 (N_22449,N_18227,N_18893);
or U22450 (N_22450,N_18082,N_18456);
and U22451 (N_22451,N_18604,N_19773);
xnor U22452 (N_22452,N_19378,N_19238);
nand U22453 (N_22453,N_17728,N_19796);
and U22454 (N_22454,N_19714,N_18341);
or U22455 (N_22455,N_18962,N_18674);
xor U22456 (N_22456,N_17724,N_19501);
or U22457 (N_22457,N_18058,N_19093);
nor U22458 (N_22458,N_18706,N_17865);
or U22459 (N_22459,N_19960,N_17564);
nor U22460 (N_22460,N_19602,N_18473);
nand U22461 (N_22461,N_17937,N_18639);
nor U22462 (N_22462,N_18036,N_17638);
and U22463 (N_22463,N_19275,N_18308);
and U22464 (N_22464,N_18989,N_19045);
or U22465 (N_22465,N_17640,N_19386);
and U22466 (N_22466,N_17555,N_19767);
and U22467 (N_22467,N_19899,N_18508);
or U22468 (N_22468,N_18524,N_19740);
nor U22469 (N_22469,N_19915,N_18325);
or U22470 (N_22470,N_19580,N_18082);
xnor U22471 (N_22471,N_18885,N_19711);
and U22472 (N_22472,N_17835,N_18583);
and U22473 (N_22473,N_18112,N_18187);
and U22474 (N_22474,N_19023,N_17546);
and U22475 (N_22475,N_18148,N_19419);
nand U22476 (N_22476,N_19144,N_18054);
and U22477 (N_22477,N_19843,N_17697);
nor U22478 (N_22478,N_18010,N_19312);
and U22479 (N_22479,N_19942,N_19902);
nor U22480 (N_22480,N_18549,N_17804);
or U22481 (N_22481,N_19686,N_19351);
or U22482 (N_22482,N_18888,N_19045);
and U22483 (N_22483,N_18298,N_18245);
nand U22484 (N_22484,N_19602,N_19628);
nand U22485 (N_22485,N_19337,N_18353);
and U22486 (N_22486,N_18361,N_17710);
or U22487 (N_22487,N_19849,N_19602);
xor U22488 (N_22488,N_18144,N_17509);
and U22489 (N_22489,N_18287,N_18348);
and U22490 (N_22490,N_18293,N_18514);
nor U22491 (N_22491,N_19506,N_18276);
or U22492 (N_22492,N_18521,N_17993);
nor U22493 (N_22493,N_18457,N_19632);
nor U22494 (N_22494,N_19944,N_17580);
nor U22495 (N_22495,N_18484,N_17622);
and U22496 (N_22496,N_17887,N_18923);
nand U22497 (N_22497,N_18231,N_19116);
nor U22498 (N_22498,N_19523,N_18221);
and U22499 (N_22499,N_19895,N_18167);
nor U22500 (N_22500,N_20725,N_21085);
nor U22501 (N_22501,N_21653,N_20738);
nor U22502 (N_22502,N_20992,N_20258);
nand U22503 (N_22503,N_22249,N_20612);
or U22504 (N_22504,N_20899,N_20650);
nor U22505 (N_22505,N_21893,N_21527);
or U22506 (N_22506,N_21853,N_20931);
and U22507 (N_22507,N_21815,N_20752);
nand U22508 (N_22508,N_20056,N_21420);
and U22509 (N_22509,N_22120,N_21160);
nor U22510 (N_22510,N_20771,N_20812);
nor U22511 (N_22511,N_20292,N_21433);
nand U22512 (N_22512,N_22124,N_21203);
or U22513 (N_22513,N_20526,N_20522);
xor U22514 (N_22514,N_21065,N_21421);
or U22515 (N_22515,N_21022,N_21621);
nor U22516 (N_22516,N_22070,N_21905);
nor U22517 (N_22517,N_20614,N_21238);
or U22518 (N_22518,N_22129,N_21775);
and U22519 (N_22519,N_21196,N_22486);
and U22520 (N_22520,N_20129,N_22349);
nand U22521 (N_22521,N_21016,N_22481);
or U22522 (N_22522,N_21828,N_20348);
nand U22523 (N_22523,N_21228,N_22004);
nand U22524 (N_22524,N_21365,N_21147);
nand U22525 (N_22525,N_20610,N_21895);
nor U22526 (N_22526,N_20722,N_22334);
or U22527 (N_22527,N_21391,N_21481);
xnor U22528 (N_22528,N_21530,N_20824);
nor U22529 (N_22529,N_22472,N_21441);
xor U22530 (N_22530,N_20030,N_20334);
nand U22531 (N_22531,N_20884,N_20418);
and U22532 (N_22532,N_21747,N_22188);
nor U22533 (N_22533,N_21865,N_22400);
xnor U22534 (N_22534,N_20822,N_21823);
or U22535 (N_22535,N_20973,N_21835);
or U22536 (N_22536,N_21353,N_22321);
and U22537 (N_22537,N_21418,N_21956);
or U22538 (N_22538,N_22235,N_20131);
or U22539 (N_22539,N_21998,N_21126);
xor U22540 (N_22540,N_21002,N_20595);
nor U22541 (N_22541,N_21807,N_21327);
or U22542 (N_22542,N_20215,N_20376);
nand U22543 (N_22543,N_20353,N_21115);
nor U22544 (N_22544,N_21920,N_22167);
nand U22545 (N_22545,N_21382,N_21061);
nand U22546 (N_22546,N_22408,N_20568);
nand U22547 (N_22547,N_22485,N_20281);
xnor U22548 (N_22548,N_20659,N_21487);
nor U22549 (N_22549,N_21681,N_20489);
and U22550 (N_22550,N_20091,N_21965);
xor U22551 (N_22551,N_21741,N_20318);
and U22552 (N_22552,N_21960,N_20816);
xor U22553 (N_22553,N_20772,N_20949);
nand U22554 (N_22554,N_22051,N_21825);
xor U22555 (N_22555,N_20905,N_20036);
nand U22556 (N_22556,N_20502,N_20354);
nand U22557 (N_22557,N_21518,N_21915);
and U22558 (N_22558,N_22148,N_20809);
nand U22559 (N_22559,N_22060,N_21068);
nor U22560 (N_22560,N_22134,N_21975);
or U22561 (N_22561,N_20068,N_20955);
nand U22562 (N_22562,N_20564,N_20803);
nand U22563 (N_22563,N_21767,N_22231);
nand U22564 (N_22564,N_20927,N_20245);
nor U22565 (N_22565,N_22115,N_22064);
nand U22566 (N_22566,N_22108,N_21885);
nor U22567 (N_22567,N_20061,N_20369);
and U22568 (N_22568,N_21523,N_21706);
or U22569 (N_22569,N_20415,N_20236);
xnor U22570 (N_22570,N_20022,N_22147);
or U22571 (N_22571,N_22384,N_21982);
nand U22572 (N_22572,N_21058,N_20073);
nand U22573 (N_22573,N_22368,N_20041);
or U22574 (N_22574,N_20575,N_20921);
nand U22575 (N_22575,N_20422,N_21964);
or U22576 (N_22576,N_20550,N_21641);
or U22577 (N_22577,N_20923,N_20984);
nor U22578 (N_22578,N_20027,N_21508);
and U22579 (N_22579,N_22047,N_22221);
or U22580 (N_22580,N_21654,N_20207);
nand U22581 (N_22581,N_21799,N_20876);
and U22582 (N_22582,N_21231,N_21473);
nand U22583 (N_22583,N_22048,N_21232);
or U22584 (N_22584,N_20565,N_21661);
nor U22585 (N_22585,N_22256,N_21243);
or U22586 (N_22586,N_21580,N_21242);
xor U22587 (N_22587,N_22431,N_20203);
xnor U22588 (N_22588,N_21038,N_22094);
or U22589 (N_22589,N_21412,N_21858);
nand U22590 (N_22590,N_20278,N_21644);
xnor U22591 (N_22591,N_21843,N_21628);
nor U22592 (N_22592,N_20101,N_21097);
or U22593 (N_22593,N_20491,N_21632);
or U22594 (N_22594,N_21648,N_22195);
or U22595 (N_22595,N_22420,N_21376);
and U22596 (N_22596,N_21652,N_20587);
and U22597 (N_22597,N_21601,N_20238);
and U22598 (N_22598,N_22117,N_20501);
or U22599 (N_22599,N_20226,N_22203);
nand U22600 (N_22600,N_22340,N_21503);
and U22601 (N_22601,N_20898,N_20753);
or U22602 (N_22602,N_22190,N_20727);
and U22603 (N_22603,N_20531,N_21875);
nor U22604 (N_22604,N_20500,N_22456);
or U22605 (N_22605,N_21897,N_20607);
and U22606 (N_22606,N_22322,N_21080);
or U22607 (N_22607,N_20558,N_21860);
or U22608 (N_22608,N_21098,N_21674);
or U22609 (N_22609,N_20189,N_20441);
xnor U22610 (N_22610,N_21261,N_21139);
nand U22611 (N_22611,N_21864,N_21151);
or U22612 (N_22612,N_20616,N_20833);
nor U22613 (N_22613,N_22437,N_22397);
nand U22614 (N_22614,N_20112,N_21223);
or U22615 (N_22615,N_22191,N_21245);
nand U22616 (N_22616,N_20970,N_22106);
or U22617 (N_22617,N_21755,N_20944);
nor U22618 (N_22618,N_20217,N_20104);
nand U22619 (N_22619,N_20434,N_20414);
or U22620 (N_22620,N_20581,N_20083);
nand U22621 (N_22621,N_21439,N_22435);
nor U22622 (N_22622,N_21230,N_21142);
nor U22623 (N_22623,N_20461,N_20031);
or U22624 (N_22624,N_22434,N_20052);
nor U22625 (N_22625,N_22404,N_20724);
or U22626 (N_22626,N_21318,N_20551);
nor U22627 (N_22627,N_20026,N_20887);
or U22628 (N_22628,N_20508,N_20473);
xnor U22629 (N_22629,N_20689,N_22197);
and U22630 (N_22630,N_20187,N_21795);
xnor U22631 (N_22631,N_21338,N_22163);
nor U22632 (N_22632,N_20947,N_21673);
and U22633 (N_22633,N_20483,N_22499);
nand U22634 (N_22634,N_20846,N_20227);
or U22635 (N_22635,N_21761,N_20696);
or U22636 (N_22636,N_22255,N_20155);
xor U22637 (N_22637,N_21409,N_21256);
and U22638 (N_22638,N_21526,N_22479);
and U22639 (N_22639,N_20065,N_21994);
nor U22640 (N_22640,N_20467,N_20021);
nor U22641 (N_22641,N_20169,N_22475);
nor U22642 (N_22642,N_20957,N_20832);
or U22643 (N_22643,N_21943,N_21346);
and U22644 (N_22644,N_21546,N_21645);
and U22645 (N_22645,N_22265,N_21449);
nor U22646 (N_22646,N_21562,N_22492);
nand U22647 (N_22647,N_20045,N_21325);
nor U22648 (N_22648,N_21286,N_22450);
xor U22649 (N_22649,N_21172,N_22263);
and U22650 (N_22650,N_20746,N_20372);
or U22651 (N_22651,N_22044,N_21406);
or U22652 (N_22652,N_20020,N_22280);
nor U22653 (N_22653,N_22429,N_21818);
and U22654 (N_22654,N_20745,N_22339);
and U22655 (N_22655,N_21600,N_21754);
and U22656 (N_22656,N_21079,N_22127);
and U22657 (N_22657,N_22457,N_20302);
nor U22658 (N_22658,N_21519,N_22385);
and U22659 (N_22659,N_20982,N_20256);
or U22660 (N_22660,N_20769,N_21572);
or U22661 (N_22661,N_22053,N_21194);
nor U22662 (N_22662,N_21703,N_20147);
or U22663 (N_22663,N_21205,N_20509);
and U22664 (N_22664,N_22013,N_21619);
nand U22665 (N_22665,N_20239,N_21395);
nor U22666 (N_22666,N_20929,N_22310);
nor U22667 (N_22667,N_20464,N_20493);
and U22668 (N_22668,N_21919,N_20795);
and U22669 (N_22669,N_20057,N_22449);
nand U22670 (N_22670,N_21783,N_20794);
or U22671 (N_22671,N_21640,N_20828);
xor U22672 (N_22672,N_21396,N_20845);
nand U22673 (N_22673,N_20181,N_21590);
nor U22674 (N_22674,N_20225,N_21564);
nand U22675 (N_22675,N_21266,N_22315);
nor U22676 (N_22676,N_21390,N_22110);
nor U22677 (N_22677,N_20210,N_20413);
and U22678 (N_22678,N_21587,N_22024);
nor U22679 (N_22679,N_20174,N_20628);
or U22680 (N_22680,N_21131,N_20760);
nor U22681 (N_22681,N_21760,N_21124);
and U22682 (N_22682,N_20471,N_22482);
xnor U22683 (N_22683,N_21350,N_21343);
and U22684 (N_22684,N_20252,N_22181);
nor U22685 (N_22685,N_21907,N_21101);
nand U22686 (N_22686,N_22058,N_20841);
nor U22687 (N_22687,N_21471,N_20907);
xor U22688 (N_22688,N_21127,N_21303);
nand U22689 (N_22689,N_20591,N_21105);
nor U22690 (N_22690,N_22411,N_20634);
and U22691 (N_22691,N_20019,N_22031);
and U22692 (N_22692,N_20578,N_20946);
nor U22693 (N_22693,N_22378,N_20934);
or U22694 (N_22694,N_20665,N_21725);
or U22695 (N_22695,N_22264,N_21272);
nor U22696 (N_22696,N_21077,N_20266);
or U22697 (N_22697,N_21557,N_21593);
and U22698 (N_22698,N_21153,N_22291);
nor U22699 (N_22699,N_21241,N_20664);
or U22700 (N_22700,N_21432,N_22209);
nand U22701 (N_22701,N_20316,N_21944);
or U22702 (N_22702,N_20865,N_21647);
nor U22703 (N_22703,N_21234,N_20685);
or U22704 (N_22704,N_21485,N_21798);
or U22705 (N_22705,N_21597,N_21890);
nand U22706 (N_22706,N_20254,N_21163);
nor U22707 (N_22707,N_20836,N_22414);
and U22708 (N_22708,N_20557,N_20098);
and U22709 (N_22709,N_20228,N_20968);
and U22710 (N_22710,N_21586,N_20494);
or U22711 (N_22711,N_22219,N_20917);
or U22712 (N_22712,N_21227,N_20244);
xnor U22713 (N_22713,N_21235,N_21870);
and U22714 (N_22714,N_21633,N_20524);
nand U22715 (N_22715,N_20247,N_21239);
nor U22716 (N_22716,N_20279,N_21214);
and U22717 (N_22717,N_21181,N_21033);
and U22718 (N_22718,N_20123,N_22307);
and U22719 (N_22719,N_21082,N_20620);
nor U22720 (N_22720,N_20343,N_21334);
nor U22721 (N_22721,N_20590,N_22158);
and U22722 (N_22722,N_22098,N_21400);
and U22723 (N_22723,N_21695,N_22443);
or U22724 (N_22724,N_21903,N_20773);
nand U22725 (N_22725,N_20511,N_20100);
nor U22726 (N_22726,N_21682,N_22401);
xor U22727 (N_22727,N_22306,N_22049);
nor U22728 (N_22728,N_22471,N_21615);
nor U22729 (N_22729,N_22377,N_22463);
or U22730 (N_22730,N_20023,N_20837);
nand U22731 (N_22731,N_20459,N_21066);
nor U22732 (N_22732,N_21307,N_22005);
nand U22733 (N_22733,N_20864,N_20149);
or U22734 (N_22734,N_20417,N_21490);
xor U22735 (N_22735,N_21934,N_21800);
nand U22736 (N_22736,N_21422,N_20867);
or U22737 (N_22737,N_21871,N_20806);
or U22738 (N_22738,N_20048,N_21697);
nor U22739 (N_22739,N_20919,N_20894);
nand U22740 (N_22740,N_20838,N_21591);
xnor U22741 (N_22741,N_20213,N_22393);
and U22742 (N_22742,N_22412,N_22067);
or U22743 (N_22743,N_21347,N_20014);
and U22744 (N_22744,N_20477,N_20719);
and U22745 (N_22745,N_21457,N_20965);
and U22746 (N_22746,N_22373,N_21083);
or U22747 (N_22747,N_21112,N_20580);
or U22748 (N_22748,N_20851,N_21824);
nor U22749 (N_22749,N_20862,N_20148);
nor U22750 (N_22750,N_22179,N_22489);
xor U22751 (N_22751,N_20054,N_20078);
xnor U22752 (N_22752,N_21474,N_21100);
or U22753 (N_22753,N_21510,N_20647);
nand U22754 (N_22754,N_20438,N_21056);
nor U22755 (N_22755,N_22097,N_21699);
nand U22756 (N_22756,N_21938,N_21972);
and U22757 (N_22757,N_22346,N_20700);
or U22758 (N_22758,N_21357,N_20920);
nand U22759 (N_22759,N_22442,N_20089);
nand U22760 (N_22760,N_20962,N_21207);
nand U22761 (N_22761,N_22017,N_20662);
nand U22762 (N_22762,N_20562,N_21442);
or U22763 (N_22763,N_20151,N_21069);
nand U22764 (N_22764,N_20111,N_22348);
nand U22765 (N_22765,N_21354,N_21846);
nor U22766 (N_22766,N_20260,N_20945);
or U22767 (N_22767,N_20287,N_21727);
nand U22768 (N_22768,N_20042,N_22079);
or U22769 (N_22769,N_21852,N_20517);
xnor U22770 (N_22770,N_20407,N_20781);
xnor U22771 (N_22771,N_20701,N_21876);
or U22772 (N_22772,N_20288,N_22016);
and U22773 (N_22773,N_22011,N_22381);
and U22774 (N_22774,N_21551,N_21678);
nand U22775 (N_22775,N_20886,N_21090);
nand U22776 (N_22776,N_20063,N_20212);
or U22777 (N_22777,N_20709,N_20704);
nand U22778 (N_22778,N_21448,N_20999);
xor U22779 (N_22779,N_21296,N_21504);
and U22780 (N_22780,N_21957,N_21847);
nor U22781 (N_22781,N_21773,N_20125);
nor U22782 (N_22782,N_22232,N_20879);
or U22783 (N_22783,N_22313,N_22374);
or U22784 (N_22784,N_20322,N_21025);
nand U22785 (N_22785,N_21009,N_21463);
nand U22786 (N_22786,N_21219,N_22239);
xor U22787 (N_22787,N_20566,N_20536);
and U22788 (N_22788,N_22359,N_22211);
or U22789 (N_22789,N_20901,N_21675);
nor U22790 (N_22790,N_21281,N_20615);
nand U22791 (N_22791,N_21001,N_22193);
nor U22792 (N_22792,N_21169,N_20544);
nand U22793 (N_22793,N_21686,N_20224);
and U22794 (N_22794,N_21381,N_22074);
or U22795 (N_22795,N_21277,N_22091);
and U22796 (N_22796,N_20788,N_22151);
nand U22797 (N_22797,N_22216,N_20191);
nand U22798 (N_22798,N_20394,N_20309);
and U22799 (N_22799,N_20485,N_21225);
or U22800 (N_22800,N_22297,N_22152);
nor U22801 (N_22801,N_21541,N_22099);
nand U22802 (N_22802,N_21348,N_22062);
or U22803 (N_22803,N_22427,N_22065);
xnor U22804 (N_22804,N_20525,N_20240);
nor U22805 (N_22805,N_20641,N_21693);
nor U22806 (N_22806,N_20644,N_21435);
nor U22807 (N_22807,N_22391,N_22498);
and U22808 (N_22808,N_21547,N_21055);
nor U22809 (N_22809,N_21556,N_21826);
nor U22810 (N_22810,N_20116,N_22462);
nand U22811 (N_22811,N_20114,N_20296);
nand U22812 (N_22812,N_21622,N_20430);
or U22813 (N_22813,N_20390,N_21466);
and U22814 (N_22814,N_20034,N_21739);
nand U22815 (N_22815,N_21469,N_21484);
or U22816 (N_22816,N_20642,N_20423);
and U22817 (N_22817,N_21866,N_21195);
xor U22818 (N_22818,N_21947,N_20363);
nor U22819 (N_22819,N_20472,N_20003);
or U22820 (N_22820,N_20675,N_22260);
nand U22821 (N_22821,N_22003,N_20231);
nor U22822 (N_22822,N_20409,N_22220);
nand U22823 (N_22823,N_20950,N_20202);
nor U22824 (N_22824,N_21293,N_22171);
or U22825 (N_22825,N_21408,N_21494);
nand U22826 (N_22826,N_20691,N_21575);
and U22827 (N_22827,N_22447,N_22465);
nor U22828 (N_22828,N_20830,N_20420);
nand U22829 (N_22829,N_21385,N_22476);
or U22830 (N_22830,N_20697,N_20000);
or U22831 (N_22831,N_21094,N_20963);
xor U22832 (N_22832,N_22363,N_22009);
nand U22833 (N_22833,N_21887,N_22236);
nand U22834 (N_22834,N_21657,N_21087);
xor U22835 (N_22835,N_20776,N_20184);
or U22836 (N_22836,N_20732,N_20756);
nand U22837 (N_22837,N_20117,N_22298);
nor U22838 (N_22838,N_22269,N_20305);
and U22839 (N_22839,N_20314,N_20142);
nor U22840 (N_22840,N_20016,N_21149);
nand U22841 (N_22841,N_20759,N_20855);
nor U22842 (N_22842,N_21283,N_22105);
nor U22843 (N_22843,N_21612,N_21255);
or U22844 (N_22844,N_20011,N_22444);
and U22845 (N_22845,N_20956,N_21176);
nor U22846 (N_22846,N_22080,N_20113);
and U22847 (N_22847,N_21446,N_21140);
or U22848 (N_22848,N_20790,N_21499);
and U22849 (N_22849,N_21561,N_20182);
nand U22850 (N_22850,N_21380,N_21788);
nor U22851 (N_22851,N_20396,N_22361);
and U22852 (N_22852,N_20345,N_20145);
nand U22853 (N_22853,N_21273,N_20718);
nor U22854 (N_22854,N_20835,N_20119);
or U22855 (N_22855,N_20969,N_22036);
nor U22856 (N_22856,N_21869,N_21425);
nand U22857 (N_22857,N_21936,N_22213);
and U22858 (N_22858,N_22273,N_22208);
nand U22859 (N_22859,N_20633,N_21260);
xnor U22860 (N_22860,N_20850,N_21121);
nor U22861 (N_22861,N_22281,N_20482);
and U22862 (N_22862,N_21766,N_21053);
nor U22863 (N_22863,N_21392,N_20938);
nand U22864 (N_22864,N_21117,N_22078);
nor U22865 (N_22865,N_20916,N_20922);
or U22866 (N_22866,N_21662,N_21049);
and U22867 (N_22867,N_21356,N_22439);
xnor U22868 (N_22868,N_20943,N_20687);
or U22869 (N_22869,N_22039,N_20271);
xnor U22870 (N_22870,N_20930,N_20975);
nand U22871 (N_22871,N_20402,N_20754);
nor U22872 (N_22872,N_20527,N_21712);
or U22873 (N_22873,N_22386,N_21596);
and U22874 (N_22874,N_20053,N_22480);
nand U22875 (N_22875,N_21922,N_20540);
or U22876 (N_22876,N_21554,N_20713);
xnor U22877 (N_22877,N_21148,N_20455);
xnor U22878 (N_22878,N_20072,N_20454);
or U22879 (N_22879,N_20342,N_21417);
nand U22880 (N_22880,N_21709,N_20044);
nor U22881 (N_22881,N_20387,N_21537);
and U22882 (N_22882,N_20802,N_22103);
and U22883 (N_22883,N_21029,N_22183);
and U22884 (N_22884,N_20810,N_22387);
or U22885 (N_22885,N_20842,N_20731);
and U22886 (N_22886,N_20115,N_21034);
nand U22887 (N_22887,N_20421,N_21040);
and U22888 (N_22888,N_21093,N_20883);
nand U22889 (N_22889,N_22246,N_20737);
nor U22890 (N_22890,N_20002,N_21208);
and U22891 (N_22891,N_20774,N_20630);
xnor U22892 (N_22892,N_21521,N_20621);
nor U22893 (N_22893,N_21777,N_21691);
or U22894 (N_22894,N_21249,N_22154);
nand U22895 (N_22895,N_20428,N_20941);
nand U22896 (N_22896,N_22248,N_20601);
and U22897 (N_22897,N_20519,N_21758);
and U22898 (N_22898,N_20286,N_20678);
or U22899 (N_22899,N_20077,N_21041);
nand U22900 (N_22900,N_22371,N_20154);
nand U22901 (N_22901,N_22304,N_20338);
and U22902 (N_22902,N_21031,N_20672);
nor U22903 (N_22903,N_22354,N_21584);
nand U22904 (N_22904,N_20029,N_20074);
and U22905 (N_22905,N_20723,N_21954);
nor U22906 (N_22906,N_22125,N_20033);
and U22907 (N_22907,N_21577,N_22112);
and U22908 (N_22908,N_20896,N_21779);
xnor U22909 (N_22909,N_20889,N_21375);
and U22910 (N_22910,N_20152,N_20495);
nand U22911 (N_22911,N_21573,N_22177);
and U22912 (N_22912,N_22076,N_20751);
and U22913 (N_22913,N_20295,N_20070);
or U22914 (N_22914,N_21458,N_20199);
or U22915 (N_22915,N_21282,N_21180);
nor U22916 (N_22916,N_21290,N_21899);
and U22917 (N_22917,N_22415,N_21827);
or U22918 (N_22918,N_20598,N_21862);
nand U22919 (N_22919,N_21339,N_20470);
nor U22920 (N_22920,N_20206,N_20677);
xor U22921 (N_22921,N_20168,N_22162);
nor U22922 (N_22922,N_21901,N_22233);
nand U22923 (N_22923,N_20503,N_22182);
and U22924 (N_22924,N_20284,N_20593);
or U22925 (N_22925,N_21088,N_22137);
and U22926 (N_22926,N_20843,N_21292);
and U22927 (N_22927,N_22460,N_21776);
or U22928 (N_22928,N_21660,N_21078);
nor U22929 (N_22929,N_21091,N_22336);
nor U22930 (N_22930,N_22285,N_20624);
or U22931 (N_22931,N_21840,N_20408);
nand U22932 (N_22932,N_21679,N_21845);
nand U22933 (N_22933,N_21752,N_20280);
nor U22934 (N_22934,N_21134,N_21789);
xnor U22935 (N_22935,N_20162,N_20577);
nor U22936 (N_22936,N_21770,N_20690);
nor U22937 (N_22937,N_21329,N_20216);
and U22938 (N_22938,N_20748,N_22464);
nand U22939 (N_22939,N_21553,N_20868);
or U22940 (N_22940,N_20561,N_21921);
nor U22941 (N_22941,N_21851,N_22376);
xnor U22942 (N_22942,N_22185,N_20733);
nand U22943 (N_22943,N_22274,N_21796);
nand U22944 (N_22944,N_20611,N_20966);
and U22945 (N_22945,N_20646,N_21206);
or U22946 (N_22946,N_22063,N_20903);
xnor U22947 (N_22947,N_20375,N_21200);
xor U22948 (N_22948,N_21162,N_21625);
xor U22949 (N_22949,N_21762,N_22253);
and U22950 (N_22950,N_22095,N_22261);
and U22951 (N_22951,N_21962,N_20613);
nor U22952 (N_22952,N_20234,N_20456);
or U22953 (N_22953,N_22165,N_20469);
nand U22954 (N_22954,N_21304,N_20859);
and U22955 (N_22955,N_21374,N_21403);
and U22956 (N_22956,N_22325,N_21413);
xnor U22957 (N_22957,N_22490,N_22228);
nor U22958 (N_22958,N_21774,N_21443);
and U22959 (N_22959,N_22319,N_21778);
nor U22960 (N_22960,N_20599,N_21387);
and U22961 (N_22961,N_20437,N_20259);
and U22962 (N_22962,N_20787,N_21438);
and U22963 (N_22963,N_20272,N_20444);
and U22964 (N_22964,N_20253,N_21585);
nor U22965 (N_22965,N_21427,N_22136);
nor U22966 (N_22966,N_22242,N_22367);
nand U22967 (N_22967,N_20386,N_20431);
nand U22968 (N_22968,N_22201,N_22335);
or U22969 (N_22969,N_21945,N_20783);
nand U22970 (N_22970,N_21880,N_20711);
nor U22971 (N_22971,N_22172,N_21589);
and U22972 (N_22972,N_20103,N_20433);
or U22973 (N_22973,N_22317,N_21459);
nand U22974 (N_22974,N_21917,N_20392);
or U22975 (N_22975,N_21174,N_21863);
or U22976 (N_22976,N_20827,N_22296);
and U22977 (N_22977,N_21440,N_20986);
or U22978 (N_22978,N_21700,N_22487);
nor U22979 (N_22979,N_21159,N_21311);
or U22980 (N_22980,N_20734,N_21616);
xnor U22981 (N_22981,N_20983,N_21737);
and U22982 (N_22982,N_20172,N_21096);
xor U22983 (N_22983,N_20312,N_20574);
and U22984 (N_22984,N_21184,N_22215);
nand U22985 (N_22985,N_21372,N_21842);
or U22986 (N_22986,N_21516,N_22075);
nor U22987 (N_22987,N_20136,N_21909);
nand U22988 (N_22988,N_20233,N_22250);
nand U22989 (N_22989,N_21992,N_21328);
and U22990 (N_22990,N_21434,N_21003);
or U22991 (N_22991,N_20506,N_20750);
and U22992 (N_22992,N_21394,N_22392);
or U22993 (N_22993,N_22175,N_21305);
and U22994 (N_22994,N_21059,N_20877);
nor U22995 (N_22995,N_20825,N_21849);
xnor U22996 (N_22996,N_22284,N_21081);
and U22997 (N_22997,N_21502,N_21896);
nor U22998 (N_22998,N_20798,N_20359);
nor U22999 (N_22999,N_20320,N_22308);
or U23000 (N_23000,N_22252,N_20398);
xor U23001 (N_23001,N_20671,N_20617);
or U23002 (N_23002,N_20608,N_20121);
nor U23003 (N_23003,N_21211,N_20171);
and U23004 (N_23004,N_21006,N_22332);
and U23005 (N_23005,N_21550,N_22012);
nor U23006 (N_23006,N_21941,N_21705);
nor U23007 (N_23007,N_20270,N_21300);
nand U23008 (N_23008,N_20736,N_20940);
or U23009 (N_23009,N_20870,N_21488);
and U23010 (N_23010,N_21658,N_20958);
or U23011 (N_23011,N_20758,N_21734);
or U23012 (N_23012,N_21341,N_22345);
and U23013 (N_23013,N_21780,N_20127);
and U23014 (N_23014,N_20261,N_21614);
nand U23015 (N_23015,N_20241,N_21419);
nand U23016 (N_23016,N_20784,N_21900);
nor U23017 (N_23017,N_21782,N_21592);
nand U23018 (N_23018,N_22350,N_21367);
nor U23019 (N_23019,N_20972,N_21017);
or U23020 (N_23020,N_20767,N_22425);
nor U23021 (N_23021,N_21386,N_20847);
nor U23022 (N_23022,N_22093,N_21405);
nor U23023 (N_23023,N_21319,N_21076);
nor U23024 (N_23024,N_20676,N_22041);
or U23025 (N_23025,N_20173,N_21216);
xor U23026 (N_23026,N_20514,N_20277);
and U23027 (N_23027,N_21460,N_21113);
nor U23028 (N_23028,N_20596,N_20282);
and U23029 (N_23029,N_20357,N_20352);
nand U23030 (N_23030,N_21465,N_21721);
and U23031 (N_23031,N_21771,N_21287);
and U23032 (N_23032,N_20635,N_21170);
nor U23033 (N_23033,N_21244,N_22069);
or U23034 (N_23034,N_21210,N_20902);
nand U23035 (N_23035,N_22022,N_21642);
nor U23036 (N_23036,N_21224,N_21110);
nor U23037 (N_23037,N_21809,N_20143);
and U23038 (N_23038,N_22406,N_20925);
nor U23039 (N_23039,N_22038,N_21209);
and U23040 (N_23040,N_21985,N_20449);
nand U23041 (N_23041,N_21804,N_21685);
nand U23042 (N_23042,N_22337,N_20761);
and U23043 (N_23043,N_21738,N_20977);
nand U23044 (N_23044,N_22417,N_20716);
or U23045 (N_23045,N_22294,N_21717);
and U23046 (N_23046,N_20668,N_21963);
and U23047 (N_23047,N_22477,N_21968);
nor U23048 (N_23048,N_21988,N_21588);
and U23049 (N_23049,N_21568,N_20051);
xnor U23050 (N_23050,N_21916,N_22204);
xor U23051 (N_23051,N_21155,N_21878);
or U23052 (N_23052,N_20443,N_21611);
and U23053 (N_23053,N_21051,N_20404);
nor U23054 (N_23054,N_21233,N_21733);
nand U23055 (N_23055,N_22085,N_20448);
xnor U23056 (N_23056,N_21102,N_21522);
nand U23057 (N_23057,N_21298,N_20328);
and U23058 (N_23058,N_20128,N_21882);
nor U23059 (N_23059,N_22369,N_20323);
and U23060 (N_23060,N_22035,N_20487);
nor U23061 (N_23061,N_20584,N_21447);
nand U23062 (N_23062,N_20450,N_20344);
and U23063 (N_23063,N_21759,N_22276);
nand U23064 (N_23064,N_20218,N_20311);
and U23065 (N_23065,N_21784,N_20012);
or U23066 (N_23066,N_21750,N_21745);
nand U23067 (N_23067,N_21315,N_21064);
nor U23068 (N_23068,N_21047,N_20710);
and U23069 (N_23069,N_20988,N_22370);
nor U23070 (N_23070,N_22357,N_20362);
xor U23071 (N_23071,N_21627,N_20707);
and U23072 (N_23072,N_22159,N_22323);
nor U23073 (N_23073,N_20885,N_20579);
or U23074 (N_23074,N_21431,N_21949);
or U23075 (N_23075,N_21769,N_22292);
or U23076 (N_23076,N_22403,N_20873);
and U23077 (N_23077,N_21525,N_22205);
or U23078 (N_23078,N_21578,N_20046);
or U23079 (N_23079,N_22241,N_21785);
nor U23080 (N_23080,N_20534,N_21811);
and U23081 (N_23081,N_21567,N_21109);
xnor U23082 (N_23082,N_21269,N_22409);
or U23083 (N_23083,N_21185,N_21125);
and U23084 (N_23084,N_20908,N_20257);
or U23085 (N_23085,N_20729,N_20214);
nor U23086 (N_23086,N_22288,N_21638);
or U23087 (N_23087,N_21345,N_20479);
xor U23088 (N_23088,N_20424,N_20381);
and U23089 (N_23089,N_20463,N_20285);
and U23090 (N_23090,N_22169,N_21335);
xnor U23091 (N_23091,N_21924,N_22453);
or U23092 (N_23092,N_21384,N_20138);
and U23093 (N_23093,N_20015,N_20913);
and U23094 (N_23094,N_20230,N_22164);
nand U23095 (N_23095,N_20706,N_21128);
and U23096 (N_23096,N_20445,N_21120);
or U23097 (N_23097,N_21714,N_21888);
and U23098 (N_23098,N_21894,N_22087);
nand U23099 (N_23099,N_22258,N_22194);
nor U23100 (N_23100,N_22166,N_20552);
nand U23101 (N_23101,N_20714,N_21461);
xnor U23102 (N_23102,N_21204,N_21740);
and U23103 (N_23103,N_22084,N_21213);
xnor U23104 (N_23104,N_20299,N_20209);
and U23105 (N_23105,N_21330,N_21822);
xnor U23106 (N_23106,N_20107,N_21698);
or U23107 (N_23107,N_20954,N_20274);
or U23108 (N_23108,N_21478,N_22000);
xnor U23109 (N_23109,N_21719,N_21144);
nor U23110 (N_23110,N_21320,N_21808);
nor U23111 (N_23111,N_20979,N_20892);
and U23112 (N_23112,N_22396,N_22077);
xnor U23113 (N_23113,N_21655,N_20403);
and U23114 (N_23114,N_21302,N_22338);
nand U23115 (N_23115,N_21999,N_21939);
nand U23116 (N_23116,N_20385,N_20484);
nand U23117 (N_23117,N_21854,N_21792);
or U23118 (N_23118,N_22007,N_21803);
and U23119 (N_23119,N_20269,N_20401);
or U23120 (N_23120,N_22114,N_21389);
nand U23121 (N_23121,N_20535,N_20429);
and U23122 (N_23122,N_20721,N_21718);
nor U23123 (N_23123,N_22495,N_22300);
or U23124 (N_23124,N_22314,N_22474);
and U23125 (N_23125,N_21794,N_20541);
xnor U23126 (N_23126,N_20188,N_20088);
nor U23127 (N_23127,N_21263,N_21251);
nor U23128 (N_23128,N_21288,N_21834);
nand U23129 (N_23129,N_22089,N_21331);
and U23130 (N_23130,N_20006,N_21253);
nand U23131 (N_23131,N_21007,N_20994);
or U23132 (N_23132,N_21529,N_21426);
nand U23133 (N_23133,N_20364,N_20680);
xnor U23134 (N_23134,N_22118,N_20582);
nor U23135 (N_23135,N_20452,N_20818);
nor U23136 (N_23136,N_20058,N_21906);
and U23137 (N_23137,N_20695,N_22229);
nor U23138 (N_23138,N_20619,N_22270);
nand U23139 (N_23139,N_21579,N_21635);
or U23140 (N_23140,N_21161,N_20351);
nand U23141 (N_23141,N_21021,N_22438);
xor U23142 (N_23142,N_20692,N_21696);
nand U23143 (N_23143,N_20661,N_22146);
or U23144 (N_23144,N_21012,N_21482);
and U23145 (N_23145,N_21368,N_21574);
or U23146 (N_23146,N_20858,N_22355);
nor U23147 (N_23147,N_21402,N_22157);
xor U23148 (N_23148,N_21542,N_20763);
xnor U23149 (N_23149,N_22131,N_20897);
and U23150 (N_23150,N_20823,N_20569);
and U23151 (N_23151,N_21602,N_21617);
and U23152 (N_23152,N_20726,N_22382);
nand U23153 (N_23153,N_20663,N_21373);
or U23154 (N_23154,N_21416,N_22293);
or U23155 (N_23155,N_21509,N_21264);
and U23156 (N_23156,N_22461,N_20179);
nand U23157 (N_23157,N_20875,N_22033);
nor U23158 (N_23158,N_21410,N_21497);
nand U23159 (N_23159,N_20273,N_21278);
nor U23160 (N_23160,N_22023,N_21991);
or U23161 (N_23161,N_21008,N_22402);
nor U23162 (N_23162,N_20549,N_21119);
or U23163 (N_23163,N_21351,N_21623);
and U23164 (N_23164,N_21048,N_20626);
or U23165 (N_23165,N_21186,N_21506);
and U23166 (N_23166,N_20640,N_20801);
and U23167 (N_23167,N_21236,N_20451);
nand U23168 (N_23168,N_21704,N_20358);
and U23169 (N_23169,N_22383,N_21855);
nor U23170 (N_23170,N_21377,N_20914);
nand U23171 (N_23171,N_20743,N_21158);
and U23172 (N_23172,N_21190,N_22329);
xor U23173 (N_23173,N_21349,N_21576);
and U23174 (N_23174,N_21528,N_21710);
or U23175 (N_23175,N_21173,N_21772);
xnor U23176 (N_23176,N_20516,N_20779);
and U23177 (N_23177,N_21285,N_22324);
nand U23178 (N_23178,N_21989,N_20405);
nor U23179 (N_23179,N_21680,N_21336);
xnor U23180 (N_23180,N_21958,N_20637);
or U23181 (N_23181,N_20513,N_21321);
nand U23182 (N_23182,N_20341,N_21722);
or U23183 (N_23183,N_21748,N_21608);
and U23184 (N_23184,N_22473,N_21950);
nor U23185 (N_23185,N_20990,N_21559);
nor U23186 (N_23186,N_21337,N_20703);
or U23187 (N_23187,N_20699,N_21116);
and U23188 (N_23188,N_21039,N_20805);
nor U23189 (N_23189,N_20505,N_21045);
or U23190 (N_23190,N_22223,N_21024);
nand U23191 (N_23191,N_20911,N_21015);
and U23192 (N_23192,N_20998,N_20055);
and U23193 (N_23193,N_20918,N_21217);
xor U23194 (N_23194,N_21814,N_20504);
nand U23195 (N_23195,N_20872,N_20118);
and U23196 (N_23196,N_21279,N_22128);
and U23197 (N_23197,N_20235,N_21948);
or U23198 (N_23198,N_22218,N_21966);
nor U23199 (N_23199,N_22302,N_21791);
nand U23200 (N_23200,N_21032,N_20684);
xnor U23201 (N_23201,N_22015,N_22025);
nor U23202 (N_23202,N_21492,N_21060);
nor U23203 (N_23203,N_22266,N_21549);
or U23204 (N_23204,N_22225,N_20882);
or U23205 (N_23205,N_21274,N_22309);
and U23206 (N_23206,N_20130,N_20249);
nand U23207 (N_23207,N_21839,N_20815);
nor U23208 (N_23208,N_20159,N_21867);
nand U23209 (N_23209,N_21157,N_21030);
or U23210 (N_23210,N_21257,N_21456);
xnor U23211 (N_23211,N_20289,N_20160);
or U23212 (N_23212,N_21026,N_20548);
xnor U23213 (N_23213,N_20890,N_21970);
nor U23214 (N_23214,N_20797,N_22424);
and U23215 (N_23215,N_21768,N_20137);
or U23216 (N_23216,N_20829,N_20361);
or U23217 (N_23217,N_20427,N_21538);
nand U23218 (N_23218,N_20537,N_20643);
nor U23219 (N_23219,N_22333,N_20377);
nand U23220 (N_23220,N_21976,N_21491);
or U23221 (N_23221,N_20997,N_21111);
or U23222 (N_23222,N_21171,N_22104);
and U23223 (N_23223,N_21467,N_22238);
nor U23224 (N_23224,N_21306,N_21581);
and U23225 (N_23225,N_21383,N_22045);
and U23226 (N_23226,N_20183,N_20820);
nand U23227 (N_23227,N_21723,N_20426);
nor U23228 (N_23228,N_21141,N_20146);
nor U23229 (N_23229,N_20995,N_21507);
or U23230 (N_23230,N_20632,N_20909);
nand U23231 (N_23231,N_21732,N_20547);
nor U23232 (N_23232,N_21046,N_20001);
nor U23233 (N_23233,N_21618,N_20478);
xnor U23234 (N_23234,N_22303,N_22410);
nand U23235 (N_23235,N_22119,N_22135);
and U23236 (N_23236,N_22139,N_21363);
or U23237 (N_23237,N_22436,N_20196);
or U23238 (N_23238,N_20087,N_20201);
and U23239 (N_23239,N_20326,N_20813);
or U23240 (N_23240,N_20980,N_22161);
nand U23241 (N_23241,N_20122,N_21708);
and U23242 (N_23242,N_20971,N_21498);
and U23243 (N_23243,N_20570,N_20157);
xnor U23244 (N_23244,N_21793,N_21477);
xnor U23245 (N_23245,N_21857,N_21073);
nand U23246 (N_23246,N_21291,N_22267);
nor U23247 (N_23247,N_20290,N_21689);
nand U23248 (N_23248,N_22452,N_22467);
nand U23249 (N_23249,N_20649,N_21000);
xor U23250 (N_23250,N_22122,N_21923);
nand U23251 (N_23251,N_20263,N_20368);
nor U23252 (N_23252,N_20800,N_20412);
and U23253 (N_23253,N_22037,N_22066);
and U23254 (N_23254,N_20009,N_21937);
and U23255 (N_23255,N_21830,N_20910);
or U23256 (N_23256,N_22214,N_20124);
xor U23257 (N_23257,N_20248,N_20631);
or U23258 (N_23258,N_21104,N_20367);
nand U23259 (N_23259,N_20032,N_20347);
nand U23260 (N_23260,N_22082,N_21891);
nand U23261 (N_23261,N_21455,N_21270);
and U23262 (N_23262,N_20480,N_21404);
and U23263 (N_23263,N_21892,N_21532);
or U23264 (N_23264,N_20037,N_22470);
and U23265 (N_23265,N_21918,N_20786);
and U23266 (N_23266,N_20826,N_20951);
and U23267 (N_23267,N_20204,N_22428);
nor U23268 (N_23268,N_21393,N_20313);
xor U23269 (N_23269,N_20139,N_21166);
nor U23270 (N_23270,N_20987,N_21129);
or U23271 (N_23271,N_21323,N_20198);
nand U23272 (N_23272,N_20932,N_20952);
nor U23273 (N_23273,N_22299,N_21831);
nand U23274 (N_23274,N_22217,N_22432);
nor U23275 (N_23275,N_21669,N_21271);
nor U23276 (N_23276,N_20243,N_22290);
nand U23277 (N_23277,N_21971,N_22282);
nor U23278 (N_23278,N_20799,N_20481);
and U23279 (N_23279,N_21052,N_20618);
nor U23280 (N_23280,N_21668,N_21927);
nand U23281 (N_23281,N_20755,N_22116);
nand U23282 (N_23282,N_21486,N_20018);
nand U23283 (N_23283,N_21610,N_21145);
nand U23284 (N_23284,N_20222,N_22418);
xor U23285 (N_23285,N_22034,N_20670);
nor U23286 (N_23286,N_20161,N_20081);
nor U23287 (N_23287,N_21607,N_22186);
and U23288 (N_23288,N_20915,N_21637);
nand U23289 (N_23289,N_21969,N_22326);
and U23290 (N_23290,N_20156,N_20040);
or U23291 (N_23291,N_21879,N_20778);
or U23292 (N_23292,N_20658,N_21787);
nand U23293 (N_23293,N_20301,N_20589);
nand U23294 (N_23294,N_20560,N_20406);
nand U23295 (N_23295,N_20765,N_20861);
or U23296 (N_23296,N_21108,N_22251);
nor U23297 (N_23297,N_20848,N_20974);
and U23298 (N_23298,N_20530,N_20667);
nand U23299 (N_23299,N_21688,N_20071);
xnor U23300 (N_23300,N_21452,N_20682);
and U23301 (N_23301,N_20712,N_22466);
and U23302 (N_23302,N_21629,N_20050);
or U23303 (N_23303,N_20365,N_20126);
and U23304 (N_23304,N_21199,N_22318);
nand U23305 (N_23305,N_20175,N_21656);
nor U23306 (N_23306,N_20874,N_21010);
or U23307 (N_23307,N_21898,N_20442);
or U23308 (N_23308,N_22029,N_21805);
nand U23309 (N_23309,N_21414,N_20331);
nor U23310 (N_23310,N_20094,N_20017);
xor U23311 (N_23311,N_21399,N_20300);
and U23312 (N_23312,N_22019,N_21872);
nand U23313 (N_23313,N_20730,N_20739);
or U23314 (N_23314,N_20717,N_21019);
and U23315 (N_23315,N_21520,N_22375);
nand U23316 (N_23316,N_20933,N_21268);
nand U23317 (N_23317,N_20796,N_20099);
nor U23318 (N_23318,N_21453,N_20229);
or U23319 (N_23319,N_22458,N_21961);
nor U23320 (N_23320,N_20953,N_21276);
or U23321 (N_23321,N_20657,N_20576);
nand U23322 (N_23322,N_20638,N_20330);
or U23323 (N_23323,N_21095,N_21980);
nand U23324 (N_23324,N_22054,N_20775);
and U23325 (N_23325,N_20639,N_21751);
nor U23326 (N_23326,N_22448,N_20976);
and U23327 (N_23327,N_20307,N_21312);
and U23328 (N_23328,N_21884,N_20583);
and U23329 (N_23329,N_21067,N_22138);
or U23330 (N_23330,N_20553,N_21694);
and U23331 (N_23331,N_21454,N_22352);
or U23332 (N_23332,N_21388,N_22469);
nor U23333 (N_23333,N_21908,N_20935);
nand U23334 (N_23334,N_21401,N_21150);
nor U23335 (N_23335,N_21308,N_22454);
nand U23336 (N_23336,N_21044,N_22407);
and U23337 (N_23337,N_21639,N_20814);
nand U23338 (N_23338,N_21967,N_22237);
nand U23339 (N_23339,N_22040,N_21512);
and U23340 (N_23340,N_20110,N_21011);
or U23341 (N_23341,N_21407,N_21836);
or U23342 (N_23342,N_22279,N_20844);
nand U23343 (N_23343,N_20194,N_22283);
and U23344 (N_23344,N_22140,N_20436);
nor U23345 (N_23345,N_20492,N_22156);
nor U23346 (N_23346,N_20891,N_22316);
nand U23347 (N_23347,N_21479,N_22244);
and U23348 (N_23348,N_21929,N_20082);
xnor U23349 (N_23349,N_20079,N_21369);
nor U23350 (N_23350,N_21952,N_22272);
nand U23351 (N_23351,N_21620,N_22390);
nor U23352 (N_23352,N_21829,N_20321);
nor U23353 (N_23353,N_20780,N_22286);
or U23354 (N_23354,N_20757,N_20766);
or U23355 (N_23355,N_20373,N_22493);
or U23356 (N_23356,N_20383,N_22416);
nand U23357 (N_23357,N_20683,N_21912);
and U23358 (N_23358,N_20900,N_21099);
and U23359 (N_23359,N_20306,N_22008);
nor U23360 (N_23360,N_21801,N_22222);
or U23361 (N_23361,N_21996,N_22068);
xor U23362 (N_23362,N_22150,N_20250);
nand U23363 (N_23363,N_21411,N_20264);
nor U23364 (N_23364,N_21299,N_21643);
or U23365 (N_23365,N_21178,N_22042);
or U23366 (N_23366,N_22090,N_20350);
nor U23367 (N_23367,N_21570,N_22327);
nand U23368 (N_23368,N_21744,N_21533);
or U23369 (N_23369,N_21424,N_20586);
nand U23370 (N_23370,N_20382,N_22192);
or U23371 (N_23371,N_21191,N_22497);
nor U23372 (N_23372,N_20108,N_21873);
and U23373 (N_23373,N_22046,N_21540);
and U23374 (N_23374,N_21667,N_21663);
and U23375 (N_23375,N_20102,N_20340);
nor U23376 (N_23376,N_22021,N_21352);
nand U23377 (N_23377,N_21167,N_22227);
nand U23378 (N_23378,N_20360,N_20180);
xnor U23379 (N_23379,N_21874,N_20465);
and U23380 (N_23380,N_21781,N_22234);
or U23381 (N_23381,N_20242,N_22422);
nand U23382 (N_23382,N_21676,N_21362);
and U23383 (N_23383,N_21951,N_20604);
and U23384 (N_23384,N_22494,N_21379);
nor U23385 (N_23385,N_21258,N_22141);
nand U23386 (N_23386,N_20275,N_22027);
and U23387 (N_23387,N_21192,N_20588);
or U23388 (N_23388,N_21018,N_22100);
nor U23389 (N_23389,N_20170,N_20446);
or U23390 (N_23390,N_21005,N_20370);
and U23391 (N_23391,N_20384,N_20978);
nand U23392 (N_23392,N_20623,N_22445);
nand U23393 (N_23393,N_20132,N_21215);
and U23394 (N_23394,N_20556,N_20096);
and U23395 (N_23395,N_22433,N_22180);
xor U23396 (N_23396,N_20936,N_21582);
or U23397 (N_23397,N_20747,N_20708);
or U23398 (N_23398,N_21437,N_21902);
nor U23399 (N_23399,N_22006,N_20319);
nor U23400 (N_23400,N_20460,N_21790);
and U23401 (N_23401,N_20339,N_21152);
and U23402 (N_23402,N_20028,N_22247);
nand U23403 (N_23403,N_20627,N_21248);
nand U23404 (N_23404,N_22268,N_21309);
nor U23405 (N_23405,N_20895,N_20066);
nor U23406 (N_23406,N_21136,N_20572);
nor U23407 (N_23407,N_21314,N_20559);
nor U23408 (N_23408,N_21983,N_20324);
nand U23409 (N_23409,N_22356,N_22320);
nor U23410 (N_23410,N_20092,N_20831);
nor U23411 (N_23411,N_20740,N_22287);
and U23412 (N_23412,N_20928,N_20490);
and U23413 (N_23413,N_21511,N_20416);
and U23414 (N_23414,N_21054,N_22328);
xor U23415 (N_23415,N_22230,N_20939);
nor U23416 (N_23416,N_21974,N_22488);
or U23417 (N_23417,N_21183,N_21913);
or U23418 (N_23418,N_20166,N_21953);
nor U23419 (N_23419,N_20924,N_20782);
and U23420 (N_23420,N_22010,N_22173);
or U23421 (N_23421,N_20609,N_22245);
nor U23422 (N_23422,N_20262,N_21179);
nand U23423 (N_23423,N_20792,N_20167);
and U23424 (N_23424,N_21817,N_20964);
xnor U23425 (N_23425,N_22289,N_21995);
xnor U23426 (N_23426,N_21715,N_20768);
nand U23427 (N_23427,N_21763,N_20881);
nand U23428 (N_23428,N_20488,N_20333);
nor U23429 (N_23429,N_20085,N_20335);
or U23430 (N_23430,N_21757,N_21177);
or U23431 (N_23431,N_22405,N_20185);
xnor U23432 (N_23432,N_21220,N_20090);
or U23433 (N_23433,N_21552,N_22380);
xnor U23434 (N_23434,N_21713,N_22057);
or U23435 (N_23435,N_22126,N_20856);
nor U23436 (N_23436,N_21707,N_20603);
and U23437 (N_23437,N_21859,N_20120);
nor U23438 (N_23438,N_21332,N_20715);
and U23439 (N_23439,N_21946,N_20105);
nor U23440 (N_23440,N_20265,N_22014);
nand U23441 (N_23441,N_20840,N_21027);
nor U23442 (N_23442,N_20084,N_21609);
or U23443 (N_23443,N_21340,N_20834);
nand U23444 (N_23444,N_20528,N_21028);
and U23445 (N_23445,N_21531,N_22155);
nand U23446 (N_23446,N_20839,N_20937);
and U23447 (N_23447,N_21889,N_21539);
nor U23448 (N_23448,N_20134,N_20510);
nor U23449 (N_23449,N_20067,N_21451);
xor U23450 (N_23450,N_21810,N_20246);
or U23451 (N_23451,N_20153,N_21137);
xnor U23452 (N_23452,N_22426,N_20602);
nand U23453 (N_23453,N_20669,N_21837);
or U23454 (N_23454,N_21092,N_21084);
nand U23455 (N_23455,N_22478,N_21063);
and U23456 (N_23456,N_21138,N_20432);
xor U23457 (N_23457,N_20654,N_21370);
or U23458 (N_23458,N_20346,N_21371);
or U23459 (N_23459,N_20329,N_20013);
and U23460 (N_23460,N_20819,N_20518);
or U23461 (N_23461,N_20688,N_21630);
and U23462 (N_23462,N_21535,N_20985);
or U23463 (N_23463,N_20961,N_21462);
or U23464 (N_23464,N_22130,N_20336);
or U23465 (N_23465,N_22344,N_20497);
nor U23466 (N_23466,N_20507,N_20397);
nand U23467 (N_23467,N_22398,N_20515);
nor U23468 (N_23468,N_20197,N_21820);
xor U23469 (N_23469,N_21848,N_20062);
and U23470 (N_23470,N_21317,N_20093);
nand U23471 (N_23471,N_20512,N_20223);
nor U23472 (N_23472,N_21743,N_22212);
xnor U23473 (N_23473,N_21361,N_21666);
or U23474 (N_23474,N_21496,N_21993);
nor U23475 (N_23475,N_21130,N_21664);
and U23476 (N_23476,N_22257,N_21035);
or U23477 (N_23477,N_20310,N_21164);
nor U23478 (N_23478,N_21524,N_20366);
and U23479 (N_23479,N_20400,N_20542);
and U23480 (N_23480,N_22187,N_21603);
or U23481 (N_23481,N_20232,N_22364);
and U23482 (N_23482,N_21514,N_21786);
or U23483 (N_23483,N_22347,N_21753);
or U23484 (N_23484,N_20379,N_21684);
nand U23485 (N_23485,N_20496,N_21468);
nor U23486 (N_23486,N_20268,N_20468);
nand U23487 (N_23487,N_20673,N_22030);
nor U23488 (N_23488,N_22254,N_21692);
or U23489 (N_23489,N_21103,N_21004);
nor U23490 (N_23490,N_22199,N_20770);
or U23491 (N_23491,N_20499,N_20546);
nor U23492 (N_23492,N_20005,N_20251);
nor U23493 (N_23493,N_20476,N_21813);
xor U23494 (N_23494,N_21175,N_22200);
nor U23495 (N_23495,N_20871,N_22451);
nor U23496 (N_23496,N_20190,N_20291);
and U23497 (N_23497,N_20317,N_22389);
nand U23498 (N_23498,N_20447,N_20388);
or U23499 (N_23499,N_22109,N_21978);
nor U23500 (N_23500,N_22028,N_21730);
and U23501 (N_23501,N_20276,N_21726);
xnor U23502 (N_23502,N_20681,N_21832);
nand U23503 (N_23503,N_22043,N_20652);
nor U23504 (N_23504,N_21886,N_20158);
xnor U23505 (N_23505,N_20742,N_20374);
nor U23506 (N_23506,N_21613,N_22198);
and U23507 (N_23507,N_20355,N_21222);
or U23508 (N_23508,N_21756,N_20622);
or U23509 (N_23509,N_21670,N_21023);
or U23510 (N_23510,N_20208,N_22202);
and U23511 (N_23511,N_21428,N_21201);
xor U23512 (N_23512,N_21193,N_21844);
nor U23513 (N_23513,N_21979,N_21973);
xor U23514 (N_23514,N_21247,N_21984);
nor U23515 (N_23515,N_21252,N_21928);
nand U23516 (N_23516,N_20010,N_21651);
nand U23517 (N_23517,N_22032,N_20150);
nor U23518 (N_23518,N_21749,N_21397);
nor U23519 (N_23519,N_21646,N_20857);
or U23520 (N_23520,N_21595,N_20532);
nand U23521 (N_23521,N_21677,N_21806);
xor U23522 (N_23522,N_21841,N_21543);
nand U23523 (N_23523,N_22259,N_20141);
nor U23524 (N_23524,N_22059,N_20135);
or U23525 (N_23525,N_21075,N_22143);
nor U23526 (N_23526,N_21254,N_20035);
or U23527 (N_23527,N_22311,N_20728);
and U23528 (N_23528,N_21833,N_21548);
and U23529 (N_23529,N_22086,N_20720);
and U23530 (N_23530,N_21475,N_21301);
or U23531 (N_23531,N_20043,N_21189);
and U23532 (N_23532,N_21483,N_20069);
xnor U23533 (N_23533,N_21106,N_20038);
nand U23534 (N_23534,N_20679,N_21560);
xor U23535 (N_23535,N_21464,N_21143);
nor U23536 (N_23536,N_20655,N_20989);
or U23537 (N_23537,N_20592,N_21188);
nand U23538 (N_23538,N_21013,N_21221);
nand U23539 (N_23539,N_21284,N_21764);
xnor U23540 (N_23540,N_20255,N_22379);
or U23541 (N_23541,N_20821,N_21072);
or U23542 (N_23542,N_21515,N_20164);
nor U23543 (N_23543,N_20804,N_20049);
or U23544 (N_23544,N_22394,N_22020);
and U23545 (N_23545,N_21558,N_20674);
nor U23546 (N_23546,N_20075,N_22341);
nor U23547 (N_23547,N_21062,N_20095);
and U23548 (N_23548,N_20097,N_22207);
nor U23549 (N_23549,N_21631,N_20391);
nor U23550 (N_23550,N_21910,N_22096);
and U23551 (N_23551,N_21650,N_21850);
nor U23552 (N_23552,N_22132,N_21911);
and U23553 (N_23553,N_20645,N_22153);
or U23554 (N_23554,N_20219,N_21505);
or U23555 (N_23555,N_22243,N_21366);
nand U23556 (N_23556,N_20475,N_22088);
nand U23557 (N_23557,N_22430,N_21450);
nor U23558 (N_23558,N_22168,N_21701);
and U23559 (N_23559,N_21517,N_20594);
xnor U23560 (N_23560,N_21932,N_21500);
nand U23561 (N_23561,N_22121,N_20777);
and U23562 (N_23562,N_21716,N_21728);
and U23563 (N_23563,N_21742,N_20571);
and U23564 (N_23564,N_22351,N_20133);
or U23565 (N_23565,N_22491,N_21043);
nand U23566 (N_23566,N_22184,N_21940);
or U23567 (N_23567,N_20297,N_22026);
nor U23568 (N_23568,N_21187,N_21883);
nand U23569 (N_23569,N_21071,N_21212);
nand U23570 (N_23570,N_20039,N_22343);
or U23571 (N_23571,N_21495,N_22178);
nand U23572 (N_23572,N_22071,N_20178);
or U23573 (N_23573,N_20304,N_20853);
and U23574 (N_23574,N_22271,N_21672);
or U23575 (N_23575,N_20462,N_20109);
nor U23576 (N_23576,N_20486,N_21074);
and U23577 (N_23577,N_20693,N_22440);
and U23578 (N_23578,N_21819,N_20888);
nand U23579 (N_23579,N_22353,N_21765);
or U23580 (N_23580,N_21925,N_22224);
or U23581 (N_23581,N_21344,N_21493);
and U23582 (N_23582,N_21711,N_22240);
nand U23583 (N_23583,N_22413,N_20294);
and U23584 (N_23584,N_21057,N_20205);
nor U23585 (N_23585,N_20789,N_21501);
and U23586 (N_23586,N_21802,N_20440);
or U23587 (N_23587,N_20024,N_20942);
nor U23588 (N_23588,N_22196,N_20793);
or U23589 (N_23589,N_21197,N_21986);
or U23590 (N_23590,N_21720,N_21316);
nor U23591 (N_23591,N_20325,N_20298);
and U23592 (N_23592,N_21259,N_21981);
and U23593 (N_23593,N_21036,N_21838);
and U23594 (N_23594,N_21736,N_21480);
and U23595 (N_23595,N_22366,N_21358);
and U23596 (N_23596,N_21250,N_22301);
and U23597 (N_23597,N_21472,N_20698);
or U23598 (N_23598,N_21430,N_22277);
or U23599 (N_23599,N_20474,N_21123);
nor U23600 (N_23600,N_21599,N_20211);
nand U23601 (N_23601,N_21571,N_21816);
nor U23602 (N_23602,N_20144,N_21360);
or U23603 (N_23603,N_20457,N_20419);
nand U23604 (N_23604,N_20912,N_21544);
nor U23605 (N_23605,N_21545,N_20741);
or U23606 (N_23606,N_21476,N_21154);
and U23607 (N_23607,N_21513,N_20163);
and U23608 (N_23608,N_20666,N_20439);
xor U23609 (N_23609,N_20303,N_21604);
and U23610 (N_23610,N_20893,N_20529);
or U23611 (N_23611,N_22210,N_22388);
and U23612 (N_23612,N_21294,N_21445);
or U23613 (N_23613,N_20025,N_21326);
or U23614 (N_23614,N_20852,N_20393);
and U23615 (N_23615,N_22149,N_22330);
xor U23616 (N_23616,N_20186,N_21295);
and U23617 (N_23617,N_20176,N_21856);
and U23618 (N_23618,N_22226,N_21146);
nand U23619 (N_23619,N_20705,N_22101);
and U23620 (N_23620,N_21489,N_21997);
or U23621 (N_23621,N_21237,N_21649);
and U23622 (N_23622,N_22002,N_21665);
nor U23623 (N_23623,N_22358,N_22331);
nand U23624 (N_23624,N_20332,N_20906);
xor U23625 (N_23625,N_20563,N_21931);
nor U23626 (N_23626,N_21020,N_20523);
and U23627 (N_23627,N_21942,N_21037);
nand U23628 (N_23628,N_21926,N_22107);
nor U23629 (N_23629,N_20315,N_20764);
and U23630 (N_23630,N_20959,N_22073);
and U23631 (N_23631,N_20545,N_21687);
nor U23632 (N_23632,N_22133,N_20200);
and U23633 (N_23633,N_20192,N_22312);
nand U23634 (N_23634,N_20904,N_21690);
and U23635 (N_23635,N_22081,N_22160);
and U23636 (N_23636,N_21229,N_21202);
or U23637 (N_23637,N_20651,N_21930);
and U23638 (N_23638,N_20686,N_21598);
and U23639 (N_23639,N_22305,N_21444);
nor U23640 (N_23640,N_21378,N_20880);
or U23641 (N_23641,N_22050,N_22052);
xor U23642 (N_23642,N_21565,N_21364);
or U23643 (N_23643,N_22113,N_21280);
and U23644 (N_23644,N_21114,N_20854);
nor U23645 (N_23645,N_20702,N_20605);
or U23646 (N_23646,N_21724,N_21868);
and U23647 (N_23647,N_21313,N_20060);
or U23648 (N_23648,N_21935,N_21423);
nand U23649 (N_23649,N_20008,N_20543);
or U23650 (N_23650,N_20656,N_20629);
and U23651 (N_23651,N_20807,N_20636);
nor U23652 (N_23652,N_21182,N_20221);
nor U23653 (N_23653,N_21198,N_20337);
and U23654 (N_23654,N_21156,N_22278);
and U23655 (N_23655,N_20817,N_20991);
nand U23656 (N_23656,N_20076,N_20521);
nor U23657 (N_23657,N_20193,N_22468);
or U23658 (N_23658,N_20585,N_20749);
nand U23659 (N_23659,N_21342,N_21797);
and U23660 (N_23660,N_20533,N_21133);
nand U23661 (N_23661,N_20660,N_21933);
or U23662 (N_23662,N_21729,N_20863);
xor U23663 (N_23663,N_20653,N_21218);
and U23664 (N_23664,N_21959,N_20349);
nor U23665 (N_23665,N_22056,N_20967);
or U23666 (N_23666,N_22170,N_21470);
and U23667 (N_23667,N_20395,N_22446);
and U23668 (N_23668,N_21594,N_21267);
or U23669 (N_23669,N_21086,N_20866);
or U23670 (N_23670,N_20948,N_20140);
xor U23671 (N_23671,N_20106,N_21289);
nand U23672 (N_23672,N_20926,N_20283);
or U23673 (N_23673,N_21671,N_22102);
nand U23674 (N_23674,N_20648,N_21821);
and U23675 (N_23675,N_22360,N_22189);
and U23676 (N_23676,N_20458,N_20064);
nand U23677 (N_23677,N_21132,N_21563);
or U23678 (N_23678,N_21042,N_20371);
nor U23679 (N_23679,N_22395,N_21659);
nor U23680 (N_23680,N_21987,N_22083);
nor U23681 (N_23681,N_21324,N_22483);
or U23682 (N_23682,N_22342,N_21881);
nor U23683 (N_23683,N_22496,N_22018);
nand U23684 (N_23684,N_22372,N_21050);
and U23685 (N_23685,N_20597,N_20435);
nand U23686 (N_23686,N_21702,N_21566);
or U23687 (N_23687,N_20981,N_21634);
xnor U23688 (N_23688,N_21955,N_21135);
nand U23689 (N_23689,N_22142,N_20869);
nor U23690 (N_23690,N_20694,N_22001);
and U23691 (N_23691,N_21977,N_20735);
and U23692 (N_23692,N_21297,N_21246);
nand U23693 (N_23693,N_21168,N_21626);
nor U23694 (N_23694,N_22365,N_22092);
nand U23695 (N_23695,N_20177,N_20520);
xnor U23696 (N_23696,N_21914,N_22144);
or U23697 (N_23697,N_21735,N_20849);
xor U23698 (N_23698,N_21275,N_22275);
nand U23699 (N_23699,N_20808,N_21122);
and U23700 (N_23700,N_20600,N_22176);
or U23701 (N_23701,N_21398,N_22423);
and U23702 (N_23702,N_21731,N_21429);
or U23703 (N_23703,N_20165,N_21904);
and U23704 (N_23704,N_20080,N_20811);
nand U23705 (N_23705,N_21014,N_21990);
nand U23706 (N_23706,N_21118,N_22295);
nor U23707 (N_23707,N_22206,N_22484);
nand U23708 (N_23708,N_22072,N_20267);
nor U23709 (N_23709,N_21415,N_22419);
nor U23710 (N_23710,N_21683,N_20555);
nor U23711 (N_23711,N_20047,N_20625);
and U23712 (N_23712,N_21070,N_20389);
and U23713 (N_23713,N_21636,N_21877);
xor U23714 (N_23714,N_21606,N_22455);
xor U23715 (N_23715,N_21355,N_21240);
nor U23716 (N_23716,N_21322,N_21861);
or U23717 (N_23717,N_21359,N_22362);
nand U23718 (N_23718,N_20425,N_21569);
and U23719 (N_23719,N_20791,N_20996);
nand U23720 (N_23720,N_22441,N_20606);
and U23721 (N_23721,N_21226,N_20960);
nor U23722 (N_23722,N_20293,N_22111);
and U23723 (N_23723,N_20059,N_22055);
xnor U23724 (N_23724,N_22061,N_21436);
or U23725 (N_23725,N_20785,N_21605);
and U23726 (N_23726,N_22123,N_20195);
xnor U23727 (N_23727,N_20327,N_22399);
or U23728 (N_23728,N_21555,N_22421);
nor U23729 (N_23729,N_21583,N_20220);
or U23730 (N_23730,N_20453,N_20308);
and U23731 (N_23731,N_21536,N_21165);
nand U23732 (N_23732,N_20554,N_20378);
nand U23733 (N_23733,N_20399,N_20538);
nand U23734 (N_23734,N_20860,N_22145);
nor U23735 (N_23735,N_20007,N_20762);
nor U23736 (N_23736,N_21265,N_21534);
and U23737 (N_23737,N_22459,N_20573);
nor U23738 (N_23738,N_20237,N_20498);
nand U23739 (N_23739,N_21624,N_20004);
or U23740 (N_23740,N_20380,N_20744);
or U23741 (N_23741,N_20539,N_20993);
nand U23742 (N_23742,N_20410,N_21812);
or U23743 (N_23743,N_20878,N_22174);
xor U23744 (N_23744,N_20411,N_20086);
nand U23745 (N_23745,N_21089,N_22262);
nand U23746 (N_23746,N_20356,N_21107);
and U23747 (N_23747,N_21333,N_21310);
nand U23748 (N_23748,N_21746,N_20466);
nand U23749 (N_23749,N_20567,N_21262);
or U23750 (N_23750,N_22354,N_20750);
and U23751 (N_23751,N_20593,N_21475);
nor U23752 (N_23752,N_21029,N_21314);
nor U23753 (N_23753,N_20085,N_21123);
xor U23754 (N_23754,N_20614,N_21568);
and U23755 (N_23755,N_22326,N_22192);
nor U23756 (N_23756,N_21034,N_21164);
or U23757 (N_23757,N_20840,N_20771);
or U23758 (N_23758,N_20289,N_21291);
nand U23759 (N_23759,N_21353,N_22192);
nor U23760 (N_23760,N_22317,N_21071);
xnor U23761 (N_23761,N_22247,N_20754);
and U23762 (N_23762,N_22166,N_20678);
or U23763 (N_23763,N_20768,N_21433);
xor U23764 (N_23764,N_22288,N_20691);
or U23765 (N_23765,N_20475,N_21451);
or U23766 (N_23766,N_20591,N_20996);
nor U23767 (N_23767,N_22091,N_21024);
nor U23768 (N_23768,N_20581,N_22013);
nand U23769 (N_23769,N_20856,N_21380);
or U23770 (N_23770,N_20748,N_21912);
nand U23771 (N_23771,N_22159,N_21961);
nand U23772 (N_23772,N_21565,N_21277);
or U23773 (N_23773,N_21434,N_21630);
and U23774 (N_23774,N_20405,N_22142);
nor U23775 (N_23775,N_20962,N_21592);
or U23776 (N_23776,N_22371,N_21929);
nor U23777 (N_23777,N_22359,N_21735);
nor U23778 (N_23778,N_21527,N_21909);
or U23779 (N_23779,N_21930,N_20936);
nor U23780 (N_23780,N_20129,N_20394);
and U23781 (N_23781,N_22283,N_21220);
nand U23782 (N_23782,N_21261,N_20763);
nor U23783 (N_23783,N_20281,N_20473);
and U23784 (N_23784,N_20835,N_22184);
and U23785 (N_23785,N_21461,N_21207);
or U23786 (N_23786,N_21073,N_21693);
or U23787 (N_23787,N_20158,N_20665);
and U23788 (N_23788,N_21358,N_20038);
or U23789 (N_23789,N_20385,N_22432);
or U23790 (N_23790,N_21638,N_21031);
and U23791 (N_23791,N_20992,N_20980);
xnor U23792 (N_23792,N_21905,N_21350);
nand U23793 (N_23793,N_21262,N_22391);
xnor U23794 (N_23794,N_20140,N_21603);
or U23795 (N_23795,N_20065,N_21826);
nand U23796 (N_23796,N_20656,N_20673);
and U23797 (N_23797,N_20092,N_20162);
and U23798 (N_23798,N_22206,N_22320);
xnor U23799 (N_23799,N_22381,N_22073);
and U23800 (N_23800,N_21096,N_21022);
xor U23801 (N_23801,N_21375,N_21357);
and U23802 (N_23802,N_20416,N_20303);
or U23803 (N_23803,N_21163,N_20192);
nand U23804 (N_23804,N_21137,N_20557);
nand U23805 (N_23805,N_21302,N_20265);
nor U23806 (N_23806,N_20294,N_22052);
and U23807 (N_23807,N_20295,N_20963);
and U23808 (N_23808,N_22348,N_21228);
nand U23809 (N_23809,N_20773,N_21483);
and U23810 (N_23810,N_20335,N_21387);
xor U23811 (N_23811,N_20223,N_20063);
and U23812 (N_23812,N_20731,N_21411);
and U23813 (N_23813,N_21106,N_21962);
nand U23814 (N_23814,N_21910,N_21334);
and U23815 (N_23815,N_21204,N_21752);
or U23816 (N_23816,N_21900,N_21976);
and U23817 (N_23817,N_21514,N_21731);
nor U23818 (N_23818,N_22422,N_21876);
nor U23819 (N_23819,N_20102,N_21048);
nor U23820 (N_23820,N_21691,N_20708);
and U23821 (N_23821,N_20801,N_20964);
and U23822 (N_23822,N_22186,N_20689);
nand U23823 (N_23823,N_21007,N_20540);
and U23824 (N_23824,N_21800,N_21011);
nor U23825 (N_23825,N_22366,N_21005);
nand U23826 (N_23826,N_20336,N_21789);
or U23827 (N_23827,N_21041,N_21949);
or U23828 (N_23828,N_22440,N_20697);
or U23829 (N_23829,N_22396,N_22408);
and U23830 (N_23830,N_20163,N_22235);
nand U23831 (N_23831,N_21980,N_21413);
or U23832 (N_23832,N_20526,N_21818);
xnor U23833 (N_23833,N_20393,N_20275);
nand U23834 (N_23834,N_21375,N_21864);
nor U23835 (N_23835,N_22258,N_20788);
nor U23836 (N_23836,N_21240,N_20179);
xor U23837 (N_23837,N_21597,N_21393);
nand U23838 (N_23838,N_21905,N_21852);
and U23839 (N_23839,N_20313,N_22097);
xor U23840 (N_23840,N_20513,N_21430);
nor U23841 (N_23841,N_21214,N_21313);
and U23842 (N_23842,N_22401,N_21090);
nand U23843 (N_23843,N_22342,N_21258);
nand U23844 (N_23844,N_21293,N_21270);
or U23845 (N_23845,N_20106,N_21259);
xor U23846 (N_23846,N_21388,N_20382);
and U23847 (N_23847,N_20271,N_21080);
nand U23848 (N_23848,N_20503,N_21247);
xor U23849 (N_23849,N_21683,N_21346);
or U23850 (N_23850,N_22280,N_22344);
and U23851 (N_23851,N_20129,N_22148);
nand U23852 (N_23852,N_20187,N_20803);
nor U23853 (N_23853,N_22204,N_21828);
and U23854 (N_23854,N_20397,N_20901);
xor U23855 (N_23855,N_21241,N_22159);
or U23856 (N_23856,N_21570,N_22193);
nand U23857 (N_23857,N_20778,N_20973);
nand U23858 (N_23858,N_20205,N_20321);
nor U23859 (N_23859,N_21689,N_20474);
and U23860 (N_23860,N_22170,N_20594);
nand U23861 (N_23861,N_21319,N_20621);
xor U23862 (N_23862,N_21516,N_20181);
or U23863 (N_23863,N_20486,N_21508);
nor U23864 (N_23864,N_21911,N_20778);
nor U23865 (N_23865,N_22189,N_20165);
or U23866 (N_23866,N_22119,N_20946);
nor U23867 (N_23867,N_20092,N_21304);
and U23868 (N_23868,N_22180,N_22229);
nor U23869 (N_23869,N_21531,N_20173);
nor U23870 (N_23870,N_21922,N_22332);
nand U23871 (N_23871,N_20335,N_20537);
nor U23872 (N_23872,N_21179,N_21222);
and U23873 (N_23873,N_21831,N_20572);
nor U23874 (N_23874,N_21919,N_21050);
xor U23875 (N_23875,N_20614,N_21352);
or U23876 (N_23876,N_22346,N_20869);
xnor U23877 (N_23877,N_20977,N_20866);
and U23878 (N_23878,N_20023,N_20157);
nor U23879 (N_23879,N_20519,N_21811);
and U23880 (N_23880,N_20856,N_20375);
and U23881 (N_23881,N_21909,N_21493);
nand U23882 (N_23882,N_20702,N_22345);
nand U23883 (N_23883,N_22437,N_21277);
or U23884 (N_23884,N_20256,N_20840);
nand U23885 (N_23885,N_21798,N_21344);
xnor U23886 (N_23886,N_20053,N_20829);
nand U23887 (N_23887,N_20467,N_20494);
nand U23888 (N_23888,N_20773,N_21468);
nor U23889 (N_23889,N_21379,N_21178);
or U23890 (N_23890,N_20199,N_20662);
nand U23891 (N_23891,N_21749,N_20161);
and U23892 (N_23892,N_21052,N_21756);
xor U23893 (N_23893,N_21754,N_22425);
or U23894 (N_23894,N_21755,N_21288);
nand U23895 (N_23895,N_22461,N_20517);
nand U23896 (N_23896,N_21341,N_21876);
nand U23897 (N_23897,N_22086,N_21370);
or U23898 (N_23898,N_20964,N_20390);
and U23899 (N_23899,N_22480,N_21670);
or U23900 (N_23900,N_22035,N_21628);
or U23901 (N_23901,N_20201,N_22131);
or U23902 (N_23902,N_21204,N_22281);
or U23903 (N_23903,N_22350,N_22252);
xor U23904 (N_23904,N_21978,N_21649);
and U23905 (N_23905,N_20125,N_22387);
nand U23906 (N_23906,N_21080,N_20697);
nand U23907 (N_23907,N_21350,N_22425);
xnor U23908 (N_23908,N_20209,N_20754);
nor U23909 (N_23909,N_22080,N_22297);
or U23910 (N_23910,N_21585,N_22291);
xnor U23911 (N_23911,N_21135,N_20388);
nand U23912 (N_23912,N_20856,N_20872);
or U23913 (N_23913,N_20849,N_21739);
xnor U23914 (N_23914,N_20489,N_22269);
nor U23915 (N_23915,N_22180,N_20525);
nand U23916 (N_23916,N_21192,N_20003);
or U23917 (N_23917,N_20702,N_21196);
or U23918 (N_23918,N_20042,N_20176);
xnor U23919 (N_23919,N_21566,N_21802);
and U23920 (N_23920,N_21219,N_21066);
and U23921 (N_23921,N_22409,N_20643);
or U23922 (N_23922,N_20513,N_21592);
nor U23923 (N_23923,N_20526,N_20102);
and U23924 (N_23924,N_20954,N_21841);
nor U23925 (N_23925,N_21604,N_21821);
nor U23926 (N_23926,N_21876,N_20563);
nor U23927 (N_23927,N_20576,N_21726);
nor U23928 (N_23928,N_20305,N_20707);
nand U23929 (N_23929,N_21695,N_21823);
nand U23930 (N_23930,N_21719,N_21427);
or U23931 (N_23931,N_21781,N_20143);
nor U23932 (N_23932,N_22400,N_22055);
nor U23933 (N_23933,N_22143,N_20672);
nor U23934 (N_23934,N_20287,N_22097);
nor U23935 (N_23935,N_21503,N_20455);
nand U23936 (N_23936,N_21046,N_21341);
nor U23937 (N_23937,N_22051,N_21949);
and U23938 (N_23938,N_21425,N_21136);
nor U23939 (N_23939,N_21001,N_20691);
and U23940 (N_23940,N_20417,N_21869);
or U23941 (N_23941,N_22395,N_22182);
and U23942 (N_23942,N_22275,N_20127);
nand U23943 (N_23943,N_22304,N_21201);
xor U23944 (N_23944,N_22385,N_22410);
nor U23945 (N_23945,N_20160,N_20103);
nor U23946 (N_23946,N_20163,N_20372);
nor U23947 (N_23947,N_21394,N_21119);
nand U23948 (N_23948,N_21296,N_21593);
or U23949 (N_23949,N_21383,N_22457);
and U23950 (N_23950,N_20352,N_20829);
nand U23951 (N_23951,N_22221,N_20572);
nand U23952 (N_23952,N_20180,N_20772);
or U23953 (N_23953,N_21698,N_20425);
and U23954 (N_23954,N_21520,N_21350);
or U23955 (N_23955,N_22306,N_22272);
nor U23956 (N_23956,N_21569,N_21518);
xnor U23957 (N_23957,N_21044,N_21358);
nand U23958 (N_23958,N_21047,N_21117);
nor U23959 (N_23959,N_21273,N_20411);
nand U23960 (N_23960,N_20234,N_22471);
nand U23961 (N_23961,N_21299,N_21933);
xnor U23962 (N_23962,N_21987,N_21400);
nand U23963 (N_23963,N_21963,N_21678);
and U23964 (N_23964,N_20408,N_21214);
nor U23965 (N_23965,N_20346,N_22158);
xor U23966 (N_23966,N_21262,N_21080);
nor U23967 (N_23967,N_21965,N_21910);
and U23968 (N_23968,N_21334,N_20968);
or U23969 (N_23969,N_20622,N_21199);
nor U23970 (N_23970,N_21729,N_20965);
nor U23971 (N_23971,N_22063,N_20571);
or U23972 (N_23972,N_22404,N_21103);
xor U23973 (N_23973,N_21250,N_22005);
nor U23974 (N_23974,N_20173,N_21546);
and U23975 (N_23975,N_20813,N_22062);
and U23976 (N_23976,N_21636,N_20951);
nor U23977 (N_23977,N_21292,N_21935);
nand U23978 (N_23978,N_22412,N_21466);
xor U23979 (N_23979,N_22409,N_22087);
nor U23980 (N_23980,N_20708,N_22214);
and U23981 (N_23981,N_22449,N_21078);
nor U23982 (N_23982,N_22497,N_22003);
and U23983 (N_23983,N_22269,N_21471);
or U23984 (N_23984,N_22321,N_20460);
and U23985 (N_23985,N_21407,N_21780);
or U23986 (N_23986,N_22203,N_21497);
nand U23987 (N_23987,N_21390,N_22257);
or U23988 (N_23988,N_21455,N_20734);
and U23989 (N_23989,N_22207,N_22150);
nor U23990 (N_23990,N_22185,N_21539);
xor U23991 (N_23991,N_21940,N_20055);
nor U23992 (N_23992,N_20335,N_20660);
xor U23993 (N_23993,N_20274,N_20042);
or U23994 (N_23994,N_21263,N_22120);
nand U23995 (N_23995,N_20420,N_21143);
xor U23996 (N_23996,N_21046,N_20765);
nand U23997 (N_23997,N_22299,N_21076);
or U23998 (N_23998,N_20762,N_21080);
nor U23999 (N_23999,N_22477,N_21456);
nor U24000 (N_24000,N_20815,N_20415);
nand U24001 (N_24001,N_20796,N_20684);
nor U24002 (N_24002,N_22376,N_22025);
and U24003 (N_24003,N_22362,N_22263);
nor U24004 (N_24004,N_21206,N_20728);
nand U24005 (N_24005,N_21970,N_20323);
or U24006 (N_24006,N_20042,N_21294);
nor U24007 (N_24007,N_20710,N_20568);
nor U24008 (N_24008,N_20410,N_21636);
and U24009 (N_24009,N_21763,N_20053);
and U24010 (N_24010,N_21812,N_21035);
nand U24011 (N_24011,N_21815,N_21480);
nor U24012 (N_24012,N_20428,N_21354);
and U24013 (N_24013,N_21804,N_21558);
nor U24014 (N_24014,N_21178,N_21961);
nand U24015 (N_24015,N_21311,N_20032);
nand U24016 (N_24016,N_22490,N_20632);
xnor U24017 (N_24017,N_20027,N_20817);
nand U24018 (N_24018,N_21460,N_22259);
and U24019 (N_24019,N_20300,N_21505);
xnor U24020 (N_24020,N_21959,N_20004);
and U24021 (N_24021,N_20971,N_20583);
nand U24022 (N_24022,N_21101,N_21294);
nor U24023 (N_24023,N_20340,N_22366);
nand U24024 (N_24024,N_21677,N_22458);
xnor U24025 (N_24025,N_20267,N_22123);
and U24026 (N_24026,N_21082,N_20200);
or U24027 (N_24027,N_22278,N_21541);
nor U24028 (N_24028,N_21730,N_20856);
nor U24029 (N_24029,N_20507,N_21747);
nand U24030 (N_24030,N_21427,N_20605);
nor U24031 (N_24031,N_20560,N_20317);
nor U24032 (N_24032,N_22124,N_20514);
nand U24033 (N_24033,N_22414,N_20506);
and U24034 (N_24034,N_21366,N_21959);
nand U24035 (N_24035,N_20451,N_21955);
and U24036 (N_24036,N_20594,N_21626);
or U24037 (N_24037,N_22119,N_20042);
nor U24038 (N_24038,N_21289,N_20516);
and U24039 (N_24039,N_21495,N_20154);
nand U24040 (N_24040,N_20033,N_21288);
nand U24041 (N_24041,N_21842,N_20303);
or U24042 (N_24042,N_21724,N_22160);
nand U24043 (N_24043,N_22455,N_20437);
and U24044 (N_24044,N_21969,N_22076);
nor U24045 (N_24045,N_21940,N_21432);
nor U24046 (N_24046,N_21285,N_20010);
and U24047 (N_24047,N_20263,N_22374);
or U24048 (N_24048,N_21661,N_21830);
and U24049 (N_24049,N_22352,N_21749);
or U24050 (N_24050,N_20271,N_20013);
nor U24051 (N_24051,N_20227,N_20600);
and U24052 (N_24052,N_21004,N_21056);
nor U24053 (N_24053,N_20018,N_21284);
and U24054 (N_24054,N_20166,N_20596);
nand U24055 (N_24055,N_22207,N_21161);
nor U24056 (N_24056,N_22137,N_22219);
nor U24057 (N_24057,N_20966,N_20140);
nand U24058 (N_24058,N_20854,N_20772);
or U24059 (N_24059,N_20661,N_22481);
nor U24060 (N_24060,N_21733,N_20177);
or U24061 (N_24061,N_21070,N_21153);
and U24062 (N_24062,N_20505,N_21327);
nand U24063 (N_24063,N_20812,N_21670);
nor U24064 (N_24064,N_22038,N_21773);
nand U24065 (N_24065,N_22295,N_20199);
or U24066 (N_24066,N_21965,N_20695);
and U24067 (N_24067,N_21951,N_20000);
xnor U24068 (N_24068,N_21810,N_20690);
nand U24069 (N_24069,N_20453,N_20708);
nand U24070 (N_24070,N_22091,N_21199);
and U24071 (N_24071,N_21175,N_21227);
nor U24072 (N_24072,N_21331,N_20430);
xor U24073 (N_24073,N_22339,N_22399);
nand U24074 (N_24074,N_21818,N_21887);
xnor U24075 (N_24075,N_20040,N_21192);
and U24076 (N_24076,N_21871,N_20647);
and U24077 (N_24077,N_22457,N_20284);
nand U24078 (N_24078,N_20521,N_21549);
xor U24079 (N_24079,N_20005,N_20971);
and U24080 (N_24080,N_20006,N_20600);
xnor U24081 (N_24081,N_22410,N_22061);
nand U24082 (N_24082,N_20937,N_22468);
or U24083 (N_24083,N_21661,N_20545);
nand U24084 (N_24084,N_21898,N_21837);
nor U24085 (N_24085,N_20655,N_22303);
nor U24086 (N_24086,N_21001,N_20206);
and U24087 (N_24087,N_22277,N_22497);
or U24088 (N_24088,N_21698,N_20702);
and U24089 (N_24089,N_20086,N_20752);
or U24090 (N_24090,N_20501,N_21610);
or U24091 (N_24091,N_20181,N_22012);
nand U24092 (N_24092,N_20567,N_21639);
and U24093 (N_24093,N_20540,N_21584);
or U24094 (N_24094,N_20986,N_20425);
nand U24095 (N_24095,N_20578,N_22170);
nor U24096 (N_24096,N_21297,N_20109);
and U24097 (N_24097,N_21739,N_21477);
and U24098 (N_24098,N_21314,N_20348);
and U24099 (N_24099,N_21166,N_20070);
or U24100 (N_24100,N_20241,N_20033);
or U24101 (N_24101,N_21421,N_20299);
nor U24102 (N_24102,N_20166,N_22069);
nor U24103 (N_24103,N_20781,N_20644);
nand U24104 (N_24104,N_21901,N_20842);
nor U24105 (N_24105,N_20871,N_20821);
and U24106 (N_24106,N_21830,N_20983);
nand U24107 (N_24107,N_22015,N_21754);
nand U24108 (N_24108,N_22089,N_21476);
nor U24109 (N_24109,N_21533,N_21291);
or U24110 (N_24110,N_20994,N_21029);
or U24111 (N_24111,N_21425,N_21471);
or U24112 (N_24112,N_21109,N_21915);
nand U24113 (N_24113,N_21828,N_21877);
and U24114 (N_24114,N_22122,N_21364);
nor U24115 (N_24115,N_20625,N_21745);
nor U24116 (N_24116,N_21749,N_20098);
nand U24117 (N_24117,N_20653,N_21871);
or U24118 (N_24118,N_20703,N_20670);
nand U24119 (N_24119,N_20594,N_21103);
or U24120 (N_24120,N_21946,N_21649);
nor U24121 (N_24121,N_20708,N_20186);
and U24122 (N_24122,N_21681,N_20525);
and U24123 (N_24123,N_20227,N_21501);
or U24124 (N_24124,N_20684,N_20007);
nor U24125 (N_24125,N_20304,N_22466);
and U24126 (N_24126,N_21773,N_21567);
and U24127 (N_24127,N_20119,N_20220);
nand U24128 (N_24128,N_20970,N_20777);
and U24129 (N_24129,N_20905,N_21572);
or U24130 (N_24130,N_20621,N_20887);
nor U24131 (N_24131,N_22481,N_22418);
and U24132 (N_24132,N_20089,N_21309);
or U24133 (N_24133,N_20543,N_20252);
nand U24134 (N_24134,N_22080,N_20973);
or U24135 (N_24135,N_20909,N_20366);
or U24136 (N_24136,N_21710,N_20857);
or U24137 (N_24137,N_20519,N_21230);
or U24138 (N_24138,N_21885,N_21162);
xor U24139 (N_24139,N_20712,N_21054);
or U24140 (N_24140,N_20140,N_21901);
and U24141 (N_24141,N_20666,N_21724);
or U24142 (N_24142,N_21530,N_20798);
xnor U24143 (N_24143,N_20125,N_21481);
nor U24144 (N_24144,N_22327,N_21771);
nor U24145 (N_24145,N_20024,N_20351);
xor U24146 (N_24146,N_20330,N_21173);
nor U24147 (N_24147,N_21700,N_20033);
nand U24148 (N_24148,N_22207,N_20841);
and U24149 (N_24149,N_22197,N_20364);
nand U24150 (N_24150,N_22424,N_21623);
or U24151 (N_24151,N_21214,N_21234);
and U24152 (N_24152,N_20556,N_20272);
and U24153 (N_24153,N_21547,N_20010);
nand U24154 (N_24154,N_20134,N_20294);
or U24155 (N_24155,N_21635,N_20411);
or U24156 (N_24156,N_20165,N_22006);
and U24157 (N_24157,N_21359,N_21460);
nand U24158 (N_24158,N_20079,N_22108);
nand U24159 (N_24159,N_20281,N_21109);
nor U24160 (N_24160,N_21314,N_20601);
or U24161 (N_24161,N_20426,N_21364);
and U24162 (N_24162,N_21319,N_22094);
nor U24163 (N_24163,N_21281,N_22096);
nand U24164 (N_24164,N_22028,N_20134);
or U24165 (N_24165,N_22434,N_21005);
or U24166 (N_24166,N_20201,N_21464);
or U24167 (N_24167,N_21370,N_20353);
or U24168 (N_24168,N_22498,N_21734);
or U24169 (N_24169,N_21735,N_22256);
and U24170 (N_24170,N_20142,N_21216);
nor U24171 (N_24171,N_21544,N_20190);
nor U24172 (N_24172,N_20375,N_22488);
and U24173 (N_24173,N_21545,N_21916);
or U24174 (N_24174,N_20196,N_21959);
or U24175 (N_24175,N_21313,N_21324);
and U24176 (N_24176,N_20406,N_20596);
xor U24177 (N_24177,N_21491,N_21379);
and U24178 (N_24178,N_21189,N_21904);
nor U24179 (N_24179,N_20324,N_20557);
nor U24180 (N_24180,N_21423,N_20765);
nand U24181 (N_24181,N_21610,N_21105);
and U24182 (N_24182,N_21743,N_22400);
nand U24183 (N_24183,N_22161,N_20496);
and U24184 (N_24184,N_22394,N_21773);
or U24185 (N_24185,N_21280,N_22351);
or U24186 (N_24186,N_20313,N_20998);
or U24187 (N_24187,N_21546,N_21046);
and U24188 (N_24188,N_20276,N_20673);
and U24189 (N_24189,N_21320,N_21979);
or U24190 (N_24190,N_20637,N_20518);
and U24191 (N_24191,N_20790,N_20438);
and U24192 (N_24192,N_22300,N_21061);
nand U24193 (N_24193,N_20101,N_21546);
nand U24194 (N_24194,N_21827,N_21497);
and U24195 (N_24195,N_20779,N_21351);
nor U24196 (N_24196,N_20698,N_22305);
xnor U24197 (N_24197,N_20321,N_20038);
nor U24198 (N_24198,N_21499,N_20141);
nand U24199 (N_24199,N_21744,N_21428);
and U24200 (N_24200,N_21680,N_20455);
or U24201 (N_24201,N_22444,N_22495);
nand U24202 (N_24202,N_22208,N_21734);
nand U24203 (N_24203,N_21771,N_22373);
nor U24204 (N_24204,N_20059,N_20713);
nor U24205 (N_24205,N_22041,N_22133);
and U24206 (N_24206,N_20094,N_20157);
nor U24207 (N_24207,N_21844,N_20981);
and U24208 (N_24208,N_22478,N_20117);
xor U24209 (N_24209,N_21557,N_22091);
nand U24210 (N_24210,N_22289,N_21513);
xor U24211 (N_24211,N_21864,N_20502);
nor U24212 (N_24212,N_21287,N_20304);
or U24213 (N_24213,N_22479,N_21559);
nor U24214 (N_24214,N_20892,N_20717);
or U24215 (N_24215,N_21704,N_20272);
xor U24216 (N_24216,N_21742,N_21602);
xor U24217 (N_24217,N_22046,N_22420);
nand U24218 (N_24218,N_20542,N_21100);
nor U24219 (N_24219,N_20228,N_20482);
and U24220 (N_24220,N_21779,N_21862);
or U24221 (N_24221,N_21282,N_21674);
nand U24222 (N_24222,N_22336,N_21119);
nand U24223 (N_24223,N_21173,N_21186);
nor U24224 (N_24224,N_21242,N_21326);
and U24225 (N_24225,N_22341,N_21946);
nand U24226 (N_24226,N_20489,N_21162);
and U24227 (N_24227,N_22042,N_21439);
nor U24228 (N_24228,N_21858,N_22044);
or U24229 (N_24229,N_20318,N_20676);
nor U24230 (N_24230,N_20619,N_21088);
nor U24231 (N_24231,N_20471,N_21393);
and U24232 (N_24232,N_22435,N_20986);
or U24233 (N_24233,N_20729,N_21624);
or U24234 (N_24234,N_20476,N_21144);
nor U24235 (N_24235,N_21769,N_22314);
nand U24236 (N_24236,N_22485,N_22192);
xnor U24237 (N_24237,N_22028,N_21773);
xnor U24238 (N_24238,N_20955,N_20067);
or U24239 (N_24239,N_22158,N_20909);
nor U24240 (N_24240,N_20172,N_20346);
nand U24241 (N_24241,N_20650,N_22039);
nand U24242 (N_24242,N_21432,N_21128);
nor U24243 (N_24243,N_20203,N_21126);
nand U24244 (N_24244,N_21597,N_21132);
or U24245 (N_24245,N_21794,N_22401);
nor U24246 (N_24246,N_20750,N_20605);
nor U24247 (N_24247,N_22162,N_20005);
nand U24248 (N_24248,N_22170,N_20767);
or U24249 (N_24249,N_21921,N_22342);
nor U24250 (N_24250,N_20305,N_20839);
and U24251 (N_24251,N_21524,N_20090);
or U24252 (N_24252,N_22001,N_20331);
and U24253 (N_24253,N_21179,N_21407);
nor U24254 (N_24254,N_22432,N_20458);
xnor U24255 (N_24255,N_21351,N_22131);
or U24256 (N_24256,N_21762,N_21945);
or U24257 (N_24257,N_22407,N_20153);
nand U24258 (N_24258,N_21359,N_21416);
nor U24259 (N_24259,N_20622,N_21421);
nor U24260 (N_24260,N_20789,N_20188);
or U24261 (N_24261,N_21404,N_20654);
xor U24262 (N_24262,N_20556,N_21179);
and U24263 (N_24263,N_22288,N_22168);
nor U24264 (N_24264,N_21677,N_21095);
or U24265 (N_24265,N_21528,N_20439);
or U24266 (N_24266,N_20857,N_21330);
nand U24267 (N_24267,N_21242,N_21112);
and U24268 (N_24268,N_21472,N_22381);
and U24269 (N_24269,N_21480,N_22019);
xnor U24270 (N_24270,N_21756,N_20874);
nor U24271 (N_24271,N_21234,N_21068);
or U24272 (N_24272,N_20265,N_22233);
nor U24273 (N_24273,N_21297,N_20508);
and U24274 (N_24274,N_21034,N_20961);
and U24275 (N_24275,N_21384,N_20480);
xor U24276 (N_24276,N_20931,N_20833);
nor U24277 (N_24277,N_20964,N_20133);
nand U24278 (N_24278,N_21957,N_21826);
and U24279 (N_24279,N_21348,N_21830);
xor U24280 (N_24280,N_22313,N_22026);
and U24281 (N_24281,N_22384,N_21440);
nor U24282 (N_24282,N_20226,N_22390);
nor U24283 (N_24283,N_21417,N_20470);
or U24284 (N_24284,N_20772,N_22043);
nor U24285 (N_24285,N_21057,N_21106);
and U24286 (N_24286,N_21941,N_22198);
nand U24287 (N_24287,N_21787,N_20299);
nand U24288 (N_24288,N_21843,N_20265);
nor U24289 (N_24289,N_20984,N_21491);
and U24290 (N_24290,N_22272,N_21073);
nor U24291 (N_24291,N_22108,N_21175);
nor U24292 (N_24292,N_22235,N_22186);
xnor U24293 (N_24293,N_20189,N_21818);
or U24294 (N_24294,N_20243,N_20572);
or U24295 (N_24295,N_21957,N_21885);
and U24296 (N_24296,N_21670,N_20273);
nand U24297 (N_24297,N_20409,N_20841);
nor U24298 (N_24298,N_21980,N_20339);
nor U24299 (N_24299,N_20068,N_20709);
nand U24300 (N_24300,N_20452,N_20123);
nor U24301 (N_24301,N_21321,N_20761);
nand U24302 (N_24302,N_20555,N_20256);
or U24303 (N_24303,N_20569,N_21290);
nor U24304 (N_24304,N_20723,N_21228);
and U24305 (N_24305,N_22142,N_20653);
or U24306 (N_24306,N_21772,N_20938);
xnor U24307 (N_24307,N_21526,N_21495);
nand U24308 (N_24308,N_21275,N_21540);
or U24309 (N_24309,N_20459,N_21544);
nand U24310 (N_24310,N_20429,N_22255);
and U24311 (N_24311,N_20029,N_20213);
xnor U24312 (N_24312,N_22474,N_21399);
nand U24313 (N_24313,N_21503,N_21080);
and U24314 (N_24314,N_21091,N_20422);
and U24315 (N_24315,N_20801,N_22250);
or U24316 (N_24316,N_20633,N_21998);
and U24317 (N_24317,N_22421,N_22274);
nor U24318 (N_24318,N_21465,N_22247);
and U24319 (N_24319,N_21304,N_20378);
nor U24320 (N_24320,N_21007,N_21575);
and U24321 (N_24321,N_20408,N_21822);
nor U24322 (N_24322,N_21327,N_20507);
nand U24323 (N_24323,N_20609,N_21461);
and U24324 (N_24324,N_21627,N_21528);
nor U24325 (N_24325,N_20750,N_21823);
nand U24326 (N_24326,N_20188,N_21877);
or U24327 (N_24327,N_21560,N_21374);
nor U24328 (N_24328,N_21550,N_21320);
or U24329 (N_24329,N_21235,N_21017);
xor U24330 (N_24330,N_21222,N_21368);
nand U24331 (N_24331,N_22494,N_20152);
or U24332 (N_24332,N_21385,N_20116);
nand U24333 (N_24333,N_22093,N_21207);
and U24334 (N_24334,N_22232,N_22346);
and U24335 (N_24335,N_21163,N_20358);
and U24336 (N_24336,N_21026,N_20295);
or U24337 (N_24337,N_22485,N_20695);
xor U24338 (N_24338,N_20365,N_21409);
nand U24339 (N_24339,N_20671,N_22401);
or U24340 (N_24340,N_20677,N_21962);
nand U24341 (N_24341,N_22159,N_20304);
or U24342 (N_24342,N_21047,N_22154);
and U24343 (N_24343,N_22362,N_21534);
nand U24344 (N_24344,N_20021,N_20479);
and U24345 (N_24345,N_22395,N_22327);
nor U24346 (N_24346,N_21341,N_22065);
nand U24347 (N_24347,N_21915,N_22326);
or U24348 (N_24348,N_20999,N_22371);
nand U24349 (N_24349,N_22192,N_21815);
nor U24350 (N_24350,N_21286,N_22451);
or U24351 (N_24351,N_20776,N_20007);
and U24352 (N_24352,N_20577,N_21790);
nand U24353 (N_24353,N_20527,N_20369);
and U24354 (N_24354,N_20967,N_22435);
nor U24355 (N_24355,N_20079,N_21567);
xor U24356 (N_24356,N_20435,N_20182);
xnor U24357 (N_24357,N_21749,N_22195);
nor U24358 (N_24358,N_20537,N_21979);
nor U24359 (N_24359,N_20345,N_20852);
or U24360 (N_24360,N_21595,N_22072);
nor U24361 (N_24361,N_20336,N_20053);
and U24362 (N_24362,N_21124,N_21549);
or U24363 (N_24363,N_20553,N_21060);
nand U24364 (N_24364,N_21682,N_21199);
and U24365 (N_24365,N_20060,N_22353);
nor U24366 (N_24366,N_20456,N_20091);
and U24367 (N_24367,N_21853,N_21427);
nor U24368 (N_24368,N_21281,N_20935);
and U24369 (N_24369,N_20188,N_21463);
and U24370 (N_24370,N_21796,N_21892);
and U24371 (N_24371,N_20550,N_21447);
or U24372 (N_24372,N_22319,N_21633);
or U24373 (N_24373,N_20558,N_21896);
nand U24374 (N_24374,N_22075,N_20875);
nor U24375 (N_24375,N_20793,N_20487);
nand U24376 (N_24376,N_21600,N_22306);
xor U24377 (N_24377,N_20774,N_21074);
and U24378 (N_24378,N_21571,N_21841);
and U24379 (N_24379,N_21695,N_20978);
and U24380 (N_24380,N_21352,N_20787);
or U24381 (N_24381,N_21675,N_22454);
and U24382 (N_24382,N_21918,N_20854);
or U24383 (N_24383,N_21067,N_20861);
nand U24384 (N_24384,N_21746,N_21731);
and U24385 (N_24385,N_22045,N_20322);
nor U24386 (N_24386,N_22485,N_21322);
and U24387 (N_24387,N_20706,N_20999);
nand U24388 (N_24388,N_21319,N_20001);
xnor U24389 (N_24389,N_20463,N_22240);
nor U24390 (N_24390,N_21402,N_20897);
nor U24391 (N_24391,N_21663,N_22003);
nor U24392 (N_24392,N_21892,N_21881);
nor U24393 (N_24393,N_21556,N_20093);
xnor U24394 (N_24394,N_21547,N_21642);
nand U24395 (N_24395,N_20857,N_22219);
nor U24396 (N_24396,N_21326,N_20724);
xor U24397 (N_24397,N_21923,N_21213);
and U24398 (N_24398,N_21317,N_20953);
or U24399 (N_24399,N_22347,N_20948);
or U24400 (N_24400,N_20235,N_20410);
nand U24401 (N_24401,N_21694,N_20045);
xnor U24402 (N_24402,N_21243,N_20806);
nand U24403 (N_24403,N_20846,N_21128);
nand U24404 (N_24404,N_20245,N_20224);
nand U24405 (N_24405,N_20869,N_20325);
and U24406 (N_24406,N_22184,N_20093);
or U24407 (N_24407,N_21565,N_22338);
nand U24408 (N_24408,N_22239,N_21731);
or U24409 (N_24409,N_20683,N_21701);
or U24410 (N_24410,N_20681,N_20574);
nor U24411 (N_24411,N_20880,N_20203);
nor U24412 (N_24412,N_22152,N_20878);
nand U24413 (N_24413,N_22054,N_22101);
xnor U24414 (N_24414,N_20494,N_20047);
and U24415 (N_24415,N_21547,N_20601);
nor U24416 (N_24416,N_20615,N_20587);
xor U24417 (N_24417,N_20419,N_21494);
or U24418 (N_24418,N_21395,N_20564);
nor U24419 (N_24419,N_21756,N_20212);
nor U24420 (N_24420,N_20613,N_22438);
nor U24421 (N_24421,N_21056,N_22367);
nand U24422 (N_24422,N_20045,N_22392);
nand U24423 (N_24423,N_21939,N_21023);
and U24424 (N_24424,N_20870,N_20801);
nand U24425 (N_24425,N_20101,N_21003);
nor U24426 (N_24426,N_22196,N_20618);
nor U24427 (N_24427,N_21783,N_21528);
and U24428 (N_24428,N_21212,N_21228);
and U24429 (N_24429,N_20321,N_20523);
or U24430 (N_24430,N_21075,N_20753);
and U24431 (N_24431,N_21743,N_22201);
xnor U24432 (N_24432,N_20545,N_20181);
and U24433 (N_24433,N_20603,N_20857);
nor U24434 (N_24434,N_20630,N_20838);
nor U24435 (N_24435,N_21513,N_21230);
or U24436 (N_24436,N_20001,N_21942);
or U24437 (N_24437,N_20255,N_20413);
and U24438 (N_24438,N_22159,N_20850);
or U24439 (N_24439,N_22263,N_20010);
nand U24440 (N_24440,N_20875,N_21155);
and U24441 (N_24441,N_21272,N_20697);
and U24442 (N_24442,N_20442,N_21881);
or U24443 (N_24443,N_21914,N_20519);
or U24444 (N_24444,N_20336,N_21523);
and U24445 (N_24445,N_21654,N_21047);
nand U24446 (N_24446,N_21027,N_22382);
nor U24447 (N_24447,N_21906,N_21881);
nand U24448 (N_24448,N_20801,N_20995);
or U24449 (N_24449,N_20486,N_21952);
and U24450 (N_24450,N_20932,N_21052);
or U24451 (N_24451,N_20842,N_21488);
nand U24452 (N_24452,N_20343,N_20026);
nor U24453 (N_24453,N_21771,N_22004);
nand U24454 (N_24454,N_22498,N_20713);
xnor U24455 (N_24455,N_21242,N_21713);
or U24456 (N_24456,N_22434,N_22311);
nor U24457 (N_24457,N_20101,N_21986);
and U24458 (N_24458,N_20400,N_21091);
nand U24459 (N_24459,N_22189,N_20561);
xor U24460 (N_24460,N_21568,N_20329);
nor U24461 (N_24461,N_21673,N_20718);
xnor U24462 (N_24462,N_21508,N_20446);
nand U24463 (N_24463,N_22437,N_21001);
xor U24464 (N_24464,N_20287,N_20684);
or U24465 (N_24465,N_21647,N_20999);
nor U24466 (N_24466,N_21943,N_20322);
or U24467 (N_24467,N_20561,N_21918);
nand U24468 (N_24468,N_20939,N_22015);
or U24469 (N_24469,N_21132,N_22362);
and U24470 (N_24470,N_20907,N_21780);
and U24471 (N_24471,N_21235,N_22117);
nand U24472 (N_24472,N_20769,N_20381);
nor U24473 (N_24473,N_22296,N_21103);
or U24474 (N_24474,N_21089,N_21898);
nor U24475 (N_24475,N_20289,N_21008);
or U24476 (N_24476,N_20660,N_20798);
and U24477 (N_24477,N_20950,N_20015);
or U24478 (N_24478,N_21808,N_20009);
or U24479 (N_24479,N_20019,N_22267);
or U24480 (N_24480,N_21506,N_20807);
nor U24481 (N_24481,N_22216,N_20696);
or U24482 (N_24482,N_22472,N_22436);
xor U24483 (N_24483,N_20475,N_21887);
or U24484 (N_24484,N_21282,N_22293);
or U24485 (N_24485,N_21292,N_20719);
xnor U24486 (N_24486,N_20181,N_21479);
xnor U24487 (N_24487,N_21441,N_20346);
nand U24488 (N_24488,N_22249,N_20579);
or U24489 (N_24489,N_22004,N_20545);
nor U24490 (N_24490,N_20109,N_21015);
nor U24491 (N_24491,N_20589,N_21324);
and U24492 (N_24492,N_20632,N_21474);
xor U24493 (N_24493,N_20461,N_20133);
or U24494 (N_24494,N_21805,N_20776);
xnor U24495 (N_24495,N_20215,N_20570);
and U24496 (N_24496,N_20778,N_20063);
and U24497 (N_24497,N_22174,N_20430);
nand U24498 (N_24498,N_20170,N_20748);
nor U24499 (N_24499,N_21743,N_20731);
nand U24500 (N_24500,N_22234,N_21108);
xnor U24501 (N_24501,N_21842,N_21795);
nor U24502 (N_24502,N_20563,N_21779);
nand U24503 (N_24503,N_21886,N_20619);
nand U24504 (N_24504,N_20910,N_21979);
or U24505 (N_24505,N_21641,N_21935);
nand U24506 (N_24506,N_20562,N_20652);
or U24507 (N_24507,N_21048,N_20501);
and U24508 (N_24508,N_20824,N_20392);
or U24509 (N_24509,N_22172,N_21106);
or U24510 (N_24510,N_20818,N_20104);
nor U24511 (N_24511,N_20290,N_22231);
nand U24512 (N_24512,N_22325,N_20937);
nor U24513 (N_24513,N_22488,N_20564);
or U24514 (N_24514,N_20206,N_21207);
nor U24515 (N_24515,N_22398,N_21440);
and U24516 (N_24516,N_20238,N_21412);
nand U24517 (N_24517,N_22212,N_20519);
or U24518 (N_24518,N_22055,N_21399);
nor U24519 (N_24519,N_20811,N_21741);
xor U24520 (N_24520,N_20850,N_22371);
nor U24521 (N_24521,N_21482,N_22345);
nor U24522 (N_24522,N_21739,N_21666);
or U24523 (N_24523,N_21102,N_20120);
nor U24524 (N_24524,N_20710,N_20026);
and U24525 (N_24525,N_21152,N_20048);
nand U24526 (N_24526,N_20808,N_21620);
nor U24527 (N_24527,N_22226,N_20485);
and U24528 (N_24528,N_21086,N_20290);
xor U24529 (N_24529,N_20993,N_20661);
or U24530 (N_24530,N_21899,N_20295);
and U24531 (N_24531,N_21180,N_20637);
xor U24532 (N_24532,N_20319,N_21135);
or U24533 (N_24533,N_21130,N_21778);
nor U24534 (N_24534,N_21345,N_20831);
and U24535 (N_24535,N_21376,N_21592);
nand U24536 (N_24536,N_21682,N_20080);
and U24537 (N_24537,N_22133,N_20402);
and U24538 (N_24538,N_22336,N_21308);
xnor U24539 (N_24539,N_20223,N_22438);
or U24540 (N_24540,N_21682,N_21641);
nor U24541 (N_24541,N_22108,N_21161);
and U24542 (N_24542,N_22119,N_20316);
or U24543 (N_24543,N_21833,N_21378);
nor U24544 (N_24544,N_20597,N_20933);
nor U24545 (N_24545,N_21920,N_20503);
xor U24546 (N_24546,N_20783,N_20604);
xnor U24547 (N_24547,N_20298,N_20156);
xor U24548 (N_24548,N_22241,N_21220);
or U24549 (N_24549,N_20965,N_21022);
or U24550 (N_24550,N_20131,N_20469);
or U24551 (N_24551,N_22125,N_21587);
xnor U24552 (N_24552,N_21871,N_20753);
nand U24553 (N_24553,N_20356,N_20146);
and U24554 (N_24554,N_21959,N_21629);
xor U24555 (N_24555,N_21785,N_20922);
nor U24556 (N_24556,N_20123,N_21066);
nand U24557 (N_24557,N_20969,N_21843);
nor U24558 (N_24558,N_20849,N_21932);
or U24559 (N_24559,N_21936,N_20115);
nor U24560 (N_24560,N_21787,N_20614);
xnor U24561 (N_24561,N_20644,N_21602);
and U24562 (N_24562,N_20058,N_20698);
and U24563 (N_24563,N_21102,N_21173);
or U24564 (N_24564,N_20171,N_22457);
or U24565 (N_24565,N_21584,N_20964);
nor U24566 (N_24566,N_21672,N_20153);
and U24567 (N_24567,N_20554,N_20546);
xor U24568 (N_24568,N_21614,N_21415);
nor U24569 (N_24569,N_20862,N_21757);
or U24570 (N_24570,N_21654,N_20100);
and U24571 (N_24571,N_21004,N_21922);
and U24572 (N_24572,N_21418,N_20013);
nand U24573 (N_24573,N_20477,N_20780);
xor U24574 (N_24574,N_21706,N_20513);
xor U24575 (N_24575,N_21729,N_20252);
nand U24576 (N_24576,N_22080,N_21545);
nor U24577 (N_24577,N_20719,N_20951);
and U24578 (N_24578,N_20118,N_21041);
or U24579 (N_24579,N_21115,N_21412);
or U24580 (N_24580,N_20355,N_20868);
xnor U24581 (N_24581,N_22056,N_21700);
or U24582 (N_24582,N_21332,N_20177);
xnor U24583 (N_24583,N_21524,N_22086);
nand U24584 (N_24584,N_21189,N_21736);
xor U24585 (N_24585,N_20964,N_22378);
nor U24586 (N_24586,N_20710,N_21627);
nor U24587 (N_24587,N_20969,N_21264);
and U24588 (N_24588,N_20585,N_21418);
nor U24589 (N_24589,N_20275,N_21792);
and U24590 (N_24590,N_22161,N_21971);
and U24591 (N_24591,N_22026,N_20909);
nand U24592 (N_24592,N_21497,N_22409);
nand U24593 (N_24593,N_20269,N_20053);
xnor U24594 (N_24594,N_20418,N_22078);
and U24595 (N_24595,N_20025,N_22387);
nor U24596 (N_24596,N_21192,N_21623);
or U24597 (N_24597,N_20023,N_22245);
xnor U24598 (N_24598,N_21275,N_20482);
nor U24599 (N_24599,N_20141,N_22023);
or U24600 (N_24600,N_21256,N_21279);
xnor U24601 (N_24601,N_20060,N_20694);
xnor U24602 (N_24602,N_20695,N_21366);
nand U24603 (N_24603,N_20032,N_21657);
nand U24604 (N_24604,N_22024,N_20649);
nor U24605 (N_24605,N_22348,N_20434);
nand U24606 (N_24606,N_21486,N_21435);
and U24607 (N_24607,N_22286,N_20898);
and U24608 (N_24608,N_21347,N_20684);
xor U24609 (N_24609,N_21488,N_21328);
nand U24610 (N_24610,N_22074,N_22236);
or U24611 (N_24611,N_20914,N_20999);
nand U24612 (N_24612,N_22344,N_21008);
nand U24613 (N_24613,N_20977,N_21469);
xnor U24614 (N_24614,N_20623,N_21141);
and U24615 (N_24615,N_22054,N_22041);
and U24616 (N_24616,N_22450,N_20067);
xor U24617 (N_24617,N_21158,N_21987);
or U24618 (N_24618,N_20516,N_21141);
or U24619 (N_24619,N_20834,N_21814);
nor U24620 (N_24620,N_21609,N_21176);
and U24621 (N_24621,N_20735,N_21891);
or U24622 (N_24622,N_20556,N_20244);
nor U24623 (N_24623,N_21584,N_20182);
nand U24624 (N_24624,N_22396,N_20109);
or U24625 (N_24625,N_21045,N_20840);
nor U24626 (N_24626,N_21095,N_21757);
or U24627 (N_24627,N_20778,N_20202);
or U24628 (N_24628,N_21994,N_20291);
or U24629 (N_24629,N_20747,N_21893);
nor U24630 (N_24630,N_20199,N_21101);
and U24631 (N_24631,N_22112,N_21374);
or U24632 (N_24632,N_22331,N_20341);
or U24633 (N_24633,N_21459,N_20330);
xnor U24634 (N_24634,N_21789,N_20567);
and U24635 (N_24635,N_21164,N_21290);
nand U24636 (N_24636,N_21924,N_22386);
and U24637 (N_24637,N_20215,N_20598);
nand U24638 (N_24638,N_20083,N_21686);
nand U24639 (N_24639,N_21338,N_20655);
nand U24640 (N_24640,N_21029,N_22247);
nand U24641 (N_24641,N_20460,N_22312);
and U24642 (N_24642,N_20688,N_21715);
or U24643 (N_24643,N_21859,N_21610);
and U24644 (N_24644,N_21707,N_22365);
and U24645 (N_24645,N_22452,N_20374);
or U24646 (N_24646,N_20130,N_20395);
and U24647 (N_24647,N_20915,N_22008);
xnor U24648 (N_24648,N_20573,N_22282);
or U24649 (N_24649,N_21663,N_20161);
nand U24650 (N_24650,N_22060,N_20709);
nand U24651 (N_24651,N_20900,N_21780);
and U24652 (N_24652,N_20956,N_20203);
and U24653 (N_24653,N_21103,N_20058);
nor U24654 (N_24654,N_21194,N_20987);
nor U24655 (N_24655,N_22083,N_20172);
xnor U24656 (N_24656,N_20833,N_20810);
nand U24657 (N_24657,N_21524,N_22497);
and U24658 (N_24658,N_22035,N_21357);
and U24659 (N_24659,N_22282,N_20692);
nor U24660 (N_24660,N_20566,N_20381);
nor U24661 (N_24661,N_21700,N_20934);
nor U24662 (N_24662,N_21220,N_22247);
nand U24663 (N_24663,N_20635,N_20864);
or U24664 (N_24664,N_20856,N_21205);
nor U24665 (N_24665,N_21340,N_20426);
nand U24666 (N_24666,N_20925,N_20332);
or U24667 (N_24667,N_21146,N_20613);
nand U24668 (N_24668,N_20495,N_22264);
or U24669 (N_24669,N_21066,N_22254);
nor U24670 (N_24670,N_20523,N_21623);
or U24671 (N_24671,N_20987,N_20741);
nor U24672 (N_24672,N_21667,N_20634);
nor U24673 (N_24673,N_20959,N_21934);
nand U24674 (N_24674,N_20733,N_21979);
or U24675 (N_24675,N_20957,N_20733);
or U24676 (N_24676,N_20809,N_21219);
nor U24677 (N_24677,N_22032,N_21529);
or U24678 (N_24678,N_20923,N_20742);
or U24679 (N_24679,N_20912,N_20532);
nor U24680 (N_24680,N_21132,N_20184);
nor U24681 (N_24681,N_21354,N_22314);
nand U24682 (N_24682,N_21059,N_20072);
nand U24683 (N_24683,N_20796,N_20206);
and U24684 (N_24684,N_20865,N_20751);
and U24685 (N_24685,N_21218,N_21605);
and U24686 (N_24686,N_20906,N_21510);
nor U24687 (N_24687,N_21374,N_22348);
or U24688 (N_24688,N_22245,N_21450);
xor U24689 (N_24689,N_21047,N_21532);
nand U24690 (N_24690,N_20122,N_20982);
nor U24691 (N_24691,N_20783,N_20311);
nand U24692 (N_24692,N_22428,N_21273);
xnor U24693 (N_24693,N_20992,N_21594);
nor U24694 (N_24694,N_21364,N_21528);
and U24695 (N_24695,N_21777,N_21280);
and U24696 (N_24696,N_21723,N_22222);
nor U24697 (N_24697,N_21689,N_21785);
and U24698 (N_24698,N_20354,N_20360);
nor U24699 (N_24699,N_20876,N_20203);
or U24700 (N_24700,N_21938,N_22475);
or U24701 (N_24701,N_20754,N_22262);
nand U24702 (N_24702,N_22078,N_20168);
nand U24703 (N_24703,N_20983,N_20544);
and U24704 (N_24704,N_21324,N_20191);
nand U24705 (N_24705,N_21138,N_20456);
and U24706 (N_24706,N_20063,N_20948);
and U24707 (N_24707,N_21791,N_21217);
and U24708 (N_24708,N_21695,N_22081);
and U24709 (N_24709,N_20120,N_20145);
nand U24710 (N_24710,N_21341,N_22475);
xor U24711 (N_24711,N_20558,N_20305);
and U24712 (N_24712,N_21817,N_22228);
xor U24713 (N_24713,N_22430,N_22025);
nor U24714 (N_24714,N_21962,N_22257);
nand U24715 (N_24715,N_20519,N_20060);
or U24716 (N_24716,N_20983,N_20272);
nand U24717 (N_24717,N_21896,N_21078);
and U24718 (N_24718,N_21134,N_22042);
nand U24719 (N_24719,N_22204,N_21183);
and U24720 (N_24720,N_22265,N_22274);
or U24721 (N_24721,N_21179,N_22280);
nand U24722 (N_24722,N_20633,N_21662);
and U24723 (N_24723,N_21421,N_20744);
xor U24724 (N_24724,N_22135,N_20701);
or U24725 (N_24725,N_20909,N_22230);
or U24726 (N_24726,N_22160,N_21008);
nor U24727 (N_24727,N_21146,N_20614);
or U24728 (N_24728,N_22098,N_21092);
nor U24729 (N_24729,N_21438,N_21892);
or U24730 (N_24730,N_20072,N_20129);
nand U24731 (N_24731,N_20847,N_21558);
or U24732 (N_24732,N_20481,N_22433);
or U24733 (N_24733,N_20101,N_20701);
nor U24734 (N_24734,N_20139,N_20452);
nand U24735 (N_24735,N_22415,N_20287);
and U24736 (N_24736,N_20574,N_21508);
and U24737 (N_24737,N_22381,N_21266);
or U24738 (N_24738,N_20492,N_21975);
and U24739 (N_24739,N_22447,N_20229);
and U24740 (N_24740,N_21289,N_21934);
nand U24741 (N_24741,N_22250,N_21673);
nor U24742 (N_24742,N_21880,N_22173);
nor U24743 (N_24743,N_20612,N_21002);
and U24744 (N_24744,N_21346,N_21743);
nor U24745 (N_24745,N_21324,N_20829);
nand U24746 (N_24746,N_20824,N_21005);
or U24747 (N_24747,N_21849,N_21673);
or U24748 (N_24748,N_20527,N_21130);
nor U24749 (N_24749,N_20042,N_22426);
nor U24750 (N_24750,N_20709,N_21467);
nand U24751 (N_24751,N_20806,N_21029);
and U24752 (N_24752,N_20841,N_22319);
or U24753 (N_24753,N_20562,N_20677);
xor U24754 (N_24754,N_20031,N_21480);
nor U24755 (N_24755,N_21759,N_21141);
nand U24756 (N_24756,N_21096,N_21539);
nand U24757 (N_24757,N_21006,N_21755);
nand U24758 (N_24758,N_21162,N_20927);
or U24759 (N_24759,N_21654,N_21593);
nor U24760 (N_24760,N_22068,N_22463);
and U24761 (N_24761,N_20818,N_21840);
or U24762 (N_24762,N_21097,N_20963);
and U24763 (N_24763,N_21769,N_21715);
and U24764 (N_24764,N_20746,N_20453);
nor U24765 (N_24765,N_22282,N_20580);
nor U24766 (N_24766,N_20637,N_20356);
or U24767 (N_24767,N_20154,N_22270);
nor U24768 (N_24768,N_20762,N_22047);
or U24769 (N_24769,N_22413,N_21426);
nand U24770 (N_24770,N_22133,N_21699);
or U24771 (N_24771,N_21762,N_21849);
nand U24772 (N_24772,N_22423,N_20999);
and U24773 (N_24773,N_21003,N_21308);
and U24774 (N_24774,N_21355,N_22429);
nand U24775 (N_24775,N_22430,N_20515);
nand U24776 (N_24776,N_20183,N_21019);
and U24777 (N_24777,N_20459,N_21403);
xor U24778 (N_24778,N_22422,N_20904);
and U24779 (N_24779,N_20492,N_21486);
xor U24780 (N_24780,N_21053,N_21825);
and U24781 (N_24781,N_20150,N_21481);
nor U24782 (N_24782,N_22135,N_21352);
nor U24783 (N_24783,N_22349,N_21206);
and U24784 (N_24784,N_20131,N_22041);
nand U24785 (N_24785,N_21139,N_21570);
or U24786 (N_24786,N_20300,N_21920);
and U24787 (N_24787,N_20136,N_21327);
nand U24788 (N_24788,N_20086,N_20535);
nor U24789 (N_24789,N_20417,N_20832);
and U24790 (N_24790,N_20119,N_21163);
and U24791 (N_24791,N_22105,N_21140);
or U24792 (N_24792,N_21017,N_20401);
nand U24793 (N_24793,N_20767,N_21237);
xor U24794 (N_24794,N_21623,N_20548);
nor U24795 (N_24795,N_21553,N_22139);
nor U24796 (N_24796,N_21161,N_21058);
or U24797 (N_24797,N_20538,N_22352);
nand U24798 (N_24798,N_21364,N_20991);
nand U24799 (N_24799,N_20341,N_21704);
or U24800 (N_24800,N_20614,N_20926);
and U24801 (N_24801,N_21301,N_20306);
nand U24802 (N_24802,N_21868,N_22266);
or U24803 (N_24803,N_21335,N_20974);
nor U24804 (N_24804,N_20334,N_22458);
nor U24805 (N_24805,N_21576,N_21949);
nor U24806 (N_24806,N_20029,N_20123);
nand U24807 (N_24807,N_21176,N_22083);
or U24808 (N_24808,N_21173,N_20952);
nor U24809 (N_24809,N_20163,N_22102);
and U24810 (N_24810,N_21865,N_21876);
xnor U24811 (N_24811,N_20893,N_21560);
nand U24812 (N_24812,N_22284,N_21614);
nor U24813 (N_24813,N_21934,N_20776);
and U24814 (N_24814,N_22185,N_21546);
nand U24815 (N_24815,N_20901,N_20533);
nand U24816 (N_24816,N_21298,N_20876);
nor U24817 (N_24817,N_21491,N_20603);
or U24818 (N_24818,N_22392,N_20272);
nor U24819 (N_24819,N_22373,N_20734);
nor U24820 (N_24820,N_20724,N_21321);
xnor U24821 (N_24821,N_21013,N_22092);
nor U24822 (N_24822,N_20710,N_21588);
nor U24823 (N_24823,N_21019,N_21039);
and U24824 (N_24824,N_20376,N_21702);
nor U24825 (N_24825,N_21918,N_22125);
and U24826 (N_24826,N_20538,N_20670);
nor U24827 (N_24827,N_21192,N_20496);
xnor U24828 (N_24828,N_21807,N_22220);
and U24829 (N_24829,N_22053,N_20427);
or U24830 (N_24830,N_20664,N_20644);
and U24831 (N_24831,N_20384,N_20218);
nor U24832 (N_24832,N_20851,N_21486);
nor U24833 (N_24833,N_22172,N_20309);
nor U24834 (N_24834,N_20964,N_22173);
nand U24835 (N_24835,N_21268,N_20549);
xor U24836 (N_24836,N_21949,N_22195);
and U24837 (N_24837,N_20402,N_21019);
nand U24838 (N_24838,N_20109,N_20407);
or U24839 (N_24839,N_21245,N_20801);
nor U24840 (N_24840,N_22261,N_22330);
xor U24841 (N_24841,N_21075,N_21944);
nand U24842 (N_24842,N_21301,N_22291);
or U24843 (N_24843,N_20220,N_20431);
nand U24844 (N_24844,N_21510,N_21729);
nor U24845 (N_24845,N_21660,N_20104);
nand U24846 (N_24846,N_21793,N_21039);
and U24847 (N_24847,N_20293,N_20056);
or U24848 (N_24848,N_21915,N_21157);
xor U24849 (N_24849,N_22040,N_20623);
nor U24850 (N_24850,N_21331,N_22194);
nand U24851 (N_24851,N_21999,N_20532);
nand U24852 (N_24852,N_21230,N_20120);
nand U24853 (N_24853,N_21432,N_21190);
xnor U24854 (N_24854,N_21244,N_21733);
or U24855 (N_24855,N_20836,N_20469);
or U24856 (N_24856,N_21044,N_21805);
nand U24857 (N_24857,N_21789,N_21937);
or U24858 (N_24858,N_20745,N_21168);
and U24859 (N_24859,N_21524,N_21083);
or U24860 (N_24860,N_22469,N_21282);
nor U24861 (N_24861,N_20428,N_21611);
or U24862 (N_24862,N_21471,N_21144);
and U24863 (N_24863,N_20519,N_21315);
and U24864 (N_24864,N_20394,N_21212);
and U24865 (N_24865,N_21697,N_21696);
or U24866 (N_24866,N_20950,N_20183);
nor U24867 (N_24867,N_21914,N_21786);
nor U24868 (N_24868,N_21437,N_20853);
xor U24869 (N_24869,N_21208,N_22273);
and U24870 (N_24870,N_20216,N_20604);
nand U24871 (N_24871,N_21132,N_20628);
nor U24872 (N_24872,N_21772,N_20831);
nor U24873 (N_24873,N_20696,N_20195);
nor U24874 (N_24874,N_20735,N_22346);
nor U24875 (N_24875,N_21269,N_21402);
and U24876 (N_24876,N_20189,N_21998);
or U24877 (N_24877,N_20773,N_21185);
or U24878 (N_24878,N_21822,N_20280);
nand U24879 (N_24879,N_20121,N_22022);
nand U24880 (N_24880,N_21104,N_21331);
xor U24881 (N_24881,N_20353,N_21431);
nand U24882 (N_24882,N_21899,N_22326);
nand U24883 (N_24883,N_20687,N_21334);
nand U24884 (N_24884,N_21764,N_22203);
nand U24885 (N_24885,N_22140,N_21298);
nand U24886 (N_24886,N_21128,N_22467);
xor U24887 (N_24887,N_20747,N_22246);
or U24888 (N_24888,N_21715,N_21110);
and U24889 (N_24889,N_22158,N_21708);
and U24890 (N_24890,N_21054,N_20772);
and U24891 (N_24891,N_21682,N_21501);
or U24892 (N_24892,N_21475,N_21828);
xor U24893 (N_24893,N_20191,N_21621);
xnor U24894 (N_24894,N_20128,N_20527);
nor U24895 (N_24895,N_21081,N_21977);
nand U24896 (N_24896,N_21760,N_20666);
nor U24897 (N_24897,N_21462,N_21216);
nand U24898 (N_24898,N_20243,N_22371);
xnor U24899 (N_24899,N_20697,N_20397);
or U24900 (N_24900,N_20407,N_21372);
nor U24901 (N_24901,N_21714,N_20351);
nor U24902 (N_24902,N_20052,N_20127);
nor U24903 (N_24903,N_21319,N_21549);
nor U24904 (N_24904,N_21084,N_21856);
nor U24905 (N_24905,N_20179,N_20866);
or U24906 (N_24906,N_21244,N_22398);
or U24907 (N_24907,N_20971,N_22103);
nand U24908 (N_24908,N_20203,N_20943);
xor U24909 (N_24909,N_20144,N_20321);
or U24910 (N_24910,N_21507,N_20574);
or U24911 (N_24911,N_20496,N_20063);
nor U24912 (N_24912,N_22032,N_20791);
or U24913 (N_24913,N_21715,N_20518);
and U24914 (N_24914,N_21388,N_20563);
nor U24915 (N_24915,N_22055,N_20270);
nor U24916 (N_24916,N_20857,N_21045);
or U24917 (N_24917,N_20979,N_22019);
xnor U24918 (N_24918,N_20472,N_20190);
and U24919 (N_24919,N_20764,N_20092);
nor U24920 (N_24920,N_20698,N_22280);
nand U24921 (N_24921,N_22415,N_20660);
and U24922 (N_24922,N_21228,N_21733);
xor U24923 (N_24923,N_20150,N_20265);
nor U24924 (N_24924,N_21646,N_22421);
and U24925 (N_24925,N_21941,N_20965);
nor U24926 (N_24926,N_21297,N_21092);
or U24927 (N_24927,N_20659,N_21499);
and U24928 (N_24928,N_21532,N_20156);
nand U24929 (N_24929,N_20616,N_20908);
nor U24930 (N_24930,N_20794,N_20258);
nor U24931 (N_24931,N_21839,N_21423);
xnor U24932 (N_24932,N_22429,N_22042);
nand U24933 (N_24933,N_22335,N_20479);
nand U24934 (N_24934,N_22257,N_20840);
nand U24935 (N_24935,N_20396,N_20000);
nand U24936 (N_24936,N_21536,N_21420);
and U24937 (N_24937,N_22098,N_20972);
nor U24938 (N_24938,N_20252,N_20016);
nor U24939 (N_24939,N_21595,N_22290);
nor U24940 (N_24940,N_20642,N_21475);
nand U24941 (N_24941,N_21802,N_20507);
nand U24942 (N_24942,N_22199,N_20720);
and U24943 (N_24943,N_21102,N_21436);
and U24944 (N_24944,N_20810,N_21591);
nand U24945 (N_24945,N_20067,N_20735);
or U24946 (N_24946,N_20434,N_20240);
or U24947 (N_24947,N_21204,N_20664);
xor U24948 (N_24948,N_20868,N_21913);
or U24949 (N_24949,N_22263,N_21188);
xnor U24950 (N_24950,N_21743,N_21124);
nor U24951 (N_24951,N_22022,N_20898);
nor U24952 (N_24952,N_20718,N_22152);
or U24953 (N_24953,N_22303,N_21540);
xor U24954 (N_24954,N_20478,N_20154);
nand U24955 (N_24955,N_20175,N_22335);
nand U24956 (N_24956,N_20356,N_20389);
nand U24957 (N_24957,N_21008,N_22292);
or U24958 (N_24958,N_22125,N_22221);
nor U24959 (N_24959,N_20096,N_20018);
nor U24960 (N_24960,N_21377,N_20127);
xnor U24961 (N_24961,N_20398,N_20777);
or U24962 (N_24962,N_22086,N_21441);
xnor U24963 (N_24963,N_20528,N_20947);
or U24964 (N_24964,N_20636,N_21311);
nand U24965 (N_24965,N_20535,N_21537);
nor U24966 (N_24966,N_22426,N_20536);
and U24967 (N_24967,N_20243,N_20941);
or U24968 (N_24968,N_21731,N_20444);
xnor U24969 (N_24969,N_21685,N_20969);
xnor U24970 (N_24970,N_22292,N_22228);
nor U24971 (N_24971,N_20155,N_22218);
nand U24972 (N_24972,N_21316,N_21664);
nand U24973 (N_24973,N_20211,N_21727);
nor U24974 (N_24974,N_21119,N_21679);
nand U24975 (N_24975,N_20277,N_21266);
nor U24976 (N_24976,N_21367,N_20500);
nor U24977 (N_24977,N_21446,N_20708);
nor U24978 (N_24978,N_20862,N_22466);
nor U24979 (N_24979,N_20596,N_21659);
and U24980 (N_24980,N_20826,N_20990);
and U24981 (N_24981,N_21463,N_20334);
xnor U24982 (N_24982,N_20783,N_20273);
nand U24983 (N_24983,N_22435,N_20990);
nand U24984 (N_24984,N_21937,N_21673);
or U24985 (N_24985,N_20003,N_20391);
nand U24986 (N_24986,N_22390,N_22312);
nand U24987 (N_24987,N_20876,N_22025);
nor U24988 (N_24988,N_20259,N_21043);
nand U24989 (N_24989,N_20672,N_22328);
and U24990 (N_24990,N_20193,N_20874);
or U24991 (N_24991,N_21032,N_20624);
nand U24992 (N_24992,N_20367,N_20689);
or U24993 (N_24993,N_20272,N_20845);
or U24994 (N_24994,N_20178,N_21946);
nand U24995 (N_24995,N_21711,N_21547);
nor U24996 (N_24996,N_22098,N_21311);
or U24997 (N_24997,N_20584,N_21415);
xor U24998 (N_24998,N_21275,N_20131);
nor U24999 (N_24999,N_21010,N_21513);
xnor UO_0 (O_0,N_24043,N_22642);
or UO_1 (O_1,N_24485,N_22822);
nor UO_2 (O_2,N_24710,N_24349);
nand UO_3 (O_3,N_23545,N_24543);
nor UO_4 (O_4,N_23023,N_22757);
and UO_5 (O_5,N_24199,N_24898);
nor UO_6 (O_6,N_22789,N_23221);
or UO_7 (O_7,N_23534,N_22674);
nor UO_8 (O_8,N_24409,N_23609);
nand UO_9 (O_9,N_23366,N_24525);
nand UO_10 (O_10,N_23590,N_23479);
or UO_11 (O_11,N_24138,N_23163);
nand UO_12 (O_12,N_23785,N_23835);
nand UO_13 (O_13,N_23076,N_23304);
nor UO_14 (O_14,N_24125,N_24445);
nor UO_15 (O_15,N_23819,N_24562);
and UO_16 (O_16,N_23034,N_22860);
nor UO_17 (O_17,N_24474,N_24900);
nand UO_18 (O_18,N_24164,N_22929);
xnor UO_19 (O_19,N_24756,N_24537);
xnor UO_20 (O_20,N_22546,N_23962);
nor UO_21 (O_21,N_22670,N_24874);
nor UO_22 (O_22,N_24890,N_24931);
xor UO_23 (O_23,N_23056,N_23311);
xnor UO_24 (O_24,N_24960,N_24886);
nor UO_25 (O_25,N_23980,N_24149);
nand UO_26 (O_26,N_24654,N_24581);
nor UO_27 (O_27,N_22570,N_23741);
xor UO_28 (O_28,N_24006,N_24820);
or UO_29 (O_29,N_24288,N_24652);
or UO_30 (O_30,N_24675,N_23910);
nor UO_31 (O_31,N_23321,N_24774);
or UO_32 (O_32,N_23569,N_22951);
and UO_33 (O_33,N_23503,N_24375);
and UO_34 (O_34,N_24056,N_24594);
and UO_35 (O_35,N_22797,N_22650);
xnor UO_36 (O_36,N_23963,N_22631);
nand UO_37 (O_37,N_23296,N_24081);
and UO_38 (O_38,N_22742,N_24992);
or UO_39 (O_39,N_24230,N_24792);
nor UO_40 (O_40,N_24294,N_22850);
nor UO_41 (O_41,N_23426,N_24722);
or UO_42 (O_42,N_23533,N_24600);
and UO_43 (O_43,N_24868,N_24996);
nand UO_44 (O_44,N_24951,N_23228);
nor UO_45 (O_45,N_24106,N_23515);
nor UO_46 (O_46,N_23816,N_24200);
nor UO_47 (O_47,N_23803,N_23710);
nand UO_48 (O_48,N_22873,N_22535);
or UO_49 (O_49,N_24546,N_24626);
or UO_50 (O_50,N_22738,N_23795);
nand UO_51 (O_51,N_24049,N_24913);
nand UO_52 (O_52,N_23331,N_24287);
and UO_53 (O_53,N_24788,N_22920);
nand UO_54 (O_54,N_24716,N_22618);
nand UO_55 (O_55,N_24887,N_23634);
and UO_56 (O_56,N_23498,N_24823);
nand UO_57 (O_57,N_24905,N_22507);
and UO_58 (O_58,N_24865,N_23755);
nand UO_59 (O_59,N_24994,N_23812);
nand UO_60 (O_60,N_23367,N_23520);
and UO_61 (O_61,N_24757,N_23011);
nand UO_62 (O_62,N_24100,N_23415);
xnor UO_63 (O_63,N_22500,N_24266);
and UO_64 (O_64,N_23390,N_24773);
or UO_65 (O_65,N_23668,N_23138);
nand UO_66 (O_66,N_23243,N_24759);
nor UO_67 (O_67,N_24233,N_22820);
or UO_68 (O_68,N_23985,N_22902);
nor UO_69 (O_69,N_23172,N_22761);
nand UO_70 (O_70,N_23645,N_22914);
or UO_71 (O_71,N_24531,N_24231);
and UO_72 (O_72,N_24143,N_24065);
nor UO_73 (O_73,N_24433,N_23414);
and UO_74 (O_74,N_24080,N_24240);
xor UO_75 (O_75,N_24393,N_23052);
nor UO_76 (O_76,N_24596,N_24037);
xnor UO_77 (O_77,N_23909,N_24893);
nand UO_78 (O_78,N_23706,N_22526);
or UO_79 (O_79,N_24320,N_23627);
or UO_80 (O_80,N_24454,N_23767);
nand UO_81 (O_81,N_24019,N_23310);
or UO_82 (O_82,N_22806,N_23689);
nor UO_83 (O_83,N_23799,N_23324);
nand UO_84 (O_84,N_24793,N_22938);
nand UO_85 (O_85,N_23975,N_23732);
nor UO_86 (O_86,N_24153,N_24567);
or UO_87 (O_87,N_23416,N_23356);
or UO_88 (O_88,N_22973,N_23912);
and UO_89 (O_89,N_22972,N_22994);
or UO_90 (O_90,N_24990,N_23670);
or UO_91 (O_91,N_23961,N_24140);
nor UO_92 (O_92,N_23920,N_22961);
nor UO_93 (O_93,N_23407,N_24361);
or UO_94 (O_94,N_24585,N_24145);
and UO_95 (O_95,N_23073,N_23192);
nor UO_96 (O_96,N_22781,N_24509);
nand UO_97 (O_97,N_24155,N_22644);
xnor UO_98 (O_98,N_23094,N_23821);
or UO_99 (O_99,N_24933,N_24502);
nand UO_100 (O_100,N_22866,N_22950);
nand UO_101 (O_101,N_23062,N_23022);
nor UO_102 (O_102,N_23919,N_23477);
nand UO_103 (O_103,N_23200,N_24306);
nor UO_104 (O_104,N_24673,N_24391);
or UO_105 (O_105,N_22949,N_24711);
nor UO_106 (O_106,N_23431,N_23487);
nand UO_107 (O_107,N_24434,N_24536);
nor UO_108 (O_108,N_23838,N_22732);
xnor UO_109 (O_109,N_23594,N_24208);
nor UO_110 (O_110,N_23804,N_22900);
nor UO_111 (O_111,N_23002,N_24246);
nor UO_112 (O_112,N_23203,N_24210);
and UO_113 (O_113,N_23420,N_22964);
nor UO_114 (O_114,N_23731,N_23169);
nor UO_115 (O_115,N_24338,N_23901);
or UO_116 (O_116,N_24250,N_23378);
and UO_117 (O_117,N_23644,N_22921);
or UO_118 (O_118,N_22672,N_24656);
nor UO_119 (O_119,N_23796,N_23990);
nand UO_120 (O_120,N_24051,N_24794);
nor UO_121 (O_121,N_24269,N_23944);
and UO_122 (O_122,N_24264,N_24787);
or UO_123 (O_123,N_24091,N_24331);
nand UO_124 (O_124,N_24571,N_23233);
nand UO_125 (O_125,N_24182,N_23623);
xor UO_126 (O_126,N_23862,N_23204);
and UO_127 (O_127,N_23016,N_24504);
nand UO_128 (O_128,N_23292,N_24623);
and UO_129 (O_129,N_22923,N_24761);
nor UO_130 (O_130,N_24460,N_23752);
or UO_131 (O_131,N_24450,N_22982);
nor UO_132 (O_132,N_23182,N_23923);
xor UO_133 (O_133,N_24755,N_23103);
nand UO_134 (O_134,N_23598,N_22617);
or UO_135 (O_135,N_23585,N_23101);
nand UO_136 (O_136,N_22651,N_23921);
nand UO_137 (O_137,N_23978,N_24408);
nand UO_138 (O_138,N_23379,N_23107);
or UO_139 (O_139,N_24684,N_23130);
nand UO_140 (O_140,N_22634,N_24777);
and UO_141 (O_141,N_22829,N_24058);
nor UO_142 (O_142,N_23165,N_23248);
or UO_143 (O_143,N_23770,N_22812);
nand UO_144 (O_144,N_24493,N_22716);
or UO_145 (O_145,N_24671,N_22848);
or UO_146 (O_146,N_24419,N_24251);
and UO_147 (O_147,N_23026,N_24625);
and UO_148 (O_148,N_23447,N_22534);
nor UO_149 (O_149,N_23854,N_23412);
xnor UO_150 (O_150,N_23509,N_23065);
and UO_151 (O_151,N_24300,N_23224);
nor UO_152 (O_152,N_24271,N_24659);
or UO_153 (O_153,N_24152,N_24701);
or UO_154 (O_154,N_23880,N_22586);
or UO_155 (O_155,N_22735,N_22804);
nor UO_156 (O_156,N_24418,N_24919);
nand UO_157 (O_157,N_23554,N_23783);
or UO_158 (O_158,N_23762,N_22518);
nand UO_159 (O_159,N_22648,N_22861);
nor UO_160 (O_160,N_24395,N_23309);
and UO_161 (O_161,N_24270,N_24323);
nor UO_162 (O_162,N_23111,N_23188);
nand UO_163 (O_163,N_24954,N_23721);
xor UO_164 (O_164,N_24752,N_23950);
or UO_165 (O_165,N_22678,N_22615);
and UO_166 (O_166,N_22522,N_24506);
and UO_167 (O_167,N_23626,N_23213);
or UO_168 (O_168,N_22912,N_23258);
or UO_169 (O_169,N_24107,N_24999);
or UO_170 (O_170,N_23703,N_24038);
nand UO_171 (O_171,N_23300,N_24841);
and UO_172 (O_172,N_23190,N_23392);
and UO_173 (O_173,N_24407,N_23465);
or UO_174 (O_174,N_23041,N_22702);
and UO_175 (O_175,N_22922,N_23858);
nand UO_176 (O_176,N_22509,N_24547);
and UO_177 (O_177,N_23144,N_22915);
xnor UO_178 (O_178,N_24598,N_23704);
nor UO_179 (O_179,N_22537,N_23380);
xor UO_180 (O_180,N_24715,N_23679);
nor UO_181 (O_181,N_24133,N_24379);
and UO_182 (O_182,N_24920,N_23466);
and UO_183 (O_183,N_23485,N_22553);
and UO_184 (O_184,N_24094,N_23012);
nand UO_185 (O_185,N_24712,N_22714);
nand UO_186 (O_186,N_23967,N_24141);
nand UO_187 (O_187,N_23049,N_24066);
nand UO_188 (O_188,N_24655,N_24627);
nor UO_189 (O_189,N_23676,N_23244);
nor UO_190 (O_190,N_24022,N_24263);
or UO_191 (O_191,N_24523,N_24750);
or UO_192 (O_192,N_23387,N_23771);
or UO_193 (O_193,N_24298,N_24204);
nand UO_194 (O_194,N_24593,N_24723);
nand UO_195 (O_195,N_24322,N_23463);
nor UO_196 (O_196,N_24579,N_23918);
and UO_197 (O_197,N_24172,N_24336);
and UO_198 (O_198,N_23446,N_24800);
and UO_199 (O_199,N_24480,N_22930);
nor UO_200 (O_200,N_24394,N_23009);
nand UO_201 (O_201,N_23707,N_24157);
xnor UO_202 (O_202,N_22776,N_22517);
and UO_203 (O_203,N_23099,N_22622);
or UO_204 (O_204,N_24902,N_24691);
xor UO_205 (O_205,N_24195,N_24550);
or UO_206 (O_206,N_22701,N_24423);
nand UO_207 (O_207,N_23110,N_23373);
nand UO_208 (O_208,N_22803,N_24003);
or UO_209 (O_209,N_24612,N_24185);
xnor UO_210 (O_210,N_24159,N_23472);
or UO_211 (O_211,N_24737,N_24526);
nand UO_212 (O_212,N_24179,N_22569);
nor UO_213 (O_213,N_23448,N_24587);
xor UO_214 (O_214,N_23451,N_24102);
nor UO_215 (O_215,N_24237,N_23652);
or UO_216 (O_216,N_23277,N_23743);
and UO_217 (O_217,N_23489,N_23050);
or UO_218 (O_218,N_24861,N_22665);
nand UO_219 (O_219,N_24437,N_23597);
nand UO_220 (O_220,N_22512,N_23075);
nor UO_221 (O_221,N_24417,N_23734);
nor UO_222 (O_222,N_23434,N_24472);
nor UO_223 (O_223,N_23863,N_24769);
and UO_224 (O_224,N_23865,N_23281);
nand UO_225 (O_225,N_22624,N_23869);
nor UO_226 (O_226,N_23374,N_23174);
or UO_227 (O_227,N_22609,N_23199);
nor UO_228 (O_228,N_23272,N_24667);
and UO_229 (O_229,N_24846,N_23377);
or UO_230 (O_230,N_22956,N_24161);
nor UO_231 (O_231,N_24220,N_24075);
or UO_232 (O_232,N_23279,N_22690);
and UO_233 (O_233,N_23772,N_24609);
nand UO_234 (O_234,N_24981,N_22613);
nor UO_235 (O_235,N_22885,N_24438);
or UO_236 (O_236,N_23084,N_23305);
nor UO_237 (O_237,N_22592,N_23019);
nor UO_238 (O_238,N_23068,N_23403);
or UO_239 (O_239,N_23563,N_24785);
xnor UO_240 (O_240,N_24462,N_22984);
xnor UO_241 (O_241,N_22807,N_23359);
xor UO_242 (O_242,N_23264,N_24441);
nand UO_243 (O_243,N_23699,N_23579);
and UO_244 (O_244,N_23587,N_24310);
nand UO_245 (O_245,N_24930,N_23715);
nand UO_246 (O_246,N_22907,N_22641);
nand UO_247 (O_247,N_24706,N_24839);
and UO_248 (O_248,N_22528,N_24897);
nand UO_249 (O_249,N_23236,N_23583);
and UO_250 (O_250,N_22706,N_24398);
and UO_251 (O_251,N_22836,N_22647);
or UO_252 (O_252,N_23547,N_23847);
or UO_253 (O_253,N_23469,N_24576);
and UO_254 (O_254,N_22538,N_24643);
nor UO_255 (O_255,N_23666,N_22870);
nor UO_256 (O_256,N_22682,N_23189);
nand UO_257 (O_257,N_23449,N_23665);
or UO_258 (O_258,N_22521,N_24901);
nor UO_259 (O_259,N_23201,N_24651);
and UO_260 (O_260,N_24085,N_23611);
nand UO_261 (O_261,N_23813,N_24685);
nor UO_262 (O_262,N_23713,N_24586);
nand UO_263 (O_263,N_23298,N_23314);
and UO_264 (O_264,N_23149,N_22800);
nand UO_265 (O_265,N_22811,N_23572);
nor UO_266 (O_266,N_23404,N_24467);
nand UO_267 (O_267,N_22604,N_22591);
nand UO_268 (O_268,N_24248,N_22573);
nor UO_269 (O_269,N_22572,N_24832);
nor UO_270 (O_270,N_22936,N_23681);
or UO_271 (O_271,N_23871,N_24640);
nand UO_272 (O_272,N_24070,N_23114);
xnor UO_273 (O_273,N_23389,N_24260);
nor UO_274 (O_274,N_23230,N_23557);
nor UO_275 (O_275,N_24489,N_23822);
nand UO_276 (O_276,N_22627,N_24446);
and UO_277 (O_277,N_23100,N_24622);
xnor UO_278 (O_278,N_22681,N_24582);
and UO_279 (O_279,N_23018,N_24144);
nand UO_280 (O_280,N_23422,N_23649);
or UO_281 (O_281,N_23947,N_24492);
or UO_282 (O_282,N_24033,N_23438);
or UO_283 (O_283,N_22988,N_24540);
nor UO_284 (O_284,N_23663,N_24223);
nor UO_285 (O_285,N_24181,N_23537);
and UO_286 (O_286,N_22532,N_24117);
or UO_287 (O_287,N_24428,N_24637);
nand UO_288 (O_288,N_22744,N_23535);
nand UO_289 (O_289,N_23486,N_23409);
and UO_290 (O_290,N_23214,N_23883);
nand UO_291 (O_291,N_24632,N_23307);
nand UO_292 (O_292,N_23067,N_24308);
xor UO_293 (O_293,N_22595,N_23617);
nand UO_294 (O_294,N_24577,N_24439);
or UO_295 (O_295,N_24936,N_24032);
nand UO_296 (O_296,N_23891,N_24218);
and UO_297 (O_297,N_23949,N_24528);
nor UO_298 (O_298,N_23417,N_24042);
and UO_299 (O_299,N_23994,N_24468);
or UO_300 (O_300,N_24374,N_23294);
nor UO_301 (O_301,N_23886,N_24993);
nand UO_302 (O_302,N_24324,N_24926);
nand UO_303 (O_303,N_23082,N_24060);
nand UO_304 (O_304,N_24872,N_22659);
and UO_305 (O_305,N_23837,N_24483);
nand UO_306 (O_306,N_24660,N_22598);
or UO_307 (O_307,N_22637,N_23290);
nor UO_308 (O_308,N_24396,N_23618);
or UO_309 (O_309,N_23556,N_23150);
and UO_310 (O_310,N_24533,N_24436);
and UO_311 (O_311,N_23982,N_22882);
nand UO_312 (O_312,N_24206,N_23239);
or UO_313 (O_313,N_24069,N_24884);
and UO_314 (O_314,N_24699,N_23368);
or UO_315 (O_315,N_24754,N_24084);
nand UO_316 (O_316,N_22916,N_23879);
and UO_317 (O_317,N_24807,N_24120);
and UO_318 (O_318,N_23013,N_22931);
nor UO_319 (O_319,N_23348,N_24073);
nor UO_320 (O_320,N_22683,N_22772);
and UO_321 (O_321,N_23476,N_23811);
and UO_322 (O_322,N_23362,N_23695);
nand UO_323 (O_323,N_22889,N_24000);
xor UO_324 (O_324,N_22838,N_23548);
nor UO_325 (O_325,N_22942,N_24293);
or UO_326 (O_326,N_24539,N_24015);
nor UO_327 (O_327,N_23104,N_24282);
and UO_328 (O_328,N_24453,N_24690);
nand UO_329 (O_329,N_23097,N_22743);
or UO_330 (O_330,N_23612,N_22710);
and UO_331 (O_331,N_24555,N_24175);
nand UO_332 (O_332,N_24628,N_24478);
and UO_333 (O_333,N_24186,N_23673);
or UO_334 (O_334,N_22635,N_22783);
xor UO_335 (O_335,N_23976,N_23004);
nand UO_336 (O_336,N_22700,N_22904);
or UO_337 (O_337,N_24697,N_24442);
xnor UO_338 (O_338,N_24205,N_24071);
or UO_339 (O_339,N_24514,N_23116);
nand UO_340 (O_340,N_23893,N_24384);
nand UO_341 (O_341,N_24565,N_24944);
or UO_342 (O_342,N_23810,N_24142);
and UO_343 (O_343,N_23220,N_24648);
or UO_344 (O_344,N_24938,N_24290);
nor UO_345 (O_345,N_23705,N_23790);
xnor UO_346 (O_346,N_24330,N_23339);
or UO_347 (O_347,N_24334,N_24512);
nor UO_348 (O_348,N_23866,N_22654);
nor UO_349 (O_349,N_24975,N_23786);
and UO_350 (O_350,N_23087,N_22625);
nor UO_351 (O_351,N_22869,N_23776);
and UO_352 (O_352,N_22919,N_24791);
nand UO_353 (O_353,N_23946,N_23133);
or UO_354 (O_354,N_23045,N_23850);
or UO_355 (O_355,N_24292,N_23030);
xor UO_356 (O_356,N_24968,N_23956);
nor UO_357 (O_357,N_24414,N_23186);
nor UO_358 (O_358,N_23855,N_22839);
nand UO_359 (O_359,N_23320,N_24744);
or UO_360 (O_360,N_23607,N_23113);
and UO_361 (O_361,N_24782,N_24849);
xnor UO_362 (O_362,N_24736,N_24564);
nor UO_363 (O_363,N_23531,N_24964);
and UO_364 (O_364,N_23411,N_24111);
or UO_365 (O_365,N_24812,N_24448);
nor UO_366 (O_366,N_24339,N_24786);
nor UO_367 (O_367,N_23086,N_23512);
nand UO_368 (O_368,N_24105,N_24128);
nor UO_369 (O_369,N_23720,N_23669);
xor UO_370 (O_370,N_23260,N_22556);
nor UO_371 (O_371,N_24174,N_24366);
nor UO_372 (O_372,N_22691,N_23071);
nor UO_373 (O_373,N_22696,N_24966);
xor UO_374 (O_374,N_23491,N_23608);
and UO_375 (O_375,N_23957,N_23526);
nand UO_376 (O_376,N_22983,N_23902);
xnor UO_377 (O_377,N_22824,N_22834);
nor UO_378 (O_378,N_24789,N_23739);
nand UO_379 (O_379,N_22842,N_23211);
nor UO_380 (O_380,N_24262,N_24278);
nor UO_381 (O_381,N_23478,N_23749);
nor UO_382 (O_382,N_23054,N_23347);
nand UO_383 (O_383,N_22536,N_23126);
and UO_384 (O_384,N_24927,N_24048);
or UO_385 (O_385,N_24915,N_22819);
nand UO_386 (O_386,N_23252,N_22796);
xor UO_387 (O_387,N_23798,N_23061);
nor UO_388 (O_388,N_22763,N_24566);
nor UO_389 (O_389,N_24718,N_22937);
nor UO_390 (O_390,N_23742,N_23341);
or UO_391 (O_391,N_24674,N_24642);
or UO_392 (O_392,N_24455,N_24479);
nand UO_393 (O_393,N_24621,N_22841);
xor UO_394 (O_394,N_23151,N_22559);
or UO_395 (O_395,N_23995,N_23170);
or UO_396 (O_396,N_23361,N_24234);
nor UO_397 (O_397,N_24299,N_24020);
nor UO_398 (O_398,N_24843,N_24803);
nor UO_399 (O_399,N_23253,N_24004);
or UO_400 (O_400,N_24921,N_23899);
nor UO_401 (O_401,N_23621,N_22809);
nand UO_402 (O_402,N_22577,N_22901);
and UO_403 (O_403,N_24881,N_24104);
or UO_404 (O_404,N_23736,N_24026);
and UO_405 (O_405,N_23005,N_24680);
and UO_406 (O_406,N_22697,N_23637);
or UO_407 (O_407,N_23800,N_23105);
and UO_408 (O_408,N_24072,N_24343);
xor UO_409 (O_409,N_22971,N_24201);
and UO_410 (O_410,N_22511,N_23455);
and UO_411 (O_411,N_23539,N_24720);
xnor UO_412 (O_412,N_23746,N_22719);
nand UO_413 (O_413,N_24911,N_24558);
xor UO_414 (O_414,N_23198,N_23674);
nor UO_415 (O_415,N_23276,N_23250);
xor UO_416 (O_416,N_22843,N_24389);
nor UO_417 (O_417,N_22717,N_24580);
xnor UO_418 (O_418,N_24376,N_24127);
nand UO_419 (O_419,N_22727,N_23913);
nand UO_420 (O_420,N_22680,N_23933);
and UO_421 (O_421,N_23826,N_22610);
nand UO_422 (O_422,N_22721,N_23915);
and UO_423 (O_423,N_23021,N_22980);
and UO_424 (O_424,N_22945,N_23059);
or UO_425 (O_425,N_22759,N_24108);
or UO_426 (O_426,N_24698,N_23815);
nor UO_427 (O_427,N_24130,N_23834);
nand UO_428 (O_428,N_23055,N_22630);
nor UO_429 (O_429,N_23565,N_23983);
xnor UO_430 (O_430,N_22867,N_22601);
or UO_431 (O_431,N_23330,N_24112);
nand UO_432 (O_432,N_23575,N_23639);
nand UO_433 (O_433,N_23971,N_24212);
nand UO_434 (O_434,N_23935,N_24273);
nor UO_435 (O_435,N_24245,N_23473);
nor UO_436 (O_436,N_22636,N_24601);
nor UO_437 (O_437,N_24272,N_24854);
and UO_438 (O_438,N_23496,N_24912);
and UO_439 (O_439,N_22758,N_22606);
nor UO_440 (O_440,N_24959,N_24035);
or UO_441 (O_441,N_22600,N_24742);
nand UO_442 (O_442,N_23508,N_23955);
xor UO_443 (O_443,N_23938,N_23355);
and UO_444 (O_444,N_24028,N_24501);
or UO_445 (O_445,N_22769,N_24093);
nand UO_446 (O_446,N_22698,N_24385);
or UO_447 (O_447,N_23223,N_24076);
nor UO_448 (O_448,N_24947,N_23079);
nand UO_449 (O_449,N_23140,N_22799);
and UO_450 (O_450,N_23313,N_22862);
nand UO_451 (O_451,N_22884,N_23143);
and UO_452 (O_452,N_23162,N_23391);
nand UO_453 (O_453,N_24544,N_24899);
and UO_454 (O_454,N_24177,N_22611);
and UO_455 (O_455,N_23842,N_24188);
nor UO_456 (O_456,N_22539,N_24748);
xor UO_457 (O_457,N_23037,N_22516);
nand UO_458 (O_458,N_23881,N_22519);
xnor UO_459 (O_459,N_23874,N_24426);
nand UO_460 (O_460,N_24099,N_23468);
nand UO_461 (O_461,N_22508,N_22728);
xnor UO_462 (O_462,N_23261,N_24511);
nor UO_463 (O_463,N_23523,N_23977);
or UO_464 (O_464,N_24956,N_22883);
nor UO_465 (O_465,N_23846,N_23954);
and UO_466 (O_466,N_23419,N_23809);
and UO_467 (O_467,N_22818,N_24729);
or UO_468 (O_468,N_22798,N_23932);
or UO_469 (O_469,N_22531,N_22813);
nand UO_470 (O_470,N_24316,N_22954);
nand UO_471 (O_471,N_24406,N_24976);
xor UO_472 (O_472,N_22955,N_24734);
and UO_473 (O_473,N_24646,N_22541);
nand UO_474 (O_474,N_24067,N_24708);
and UO_475 (O_475,N_23332,N_24430);
nand UO_476 (O_476,N_23769,N_23929);
nand UO_477 (O_477,N_24688,N_24347);
or UO_478 (O_478,N_23283,N_24165);
nor UO_479 (O_479,N_22745,N_22677);
or UO_480 (O_480,N_23504,N_23925);
nand UO_481 (O_481,N_23641,N_23525);
nand UO_482 (O_482,N_23553,N_22941);
xor UO_483 (O_483,N_23780,N_23787);
nor UO_484 (O_484,N_23441,N_24192);
xor UO_485 (O_485,N_23247,N_23788);
nand UO_486 (O_486,N_24707,N_24764);
xnor UO_487 (O_487,N_22981,N_23958);
and UO_488 (O_488,N_24765,N_22913);
and UO_489 (O_489,N_23179,N_22639);
or UO_490 (O_490,N_24217,N_22726);
nand UO_491 (O_491,N_23218,N_22924);
xnor UO_492 (O_492,N_24477,N_24840);
nor UO_493 (O_493,N_24129,N_23217);
or UO_494 (O_494,N_23824,N_24862);
nor UO_495 (O_495,N_22756,N_24634);
nor UO_496 (O_496,N_22557,N_24645);
or UO_497 (O_497,N_23725,N_22855);
nand UO_498 (O_498,N_23999,N_23969);
or UO_499 (O_499,N_24435,N_23584);
nor UO_500 (O_500,N_24524,N_23440);
nor UO_501 (O_501,N_24424,N_23057);
nor UO_502 (O_502,N_24180,N_24132);
nand UO_503 (O_503,N_23315,N_23234);
and UO_504 (O_504,N_24447,N_24746);
nor UO_505 (O_505,N_24007,N_24986);
and UO_506 (O_506,N_23108,N_22655);
and UO_507 (O_507,N_23694,N_24355);
and UO_508 (O_508,N_24340,N_24694);
or UO_509 (O_509,N_22652,N_23848);
nand UO_510 (O_510,N_23000,N_24767);
nand UO_511 (O_511,N_22755,N_24052);
and UO_512 (O_512,N_24416,N_23413);
or UO_513 (O_513,N_23890,N_23338);
or UO_514 (O_514,N_22817,N_22524);
nor UO_515 (O_515,N_24471,N_23593);
nand UO_516 (O_516,N_22777,N_23708);
nand UO_517 (O_517,N_23516,N_22679);
nor UO_518 (O_518,N_23832,N_22925);
and UO_519 (O_519,N_23632,N_24778);
and UO_520 (O_520,N_23077,N_24505);
or UO_521 (O_521,N_24258,N_22778);
or UO_522 (O_522,N_24575,N_24863);
nor UO_523 (O_523,N_24738,N_24871);
or UO_524 (O_524,N_24836,N_23329);
and UO_525 (O_525,N_24768,N_24924);
nand UO_526 (O_526,N_24012,N_24082);
xnor UO_527 (O_527,N_24530,N_23601);
nand UO_528 (O_528,N_24103,N_24545);
nand UO_529 (O_529,N_23069,N_23155);
and UO_530 (O_530,N_23318,N_22962);
or UO_531 (O_531,N_23360,N_22952);
and UO_532 (O_532,N_24275,N_24429);
or UO_533 (O_533,N_23095,N_23603);
or UO_534 (O_534,N_23936,N_23129);
xnor UO_535 (O_535,N_23636,N_22943);
or UO_536 (O_536,N_24412,N_24124);
nor UO_537 (O_537,N_23613,N_23635);
xor UO_538 (O_538,N_24852,N_23737);
nand UO_539 (O_539,N_22897,N_23830);
nor UO_540 (O_540,N_22657,N_23945);
and UO_541 (O_541,N_24486,N_23275);
nand UO_542 (O_542,N_23255,N_24280);
or UO_543 (O_543,N_22668,N_22899);
and UO_544 (O_544,N_22566,N_23561);
nor UO_545 (O_545,N_23123,N_24572);
or UO_546 (O_546,N_23405,N_24303);
nand UO_547 (O_547,N_23467,N_22623);
or UO_548 (O_548,N_24745,N_24139);
and UO_549 (O_549,N_24341,N_22785);
and UO_550 (O_550,N_24315,N_24513);
nand UO_551 (O_551,N_23128,N_23212);
and UO_552 (O_552,N_24989,N_24225);
nor UO_553 (O_553,N_23402,N_22725);
nand UO_554 (O_554,N_22547,N_24624);
and UO_555 (O_555,N_23505,N_22621);
xor UO_556 (O_556,N_24371,N_23432);
and UO_557 (O_557,N_22852,N_23852);
or UO_558 (O_558,N_24827,N_23288);
xnor UO_559 (O_559,N_23371,N_22709);
or UO_560 (O_560,N_23345,N_24503);
nand UO_561 (O_561,N_22514,N_22736);
nor UO_562 (O_562,N_23817,N_24835);
or UO_563 (O_563,N_22933,N_23278);
nor UO_564 (O_564,N_23238,N_22911);
nand UO_565 (O_565,N_22791,N_24616);
or UO_566 (O_566,N_24906,N_24907);
nor UO_567 (O_567,N_23763,N_22540);
nor UO_568 (O_568,N_24844,N_22675);
xnor UO_569 (O_569,N_23142,N_24978);
xnor UO_570 (O_570,N_23841,N_24681);
nand UO_571 (O_571,N_23483,N_23624);
or UO_572 (O_572,N_24226,N_24943);
or UO_573 (O_573,N_23488,N_24291);
nand UO_574 (O_574,N_24928,N_24726);
nor UO_575 (O_575,N_24279,N_23462);
or UO_576 (O_576,N_24044,N_23643);
and UO_577 (O_577,N_24259,N_23375);
xor UO_578 (O_578,N_24638,N_23316);
and UO_579 (O_579,N_23202,N_24965);
and UO_580 (O_580,N_23425,N_22552);
nand UO_581 (O_581,N_24254,N_23381);
or UO_582 (O_582,N_24798,N_24535);
nor UO_583 (O_583,N_22996,N_23986);
and UO_584 (O_584,N_22578,N_24097);
or UO_585 (O_585,N_23167,N_22854);
nor UO_586 (O_586,N_24420,N_24224);
xnor UO_587 (O_587,N_24228,N_23744);
nand UO_588 (O_588,N_22991,N_24713);
and UO_589 (O_589,N_22917,N_24805);
or UO_590 (O_590,N_24122,N_24367);
nor UO_591 (O_591,N_22944,N_24463);
and UO_592 (O_592,N_24641,N_24864);
and UO_593 (O_593,N_24404,N_22774);
xnor UO_594 (O_594,N_23197,N_24647);
nand UO_595 (O_595,N_23840,N_23040);
and UO_596 (O_596,N_23610,N_22906);
and UO_597 (O_597,N_24534,N_23552);
xor UO_598 (O_598,N_24168,N_24942);
nor UO_599 (O_599,N_23653,N_23555);
xnor UO_600 (O_600,N_23916,N_23843);
xor UO_601 (O_601,N_24047,N_23456);
and UO_602 (O_602,N_22840,N_24305);
xnor UO_603 (O_603,N_24538,N_24295);
or UO_604 (O_604,N_24549,N_24383);
nand UO_605 (O_605,N_24173,N_23697);
and UO_606 (O_606,N_23718,N_23536);
and UO_607 (O_607,N_23171,N_23014);
nand UO_608 (O_608,N_24190,N_23401);
or UO_609 (O_609,N_24083,N_22545);
nand UO_610 (O_610,N_23633,N_23060);
or UO_611 (O_611,N_22502,N_23867);
and UO_612 (O_612,N_24876,N_23538);
and UO_613 (O_613,N_24977,N_23908);
and UO_614 (O_614,N_22530,N_24431);
and UO_615 (O_615,N_24830,N_23117);
or UO_616 (O_616,N_22584,N_24693);
or UO_617 (O_617,N_23388,N_23693);
nand UO_618 (O_618,N_24079,N_24845);
nand UO_619 (O_619,N_22589,N_24584);
and UO_620 (O_620,N_23291,N_24222);
and UO_621 (O_621,N_24650,N_24005);
xor UO_622 (O_622,N_23589,N_24630);
or UO_623 (O_623,N_24363,N_24866);
nand UO_624 (O_624,N_23042,N_23344);
nor UO_625 (O_625,N_24283,N_23029);
xor UO_626 (O_626,N_23773,N_24247);
and UO_627 (O_627,N_23941,N_24166);
and UO_628 (O_628,N_23828,N_22830);
xor UO_629 (O_629,N_22575,N_22767);
or UO_630 (O_630,N_24909,N_24838);
nand UO_631 (O_631,N_23231,N_23524);
and UO_632 (O_632,N_24617,N_24856);
and UO_633 (O_633,N_23581,N_24686);
and UO_634 (O_634,N_22821,N_23033);
nand UO_635 (O_635,N_23559,N_23470);
xnor UO_636 (O_636,N_22571,N_23654);
nand UO_637 (O_637,N_23263,N_24352);
or UO_638 (O_638,N_22815,N_23363);
or UO_639 (O_639,N_23926,N_24940);
nor UO_640 (O_640,N_22934,N_23173);
and UO_641 (O_641,N_22663,N_24703);
nand UO_642 (O_642,N_22999,N_24034);
or UO_643 (O_643,N_23839,N_22686);
and UO_644 (O_644,N_22849,N_23530);
nor UO_645 (O_645,N_23661,N_23606);
and UO_646 (O_646,N_24126,N_22977);
or UO_647 (O_647,N_23135,N_23775);
and UO_648 (O_648,N_23542,N_24747);
and UO_649 (O_649,N_24877,N_24518);
or UO_650 (O_650,N_24045,N_23779);
nor UO_651 (O_651,N_23048,N_24644);
and UO_652 (O_652,N_23758,N_24772);
xor UO_653 (O_653,N_24988,N_24665);
and UO_654 (O_654,N_24196,N_22888);
nor UO_655 (O_655,N_23930,N_23349);
and UO_656 (O_656,N_23730,N_24265);
or UO_657 (O_657,N_24057,N_22868);
and UO_658 (O_658,N_23043,N_23051);
nor UO_659 (O_659,N_23934,N_22833);
and UO_660 (O_660,N_24221,N_24904);
and UO_661 (O_661,N_22733,N_23667);
xor UO_662 (O_662,N_24449,N_22857);
nand UO_663 (O_663,N_23437,N_23265);
and UO_664 (O_664,N_24882,N_23896);
nand UO_665 (O_665,N_22560,N_22935);
and UO_666 (O_666,N_24203,N_22632);
and UO_667 (O_667,N_23353,N_22580);
xor UO_668 (O_668,N_23656,N_23541);
or UO_669 (O_669,N_24743,N_24850);
and UO_670 (O_670,N_23709,N_23216);
nand UO_671 (O_671,N_23124,N_23658);
and UO_672 (O_672,N_24678,N_24202);
or UO_673 (O_673,N_23158,N_23517);
nor UO_674 (O_674,N_24319,N_23429);
and UO_675 (O_675,N_23882,N_22948);
or UO_676 (O_676,N_22705,N_22581);
nor UO_677 (O_677,N_24123,N_24194);
or UO_678 (O_678,N_23146,N_22895);
nor UO_679 (O_679,N_23651,N_24121);
nor UO_680 (O_680,N_24529,N_24148);
or UO_681 (O_681,N_23684,N_23529);
or UO_682 (O_682,N_22975,N_24657);
nand UO_683 (O_683,N_24326,N_23549);
xnor UO_684 (O_684,N_22554,N_23148);
nand UO_685 (O_685,N_24284,N_24984);
or UO_686 (O_686,N_24023,N_24740);
and UO_687 (O_687,N_24962,N_24377);
nor UO_688 (O_688,N_24207,N_24795);
and UO_689 (O_689,N_24297,N_22708);
nor UO_690 (O_690,N_23141,N_23992);
and UO_691 (O_691,N_22832,N_23088);
and UO_692 (O_692,N_22520,N_23227);
and UO_693 (O_693,N_24808,N_23972);
xor UO_694 (O_694,N_24329,N_23326);
and UO_695 (O_695,N_22825,N_23225);
or UO_696 (O_696,N_22723,N_23164);
and UO_697 (O_697,N_24666,N_23596);
nor UO_698 (O_698,N_24613,N_23564);
nand UO_699 (O_699,N_23006,N_22501);
nand UO_700 (O_700,N_22871,N_24521);
and UO_701 (O_701,N_23112,N_23791);
nand UO_702 (O_702,N_23630,N_23889);
or UO_703 (O_703,N_24286,N_23089);
and UO_704 (O_704,N_24031,N_24002);
nand UO_705 (O_705,N_23418,N_22970);
nand UO_706 (O_706,N_22646,N_23333);
nand UO_707 (O_707,N_24608,N_24163);
xor UO_708 (O_708,N_23397,N_24088);
or UO_709 (O_709,N_24735,N_23671);
and UO_710 (O_710,N_24831,N_24553);
or UO_711 (O_711,N_22891,N_24910);
nor UO_712 (O_712,N_23970,N_22748);
nand UO_713 (O_713,N_23748,N_23735);
or UO_714 (O_714,N_24961,N_23266);
nor UO_715 (O_715,N_22782,N_24589);
nor UO_716 (O_716,N_23711,N_24847);
nor UO_717 (O_717,N_23953,N_23493);
or UO_718 (O_718,N_24819,N_22692);
or UO_719 (O_719,N_22671,N_23700);
nor UO_720 (O_720,N_22764,N_23943);
nand UO_721 (O_721,N_22510,N_23299);
xor UO_722 (O_722,N_23723,N_24311);
or UO_723 (O_723,N_23445,N_22746);
and UO_724 (O_724,N_24728,N_24811);
nand UO_725 (O_725,N_24860,N_24368);
nor UO_726 (O_726,N_24392,N_22880);
nand UO_727 (O_727,N_24131,N_23778);
and UO_728 (O_728,N_23987,N_23519);
nand UO_729 (O_729,N_24953,N_22676);
and UO_730 (O_730,N_24214,N_24342);
and UO_731 (O_731,N_24089,N_23396);
or UO_732 (O_732,N_23351,N_24602);
nor UO_733 (O_733,N_24359,N_24238);
nand UO_734 (O_734,N_23370,N_23696);
and UO_735 (O_735,N_22794,N_23857);
or UO_736 (O_736,N_23160,N_22872);
or UO_737 (O_737,N_24495,N_24932);
nand UO_738 (O_738,N_23728,N_23761);
nor UO_739 (O_739,N_23939,N_23712);
and UO_740 (O_740,N_23183,N_23906);
nand UO_741 (O_741,N_23522,N_22568);
nand UO_742 (O_742,N_23756,N_22787);
nor UO_743 (O_743,N_23997,N_23688);
or UO_744 (O_744,N_23308,N_23844);
and UO_745 (O_745,N_24242,N_24309);
and UO_746 (O_746,N_24285,N_23682);
nor UO_747 (O_747,N_24520,N_23868);
and UO_748 (O_748,N_24317,N_22666);
and UO_749 (O_749,N_22846,N_22551);
nor UO_750 (O_750,N_23191,N_23692);
nor UO_751 (O_751,N_23640,N_22558);
or UO_752 (O_752,N_24879,N_24459);
nand UO_753 (O_753,N_24137,N_23237);
nor UO_754 (O_754,N_22865,N_23860);
xor UO_755 (O_755,N_24799,N_23789);
nand UO_756 (O_756,N_24607,N_24470);
and UO_757 (O_757,N_24682,N_24354);
and UO_758 (O_758,N_24146,N_23340);
nand UO_759 (O_759,N_22515,N_23439);
nand UO_760 (O_760,N_23495,N_23701);
or UO_761 (O_761,N_23808,N_24870);
xnor UO_762 (O_762,N_23499,N_24603);
or UO_763 (O_763,N_22669,N_23591);
nand UO_764 (O_764,N_22593,N_24357);
or UO_765 (O_765,N_24397,N_23966);
nand UO_766 (O_766,N_24092,N_24425);
and UO_767 (O_767,N_23685,N_23960);
xor UO_768 (O_768,N_23507,N_23586);
nand UO_769 (O_769,N_24760,N_22979);
nor UO_770 (O_770,N_23336,N_22585);
nor UO_771 (O_771,N_22703,N_24955);
nor UO_772 (O_772,N_23127,N_22890);
and UO_773 (O_773,N_23393,N_24444);
or UO_774 (O_774,N_24098,N_23793);
or UO_775 (O_775,N_24510,N_24219);
nor UO_776 (O_776,N_24268,N_24151);
or UO_777 (O_777,N_24276,N_24046);
xnor UO_778 (O_778,N_24243,N_23074);
nor UO_779 (O_779,N_23118,N_24779);
nand UO_780 (O_780,N_23001,N_22801);
nor UO_781 (O_781,N_23528,N_24578);
xnor UO_782 (O_782,N_22886,N_23196);
nand UO_783 (O_783,N_23193,N_22894);
nand UO_784 (O_784,N_23053,N_23628);
and UO_785 (O_785,N_23806,N_23614);
and UO_786 (O_786,N_24213,N_23350);
nand UO_787 (O_787,N_22814,N_23301);
and UO_788 (O_788,N_22989,N_23833);
nor UO_789 (O_789,N_22875,N_23092);
nand UO_790 (O_790,N_23383,N_23973);
and UO_791 (O_791,N_23861,N_24135);
and UO_792 (O_792,N_23136,N_23251);
or UO_793 (O_793,N_23153,N_23436);
nand UO_794 (O_794,N_22715,N_22685);
and UO_795 (O_795,N_22887,N_24014);
or UO_796 (O_796,N_24469,N_24974);
and UO_797 (O_797,N_22856,N_22729);
or UO_798 (O_798,N_22616,N_23942);
nor UO_799 (O_799,N_22739,N_23346);
nor UO_800 (O_800,N_22607,N_23269);
nand UO_801 (O_801,N_24086,N_23474);
and UO_802 (O_802,N_23335,N_23905);
xnor UO_803 (O_803,N_24869,N_24318);
and UO_804 (O_804,N_23271,N_22918);
and UO_805 (O_805,N_24669,N_23394);
or UO_806 (O_806,N_24183,N_24191);
nand UO_807 (O_807,N_22864,N_23677);
nor UO_808 (O_808,N_24801,N_23856);
nor UO_809 (O_809,N_23482,N_24762);
nor UO_810 (O_810,N_23070,N_23464);
nand UO_811 (O_811,N_22995,N_22754);
nor UO_812 (O_812,N_24721,N_23988);
nand UO_813 (O_813,N_23210,N_22969);
nand UO_814 (O_814,N_22978,N_23917);
nor UO_815 (O_815,N_22564,N_24496);
or UO_816 (O_816,N_23662,N_23543);
nand UO_817 (O_817,N_24658,N_24344);
and UO_818 (O_818,N_23072,N_22878);
xor UO_819 (O_819,N_22992,N_23660);
nor UO_820 (O_820,N_23125,N_22741);
and UO_821 (O_821,N_22784,N_22960);
nand UO_822 (O_822,N_24809,N_23132);
xor UO_823 (O_823,N_22753,N_23177);
and UO_824 (O_824,N_23256,N_24833);
nor UO_825 (O_825,N_23372,N_23063);
and UO_826 (O_826,N_22740,N_24971);
or UO_827 (O_827,N_23442,N_24150);
and UO_828 (O_828,N_23616,N_24451);
nor UO_829 (O_829,N_22790,N_24679);
and UO_830 (O_830,N_23638,N_24570);
xnor UO_831 (O_831,N_24364,N_23302);
and UO_832 (O_832,N_23376,N_23137);
nor UO_833 (O_833,N_24011,N_23727);
and UO_834 (O_834,N_23027,N_23267);
or UO_835 (O_835,N_22770,N_24776);
nor UO_836 (O_836,N_24552,N_22752);
nor UO_837 (O_837,N_22550,N_24948);
nand UO_838 (O_838,N_24147,N_24010);
and UO_839 (O_839,N_23998,N_24732);
and UO_840 (O_840,N_24256,N_22689);
nand UO_841 (O_841,N_24618,N_23475);
nand UO_842 (O_842,N_23080,N_23492);
or UO_843 (O_843,N_23802,N_23284);
and UO_844 (O_844,N_22602,N_24560);
and UO_845 (O_845,N_24312,N_24946);
and UO_846 (O_846,N_23015,N_23147);
and UO_847 (O_847,N_23979,N_23687);
nand UO_848 (O_848,N_22967,N_23544);
nand UO_849 (O_849,N_24257,N_24696);
xnor UO_850 (O_850,N_24443,N_24804);
and UO_851 (O_851,N_23968,N_23620);
and UO_852 (O_852,N_23678,N_23159);
or UO_853 (O_853,N_22898,N_24413);
xnor UO_854 (O_854,N_23506,N_24403);
or UO_855 (O_855,N_22747,N_24790);
nor UO_856 (O_856,N_24170,N_24895);
nor UO_857 (O_857,N_23805,N_24491);
and UO_858 (O_858,N_24464,N_22837);
xor UO_859 (O_859,N_22684,N_22661);
and UO_860 (O_860,N_24473,N_23245);
nor UO_861 (O_861,N_24381,N_24662);
and UO_862 (O_862,N_24162,N_23823);
or UO_863 (O_863,N_23532,N_22579);
nand UO_864 (O_864,N_23323,N_22844);
and UO_865 (O_865,N_23629,N_23683);
nor UO_866 (O_866,N_24574,N_23430);
and UO_867 (O_867,N_23864,N_23794);
and UO_868 (O_868,N_23719,N_23322);
or UO_869 (O_869,N_24822,N_24466);
or UO_870 (O_870,N_24925,N_24611);
or UO_871 (O_871,N_23497,N_22619);
nand UO_872 (O_872,N_24880,N_23831);
and UO_873 (O_873,N_23851,N_22588);
and UO_874 (O_874,N_24313,N_23642);
nor UO_875 (O_875,N_24215,N_24178);
and UO_876 (O_876,N_24333,N_22974);
nand UO_877 (O_877,N_23750,N_24253);
nor UO_878 (O_878,N_23884,N_24227);
nor UO_879 (O_879,N_23134,N_24176);
or UO_880 (O_880,N_23286,N_23427);
xor UO_881 (O_881,N_24041,N_22909);
nor UO_882 (O_882,N_22664,N_23753);
nand UO_883 (O_883,N_22722,N_24348);
or UO_884 (O_884,N_23003,N_23717);
nor UO_885 (O_885,N_24432,N_24017);
and UO_886 (O_886,N_23287,N_24821);
nand UO_887 (O_887,N_22695,N_23365);
or UO_888 (O_888,N_24653,N_24916);
nand UO_889 (O_889,N_23066,N_23582);
nand UO_890 (O_890,N_24113,N_22926);
and UO_891 (O_891,N_24614,N_23774);
and UO_892 (O_892,N_24751,N_23031);
or UO_893 (O_893,N_22614,N_24606);
and UO_894 (O_894,N_22788,N_23511);
nor UO_895 (O_895,N_24551,N_23948);
and UO_896 (O_896,N_24136,N_23514);
and UO_897 (O_897,N_23270,N_23740);
or UO_898 (O_898,N_23364,N_24784);
and UO_899 (O_899,N_24875,N_24700);
or UO_900 (O_900,N_24937,N_24825);
nor UO_901 (O_901,N_23343,N_22768);
nand UO_902 (O_902,N_23698,N_24676);
and UO_903 (O_903,N_23139,N_23036);
xnor UO_904 (O_904,N_24078,N_24683);
nand UO_905 (O_905,N_24516,N_23646);
or UO_906 (O_906,N_23249,N_22827);
and UO_907 (O_907,N_23578,N_23892);
and UO_908 (O_908,N_23039,N_24770);
nor UO_909 (O_909,N_24360,N_23044);
xnor UO_910 (O_910,N_24727,N_24345);
or UO_911 (O_911,N_23922,N_24619);
nor UO_912 (O_912,N_23337,N_24842);
and UO_913 (O_913,N_24036,N_24030);
or UO_914 (O_914,N_23398,N_23452);
nand UO_915 (O_915,N_24039,N_23501);
nand UO_916 (O_916,N_22946,N_23546);
nor UO_917 (O_917,N_22905,N_22645);
nand UO_918 (O_918,N_24816,N_22629);
nand UO_919 (O_919,N_23827,N_23984);
nand UO_920 (O_920,N_23091,N_22958);
nor UO_921 (O_921,N_24402,N_23604);
or UO_922 (O_922,N_24465,N_22874);
and UO_923 (O_923,N_24209,N_24507);
and UO_924 (O_924,N_24687,N_23959);
and UO_925 (O_925,N_24456,N_22640);
or UO_926 (O_926,N_23566,N_23751);
and UO_927 (O_927,N_24301,N_24813);
and UO_928 (O_928,N_23131,N_24605);
nand UO_929 (O_929,N_23952,N_22828);
or UO_930 (O_930,N_23550,N_23342);
and UO_931 (O_931,N_22628,N_24945);
nor UO_932 (O_932,N_23328,N_24664);
nand UO_933 (O_933,N_23035,N_23766);
nor UO_934 (O_934,N_23327,N_24979);
nand UO_935 (O_935,N_23759,N_24997);
xnor UO_936 (O_936,N_23215,N_24670);
and UO_937 (O_937,N_24411,N_23274);
nand UO_938 (O_938,N_24115,N_24952);
nor UO_939 (O_939,N_24110,N_23768);
nand UO_940 (O_940,N_24677,N_22724);
or UO_941 (O_941,N_23577,N_24663);
nor UO_942 (O_942,N_24970,N_23096);
nor UO_943 (O_943,N_23161,N_24169);
nand UO_944 (O_944,N_24457,N_23122);
xnor UO_945 (O_945,N_22544,N_22658);
nand UO_946 (O_946,N_22877,N_23317);
nor UO_947 (O_947,N_24563,N_22590);
or UO_948 (O_948,N_22587,N_23765);
nor UO_949 (O_949,N_23777,N_22693);
or UO_950 (O_950,N_23098,N_24461);
nand UO_951 (O_951,N_24753,N_24517);
nor UO_952 (O_952,N_22965,N_22908);
and UO_953 (O_953,N_22927,N_23166);
nand UO_954 (O_954,N_23928,N_24610);
and UO_955 (O_955,N_24888,N_24050);
or UO_956 (O_956,N_22562,N_22643);
xnor UO_957 (O_957,N_24458,N_23859);
or UO_958 (O_958,N_24021,N_23058);
nand UO_959 (O_959,N_24353,N_24399);
and UO_960 (O_960,N_24494,N_22976);
and UO_961 (O_961,N_23032,N_24725);
and UO_962 (O_962,N_24171,N_23580);
nor UO_963 (O_963,N_22858,N_24724);
or UO_964 (O_964,N_23453,N_23567);
or UO_965 (O_965,N_24763,N_24118);
and UO_966 (O_966,N_24421,N_23285);
and UO_967 (O_967,N_22845,N_24241);
xor UO_968 (O_968,N_23083,N_22576);
nand UO_969 (O_969,N_22549,N_22985);
nand UO_970 (O_970,N_23423,N_24826);
or UO_971 (O_971,N_23384,N_23240);
xor UO_972 (O_972,N_23209,N_23406);
nor UO_973 (O_973,N_24692,N_22525);
or UO_974 (O_974,N_24484,N_24983);
and UO_975 (O_975,N_24244,N_23232);
or UO_976 (O_976,N_23102,N_23878);
nand UO_977 (O_977,N_23119,N_23724);
and UO_978 (O_978,N_23904,N_24119);
nand UO_979 (O_979,N_23900,N_23024);
nand UO_980 (O_980,N_23870,N_24806);
nor UO_981 (O_981,N_22779,N_23156);
nor UO_982 (O_982,N_23121,N_23184);
nand UO_983 (O_983,N_23386,N_23458);
xnor UO_984 (O_984,N_23500,N_23257);
nor UO_985 (O_985,N_23690,N_24235);
nor UO_986 (O_986,N_23229,N_24985);
or UO_987 (O_987,N_23745,N_23259);
and UO_988 (O_988,N_23853,N_22694);
nand UO_989 (O_989,N_23784,N_23875);
nand UO_990 (O_990,N_22506,N_24599);
nand UO_991 (O_991,N_24400,N_24796);
and UO_992 (O_992,N_23560,N_23289);
or UO_993 (O_993,N_23145,N_23574);
nand UO_994 (O_994,N_23007,N_24705);
nor UO_995 (O_995,N_24973,N_23940);
and UO_996 (O_996,N_23176,N_24810);
or UO_997 (O_997,N_24739,N_24382);
nor UO_998 (O_998,N_24074,N_23481);
or UO_999 (O_999,N_23792,N_24499);
nand UO_1000 (O_1000,N_23818,N_23280);
and UO_1001 (O_1001,N_23028,N_22762);
nor UO_1002 (O_1002,N_24362,N_24527);
nor UO_1003 (O_1003,N_23814,N_24668);
nand UO_1004 (O_1004,N_24967,N_24568);
or UO_1005 (O_1005,N_22612,N_22563);
nand UO_1006 (O_1006,N_23471,N_24749);
or UO_1007 (O_1007,N_23602,N_23672);
and UO_1008 (O_1008,N_22704,N_23428);
nor UO_1009 (O_1009,N_22966,N_24261);
nand UO_1010 (O_1010,N_23600,N_23914);
xnor UO_1011 (O_1011,N_24991,N_24167);
or UO_1012 (O_1012,N_23664,N_24410);
and UO_1013 (O_1013,N_24903,N_23242);
nor UO_1014 (O_1014,N_24922,N_23568);
xnor UO_1015 (O_1015,N_24189,N_23981);
and UO_1016 (O_1016,N_24855,N_24635);
nand UO_1017 (O_1017,N_22792,N_24620);
xor UO_1018 (O_1018,N_23334,N_24274);
nor UO_1019 (O_1019,N_22620,N_23047);
nand UO_1020 (O_1020,N_22802,N_24350);
nor UO_1021 (O_1021,N_22750,N_23836);
nor UO_1022 (O_1022,N_22876,N_23927);
and UO_1023 (O_1023,N_24387,N_24325);
nor UO_1024 (O_1024,N_23716,N_24982);
nor UO_1025 (O_1025,N_23576,N_22903);
and UO_1026 (O_1026,N_23675,N_24255);
and UO_1027 (O_1027,N_22816,N_23273);
nand UO_1028 (O_1028,N_22605,N_24797);
xnor UO_1029 (O_1029,N_23754,N_24211);
or UO_1030 (O_1030,N_24365,N_24591);
or UO_1031 (O_1031,N_24328,N_24018);
and UO_1032 (O_1032,N_24388,N_23312);
or UO_1033 (O_1033,N_24592,N_23911);
nand UO_1034 (O_1034,N_23993,N_22597);
nor UO_1035 (O_1035,N_24583,N_23764);
nor UO_1036 (O_1036,N_24848,N_22957);
and UO_1037 (O_1037,N_24969,N_24008);
nor UO_1038 (O_1038,N_23235,N_22968);
or UO_1039 (O_1039,N_24025,N_24958);
and UO_1040 (O_1040,N_22932,N_23965);
or UO_1041 (O_1041,N_23573,N_23254);
nor UO_1042 (O_1042,N_24802,N_24109);
xor UO_1043 (O_1043,N_23845,N_24554);
or UO_1044 (O_1044,N_22940,N_24372);
and UO_1045 (O_1045,N_22561,N_24358);
or UO_1046 (O_1046,N_24476,N_23226);
nand UO_1047 (O_1047,N_24889,N_23185);
and UO_1048 (O_1048,N_24783,N_24095);
nand UO_1049 (O_1049,N_22734,N_24815);
nor UO_1050 (O_1050,N_22548,N_23168);
xor UO_1051 (O_1051,N_23599,N_24193);
nor UO_1052 (O_1052,N_22793,N_23459);
nor UO_1053 (O_1053,N_23686,N_23303);
xnor UO_1054 (O_1054,N_24629,N_23085);
and UO_1055 (O_1055,N_24541,N_23297);
and UO_1056 (O_1056,N_24061,N_22775);
and UO_1057 (O_1057,N_23352,N_23181);
or UO_1058 (O_1058,N_24184,N_24267);
and UO_1059 (O_1059,N_24894,N_24160);
xor UO_1060 (O_1060,N_23325,N_23194);
or UO_1061 (O_1061,N_24639,N_22805);
and UO_1062 (O_1062,N_23650,N_23989);
nand UO_1063 (O_1063,N_24853,N_22720);
and UO_1064 (O_1064,N_22835,N_24281);
nor UO_1065 (O_1065,N_23820,N_23484);
and UO_1066 (O_1066,N_24487,N_23400);
and UO_1067 (O_1067,N_23657,N_24380);
xor UO_1068 (O_1068,N_23937,N_23551);
or UO_1069 (O_1069,N_23435,N_22893);
and UO_1070 (O_1070,N_23319,N_24482);
nor UO_1071 (O_1071,N_22688,N_24327);
and UO_1072 (O_1072,N_24229,N_22881);
and UO_1073 (O_1073,N_23622,N_23631);
and UO_1074 (O_1074,N_24351,N_22773);
or UO_1075 (O_1075,N_24949,N_22730);
and UO_1076 (O_1076,N_23219,N_23592);
or UO_1077 (O_1077,N_24995,N_22503);
xor UO_1078 (O_1078,N_24296,N_24101);
or UO_1079 (O_1079,N_24332,N_22660);
nand UO_1080 (O_1080,N_24422,N_24980);
and UO_1081 (O_1081,N_23888,N_23849);
nor UO_1082 (O_1082,N_23444,N_23991);
or UO_1083 (O_1083,N_23246,N_23421);
and UO_1084 (O_1084,N_23207,N_24252);
nor UO_1085 (O_1085,N_24198,N_23747);
xor UO_1086 (O_1086,N_24818,N_24401);
and UO_1087 (O_1087,N_24154,N_22713);
xnor UO_1088 (O_1088,N_24873,N_23385);
xnor UO_1089 (O_1089,N_24346,N_23885);
nand UO_1090 (O_1090,N_22990,N_23659);
and UO_1091 (O_1091,N_23876,N_24053);
or UO_1092 (O_1092,N_24569,N_23295);
nor UO_1093 (O_1093,N_23887,N_24908);
nand UO_1094 (O_1094,N_22766,N_24604);
and UO_1095 (O_1095,N_23178,N_23895);
or UO_1096 (O_1096,N_22542,N_23595);
nand UO_1097 (O_1097,N_24731,N_24817);
nand UO_1098 (O_1098,N_22986,N_23964);
xnor UO_1099 (O_1099,N_23872,N_23461);
nor UO_1100 (O_1100,N_24633,N_24775);
nand UO_1101 (O_1101,N_23996,N_23152);
nand UO_1102 (O_1102,N_24780,N_22859);
nand UO_1103 (O_1103,N_23615,N_24415);
and UO_1104 (O_1104,N_24187,N_23625);
nor UO_1105 (O_1105,N_24636,N_24556);
nand UO_1106 (O_1106,N_23691,N_24781);
and UO_1107 (O_1107,N_24515,N_24631);
nand UO_1108 (O_1108,N_22543,N_24239);
nor UO_1109 (O_1109,N_22523,N_24730);
nor UO_1110 (O_1110,N_24998,N_24114);
or UO_1111 (O_1111,N_24386,N_22513);
nand UO_1112 (O_1112,N_24508,N_23494);
and UO_1113 (O_1113,N_23502,N_24059);
and UO_1114 (O_1114,N_23154,N_22810);
nor UO_1115 (O_1115,N_24878,N_24914);
nor UO_1116 (O_1116,N_22699,N_24649);
nor UO_1117 (O_1117,N_24950,N_22608);
and UO_1118 (O_1118,N_23903,N_22653);
xnor UO_1119 (O_1119,N_22667,N_23894);
or UO_1120 (O_1120,N_22853,N_23480);
xnor UO_1121 (O_1121,N_23017,N_22505);
or UO_1122 (O_1122,N_23807,N_24197);
nor UO_1123 (O_1123,N_23510,N_23424);
nor UO_1124 (O_1124,N_24029,N_24427);
or UO_1125 (O_1125,N_22795,N_23205);
and UO_1126 (O_1126,N_23907,N_22596);
and UO_1127 (O_1127,N_24559,N_24063);
or UO_1128 (O_1128,N_24304,N_24939);
nand UO_1129 (O_1129,N_23241,N_23090);
nand UO_1130 (O_1130,N_23797,N_24828);
nor UO_1131 (O_1131,N_24321,N_23757);
or UO_1132 (O_1132,N_24595,N_24758);
and UO_1133 (O_1133,N_23410,N_24957);
nand UO_1134 (O_1134,N_24935,N_22947);
and UO_1135 (O_1135,N_23187,N_22737);
and UO_1136 (O_1136,N_22599,N_23382);
and UO_1137 (O_1137,N_23898,N_22896);
and UO_1138 (O_1138,N_22851,N_23760);
and UO_1139 (O_1139,N_23395,N_23829);
nand UO_1140 (O_1140,N_22786,N_22504);
nand UO_1141 (O_1141,N_22638,N_22997);
or UO_1142 (O_1142,N_24001,N_24672);
or UO_1143 (O_1143,N_24481,N_23457);
xnor UO_1144 (O_1144,N_23433,N_24532);
and UO_1145 (O_1145,N_23605,N_24490);
or UO_1146 (O_1146,N_22939,N_24963);
nor UO_1147 (O_1147,N_22751,N_23781);
or UO_1148 (O_1148,N_24068,N_24370);
or UO_1149 (O_1149,N_24719,N_23974);
nand UO_1150 (O_1150,N_22662,N_24087);
nor UO_1151 (O_1151,N_23046,N_24557);
or UO_1152 (O_1152,N_23588,N_23729);
and UO_1153 (O_1153,N_22718,N_23655);
xor UO_1154 (O_1154,N_24857,N_23513);
nand UO_1155 (O_1155,N_24837,N_22765);
xor UO_1156 (O_1156,N_22823,N_23733);
nand UO_1157 (O_1157,N_24885,N_24917);
and UO_1158 (O_1158,N_24302,N_24972);
nand UO_1159 (O_1159,N_23268,N_23527);
or UO_1160 (O_1160,N_23157,N_24918);
xnor UO_1161 (O_1161,N_23460,N_23619);
xor UO_1162 (O_1162,N_24522,N_23540);
nor UO_1163 (O_1163,N_24519,N_24814);
nor UO_1164 (O_1164,N_22567,N_22987);
and UO_1165 (O_1165,N_23064,N_22928);
or UO_1166 (O_1166,N_24452,N_22574);
or UO_1167 (O_1167,N_22879,N_23825);
nor UO_1168 (O_1168,N_22565,N_22863);
and UO_1169 (O_1169,N_24867,N_23115);
nand UO_1170 (O_1170,N_22892,N_24892);
or UO_1171 (O_1171,N_24858,N_23454);
nor UO_1172 (O_1172,N_24216,N_22594);
or UO_1173 (O_1173,N_23357,N_24859);
or UO_1174 (O_1174,N_24335,N_24236);
or UO_1175 (O_1175,N_24891,N_22529);
nand UO_1176 (O_1176,N_22963,N_23293);
nand UO_1177 (O_1177,N_23648,N_22760);
or UO_1178 (O_1178,N_23078,N_23570);
or UO_1179 (O_1179,N_23924,N_24851);
and UO_1180 (O_1180,N_24488,N_24249);
xnor UO_1181 (O_1181,N_23008,N_22656);
and UO_1182 (O_1182,N_22910,N_24733);
nor UO_1183 (O_1183,N_24702,N_23262);
and UO_1184 (O_1184,N_23180,N_22959);
or UO_1185 (O_1185,N_24590,N_23702);
or UO_1186 (O_1186,N_24824,N_23093);
nand UO_1187 (O_1187,N_24987,N_24027);
nand UO_1188 (O_1188,N_24498,N_24024);
nand UO_1189 (O_1189,N_23680,N_24356);
and UO_1190 (O_1190,N_23358,N_24548);
nand UO_1191 (O_1191,N_22707,N_23931);
and UO_1192 (O_1192,N_24062,N_23782);
or UO_1193 (O_1193,N_22749,N_24941);
and UO_1194 (O_1194,N_24134,N_22582);
nand UO_1195 (O_1195,N_23722,N_24661);
nor UO_1196 (O_1196,N_23282,N_22533);
and UO_1197 (O_1197,N_22712,N_24307);
nor UO_1198 (O_1198,N_22527,N_22808);
nor UO_1199 (O_1199,N_23206,N_24077);
xor UO_1200 (O_1200,N_24717,N_22555);
xnor UO_1201 (O_1201,N_24766,N_22649);
or UO_1202 (O_1202,N_22998,N_24475);
nor UO_1203 (O_1203,N_23369,N_24695);
nor UO_1204 (O_1204,N_22583,N_24771);
xor UO_1205 (O_1205,N_24116,N_23222);
and UO_1206 (O_1206,N_23558,N_24834);
or UO_1207 (O_1207,N_23877,N_23208);
nor UO_1208 (O_1208,N_22626,N_24542);
and UO_1209 (O_1209,N_24277,N_22993);
or UO_1210 (O_1210,N_23450,N_22603);
xnor UO_1211 (O_1211,N_24440,N_23738);
and UO_1212 (O_1212,N_24232,N_23306);
nand UO_1213 (O_1213,N_23726,N_24573);
nor UO_1214 (O_1214,N_23354,N_22847);
nand UO_1215 (O_1215,N_24923,N_24704);
or UO_1216 (O_1216,N_24561,N_22953);
or UO_1217 (O_1217,N_23562,N_22780);
and UO_1218 (O_1218,N_24158,N_23038);
nor UO_1219 (O_1219,N_23873,N_24597);
xnor UO_1220 (O_1220,N_24741,N_23081);
nor UO_1221 (O_1221,N_24156,N_24369);
nor UO_1222 (O_1222,N_24829,N_23951);
nor UO_1223 (O_1223,N_23490,N_24314);
nor UO_1224 (O_1224,N_23109,N_22731);
and UO_1225 (O_1225,N_24405,N_22673);
or UO_1226 (O_1226,N_24714,N_24689);
nand UO_1227 (O_1227,N_24896,N_23195);
and UO_1228 (O_1228,N_23399,N_24289);
or UO_1229 (O_1229,N_23521,N_24054);
or UO_1230 (O_1230,N_24883,N_24096);
xor UO_1231 (O_1231,N_24016,N_22831);
and UO_1232 (O_1232,N_24090,N_24500);
or UO_1233 (O_1233,N_24040,N_24013);
nor UO_1234 (O_1234,N_23025,N_22687);
nand UO_1235 (O_1235,N_22633,N_23106);
and UO_1236 (O_1236,N_23801,N_24615);
xor UO_1237 (O_1237,N_24378,N_23647);
xnor UO_1238 (O_1238,N_24934,N_23897);
and UO_1239 (O_1239,N_23010,N_23020);
and UO_1240 (O_1240,N_24709,N_23408);
and UO_1241 (O_1241,N_23714,N_24337);
and UO_1242 (O_1242,N_22771,N_22711);
or UO_1243 (O_1243,N_24055,N_23443);
nor UO_1244 (O_1244,N_24929,N_24390);
nand UO_1245 (O_1245,N_23518,N_23175);
nor UO_1246 (O_1246,N_24373,N_22826);
or UO_1247 (O_1247,N_23571,N_24497);
nor UO_1248 (O_1248,N_23120,N_24064);
nand UO_1249 (O_1249,N_24009,N_24588);
nand UO_1250 (O_1250,N_23379,N_24409);
or UO_1251 (O_1251,N_24635,N_23211);
nor UO_1252 (O_1252,N_22657,N_23343);
xnor UO_1253 (O_1253,N_24399,N_23921);
nand UO_1254 (O_1254,N_23932,N_24740);
nor UO_1255 (O_1255,N_22926,N_24035);
and UO_1256 (O_1256,N_24919,N_24739);
nand UO_1257 (O_1257,N_22560,N_24396);
nor UO_1258 (O_1258,N_24741,N_23125);
or UO_1259 (O_1259,N_24539,N_23823);
nand UO_1260 (O_1260,N_24486,N_23502);
xor UO_1261 (O_1261,N_22770,N_22743);
and UO_1262 (O_1262,N_23018,N_23902);
and UO_1263 (O_1263,N_22791,N_24075);
nand UO_1264 (O_1264,N_24161,N_23574);
or UO_1265 (O_1265,N_24935,N_24585);
nand UO_1266 (O_1266,N_23728,N_23034);
and UO_1267 (O_1267,N_23616,N_24655);
xor UO_1268 (O_1268,N_24644,N_23232);
nand UO_1269 (O_1269,N_23960,N_23928);
nand UO_1270 (O_1270,N_23938,N_23842);
and UO_1271 (O_1271,N_23010,N_24546);
nor UO_1272 (O_1272,N_23057,N_24414);
and UO_1273 (O_1273,N_22766,N_23277);
xnor UO_1274 (O_1274,N_24296,N_23799);
nor UO_1275 (O_1275,N_22994,N_23860);
nand UO_1276 (O_1276,N_22911,N_24153);
nand UO_1277 (O_1277,N_23446,N_24758);
xnor UO_1278 (O_1278,N_24839,N_23972);
nor UO_1279 (O_1279,N_23961,N_24136);
or UO_1280 (O_1280,N_24254,N_22524);
nand UO_1281 (O_1281,N_23962,N_23057);
and UO_1282 (O_1282,N_24561,N_23671);
nor UO_1283 (O_1283,N_24367,N_24216);
or UO_1284 (O_1284,N_23461,N_23302);
nand UO_1285 (O_1285,N_22675,N_24419);
xnor UO_1286 (O_1286,N_24744,N_24798);
nand UO_1287 (O_1287,N_23214,N_23786);
nand UO_1288 (O_1288,N_23521,N_24563);
nor UO_1289 (O_1289,N_24519,N_24327);
nor UO_1290 (O_1290,N_22647,N_23801);
or UO_1291 (O_1291,N_24126,N_24697);
or UO_1292 (O_1292,N_24862,N_22883);
nor UO_1293 (O_1293,N_23000,N_23233);
nor UO_1294 (O_1294,N_23359,N_23947);
or UO_1295 (O_1295,N_23028,N_23824);
and UO_1296 (O_1296,N_22688,N_23039);
nand UO_1297 (O_1297,N_24153,N_24313);
or UO_1298 (O_1298,N_22603,N_24462);
nand UO_1299 (O_1299,N_24625,N_22585);
or UO_1300 (O_1300,N_24316,N_22717);
or UO_1301 (O_1301,N_23985,N_24645);
xor UO_1302 (O_1302,N_22567,N_22884);
xor UO_1303 (O_1303,N_24951,N_23527);
or UO_1304 (O_1304,N_24575,N_23770);
nand UO_1305 (O_1305,N_24531,N_23365);
nor UO_1306 (O_1306,N_24502,N_22602);
and UO_1307 (O_1307,N_24646,N_24498);
xnor UO_1308 (O_1308,N_24054,N_24906);
and UO_1309 (O_1309,N_24945,N_23716);
nand UO_1310 (O_1310,N_24627,N_24114);
nor UO_1311 (O_1311,N_24224,N_23447);
and UO_1312 (O_1312,N_23702,N_23045);
and UO_1313 (O_1313,N_23090,N_24851);
and UO_1314 (O_1314,N_24837,N_24188);
and UO_1315 (O_1315,N_24535,N_24924);
nor UO_1316 (O_1316,N_23795,N_24590);
and UO_1317 (O_1317,N_23079,N_23616);
or UO_1318 (O_1318,N_23656,N_23665);
nor UO_1319 (O_1319,N_24676,N_24006);
and UO_1320 (O_1320,N_23375,N_23444);
nor UO_1321 (O_1321,N_22994,N_22527);
or UO_1322 (O_1322,N_24874,N_23144);
nor UO_1323 (O_1323,N_24777,N_22624);
and UO_1324 (O_1324,N_23551,N_24969);
or UO_1325 (O_1325,N_24052,N_22736);
or UO_1326 (O_1326,N_23834,N_24094);
or UO_1327 (O_1327,N_23407,N_23528);
xor UO_1328 (O_1328,N_23825,N_22731);
xnor UO_1329 (O_1329,N_23367,N_23310);
nor UO_1330 (O_1330,N_22732,N_24293);
or UO_1331 (O_1331,N_23612,N_22512);
and UO_1332 (O_1332,N_24766,N_24472);
xnor UO_1333 (O_1333,N_24090,N_23262);
nor UO_1334 (O_1334,N_23696,N_24133);
nor UO_1335 (O_1335,N_23599,N_23951);
xor UO_1336 (O_1336,N_23588,N_24335);
and UO_1337 (O_1337,N_24582,N_24986);
nor UO_1338 (O_1338,N_23513,N_23663);
nand UO_1339 (O_1339,N_23093,N_24743);
xnor UO_1340 (O_1340,N_23319,N_24716);
nor UO_1341 (O_1341,N_23725,N_24864);
or UO_1342 (O_1342,N_22652,N_23850);
xor UO_1343 (O_1343,N_22504,N_23015);
nand UO_1344 (O_1344,N_23845,N_23367);
nor UO_1345 (O_1345,N_23397,N_24508);
nor UO_1346 (O_1346,N_24322,N_24310);
or UO_1347 (O_1347,N_22849,N_24729);
nor UO_1348 (O_1348,N_23672,N_24978);
or UO_1349 (O_1349,N_24264,N_22736);
and UO_1350 (O_1350,N_24232,N_22802);
nand UO_1351 (O_1351,N_23756,N_24170);
and UO_1352 (O_1352,N_22690,N_24005);
nand UO_1353 (O_1353,N_23831,N_24019);
nand UO_1354 (O_1354,N_22689,N_24518);
or UO_1355 (O_1355,N_24575,N_23935);
nor UO_1356 (O_1356,N_24652,N_22982);
and UO_1357 (O_1357,N_22695,N_23611);
and UO_1358 (O_1358,N_24820,N_23531);
xnor UO_1359 (O_1359,N_24729,N_24314);
nor UO_1360 (O_1360,N_24296,N_23457);
or UO_1361 (O_1361,N_24892,N_24514);
nand UO_1362 (O_1362,N_24528,N_24596);
or UO_1363 (O_1363,N_23114,N_23680);
nor UO_1364 (O_1364,N_23090,N_23622);
or UO_1365 (O_1365,N_24349,N_24371);
and UO_1366 (O_1366,N_24877,N_24424);
and UO_1367 (O_1367,N_24876,N_22838);
nand UO_1368 (O_1368,N_23329,N_24775);
nand UO_1369 (O_1369,N_24719,N_23518);
nand UO_1370 (O_1370,N_24742,N_24868);
nor UO_1371 (O_1371,N_24157,N_23864);
nor UO_1372 (O_1372,N_23062,N_23369);
or UO_1373 (O_1373,N_22633,N_22508);
and UO_1374 (O_1374,N_22734,N_22570);
nor UO_1375 (O_1375,N_22683,N_23305);
or UO_1376 (O_1376,N_22720,N_23439);
nand UO_1377 (O_1377,N_23391,N_23275);
nor UO_1378 (O_1378,N_24395,N_24979);
or UO_1379 (O_1379,N_23805,N_24353);
nor UO_1380 (O_1380,N_22858,N_24460);
nor UO_1381 (O_1381,N_22874,N_23279);
nor UO_1382 (O_1382,N_24099,N_23099);
nor UO_1383 (O_1383,N_24064,N_24770);
nor UO_1384 (O_1384,N_22535,N_24808);
or UO_1385 (O_1385,N_24666,N_23654);
or UO_1386 (O_1386,N_23251,N_24705);
nand UO_1387 (O_1387,N_22647,N_23988);
and UO_1388 (O_1388,N_23831,N_22820);
or UO_1389 (O_1389,N_24434,N_23316);
or UO_1390 (O_1390,N_24356,N_23334);
or UO_1391 (O_1391,N_23699,N_23232);
nor UO_1392 (O_1392,N_22749,N_24028);
nand UO_1393 (O_1393,N_23488,N_23675);
nand UO_1394 (O_1394,N_24151,N_24615);
nor UO_1395 (O_1395,N_24154,N_24548);
nand UO_1396 (O_1396,N_24843,N_22999);
nand UO_1397 (O_1397,N_23031,N_23574);
nor UO_1398 (O_1398,N_22698,N_24408);
xor UO_1399 (O_1399,N_23881,N_24811);
or UO_1400 (O_1400,N_24073,N_24846);
nand UO_1401 (O_1401,N_23749,N_23068);
nand UO_1402 (O_1402,N_24596,N_24760);
nand UO_1403 (O_1403,N_23932,N_23471);
nand UO_1404 (O_1404,N_24652,N_23382);
nand UO_1405 (O_1405,N_24133,N_22540);
nand UO_1406 (O_1406,N_24489,N_24508);
nand UO_1407 (O_1407,N_24945,N_24015);
or UO_1408 (O_1408,N_23178,N_22973);
nor UO_1409 (O_1409,N_24084,N_22918);
nand UO_1410 (O_1410,N_22877,N_23597);
or UO_1411 (O_1411,N_24806,N_23275);
nor UO_1412 (O_1412,N_23761,N_23353);
nand UO_1413 (O_1413,N_24987,N_24920);
xor UO_1414 (O_1414,N_23938,N_24587);
and UO_1415 (O_1415,N_24806,N_23992);
xnor UO_1416 (O_1416,N_24053,N_24775);
and UO_1417 (O_1417,N_23450,N_24091);
and UO_1418 (O_1418,N_23436,N_22798);
or UO_1419 (O_1419,N_22800,N_24531);
and UO_1420 (O_1420,N_24709,N_24876);
nor UO_1421 (O_1421,N_23981,N_24786);
nor UO_1422 (O_1422,N_24540,N_22966);
nor UO_1423 (O_1423,N_24318,N_24238);
nor UO_1424 (O_1424,N_22960,N_24558);
and UO_1425 (O_1425,N_23210,N_23327);
nand UO_1426 (O_1426,N_24595,N_24766);
nor UO_1427 (O_1427,N_23967,N_22887);
or UO_1428 (O_1428,N_23103,N_23802);
nand UO_1429 (O_1429,N_22720,N_22967);
or UO_1430 (O_1430,N_23795,N_22818);
nand UO_1431 (O_1431,N_24591,N_24201);
and UO_1432 (O_1432,N_23754,N_23722);
nor UO_1433 (O_1433,N_22996,N_23805);
and UO_1434 (O_1434,N_24262,N_22770);
or UO_1435 (O_1435,N_22545,N_22912);
nor UO_1436 (O_1436,N_23393,N_24467);
nor UO_1437 (O_1437,N_23987,N_23433);
or UO_1438 (O_1438,N_23827,N_23234);
nor UO_1439 (O_1439,N_24504,N_23748);
nand UO_1440 (O_1440,N_22777,N_23457);
nand UO_1441 (O_1441,N_22722,N_22832);
nand UO_1442 (O_1442,N_23236,N_23066);
and UO_1443 (O_1443,N_23073,N_24028);
nor UO_1444 (O_1444,N_24508,N_23893);
nand UO_1445 (O_1445,N_23477,N_24156);
and UO_1446 (O_1446,N_23874,N_22820);
xor UO_1447 (O_1447,N_23571,N_22972);
nor UO_1448 (O_1448,N_22807,N_22818);
or UO_1449 (O_1449,N_24775,N_22573);
and UO_1450 (O_1450,N_24307,N_24838);
nand UO_1451 (O_1451,N_23432,N_24343);
nand UO_1452 (O_1452,N_23366,N_24698);
or UO_1453 (O_1453,N_23377,N_23035);
or UO_1454 (O_1454,N_24610,N_22785);
nand UO_1455 (O_1455,N_23153,N_23113);
or UO_1456 (O_1456,N_22740,N_22952);
nor UO_1457 (O_1457,N_22618,N_24250);
nand UO_1458 (O_1458,N_22581,N_24194);
xor UO_1459 (O_1459,N_24396,N_24701);
and UO_1460 (O_1460,N_24050,N_23250);
nand UO_1461 (O_1461,N_24834,N_24273);
nor UO_1462 (O_1462,N_23459,N_23517);
or UO_1463 (O_1463,N_23714,N_23975);
nor UO_1464 (O_1464,N_23239,N_24327);
and UO_1465 (O_1465,N_23204,N_23147);
or UO_1466 (O_1466,N_23297,N_23809);
and UO_1467 (O_1467,N_23571,N_24529);
and UO_1468 (O_1468,N_22616,N_23237);
xor UO_1469 (O_1469,N_23777,N_23948);
xnor UO_1470 (O_1470,N_23107,N_24917);
nor UO_1471 (O_1471,N_23750,N_23451);
and UO_1472 (O_1472,N_24590,N_23489);
or UO_1473 (O_1473,N_22831,N_22924);
nand UO_1474 (O_1474,N_23173,N_24156);
or UO_1475 (O_1475,N_23715,N_24602);
nand UO_1476 (O_1476,N_23465,N_24057);
nand UO_1477 (O_1477,N_24031,N_23136);
nand UO_1478 (O_1478,N_24859,N_22820);
and UO_1479 (O_1479,N_23333,N_23262);
or UO_1480 (O_1480,N_23923,N_24904);
nor UO_1481 (O_1481,N_22725,N_23877);
nand UO_1482 (O_1482,N_23878,N_23604);
nand UO_1483 (O_1483,N_23434,N_24727);
and UO_1484 (O_1484,N_23535,N_22800);
nand UO_1485 (O_1485,N_23312,N_24714);
nand UO_1486 (O_1486,N_23115,N_24081);
nand UO_1487 (O_1487,N_22594,N_24720);
xor UO_1488 (O_1488,N_22608,N_22749);
nor UO_1489 (O_1489,N_24374,N_24402);
or UO_1490 (O_1490,N_23851,N_22656);
and UO_1491 (O_1491,N_23112,N_23679);
xnor UO_1492 (O_1492,N_24408,N_22831);
nand UO_1493 (O_1493,N_22836,N_24509);
or UO_1494 (O_1494,N_24465,N_23494);
and UO_1495 (O_1495,N_24944,N_24163);
and UO_1496 (O_1496,N_23026,N_23182);
xor UO_1497 (O_1497,N_22912,N_24913);
nor UO_1498 (O_1498,N_24848,N_24835);
nand UO_1499 (O_1499,N_24838,N_23470);
nand UO_1500 (O_1500,N_23241,N_23396);
or UO_1501 (O_1501,N_24541,N_24497);
nor UO_1502 (O_1502,N_24636,N_24942);
and UO_1503 (O_1503,N_23583,N_23461);
or UO_1504 (O_1504,N_23747,N_23901);
or UO_1505 (O_1505,N_24012,N_24471);
and UO_1506 (O_1506,N_24767,N_22953);
nand UO_1507 (O_1507,N_24253,N_24687);
or UO_1508 (O_1508,N_24193,N_23484);
or UO_1509 (O_1509,N_23379,N_24398);
and UO_1510 (O_1510,N_24019,N_22733);
xnor UO_1511 (O_1511,N_22860,N_24859);
and UO_1512 (O_1512,N_24153,N_23201);
nor UO_1513 (O_1513,N_24538,N_24039);
or UO_1514 (O_1514,N_24273,N_22770);
nand UO_1515 (O_1515,N_24693,N_22778);
nand UO_1516 (O_1516,N_22810,N_23354);
or UO_1517 (O_1517,N_22809,N_24779);
xor UO_1518 (O_1518,N_24032,N_24445);
or UO_1519 (O_1519,N_24454,N_24043);
nand UO_1520 (O_1520,N_24951,N_23274);
xor UO_1521 (O_1521,N_24661,N_24111);
or UO_1522 (O_1522,N_23490,N_23833);
and UO_1523 (O_1523,N_23523,N_22952);
nand UO_1524 (O_1524,N_23358,N_23958);
nor UO_1525 (O_1525,N_23174,N_22819);
and UO_1526 (O_1526,N_23688,N_22885);
and UO_1527 (O_1527,N_24281,N_22763);
nor UO_1528 (O_1528,N_22618,N_23369);
nand UO_1529 (O_1529,N_23531,N_23347);
nor UO_1530 (O_1530,N_24323,N_24347);
nor UO_1531 (O_1531,N_24602,N_24769);
nor UO_1532 (O_1532,N_23157,N_24838);
or UO_1533 (O_1533,N_22841,N_24823);
nor UO_1534 (O_1534,N_24998,N_23740);
xor UO_1535 (O_1535,N_24723,N_23272);
xnor UO_1536 (O_1536,N_24256,N_23713);
nand UO_1537 (O_1537,N_24825,N_23251);
nand UO_1538 (O_1538,N_22899,N_24431);
or UO_1539 (O_1539,N_24843,N_23795);
xnor UO_1540 (O_1540,N_23571,N_22530);
or UO_1541 (O_1541,N_23332,N_24038);
or UO_1542 (O_1542,N_24656,N_22838);
nand UO_1543 (O_1543,N_23584,N_22801);
nor UO_1544 (O_1544,N_24654,N_24030);
or UO_1545 (O_1545,N_24786,N_24951);
nor UO_1546 (O_1546,N_23754,N_22797);
and UO_1547 (O_1547,N_24588,N_22680);
or UO_1548 (O_1548,N_23954,N_24734);
or UO_1549 (O_1549,N_22905,N_22777);
xor UO_1550 (O_1550,N_23878,N_23631);
or UO_1551 (O_1551,N_24055,N_24251);
or UO_1552 (O_1552,N_24469,N_24188);
nor UO_1553 (O_1553,N_23108,N_24630);
or UO_1554 (O_1554,N_22854,N_24553);
and UO_1555 (O_1555,N_24577,N_24827);
nor UO_1556 (O_1556,N_24932,N_24547);
or UO_1557 (O_1557,N_24442,N_24810);
nor UO_1558 (O_1558,N_24267,N_24538);
nand UO_1559 (O_1559,N_23532,N_22802);
nor UO_1560 (O_1560,N_22617,N_24508);
xnor UO_1561 (O_1561,N_24256,N_24684);
nand UO_1562 (O_1562,N_23683,N_22850);
and UO_1563 (O_1563,N_23863,N_24874);
or UO_1564 (O_1564,N_24165,N_24435);
nor UO_1565 (O_1565,N_23342,N_24447);
xor UO_1566 (O_1566,N_23729,N_23553);
and UO_1567 (O_1567,N_23503,N_23466);
and UO_1568 (O_1568,N_22883,N_23175);
and UO_1569 (O_1569,N_23929,N_23694);
nor UO_1570 (O_1570,N_24564,N_24526);
xor UO_1571 (O_1571,N_23955,N_24692);
or UO_1572 (O_1572,N_24723,N_24362);
xnor UO_1573 (O_1573,N_23372,N_23415);
or UO_1574 (O_1574,N_23390,N_24087);
xnor UO_1575 (O_1575,N_24246,N_22763);
and UO_1576 (O_1576,N_22619,N_24439);
or UO_1577 (O_1577,N_23661,N_24661);
nor UO_1578 (O_1578,N_23033,N_24747);
or UO_1579 (O_1579,N_22877,N_22868);
and UO_1580 (O_1580,N_24841,N_23819);
nor UO_1581 (O_1581,N_23673,N_22826);
or UO_1582 (O_1582,N_24970,N_23293);
and UO_1583 (O_1583,N_22655,N_24630);
and UO_1584 (O_1584,N_22526,N_24586);
nand UO_1585 (O_1585,N_24884,N_24779);
and UO_1586 (O_1586,N_22572,N_23757);
nand UO_1587 (O_1587,N_23846,N_22510);
or UO_1588 (O_1588,N_23902,N_24230);
or UO_1589 (O_1589,N_23138,N_23759);
and UO_1590 (O_1590,N_24569,N_23859);
or UO_1591 (O_1591,N_24865,N_23475);
and UO_1592 (O_1592,N_23966,N_24617);
and UO_1593 (O_1593,N_24052,N_22786);
or UO_1594 (O_1594,N_23314,N_24051);
nand UO_1595 (O_1595,N_24747,N_23598);
nand UO_1596 (O_1596,N_24793,N_22807);
or UO_1597 (O_1597,N_23435,N_24490);
nor UO_1598 (O_1598,N_24433,N_23537);
or UO_1599 (O_1599,N_24033,N_23354);
or UO_1600 (O_1600,N_24768,N_23384);
and UO_1601 (O_1601,N_24776,N_23846);
and UO_1602 (O_1602,N_22858,N_23303);
nor UO_1603 (O_1603,N_22752,N_22543);
nand UO_1604 (O_1604,N_23304,N_24219);
and UO_1605 (O_1605,N_24903,N_24095);
or UO_1606 (O_1606,N_23349,N_23937);
xnor UO_1607 (O_1607,N_24904,N_22755);
or UO_1608 (O_1608,N_24153,N_24697);
or UO_1609 (O_1609,N_24696,N_24873);
nand UO_1610 (O_1610,N_24122,N_23107);
nand UO_1611 (O_1611,N_23393,N_24657);
xor UO_1612 (O_1612,N_24222,N_22987);
nand UO_1613 (O_1613,N_24610,N_24578);
and UO_1614 (O_1614,N_23868,N_23546);
nor UO_1615 (O_1615,N_24994,N_23576);
nand UO_1616 (O_1616,N_22970,N_22642);
xor UO_1617 (O_1617,N_24096,N_23366);
or UO_1618 (O_1618,N_23476,N_24632);
nor UO_1619 (O_1619,N_24057,N_23013);
xnor UO_1620 (O_1620,N_23541,N_24992);
nand UO_1621 (O_1621,N_24929,N_23932);
xor UO_1622 (O_1622,N_23903,N_24802);
and UO_1623 (O_1623,N_23982,N_23053);
or UO_1624 (O_1624,N_24615,N_23101);
and UO_1625 (O_1625,N_24971,N_24420);
nand UO_1626 (O_1626,N_23445,N_24463);
and UO_1627 (O_1627,N_22611,N_23255);
nand UO_1628 (O_1628,N_22855,N_23943);
or UO_1629 (O_1629,N_24602,N_23932);
or UO_1630 (O_1630,N_24432,N_24976);
nor UO_1631 (O_1631,N_24363,N_22567);
xor UO_1632 (O_1632,N_24686,N_22918);
or UO_1633 (O_1633,N_24257,N_24394);
nand UO_1634 (O_1634,N_23986,N_22888);
xor UO_1635 (O_1635,N_24400,N_24346);
nand UO_1636 (O_1636,N_22859,N_23959);
and UO_1637 (O_1637,N_23758,N_23143);
nor UO_1638 (O_1638,N_22829,N_24065);
or UO_1639 (O_1639,N_24808,N_24424);
and UO_1640 (O_1640,N_23112,N_24398);
nor UO_1641 (O_1641,N_22695,N_24425);
nor UO_1642 (O_1642,N_24618,N_24753);
or UO_1643 (O_1643,N_23864,N_24194);
or UO_1644 (O_1644,N_22856,N_23742);
and UO_1645 (O_1645,N_23081,N_23664);
nand UO_1646 (O_1646,N_23115,N_24875);
or UO_1647 (O_1647,N_23761,N_23948);
and UO_1648 (O_1648,N_24026,N_23067);
nand UO_1649 (O_1649,N_24324,N_23307);
nor UO_1650 (O_1650,N_22571,N_24216);
nor UO_1651 (O_1651,N_22636,N_22986);
nand UO_1652 (O_1652,N_23641,N_23390);
or UO_1653 (O_1653,N_23446,N_24360);
nor UO_1654 (O_1654,N_23779,N_24632);
xnor UO_1655 (O_1655,N_24481,N_24716);
nor UO_1656 (O_1656,N_22996,N_24248);
and UO_1657 (O_1657,N_23810,N_23538);
and UO_1658 (O_1658,N_24942,N_22886);
and UO_1659 (O_1659,N_24668,N_22954);
and UO_1660 (O_1660,N_22686,N_22648);
or UO_1661 (O_1661,N_23708,N_23174);
and UO_1662 (O_1662,N_23209,N_24559);
and UO_1663 (O_1663,N_22854,N_24449);
nor UO_1664 (O_1664,N_24990,N_22753);
nand UO_1665 (O_1665,N_24859,N_24270);
xnor UO_1666 (O_1666,N_22554,N_24492);
nor UO_1667 (O_1667,N_23787,N_23858);
and UO_1668 (O_1668,N_24495,N_23867);
or UO_1669 (O_1669,N_22600,N_24855);
and UO_1670 (O_1670,N_24558,N_22748);
and UO_1671 (O_1671,N_23944,N_24675);
nand UO_1672 (O_1672,N_22670,N_23156);
and UO_1673 (O_1673,N_24942,N_23383);
nand UO_1674 (O_1674,N_23844,N_23628);
xor UO_1675 (O_1675,N_22867,N_23512);
xor UO_1676 (O_1676,N_24721,N_22824);
nand UO_1677 (O_1677,N_24843,N_22739);
xor UO_1678 (O_1678,N_23982,N_24962);
or UO_1679 (O_1679,N_23981,N_24459);
and UO_1680 (O_1680,N_24168,N_24762);
nor UO_1681 (O_1681,N_23739,N_24159);
nor UO_1682 (O_1682,N_24245,N_24655);
xor UO_1683 (O_1683,N_23160,N_24109);
or UO_1684 (O_1684,N_24108,N_23805);
or UO_1685 (O_1685,N_22813,N_24048);
xnor UO_1686 (O_1686,N_24099,N_23737);
or UO_1687 (O_1687,N_23320,N_24174);
nand UO_1688 (O_1688,N_23721,N_24252);
nand UO_1689 (O_1689,N_24134,N_23839);
xor UO_1690 (O_1690,N_23337,N_24945);
or UO_1691 (O_1691,N_22633,N_23516);
and UO_1692 (O_1692,N_23008,N_23044);
nor UO_1693 (O_1693,N_24299,N_23969);
or UO_1694 (O_1694,N_22710,N_23450);
nand UO_1695 (O_1695,N_24095,N_23663);
nor UO_1696 (O_1696,N_24608,N_23979);
or UO_1697 (O_1697,N_24486,N_24646);
or UO_1698 (O_1698,N_24124,N_23566);
or UO_1699 (O_1699,N_23378,N_24014);
nor UO_1700 (O_1700,N_24783,N_22658);
or UO_1701 (O_1701,N_22610,N_22989);
nand UO_1702 (O_1702,N_23923,N_23734);
and UO_1703 (O_1703,N_22727,N_24683);
nor UO_1704 (O_1704,N_24075,N_23854);
xnor UO_1705 (O_1705,N_24397,N_24119);
nand UO_1706 (O_1706,N_24604,N_24741);
or UO_1707 (O_1707,N_24560,N_22986);
nor UO_1708 (O_1708,N_24551,N_23343);
and UO_1709 (O_1709,N_24974,N_22989);
nor UO_1710 (O_1710,N_24062,N_22503);
nand UO_1711 (O_1711,N_24630,N_22842);
and UO_1712 (O_1712,N_22811,N_23677);
nand UO_1713 (O_1713,N_23697,N_22724);
xnor UO_1714 (O_1714,N_24008,N_23459);
nor UO_1715 (O_1715,N_24741,N_24545);
or UO_1716 (O_1716,N_22954,N_23990);
and UO_1717 (O_1717,N_24841,N_22668);
and UO_1718 (O_1718,N_23242,N_23425);
or UO_1719 (O_1719,N_23073,N_24815);
or UO_1720 (O_1720,N_22984,N_24989);
or UO_1721 (O_1721,N_24226,N_23787);
nand UO_1722 (O_1722,N_23935,N_24605);
nand UO_1723 (O_1723,N_22619,N_24063);
nor UO_1724 (O_1724,N_23176,N_24856);
nand UO_1725 (O_1725,N_23181,N_24373);
xnor UO_1726 (O_1726,N_23272,N_24348);
or UO_1727 (O_1727,N_23934,N_24966);
nand UO_1728 (O_1728,N_23780,N_22942);
nand UO_1729 (O_1729,N_24363,N_24773);
nand UO_1730 (O_1730,N_23676,N_23646);
nand UO_1731 (O_1731,N_22521,N_23322);
or UO_1732 (O_1732,N_24385,N_23380);
and UO_1733 (O_1733,N_22957,N_23727);
nand UO_1734 (O_1734,N_24975,N_22637);
nand UO_1735 (O_1735,N_23888,N_23686);
nand UO_1736 (O_1736,N_24922,N_24819);
nand UO_1737 (O_1737,N_23448,N_24569);
or UO_1738 (O_1738,N_23400,N_24363);
nand UO_1739 (O_1739,N_22651,N_24589);
or UO_1740 (O_1740,N_24557,N_23500);
nand UO_1741 (O_1741,N_23719,N_23788);
or UO_1742 (O_1742,N_23766,N_23520);
and UO_1743 (O_1743,N_24460,N_24931);
and UO_1744 (O_1744,N_23949,N_23977);
nor UO_1745 (O_1745,N_23857,N_22652);
or UO_1746 (O_1746,N_22563,N_23001);
nor UO_1747 (O_1747,N_24384,N_22738);
or UO_1748 (O_1748,N_24630,N_23001);
nand UO_1749 (O_1749,N_23840,N_23032);
or UO_1750 (O_1750,N_22786,N_23587);
or UO_1751 (O_1751,N_23898,N_24834);
and UO_1752 (O_1752,N_23792,N_23093);
or UO_1753 (O_1753,N_23141,N_24750);
nor UO_1754 (O_1754,N_22867,N_24846);
nand UO_1755 (O_1755,N_23869,N_22765);
and UO_1756 (O_1756,N_22580,N_23179);
nor UO_1757 (O_1757,N_23257,N_22591);
or UO_1758 (O_1758,N_24785,N_24777);
nand UO_1759 (O_1759,N_22559,N_23717);
nand UO_1760 (O_1760,N_24389,N_22609);
nor UO_1761 (O_1761,N_24729,N_23685);
nor UO_1762 (O_1762,N_23837,N_23625);
nor UO_1763 (O_1763,N_23917,N_24231);
and UO_1764 (O_1764,N_22649,N_22710);
nand UO_1765 (O_1765,N_24832,N_23512);
xor UO_1766 (O_1766,N_22562,N_22518);
and UO_1767 (O_1767,N_24828,N_24911);
or UO_1768 (O_1768,N_24572,N_23363);
nand UO_1769 (O_1769,N_23038,N_24637);
nand UO_1770 (O_1770,N_23166,N_22617);
nand UO_1771 (O_1771,N_23084,N_23062);
nor UO_1772 (O_1772,N_24305,N_24332);
nand UO_1773 (O_1773,N_22643,N_24201);
and UO_1774 (O_1774,N_22760,N_23459);
or UO_1775 (O_1775,N_24542,N_24842);
nand UO_1776 (O_1776,N_24662,N_23294);
or UO_1777 (O_1777,N_23598,N_23173);
nor UO_1778 (O_1778,N_23177,N_22760);
and UO_1779 (O_1779,N_24470,N_24694);
nand UO_1780 (O_1780,N_23024,N_22688);
nand UO_1781 (O_1781,N_23119,N_24573);
nor UO_1782 (O_1782,N_23642,N_23870);
and UO_1783 (O_1783,N_22577,N_24863);
and UO_1784 (O_1784,N_23866,N_22922);
or UO_1785 (O_1785,N_23931,N_22786);
nor UO_1786 (O_1786,N_24503,N_24679);
or UO_1787 (O_1787,N_23863,N_24017);
nand UO_1788 (O_1788,N_22771,N_24114);
nor UO_1789 (O_1789,N_22690,N_23461);
nor UO_1790 (O_1790,N_24252,N_23778);
and UO_1791 (O_1791,N_23406,N_24770);
nor UO_1792 (O_1792,N_24807,N_24385);
and UO_1793 (O_1793,N_24453,N_24101);
and UO_1794 (O_1794,N_24376,N_24982);
or UO_1795 (O_1795,N_23308,N_24014);
or UO_1796 (O_1796,N_24287,N_24314);
nor UO_1797 (O_1797,N_24423,N_24649);
or UO_1798 (O_1798,N_22824,N_23617);
or UO_1799 (O_1799,N_24367,N_24331);
nand UO_1800 (O_1800,N_23529,N_23840);
nand UO_1801 (O_1801,N_23307,N_23065);
and UO_1802 (O_1802,N_24415,N_24504);
nor UO_1803 (O_1803,N_23406,N_24434);
nor UO_1804 (O_1804,N_24623,N_24151);
or UO_1805 (O_1805,N_24196,N_22642);
or UO_1806 (O_1806,N_23431,N_22573);
nor UO_1807 (O_1807,N_23135,N_24564);
or UO_1808 (O_1808,N_23630,N_22620);
nand UO_1809 (O_1809,N_22770,N_24595);
and UO_1810 (O_1810,N_24626,N_24985);
nor UO_1811 (O_1811,N_23165,N_23366);
nor UO_1812 (O_1812,N_22761,N_24613);
and UO_1813 (O_1813,N_23836,N_24645);
or UO_1814 (O_1814,N_23268,N_24876);
and UO_1815 (O_1815,N_24290,N_22717);
xnor UO_1816 (O_1816,N_23451,N_24295);
xnor UO_1817 (O_1817,N_23316,N_24508);
nand UO_1818 (O_1818,N_24893,N_24837);
xnor UO_1819 (O_1819,N_24406,N_23222);
nor UO_1820 (O_1820,N_23215,N_23609);
nand UO_1821 (O_1821,N_22841,N_22979);
xor UO_1822 (O_1822,N_23320,N_22988);
nand UO_1823 (O_1823,N_23257,N_23269);
and UO_1824 (O_1824,N_24668,N_24078);
nand UO_1825 (O_1825,N_23377,N_22516);
or UO_1826 (O_1826,N_23513,N_24864);
or UO_1827 (O_1827,N_23501,N_23530);
nor UO_1828 (O_1828,N_22724,N_24288);
and UO_1829 (O_1829,N_23985,N_23081);
or UO_1830 (O_1830,N_24551,N_23541);
nand UO_1831 (O_1831,N_23341,N_24939);
and UO_1832 (O_1832,N_22689,N_23556);
and UO_1833 (O_1833,N_22755,N_24881);
nand UO_1834 (O_1834,N_24067,N_24064);
and UO_1835 (O_1835,N_24996,N_23351);
and UO_1836 (O_1836,N_23883,N_22587);
and UO_1837 (O_1837,N_24032,N_23935);
xnor UO_1838 (O_1838,N_22889,N_24730);
nor UO_1839 (O_1839,N_24923,N_22987);
or UO_1840 (O_1840,N_23976,N_24527);
and UO_1841 (O_1841,N_24235,N_23968);
and UO_1842 (O_1842,N_24542,N_24806);
or UO_1843 (O_1843,N_23719,N_24044);
nor UO_1844 (O_1844,N_22537,N_23415);
nor UO_1845 (O_1845,N_23191,N_24888);
nor UO_1846 (O_1846,N_24090,N_24613);
nor UO_1847 (O_1847,N_24686,N_24088);
nand UO_1848 (O_1848,N_22622,N_23395);
nand UO_1849 (O_1849,N_23917,N_24811);
nand UO_1850 (O_1850,N_23849,N_22620);
nand UO_1851 (O_1851,N_24377,N_24823);
and UO_1852 (O_1852,N_24551,N_23250);
nand UO_1853 (O_1853,N_24887,N_23902);
or UO_1854 (O_1854,N_24090,N_23909);
nand UO_1855 (O_1855,N_23216,N_23338);
and UO_1856 (O_1856,N_22973,N_22518);
or UO_1857 (O_1857,N_22707,N_24492);
nor UO_1858 (O_1858,N_23180,N_22920);
nand UO_1859 (O_1859,N_22621,N_24819);
nand UO_1860 (O_1860,N_24100,N_23666);
or UO_1861 (O_1861,N_24204,N_23120);
or UO_1862 (O_1862,N_24417,N_24626);
nor UO_1863 (O_1863,N_23674,N_23510);
xnor UO_1864 (O_1864,N_24959,N_23457);
and UO_1865 (O_1865,N_23959,N_24995);
nand UO_1866 (O_1866,N_22613,N_22666);
and UO_1867 (O_1867,N_23431,N_22696);
nand UO_1868 (O_1868,N_22623,N_23157);
nand UO_1869 (O_1869,N_23476,N_23407);
xor UO_1870 (O_1870,N_23181,N_24023);
nor UO_1871 (O_1871,N_24462,N_24934);
and UO_1872 (O_1872,N_24448,N_24783);
nor UO_1873 (O_1873,N_23580,N_24699);
nor UO_1874 (O_1874,N_23594,N_23270);
or UO_1875 (O_1875,N_24082,N_22732);
nand UO_1876 (O_1876,N_23895,N_22957);
or UO_1877 (O_1877,N_22670,N_23401);
nor UO_1878 (O_1878,N_22979,N_24220);
nor UO_1879 (O_1879,N_22536,N_24734);
and UO_1880 (O_1880,N_24277,N_23828);
and UO_1881 (O_1881,N_22900,N_23253);
nor UO_1882 (O_1882,N_22761,N_22899);
xnor UO_1883 (O_1883,N_24976,N_24196);
nor UO_1884 (O_1884,N_24175,N_24270);
or UO_1885 (O_1885,N_24777,N_23376);
nor UO_1886 (O_1886,N_23191,N_24238);
or UO_1887 (O_1887,N_23614,N_23710);
nand UO_1888 (O_1888,N_24649,N_23442);
nand UO_1889 (O_1889,N_23526,N_24648);
and UO_1890 (O_1890,N_24830,N_24787);
nor UO_1891 (O_1891,N_24967,N_24981);
and UO_1892 (O_1892,N_23578,N_24712);
and UO_1893 (O_1893,N_22594,N_23944);
and UO_1894 (O_1894,N_24131,N_24309);
or UO_1895 (O_1895,N_24616,N_24047);
or UO_1896 (O_1896,N_23919,N_22553);
nor UO_1897 (O_1897,N_24958,N_23518);
nand UO_1898 (O_1898,N_22750,N_22864);
xor UO_1899 (O_1899,N_22571,N_24503);
nor UO_1900 (O_1900,N_24577,N_23710);
or UO_1901 (O_1901,N_24013,N_23456);
and UO_1902 (O_1902,N_23862,N_24076);
nand UO_1903 (O_1903,N_24397,N_24773);
nor UO_1904 (O_1904,N_22673,N_23285);
or UO_1905 (O_1905,N_24999,N_23082);
nor UO_1906 (O_1906,N_24429,N_23785);
nor UO_1907 (O_1907,N_24843,N_24909);
and UO_1908 (O_1908,N_22514,N_24088);
and UO_1909 (O_1909,N_24908,N_24286);
or UO_1910 (O_1910,N_24779,N_22873);
nor UO_1911 (O_1911,N_23361,N_22955);
and UO_1912 (O_1912,N_22607,N_23896);
or UO_1913 (O_1913,N_23271,N_24204);
and UO_1914 (O_1914,N_22646,N_23775);
and UO_1915 (O_1915,N_22886,N_23595);
or UO_1916 (O_1916,N_23732,N_24253);
and UO_1917 (O_1917,N_23561,N_22835);
and UO_1918 (O_1918,N_24364,N_24228);
and UO_1919 (O_1919,N_22871,N_24689);
nand UO_1920 (O_1920,N_24259,N_23837);
or UO_1921 (O_1921,N_23301,N_22565);
and UO_1922 (O_1922,N_24572,N_24556);
or UO_1923 (O_1923,N_24502,N_22973);
nor UO_1924 (O_1924,N_23575,N_24251);
nor UO_1925 (O_1925,N_24770,N_24037);
or UO_1926 (O_1926,N_23482,N_22795);
nand UO_1927 (O_1927,N_23126,N_23590);
and UO_1928 (O_1928,N_22523,N_23906);
or UO_1929 (O_1929,N_23530,N_24227);
nand UO_1930 (O_1930,N_23995,N_22643);
or UO_1931 (O_1931,N_24905,N_23122);
or UO_1932 (O_1932,N_23046,N_24433);
or UO_1933 (O_1933,N_24381,N_24656);
nor UO_1934 (O_1934,N_24244,N_22930);
and UO_1935 (O_1935,N_24760,N_23910);
or UO_1936 (O_1936,N_23245,N_24256);
or UO_1937 (O_1937,N_22528,N_23251);
or UO_1938 (O_1938,N_24866,N_23855);
nand UO_1939 (O_1939,N_24559,N_22718);
or UO_1940 (O_1940,N_24040,N_24325);
nor UO_1941 (O_1941,N_24791,N_22503);
nand UO_1942 (O_1942,N_23169,N_24160);
nand UO_1943 (O_1943,N_23787,N_22885);
nand UO_1944 (O_1944,N_24863,N_24132);
or UO_1945 (O_1945,N_24557,N_23426);
nor UO_1946 (O_1946,N_24597,N_23537);
or UO_1947 (O_1947,N_23809,N_22996);
nand UO_1948 (O_1948,N_24455,N_22813);
nor UO_1949 (O_1949,N_24975,N_24409);
nor UO_1950 (O_1950,N_23975,N_22888);
nand UO_1951 (O_1951,N_23896,N_22881);
and UO_1952 (O_1952,N_22837,N_22923);
and UO_1953 (O_1953,N_23117,N_24034);
nor UO_1954 (O_1954,N_24475,N_23182);
nor UO_1955 (O_1955,N_24256,N_23074);
and UO_1956 (O_1956,N_24536,N_24096);
nor UO_1957 (O_1957,N_24674,N_24689);
or UO_1958 (O_1958,N_23304,N_22514);
nor UO_1959 (O_1959,N_22989,N_24850);
xnor UO_1960 (O_1960,N_23254,N_24468);
nor UO_1961 (O_1961,N_23900,N_23076);
or UO_1962 (O_1962,N_24610,N_24016);
nand UO_1963 (O_1963,N_22572,N_23293);
or UO_1964 (O_1964,N_23732,N_24604);
nor UO_1965 (O_1965,N_23230,N_24418);
nor UO_1966 (O_1966,N_24006,N_23012);
nor UO_1967 (O_1967,N_23322,N_24352);
and UO_1968 (O_1968,N_24026,N_24077);
or UO_1969 (O_1969,N_24529,N_23572);
nand UO_1970 (O_1970,N_24287,N_23302);
nor UO_1971 (O_1971,N_24770,N_24508);
xor UO_1972 (O_1972,N_24543,N_22568);
nor UO_1973 (O_1973,N_23389,N_23788);
or UO_1974 (O_1974,N_22787,N_24856);
and UO_1975 (O_1975,N_24966,N_23012);
nand UO_1976 (O_1976,N_24442,N_24690);
xnor UO_1977 (O_1977,N_23210,N_23569);
and UO_1978 (O_1978,N_23284,N_23777);
or UO_1979 (O_1979,N_23883,N_23247);
nand UO_1980 (O_1980,N_24150,N_24456);
and UO_1981 (O_1981,N_22871,N_22958);
and UO_1982 (O_1982,N_24352,N_23579);
nand UO_1983 (O_1983,N_24551,N_23170);
nor UO_1984 (O_1984,N_23664,N_24144);
or UO_1985 (O_1985,N_22501,N_23750);
or UO_1986 (O_1986,N_23081,N_24499);
and UO_1987 (O_1987,N_23283,N_23975);
and UO_1988 (O_1988,N_22609,N_23158);
nand UO_1989 (O_1989,N_24767,N_24053);
xnor UO_1990 (O_1990,N_22569,N_23536);
and UO_1991 (O_1991,N_23115,N_23684);
nand UO_1992 (O_1992,N_23253,N_24053);
or UO_1993 (O_1993,N_23719,N_23537);
or UO_1994 (O_1994,N_23613,N_22676);
and UO_1995 (O_1995,N_22854,N_24315);
or UO_1996 (O_1996,N_23564,N_24153);
nor UO_1997 (O_1997,N_24890,N_24785);
nand UO_1998 (O_1998,N_22532,N_24936);
and UO_1999 (O_1999,N_22950,N_24210);
nor UO_2000 (O_2000,N_22806,N_23029);
or UO_2001 (O_2001,N_23142,N_24152);
or UO_2002 (O_2002,N_24017,N_24121);
or UO_2003 (O_2003,N_24159,N_24641);
nor UO_2004 (O_2004,N_22507,N_23631);
and UO_2005 (O_2005,N_22778,N_24320);
and UO_2006 (O_2006,N_24634,N_24601);
nand UO_2007 (O_2007,N_24882,N_23054);
or UO_2008 (O_2008,N_22706,N_23312);
xor UO_2009 (O_2009,N_23360,N_23873);
nand UO_2010 (O_2010,N_24808,N_24798);
nor UO_2011 (O_2011,N_24967,N_22884);
xnor UO_2012 (O_2012,N_24152,N_24893);
nand UO_2013 (O_2013,N_24905,N_23415);
nand UO_2014 (O_2014,N_24066,N_23980);
and UO_2015 (O_2015,N_22944,N_23113);
nand UO_2016 (O_2016,N_24889,N_22799);
nand UO_2017 (O_2017,N_23678,N_24603);
and UO_2018 (O_2018,N_22573,N_23405);
or UO_2019 (O_2019,N_24378,N_24035);
nor UO_2020 (O_2020,N_22994,N_24684);
and UO_2021 (O_2021,N_22963,N_23668);
or UO_2022 (O_2022,N_23644,N_22926);
xnor UO_2023 (O_2023,N_23045,N_24686);
or UO_2024 (O_2024,N_24072,N_23668);
and UO_2025 (O_2025,N_24686,N_23491);
xor UO_2026 (O_2026,N_23847,N_23073);
nand UO_2027 (O_2027,N_23835,N_23125);
or UO_2028 (O_2028,N_24806,N_22974);
and UO_2029 (O_2029,N_23764,N_24968);
and UO_2030 (O_2030,N_24601,N_22564);
and UO_2031 (O_2031,N_24032,N_24223);
nand UO_2032 (O_2032,N_22992,N_24959);
nor UO_2033 (O_2033,N_23377,N_24090);
xor UO_2034 (O_2034,N_24027,N_23003);
or UO_2035 (O_2035,N_24816,N_24543);
nor UO_2036 (O_2036,N_24677,N_24177);
xnor UO_2037 (O_2037,N_23599,N_24300);
xnor UO_2038 (O_2038,N_23449,N_24890);
nor UO_2039 (O_2039,N_24673,N_23732);
and UO_2040 (O_2040,N_23032,N_24217);
and UO_2041 (O_2041,N_23235,N_23854);
and UO_2042 (O_2042,N_22586,N_22519);
xnor UO_2043 (O_2043,N_24650,N_24166);
nand UO_2044 (O_2044,N_22527,N_23932);
nor UO_2045 (O_2045,N_23436,N_24983);
or UO_2046 (O_2046,N_23778,N_24377);
or UO_2047 (O_2047,N_22828,N_24405);
xor UO_2048 (O_2048,N_22768,N_23091);
and UO_2049 (O_2049,N_23949,N_22642);
or UO_2050 (O_2050,N_23952,N_23023);
nor UO_2051 (O_2051,N_24677,N_24105);
or UO_2052 (O_2052,N_24461,N_23794);
nand UO_2053 (O_2053,N_24254,N_24174);
nor UO_2054 (O_2054,N_23592,N_22784);
or UO_2055 (O_2055,N_24864,N_24949);
nor UO_2056 (O_2056,N_24818,N_22984);
nand UO_2057 (O_2057,N_23599,N_22605);
nand UO_2058 (O_2058,N_24193,N_22884);
and UO_2059 (O_2059,N_24696,N_23540);
or UO_2060 (O_2060,N_23363,N_24729);
xor UO_2061 (O_2061,N_23643,N_22590);
xnor UO_2062 (O_2062,N_23421,N_24307);
nor UO_2063 (O_2063,N_22764,N_23141);
and UO_2064 (O_2064,N_24252,N_24056);
nor UO_2065 (O_2065,N_24003,N_22623);
or UO_2066 (O_2066,N_23143,N_22610);
nand UO_2067 (O_2067,N_24316,N_24694);
nor UO_2068 (O_2068,N_22937,N_24911);
nand UO_2069 (O_2069,N_23245,N_24176);
nand UO_2070 (O_2070,N_22629,N_23101);
or UO_2071 (O_2071,N_24122,N_23790);
and UO_2072 (O_2072,N_23341,N_23805);
nand UO_2073 (O_2073,N_22691,N_22963);
nand UO_2074 (O_2074,N_24857,N_24530);
nor UO_2075 (O_2075,N_24631,N_23789);
nand UO_2076 (O_2076,N_24369,N_24300);
or UO_2077 (O_2077,N_24344,N_23581);
nor UO_2078 (O_2078,N_23770,N_24613);
xnor UO_2079 (O_2079,N_24497,N_23745);
and UO_2080 (O_2080,N_23737,N_24991);
xnor UO_2081 (O_2081,N_24716,N_23771);
nor UO_2082 (O_2082,N_24622,N_24558);
and UO_2083 (O_2083,N_24136,N_23135);
or UO_2084 (O_2084,N_23087,N_24448);
or UO_2085 (O_2085,N_24228,N_23455);
and UO_2086 (O_2086,N_23185,N_24477);
xnor UO_2087 (O_2087,N_23356,N_22732);
nand UO_2088 (O_2088,N_23449,N_24885);
nand UO_2089 (O_2089,N_24506,N_23743);
nand UO_2090 (O_2090,N_22730,N_24979);
nand UO_2091 (O_2091,N_23289,N_24427);
or UO_2092 (O_2092,N_22789,N_22866);
nand UO_2093 (O_2093,N_22799,N_24942);
nand UO_2094 (O_2094,N_23710,N_24376);
or UO_2095 (O_2095,N_22610,N_23808);
nor UO_2096 (O_2096,N_23560,N_22590);
or UO_2097 (O_2097,N_24343,N_22527);
and UO_2098 (O_2098,N_23600,N_23569);
or UO_2099 (O_2099,N_24682,N_23338);
or UO_2100 (O_2100,N_23031,N_23359);
nor UO_2101 (O_2101,N_24418,N_22817);
or UO_2102 (O_2102,N_23173,N_23744);
or UO_2103 (O_2103,N_23712,N_24474);
and UO_2104 (O_2104,N_24273,N_23204);
nor UO_2105 (O_2105,N_22687,N_23070);
nand UO_2106 (O_2106,N_23350,N_24154);
nor UO_2107 (O_2107,N_24135,N_24792);
or UO_2108 (O_2108,N_22560,N_24253);
and UO_2109 (O_2109,N_23558,N_23806);
and UO_2110 (O_2110,N_24717,N_24014);
or UO_2111 (O_2111,N_24437,N_24146);
and UO_2112 (O_2112,N_24223,N_23144);
and UO_2113 (O_2113,N_22889,N_24319);
nor UO_2114 (O_2114,N_24995,N_23499);
nor UO_2115 (O_2115,N_24209,N_23806);
xor UO_2116 (O_2116,N_23507,N_24728);
and UO_2117 (O_2117,N_23066,N_23024);
and UO_2118 (O_2118,N_22553,N_23042);
nand UO_2119 (O_2119,N_23266,N_24847);
nor UO_2120 (O_2120,N_24743,N_22696);
xor UO_2121 (O_2121,N_22928,N_23176);
and UO_2122 (O_2122,N_22785,N_23944);
nand UO_2123 (O_2123,N_24138,N_22851);
nor UO_2124 (O_2124,N_24314,N_22974);
nand UO_2125 (O_2125,N_24035,N_22798);
nand UO_2126 (O_2126,N_24812,N_23025);
nand UO_2127 (O_2127,N_24729,N_23161);
nand UO_2128 (O_2128,N_22902,N_23632);
nor UO_2129 (O_2129,N_23116,N_24515);
or UO_2130 (O_2130,N_24238,N_24354);
or UO_2131 (O_2131,N_24383,N_24996);
nor UO_2132 (O_2132,N_23314,N_23036);
nand UO_2133 (O_2133,N_24798,N_23840);
and UO_2134 (O_2134,N_22643,N_24789);
and UO_2135 (O_2135,N_24640,N_23630);
and UO_2136 (O_2136,N_23574,N_22738);
or UO_2137 (O_2137,N_23212,N_24676);
and UO_2138 (O_2138,N_22561,N_22637);
nand UO_2139 (O_2139,N_24237,N_23202);
nand UO_2140 (O_2140,N_23952,N_24727);
or UO_2141 (O_2141,N_24331,N_23425);
and UO_2142 (O_2142,N_23939,N_24887);
nand UO_2143 (O_2143,N_22855,N_22994);
nor UO_2144 (O_2144,N_22924,N_24892);
nand UO_2145 (O_2145,N_23824,N_24695);
or UO_2146 (O_2146,N_24993,N_23147);
and UO_2147 (O_2147,N_23992,N_22570);
nand UO_2148 (O_2148,N_23448,N_24065);
and UO_2149 (O_2149,N_24303,N_22732);
nand UO_2150 (O_2150,N_24569,N_24628);
and UO_2151 (O_2151,N_22878,N_23704);
and UO_2152 (O_2152,N_22779,N_22995);
and UO_2153 (O_2153,N_24530,N_24495);
nand UO_2154 (O_2154,N_24739,N_24780);
or UO_2155 (O_2155,N_22694,N_24278);
or UO_2156 (O_2156,N_22648,N_24578);
and UO_2157 (O_2157,N_22867,N_23118);
nand UO_2158 (O_2158,N_24932,N_24082);
or UO_2159 (O_2159,N_24512,N_23963);
or UO_2160 (O_2160,N_23584,N_24648);
and UO_2161 (O_2161,N_24034,N_22635);
and UO_2162 (O_2162,N_23766,N_23611);
or UO_2163 (O_2163,N_24943,N_23356);
and UO_2164 (O_2164,N_23519,N_24545);
and UO_2165 (O_2165,N_23387,N_24034);
nand UO_2166 (O_2166,N_23973,N_23205);
or UO_2167 (O_2167,N_22681,N_24863);
and UO_2168 (O_2168,N_24791,N_23803);
nand UO_2169 (O_2169,N_24680,N_24182);
nand UO_2170 (O_2170,N_24236,N_22584);
nor UO_2171 (O_2171,N_23952,N_23613);
and UO_2172 (O_2172,N_23305,N_23853);
nor UO_2173 (O_2173,N_24816,N_23209);
and UO_2174 (O_2174,N_24863,N_24189);
nor UO_2175 (O_2175,N_23187,N_24888);
nand UO_2176 (O_2176,N_24733,N_24341);
nand UO_2177 (O_2177,N_23625,N_24861);
and UO_2178 (O_2178,N_24347,N_24423);
nor UO_2179 (O_2179,N_22640,N_23033);
or UO_2180 (O_2180,N_22554,N_22744);
or UO_2181 (O_2181,N_24628,N_24159);
nor UO_2182 (O_2182,N_23614,N_22631);
nand UO_2183 (O_2183,N_24259,N_24866);
and UO_2184 (O_2184,N_22974,N_23301);
and UO_2185 (O_2185,N_23116,N_22716);
nor UO_2186 (O_2186,N_24032,N_23214);
nand UO_2187 (O_2187,N_23874,N_24421);
and UO_2188 (O_2188,N_23722,N_23340);
and UO_2189 (O_2189,N_24989,N_23728);
or UO_2190 (O_2190,N_22593,N_23505);
nand UO_2191 (O_2191,N_24739,N_23902);
nor UO_2192 (O_2192,N_24014,N_24934);
and UO_2193 (O_2193,N_24292,N_24357);
or UO_2194 (O_2194,N_23962,N_23736);
nand UO_2195 (O_2195,N_22504,N_24710);
or UO_2196 (O_2196,N_24135,N_22888);
nand UO_2197 (O_2197,N_22914,N_24093);
and UO_2198 (O_2198,N_22505,N_23778);
nor UO_2199 (O_2199,N_23955,N_22868);
or UO_2200 (O_2200,N_22527,N_24884);
and UO_2201 (O_2201,N_24175,N_22630);
nor UO_2202 (O_2202,N_22843,N_22842);
nand UO_2203 (O_2203,N_24765,N_23266);
or UO_2204 (O_2204,N_23182,N_23378);
and UO_2205 (O_2205,N_22926,N_23359);
and UO_2206 (O_2206,N_22833,N_24934);
nand UO_2207 (O_2207,N_24066,N_23063);
or UO_2208 (O_2208,N_24229,N_24686);
or UO_2209 (O_2209,N_24427,N_23884);
nor UO_2210 (O_2210,N_24944,N_23705);
and UO_2211 (O_2211,N_23977,N_23951);
nor UO_2212 (O_2212,N_23611,N_23519);
nor UO_2213 (O_2213,N_23379,N_22821);
or UO_2214 (O_2214,N_22902,N_24036);
or UO_2215 (O_2215,N_23512,N_22690);
nor UO_2216 (O_2216,N_24855,N_24359);
nor UO_2217 (O_2217,N_23111,N_23420);
nor UO_2218 (O_2218,N_24050,N_24526);
nand UO_2219 (O_2219,N_22679,N_23480);
and UO_2220 (O_2220,N_22651,N_24871);
or UO_2221 (O_2221,N_23876,N_22854);
nor UO_2222 (O_2222,N_23750,N_23464);
nand UO_2223 (O_2223,N_23184,N_24830);
and UO_2224 (O_2224,N_24654,N_24641);
nand UO_2225 (O_2225,N_23672,N_24728);
nand UO_2226 (O_2226,N_22598,N_23294);
or UO_2227 (O_2227,N_22754,N_22943);
nor UO_2228 (O_2228,N_22699,N_24674);
and UO_2229 (O_2229,N_23780,N_23129);
nor UO_2230 (O_2230,N_24048,N_23931);
xor UO_2231 (O_2231,N_24023,N_22568);
or UO_2232 (O_2232,N_24573,N_24479);
xnor UO_2233 (O_2233,N_24763,N_23878);
xor UO_2234 (O_2234,N_24039,N_24462);
nor UO_2235 (O_2235,N_23330,N_24413);
and UO_2236 (O_2236,N_22562,N_23508);
and UO_2237 (O_2237,N_23880,N_23711);
nor UO_2238 (O_2238,N_23259,N_23249);
nand UO_2239 (O_2239,N_22821,N_24570);
and UO_2240 (O_2240,N_22899,N_24883);
nor UO_2241 (O_2241,N_24037,N_24558);
nor UO_2242 (O_2242,N_24422,N_22846);
nor UO_2243 (O_2243,N_23170,N_23376);
and UO_2244 (O_2244,N_23214,N_22642);
nand UO_2245 (O_2245,N_24392,N_23072);
nor UO_2246 (O_2246,N_23675,N_22512);
nor UO_2247 (O_2247,N_24245,N_24318);
and UO_2248 (O_2248,N_24434,N_22581);
or UO_2249 (O_2249,N_24105,N_23450);
or UO_2250 (O_2250,N_23309,N_24558);
nor UO_2251 (O_2251,N_24068,N_23425);
nor UO_2252 (O_2252,N_22506,N_23417);
xnor UO_2253 (O_2253,N_23060,N_24826);
xor UO_2254 (O_2254,N_23828,N_24885);
nor UO_2255 (O_2255,N_24716,N_24816);
nand UO_2256 (O_2256,N_22628,N_22656);
nor UO_2257 (O_2257,N_22986,N_23530);
nor UO_2258 (O_2258,N_24677,N_23013);
or UO_2259 (O_2259,N_24264,N_24001);
xor UO_2260 (O_2260,N_24937,N_22982);
nand UO_2261 (O_2261,N_24832,N_23969);
nor UO_2262 (O_2262,N_23850,N_23376);
or UO_2263 (O_2263,N_23355,N_24462);
nand UO_2264 (O_2264,N_24990,N_22897);
nand UO_2265 (O_2265,N_24011,N_23368);
or UO_2266 (O_2266,N_24906,N_23408);
or UO_2267 (O_2267,N_22895,N_24987);
nand UO_2268 (O_2268,N_24284,N_22530);
nand UO_2269 (O_2269,N_22745,N_23129);
and UO_2270 (O_2270,N_23165,N_24855);
and UO_2271 (O_2271,N_24569,N_23375);
or UO_2272 (O_2272,N_22999,N_22930);
and UO_2273 (O_2273,N_24370,N_24719);
nand UO_2274 (O_2274,N_23773,N_23575);
and UO_2275 (O_2275,N_23177,N_23757);
nand UO_2276 (O_2276,N_24753,N_23552);
and UO_2277 (O_2277,N_22756,N_23806);
nand UO_2278 (O_2278,N_24811,N_23000);
nor UO_2279 (O_2279,N_24393,N_23660);
nor UO_2280 (O_2280,N_23947,N_24559);
nand UO_2281 (O_2281,N_24475,N_24673);
nor UO_2282 (O_2282,N_23546,N_24503);
or UO_2283 (O_2283,N_24829,N_23310);
nor UO_2284 (O_2284,N_23538,N_24344);
nand UO_2285 (O_2285,N_24200,N_23538);
or UO_2286 (O_2286,N_22925,N_23661);
and UO_2287 (O_2287,N_22726,N_22903);
and UO_2288 (O_2288,N_22878,N_22645);
nand UO_2289 (O_2289,N_23980,N_23193);
nor UO_2290 (O_2290,N_23340,N_23456);
nor UO_2291 (O_2291,N_22670,N_24471);
xnor UO_2292 (O_2292,N_22665,N_22978);
or UO_2293 (O_2293,N_23905,N_22803);
or UO_2294 (O_2294,N_24560,N_24576);
or UO_2295 (O_2295,N_24389,N_24563);
and UO_2296 (O_2296,N_23817,N_23092);
or UO_2297 (O_2297,N_24118,N_23489);
or UO_2298 (O_2298,N_23367,N_24947);
xor UO_2299 (O_2299,N_24519,N_23758);
nand UO_2300 (O_2300,N_22537,N_23861);
nand UO_2301 (O_2301,N_22502,N_24694);
or UO_2302 (O_2302,N_24713,N_23947);
or UO_2303 (O_2303,N_22993,N_23356);
or UO_2304 (O_2304,N_22779,N_24300);
nand UO_2305 (O_2305,N_23441,N_23386);
or UO_2306 (O_2306,N_24348,N_24318);
or UO_2307 (O_2307,N_24183,N_23037);
and UO_2308 (O_2308,N_23340,N_24686);
and UO_2309 (O_2309,N_24199,N_24548);
nor UO_2310 (O_2310,N_22628,N_24250);
or UO_2311 (O_2311,N_24147,N_23070);
or UO_2312 (O_2312,N_23971,N_23905);
xnor UO_2313 (O_2313,N_22646,N_23589);
nor UO_2314 (O_2314,N_24037,N_24532);
and UO_2315 (O_2315,N_23273,N_23436);
nand UO_2316 (O_2316,N_23717,N_24296);
nand UO_2317 (O_2317,N_23740,N_23887);
nor UO_2318 (O_2318,N_24995,N_22668);
or UO_2319 (O_2319,N_22703,N_24282);
nand UO_2320 (O_2320,N_22683,N_23439);
or UO_2321 (O_2321,N_24377,N_23271);
and UO_2322 (O_2322,N_23717,N_24372);
nand UO_2323 (O_2323,N_23782,N_23548);
nor UO_2324 (O_2324,N_24752,N_24620);
nand UO_2325 (O_2325,N_23017,N_23212);
or UO_2326 (O_2326,N_22843,N_23765);
and UO_2327 (O_2327,N_23187,N_23802);
and UO_2328 (O_2328,N_22718,N_23573);
nand UO_2329 (O_2329,N_24479,N_22923);
nor UO_2330 (O_2330,N_23683,N_22813);
or UO_2331 (O_2331,N_23059,N_23840);
nor UO_2332 (O_2332,N_23185,N_24160);
nand UO_2333 (O_2333,N_22810,N_23355);
nor UO_2334 (O_2334,N_22846,N_24274);
nor UO_2335 (O_2335,N_23014,N_24157);
and UO_2336 (O_2336,N_23926,N_24547);
xor UO_2337 (O_2337,N_24156,N_22612);
nand UO_2338 (O_2338,N_22995,N_24831);
xnor UO_2339 (O_2339,N_22557,N_23641);
xor UO_2340 (O_2340,N_23840,N_23528);
and UO_2341 (O_2341,N_23027,N_24467);
nand UO_2342 (O_2342,N_24098,N_24285);
and UO_2343 (O_2343,N_24041,N_24882);
or UO_2344 (O_2344,N_24790,N_23076);
nand UO_2345 (O_2345,N_23855,N_22792);
xnor UO_2346 (O_2346,N_22935,N_23894);
xnor UO_2347 (O_2347,N_24138,N_22625);
and UO_2348 (O_2348,N_22814,N_23021);
nor UO_2349 (O_2349,N_23715,N_23192);
or UO_2350 (O_2350,N_23071,N_24302);
nor UO_2351 (O_2351,N_23291,N_23345);
nand UO_2352 (O_2352,N_23447,N_24558);
or UO_2353 (O_2353,N_23930,N_23588);
or UO_2354 (O_2354,N_22961,N_24693);
or UO_2355 (O_2355,N_24767,N_23552);
nand UO_2356 (O_2356,N_23924,N_24254);
and UO_2357 (O_2357,N_22607,N_23777);
and UO_2358 (O_2358,N_24682,N_22946);
xor UO_2359 (O_2359,N_24988,N_24336);
or UO_2360 (O_2360,N_23208,N_24535);
nand UO_2361 (O_2361,N_24615,N_24544);
or UO_2362 (O_2362,N_23740,N_23844);
xnor UO_2363 (O_2363,N_24386,N_22825);
or UO_2364 (O_2364,N_24092,N_24721);
nor UO_2365 (O_2365,N_22989,N_22666);
nand UO_2366 (O_2366,N_22913,N_22576);
and UO_2367 (O_2367,N_24042,N_24745);
nand UO_2368 (O_2368,N_24314,N_23702);
and UO_2369 (O_2369,N_22902,N_24092);
nor UO_2370 (O_2370,N_23160,N_24575);
or UO_2371 (O_2371,N_23918,N_23149);
nand UO_2372 (O_2372,N_24639,N_23763);
nand UO_2373 (O_2373,N_24298,N_24009);
nand UO_2374 (O_2374,N_23660,N_23160);
nand UO_2375 (O_2375,N_24728,N_23610);
and UO_2376 (O_2376,N_24817,N_24844);
xnor UO_2377 (O_2377,N_24079,N_23355);
nand UO_2378 (O_2378,N_23067,N_23576);
and UO_2379 (O_2379,N_24167,N_22855);
or UO_2380 (O_2380,N_22808,N_22900);
xor UO_2381 (O_2381,N_24349,N_24393);
nor UO_2382 (O_2382,N_23923,N_23748);
nor UO_2383 (O_2383,N_24338,N_23647);
nand UO_2384 (O_2384,N_24556,N_24496);
xnor UO_2385 (O_2385,N_23045,N_23057);
and UO_2386 (O_2386,N_23941,N_24086);
or UO_2387 (O_2387,N_24099,N_23236);
and UO_2388 (O_2388,N_23504,N_24314);
and UO_2389 (O_2389,N_24670,N_24779);
nand UO_2390 (O_2390,N_23908,N_23966);
xor UO_2391 (O_2391,N_24880,N_23592);
or UO_2392 (O_2392,N_24886,N_24020);
and UO_2393 (O_2393,N_23921,N_23686);
or UO_2394 (O_2394,N_24136,N_24389);
nand UO_2395 (O_2395,N_23048,N_24127);
or UO_2396 (O_2396,N_23909,N_23516);
nand UO_2397 (O_2397,N_22894,N_23707);
nor UO_2398 (O_2398,N_22753,N_24014);
nor UO_2399 (O_2399,N_23469,N_23688);
nor UO_2400 (O_2400,N_24414,N_23536);
or UO_2401 (O_2401,N_23162,N_22913);
and UO_2402 (O_2402,N_22977,N_24396);
or UO_2403 (O_2403,N_24870,N_24194);
and UO_2404 (O_2404,N_24346,N_23127);
and UO_2405 (O_2405,N_22669,N_24079);
or UO_2406 (O_2406,N_24238,N_24700);
and UO_2407 (O_2407,N_24681,N_22704);
and UO_2408 (O_2408,N_23510,N_24743);
and UO_2409 (O_2409,N_24214,N_22933);
xnor UO_2410 (O_2410,N_22893,N_24146);
or UO_2411 (O_2411,N_24972,N_24823);
xor UO_2412 (O_2412,N_22575,N_23733);
and UO_2413 (O_2413,N_22569,N_22787);
or UO_2414 (O_2414,N_24790,N_24667);
xor UO_2415 (O_2415,N_24060,N_24843);
or UO_2416 (O_2416,N_22892,N_22751);
or UO_2417 (O_2417,N_24778,N_24645);
or UO_2418 (O_2418,N_22975,N_23643);
and UO_2419 (O_2419,N_23355,N_24256);
nor UO_2420 (O_2420,N_23472,N_23482);
and UO_2421 (O_2421,N_23336,N_24289);
and UO_2422 (O_2422,N_24747,N_22605);
nand UO_2423 (O_2423,N_24700,N_22982);
and UO_2424 (O_2424,N_24850,N_24475);
or UO_2425 (O_2425,N_23271,N_24387);
and UO_2426 (O_2426,N_24362,N_24211);
and UO_2427 (O_2427,N_22931,N_23934);
and UO_2428 (O_2428,N_23181,N_24077);
or UO_2429 (O_2429,N_23290,N_24771);
nand UO_2430 (O_2430,N_23130,N_23329);
nor UO_2431 (O_2431,N_23634,N_23077);
and UO_2432 (O_2432,N_24334,N_24625);
and UO_2433 (O_2433,N_23187,N_24917);
nand UO_2434 (O_2434,N_24372,N_24167);
xor UO_2435 (O_2435,N_24464,N_23411);
xnor UO_2436 (O_2436,N_24561,N_23003);
or UO_2437 (O_2437,N_23177,N_24195);
nand UO_2438 (O_2438,N_22515,N_24150);
nand UO_2439 (O_2439,N_22535,N_22932);
nor UO_2440 (O_2440,N_23204,N_24051);
and UO_2441 (O_2441,N_22874,N_24063);
nor UO_2442 (O_2442,N_22655,N_22811);
or UO_2443 (O_2443,N_24232,N_24737);
nand UO_2444 (O_2444,N_22731,N_23542);
and UO_2445 (O_2445,N_23921,N_23100);
nand UO_2446 (O_2446,N_24268,N_23758);
and UO_2447 (O_2447,N_22674,N_23299);
and UO_2448 (O_2448,N_22975,N_23479);
nor UO_2449 (O_2449,N_23316,N_24285);
or UO_2450 (O_2450,N_24865,N_24073);
xor UO_2451 (O_2451,N_24142,N_24991);
nor UO_2452 (O_2452,N_24024,N_22516);
or UO_2453 (O_2453,N_24661,N_24362);
or UO_2454 (O_2454,N_22866,N_24867);
or UO_2455 (O_2455,N_22501,N_22667);
or UO_2456 (O_2456,N_22701,N_23335);
or UO_2457 (O_2457,N_23703,N_24771);
nand UO_2458 (O_2458,N_23521,N_22725);
and UO_2459 (O_2459,N_24316,N_22997);
nand UO_2460 (O_2460,N_23819,N_23885);
and UO_2461 (O_2461,N_23750,N_24568);
nand UO_2462 (O_2462,N_23613,N_23322);
nand UO_2463 (O_2463,N_24240,N_22936);
and UO_2464 (O_2464,N_24511,N_24355);
or UO_2465 (O_2465,N_23896,N_22553);
or UO_2466 (O_2466,N_24686,N_22685);
nor UO_2467 (O_2467,N_23574,N_23820);
and UO_2468 (O_2468,N_24209,N_22886);
and UO_2469 (O_2469,N_24719,N_23709);
and UO_2470 (O_2470,N_23230,N_23687);
nand UO_2471 (O_2471,N_24346,N_22923);
and UO_2472 (O_2472,N_24983,N_23617);
nand UO_2473 (O_2473,N_24387,N_22516);
and UO_2474 (O_2474,N_23777,N_23075);
or UO_2475 (O_2475,N_23015,N_24811);
or UO_2476 (O_2476,N_22966,N_23866);
nor UO_2477 (O_2477,N_23033,N_23930);
or UO_2478 (O_2478,N_24822,N_23864);
and UO_2479 (O_2479,N_24064,N_24708);
xor UO_2480 (O_2480,N_24397,N_23940);
or UO_2481 (O_2481,N_24692,N_24191);
nor UO_2482 (O_2482,N_24353,N_22980);
nand UO_2483 (O_2483,N_23827,N_24593);
or UO_2484 (O_2484,N_24676,N_23234);
nand UO_2485 (O_2485,N_23379,N_24200);
xor UO_2486 (O_2486,N_23669,N_24064);
or UO_2487 (O_2487,N_22680,N_24420);
and UO_2488 (O_2488,N_22745,N_24258);
nand UO_2489 (O_2489,N_24328,N_24692);
and UO_2490 (O_2490,N_23515,N_24182);
or UO_2491 (O_2491,N_22799,N_23019);
nand UO_2492 (O_2492,N_24730,N_24353);
and UO_2493 (O_2493,N_23257,N_22547);
nor UO_2494 (O_2494,N_22509,N_24918);
nand UO_2495 (O_2495,N_22861,N_24021);
nand UO_2496 (O_2496,N_23933,N_22849);
or UO_2497 (O_2497,N_23467,N_23729);
and UO_2498 (O_2498,N_23069,N_23388);
and UO_2499 (O_2499,N_24324,N_22664);
nand UO_2500 (O_2500,N_24331,N_24324);
and UO_2501 (O_2501,N_24619,N_24333);
and UO_2502 (O_2502,N_24188,N_22893);
and UO_2503 (O_2503,N_23297,N_23681);
nand UO_2504 (O_2504,N_24560,N_23376);
or UO_2505 (O_2505,N_23767,N_23228);
and UO_2506 (O_2506,N_23644,N_22969);
or UO_2507 (O_2507,N_24374,N_23876);
and UO_2508 (O_2508,N_23319,N_23915);
nor UO_2509 (O_2509,N_24095,N_24848);
and UO_2510 (O_2510,N_24052,N_23503);
nand UO_2511 (O_2511,N_24625,N_24955);
or UO_2512 (O_2512,N_22691,N_23455);
and UO_2513 (O_2513,N_23236,N_23588);
nor UO_2514 (O_2514,N_24161,N_23281);
and UO_2515 (O_2515,N_23361,N_22799);
or UO_2516 (O_2516,N_22547,N_22592);
nor UO_2517 (O_2517,N_24012,N_23317);
nor UO_2518 (O_2518,N_23483,N_24708);
nand UO_2519 (O_2519,N_22631,N_24044);
nand UO_2520 (O_2520,N_24077,N_24734);
or UO_2521 (O_2521,N_24733,N_24389);
nor UO_2522 (O_2522,N_24078,N_22859);
or UO_2523 (O_2523,N_24889,N_23909);
and UO_2524 (O_2524,N_22810,N_22563);
nand UO_2525 (O_2525,N_23450,N_24005);
or UO_2526 (O_2526,N_22608,N_23960);
and UO_2527 (O_2527,N_23403,N_24343);
nor UO_2528 (O_2528,N_23078,N_24044);
or UO_2529 (O_2529,N_23822,N_24808);
nor UO_2530 (O_2530,N_24720,N_22915);
or UO_2531 (O_2531,N_24154,N_23472);
and UO_2532 (O_2532,N_24752,N_24717);
or UO_2533 (O_2533,N_24942,N_23044);
nand UO_2534 (O_2534,N_22746,N_24849);
nor UO_2535 (O_2535,N_23589,N_22819);
xor UO_2536 (O_2536,N_24187,N_24678);
and UO_2537 (O_2537,N_23452,N_24977);
and UO_2538 (O_2538,N_23558,N_22850);
nand UO_2539 (O_2539,N_24106,N_24782);
nand UO_2540 (O_2540,N_22566,N_23289);
nand UO_2541 (O_2541,N_24377,N_22835);
xnor UO_2542 (O_2542,N_23470,N_23143);
nand UO_2543 (O_2543,N_23194,N_24409);
and UO_2544 (O_2544,N_22782,N_24494);
and UO_2545 (O_2545,N_23568,N_24426);
nand UO_2546 (O_2546,N_23177,N_24847);
or UO_2547 (O_2547,N_24384,N_24400);
nand UO_2548 (O_2548,N_22504,N_23892);
or UO_2549 (O_2549,N_23313,N_22731);
nand UO_2550 (O_2550,N_24160,N_23663);
and UO_2551 (O_2551,N_23700,N_24042);
or UO_2552 (O_2552,N_22532,N_24515);
nor UO_2553 (O_2553,N_24383,N_24538);
nand UO_2554 (O_2554,N_23221,N_22885);
and UO_2555 (O_2555,N_23493,N_24437);
nor UO_2556 (O_2556,N_23584,N_24402);
nand UO_2557 (O_2557,N_23245,N_23738);
nor UO_2558 (O_2558,N_22845,N_24590);
or UO_2559 (O_2559,N_23162,N_22985);
nor UO_2560 (O_2560,N_22811,N_22983);
or UO_2561 (O_2561,N_23076,N_22985);
nor UO_2562 (O_2562,N_23008,N_24520);
xnor UO_2563 (O_2563,N_23643,N_23489);
nand UO_2564 (O_2564,N_23203,N_23972);
nand UO_2565 (O_2565,N_24134,N_24348);
xnor UO_2566 (O_2566,N_22715,N_22874);
nand UO_2567 (O_2567,N_22795,N_23437);
nor UO_2568 (O_2568,N_23201,N_23651);
nor UO_2569 (O_2569,N_24079,N_23613);
and UO_2570 (O_2570,N_23974,N_24652);
or UO_2571 (O_2571,N_24964,N_24147);
nand UO_2572 (O_2572,N_22722,N_24279);
and UO_2573 (O_2573,N_23637,N_22685);
and UO_2574 (O_2574,N_24658,N_24519);
and UO_2575 (O_2575,N_22711,N_24583);
or UO_2576 (O_2576,N_23675,N_22522);
nand UO_2577 (O_2577,N_23022,N_24230);
and UO_2578 (O_2578,N_23779,N_23133);
or UO_2579 (O_2579,N_24474,N_23213);
nand UO_2580 (O_2580,N_23292,N_24020);
or UO_2581 (O_2581,N_24387,N_23315);
or UO_2582 (O_2582,N_24378,N_22783);
or UO_2583 (O_2583,N_22507,N_23132);
or UO_2584 (O_2584,N_23089,N_23752);
and UO_2585 (O_2585,N_22880,N_23856);
nor UO_2586 (O_2586,N_24684,N_22945);
xor UO_2587 (O_2587,N_23710,N_22673);
nand UO_2588 (O_2588,N_24304,N_24816);
nor UO_2589 (O_2589,N_23440,N_22868);
and UO_2590 (O_2590,N_24853,N_23079);
or UO_2591 (O_2591,N_23267,N_23141);
nor UO_2592 (O_2592,N_24649,N_24954);
nand UO_2593 (O_2593,N_23053,N_22959);
nor UO_2594 (O_2594,N_23950,N_24121);
and UO_2595 (O_2595,N_22846,N_23220);
and UO_2596 (O_2596,N_22758,N_24870);
and UO_2597 (O_2597,N_24361,N_22500);
xor UO_2598 (O_2598,N_23351,N_23278);
or UO_2599 (O_2599,N_23977,N_23553);
and UO_2600 (O_2600,N_23942,N_23708);
nand UO_2601 (O_2601,N_23407,N_24439);
xor UO_2602 (O_2602,N_24790,N_24797);
xnor UO_2603 (O_2603,N_24274,N_23331);
or UO_2604 (O_2604,N_23086,N_24289);
and UO_2605 (O_2605,N_22773,N_22821);
or UO_2606 (O_2606,N_24388,N_24795);
nor UO_2607 (O_2607,N_23884,N_22613);
and UO_2608 (O_2608,N_24016,N_23697);
nand UO_2609 (O_2609,N_24903,N_24191);
nor UO_2610 (O_2610,N_23389,N_23821);
and UO_2611 (O_2611,N_24326,N_23949);
nand UO_2612 (O_2612,N_22961,N_24939);
and UO_2613 (O_2613,N_23794,N_23599);
nor UO_2614 (O_2614,N_23514,N_22711);
nor UO_2615 (O_2615,N_24082,N_23050);
and UO_2616 (O_2616,N_22944,N_24506);
and UO_2617 (O_2617,N_24707,N_23768);
and UO_2618 (O_2618,N_23528,N_23138);
xor UO_2619 (O_2619,N_23998,N_23301);
and UO_2620 (O_2620,N_23448,N_24255);
xnor UO_2621 (O_2621,N_24019,N_23030);
nor UO_2622 (O_2622,N_22619,N_22648);
and UO_2623 (O_2623,N_23846,N_23813);
nand UO_2624 (O_2624,N_24960,N_23923);
nand UO_2625 (O_2625,N_24502,N_24225);
nor UO_2626 (O_2626,N_23318,N_22794);
or UO_2627 (O_2627,N_23809,N_22735);
or UO_2628 (O_2628,N_22807,N_24889);
nand UO_2629 (O_2629,N_23490,N_22684);
or UO_2630 (O_2630,N_23852,N_23025);
xnor UO_2631 (O_2631,N_22565,N_23607);
and UO_2632 (O_2632,N_24075,N_22666);
nand UO_2633 (O_2633,N_24776,N_22815);
nand UO_2634 (O_2634,N_23757,N_23225);
nor UO_2635 (O_2635,N_23609,N_23409);
xor UO_2636 (O_2636,N_24717,N_23662);
nor UO_2637 (O_2637,N_24661,N_23071);
nand UO_2638 (O_2638,N_22961,N_22553);
nor UO_2639 (O_2639,N_23546,N_24065);
or UO_2640 (O_2640,N_24342,N_22542);
nor UO_2641 (O_2641,N_24643,N_23471);
xnor UO_2642 (O_2642,N_23829,N_22501);
or UO_2643 (O_2643,N_23734,N_24694);
and UO_2644 (O_2644,N_24812,N_24189);
or UO_2645 (O_2645,N_24951,N_23448);
and UO_2646 (O_2646,N_23925,N_23012);
xnor UO_2647 (O_2647,N_22699,N_23682);
nor UO_2648 (O_2648,N_23813,N_24795);
nand UO_2649 (O_2649,N_22504,N_22526);
and UO_2650 (O_2650,N_23361,N_23522);
nand UO_2651 (O_2651,N_23396,N_23328);
nor UO_2652 (O_2652,N_22696,N_24449);
or UO_2653 (O_2653,N_24777,N_24156);
nor UO_2654 (O_2654,N_23670,N_24218);
nand UO_2655 (O_2655,N_22754,N_24066);
nand UO_2656 (O_2656,N_23183,N_24398);
or UO_2657 (O_2657,N_24366,N_23349);
and UO_2658 (O_2658,N_23630,N_24890);
or UO_2659 (O_2659,N_22814,N_24663);
or UO_2660 (O_2660,N_23374,N_23461);
nor UO_2661 (O_2661,N_23515,N_23561);
and UO_2662 (O_2662,N_24216,N_23486);
or UO_2663 (O_2663,N_23634,N_24538);
nand UO_2664 (O_2664,N_24396,N_23417);
nor UO_2665 (O_2665,N_24980,N_24564);
and UO_2666 (O_2666,N_24139,N_23931);
or UO_2667 (O_2667,N_24362,N_24906);
or UO_2668 (O_2668,N_24647,N_24481);
nand UO_2669 (O_2669,N_23438,N_22690);
nor UO_2670 (O_2670,N_22732,N_22739);
and UO_2671 (O_2671,N_22825,N_23856);
nand UO_2672 (O_2672,N_24827,N_22526);
or UO_2673 (O_2673,N_24669,N_24389);
or UO_2674 (O_2674,N_23414,N_24797);
or UO_2675 (O_2675,N_22593,N_22619);
nor UO_2676 (O_2676,N_22573,N_23066);
and UO_2677 (O_2677,N_23713,N_24982);
or UO_2678 (O_2678,N_24118,N_24124);
and UO_2679 (O_2679,N_23885,N_24532);
nor UO_2680 (O_2680,N_24854,N_23228);
nand UO_2681 (O_2681,N_23018,N_23319);
nor UO_2682 (O_2682,N_22672,N_22954);
nand UO_2683 (O_2683,N_24281,N_23884);
xor UO_2684 (O_2684,N_23312,N_24744);
and UO_2685 (O_2685,N_23415,N_23867);
or UO_2686 (O_2686,N_22578,N_22501);
nor UO_2687 (O_2687,N_23895,N_23981);
or UO_2688 (O_2688,N_24395,N_24005);
nor UO_2689 (O_2689,N_22538,N_24364);
nand UO_2690 (O_2690,N_24284,N_23312);
nor UO_2691 (O_2691,N_24625,N_22927);
or UO_2692 (O_2692,N_22880,N_23981);
nand UO_2693 (O_2693,N_24459,N_24331);
xor UO_2694 (O_2694,N_22837,N_24564);
and UO_2695 (O_2695,N_23832,N_23982);
nand UO_2696 (O_2696,N_24942,N_22758);
or UO_2697 (O_2697,N_23419,N_23641);
nand UO_2698 (O_2698,N_22965,N_22506);
and UO_2699 (O_2699,N_24381,N_23806);
and UO_2700 (O_2700,N_22759,N_24564);
and UO_2701 (O_2701,N_24790,N_23857);
and UO_2702 (O_2702,N_23887,N_24682);
xor UO_2703 (O_2703,N_24067,N_23304);
nor UO_2704 (O_2704,N_24546,N_24819);
nor UO_2705 (O_2705,N_24849,N_23848);
nor UO_2706 (O_2706,N_23068,N_24893);
nor UO_2707 (O_2707,N_24083,N_24405);
or UO_2708 (O_2708,N_23793,N_23556);
nor UO_2709 (O_2709,N_24355,N_24144);
or UO_2710 (O_2710,N_23581,N_23368);
nor UO_2711 (O_2711,N_23993,N_23185);
nor UO_2712 (O_2712,N_23936,N_23251);
and UO_2713 (O_2713,N_24941,N_22573);
nor UO_2714 (O_2714,N_23686,N_24129);
or UO_2715 (O_2715,N_22740,N_23300);
and UO_2716 (O_2716,N_24251,N_24576);
or UO_2717 (O_2717,N_22806,N_23992);
and UO_2718 (O_2718,N_23532,N_24328);
xor UO_2719 (O_2719,N_23413,N_24962);
and UO_2720 (O_2720,N_23143,N_23139);
and UO_2721 (O_2721,N_24220,N_22704);
and UO_2722 (O_2722,N_22831,N_24444);
and UO_2723 (O_2723,N_22875,N_24392);
xnor UO_2724 (O_2724,N_23857,N_24817);
nor UO_2725 (O_2725,N_24997,N_23730);
and UO_2726 (O_2726,N_23272,N_23827);
nor UO_2727 (O_2727,N_24866,N_23699);
and UO_2728 (O_2728,N_23623,N_23011);
and UO_2729 (O_2729,N_24428,N_24278);
nor UO_2730 (O_2730,N_22715,N_23957);
nor UO_2731 (O_2731,N_23537,N_23696);
or UO_2732 (O_2732,N_24357,N_22929);
nor UO_2733 (O_2733,N_22555,N_24367);
or UO_2734 (O_2734,N_23444,N_23425);
nand UO_2735 (O_2735,N_24869,N_24347);
nand UO_2736 (O_2736,N_23173,N_24392);
xnor UO_2737 (O_2737,N_23408,N_22962);
or UO_2738 (O_2738,N_23493,N_22969);
and UO_2739 (O_2739,N_22763,N_23425);
and UO_2740 (O_2740,N_23505,N_24198);
nand UO_2741 (O_2741,N_22689,N_23257);
xor UO_2742 (O_2742,N_23207,N_24446);
and UO_2743 (O_2743,N_23359,N_23662);
or UO_2744 (O_2744,N_24995,N_24273);
nor UO_2745 (O_2745,N_22663,N_24130);
and UO_2746 (O_2746,N_23582,N_24524);
nor UO_2747 (O_2747,N_23035,N_22967);
and UO_2748 (O_2748,N_24594,N_24911);
nand UO_2749 (O_2749,N_24126,N_24528);
and UO_2750 (O_2750,N_22936,N_23204);
nor UO_2751 (O_2751,N_23190,N_22621);
or UO_2752 (O_2752,N_24911,N_22897);
nor UO_2753 (O_2753,N_24997,N_23533);
and UO_2754 (O_2754,N_23533,N_24701);
nand UO_2755 (O_2755,N_23406,N_24889);
nor UO_2756 (O_2756,N_23362,N_22516);
or UO_2757 (O_2757,N_23759,N_23767);
xor UO_2758 (O_2758,N_23114,N_22892);
and UO_2759 (O_2759,N_23781,N_24101);
xnor UO_2760 (O_2760,N_24680,N_24836);
or UO_2761 (O_2761,N_22768,N_23771);
xnor UO_2762 (O_2762,N_24139,N_23073);
nor UO_2763 (O_2763,N_23978,N_22842);
nor UO_2764 (O_2764,N_24447,N_22865);
or UO_2765 (O_2765,N_23623,N_22968);
and UO_2766 (O_2766,N_24482,N_24071);
and UO_2767 (O_2767,N_24871,N_23894);
and UO_2768 (O_2768,N_23106,N_23441);
nand UO_2769 (O_2769,N_23285,N_23944);
or UO_2770 (O_2770,N_24670,N_22782);
or UO_2771 (O_2771,N_22968,N_23873);
or UO_2772 (O_2772,N_22502,N_23174);
nand UO_2773 (O_2773,N_23447,N_22989);
and UO_2774 (O_2774,N_24515,N_24598);
nor UO_2775 (O_2775,N_24650,N_24323);
xor UO_2776 (O_2776,N_23853,N_24743);
and UO_2777 (O_2777,N_24504,N_23283);
and UO_2778 (O_2778,N_23534,N_23995);
nor UO_2779 (O_2779,N_22545,N_24416);
nand UO_2780 (O_2780,N_24431,N_24333);
or UO_2781 (O_2781,N_23550,N_24868);
nor UO_2782 (O_2782,N_23775,N_24455);
and UO_2783 (O_2783,N_24158,N_24746);
and UO_2784 (O_2784,N_24043,N_23831);
or UO_2785 (O_2785,N_24787,N_24248);
nand UO_2786 (O_2786,N_23573,N_22958);
nor UO_2787 (O_2787,N_23010,N_23003);
or UO_2788 (O_2788,N_23578,N_24635);
nand UO_2789 (O_2789,N_24966,N_23377);
xor UO_2790 (O_2790,N_24495,N_24861);
nor UO_2791 (O_2791,N_24623,N_24556);
and UO_2792 (O_2792,N_23398,N_23315);
and UO_2793 (O_2793,N_24909,N_23266);
xnor UO_2794 (O_2794,N_22998,N_23674);
xor UO_2795 (O_2795,N_23079,N_23154);
or UO_2796 (O_2796,N_23861,N_24833);
or UO_2797 (O_2797,N_23893,N_22653);
and UO_2798 (O_2798,N_23077,N_22911);
or UO_2799 (O_2799,N_24317,N_24376);
or UO_2800 (O_2800,N_23460,N_24115);
nand UO_2801 (O_2801,N_24680,N_24408);
xnor UO_2802 (O_2802,N_22763,N_22609);
nand UO_2803 (O_2803,N_24513,N_24668);
xnor UO_2804 (O_2804,N_24139,N_23071);
nand UO_2805 (O_2805,N_22609,N_23445);
and UO_2806 (O_2806,N_23018,N_22573);
nor UO_2807 (O_2807,N_22582,N_22742);
xnor UO_2808 (O_2808,N_24210,N_23832);
nand UO_2809 (O_2809,N_24059,N_24867);
nand UO_2810 (O_2810,N_24619,N_24885);
xor UO_2811 (O_2811,N_22791,N_24024);
nor UO_2812 (O_2812,N_23816,N_23194);
nor UO_2813 (O_2813,N_23087,N_24063);
nor UO_2814 (O_2814,N_23686,N_23637);
nor UO_2815 (O_2815,N_22762,N_22536);
nand UO_2816 (O_2816,N_24637,N_24249);
nand UO_2817 (O_2817,N_24867,N_23999);
nand UO_2818 (O_2818,N_24361,N_24725);
xor UO_2819 (O_2819,N_22518,N_23633);
and UO_2820 (O_2820,N_22804,N_24260);
and UO_2821 (O_2821,N_23417,N_23093);
and UO_2822 (O_2822,N_24508,N_23548);
and UO_2823 (O_2823,N_24523,N_24781);
xor UO_2824 (O_2824,N_24410,N_24431);
nor UO_2825 (O_2825,N_23795,N_24379);
nand UO_2826 (O_2826,N_23462,N_24783);
nand UO_2827 (O_2827,N_22614,N_23479);
nor UO_2828 (O_2828,N_23304,N_24811);
nor UO_2829 (O_2829,N_23374,N_22525);
and UO_2830 (O_2830,N_24908,N_24833);
or UO_2831 (O_2831,N_23859,N_24340);
or UO_2832 (O_2832,N_23059,N_24602);
or UO_2833 (O_2833,N_23347,N_23835);
xnor UO_2834 (O_2834,N_24311,N_23728);
nor UO_2835 (O_2835,N_24882,N_24699);
and UO_2836 (O_2836,N_24780,N_23167);
xnor UO_2837 (O_2837,N_23689,N_24648);
nand UO_2838 (O_2838,N_24917,N_22905);
or UO_2839 (O_2839,N_24902,N_24989);
nand UO_2840 (O_2840,N_24978,N_23532);
nor UO_2841 (O_2841,N_24107,N_24882);
and UO_2842 (O_2842,N_24242,N_24034);
nor UO_2843 (O_2843,N_23972,N_23665);
or UO_2844 (O_2844,N_24179,N_22827);
or UO_2845 (O_2845,N_22578,N_24339);
and UO_2846 (O_2846,N_23793,N_22525);
and UO_2847 (O_2847,N_24629,N_22600);
or UO_2848 (O_2848,N_24059,N_22627);
and UO_2849 (O_2849,N_24014,N_23396);
and UO_2850 (O_2850,N_24046,N_23812);
nor UO_2851 (O_2851,N_23050,N_22970);
or UO_2852 (O_2852,N_22852,N_22564);
and UO_2853 (O_2853,N_24581,N_23916);
nand UO_2854 (O_2854,N_23634,N_22751);
nor UO_2855 (O_2855,N_24708,N_22504);
nand UO_2856 (O_2856,N_24898,N_24128);
nor UO_2857 (O_2857,N_22737,N_22953);
and UO_2858 (O_2858,N_22992,N_24925);
or UO_2859 (O_2859,N_24215,N_23796);
or UO_2860 (O_2860,N_23391,N_24405);
xnor UO_2861 (O_2861,N_23332,N_22656);
xor UO_2862 (O_2862,N_24810,N_24766);
nand UO_2863 (O_2863,N_24700,N_23250);
xnor UO_2864 (O_2864,N_22519,N_23076);
nor UO_2865 (O_2865,N_24781,N_24342);
nand UO_2866 (O_2866,N_22960,N_24549);
and UO_2867 (O_2867,N_23127,N_22867);
or UO_2868 (O_2868,N_23581,N_22999);
or UO_2869 (O_2869,N_22707,N_23104);
and UO_2870 (O_2870,N_23985,N_23466);
nand UO_2871 (O_2871,N_23943,N_23575);
nor UO_2872 (O_2872,N_23104,N_24749);
nor UO_2873 (O_2873,N_23666,N_24049);
nand UO_2874 (O_2874,N_24812,N_23336);
nand UO_2875 (O_2875,N_24757,N_23829);
nor UO_2876 (O_2876,N_24376,N_22922);
nor UO_2877 (O_2877,N_23610,N_23062);
nand UO_2878 (O_2878,N_24984,N_23494);
xnor UO_2879 (O_2879,N_22796,N_23549);
xnor UO_2880 (O_2880,N_24795,N_22783);
nand UO_2881 (O_2881,N_22736,N_23003);
and UO_2882 (O_2882,N_23484,N_23923);
or UO_2883 (O_2883,N_23077,N_23248);
nor UO_2884 (O_2884,N_22756,N_24149);
nand UO_2885 (O_2885,N_22886,N_22713);
or UO_2886 (O_2886,N_24367,N_22612);
and UO_2887 (O_2887,N_24322,N_23720);
nand UO_2888 (O_2888,N_23055,N_23405);
or UO_2889 (O_2889,N_22913,N_23890);
and UO_2890 (O_2890,N_24429,N_23660);
or UO_2891 (O_2891,N_24627,N_23691);
and UO_2892 (O_2892,N_24301,N_22629);
or UO_2893 (O_2893,N_23243,N_22656);
or UO_2894 (O_2894,N_23475,N_22604);
and UO_2895 (O_2895,N_24137,N_22845);
nand UO_2896 (O_2896,N_24509,N_24895);
nor UO_2897 (O_2897,N_24418,N_23278);
and UO_2898 (O_2898,N_24579,N_24157);
nand UO_2899 (O_2899,N_23679,N_23067);
nor UO_2900 (O_2900,N_24672,N_24962);
nand UO_2901 (O_2901,N_23524,N_24358);
nand UO_2902 (O_2902,N_23093,N_22739);
and UO_2903 (O_2903,N_23321,N_23489);
and UO_2904 (O_2904,N_22728,N_23678);
nand UO_2905 (O_2905,N_23218,N_22879);
xnor UO_2906 (O_2906,N_24781,N_23162);
or UO_2907 (O_2907,N_23206,N_23006);
nor UO_2908 (O_2908,N_23851,N_23808);
nor UO_2909 (O_2909,N_24909,N_23468);
nor UO_2910 (O_2910,N_23276,N_24974);
or UO_2911 (O_2911,N_23772,N_22686);
or UO_2912 (O_2912,N_24099,N_22942);
and UO_2913 (O_2913,N_23033,N_24832);
nor UO_2914 (O_2914,N_23738,N_24466);
and UO_2915 (O_2915,N_24460,N_24971);
and UO_2916 (O_2916,N_23890,N_24107);
nor UO_2917 (O_2917,N_24040,N_23191);
nor UO_2918 (O_2918,N_22758,N_24520);
nand UO_2919 (O_2919,N_22839,N_24454);
and UO_2920 (O_2920,N_24186,N_24361);
or UO_2921 (O_2921,N_24276,N_24219);
and UO_2922 (O_2922,N_23977,N_23759);
or UO_2923 (O_2923,N_23095,N_24460);
nand UO_2924 (O_2924,N_24176,N_22812);
and UO_2925 (O_2925,N_24145,N_23904);
or UO_2926 (O_2926,N_22728,N_24640);
nor UO_2927 (O_2927,N_23927,N_23392);
nand UO_2928 (O_2928,N_24209,N_24900);
and UO_2929 (O_2929,N_23170,N_24350);
and UO_2930 (O_2930,N_22689,N_24784);
nand UO_2931 (O_2931,N_23607,N_22601);
xnor UO_2932 (O_2932,N_24940,N_23196);
nor UO_2933 (O_2933,N_23472,N_23370);
and UO_2934 (O_2934,N_23495,N_24504);
xor UO_2935 (O_2935,N_22636,N_23254);
and UO_2936 (O_2936,N_24254,N_24140);
or UO_2937 (O_2937,N_24173,N_23728);
and UO_2938 (O_2938,N_22556,N_24264);
xor UO_2939 (O_2939,N_23659,N_24340);
nand UO_2940 (O_2940,N_24452,N_22584);
nor UO_2941 (O_2941,N_24995,N_23573);
or UO_2942 (O_2942,N_23002,N_23502);
or UO_2943 (O_2943,N_22942,N_23948);
nor UO_2944 (O_2944,N_24548,N_23426);
or UO_2945 (O_2945,N_24410,N_23517);
and UO_2946 (O_2946,N_24889,N_22794);
nand UO_2947 (O_2947,N_22747,N_23700);
and UO_2948 (O_2948,N_23349,N_22533);
nand UO_2949 (O_2949,N_22853,N_23501);
nand UO_2950 (O_2950,N_24014,N_22798);
or UO_2951 (O_2951,N_23166,N_22730);
or UO_2952 (O_2952,N_23531,N_23192);
nand UO_2953 (O_2953,N_23512,N_23945);
nand UO_2954 (O_2954,N_24408,N_23576);
xnor UO_2955 (O_2955,N_23507,N_23953);
xor UO_2956 (O_2956,N_23661,N_24675);
or UO_2957 (O_2957,N_23720,N_24872);
nand UO_2958 (O_2958,N_24960,N_23251);
nand UO_2959 (O_2959,N_24830,N_24844);
and UO_2960 (O_2960,N_22508,N_24821);
xnor UO_2961 (O_2961,N_23088,N_22854);
nor UO_2962 (O_2962,N_23385,N_22909);
nand UO_2963 (O_2963,N_22567,N_23573);
xor UO_2964 (O_2964,N_24590,N_24612);
nand UO_2965 (O_2965,N_24075,N_24791);
nor UO_2966 (O_2966,N_24483,N_24668);
or UO_2967 (O_2967,N_23867,N_23706);
nor UO_2968 (O_2968,N_22733,N_24191);
nand UO_2969 (O_2969,N_23658,N_22878);
nand UO_2970 (O_2970,N_24083,N_24345);
nand UO_2971 (O_2971,N_24805,N_23646);
nand UO_2972 (O_2972,N_24901,N_22562);
xnor UO_2973 (O_2973,N_23499,N_23551);
or UO_2974 (O_2974,N_23305,N_24632);
or UO_2975 (O_2975,N_24383,N_24040);
or UO_2976 (O_2976,N_23945,N_23041);
and UO_2977 (O_2977,N_22616,N_24965);
or UO_2978 (O_2978,N_23444,N_23511);
nor UO_2979 (O_2979,N_23913,N_22887);
or UO_2980 (O_2980,N_24283,N_23351);
or UO_2981 (O_2981,N_23632,N_23605);
or UO_2982 (O_2982,N_24537,N_22720);
xnor UO_2983 (O_2983,N_24676,N_24334);
nor UO_2984 (O_2984,N_22725,N_24701);
and UO_2985 (O_2985,N_23287,N_23842);
or UO_2986 (O_2986,N_23670,N_23530);
nand UO_2987 (O_2987,N_22825,N_23746);
and UO_2988 (O_2988,N_23489,N_24116);
nor UO_2989 (O_2989,N_22815,N_24339);
and UO_2990 (O_2990,N_24169,N_24794);
or UO_2991 (O_2991,N_22657,N_23969);
nand UO_2992 (O_2992,N_23775,N_23875);
nor UO_2993 (O_2993,N_23228,N_22917);
nor UO_2994 (O_2994,N_22717,N_24173);
nor UO_2995 (O_2995,N_23144,N_23854);
nand UO_2996 (O_2996,N_24830,N_23574);
or UO_2997 (O_2997,N_23889,N_22549);
and UO_2998 (O_2998,N_24701,N_22506);
and UO_2999 (O_2999,N_24823,N_24965);
endmodule