module basic_1000_10000_1500_10_levels_2xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
and U0 (N_0,In_110,In_233);
nand U1 (N_1,In_886,In_977);
nand U2 (N_2,In_789,In_706);
and U3 (N_3,In_83,In_989);
nor U4 (N_4,In_826,In_30);
nand U5 (N_5,In_304,In_61);
or U6 (N_6,In_950,In_218);
xnor U7 (N_7,In_139,In_740);
and U8 (N_8,In_857,In_987);
nand U9 (N_9,In_253,In_902);
xnor U10 (N_10,In_667,In_644);
nor U11 (N_11,In_479,In_847);
or U12 (N_12,In_311,In_585);
or U13 (N_13,In_582,In_124);
and U14 (N_14,In_484,In_143);
nand U15 (N_15,In_406,In_806);
nand U16 (N_16,In_637,In_410);
and U17 (N_17,In_382,In_100);
nor U18 (N_18,In_547,In_595);
nor U19 (N_19,In_846,In_424);
and U20 (N_20,In_549,In_899);
nor U21 (N_21,In_421,In_995);
xnor U22 (N_22,In_542,In_467);
and U23 (N_23,In_300,In_296);
nor U24 (N_24,In_701,In_809);
and U25 (N_25,In_29,In_960);
or U26 (N_26,In_272,In_281);
nor U27 (N_27,In_142,In_873);
nand U28 (N_28,In_648,In_640);
or U29 (N_29,In_224,In_279);
or U30 (N_30,In_691,In_622);
and U31 (N_31,In_752,In_793);
nand U32 (N_32,In_299,In_22);
or U33 (N_33,In_580,In_610);
nor U34 (N_34,In_444,In_791);
and U35 (N_35,In_92,In_502);
or U36 (N_36,In_699,In_482);
nand U37 (N_37,In_919,In_732);
nor U38 (N_38,In_134,In_438);
nor U39 (N_39,In_18,In_744);
nand U40 (N_40,In_745,In_932);
nor U41 (N_41,In_356,In_604);
nor U42 (N_42,In_660,In_653);
nand U43 (N_43,In_680,In_230);
or U44 (N_44,In_36,In_958);
nor U45 (N_45,In_551,In_11);
and U46 (N_46,In_850,In_41);
nor U47 (N_47,In_803,In_761);
nor U48 (N_48,In_844,In_123);
nand U49 (N_49,In_27,In_239);
nor U50 (N_50,In_469,In_900);
nand U51 (N_51,In_824,In_676);
nor U52 (N_52,In_603,In_627);
nor U53 (N_53,In_816,In_992);
nor U54 (N_54,In_657,In_565);
nor U55 (N_55,In_292,In_7);
and U56 (N_56,In_297,In_853);
nor U57 (N_57,In_669,In_500);
nor U58 (N_58,In_372,In_387);
or U59 (N_59,In_215,In_998);
and U60 (N_60,In_418,In_859);
nor U61 (N_61,In_544,In_133);
nand U62 (N_62,In_925,In_481);
nand U63 (N_63,In_156,In_489);
xnor U64 (N_64,In_914,In_33);
nor U65 (N_65,In_154,In_738);
and U66 (N_66,In_875,In_68);
or U67 (N_67,In_843,In_115);
nor U68 (N_68,In_711,In_633);
xnor U69 (N_69,In_270,In_125);
nand U70 (N_70,In_739,In_363);
nor U71 (N_71,In_755,In_804);
and U72 (N_72,In_629,In_635);
nand U73 (N_73,In_194,In_876);
or U74 (N_74,In_910,In_709);
or U75 (N_75,In_399,In_463);
xor U76 (N_76,In_885,In_474);
nand U77 (N_77,In_666,In_232);
or U78 (N_78,In_248,In_345);
nor U79 (N_79,In_184,In_211);
nand U80 (N_80,In_338,In_54);
nor U81 (N_81,In_283,In_548);
and U82 (N_82,In_874,In_815);
and U83 (N_83,In_730,In_274);
nor U84 (N_84,In_763,In_390);
or U85 (N_85,In_955,In_371);
and U86 (N_86,In_389,In_97);
nor U87 (N_87,In_331,In_636);
and U88 (N_88,In_678,In_999);
or U89 (N_89,In_89,In_715);
nand U90 (N_90,In_727,In_433);
nand U91 (N_91,In_312,In_831);
nand U92 (N_92,In_820,In_122);
nor U93 (N_93,In_349,In_956);
xnor U94 (N_94,In_81,In_466);
nor U95 (N_95,In_188,In_499);
nand U96 (N_96,In_206,In_975);
nor U97 (N_97,In_392,In_289);
and U98 (N_98,In_788,In_722);
or U99 (N_99,In_119,In_609);
or U100 (N_100,In_12,In_976);
and U101 (N_101,In_405,In_725);
and U102 (N_102,In_265,In_77);
nand U103 (N_103,In_923,In_769);
nand U104 (N_104,In_756,In_225);
xnor U105 (N_105,In_367,In_385);
nor U106 (N_106,In_323,In_497);
nor U107 (N_107,In_94,In_429);
and U108 (N_108,In_533,In_452);
nand U109 (N_109,In_777,In_796);
or U110 (N_110,In_584,In_887);
and U111 (N_111,In_483,In_415);
or U112 (N_112,In_797,In_167);
nand U113 (N_113,In_959,In_103);
nand U114 (N_114,In_984,In_116);
or U115 (N_115,In_736,In_85);
nor U116 (N_116,In_447,In_186);
nand U117 (N_117,In_654,In_197);
nor U118 (N_118,In_927,In_287);
or U119 (N_119,In_618,In_73);
or U120 (N_120,In_832,In_377);
nand U121 (N_121,In_164,In_579);
or U122 (N_122,In_471,In_827);
and U123 (N_123,In_835,In_778);
nand U124 (N_124,In_511,In_343);
nor U125 (N_125,In_196,In_384);
and U126 (N_126,In_612,In_868);
nand U127 (N_127,In_978,In_180);
nor U128 (N_128,In_712,In_91);
and U129 (N_129,In_598,In_16);
or U130 (N_130,In_535,In_808);
or U131 (N_131,In_737,In_829);
nand U132 (N_132,In_504,In_628);
nor U133 (N_133,In_605,In_344);
nand U134 (N_134,In_314,In_370);
or U135 (N_135,In_681,In_907);
nand U136 (N_136,In_404,In_921);
nor U137 (N_137,In_468,In_563);
nor U138 (N_138,In_257,In_420);
nand U139 (N_139,In_781,In_46);
or U140 (N_140,In_207,In_288);
and U141 (N_141,In_554,In_718);
nor U142 (N_142,In_785,In_767);
and U143 (N_143,In_822,In_509);
nor U144 (N_144,In_555,In_255);
nand U145 (N_145,In_567,In_790);
and U146 (N_146,In_645,In_607);
nor U147 (N_147,In_90,In_357);
or U148 (N_148,In_674,In_571);
or U149 (N_149,In_0,In_425);
nor U150 (N_150,In_498,In_606);
nor U151 (N_151,In_710,In_491);
or U152 (N_152,In_21,In_105);
or U153 (N_153,In_332,In_47);
and U154 (N_154,In_79,In_780);
nor U155 (N_155,In_505,In_231);
nand U156 (N_156,In_946,In_56);
nand U157 (N_157,In_677,In_953);
nor U158 (N_158,In_825,In_634);
or U159 (N_159,In_38,In_558);
nand U160 (N_160,In_583,In_132);
nor U161 (N_161,In_456,In_707);
nand U162 (N_162,In_774,In_772);
nand U163 (N_163,In_979,In_307);
nand U164 (N_164,In_168,In_684);
nor U165 (N_165,In_540,In_52);
and U166 (N_166,In_541,In_714);
nand U167 (N_167,In_728,In_63);
nand U168 (N_168,In_347,In_457);
or U169 (N_169,In_86,In_409);
and U170 (N_170,In_890,In_852);
and U171 (N_171,In_668,In_416);
and U172 (N_172,In_526,In_348);
and U173 (N_173,In_798,In_490);
xnor U174 (N_174,In_198,In_459);
nor U175 (N_175,In_717,In_938);
or U176 (N_176,In_6,In_673);
nand U177 (N_177,In_762,In_319);
nand U178 (N_178,In_974,In_379);
nor U179 (N_179,In_126,In_195);
nor U180 (N_180,In_775,In_432);
nand U181 (N_181,In_833,In_219);
and U182 (N_182,In_109,In_599);
nor U183 (N_183,In_10,In_203);
and U184 (N_184,In_812,In_325);
nand U185 (N_185,In_861,In_517);
nand U186 (N_186,In_104,In_414);
nor U187 (N_187,In_911,In_906);
nor U188 (N_188,In_49,In_366);
and U189 (N_189,In_939,In_501);
nand U190 (N_190,In_318,In_93);
and U191 (N_191,In_151,In_179);
nand U192 (N_192,In_1,In_903);
nor U193 (N_193,In_894,In_795);
nor U194 (N_194,In_532,In_621);
and U195 (N_195,In_746,In_968);
and U196 (N_196,In_631,In_700);
and U197 (N_197,In_695,In_776);
xnor U198 (N_198,In_2,In_40);
and U199 (N_199,In_687,In_726);
nand U200 (N_200,In_748,In_315);
or U201 (N_201,In_342,In_64);
and U202 (N_202,In_940,In_856);
and U203 (N_203,In_295,In_329);
nand U204 (N_204,In_448,In_661);
nand U205 (N_205,In_639,In_965);
and U206 (N_206,In_792,In_649);
nand U207 (N_207,In_200,In_750);
or U208 (N_208,In_155,In_993);
nor U209 (N_209,In_920,In_496);
nand U210 (N_210,In_174,In_908);
and U211 (N_211,In_23,In_84);
or U212 (N_212,In_191,In_252);
and U213 (N_213,In_39,In_422);
or U214 (N_214,In_221,In_146);
nand U215 (N_215,In_82,In_836);
and U216 (N_216,In_536,In_729);
or U217 (N_217,In_241,In_513);
nand U218 (N_218,In_177,In_690);
and U219 (N_219,In_952,In_638);
and U220 (N_220,In_381,In_487);
and U221 (N_221,In_401,In_204);
or U222 (N_222,In_80,In_596);
or U223 (N_223,In_277,In_572);
or U224 (N_224,In_340,In_413);
xor U225 (N_225,In_461,In_361);
nor U226 (N_226,In_757,In_136);
nor U227 (N_227,In_869,In_698);
and U228 (N_228,In_396,In_658);
and U229 (N_229,In_284,In_165);
or U230 (N_230,In_983,In_538);
or U231 (N_231,In_884,In_310);
or U232 (N_232,In_864,In_298);
and U233 (N_233,In_516,In_402);
nor U234 (N_234,In_904,In_145);
nor U235 (N_235,In_346,In_753);
or U236 (N_236,In_170,In_916);
nor U237 (N_237,In_670,In_427);
xor U238 (N_238,In_320,In_368);
and U239 (N_239,In_839,In_764);
or U240 (N_240,In_408,In_59);
and U241 (N_241,In_877,In_326);
nor U242 (N_242,In_129,In_20);
nor U243 (N_243,In_564,In_364);
or U244 (N_244,In_672,In_291);
or U245 (N_245,In_375,In_849);
or U246 (N_246,In_840,In_25);
or U247 (N_247,In_182,In_493);
nor U248 (N_248,In_321,In_895);
nor U249 (N_249,In_131,In_193);
or U250 (N_250,In_759,In_988);
nand U251 (N_251,In_924,In_365);
nand U252 (N_252,In_261,In_862);
nand U253 (N_253,In_28,In_529);
nand U254 (N_254,In_592,In_458);
nor U255 (N_255,In_515,In_854);
and U256 (N_256,In_477,In_293);
and U257 (N_257,In_480,In_111);
or U258 (N_258,In_334,In_148);
and U259 (N_259,In_937,In_227);
nor U260 (N_260,In_178,In_303);
nor U261 (N_261,In_117,In_512);
nor U262 (N_262,In_465,In_439);
and U263 (N_263,In_751,In_37);
nor U264 (N_264,In_341,In_216);
nand U265 (N_265,In_138,In_845);
nor U266 (N_266,In_613,In_786);
and U267 (N_267,In_66,In_214);
nor U268 (N_268,In_814,In_970);
and U269 (N_269,In_434,In_19);
nand U270 (N_270,In_525,In_358);
nand U271 (N_271,In_158,In_285);
or U272 (N_272,In_436,In_118);
and U273 (N_273,In_766,In_758);
and U274 (N_274,In_144,In_238);
nor U275 (N_275,In_235,In_819);
xor U276 (N_276,In_441,In_980);
xnor U277 (N_277,In_226,In_561);
and U278 (N_278,In_395,In_537);
or U279 (N_279,In_127,In_619);
or U280 (N_280,In_588,In_768);
nand U281 (N_281,In_830,In_309);
nor U282 (N_282,In_659,In_704);
and U283 (N_283,In_55,In_616);
or U284 (N_284,In_963,In_624);
or U285 (N_285,In_445,In_724);
or U286 (N_286,In_275,In_747);
and U287 (N_287,In_817,In_552);
and U288 (N_288,In_282,In_705);
and U289 (N_289,In_205,In_973);
nand U290 (N_290,In_962,In_679);
or U291 (N_291,In_794,In_945);
or U292 (N_292,In_573,In_212);
nand U293 (N_293,In_647,In_721);
nor U294 (N_294,In_453,In_286);
or U295 (N_295,In_883,In_581);
nor U296 (N_296,In_575,In_696);
nand U297 (N_297,In_615,In_734);
nand U298 (N_298,In_742,In_770);
nand U299 (N_299,In_848,In_256);
nor U300 (N_300,In_985,In_694);
nor U301 (N_301,In_400,In_333);
nor U302 (N_302,In_799,In_169);
and U303 (N_303,In_929,In_546);
and U304 (N_304,In_578,In_183);
or U305 (N_305,In_175,In_316);
and U306 (N_306,In_140,In_69);
nand U307 (N_307,In_866,In_842);
and U308 (N_308,In_943,In_574);
nor U309 (N_309,In_642,In_171);
and U310 (N_310,In_917,In_878);
or U311 (N_311,In_271,In_449);
nand U312 (N_312,In_419,In_841);
nand U313 (N_313,In_78,In_201);
nor U314 (N_314,In_190,In_528);
or U315 (N_315,In_250,In_863);
nand U316 (N_316,In_813,In_508);
nand U317 (N_317,In_760,In_4);
and U318 (N_318,In_435,In_527);
and U319 (N_319,In_787,In_128);
nand U320 (N_320,In_407,In_101);
nor U321 (N_321,In_893,In_855);
and U322 (N_322,In_373,In_397);
nor U323 (N_323,In_51,In_783);
nand U324 (N_324,In_683,In_234);
or U325 (N_325,In_663,In_643);
nand U326 (N_326,In_388,In_62);
or U327 (N_327,In_150,In_543);
or U328 (N_328,In_662,In_782);
nand U329 (N_329,In_327,In_15);
nor U330 (N_330,In_313,In_460);
and U331 (N_331,In_702,In_244);
nand U332 (N_332,In_703,In_870);
nor U333 (N_333,In_823,In_997);
or U334 (N_334,In_113,In_773);
nor U335 (N_335,In_222,In_942);
or U336 (N_336,In_267,In_858);
nor U337 (N_337,In_393,In_928);
nand U338 (N_338,In_593,In_488);
xnor U339 (N_339,In_217,In_591);
nand U340 (N_340,In_996,In_446);
and U341 (N_341,In_251,In_269);
or U342 (N_342,In_254,In_971);
nand U343 (N_343,In_811,In_454);
nand U344 (N_344,In_189,In_765);
nand U345 (N_345,In_48,In_994);
or U346 (N_346,In_913,In_273);
or U347 (N_347,In_733,In_898);
xor U348 (N_348,In_278,In_521);
nand U349 (N_349,In_986,In_24);
nor U350 (N_350,In_523,In_476);
xor U351 (N_351,In_95,In_8);
or U352 (N_352,In_602,In_147);
nor U353 (N_353,In_577,In_322);
or U354 (N_354,In_731,In_9);
and U355 (N_355,In_43,In_594);
nand U356 (N_356,In_623,In_26);
nor U357 (N_357,In_249,In_743);
nor U358 (N_358,In_518,In_403);
nand U359 (N_359,In_881,In_213);
nand U360 (N_360,In_779,In_130);
nor U361 (N_361,In_236,In_172);
and U362 (N_362,In_964,In_784);
and U363 (N_363,In_185,In_398);
nand U364 (N_364,In_949,In_539);
nor U365 (N_365,In_411,In_242);
or U366 (N_366,In_106,In_837);
and U367 (N_367,In_632,In_324);
or U368 (N_368,In_626,In_259);
xnor U369 (N_369,In_961,In_867);
and U370 (N_370,In_306,In_557);
or U371 (N_371,In_354,In_896);
xor U372 (N_372,In_374,In_569);
nor U373 (N_373,In_376,In_470);
nor U374 (N_374,In_208,In_838);
and U375 (N_375,In_161,In_74);
nand U376 (N_376,In_423,In_590);
nand U377 (N_377,In_350,In_245);
or U378 (N_378,In_162,In_263);
or U379 (N_379,In_934,In_247);
nand U380 (N_380,In_982,In_944);
or U381 (N_381,In_220,In_915);
nand U382 (N_382,In_646,In_114);
nand U383 (N_383,In_262,In_163);
nor U384 (N_384,In_121,In_60);
and U385 (N_385,In_486,In_192);
or U386 (N_386,In_229,In_909);
nor U387 (N_387,In_545,In_957);
and U388 (N_388,In_948,In_50);
or U389 (N_389,In_264,In_67);
and U390 (N_390,In_102,In_889);
or U391 (N_391,In_720,In_112);
or U392 (N_392,In_369,In_352);
and U393 (N_393,In_160,In_872);
nand U394 (N_394,In_735,In_380);
and U395 (N_395,In_930,In_947);
nor U396 (N_396,In_280,In_522);
nand U397 (N_397,In_3,In_276);
and U398 (N_398,In_473,In_290);
and U399 (N_399,In_918,In_96);
xnor U400 (N_400,In_157,In_566);
and U401 (N_401,In_597,In_936);
or U402 (N_402,In_912,In_437);
and U403 (N_403,In_802,In_353);
or U404 (N_404,In_689,In_951);
and U405 (N_405,In_879,In_990);
nor U406 (N_406,In_559,In_317);
xor U407 (N_407,In_34,In_87);
or U408 (N_408,In_335,In_954);
or U409 (N_409,In_258,In_754);
nand U410 (N_410,In_412,In_905);
nor U411 (N_411,In_800,In_351);
or U412 (N_412,In_475,In_865);
or U413 (N_413,In_58,In_671);
and U414 (N_414,In_600,In_485);
or U415 (N_415,In_818,In_828);
or U416 (N_416,In_44,In_805);
nor U417 (N_417,In_339,In_697);
nand U418 (N_418,In_601,In_933);
nand U419 (N_419,In_243,In_708);
and U420 (N_420,In_266,In_664);
or U421 (N_421,In_553,In_931);
and U422 (N_422,In_260,In_495);
and U423 (N_423,In_141,In_336);
and U424 (N_424,In_440,In_72);
or U425 (N_425,In_228,In_35);
or U426 (N_426,In_31,In_337);
and U427 (N_427,In_159,In_152);
and U428 (N_428,In_99,In_570);
nand U429 (N_429,In_506,In_614);
and U430 (N_430,In_472,In_688);
nand U431 (N_431,In_65,In_246);
nor U432 (N_432,In_430,In_514);
nor U433 (N_433,In_187,In_935);
nand U434 (N_434,In_88,In_359);
nor U435 (N_435,In_534,In_135);
nor U436 (N_436,In_149,In_586);
and U437 (N_437,In_807,In_560);
nor U438 (N_438,In_305,In_901);
or U439 (N_439,In_362,In_378);
nand U440 (N_440,In_576,In_589);
nand U441 (N_441,In_665,In_871);
or U442 (N_442,In_308,In_442);
or U443 (N_443,In_655,In_383);
xnor U444 (N_444,In_492,In_443);
and U445 (N_445,In_969,In_107);
or U446 (N_446,In_428,In_237);
or U447 (N_447,In_75,In_426);
nand U448 (N_448,In_991,In_749);
nor U449 (N_449,In_202,In_294);
or U450 (N_450,In_520,In_568);
and U451 (N_451,In_166,In_651);
nor U452 (N_452,In_455,In_98);
or U453 (N_453,In_153,In_210);
nor U454 (N_454,In_608,In_531);
nand U455 (N_455,In_181,In_692);
or U456 (N_456,In_32,In_223);
nand U457 (N_457,In_686,In_972);
nor U458 (N_458,In_834,In_926);
or U459 (N_459,In_981,In_630);
nor U460 (N_460,In_611,In_45);
nand U461 (N_461,In_556,In_53);
or U462 (N_462,In_302,In_120);
nor U463 (N_463,In_967,In_391);
and U464 (N_464,In_650,In_330);
xor U465 (N_465,In_360,In_587);
or U466 (N_466,In_71,In_713);
xor U467 (N_467,In_268,In_394);
and U468 (N_468,In_510,In_462);
or U469 (N_469,In_891,In_14);
and U470 (N_470,In_386,In_656);
nand U471 (N_471,In_693,In_620);
or U472 (N_472,In_652,In_880);
or U473 (N_473,In_42,In_451);
or U474 (N_474,In_301,In_450);
or U475 (N_475,In_892,In_966);
nor U476 (N_476,In_550,In_897);
and U477 (N_477,In_173,In_17);
and U478 (N_478,In_617,In_240);
nand U479 (N_479,In_771,In_723);
nor U480 (N_480,In_882,In_821);
xnor U481 (N_481,In_328,In_716);
and U482 (N_482,In_922,In_494);
nand U483 (N_483,In_625,In_685);
and U484 (N_484,In_137,In_5);
and U485 (N_485,In_503,In_810);
and U486 (N_486,In_675,In_682);
and U487 (N_487,In_741,In_199);
nand U488 (N_488,In_801,In_851);
nor U489 (N_489,In_464,In_562);
or U490 (N_490,In_860,In_13);
or U491 (N_491,In_530,In_888);
and U492 (N_492,In_76,In_478);
or U493 (N_493,In_70,In_355);
or U494 (N_494,In_941,In_417);
or U495 (N_495,In_431,In_641);
nand U496 (N_496,In_524,In_176);
or U497 (N_497,In_57,In_507);
and U498 (N_498,In_719,In_519);
nand U499 (N_499,In_108,In_209);
and U500 (N_500,In_163,In_683);
nor U501 (N_501,In_482,In_421);
nand U502 (N_502,In_754,In_958);
or U503 (N_503,In_407,In_29);
or U504 (N_504,In_284,In_861);
nand U505 (N_505,In_369,In_313);
nor U506 (N_506,In_318,In_419);
nor U507 (N_507,In_6,In_93);
or U508 (N_508,In_451,In_599);
nor U509 (N_509,In_31,In_814);
nand U510 (N_510,In_77,In_351);
xnor U511 (N_511,In_574,In_502);
and U512 (N_512,In_356,In_185);
nor U513 (N_513,In_298,In_511);
nand U514 (N_514,In_875,In_762);
and U515 (N_515,In_728,In_24);
and U516 (N_516,In_940,In_800);
nor U517 (N_517,In_992,In_832);
or U518 (N_518,In_611,In_853);
nor U519 (N_519,In_977,In_368);
nand U520 (N_520,In_953,In_143);
nor U521 (N_521,In_208,In_47);
and U522 (N_522,In_686,In_266);
nor U523 (N_523,In_230,In_811);
nor U524 (N_524,In_920,In_424);
nor U525 (N_525,In_900,In_965);
and U526 (N_526,In_192,In_496);
nand U527 (N_527,In_59,In_898);
nand U528 (N_528,In_365,In_692);
and U529 (N_529,In_707,In_414);
or U530 (N_530,In_490,In_434);
xor U531 (N_531,In_149,In_579);
nor U532 (N_532,In_632,In_312);
and U533 (N_533,In_332,In_935);
nand U534 (N_534,In_278,In_970);
or U535 (N_535,In_430,In_338);
nor U536 (N_536,In_317,In_260);
nor U537 (N_537,In_760,In_32);
nand U538 (N_538,In_98,In_58);
nand U539 (N_539,In_941,In_704);
nand U540 (N_540,In_269,In_312);
nand U541 (N_541,In_99,In_59);
nand U542 (N_542,In_364,In_515);
and U543 (N_543,In_309,In_386);
or U544 (N_544,In_81,In_698);
and U545 (N_545,In_509,In_986);
nand U546 (N_546,In_501,In_735);
and U547 (N_547,In_546,In_364);
and U548 (N_548,In_827,In_478);
nand U549 (N_549,In_782,In_814);
and U550 (N_550,In_288,In_362);
nor U551 (N_551,In_199,In_312);
xnor U552 (N_552,In_261,In_489);
nand U553 (N_553,In_62,In_830);
nor U554 (N_554,In_562,In_322);
and U555 (N_555,In_576,In_365);
nand U556 (N_556,In_297,In_601);
nand U557 (N_557,In_194,In_355);
nand U558 (N_558,In_952,In_81);
nand U559 (N_559,In_938,In_975);
nor U560 (N_560,In_601,In_36);
and U561 (N_561,In_508,In_867);
or U562 (N_562,In_23,In_340);
and U563 (N_563,In_953,In_386);
nand U564 (N_564,In_521,In_57);
or U565 (N_565,In_405,In_506);
nor U566 (N_566,In_83,In_393);
or U567 (N_567,In_6,In_371);
nor U568 (N_568,In_734,In_353);
xor U569 (N_569,In_215,In_944);
nand U570 (N_570,In_535,In_349);
nand U571 (N_571,In_711,In_665);
and U572 (N_572,In_21,In_446);
nor U573 (N_573,In_757,In_942);
nand U574 (N_574,In_3,In_214);
nand U575 (N_575,In_921,In_991);
and U576 (N_576,In_359,In_142);
xnor U577 (N_577,In_255,In_708);
and U578 (N_578,In_583,In_540);
and U579 (N_579,In_606,In_541);
nand U580 (N_580,In_164,In_94);
nor U581 (N_581,In_724,In_316);
nand U582 (N_582,In_299,In_668);
or U583 (N_583,In_687,In_954);
or U584 (N_584,In_166,In_755);
nand U585 (N_585,In_738,In_250);
or U586 (N_586,In_191,In_838);
and U587 (N_587,In_527,In_873);
or U588 (N_588,In_105,In_545);
nand U589 (N_589,In_546,In_493);
nor U590 (N_590,In_520,In_307);
and U591 (N_591,In_659,In_915);
nand U592 (N_592,In_137,In_779);
and U593 (N_593,In_686,In_238);
and U594 (N_594,In_310,In_604);
and U595 (N_595,In_297,In_785);
or U596 (N_596,In_208,In_79);
and U597 (N_597,In_268,In_891);
nor U598 (N_598,In_762,In_979);
nand U599 (N_599,In_358,In_427);
and U600 (N_600,In_580,In_345);
or U601 (N_601,In_815,In_353);
and U602 (N_602,In_980,In_954);
and U603 (N_603,In_791,In_239);
or U604 (N_604,In_661,In_982);
or U605 (N_605,In_713,In_905);
and U606 (N_606,In_342,In_712);
and U607 (N_607,In_636,In_259);
nor U608 (N_608,In_90,In_382);
nor U609 (N_609,In_331,In_224);
and U610 (N_610,In_161,In_773);
nor U611 (N_611,In_50,In_831);
nand U612 (N_612,In_857,In_348);
nor U613 (N_613,In_480,In_819);
nand U614 (N_614,In_177,In_779);
and U615 (N_615,In_607,In_989);
nand U616 (N_616,In_407,In_353);
nand U617 (N_617,In_555,In_635);
and U618 (N_618,In_191,In_463);
and U619 (N_619,In_280,In_829);
xnor U620 (N_620,In_963,In_162);
and U621 (N_621,In_128,In_617);
or U622 (N_622,In_518,In_189);
xnor U623 (N_623,In_892,In_345);
nor U624 (N_624,In_597,In_225);
nor U625 (N_625,In_626,In_609);
nor U626 (N_626,In_194,In_536);
nor U627 (N_627,In_165,In_845);
nor U628 (N_628,In_823,In_814);
nand U629 (N_629,In_205,In_87);
or U630 (N_630,In_712,In_858);
nand U631 (N_631,In_121,In_763);
or U632 (N_632,In_550,In_996);
or U633 (N_633,In_93,In_887);
or U634 (N_634,In_963,In_432);
and U635 (N_635,In_329,In_858);
nor U636 (N_636,In_341,In_447);
nor U637 (N_637,In_941,In_246);
and U638 (N_638,In_838,In_179);
or U639 (N_639,In_396,In_620);
nor U640 (N_640,In_544,In_317);
or U641 (N_641,In_392,In_849);
nand U642 (N_642,In_832,In_116);
nor U643 (N_643,In_294,In_227);
or U644 (N_644,In_593,In_133);
nor U645 (N_645,In_900,In_939);
nor U646 (N_646,In_71,In_34);
nand U647 (N_647,In_900,In_711);
or U648 (N_648,In_831,In_90);
nor U649 (N_649,In_934,In_396);
and U650 (N_650,In_310,In_490);
nor U651 (N_651,In_81,In_192);
or U652 (N_652,In_899,In_418);
nand U653 (N_653,In_641,In_629);
nand U654 (N_654,In_326,In_733);
nand U655 (N_655,In_346,In_549);
xnor U656 (N_656,In_807,In_537);
and U657 (N_657,In_273,In_509);
nand U658 (N_658,In_85,In_140);
and U659 (N_659,In_218,In_14);
or U660 (N_660,In_770,In_189);
nor U661 (N_661,In_446,In_483);
nand U662 (N_662,In_527,In_124);
or U663 (N_663,In_935,In_266);
or U664 (N_664,In_644,In_420);
nand U665 (N_665,In_32,In_605);
and U666 (N_666,In_43,In_693);
or U667 (N_667,In_763,In_63);
nand U668 (N_668,In_318,In_883);
nand U669 (N_669,In_794,In_847);
xor U670 (N_670,In_942,In_654);
nor U671 (N_671,In_665,In_16);
and U672 (N_672,In_319,In_543);
nand U673 (N_673,In_204,In_600);
nand U674 (N_674,In_418,In_683);
nand U675 (N_675,In_432,In_416);
and U676 (N_676,In_717,In_594);
nand U677 (N_677,In_890,In_469);
nand U678 (N_678,In_366,In_668);
and U679 (N_679,In_21,In_138);
or U680 (N_680,In_808,In_943);
nor U681 (N_681,In_935,In_545);
and U682 (N_682,In_462,In_883);
and U683 (N_683,In_172,In_857);
nor U684 (N_684,In_700,In_572);
or U685 (N_685,In_389,In_830);
or U686 (N_686,In_207,In_216);
and U687 (N_687,In_180,In_16);
or U688 (N_688,In_657,In_636);
or U689 (N_689,In_650,In_501);
and U690 (N_690,In_546,In_78);
nor U691 (N_691,In_697,In_964);
nor U692 (N_692,In_797,In_445);
nor U693 (N_693,In_2,In_126);
nor U694 (N_694,In_337,In_123);
or U695 (N_695,In_877,In_132);
xnor U696 (N_696,In_453,In_865);
or U697 (N_697,In_911,In_552);
nor U698 (N_698,In_537,In_170);
and U699 (N_699,In_115,In_902);
and U700 (N_700,In_231,In_23);
or U701 (N_701,In_21,In_659);
and U702 (N_702,In_436,In_715);
nor U703 (N_703,In_118,In_447);
and U704 (N_704,In_985,In_678);
nor U705 (N_705,In_259,In_378);
nor U706 (N_706,In_357,In_234);
nand U707 (N_707,In_383,In_607);
xor U708 (N_708,In_496,In_257);
nand U709 (N_709,In_939,In_265);
nand U710 (N_710,In_111,In_948);
nand U711 (N_711,In_337,In_536);
nor U712 (N_712,In_129,In_21);
nor U713 (N_713,In_946,In_631);
nor U714 (N_714,In_94,In_827);
nand U715 (N_715,In_667,In_57);
or U716 (N_716,In_872,In_561);
or U717 (N_717,In_981,In_255);
and U718 (N_718,In_267,In_642);
nand U719 (N_719,In_821,In_37);
nand U720 (N_720,In_122,In_769);
or U721 (N_721,In_72,In_456);
nand U722 (N_722,In_322,In_236);
nor U723 (N_723,In_303,In_73);
xnor U724 (N_724,In_962,In_935);
nand U725 (N_725,In_127,In_228);
nand U726 (N_726,In_156,In_305);
nor U727 (N_727,In_384,In_442);
and U728 (N_728,In_980,In_426);
nor U729 (N_729,In_437,In_712);
or U730 (N_730,In_138,In_178);
nand U731 (N_731,In_111,In_411);
nor U732 (N_732,In_701,In_254);
or U733 (N_733,In_932,In_893);
xnor U734 (N_734,In_840,In_369);
nand U735 (N_735,In_884,In_584);
nand U736 (N_736,In_467,In_398);
or U737 (N_737,In_212,In_252);
nand U738 (N_738,In_835,In_512);
or U739 (N_739,In_492,In_688);
xor U740 (N_740,In_426,In_759);
nor U741 (N_741,In_825,In_773);
nor U742 (N_742,In_365,In_189);
nand U743 (N_743,In_69,In_249);
nor U744 (N_744,In_774,In_211);
nand U745 (N_745,In_895,In_891);
and U746 (N_746,In_42,In_867);
nand U747 (N_747,In_639,In_540);
and U748 (N_748,In_11,In_948);
or U749 (N_749,In_53,In_753);
nand U750 (N_750,In_215,In_200);
nor U751 (N_751,In_552,In_766);
nand U752 (N_752,In_158,In_799);
and U753 (N_753,In_655,In_527);
and U754 (N_754,In_730,In_627);
nand U755 (N_755,In_567,In_888);
or U756 (N_756,In_517,In_399);
or U757 (N_757,In_244,In_768);
nand U758 (N_758,In_653,In_348);
nand U759 (N_759,In_630,In_862);
or U760 (N_760,In_186,In_25);
nand U761 (N_761,In_348,In_915);
and U762 (N_762,In_89,In_718);
nor U763 (N_763,In_842,In_264);
and U764 (N_764,In_159,In_226);
xor U765 (N_765,In_55,In_582);
nor U766 (N_766,In_681,In_441);
and U767 (N_767,In_79,In_771);
nand U768 (N_768,In_293,In_143);
nand U769 (N_769,In_773,In_418);
and U770 (N_770,In_314,In_890);
and U771 (N_771,In_15,In_222);
and U772 (N_772,In_818,In_330);
nand U773 (N_773,In_949,In_799);
nand U774 (N_774,In_870,In_641);
nor U775 (N_775,In_273,In_45);
or U776 (N_776,In_229,In_613);
nor U777 (N_777,In_154,In_606);
nand U778 (N_778,In_217,In_696);
xnor U779 (N_779,In_292,In_542);
or U780 (N_780,In_86,In_22);
and U781 (N_781,In_469,In_775);
nand U782 (N_782,In_113,In_941);
nand U783 (N_783,In_804,In_629);
nand U784 (N_784,In_288,In_212);
nor U785 (N_785,In_200,In_473);
nor U786 (N_786,In_107,In_198);
nand U787 (N_787,In_953,In_765);
nand U788 (N_788,In_354,In_439);
nor U789 (N_789,In_77,In_654);
nor U790 (N_790,In_198,In_676);
nand U791 (N_791,In_879,In_631);
and U792 (N_792,In_989,In_640);
and U793 (N_793,In_304,In_695);
or U794 (N_794,In_964,In_693);
nor U795 (N_795,In_787,In_320);
nand U796 (N_796,In_278,In_541);
nor U797 (N_797,In_5,In_981);
nor U798 (N_798,In_763,In_359);
nor U799 (N_799,In_58,In_268);
and U800 (N_800,In_476,In_251);
nor U801 (N_801,In_605,In_921);
nor U802 (N_802,In_625,In_387);
and U803 (N_803,In_949,In_697);
and U804 (N_804,In_124,In_326);
nand U805 (N_805,In_191,In_44);
nor U806 (N_806,In_234,In_324);
nand U807 (N_807,In_221,In_91);
nor U808 (N_808,In_573,In_576);
and U809 (N_809,In_624,In_967);
nand U810 (N_810,In_402,In_720);
and U811 (N_811,In_467,In_991);
and U812 (N_812,In_400,In_49);
and U813 (N_813,In_10,In_116);
nor U814 (N_814,In_623,In_334);
nor U815 (N_815,In_999,In_250);
and U816 (N_816,In_704,In_856);
or U817 (N_817,In_731,In_443);
or U818 (N_818,In_329,In_500);
or U819 (N_819,In_353,In_259);
nand U820 (N_820,In_589,In_532);
and U821 (N_821,In_677,In_792);
nand U822 (N_822,In_72,In_325);
and U823 (N_823,In_834,In_752);
nand U824 (N_824,In_12,In_848);
nand U825 (N_825,In_810,In_211);
and U826 (N_826,In_89,In_81);
or U827 (N_827,In_554,In_412);
and U828 (N_828,In_986,In_827);
xor U829 (N_829,In_388,In_154);
or U830 (N_830,In_356,In_243);
nand U831 (N_831,In_494,In_565);
nand U832 (N_832,In_279,In_116);
or U833 (N_833,In_39,In_609);
or U834 (N_834,In_926,In_128);
or U835 (N_835,In_551,In_179);
or U836 (N_836,In_854,In_422);
and U837 (N_837,In_652,In_21);
nor U838 (N_838,In_486,In_827);
nor U839 (N_839,In_592,In_738);
and U840 (N_840,In_600,In_356);
nor U841 (N_841,In_810,In_818);
nand U842 (N_842,In_28,In_273);
nor U843 (N_843,In_490,In_401);
nor U844 (N_844,In_49,In_220);
nand U845 (N_845,In_523,In_932);
nor U846 (N_846,In_882,In_391);
or U847 (N_847,In_117,In_580);
nand U848 (N_848,In_581,In_113);
xor U849 (N_849,In_613,In_819);
or U850 (N_850,In_15,In_626);
nor U851 (N_851,In_699,In_964);
or U852 (N_852,In_77,In_750);
and U853 (N_853,In_907,In_594);
and U854 (N_854,In_152,In_708);
and U855 (N_855,In_570,In_842);
or U856 (N_856,In_90,In_924);
or U857 (N_857,In_504,In_793);
and U858 (N_858,In_961,In_516);
or U859 (N_859,In_590,In_146);
nand U860 (N_860,In_358,In_937);
and U861 (N_861,In_395,In_747);
and U862 (N_862,In_936,In_805);
and U863 (N_863,In_646,In_817);
nand U864 (N_864,In_89,In_886);
and U865 (N_865,In_929,In_647);
or U866 (N_866,In_550,In_458);
nor U867 (N_867,In_176,In_701);
nor U868 (N_868,In_262,In_344);
or U869 (N_869,In_543,In_857);
nand U870 (N_870,In_73,In_262);
nor U871 (N_871,In_521,In_520);
nor U872 (N_872,In_652,In_347);
or U873 (N_873,In_664,In_981);
or U874 (N_874,In_908,In_826);
and U875 (N_875,In_578,In_219);
nor U876 (N_876,In_214,In_413);
and U877 (N_877,In_340,In_38);
or U878 (N_878,In_777,In_461);
and U879 (N_879,In_522,In_818);
nand U880 (N_880,In_971,In_176);
or U881 (N_881,In_540,In_606);
nor U882 (N_882,In_644,In_475);
and U883 (N_883,In_393,In_15);
and U884 (N_884,In_480,In_329);
and U885 (N_885,In_715,In_993);
and U886 (N_886,In_958,In_604);
nand U887 (N_887,In_906,In_619);
and U888 (N_888,In_281,In_342);
nand U889 (N_889,In_43,In_109);
or U890 (N_890,In_645,In_609);
or U891 (N_891,In_66,In_508);
nor U892 (N_892,In_467,In_24);
and U893 (N_893,In_92,In_678);
nor U894 (N_894,In_949,In_423);
nor U895 (N_895,In_666,In_367);
or U896 (N_896,In_890,In_228);
or U897 (N_897,In_728,In_317);
and U898 (N_898,In_959,In_741);
and U899 (N_899,In_527,In_206);
xnor U900 (N_900,In_767,In_741);
or U901 (N_901,In_738,In_128);
and U902 (N_902,In_741,In_641);
nand U903 (N_903,In_141,In_558);
nand U904 (N_904,In_966,In_695);
and U905 (N_905,In_513,In_911);
and U906 (N_906,In_327,In_930);
nor U907 (N_907,In_615,In_497);
or U908 (N_908,In_588,In_130);
nand U909 (N_909,In_227,In_107);
and U910 (N_910,In_17,In_843);
or U911 (N_911,In_574,In_705);
nor U912 (N_912,In_129,In_503);
and U913 (N_913,In_824,In_468);
or U914 (N_914,In_849,In_933);
and U915 (N_915,In_400,In_43);
nand U916 (N_916,In_88,In_416);
nand U917 (N_917,In_306,In_764);
or U918 (N_918,In_112,In_790);
or U919 (N_919,In_484,In_674);
or U920 (N_920,In_188,In_108);
nor U921 (N_921,In_622,In_184);
or U922 (N_922,In_601,In_196);
nor U923 (N_923,In_667,In_202);
nand U924 (N_924,In_896,In_673);
or U925 (N_925,In_27,In_684);
or U926 (N_926,In_429,In_981);
and U927 (N_927,In_864,In_974);
or U928 (N_928,In_190,In_281);
nand U929 (N_929,In_218,In_281);
and U930 (N_930,In_995,In_798);
nor U931 (N_931,In_949,In_841);
nand U932 (N_932,In_705,In_119);
or U933 (N_933,In_337,In_386);
and U934 (N_934,In_781,In_888);
nand U935 (N_935,In_774,In_548);
nand U936 (N_936,In_814,In_966);
and U937 (N_937,In_663,In_939);
or U938 (N_938,In_264,In_57);
nor U939 (N_939,In_601,In_745);
or U940 (N_940,In_153,In_730);
or U941 (N_941,In_794,In_553);
and U942 (N_942,In_443,In_404);
and U943 (N_943,In_199,In_816);
nand U944 (N_944,In_122,In_488);
or U945 (N_945,In_822,In_706);
and U946 (N_946,In_307,In_157);
or U947 (N_947,In_210,In_352);
or U948 (N_948,In_939,In_545);
nor U949 (N_949,In_627,In_279);
nor U950 (N_950,In_557,In_284);
or U951 (N_951,In_559,In_348);
and U952 (N_952,In_202,In_6);
or U953 (N_953,In_862,In_32);
or U954 (N_954,In_486,In_216);
nor U955 (N_955,In_694,In_374);
nand U956 (N_956,In_741,In_875);
nor U957 (N_957,In_255,In_540);
and U958 (N_958,In_24,In_750);
and U959 (N_959,In_939,In_161);
or U960 (N_960,In_834,In_708);
nand U961 (N_961,In_206,In_820);
nor U962 (N_962,In_835,In_100);
nor U963 (N_963,In_106,In_550);
nor U964 (N_964,In_339,In_439);
and U965 (N_965,In_48,In_220);
nor U966 (N_966,In_450,In_840);
or U967 (N_967,In_985,In_913);
and U968 (N_968,In_123,In_191);
or U969 (N_969,In_136,In_987);
and U970 (N_970,In_144,In_284);
nand U971 (N_971,In_0,In_144);
or U972 (N_972,In_751,In_258);
and U973 (N_973,In_324,In_544);
nand U974 (N_974,In_378,In_421);
or U975 (N_975,In_534,In_513);
nor U976 (N_976,In_353,In_892);
nor U977 (N_977,In_850,In_129);
and U978 (N_978,In_513,In_442);
or U979 (N_979,In_655,In_592);
or U980 (N_980,In_855,In_985);
nand U981 (N_981,In_376,In_380);
nor U982 (N_982,In_49,In_273);
or U983 (N_983,In_519,In_669);
and U984 (N_984,In_849,In_68);
nand U985 (N_985,In_284,In_207);
or U986 (N_986,In_90,In_361);
nand U987 (N_987,In_816,In_538);
and U988 (N_988,In_882,In_5);
or U989 (N_989,In_506,In_105);
or U990 (N_990,In_550,In_836);
nor U991 (N_991,In_758,In_673);
nand U992 (N_992,In_737,In_186);
nor U993 (N_993,In_680,In_184);
and U994 (N_994,In_167,In_631);
nor U995 (N_995,In_218,In_66);
and U996 (N_996,In_566,In_10);
nand U997 (N_997,In_897,In_607);
nand U998 (N_998,In_247,In_376);
and U999 (N_999,In_220,In_904);
nor U1000 (N_1000,N_803,N_576);
and U1001 (N_1001,N_126,N_880);
or U1002 (N_1002,N_608,N_638);
nand U1003 (N_1003,N_781,N_312);
and U1004 (N_1004,N_481,N_221);
or U1005 (N_1005,N_814,N_611);
nand U1006 (N_1006,N_977,N_67);
nor U1007 (N_1007,N_345,N_805);
nor U1008 (N_1008,N_914,N_228);
or U1009 (N_1009,N_199,N_770);
or U1010 (N_1010,N_112,N_734);
nand U1011 (N_1011,N_419,N_782);
nand U1012 (N_1012,N_148,N_704);
and U1013 (N_1013,N_139,N_716);
and U1014 (N_1014,N_722,N_999);
nor U1015 (N_1015,N_754,N_203);
nand U1016 (N_1016,N_122,N_788);
nor U1017 (N_1017,N_687,N_108);
or U1018 (N_1018,N_653,N_769);
or U1019 (N_1019,N_86,N_322);
nor U1020 (N_1020,N_615,N_629);
nand U1021 (N_1021,N_462,N_568);
nor U1022 (N_1022,N_171,N_390);
or U1023 (N_1023,N_65,N_170);
nand U1024 (N_1024,N_23,N_969);
or U1025 (N_1025,N_52,N_229);
or U1026 (N_1026,N_226,N_428);
nor U1027 (N_1027,N_516,N_91);
nand U1028 (N_1028,N_667,N_246);
or U1029 (N_1029,N_938,N_966);
nor U1030 (N_1030,N_301,N_726);
or U1031 (N_1031,N_719,N_15);
or U1032 (N_1032,N_949,N_937);
or U1033 (N_1033,N_299,N_596);
and U1034 (N_1034,N_383,N_832);
nor U1035 (N_1035,N_41,N_696);
and U1036 (N_1036,N_924,N_297);
or U1037 (N_1037,N_705,N_910);
and U1038 (N_1038,N_386,N_800);
nand U1039 (N_1039,N_980,N_265);
and U1040 (N_1040,N_442,N_842);
nor U1041 (N_1041,N_406,N_375);
nor U1042 (N_1042,N_374,N_304);
and U1043 (N_1043,N_378,N_731);
nand U1044 (N_1044,N_616,N_495);
nand U1045 (N_1045,N_56,N_85);
xnor U1046 (N_1046,N_556,N_703);
xnor U1047 (N_1047,N_467,N_780);
and U1048 (N_1048,N_167,N_790);
or U1049 (N_1049,N_876,N_786);
nor U1050 (N_1050,N_119,N_166);
nor U1051 (N_1051,N_518,N_929);
nor U1052 (N_1052,N_522,N_371);
and U1053 (N_1053,N_831,N_453);
nor U1054 (N_1054,N_848,N_225);
nand U1055 (N_1055,N_733,N_279);
and U1056 (N_1056,N_163,N_593);
nor U1057 (N_1057,N_164,N_373);
or U1058 (N_1058,N_735,N_196);
or U1059 (N_1059,N_872,N_998);
or U1060 (N_1060,N_422,N_338);
nand U1061 (N_1061,N_305,N_101);
or U1062 (N_1062,N_114,N_271);
nand U1063 (N_1063,N_845,N_923);
and U1064 (N_1064,N_544,N_895);
nand U1065 (N_1065,N_81,N_451);
xnor U1066 (N_1066,N_124,N_524);
or U1067 (N_1067,N_247,N_44);
xnor U1068 (N_1068,N_702,N_72);
nor U1069 (N_1069,N_686,N_652);
and U1070 (N_1070,N_597,N_361);
or U1071 (N_1071,N_478,N_380);
nand U1072 (N_1072,N_477,N_985);
nor U1073 (N_1073,N_943,N_626);
nor U1074 (N_1074,N_835,N_963);
or U1075 (N_1075,N_22,N_517);
and U1076 (N_1076,N_62,N_490);
xnor U1077 (N_1077,N_257,N_793);
and U1078 (N_1078,N_314,N_992);
and U1079 (N_1079,N_765,N_210);
and U1080 (N_1080,N_384,N_70);
or U1081 (N_1081,N_717,N_801);
and U1082 (N_1082,N_309,N_752);
nand U1083 (N_1083,N_492,N_715);
or U1084 (N_1084,N_349,N_244);
nand U1085 (N_1085,N_179,N_713);
and U1086 (N_1086,N_681,N_526);
or U1087 (N_1087,N_655,N_824);
or U1088 (N_1088,N_856,N_212);
nor U1089 (N_1089,N_973,N_446);
nor U1090 (N_1090,N_63,N_673);
and U1091 (N_1091,N_989,N_181);
and U1092 (N_1092,N_77,N_818);
nor U1093 (N_1093,N_987,N_3);
and U1094 (N_1094,N_511,N_891);
or U1095 (N_1095,N_443,N_435);
nand U1096 (N_1096,N_946,N_636);
and U1097 (N_1097,N_887,N_609);
and U1098 (N_1098,N_767,N_382);
or U1099 (N_1099,N_188,N_359);
xor U1100 (N_1100,N_874,N_828);
nand U1101 (N_1101,N_9,N_316);
or U1102 (N_1102,N_587,N_589);
nand U1103 (N_1103,N_941,N_337);
nand U1104 (N_1104,N_591,N_857);
and U1105 (N_1105,N_395,N_209);
and U1106 (N_1106,N_925,N_127);
and U1107 (N_1107,N_557,N_951);
and U1108 (N_1108,N_303,N_54);
and U1109 (N_1109,N_808,N_965);
and U1110 (N_1110,N_952,N_764);
nor U1111 (N_1111,N_506,N_459);
or U1112 (N_1112,N_336,N_829);
nand U1113 (N_1113,N_68,N_649);
nor U1114 (N_1114,N_707,N_956);
xor U1115 (N_1115,N_894,N_330);
nor U1116 (N_1116,N_975,N_281);
and U1117 (N_1117,N_513,N_817);
nand U1118 (N_1118,N_236,N_414);
nand U1119 (N_1119,N_551,N_485);
nor U1120 (N_1120,N_892,N_353);
nand U1121 (N_1121,N_538,N_307);
nand U1122 (N_1122,N_133,N_635);
and U1123 (N_1123,N_493,N_860);
nand U1124 (N_1124,N_791,N_675);
and U1125 (N_1125,N_919,N_525);
nor U1126 (N_1126,N_574,N_683);
or U1127 (N_1127,N_700,N_515);
or U1128 (N_1128,N_457,N_147);
and U1129 (N_1129,N_529,N_291);
and U1130 (N_1130,N_315,N_740);
and U1131 (N_1131,N_473,N_751);
nand U1132 (N_1132,N_233,N_785);
or U1133 (N_1133,N_282,N_376);
and U1134 (N_1134,N_935,N_121);
nand U1135 (N_1135,N_146,N_745);
nor U1136 (N_1136,N_913,N_193);
nand U1137 (N_1137,N_758,N_555);
or U1138 (N_1138,N_420,N_862);
and U1139 (N_1139,N_18,N_908);
nor U1140 (N_1140,N_363,N_311);
xor U1141 (N_1141,N_864,N_253);
nand U1142 (N_1142,N_933,N_886);
nand U1143 (N_1143,N_614,N_184);
nor U1144 (N_1144,N_151,N_932);
nand U1145 (N_1145,N_200,N_332);
nor U1146 (N_1146,N_125,N_415);
xnor U1147 (N_1147,N_631,N_218);
or U1148 (N_1148,N_942,N_501);
and U1149 (N_1149,N_604,N_333);
nor U1150 (N_1150,N_177,N_152);
nand U1151 (N_1151,N_392,N_601);
nor U1152 (N_1152,N_458,N_508);
and U1153 (N_1153,N_639,N_882);
nand U1154 (N_1154,N_662,N_192);
nor U1155 (N_1155,N_429,N_342);
or U1156 (N_1156,N_340,N_520);
and U1157 (N_1157,N_504,N_656);
and U1158 (N_1158,N_438,N_476);
and U1159 (N_1159,N_73,N_772);
and U1160 (N_1160,N_400,N_798);
and U1161 (N_1161,N_996,N_205);
nand U1162 (N_1162,N_640,N_208);
or U1163 (N_1163,N_198,N_439);
nor U1164 (N_1164,N_674,N_69);
nor U1165 (N_1165,N_632,N_335);
nor U1166 (N_1166,N_401,N_721);
nand U1167 (N_1167,N_302,N_534);
or U1168 (N_1168,N_671,N_778);
or U1169 (N_1169,N_581,N_118);
nor U1170 (N_1170,N_387,N_404);
or U1171 (N_1171,N_447,N_663);
nor U1172 (N_1172,N_795,N_417);
nor U1173 (N_1173,N_792,N_317);
or U1174 (N_1174,N_402,N_79);
nand U1175 (N_1175,N_36,N_960);
and U1176 (N_1176,N_405,N_658);
and U1177 (N_1177,N_452,N_92);
nor U1178 (N_1178,N_89,N_248);
and U1179 (N_1179,N_245,N_619);
xnor U1180 (N_1180,N_796,N_427);
nor U1181 (N_1181,N_742,N_98);
or U1182 (N_1182,N_621,N_283);
or U1183 (N_1183,N_99,N_123);
or U1184 (N_1184,N_165,N_558);
nand U1185 (N_1185,N_741,N_49);
nor U1186 (N_1186,N_928,N_947);
and U1187 (N_1187,N_761,N_870);
and U1188 (N_1188,N_454,N_915);
xnor U1189 (N_1189,N_318,N_809);
or U1190 (N_1190,N_34,N_261);
or U1191 (N_1191,N_836,N_145);
and U1192 (N_1192,N_252,N_554);
and U1193 (N_1193,N_699,N_60);
nand U1194 (N_1194,N_777,N_17);
and U1195 (N_1195,N_313,N_143);
nor U1196 (N_1196,N_564,N_714);
nand U1197 (N_1197,N_861,N_103);
or U1198 (N_1198,N_579,N_553);
or U1199 (N_1199,N_606,N_308);
and U1200 (N_1200,N_409,N_42);
nor U1201 (N_1201,N_250,N_364);
or U1202 (N_1202,N_66,N_142);
nor U1203 (N_1203,N_241,N_900);
nand U1204 (N_1204,N_979,N_744);
and U1205 (N_1205,N_659,N_189);
nor U1206 (N_1206,N_633,N_762);
or U1207 (N_1207,N_134,N_905);
and U1208 (N_1208,N_853,N_217);
nand U1209 (N_1209,N_347,N_569);
or U1210 (N_1210,N_496,N_917);
nand U1211 (N_1211,N_903,N_695);
nand U1212 (N_1212,N_37,N_768);
or U1213 (N_1213,N_676,N_665);
or U1214 (N_1214,N_61,N_821);
nand U1215 (N_1215,N_78,N_990);
nand U1216 (N_1216,N_75,N_183);
and U1217 (N_1217,N_201,N_31);
xnor U1218 (N_1218,N_488,N_970);
nor U1219 (N_1219,N_76,N_623);
nor U1220 (N_1220,N_185,N_190);
and U1221 (N_1221,N_827,N_546);
nor U1222 (N_1222,N_377,N_162);
or U1223 (N_1223,N_953,N_502);
nor U1224 (N_1224,N_270,N_156);
nor U1225 (N_1225,N_865,N_819);
or U1226 (N_1226,N_595,N_296);
nor U1227 (N_1227,N_412,N_605);
nor U1228 (N_1228,N_637,N_904);
or U1229 (N_1229,N_219,N_276);
nor U1230 (N_1230,N_617,N_749);
nand U1231 (N_1231,N_945,N_465);
and U1232 (N_1232,N_355,N_242);
or U1233 (N_1233,N_784,N_691);
or U1234 (N_1234,N_955,N_214);
and U1235 (N_1235,N_560,N_434);
and U1236 (N_1236,N_433,N_48);
or U1237 (N_1237,N_565,N_231);
or U1238 (N_1238,N_815,N_756);
nand U1239 (N_1239,N_25,N_11);
or U1240 (N_1240,N_223,N_584);
xnor U1241 (N_1241,N_890,N_96);
and U1242 (N_1242,N_852,N_144);
nor U1243 (N_1243,N_24,N_487);
nor U1244 (N_1244,N_110,N_612);
nand U1245 (N_1245,N_295,N_540);
and U1246 (N_1246,N_263,N_7);
and U1247 (N_1247,N_549,N_95);
or U1248 (N_1248,N_550,N_986);
and U1249 (N_1249,N_881,N_366);
nor U1250 (N_1250,N_779,N_875);
nor U1251 (N_1251,N_413,N_350);
or U1252 (N_1252,N_878,N_491);
and U1253 (N_1253,N_255,N_149);
nand U1254 (N_1254,N_213,N_883);
nor U1255 (N_1255,N_826,N_918);
nand U1256 (N_1256,N_503,N_13);
or U1257 (N_1257,N_39,N_570);
or U1258 (N_1258,N_463,N_607);
nor U1259 (N_1259,N_358,N_227);
or U1260 (N_1260,N_645,N_512);
nand U1261 (N_1261,N_537,N_160);
and U1262 (N_1262,N_927,N_186);
and U1263 (N_1263,N_258,N_293);
nand U1264 (N_1264,N_922,N_470);
or U1265 (N_1265,N_460,N_837);
and U1266 (N_1266,N_855,N_718);
nand U1267 (N_1267,N_50,N_562);
nand U1268 (N_1268,N_911,N_893);
or U1269 (N_1269,N_590,N_399);
or U1270 (N_1270,N_622,N_578);
and U1271 (N_1271,N_907,N_425);
nand U1272 (N_1272,N_624,N_176);
nor U1273 (N_1273,N_141,N_379);
or U1274 (N_1274,N_360,N_321);
and U1275 (N_1275,N_306,N_53);
nor U1276 (N_1276,N_902,N_958);
and U1277 (N_1277,N_320,N_266);
nor U1278 (N_1278,N_725,N_489);
nand U1279 (N_1279,N_220,N_885);
nor U1280 (N_1280,N_240,N_230);
nand U1281 (N_1281,N_899,N_732);
nand U1282 (N_1282,N_479,N_535);
nor U1283 (N_1283,N_961,N_117);
nand U1284 (N_1284,N_339,N_294);
or U1285 (N_1285,N_251,N_794);
nand U1286 (N_1286,N_968,N_129);
nand U1287 (N_1287,N_421,N_354);
nand U1288 (N_1288,N_329,N_243);
or U1289 (N_1289,N_344,N_692);
or U1290 (N_1290,N_71,N_328);
nand U1291 (N_1291,N_706,N_416);
and U1292 (N_1292,N_547,N_59);
nor U1293 (N_1293,N_367,N_753);
or U1294 (N_1294,N_84,N_51);
and U1295 (N_1295,N_131,N_100);
nor U1296 (N_1296,N_690,N_563);
or U1297 (N_1297,N_672,N_277);
and U1298 (N_1298,N_33,N_484);
nor U1299 (N_1299,N_444,N_499);
nor U1300 (N_1300,N_341,N_369);
nand U1301 (N_1301,N_430,N_527);
nor U1302 (N_1302,N_838,N_161);
and U1303 (N_1303,N_536,N_411);
nand U1304 (N_1304,N_259,N_850);
and U1305 (N_1305,N_682,N_825);
and U1306 (N_1306,N_300,N_763);
nor U1307 (N_1307,N_356,N_278);
or U1308 (N_1308,N_224,N_351);
nand U1309 (N_1309,N_543,N_567);
nand U1310 (N_1310,N_841,N_869);
or U1311 (N_1311,N_153,N_58);
nand U1312 (N_1312,N_994,N_995);
nand U1313 (N_1313,N_74,N_115);
or U1314 (N_1314,N_464,N_884);
or U1315 (N_1315,N_747,N_720);
nor U1316 (N_1316,N_743,N_254);
and U1317 (N_1317,N_710,N_195);
and U1318 (N_1318,N_173,N_594);
or U1319 (N_1319,N_172,N_140);
or U1320 (N_1320,N_936,N_909);
or U1321 (N_1321,N_35,N_106);
nor U1322 (N_1322,N_847,N_976);
nand U1323 (N_1323,N_272,N_776);
nand U1324 (N_1324,N_158,N_934);
and U1325 (N_1325,N_4,N_8);
nand U1326 (N_1326,N_206,N_204);
and U1327 (N_1327,N_510,N_432);
or U1328 (N_1328,N_993,N_40);
nor U1329 (N_1329,N_222,N_483);
or U1330 (N_1330,N_709,N_810);
or U1331 (N_1331,N_482,N_249);
nor U1332 (N_1332,N_239,N_577);
and U1333 (N_1333,N_868,N_531);
nor U1334 (N_1334,N_461,N_583);
or U1335 (N_1335,N_967,N_334);
nand U1336 (N_1336,N_135,N_984);
nor U1337 (N_1337,N_269,N_46);
nand U1338 (N_1338,N_552,N_175);
nand U1339 (N_1339,N_468,N_262);
or U1340 (N_1340,N_739,N_55);
and U1341 (N_1341,N_613,N_102);
and U1342 (N_1342,N_728,N_654);
or U1343 (N_1343,N_618,N_324);
xnor U1344 (N_1344,N_685,N_711);
and U1345 (N_1345,N_668,N_723);
nand U1346 (N_1346,N_991,N_187);
nand U1347 (N_1347,N_851,N_174);
nor U1348 (N_1348,N_64,N_603);
or U1349 (N_1349,N_440,N_275);
nand U1350 (N_1350,N_448,N_90);
or U1351 (N_1351,N_310,N_548);
nor U1352 (N_1352,N_916,N_274);
nand U1353 (N_1353,N_298,N_456);
nand U1354 (N_1354,N_43,N_804);
xor U1355 (N_1355,N_766,N_729);
nand U1356 (N_1356,N_388,N_641);
nand U1357 (N_1357,N_2,N_698);
or U1358 (N_1358,N_530,N_789);
and U1359 (N_1359,N_580,N_82);
and U1360 (N_1360,N_394,N_787);
and U1361 (N_1361,N_666,N_684);
or U1362 (N_1362,N_811,N_475);
xnor U1363 (N_1363,N_888,N_498);
and U1364 (N_1364,N_357,N_450);
nor U1365 (N_1365,N_634,N_5);
or U1366 (N_1366,N_507,N_211);
nor U1367 (N_1367,N_45,N_974);
or U1368 (N_1368,N_844,N_136);
and U1369 (N_1369,N_441,N_866);
and U1370 (N_1370,N_849,N_396);
nor U1371 (N_1371,N_625,N_113);
and U1372 (N_1372,N_207,N_712);
nand U1373 (N_1373,N_830,N_32);
nand U1374 (N_1374,N_418,N_182);
and U1375 (N_1375,N_27,N_783);
and U1376 (N_1376,N_571,N_287);
or U1377 (N_1377,N_197,N_403);
or U1378 (N_1378,N_846,N_839);
nor U1379 (N_1379,N_10,N_16);
xnor U1380 (N_1380,N_87,N_325);
or U1381 (N_1381,N_964,N_650);
or U1382 (N_1382,N_109,N_694);
or U1383 (N_1383,N_738,N_408);
or U1384 (N_1384,N_981,N_867);
xnor U1385 (N_1385,N_661,N_627);
nor U1386 (N_1386,N_268,N_948);
nand U1387 (N_1387,N_748,N_954);
nand U1388 (N_1388,N_107,N_533);
and U1389 (N_1389,N_545,N_120);
nand U1390 (N_1390,N_348,N_234);
nand U1391 (N_1391,N_391,N_47);
or U1392 (N_1392,N_859,N_760);
and U1393 (N_1393,N_863,N_437);
nor U1394 (N_1394,N_191,N_858);
and U1395 (N_1395,N_877,N_727);
xor U1396 (N_1396,N_630,N_497);
nor U1397 (N_1397,N_372,N_21);
and U1398 (N_1398,N_202,N_128);
nor U1399 (N_1399,N_813,N_284);
or U1400 (N_1400,N_931,N_843);
or U1401 (N_1401,N_137,N_29);
nand U1402 (N_1402,N_940,N_424);
or U1403 (N_1403,N_326,N_155);
nand U1404 (N_1404,N_944,N_921);
nand U1405 (N_1405,N_971,N_235);
nand U1406 (N_1406,N_802,N_26);
nor U1407 (N_1407,N_180,N_346);
and U1408 (N_1408,N_708,N_730);
nor U1409 (N_1409,N_678,N_930);
nand U1410 (N_1410,N_598,N_610);
nor U1411 (N_1411,N_178,N_288);
nand U1412 (N_1412,N_343,N_644);
or U1413 (N_1413,N_912,N_573);
or U1414 (N_1414,N_959,N_697);
nor U1415 (N_1415,N_988,N_651);
nor U1416 (N_1416,N_154,N_519);
nand U1417 (N_1417,N_474,N_559);
and U1418 (N_1418,N_449,N_0);
and U1419 (N_1419,N_6,N_736);
and U1420 (N_1420,N_680,N_292);
nor U1421 (N_1421,N_600,N_397);
or U1422 (N_1422,N_471,N_12);
and U1423 (N_1423,N_585,N_806);
nand U1424 (N_1424,N_168,N_57);
and U1425 (N_1425,N_539,N_331);
or U1426 (N_1426,N_664,N_628);
or U1427 (N_1427,N_509,N_472);
nand U1428 (N_1428,N_897,N_407);
xnor U1429 (N_1429,N_939,N_657);
and U1430 (N_1430,N_646,N_398);
nor U1431 (N_1431,N_582,N_393);
nor U1432 (N_1432,N_820,N_642);
or U1433 (N_1433,N_799,N_445);
or U1434 (N_1434,N_327,N_14);
or U1435 (N_1435,N_28,N_486);
nand U1436 (N_1436,N_104,N_822);
nor U1437 (N_1437,N_572,N_370);
nand U1438 (N_1438,N_431,N_647);
nand U1439 (N_1439,N_215,N_669);
nand U1440 (N_1440,N_352,N_232);
nor U1441 (N_1441,N_812,N_873);
nand U1442 (N_1442,N_19,N_514);
nand U1443 (N_1443,N_586,N_602);
and U1444 (N_1444,N_286,N_194);
or U1445 (N_1445,N_494,N_643);
nor U1446 (N_1446,N_528,N_797);
and U1447 (N_1447,N_256,N_264);
or U1448 (N_1448,N_532,N_410);
nor U1449 (N_1449,N_833,N_840);
or U1450 (N_1450,N_901,N_521);
and U1451 (N_1451,N_130,N_365);
and U1452 (N_1452,N_648,N_169);
nor U1453 (N_1453,N_620,N_542);
and U1454 (N_1454,N_724,N_896);
and U1455 (N_1455,N_426,N_926);
or U1456 (N_1456,N_93,N_323);
or U1457 (N_1457,N_816,N_920);
nand U1458 (N_1458,N_138,N_290);
nor U1459 (N_1459,N_1,N_997);
xor U1460 (N_1460,N_561,N_20);
nand U1461 (N_1461,N_957,N_962);
or U1462 (N_1462,N_80,N_746);
and U1463 (N_1463,N_807,N_30);
or U1464 (N_1464,N_660,N_116);
nor U1465 (N_1465,N_775,N_319);
and U1466 (N_1466,N_469,N_950);
or U1467 (N_1467,N_906,N_774);
nand U1468 (N_1468,N_834,N_105);
nor U1469 (N_1469,N_679,N_588);
or U1470 (N_1470,N_750,N_677);
and U1471 (N_1471,N_83,N_982);
nand U1472 (N_1472,N_280,N_879);
nor U1473 (N_1473,N_455,N_368);
and U1474 (N_1474,N_566,N_94);
nor U1475 (N_1475,N_436,N_500);
and U1476 (N_1476,N_523,N_983);
nor U1477 (N_1477,N_385,N_898);
nand U1478 (N_1478,N_132,N_150);
nor U1479 (N_1479,N_889,N_541);
xor U1480 (N_1480,N_689,N_260);
nor U1481 (N_1481,N_389,N_688);
nor U1482 (N_1482,N_670,N_771);
nor U1483 (N_1483,N_267,N_423);
nand U1484 (N_1484,N_823,N_755);
nand U1485 (N_1485,N_592,N_88);
nand U1486 (N_1486,N_773,N_757);
nand U1487 (N_1487,N_978,N_599);
xor U1488 (N_1488,N_693,N_111);
nor U1489 (N_1489,N_701,N_159);
nand U1490 (N_1490,N_854,N_237);
nor U1491 (N_1491,N_285,N_575);
or U1492 (N_1492,N_362,N_480);
nor U1493 (N_1493,N_466,N_505);
nor U1494 (N_1494,N_871,N_216);
and U1495 (N_1495,N_97,N_972);
nand U1496 (N_1496,N_273,N_289);
and U1497 (N_1497,N_38,N_157);
nand U1498 (N_1498,N_381,N_759);
and U1499 (N_1499,N_737,N_238);
and U1500 (N_1500,N_356,N_349);
nand U1501 (N_1501,N_152,N_396);
nand U1502 (N_1502,N_477,N_761);
nor U1503 (N_1503,N_475,N_745);
or U1504 (N_1504,N_970,N_865);
and U1505 (N_1505,N_426,N_40);
nor U1506 (N_1506,N_913,N_623);
nor U1507 (N_1507,N_65,N_243);
nor U1508 (N_1508,N_667,N_64);
and U1509 (N_1509,N_184,N_413);
or U1510 (N_1510,N_216,N_268);
nand U1511 (N_1511,N_269,N_640);
and U1512 (N_1512,N_349,N_879);
and U1513 (N_1513,N_341,N_818);
nand U1514 (N_1514,N_394,N_740);
and U1515 (N_1515,N_775,N_480);
and U1516 (N_1516,N_968,N_736);
nor U1517 (N_1517,N_354,N_444);
nor U1518 (N_1518,N_294,N_432);
nor U1519 (N_1519,N_812,N_41);
or U1520 (N_1520,N_543,N_711);
nor U1521 (N_1521,N_577,N_339);
nand U1522 (N_1522,N_405,N_36);
nor U1523 (N_1523,N_239,N_613);
and U1524 (N_1524,N_366,N_146);
nand U1525 (N_1525,N_503,N_123);
and U1526 (N_1526,N_495,N_380);
nor U1527 (N_1527,N_239,N_370);
nor U1528 (N_1528,N_183,N_531);
or U1529 (N_1529,N_975,N_416);
and U1530 (N_1530,N_677,N_430);
nand U1531 (N_1531,N_423,N_904);
and U1532 (N_1532,N_350,N_504);
nand U1533 (N_1533,N_623,N_759);
nand U1534 (N_1534,N_909,N_186);
and U1535 (N_1535,N_367,N_755);
nand U1536 (N_1536,N_400,N_173);
or U1537 (N_1537,N_863,N_747);
and U1538 (N_1538,N_927,N_905);
and U1539 (N_1539,N_409,N_683);
nor U1540 (N_1540,N_671,N_24);
and U1541 (N_1541,N_857,N_371);
nor U1542 (N_1542,N_67,N_515);
or U1543 (N_1543,N_827,N_318);
or U1544 (N_1544,N_242,N_108);
and U1545 (N_1545,N_759,N_898);
or U1546 (N_1546,N_981,N_276);
and U1547 (N_1547,N_260,N_699);
nand U1548 (N_1548,N_351,N_176);
or U1549 (N_1549,N_966,N_188);
or U1550 (N_1550,N_81,N_931);
and U1551 (N_1551,N_47,N_240);
nand U1552 (N_1552,N_933,N_18);
nor U1553 (N_1553,N_455,N_153);
nand U1554 (N_1554,N_278,N_712);
nor U1555 (N_1555,N_403,N_310);
and U1556 (N_1556,N_750,N_129);
nand U1557 (N_1557,N_346,N_519);
nand U1558 (N_1558,N_119,N_64);
nor U1559 (N_1559,N_305,N_855);
nand U1560 (N_1560,N_853,N_419);
and U1561 (N_1561,N_370,N_469);
or U1562 (N_1562,N_472,N_222);
nor U1563 (N_1563,N_701,N_48);
or U1564 (N_1564,N_142,N_769);
or U1565 (N_1565,N_490,N_417);
and U1566 (N_1566,N_599,N_607);
nor U1567 (N_1567,N_576,N_479);
or U1568 (N_1568,N_479,N_277);
nand U1569 (N_1569,N_773,N_192);
or U1570 (N_1570,N_78,N_625);
or U1571 (N_1571,N_883,N_276);
and U1572 (N_1572,N_945,N_348);
nand U1573 (N_1573,N_81,N_310);
nand U1574 (N_1574,N_793,N_889);
nor U1575 (N_1575,N_132,N_889);
nor U1576 (N_1576,N_639,N_689);
and U1577 (N_1577,N_862,N_584);
nor U1578 (N_1578,N_28,N_395);
nor U1579 (N_1579,N_509,N_122);
and U1580 (N_1580,N_424,N_36);
and U1581 (N_1581,N_163,N_332);
nand U1582 (N_1582,N_127,N_467);
nand U1583 (N_1583,N_334,N_261);
or U1584 (N_1584,N_570,N_580);
nand U1585 (N_1585,N_558,N_304);
or U1586 (N_1586,N_880,N_557);
nor U1587 (N_1587,N_393,N_921);
nand U1588 (N_1588,N_746,N_125);
nor U1589 (N_1589,N_184,N_46);
nand U1590 (N_1590,N_273,N_664);
or U1591 (N_1591,N_49,N_730);
nand U1592 (N_1592,N_714,N_252);
and U1593 (N_1593,N_181,N_623);
or U1594 (N_1594,N_148,N_114);
or U1595 (N_1595,N_573,N_474);
nor U1596 (N_1596,N_415,N_971);
and U1597 (N_1597,N_892,N_458);
or U1598 (N_1598,N_797,N_519);
xor U1599 (N_1599,N_91,N_635);
nand U1600 (N_1600,N_553,N_320);
nand U1601 (N_1601,N_752,N_754);
nand U1602 (N_1602,N_791,N_0);
or U1603 (N_1603,N_570,N_866);
nor U1604 (N_1604,N_657,N_220);
xnor U1605 (N_1605,N_901,N_891);
xnor U1606 (N_1606,N_399,N_204);
and U1607 (N_1607,N_952,N_282);
and U1608 (N_1608,N_695,N_904);
and U1609 (N_1609,N_380,N_906);
and U1610 (N_1610,N_420,N_748);
or U1611 (N_1611,N_969,N_805);
and U1612 (N_1612,N_597,N_889);
nand U1613 (N_1613,N_909,N_25);
and U1614 (N_1614,N_82,N_459);
nor U1615 (N_1615,N_252,N_386);
or U1616 (N_1616,N_202,N_686);
nor U1617 (N_1617,N_447,N_925);
or U1618 (N_1618,N_979,N_660);
and U1619 (N_1619,N_478,N_214);
nand U1620 (N_1620,N_15,N_700);
and U1621 (N_1621,N_775,N_743);
or U1622 (N_1622,N_800,N_261);
or U1623 (N_1623,N_826,N_449);
nand U1624 (N_1624,N_149,N_673);
or U1625 (N_1625,N_456,N_337);
nand U1626 (N_1626,N_227,N_947);
or U1627 (N_1627,N_557,N_765);
nor U1628 (N_1628,N_138,N_414);
or U1629 (N_1629,N_468,N_529);
nor U1630 (N_1630,N_316,N_247);
nor U1631 (N_1631,N_317,N_408);
or U1632 (N_1632,N_703,N_285);
or U1633 (N_1633,N_476,N_205);
nor U1634 (N_1634,N_902,N_202);
xor U1635 (N_1635,N_61,N_3);
nand U1636 (N_1636,N_819,N_72);
or U1637 (N_1637,N_286,N_56);
and U1638 (N_1638,N_971,N_786);
or U1639 (N_1639,N_10,N_250);
nand U1640 (N_1640,N_287,N_54);
and U1641 (N_1641,N_394,N_549);
nor U1642 (N_1642,N_824,N_918);
or U1643 (N_1643,N_835,N_54);
and U1644 (N_1644,N_828,N_344);
nor U1645 (N_1645,N_147,N_933);
nor U1646 (N_1646,N_537,N_75);
nand U1647 (N_1647,N_514,N_326);
nor U1648 (N_1648,N_869,N_477);
nand U1649 (N_1649,N_87,N_134);
nand U1650 (N_1650,N_566,N_493);
nor U1651 (N_1651,N_839,N_704);
or U1652 (N_1652,N_425,N_210);
nor U1653 (N_1653,N_836,N_577);
nor U1654 (N_1654,N_155,N_456);
nand U1655 (N_1655,N_738,N_604);
nand U1656 (N_1656,N_889,N_809);
or U1657 (N_1657,N_68,N_245);
and U1658 (N_1658,N_860,N_782);
or U1659 (N_1659,N_352,N_428);
or U1660 (N_1660,N_790,N_65);
and U1661 (N_1661,N_816,N_198);
and U1662 (N_1662,N_297,N_860);
nor U1663 (N_1663,N_183,N_345);
nand U1664 (N_1664,N_86,N_925);
nor U1665 (N_1665,N_782,N_992);
or U1666 (N_1666,N_540,N_98);
and U1667 (N_1667,N_508,N_855);
nor U1668 (N_1668,N_811,N_279);
or U1669 (N_1669,N_148,N_944);
or U1670 (N_1670,N_47,N_596);
and U1671 (N_1671,N_956,N_839);
nand U1672 (N_1672,N_426,N_894);
and U1673 (N_1673,N_923,N_640);
or U1674 (N_1674,N_661,N_674);
or U1675 (N_1675,N_755,N_814);
nor U1676 (N_1676,N_551,N_534);
or U1677 (N_1677,N_812,N_312);
and U1678 (N_1678,N_616,N_104);
and U1679 (N_1679,N_371,N_577);
and U1680 (N_1680,N_511,N_313);
nor U1681 (N_1681,N_978,N_757);
nor U1682 (N_1682,N_857,N_653);
nor U1683 (N_1683,N_755,N_784);
nor U1684 (N_1684,N_880,N_505);
and U1685 (N_1685,N_334,N_201);
nand U1686 (N_1686,N_89,N_905);
and U1687 (N_1687,N_182,N_196);
nand U1688 (N_1688,N_876,N_161);
nor U1689 (N_1689,N_284,N_683);
and U1690 (N_1690,N_969,N_391);
and U1691 (N_1691,N_710,N_552);
nor U1692 (N_1692,N_455,N_717);
nor U1693 (N_1693,N_944,N_236);
nand U1694 (N_1694,N_290,N_958);
nand U1695 (N_1695,N_412,N_562);
and U1696 (N_1696,N_999,N_514);
nor U1697 (N_1697,N_94,N_606);
nand U1698 (N_1698,N_665,N_892);
nand U1699 (N_1699,N_989,N_361);
nand U1700 (N_1700,N_281,N_254);
and U1701 (N_1701,N_78,N_641);
nand U1702 (N_1702,N_830,N_456);
and U1703 (N_1703,N_475,N_656);
nand U1704 (N_1704,N_238,N_755);
nor U1705 (N_1705,N_765,N_550);
and U1706 (N_1706,N_635,N_125);
xor U1707 (N_1707,N_968,N_482);
and U1708 (N_1708,N_754,N_362);
and U1709 (N_1709,N_564,N_58);
nor U1710 (N_1710,N_577,N_950);
nor U1711 (N_1711,N_235,N_90);
nand U1712 (N_1712,N_943,N_424);
or U1713 (N_1713,N_860,N_234);
nand U1714 (N_1714,N_949,N_570);
or U1715 (N_1715,N_709,N_252);
and U1716 (N_1716,N_72,N_805);
and U1717 (N_1717,N_847,N_715);
or U1718 (N_1718,N_52,N_314);
nor U1719 (N_1719,N_883,N_595);
and U1720 (N_1720,N_850,N_856);
nand U1721 (N_1721,N_327,N_852);
and U1722 (N_1722,N_745,N_961);
nand U1723 (N_1723,N_620,N_33);
and U1724 (N_1724,N_544,N_652);
or U1725 (N_1725,N_519,N_753);
and U1726 (N_1726,N_805,N_547);
nor U1727 (N_1727,N_826,N_381);
and U1728 (N_1728,N_712,N_808);
nand U1729 (N_1729,N_147,N_967);
and U1730 (N_1730,N_93,N_508);
and U1731 (N_1731,N_92,N_987);
xnor U1732 (N_1732,N_673,N_774);
or U1733 (N_1733,N_495,N_195);
nor U1734 (N_1734,N_85,N_133);
nand U1735 (N_1735,N_884,N_907);
nor U1736 (N_1736,N_804,N_16);
nor U1737 (N_1737,N_127,N_661);
nor U1738 (N_1738,N_128,N_252);
nor U1739 (N_1739,N_709,N_437);
or U1740 (N_1740,N_497,N_809);
nand U1741 (N_1741,N_7,N_718);
nor U1742 (N_1742,N_807,N_658);
nand U1743 (N_1743,N_674,N_295);
nor U1744 (N_1744,N_818,N_357);
nand U1745 (N_1745,N_507,N_368);
nor U1746 (N_1746,N_336,N_840);
and U1747 (N_1747,N_328,N_359);
xor U1748 (N_1748,N_129,N_730);
nor U1749 (N_1749,N_735,N_354);
and U1750 (N_1750,N_605,N_692);
and U1751 (N_1751,N_350,N_241);
nor U1752 (N_1752,N_82,N_855);
nor U1753 (N_1753,N_393,N_821);
nand U1754 (N_1754,N_892,N_619);
nand U1755 (N_1755,N_168,N_989);
and U1756 (N_1756,N_739,N_40);
nand U1757 (N_1757,N_99,N_274);
nor U1758 (N_1758,N_156,N_672);
nor U1759 (N_1759,N_37,N_254);
nor U1760 (N_1760,N_437,N_668);
or U1761 (N_1761,N_382,N_701);
or U1762 (N_1762,N_927,N_644);
and U1763 (N_1763,N_87,N_583);
nand U1764 (N_1764,N_315,N_196);
or U1765 (N_1765,N_187,N_392);
nand U1766 (N_1766,N_279,N_928);
nand U1767 (N_1767,N_852,N_690);
nand U1768 (N_1768,N_741,N_813);
and U1769 (N_1769,N_100,N_228);
and U1770 (N_1770,N_641,N_356);
and U1771 (N_1771,N_358,N_496);
and U1772 (N_1772,N_947,N_666);
and U1773 (N_1773,N_486,N_242);
nand U1774 (N_1774,N_567,N_835);
and U1775 (N_1775,N_528,N_646);
or U1776 (N_1776,N_779,N_871);
and U1777 (N_1777,N_570,N_612);
and U1778 (N_1778,N_964,N_246);
and U1779 (N_1779,N_858,N_847);
nor U1780 (N_1780,N_179,N_454);
and U1781 (N_1781,N_754,N_561);
or U1782 (N_1782,N_60,N_838);
nand U1783 (N_1783,N_235,N_229);
nor U1784 (N_1784,N_890,N_123);
and U1785 (N_1785,N_511,N_659);
and U1786 (N_1786,N_762,N_862);
and U1787 (N_1787,N_75,N_640);
and U1788 (N_1788,N_481,N_107);
nand U1789 (N_1789,N_165,N_993);
nand U1790 (N_1790,N_242,N_60);
or U1791 (N_1791,N_68,N_386);
nor U1792 (N_1792,N_176,N_778);
nand U1793 (N_1793,N_330,N_27);
nand U1794 (N_1794,N_48,N_422);
nor U1795 (N_1795,N_877,N_99);
or U1796 (N_1796,N_830,N_45);
nor U1797 (N_1797,N_105,N_264);
and U1798 (N_1798,N_711,N_177);
nand U1799 (N_1799,N_530,N_81);
or U1800 (N_1800,N_883,N_165);
and U1801 (N_1801,N_371,N_940);
nand U1802 (N_1802,N_20,N_681);
or U1803 (N_1803,N_475,N_611);
xor U1804 (N_1804,N_475,N_957);
nand U1805 (N_1805,N_807,N_761);
and U1806 (N_1806,N_479,N_132);
nand U1807 (N_1807,N_398,N_534);
and U1808 (N_1808,N_575,N_398);
and U1809 (N_1809,N_97,N_435);
or U1810 (N_1810,N_860,N_960);
xor U1811 (N_1811,N_877,N_531);
nand U1812 (N_1812,N_297,N_780);
nand U1813 (N_1813,N_799,N_364);
and U1814 (N_1814,N_296,N_938);
nor U1815 (N_1815,N_522,N_844);
and U1816 (N_1816,N_593,N_279);
nor U1817 (N_1817,N_144,N_982);
or U1818 (N_1818,N_659,N_841);
nor U1819 (N_1819,N_977,N_795);
or U1820 (N_1820,N_501,N_186);
nor U1821 (N_1821,N_979,N_719);
nand U1822 (N_1822,N_986,N_759);
and U1823 (N_1823,N_429,N_64);
xnor U1824 (N_1824,N_738,N_780);
and U1825 (N_1825,N_987,N_755);
or U1826 (N_1826,N_698,N_397);
or U1827 (N_1827,N_121,N_771);
and U1828 (N_1828,N_452,N_254);
nand U1829 (N_1829,N_510,N_232);
or U1830 (N_1830,N_965,N_378);
and U1831 (N_1831,N_73,N_46);
nand U1832 (N_1832,N_399,N_28);
and U1833 (N_1833,N_559,N_66);
or U1834 (N_1834,N_840,N_724);
nor U1835 (N_1835,N_202,N_593);
nor U1836 (N_1836,N_251,N_328);
and U1837 (N_1837,N_557,N_370);
and U1838 (N_1838,N_521,N_971);
nand U1839 (N_1839,N_199,N_406);
or U1840 (N_1840,N_602,N_57);
nor U1841 (N_1841,N_744,N_521);
nand U1842 (N_1842,N_751,N_387);
and U1843 (N_1843,N_399,N_242);
nand U1844 (N_1844,N_424,N_412);
xor U1845 (N_1845,N_596,N_114);
nor U1846 (N_1846,N_128,N_223);
nor U1847 (N_1847,N_697,N_426);
or U1848 (N_1848,N_826,N_312);
xnor U1849 (N_1849,N_551,N_606);
nand U1850 (N_1850,N_204,N_999);
nand U1851 (N_1851,N_761,N_308);
and U1852 (N_1852,N_183,N_522);
and U1853 (N_1853,N_998,N_863);
nand U1854 (N_1854,N_303,N_729);
nand U1855 (N_1855,N_964,N_861);
nor U1856 (N_1856,N_845,N_546);
nand U1857 (N_1857,N_669,N_169);
or U1858 (N_1858,N_246,N_488);
nand U1859 (N_1859,N_418,N_280);
or U1860 (N_1860,N_862,N_31);
or U1861 (N_1861,N_198,N_56);
or U1862 (N_1862,N_611,N_524);
or U1863 (N_1863,N_498,N_403);
or U1864 (N_1864,N_68,N_819);
or U1865 (N_1865,N_981,N_618);
nand U1866 (N_1866,N_521,N_767);
nor U1867 (N_1867,N_70,N_957);
xor U1868 (N_1868,N_554,N_309);
or U1869 (N_1869,N_267,N_756);
and U1870 (N_1870,N_285,N_247);
or U1871 (N_1871,N_54,N_977);
nor U1872 (N_1872,N_153,N_595);
nor U1873 (N_1873,N_515,N_175);
nand U1874 (N_1874,N_749,N_682);
nand U1875 (N_1875,N_868,N_163);
nor U1876 (N_1876,N_410,N_920);
nor U1877 (N_1877,N_420,N_70);
or U1878 (N_1878,N_199,N_22);
or U1879 (N_1879,N_403,N_75);
nor U1880 (N_1880,N_96,N_919);
nand U1881 (N_1881,N_709,N_53);
or U1882 (N_1882,N_97,N_825);
and U1883 (N_1883,N_117,N_723);
xnor U1884 (N_1884,N_47,N_616);
or U1885 (N_1885,N_873,N_167);
nand U1886 (N_1886,N_315,N_546);
nor U1887 (N_1887,N_947,N_766);
or U1888 (N_1888,N_151,N_902);
nor U1889 (N_1889,N_322,N_922);
or U1890 (N_1890,N_749,N_639);
and U1891 (N_1891,N_154,N_953);
nand U1892 (N_1892,N_386,N_493);
or U1893 (N_1893,N_504,N_753);
nor U1894 (N_1894,N_451,N_426);
nor U1895 (N_1895,N_980,N_408);
and U1896 (N_1896,N_463,N_31);
and U1897 (N_1897,N_366,N_208);
nor U1898 (N_1898,N_625,N_277);
or U1899 (N_1899,N_650,N_470);
nand U1900 (N_1900,N_519,N_392);
nor U1901 (N_1901,N_469,N_189);
nand U1902 (N_1902,N_554,N_862);
nor U1903 (N_1903,N_146,N_312);
and U1904 (N_1904,N_272,N_297);
xor U1905 (N_1905,N_65,N_548);
or U1906 (N_1906,N_597,N_645);
or U1907 (N_1907,N_120,N_147);
or U1908 (N_1908,N_327,N_952);
and U1909 (N_1909,N_840,N_648);
or U1910 (N_1910,N_907,N_657);
nor U1911 (N_1911,N_443,N_659);
nand U1912 (N_1912,N_242,N_769);
and U1913 (N_1913,N_949,N_831);
nand U1914 (N_1914,N_891,N_683);
and U1915 (N_1915,N_863,N_14);
and U1916 (N_1916,N_680,N_301);
nor U1917 (N_1917,N_617,N_159);
nor U1918 (N_1918,N_88,N_967);
nand U1919 (N_1919,N_387,N_436);
or U1920 (N_1920,N_754,N_799);
nand U1921 (N_1921,N_307,N_714);
and U1922 (N_1922,N_222,N_132);
nand U1923 (N_1923,N_228,N_409);
or U1924 (N_1924,N_682,N_545);
and U1925 (N_1925,N_844,N_970);
nand U1926 (N_1926,N_688,N_250);
nand U1927 (N_1927,N_905,N_873);
or U1928 (N_1928,N_613,N_219);
nor U1929 (N_1929,N_621,N_940);
nand U1930 (N_1930,N_320,N_944);
nor U1931 (N_1931,N_235,N_27);
nor U1932 (N_1932,N_282,N_55);
and U1933 (N_1933,N_426,N_115);
nand U1934 (N_1934,N_737,N_333);
or U1935 (N_1935,N_193,N_694);
nor U1936 (N_1936,N_720,N_696);
nor U1937 (N_1937,N_540,N_223);
nand U1938 (N_1938,N_919,N_216);
nand U1939 (N_1939,N_772,N_359);
and U1940 (N_1940,N_636,N_177);
or U1941 (N_1941,N_473,N_21);
and U1942 (N_1942,N_540,N_968);
and U1943 (N_1943,N_510,N_996);
nand U1944 (N_1944,N_116,N_233);
and U1945 (N_1945,N_786,N_233);
or U1946 (N_1946,N_986,N_346);
xor U1947 (N_1947,N_614,N_47);
nor U1948 (N_1948,N_101,N_835);
and U1949 (N_1949,N_428,N_243);
nor U1950 (N_1950,N_608,N_141);
nand U1951 (N_1951,N_705,N_622);
or U1952 (N_1952,N_812,N_217);
nor U1953 (N_1953,N_910,N_855);
nor U1954 (N_1954,N_102,N_31);
and U1955 (N_1955,N_627,N_568);
and U1956 (N_1956,N_580,N_46);
and U1957 (N_1957,N_342,N_692);
nor U1958 (N_1958,N_554,N_588);
or U1959 (N_1959,N_790,N_223);
or U1960 (N_1960,N_356,N_145);
and U1961 (N_1961,N_322,N_4);
or U1962 (N_1962,N_23,N_979);
nand U1963 (N_1963,N_488,N_932);
and U1964 (N_1964,N_210,N_750);
and U1965 (N_1965,N_435,N_511);
nor U1966 (N_1966,N_343,N_367);
and U1967 (N_1967,N_545,N_777);
and U1968 (N_1968,N_15,N_403);
and U1969 (N_1969,N_293,N_175);
and U1970 (N_1970,N_256,N_66);
or U1971 (N_1971,N_680,N_393);
nor U1972 (N_1972,N_168,N_746);
or U1973 (N_1973,N_30,N_778);
and U1974 (N_1974,N_261,N_417);
nand U1975 (N_1975,N_851,N_905);
nor U1976 (N_1976,N_68,N_834);
and U1977 (N_1977,N_288,N_38);
and U1978 (N_1978,N_97,N_101);
or U1979 (N_1979,N_130,N_602);
or U1980 (N_1980,N_20,N_677);
or U1981 (N_1981,N_140,N_256);
nand U1982 (N_1982,N_150,N_111);
and U1983 (N_1983,N_221,N_409);
or U1984 (N_1984,N_319,N_686);
and U1985 (N_1985,N_242,N_799);
and U1986 (N_1986,N_912,N_730);
and U1987 (N_1987,N_445,N_344);
nor U1988 (N_1988,N_480,N_382);
nor U1989 (N_1989,N_852,N_977);
or U1990 (N_1990,N_128,N_347);
nor U1991 (N_1991,N_102,N_640);
nand U1992 (N_1992,N_407,N_922);
nand U1993 (N_1993,N_762,N_134);
and U1994 (N_1994,N_482,N_43);
nor U1995 (N_1995,N_765,N_724);
or U1996 (N_1996,N_42,N_753);
nand U1997 (N_1997,N_175,N_869);
nand U1998 (N_1998,N_135,N_326);
and U1999 (N_1999,N_835,N_201);
and U2000 (N_2000,N_1940,N_1474);
nor U2001 (N_2001,N_1883,N_1828);
nand U2002 (N_2002,N_1979,N_1838);
and U2003 (N_2003,N_1622,N_1157);
or U2004 (N_2004,N_1894,N_1261);
nand U2005 (N_2005,N_1668,N_1025);
nor U2006 (N_2006,N_1341,N_1333);
nor U2007 (N_2007,N_1275,N_1397);
nand U2008 (N_2008,N_1877,N_1980);
nor U2009 (N_2009,N_1825,N_1430);
or U2010 (N_2010,N_1888,N_1370);
nand U2011 (N_2011,N_1433,N_1133);
nand U2012 (N_2012,N_1608,N_1308);
nand U2013 (N_2013,N_1209,N_1478);
or U2014 (N_2014,N_1052,N_1540);
or U2015 (N_2015,N_1935,N_1394);
or U2016 (N_2016,N_1956,N_1099);
and U2017 (N_2017,N_1497,N_1039);
and U2018 (N_2018,N_1444,N_1831);
nand U2019 (N_2019,N_1607,N_1896);
nand U2020 (N_2020,N_1899,N_1205);
nand U2021 (N_2021,N_1734,N_1619);
nand U2022 (N_2022,N_1794,N_1897);
nor U2023 (N_2023,N_1826,N_1097);
or U2024 (N_2024,N_1530,N_1024);
or U2025 (N_2025,N_1799,N_1732);
nor U2026 (N_2026,N_1775,N_1447);
nor U2027 (N_2027,N_1198,N_1148);
nor U2028 (N_2028,N_1352,N_1919);
or U2029 (N_2029,N_1698,N_1222);
or U2030 (N_2030,N_1448,N_1504);
or U2031 (N_2031,N_1297,N_1639);
nor U2032 (N_2032,N_1944,N_1191);
nor U2033 (N_2033,N_1957,N_1458);
nand U2034 (N_2034,N_1455,N_1230);
nor U2035 (N_2035,N_1911,N_1409);
nand U2036 (N_2036,N_1118,N_1836);
or U2037 (N_2037,N_1364,N_1131);
nand U2038 (N_2038,N_1396,N_1660);
or U2039 (N_2039,N_1724,N_1163);
nand U2040 (N_2040,N_1987,N_1225);
xnor U2041 (N_2041,N_1250,N_1853);
or U2042 (N_2042,N_1889,N_1511);
nor U2043 (N_2043,N_1598,N_1676);
or U2044 (N_2044,N_1968,N_1087);
and U2045 (N_2045,N_1164,N_1907);
and U2046 (N_2046,N_1064,N_1545);
xor U2047 (N_2047,N_1602,N_1927);
or U2048 (N_2048,N_1730,N_1757);
nor U2049 (N_2049,N_1151,N_1477);
nand U2050 (N_2050,N_1938,N_1103);
nor U2051 (N_2051,N_1976,N_1638);
and U2052 (N_2052,N_1606,N_1385);
nand U2053 (N_2053,N_1661,N_1324);
and U2054 (N_2054,N_1130,N_1321);
and U2055 (N_2055,N_1900,N_1780);
or U2056 (N_2056,N_1658,N_1193);
or U2057 (N_2057,N_1013,N_1053);
nor U2058 (N_2058,N_1588,N_1147);
and U2059 (N_2059,N_1893,N_1363);
and U2060 (N_2060,N_1247,N_1177);
nor U2061 (N_2061,N_1578,N_1381);
nand U2062 (N_2062,N_1281,N_1837);
nand U2063 (N_2063,N_1008,N_1467);
nand U2064 (N_2064,N_1549,N_1641);
or U2065 (N_2065,N_1821,N_1946);
nor U2066 (N_2066,N_1531,N_1055);
xnor U2067 (N_2067,N_1128,N_1279);
nand U2068 (N_2068,N_1594,N_1239);
xnor U2069 (N_2069,N_1366,N_1743);
nor U2070 (N_2070,N_1656,N_1375);
and U2071 (N_2071,N_1400,N_1180);
nand U2072 (N_2072,N_1586,N_1206);
nand U2073 (N_2073,N_1993,N_1390);
and U2074 (N_2074,N_1604,N_1521);
or U2075 (N_2075,N_1937,N_1181);
nand U2076 (N_2076,N_1078,N_1716);
nor U2077 (N_2077,N_1288,N_1959);
or U2078 (N_2078,N_1355,N_1923);
or U2079 (N_2079,N_1655,N_1582);
nor U2080 (N_2080,N_1751,N_1867);
nand U2081 (N_2081,N_1871,N_1762);
or U2082 (N_2082,N_1978,N_1334);
or U2083 (N_2083,N_1731,N_1260);
nor U2084 (N_2084,N_1313,N_1568);
or U2085 (N_2085,N_1007,N_1705);
and U2086 (N_2086,N_1590,N_1489);
nand U2087 (N_2087,N_1692,N_1989);
xor U2088 (N_2088,N_1422,N_1171);
nor U2089 (N_2089,N_1091,N_1718);
and U2090 (N_2090,N_1844,N_1139);
and U2091 (N_2091,N_1814,N_1016);
nor U2092 (N_2092,N_1067,N_1952);
nor U2093 (N_2093,N_1112,N_1041);
and U2094 (N_2094,N_1136,N_1964);
and U2095 (N_2095,N_1357,N_1028);
nand U2096 (N_2096,N_1450,N_1382);
nand U2097 (N_2097,N_1726,N_1537);
nand U2098 (N_2098,N_1977,N_1207);
or U2099 (N_2099,N_1124,N_1309);
nor U2100 (N_2100,N_1253,N_1407);
nor U2101 (N_2101,N_1150,N_1211);
nand U2102 (N_2102,N_1847,N_1083);
and U2103 (N_2103,N_1141,N_1519);
nor U2104 (N_2104,N_1476,N_1102);
nor U2105 (N_2105,N_1411,N_1542);
nor U2106 (N_2106,N_1802,N_1885);
nor U2107 (N_2107,N_1340,N_1872);
nand U2108 (N_2108,N_1713,N_1882);
or U2109 (N_2109,N_1930,N_1566);
or U2110 (N_2110,N_1416,N_1452);
or U2111 (N_2111,N_1522,N_1190);
or U2112 (N_2112,N_1833,N_1966);
nand U2113 (N_2113,N_1328,N_1246);
and U2114 (N_2114,N_1969,N_1256);
nand U2115 (N_2115,N_1307,N_1753);
and U2116 (N_2116,N_1574,N_1868);
nor U2117 (N_2117,N_1983,N_1495);
or U2118 (N_2118,N_1787,N_1525);
nand U2119 (N_2119,N_1264,N_1415);
nand U2120 (N_2120,N_1740,N_1453);
or U2121 (N_2121,N_1406,N_1999);
or U2122 (N_2122,N_1388,N_1673);
nor U2123 (N_2123,N_1675,N_1047);
or U2124 (N_2124,N_1173,N_1902);
and U2125 (N_2125,N_1647,N_1581);
nand U2126 (N_2126,N_1842,N_1955);
and U2127 (N_2127,N_1305,N_1565);
and U2128 (N_2128,N_1258,N_1652);
and U2129 (N_2129,N_1817,N_1270);
nand U2130 (N_2130,N_1903,N_1104);
nor U2131 (N_2131,N_1696,N_1295);
and U2132 (N_2132,N_1096,N_1666);
nor U2133 (N_2133,N_1241,N_1348);
nand U2134 (N_2134,N_1315,N_1482);
nor U2135 (N_2135,N_1697,N_1689);
or U2136 (N_2136,N_1789,N_1040);
or U2137 (N_2137,N_1851,N_1600);
nand U2138 (N_2138,N_1259,N_1709);
nor U2139 (N_2139,N_1304,N_1018);
nor U2140 (N_2140,N_1353,N_1459);
nor U2141 (N_2141,N_1142,N_1000);
and U2142 (N_2142,N_1446,N_1950);
xor U2143 (N_2143,N_1630,N_1123);
nand U2144 (N_2144,N_1928,N_1788);
xnor U2145 (N_2145,N_1371,N_1832);
nand U2146 (N_2146,N_1332,N_1918);
nand U2147 (N_2147,N_1419,N_1032);
nor U2148 (N_2148,N_1350,N_1351);
and U2149 (N_2149,N_1764,N_1684);
nor U2150 (N_2150,N_1856,N_1105);
nor U2151 (N_2151,N_1687,N_1564);
and U2152 (N_2152,N_1187,N_1524);
or U2153 (N_2153,N_1514,N_1202);
or U2154 (N_2154,N_1634,N_1505);
nand U2155 (N_2155,N_1553,N_1848);
nand U2156 (N_2156,N_1529,N_1644);
or U2157 (N_2157,N_1575,N_1006);
or U2158 (N_2158,N_1109,N_1806);
nand U2159 (N_2159,N_1895,N_1958);
and U2160 (N_2160,N_1621,N_1266);
nand U2161 (N_2161,N_1162,N_1170);
nor U2162 (N_2162,N_1801,N_1428);
nand U2163 (N_2163,N_1890,N_1046);
or U2164 (N_2164,N_1010,N_1318);
or U2165 (N_2165,N_1770,N_1820);
and U2166 (N_2166,N_1558,N_1991);
xnor U2167 (N_2167,N_1242,N_1084);
nor U2168 (N_2168,N_1143,N_1862);
nor U2169 (N_2169,N_1500,N_1175);
nand U2170 (N_2170,N_1042,N_1376);
or U2171 (N_2171,N_1601,N_1921);
or U2172 (N_2172,N_1733,N_1792);
nor U2173 (N_2173,N_1997,N_1249);
and U2174 (N_2174,N_1533,N_1784);
and U2175 (N_2175,N_1998,N_1485);
or U2176 (N_2176,N_1822,N_1922);
and U2177 (N_2177,N_1145,N_1917);
and U2178 (N_2178,N_1613,N_1996);
and U2179 (N_2179,N_1985,N_1612);
or U2180 (N_2180,N_1057,N_1404);
or U2181 (N_2181,N_1300,N_1059);
or U2182 (N_2182,N_1589,N_1272);
and U2183 (N_2183,N_1651,N_1329);
and U2184 (N_2184,N_1383,N_1569);
nor U2185 (N_2185,N_1238,N_1912);
or U2186 (N_2186,N_1475,N_1701);
and U2187 (N_2187,N_1081,N_1101);
nand U2188 (N_2188,N_1271,N_1073);
nand U2189 (N_2189,N_1345,N_1981);
and U2190 (N_2190,N_1255,N_1623);
nand U2191 (N_2191,N_1033,N_1113);
and U2192 (N_2192,N_1712,N_1335);
or U2193 (N_2193,N_1653,N_1779);
nor U2194 (N_2194,N_1532,N_1146);
nor U2195 (N_2195,N_1793,N_1869);
nand U2196 (N_2196,N_1798,N_1050);
nor U2197 (N_2197,N_1036,N_1429);
or U2198 (N_2198,N_1481,N_1484);
or U2199 (N_2199,N_1359,N_1681);
and U2200 (N_2200,N_1325,N_1449);
or U2201 (N_2201,N_1274,N_1369);
and U2202 (N_2202,N_1499,N_1116);
nor U2203 (N_2203,N_1461,N_1488);
or U2204 (N_2204,N_1294,N_1306);
nand U2205 (N_2205,N_1496,N_1849);
or U2206 (N_2206,N_1631,N_1664);
or U2207 (N_2207,N_1587,N_1115);
nand U2208 (N_2208,N_1554,N_1001);
and U2209 (N_2209,N_1559,N_1597);
or U2210 (N_2210,N_1389,N_1337);
nor U2211 (N_2211,N_1188,N_1766);
nor U2212 (N_2212,N_1437,N_1074);
nor U2213 (N_2213,N_1346,N_1616);
nand U2214 (N_2214,N_1859,N_1121);
and U2215 (N_2215,N_1570,N_1031);
nand U2216 (N_2216,N_1649,N_1417);
nor U2217 (N_2217,N_1509,N_1440);
or U2218 (N_2218,N_1772,N_1424);
and U2219 (N_2219,N_1700,N_1551);
and U2220 (N_2220,N_1626,N_1088);
and U2221 (N_2221,N_1702,N_1614);
and U2222 (N_2222,N_1159,N_1547);
nand U2223 (N_2223,N_1398,N_1878);
or U2224 (N_2224,N_1541,N_1576);
or U2225 (N_2225,N_1285,N_1536);
or U2226 (N_2226,N_1796,N_1876);
nand U2227 (N_2227,N_1227,N_1487);
and U2228 (N_2228,N_1265,N_1322);
or U2229 (N_2229,N_1517,N_1508);
and U2230 (N_2230,N_1665,N_1286);
nand U2231 (N_2231,N_1377,N_1808);
nand U2232 (N_2232,N_1117,N_1257);
or U2233 (N_2233,N_1829,N_1620);
nor U2234 (N_2234,N_1319,N_1768);
or U2235 (N_2235,N_1004,N_1093);
and U2236 (N_2236,N_1423,N_1195);
or U2237 (N_2237,N_1220,N_1617);
or U2238 (N_2238,N_1072,N_1534);
and U2239 (N_2239,N_1628,N_1967);
or U2240 (N_2240,N_1326,N_1431);
nand U2241 (N_2241,N_1401,N_1816);
and U2242 (N_2242,N_1178,N_1526);
nor U2243 (N_2243,N_1254,N_1323);
or U2244 (N_2244,N_1672,N_1462);
or U2245 (N_2245,N_1427,N_1790);
or U2246 (N_2246,N_1432,N_1506);
nor U2247 (N_2247,N_1282,N_1627);
or U2248 (N_2248,N_1925,N_1502);
nor U2249 (N_2249,N_1212,N_1126);
xnor U2250 (N_2250,N_1169,N_1637);
nor U2251 (N_2251,N_1068,N_1722);
and U2252 (N_2252,N_1642,N_1374);
or U2253 (N_2253,N_1695,N_1208);
nor U2254 (N_2254,N_1807,N_1441);
nor U2255 (N_2255,N_1786,N_1715);
nor U2256 (N_2256,N_1906,N_1562);
and U2257 (N_2257,N_1943,N_1296);
or U2258 (N_2258,N_1717,N_1009);
and U2259 (N_2259,N_1111,N_1035);
nand U2260 (N_2260,N_1800,N_1420);
and U2261 (N_2261,N_1216,N_1579);
or U2262 (N_2262,N_1603,N_1284);
nand U2263 (N_2263,N_1763,N_1122);
nor U2264 (N_2264,N_1491,N_1120);
nor U2265 (N_2265,N_1435,N_1823);
xnor U2266 (N_2266,N_1916,N_1092);
xor U2267 (N_2267,N_1543,N_1742);
xor U2268 (N_2268,N_1683,N_1913);
nand U2269 (N_2269,N_1804,N_1992);
or U2270 (N_2270,N_1015,N_1386);
xnor U2271 (N_2271,N_1045,N_1290);
nor U2272 (N_2272,N_1314,N_1330);
nor U2273 (N_2273,N_1677,N_1303);
nor U2274 (N_2274,N_1791,N_1454);
or U2275 (N_2275,N_1707,N_1861);
nand U2276 (N_2276,N_1942,N_1155);
or U2277 (N_2277,N_1984,N_1931);
nor U2278 (N_2278,N_1745,N_1043);
or U2279 (N_2279,N_1368,N_1812);
xor U2280 (N_2280,N_1214,N_1086);
nand U2281 (N_2281,N_1563,N_1744);
nor U2282 (N_2282,N_1240,N_1739);
nor U2283 (N_2283,N_1469,N_1669);
or U2284 (N_2284,N_1645,N_1372);
nor U2285 (N_2285,N_1005,N_1395);
nand U2286 (N_2286,N_1012,N_1591);
nor U2287 (N_2287,N_1908,N_1926);
xor U2288 (N_2288,N_1197,N_1356);
nand U2289 (N_2289,N_1749,N_1593);
and U2290 (N_2290,N_1291,N_1165);
and U2291 (N_2291,N_1228,N_1699);
and U2292 (N_2292,N_1605,N_1049);
nor U2293 (N_2293,N_1960,N_1134);
nand U2294 (N_2294,N_1557,N_1244);
and U2295 (N_2295,N_1234,N_1855);
and U2296 (N_2296,N_1609,N_1125);
and U2297 (N_2297,N_1203,N_1152);
nor U2298 (N_2298,N_1571,N_1172);
and U2299 (N_2299,N_1034,N_1972);
or U2300 (N_2300,N_1223,N_1338);
nor U2301 (N_2301,N_1741,N_1640);
nand U2302 (N_2302,N_1954,N_1166);
and U2303 (N_2303,N_1161,N_1596);
and U2304 (N_2304,N_1480,N_1472);
or U2305 (N_2305,N_1881,N_1752);
nand U2306 (N_2306,N_1845,N_1347);
and U2307 (N_2307,N_1344,N_1479);
nand U2308 (N_2308,N_1443,N_1235);
or U2309 (N_2309,N_1378,N_1199);
nand U2310 (N_2310,N_1466,N_1523);
nand U2311 (N_2311,N_1457,N_1327);
nand U2312 (N_2312,N_1367,N_1463);
nor U2313 (N_2313,N_1445,N_1657);
nand U2314 (N_2314,N_1160,N_1965);
or U2315 (N_2315,N_1694,N_1464);
and U2316 (N_2316,N_1425,N_1183);
nand U2317 (N_2317,N_1948,N_1988);
nor U2318 (N_2318,N_1438,N_1904);
nor U2319 (N_2319,N_1029,N_1158);
nor U2320 (N_2320,N_1129,N_1555);
or U2321 (N_2321,N_1107,N_1650);
or U2322 (N_2322,N_1060,N_1824);
and U2323 (N_2323,N_1611,N_1750);
nor U2324 (N_2324,N_1098,N_1301);
and U2325 (N_2325,N_1830,N_1135);
or U2326 (N_2326,N_1224,N_1292);
nor U2327 (N_2327,N_1358,N_1773);
and U2328 (N_2328,N_1269,N_1391);
nand U2329 (N_2329,N_1215,N_1439);
and U2330 (N_2330,N_1251,N_1030);
and U2331 (N_2331,N_1809,N_1879);
nor U2332 (N_2332,N_1818,N_1819);
nand U2333 (N_2333,N_1920,N_1778);
nand U2334 (N_2334,N_1317,N_1137);
and U2335 (N_2335,N_1293,N_1834);
nand U2336 (N_2336,N_1302,N_1725);
nand U2337 (N_2337,N_1729,N_1515);
and U2338 (N_2338,N_1027,N_1690);
nor U2339 (N_2339,N_1827,N_1548);
nor U2340 (N_2340,N_1414,N_1312);
and U2341 (N_2341,N_1217,N_1805);
and U2342 (N_2342,N_1840,N_1077);
nand U2343 (N_2343,N_1268,N_1755);
nand U2344 (N_2344,N_1512,N_1520);
and U2345 (N_2345,N_1528,N_1154);
or U2346 (N_2346,N_1156,N_1560);
or U2347 (N_2347,N_1237,N_1310);
and U2348 (N_2348,N_1970,N_1192);
or U2349 (N_2349,N_1280,N_1076);
nor U2350 (N_2350,N_1648,N_1636);
nand U2351 (N_2351,N_1624,N_1311);
nand U2352 (N_2352,N_1070,N_1756);
and U2353 (N_2353,N_1561,N_1864);
or U2354 (N_2354,N_1783,N_1552);
nor U2355 (N_2355,N_1580,N_1379);
nor U2356 (N_2356,N_1094,N_1905);
nor U2357 (N_2357,N_1720,N_1287);
or U2358 (N_2358,N_1493,N_1901);
nand U2359 (N_2359,N_1719,N_1962);
or U2360 (N_2360,N_1392,N_1408);
or U2361 (N_2361,N_1380,N_1153);
xnor U2362 (N_2362,N_1174,N_1693);
and U2363 (N_2363,N_1754,N_1982);
nor U2364 (N_2364,N_1610,N_1516);
nand U2365 (N_2365,N_1573,N_1785);
nand U2366 (N_2366,N_1852,N_1513);
or U2367 (N_2367,N_1470,N_1884);
nand U2368 (N_2368,N_1518,N_1854);
nor U2369 (N_2369,N_1510,N_1674);
or U2370 (N_2370,N_1846,N_1085);
and U2371 (N_2371,N_1393,N_1267);
nand U2372 (N_2372,N_1184,N_1289);
nand U2373 (N_2373,N_1201,N_1194);
nand U2374 (N_2374,N_1442,N_1728);
and U2375 (N_2375,N_1951,N_1063);
nor U2376 (N_2376,N_1706,N_1841);
or U2377 (N_2377,N_1646,N_1932);
and U2378 (N_2378,N_1662,N_1874);
and U2379 (N_2379,N_1021,N_1746);
nand U2380 (N_2380,N_1054,N_1373);
nand U2381 (N_2381,N_1858,N_1069);
or U2382 (N_2382,N_1760,N_1670);
and U2383 (N_2383,N_1252,N_1738);
or U2384 (N_2384,N_1185,N_1051);
or U2385 (N_2385,N_1583,N_1248);
nor U2386 (N_2386,N_1119,N_1200);
nand U2387 (N_2387,N_1402,N_1949);
and U2388 (N_2388,N_1410,N_1618);
or U2389 (N_2389,N_1168,N_1663);
and U2390 (N_2390,N_1671,N_1711);
or U2391 (N_2391,N_1298,N_1686);
nor U2392 (N_2392,N_1219,N_1132);
and U2393 (N_2393,N_1079,N_1863);
or U2394 (N_2394,N_1986,N_1704);
nor U2395 (N_2395,N_1941,N_1062);
and U2396 (N_2396,N_1924,N_1167);
nor U2397 (N_2397,N_1436,N_1492);
nand U2398 (N_2398,N_1546,N_1934);
or U2399 (N_2399,N_1995,N_1909);
nor U2400 (N_2400,N_1795,N_1811);
nor U2401 (N_2401,N_1138,N_1737);
and U2402 (N_2402,N_1262,N_1947);
or U2403 (N_2403,N_1232,N_1245);
or U2404 (N_2404,N_1887,N_1736);
or U2405 (N_2405,N_1460,N_1735);
nand U2406 (N_2406,N_1221,N_1362);
nand U2407 (N_2407,N_1629,N_1680);
and U2408 (N_2408,N_1231,N_1213);
and U2409 (N_2409,N_1572,N_1810);
and U2410 (N_2410,N_1186,N_1860);
or U2411 (N_2411,N_1149,N_1781);
and U2412 (N_2412,N_1038,N_1592);
or U2413 (N_2413,N_1144,N_1090);
or U2414 (N_2414,N_1761,N_1865);
nand U2415 (N_2415,N_1468,N_1048);
nor U2416 (N_2416,N_1490,N_1963);
nand U2417 (N_2417,N_1014,N_1421);
nand U2418 (N_2418,N_1782,N_1503);
nor U2419 (N_2419,N_1933,N_1365);
nor U2420 (N_2420,N_1774,N_1486);
nor U2421 (N_2421,N_1498,N_1803);
and U2422 (N_2422,N_1011,N_1507);
or U2423 (N_2423,N_1273,N_1339);
nor U2424 (N_2424,N_1065,N_1003);
or U2425 (N_2425,N_1095,N_1434);
and U2426 (N_2426,N_1797,N_1567);
nand U2427 (N_2427,N_1815,N_1667);
nand U2428 (N_2428,N_1813,N_1850);
and U2429 (N_2429,N_1679,N_1678);
or U2430 (N_2430,N_1714,N_1387);
or U2431 (N_2431,N_1975,N_1839);
nor U2432 (N_2432,N_1140,N_1723);
or U2433 (N_2433,N_1179,N_1451);
or U2434 (N_2434,N_1915,N_1539);
nand U2435 (N_2435,N_1721,N_1413);
and U2436 (N_2436,N_1577,N_1914);
and U2437 (N_2437,N_1236,N_1767);
nand U2438 (N_2438,N_1776,N_1759);
nor U2439 (N_2439,N_1974,N_1929);
nand U2440 (N_2440,N_1020,N_1361);
nand U2441 (N_2441,N_1973,N_1002);
nand U2442 (N_2442,N_1058,N_1710);
nand U2443 (N_2443,N_1108,N_1843);
xnor U2444 (N_2444,N_1777,N_1691);
nand U2445 (N_2445,N_1218,N_1682);
nand U2446 (N_2446,N_1654,N_1659);
or U2447 (N_2447,N_1360,N_1910);
or U2448 (N_2448,N_1089,N_1688);
nor U2449 (N_2449,N_1277,N_1866);
nand U2450 (N_2450,N_1535,N_1873);
or U2451 (N_2451,N_1892,N_1643);
and U2452 (N_2452,N_1875,N_1022);
and U2453 (N_2453,N_1399,N_1870);
or U2454 (N_2454,N_1384,N_1456);
or U2455 (N_2455,N_1342,N_1615);
nand U2456 (N_2456,N_1538,N_1316);
nor U2457 (N_2457,N_1599,N_1061);
nor U2458 (N_2458,N_1465,N_1758);
nand U2459 (N_2459,N_1080,N_1747);
nand U2460 (N_2460,N_1066,N_1765);
nor U2461 (N_2461,N_1204,N_1343);
or U2462 (N_2462,N_1994,N_1418);
or U2463 (N_2463,N_1075,N_1501);
nor U2464 (N_2464,N_1483,N_1727);
and U2465 (N_2465,N_1494,N_1176);
and U2466 (N_2466,N_1110,N_1835);
or U2467 (N_2467,N_1961,N_1189);
and U2468 (N_2468,N_1403,N_1771);
or U2469 (N_2469,N_1898,N_1331);
nand U2470 (N_2470,N_1037,N_1336);
nand U2471 (N_2471,N_1748,N_1100);
or U2472 (N_2472,N_1886,N_1017);
nand U2473 (N_2473,N_1044,N_1114);
or U2474 (N_2474,N_1584,N_1527);
or U2475 (N_2475,N_1550,N_1595);
nor U2476 (N_2476,N_1026,N_1019);
or U2477 (N_2477,N_1703,N_1182);
nand U2478 (N_2478,N_1106,N_1229);
nor U2479 (N_2479,N_1632,N_1880);
nor U2480 (N_2480,N_1891,N_1971);
nand U2481 (N_2481,N_1625,N_1936);
or U2482 (N_2482,N_1071,N_1243);
or U2483 (N_2483,N_1226,N_1210);
nand U2484 (N_2484,N_1233,N_1056);
or U2485 (N_2485,N_1405,N_1635);
nor U2486 (N_2486,N_1283,N_1708);
or U2487 (N_2487,N_1556,N_1685);
nand U2488 (N_2488,N_1263,N_1354);
nor U2489 (N_2489,N_1473,N_1953);
nand U2490 (N_2490,N_1349,N_1544);
or U2491 (N_2491,N_1990,N_1412);
or U2492 (N_2492,N_1127,N_1196);
xor U2493 (N_2493,N_1857,N_1633);
nand U2494 (N_2494,N_1426,N_1276);
and U2495 (N_2495,N_1023,N_1082);
and U2496 (N_2496,N_1939,N_1471);
or U2497 (N_2497,N_1945,N_1278);
or U2498 (N_2498,N_1585,N_1299);
and U2499 (N_2499,N_1320,N_1769);
or U2500 (N_2500,N_1731,N_1324);
nor U2501 (N_2501,N_1313,N_1336);
or U2502 (N_2502,N_1033,N_1323);
nor U2503 (N_2503,N_1843,N_1774);
nand U2504 (N_2504,N_1784,N_1704);
and U2505 (N_2505,N_1388,N_1617);
or U2506 (N_2506,N_1782,N_1216);
xnor U2507 (N_2507,N_1574,N_1907);
or U2508 (N_2508,N_1537,N_1662);
nor U2509 (N_2509,N_1699,N_1269);
and U2510 (N_2510,N_1774,N_1212);
and U2511 (N_2511,N_1063,N_1390);
or U2512 (N_2512,N_1323,N_1979);
nor U2513 (N_2513,N_1617,N_1991);
or U2514 (N_2514,N_1566,N_1984);
and U2515 (N_2515,N_1239,N_1285);
nor U2516 (N_2516,N_1896,N_1198);
and U2517 (N_2517,N_1747,N_1697);
and U2518 (N_2518,N_1168,N_1807);
nor U2519 (N_2519,N_1887,N_1498);
nand U2520 (N_2520,N_1643,N_1966);
or U2521 (N_2521,N_1633,N_1371);
nor U2522 (N_2522,N_1418,N_1993);
nor U2523 (N_2523,N_1138,N_1427);
and U2524 (N_2524,N_1445,N_1520);
or U2525 (N_2525,N_1115,N_1165);
nand U2526 (N_2526,N_1804,N_1740);
and U2527 (N_2527,N_1240,N_1668);
or U2528 (N_2528,N_1485,N_1839);
nor U2529 (N_2529,N_1949,N_1597);
or U2530 (N_2530,N_1236,N_1899);
or U2531 (N_2531,N_1357,N_1580);
and U2532 (N_2532,N_1286,N_1605);
nand U2533 (N_2533,N_1141,N_1277);
or U2534 (N_2534,N_1421,N_1925);
and U2535 (N_2535,N_1142,N_1127);
nor U2536 (N_2536,N_1699,N_1615);
nor U2537 (N_2537,N_1479,N_1063);
nor U2538 (N_2538,N_1438,N_1177);
nor U2539 (N_2539,N_1641,N_1492);
or U2540 (N_2540,N_1801,N_1761);
or U2541 (N_2541,N_1538,N_1869);
xor U2542 (N_2542,N_1498,N_1506);
and U2543 (N_2543,N_1748,N_1496);
and U2544 (N_2544,N_1995,N_1879);
xor U2545 (N_2545,N_1279,N_1483);
and U2546 (N_2546,N_1790,N_1561);
nor U2547 (N_2547,N_1708,N_1044);
nor U2548 (N_2548,N_1265,N_1210);
and U2549 (N_2549,N_1421,N_1259);
nor U2550 (N_2550,N_1121,N_1060);
nor U2551 (N_2551,N_1009,N_1025);
and U2552 (N_2552,N_1716,N_1291);
nand U2553 (N_2553,N_1980,N_1907);
nand U2554 (N_2554,N_1418,N_1636);
nor U2555 (N_2555,N_1153,N_1700);
nor U2556 (N_2556,N_1036,N_1332);
or U2557 (N_2557,N_1290,N_1224);
nor U2558 (N_2558,N_1169,N_1639);
and U2559 (N_2559,N_1584,N_1757);
nand U2560 (N_2560,N_1971,N_1354);
and U2561 (N_2561,N_1971,N_1492);
or U2562 (N_2562,N_1560,N_1905);
and U2563 (N_2563,N_1883,N_1240);
or U2564 (N_2564,N_1106,N_1024);
or U2565 (N_2565,N_1919,N_1000);
and U2566 (N_2566,N_1425,N_1745);
and U2567 (N_2567,N_1337,N_1905);
or U2568 (N_2568,N_1671,N_1817);
nand U2569 (N_2569,N_1646,N_1875);
or U2570 (N_2570,N_1431,N_1638);
and U2571 (N_2571,N_1928,N_1855);
and U2572 (N_2572,N_1254,N_1585);
and U2573 (N_2573,N_1374,N_1559);
or U2574 (N_2574,N_1739,N_1911);
and U2575 (N_2575,N_1414,N_1722);
xnor U2576 (N_2576,N_1459,N_1962);
nand U2577 (N_2577,N_1724,N_1572);
and U2578 (N_2578,N_1298,N_1929);
nand U2579 (N_2579,N_1388,N_1766);
and U2580 (N_2580,N_1726,N_1684);
nand U2581 (N_2581,N_1730,N_1116);
or U2582 (N_2582,N_1291,N_1489);
or U2583 (N_2583,N_1452,N_1946);
nand U2584 (N_2584,N_1966,N_1905);
nand U2585 (N_2585,N_1533,N_1944);
or U2586 (N_2586,N_1915,N_1837);
nor U2587 (N_2587,N_1927,N_1547);
nand U2588 (N_2588,N_1084,N_1092);
and U2589 (N_2589,N_1261,N_1610);
or U2590 (N_2590,N_1080,N_1003);
nand U2591 (N_2591,N_1165,N_1145);
nor U2592 (N_2592,N_1252,N_1824);
nor U2593 (N_2593,N_1694,N_1654);
xor U2594 (N_2594,N_1030,N_1392);
and U2595 (N_2595,N_1048,N_1000);
nand U2596 (N_2596,N_1087,N_1348);
nor U2597 (N_2597,N_1178,N_1286);
nor U2598 (N_2598,N_1958,N_1047);
nand U2599 (N_2599,N_1748,N_1858);
nor U2600 (N_2600,N_1396,N_1944);
nand U2601 (N_2601,N_1984,N_1130);
nor U2602 (N_2602,N_1718,N_1617);
and U2603 (N_2603,N_1770,N_1718);
or U2604 (N_2604,N_1599,N_1122);
nor U2605 (N_2605,N_1326,N_1178);
nand U2606 (N_2606,N_1889,N_1478);
nand U2607 (N_2607,N_1273,N_1866);
and U2608 (N_2608,N_1499,N_1045);
nor U2609 (N_2609,N_1719,N_1310);
nand U2610 (N_2610,N_1638,N_1818);
nand U2611 (N_2611,N_1466,N_1994);
xor U2612 (N_2612,N_1155,N_1076);
and U2613 (N_2613,N_1431,N_1113);
and U2614 (N_2614,N_1125,N_1393);
or U2615 (N_2615,N_1589,N_1897);
and U2616 (N_2616,N_1516,N_1688);
nor U2617 (N_2617,N_1892,N_1445);
xor U2618 (N_2618,N_1486,N_1533);
and U2619 (N_2619,N_1302,N_1505);
and U2620 (N_2620,N_1702,N_1746);
or U2621 (N_2621,N_1030,N_1497);
or U2622 (N_2622,N_1369,N_1480);
xor U2623 (N_2623,N_1878,N_1339);
nand U2624 (N_2624,N_1496,N_1845);
nor U2625 (N_2625,N_1136,N_1846);
nor U2626 (N_2626,N_1808,N_1838);
nand U2627 (N_2627,N_1475,N_1990);
nand U2628 (N_2628,N_1580,N_1751);
nor U2629 (N_2629,N_1480,N_1620);
nand U2630 (N_2630,N_1002,N_1758);
or U2631 (N_2631,N_1608,N_1066);
and U2632 (N_2632,N_1699,N_1511);
xnor U2633 (N_2633,N_1949,N_1598);
or U2634 (N_2634,N_1632,N_1448);
nand U2635 (N_2635,N_1534,N_1809);
or U2636 (N_2636,N_1012,N_1701);
nand U2637 (N_2637,N_1366,N_1012);
nand U2638 (N_2638,N_1467,N_1106);
nand U2639 (N_2639,N_1020,N_1390);
nand U2640 (N_2640,N_1208,N_1940);
nand U2641 (N_2641,N_1943,N_1322);
or U2642 (N_2642,N_1503,N_1847);
and U2643 (N_2643,N_1974,N_1101);
or U2644 (N_2644,N_1236,N_1158);
nor U2645 (N_2645,N_1555,N_1659);
or U2646 (N_2646,N_1969,N_1147);
nand U2647 (N_2647,N_1312,N_1576);
or U2648 (N_2648,N_1241,N_1772);
and U2649 (N_2649,N_1556,N_1971);
and U2650 (N_2650,N_1114,N_1771);
xor U2651 (N_2651,N_1596,N_1745);
or U2652 (N_2652,N_1042,N_1201);
or U2653 (N_2653,N_1754,N_1035);
and U2654 (N_2654,N_1039,N_1200);
and U2655 (N_2655,N_1160,N_1940);
nor U2656 (N_2656,N_1714,N_1470);
nand U2657 (N_2657,N_1093,N_1697);
or U2658 (N_2658,N_1307,N_1756);
and U2659 (N_2659,N_1271,N_1413);
and U2660 (N_2660,N_1260,N_1249);
nand U2661 (N_2661,N_1457,N_1723);
nand U2662 (N_2662,N_1388,N_1993);
or U2663 (N_2663,N_1178,N_1208);
and U2664 (N_2664,N_1780,N_1422);
nor U2665 (N_2665,N_1053,N_1450);
nor U2666 (N_2666,N_1773,N_1464);
and U2667 (N_2667,N_1045,N_1233);
and U2668 (N_2668,N_1173,N_1477);
or U2669 (N_2669,N_1939,N_1798);
and U2670 (N_2670,N_1131,N_1871);
nor U2671 (N_2671,N_1386,N_1134);
nand U2672 (N_2672,N_1630,N_1462);
and U2673 (N_2673,N_1018,N_1345);
and U2674 (N_2674,N_1246,N_1953);
xor U2675 (N_2675,N_1098,N_1779);
and U2676 (N_2676,N_1307,N_1721);
nor U2677 (N_2677,N_1719,N_1530);
and U2678 (N_2678,N_1918,N_1966);
nor U2679 (N_2679,N_1049,N_1533);
nand U2680 (N_2680,N_1764,N_1572);
nor U2681 (N_2681,N_1507,N_1589);
nor U2682 (N_2682,N_1594,N_1080);
nor U2683 (N_2683,N_1567,N_1785);
nand U2684 (N_2684,N_1666,N_1562);
and U2685 (N_2685,N_1491,N_1062);
nor U2686 (N_2686,N_1167,N_1620);
nor U2687 (N_2687,N_1485,N_1451);
or U2688 (N_2688,N_1206,N_1137);
nor U2689 (N_2689,N_1067,N_1737);
and U2690 (N_2690,N_1407,N_1274);
or U2691 (N_2691,N_1578,N_1659);
nor U2692 (N_2692,N_1508,N_1886);
and U2693 (N_2693,N_1721,N_1301);
or U2694 (N_2694,N_1376,N_1513);
nor U2695 (N_2695,N_1535,N_1502);
nand U2696 (N_2696,N_1969,N_1498);
nor U2697 (N_2697,N_1300,N_1880);
nor U2698 (N_2698,N_1621,N_1335);
nand U2699 (N_2699,N_1674,N_1295);
or U2700 (N_2700,N_1847,N_1711);
or U2701 (N_2701,N_1587,N_1469);
xor U2702 (N_2702,N_1116,N_1859);
or U2703 (N_2703,N_1369,N_1149);
or U2704 (N_2704,N_1654,N_1598);
nor U2705 (N_2705,N_1050,N_1341);
or U2706 (N_2706,N_1897,N_1844);
nand U2707 (N_2707,N_1455,N_1804);
nand U2708 (N_2708,N_1709,N_1459);
or U2709 (N_2709,N_1506,N_1996);
nand U2710 (N_2710,N_1075,N_1498);
and U2711 (N_2711,N_1533,N_1959);
or U2712 (N_2712,N_1164,N_1279);
and U2713 (N_2713,N_1229,N_1446);
nor U2714 (N_2714,N_1297,N_1355);
nor U2715 (N_2715,N_1259,N_1083);
and U2716 (N_2716,N_1181,N_1981);
nor U2717 (N_2717,N_1536,N_1542);
and U2718 (N_2718,N_1408,N_1553);
or U2719 (N_2719,N_1108,N_1543);
and U2720 (N_2720,N_1203,N_1855);
and U2721 (N_2721,N_1584,N_1689);
nand U2722 (N_2722,N_1654,N_1978);
nor U2723 (N_2723,N_1274,N_1559);
nand U2724 (N_2724,N_1835,N_1545);
and U2725 (N_2725,N_1225,N_1896);
nand U2726 (N_2726,N_1494,N_1192);
nand U2727 (N_2727,N_1525,N_1055);
nor U2728 (N_2728,N_1047,N_1625);
nor U2729 (N_2729,N_1315,N_1304);
or U2730 (N_2730,N_1647,N_1935);
nor U2731 (N_2731,N_1659,N_1791);
nor U2732 (N_2732,N_1962,N_1495);
xnor U2733 (N_2733,N_1050,N_1364);
or U2734 (N_2734,N_1450,N_1846);
and U2735 (N_2735,N_1297,N_1269);
or U2736 (N_2736,N_1304,N_1615);
nand U2737 (N_2737,N_1224,N_1484);
or U2738 (N_2738,N_1277,N_1313);
nand U2739 (N_2739,N_1077,N_1813);
xnor U2740 (N_2740,N_1383,N_1164);
nand U2741 (N_2741,N_1083,N_1792);
nor U2742 (N_2742,N_1486,N_1094);
or U2743 (N_2743,N_1983,N_1489);
or U2744 (N_2744,N_1552,N_1101);
nand U2745 (N_2745,N_1365,N_1636);
nor U2746 (N_2746,N_1054,N_1547);
nor U2747 (N_2747,N_1262,N_1072);
or U2748 (N_2748,N_1713,N_1522);
or U2749 (N_2749,N_1431,N_1117);
and U2750 (N_2750,N_1049,N_1846);
nand U2751 (N_2751,N_1967,N_1744);
nor U2752 (N_2752,N_1422,N_1228);
nor U2753 (N_2753,N_1681,N_1381);
or U2754 (N_2754,N_1824,N_1377);
nand U2755 (N_2755,N_1958,N_1064);
nand U2756 (N_2756,N_1915,N_1796);
nor U2757 (N_2757,N_1553,N_1439);
nand U2758 (N_2758,N_1255,N_1843);
xor U2759 (N_2759,N_1893,N_1444);
and U2760 (N_2760,N_1695,N_1623);
nor U2761 (N_2761,N_1234,N_1286);
or U2762 (N_2762,N_1999,N_1755);
or U2763 (N_2763,N_1880,N_1933);
or U2764 (N_2764,N_1386,N_1373);
or U2765 (N_2765,N_1793,N_1077);
nand U2766 (N_2766,N_1018,N_1169);
nor U2767 (N_2767,N_1843,N_1984);
and U2768 (N_2768,N_1914,N_1466);
nand U2769 (N_2769,N_1143,N_1960);
and U2770 (N_2770,N_1096,N_1799);
and U2771 (N_2771,N_1715,N_1108);
nor U2772 (N_2772,N_1248,N_1474);
or U2773 (N_2773,N_1463,N_1971);
or U2774 (N_2774,N_1901,N_1600);
nor U2775 (N_2775,N_1021,N_1603);
and U2776 (N_2776,N_1117,N_1184);
nand U2777 (N_2777,N_1689,N_1646);
or U2778 (N_2778,N_1764,N_1562);
and U2779 (N_2779,N_1510,N_1214);
nand U2780 (N_2780,N_1592,N_1321);
nor U2781 (N_2781,N_1332,N_1543);
nand U2782 (N_2782,N_1492,N_1793);
nor U2783 (N_2783,N_1725,N_1964);
nand U2784 (N_2784,N_1916,N_1302);
and U2785 (N_2785,N_1792,N_1529);
nand U2786 (N_2786,N_1127,N_1404);
nand U2787 (N_2787,N_1406,N_1967);
or U2788 (N_2788,N_1377,N_1093);
and U2789 (N_2789,N_1139,N_1433);
nor U2790 (N_2790,N_1035,N_1381);
nor U2791 (N_2791,N_1352,N_1864);
or U2792 (N_2792,N_1882,N_1704);
or U2793 (N_2793,N_1041,N_1192);
nor U2794 (N_2794,N_1432,N_1437);
or U2795 (N_2795,N_1269,N_1962);
or U2796 (N_2796,N_1982,N_1039);
nor U2797 (N_2797,N_1409,N_1416);
or U2798 (N_2798,N_1079,N_1716);
or U2799 (N_2799,N_1974,N_1165);
nand U2800 (N_2800,N_1760,N_1585);
nor U2801 (N_2801,N_1492,N_1987);
nor U2802 (N_2802,N_1647,N_1387);
nand U2803 (N_2803,N_1971,N_1790);
and U2804 (N_2804,N_1837,N_1641);
and U2805 (N_2805,N_1362,N_1274);
nor U2806 (N_2806,N_1593,N_1294);
and U2807 (N_2807,N_1479,N_1999);
or U2808 (N_2808,N_1207,N_1219);
or U2809 (N_2809,N_1719,N_1495);
or U2810 (N_2810,N_1913,N_1614);
or U2811 (N_2811,N_1740,N_1044);
or U2812 (N_2812,N_1476,N_1368);
and U2813 (N_2813,N_1653,N_1027);
and U2814 (N_2814,N_1754,N_1398);
nand U2815 (N_2815,N_1615,N_1015);
and U2816 (N_2816,N_1292,N_1971);
and U2817 (N_2817,N_1286,N_1213);
nor U2818 (N_2818,N_1611,N_1944);
and U2819 (N_2819,N_1945,N_1691);
nor U2820 (N_2820,N_1650,N_1255);
or U2821 (N_2821,N_1013,N_1113);
and U2822 (N_2822,N_1878,N_1328);
nor U2823 (N_2823,N_1031,N_1336);
or U2824 (N_2824,N_1291,N_1069);
or U2825 (N_2825,N_1370,N_1675);
and U2826 (N_2826,N_1138,N_1194);
and U2827 (N_2827,N_1755,N_1056);
nand U2828 (N_2828,N_1721,N_1068);
and U2829 (N_2829,N_1563,N_1378);
nor U2830 (N_2830,N_1798,N_1650);
xor U2831 (N_2831,N_1529,N_1947);
and U2832 (N_2832,N_1570,N_1531);
or U2833 (N_2833,N_1143,N_1159);
nand U2834 (N_2834,N_1295,N_1098);
nand U2835 (N_2835,N_1359,N_1494);
nor U2836 (N_2836,N_1231,N_1544);
nand U2837 (N_2837,N_1430,N_1526);
nor U2838 (N_2838,N_1122,N_1293);
or U2839 (N_2839,N_1378,N_1722);
and U2840 (N_2840,N_1290,N_1164);
nor U2841 (N_2841,N_1336,N_1502);
and U2842 (N_2842,N_1960,N_1916);
and U2843 (N_2843,N_1755,N_1665);
nor U2844 (N_2844,N_1324,N_1678);
xnor U2845 (N_2845,N_1625,N_1925);
and U2846 (N_2846,N_1502,N_1058);
nor U2847 (N_2847,N_1108,N_1848);
nand U2848 (N_2848,N_1083,N_1528);
and U2849 (N_2849,N_1566,N_1364);
nand U2850 (N_2850,N_1349,N_1464);
or U2851 (N_2851,N_1477,N_1907);
nand U2852 (N_2852,N_1059,N_1208);
and U2853 (N_2853,N_1775,N_1579);
or U2854 (N_2854,N_1713,N_1697);
nor U2855 (N_2855,N_1805,N_1439);
or U2856 (N_2856,N_1653,N_1061);
and U2857 (N_2857,N_1878,N_1245);
or U2858 (N_2858,N_1469,N_1623);
or U2859 (N_2859,N_1721,N_1659);
nor U2860 (N_2860,N_1633,N_1790);
nand U2861 (N_2861,N_1052,N_1130);
nor U2862 (N_2862,N_1145,N_1184);
nand U2863 (N_2863,N_1032,N_1244);
and U2864 (N_2864,N_1553,N_1131);
nor U2865 (N_2865,N_1959,N_1816);
and U2866 (N_2866,N_1821,N_1396);
or U2867 (N_2867,N_1134,N_1593);
and U2868 (N_2868,N_1486,N_1567);
and U2869 (N_2869,N_1998,N_1867);
nor U2870 (N_2870,N_1699,N_1477);
or U2871 (N_2871,N_1145,N_1304);
xor U2872 (N_2872,N_1526,N_1772);
nor U2873 (N_2873,N_1106,N_1196);
nor U2874 (N_2874,N_1335,N_1457);
nor U2875 (N_2875,N_1283,N_1662);
nor U2876 (N_2876,N_1652,N_1718);
and U2877 (N_2877,N_1470,N_1698);
xnor U2878 (N_2878,N_1727,N_1304);
nand U2879 (N_2879,N_1948,N_1610);
nand U2880 (N_2880,N_1917,N_1246);
and U2881 (N_2881,N_1138,N_1304);
xnor U2882 (N_2882,N_1337,N_1873);
or U2883 (N_2883,N_1924,N_1169);
nor U2884 (N_2884,N_1583,N_1737);
nand U2885 (N_2885,N_1346,N_1037);
or U2886 (N_2886,N_1057,N_1118);
or U2887 (N_2887,N_1600,N_1228);
nor U2888 (N_2888,N_1091,N_1269);
and U2889 (N_2889,N_1012,N_1853);
nand U2890 (N_2890,N_1253,N_1440);
and U2891 (N_2891,N_1526,N_1895);
nand U2892 (N_2892,N_1701,N_1065);
or U2893 (N_2893,N_1385,N_1973);
nor U2894 (N_2894,N_1441,N_1382);
and U2895 (N_2895,N_1273,N_1222);
nor U2896 (N_2896,N_1253,N_1272);
or U2897 (N_2897,N_1280,N_1273);
nor U2898 (N_2898,N_1944,N_1283);
or U2899 (N_2899,N_1172,N_1754);
or U2900 (N_2900,N_1178,N_1985);
and U2901 (N_2901,N_1853,N_1003);
nor U2902 (N_2902,N_1475,N_1420);
nor U2903 (N_2903,N_1101,N_1137);
nand U2904 (N_2904,N_1230,N_1078);
nand U2905 (N_2905,N_1030,N_1193);
xor U2906 (N_2906,N_1980,N_1463);
and U2907 (N_2907,N_1582,N_1206);
and U2908 (N_2908,N_1365,N_1193);
nand U2909 (N_2909,N_1053,N_1137);
or U2910 (N_2910,N_1196,N_1972);
or U2911 (N_2911,N_1042,N_1909);
nand U2912 (N_2912,N_1915,N_1567);
nand U2913 (N_2913,N_1717,N_1953);
or U2914 (N_2914,N_1107,N_1158);
and U2915 (N_2915,N_1552,N_1059);
nor U2916 (N_2916,N_1505,N_1721);
and U2917 (N_2917,N_1153,N_1420);
or U2918 (N_2918,N_1444,N_1549);
and U2919 (N_2919,N_1766,N_1773);
or U2920 (N_2920,N_1900,N_1627);
nor U2921 (N_2921,N_1787,N_1329);
or U2922 (N_2922,N_1720,N_1088);
nand U2923 (N_2923,N_1229,N_1533);
nand U2924 (N_2924,N_1000,N_1044);
or U2925 (N_2925,N_1131,N_1024);
nor U2926 (N_2926,N_1223,N_1065);
nor U2927 (N_2927,N_1783,N_1277);
nand U2928 (N_2928,N_1702,N_1421);
or U2929 (N_2929,N_1738,N_1867);
and U2930 (N_2930,N_1602,N_1070);
nand U2931 (N_2931,N_1684,N_1145);
nand U2932 (N_2932,N_1699,N_1563);
or U2933 (N_2933,N_1653,N_1812);
nor U2934 (N_2934,N_1427,N_1098);
or U2935 (N_2935,N_1297,N_1798);
nand U2936 (N_2936,N_1905,N_1018);
or U2937 (N_2937,N_1906,N_1733);
nor U2938 (N_2938,N_1272,N_1855);
or U2939 (N_2939,N_1837,N_1815);
and U2940 (N_2940,N_1959,N_1941);
nor U2941 (N_2941,N_1148,N_1900);
nand U2942 (N_2942,N_1900,N_1149);
or U2943 (N_2943,N_1898,N_1192);
or U2944 (N_2944,N_1293,N_1963);
and U2945 (N_2945,N_1946,N_1097);
and U2946 (N_2946,N_1364,N_1034);
nand U2947 (N_2947,N_1109,N_1553);
nand U2948 (N_2948,N_1561,N_1711);
nand U2949 (N_2949,N_1459,N_1556);
nand U2950 (N_2950,N_1655,N_1554);
or U2951 (N_2951,N_1645,N_1752);
nor U2952 (N_2952,N_1014,N_1971);
nand U2953 (N_2953,N_1202,N_1845);
or U2954 (N_2954,N_1846,N_1630);
and U2955 (N_2955,N_1449,N_1815);
nor U2956 (N_2956,N_1290,N_1488);
and U2957 (N_2957,N_1238,N_1057);
nor U2958 (N_2958,N_1150,N_1619);
and U2959 (N_2959,N_1111,N_1678);
or U2960 (N_2960,N_1672,N_1569);
nand U2961 (N_2961,N_1357,N_1088);
nand U2962 (N_2962,N_1200,N_1604);
nand U2963 (N_2963,N_1681,N_1048);
and U2964 (N_2964,N_1057,N_1017);
nor U2965 (N_2965,N_1386,N_1350);
or U2966 (N_2966,N_1016,N_1923);
and U2967 (N_2967,N_1376,N_1255);
nand U2968 (N_2968,N_1006,N_1804);
or U2969 (N_2969,N_1186,N_1361);
or U2970 (N_2970,N_1758,N_1609);
nor U2971 (N_2971,N_1385,N_1430);
nand U2972 (N_2972,N_1102,N_1950);
nor U2973 (N_2973,N_1893,N_1668);
or U2974 (N_2974,N_1274,N_1138);
nand U2975 (N_2975,N_1233,N_1789);
nor U2976 (N_2976,N_1688,N_1197);
nor U2977 (N_2977,N_1798,N_1043);
nand U2978 (N_2978,N_1154,N_1823);
and U2979 (N_2979,N_1321,N_1239);
and U2980 (N_2980,N_1406,N_1206);
or U2981 (N_2981,N_1067,N_1979);
nor U2982 (N_2982,N_1425,N_1943);
or U2983 (N_2983,N_1971,N_1296);
and U2984 (N_2984,N_1120,N_1780);
nor U2985 (N_2985,N_1426,N_1505);
nand U2986 (N_2986,N_1081,N_1236);
or U2987 (N_2987,N_1097,N_1315);
nor U2988 (N_2988,N_1822,N_1115);
nor U2989 (N_2989,N_1061,N_1912);
nor U2990 (N_2990,N_1813,N_1838);
nand U2991 (N_2991,N_1019,N_1563);
nor U2992 (N_2992,N_1402,N_1699);
nand U2993 (N_2993,N_1831,N_1472);
nor U2994 (N_2994,N_1933,N_1992);
and U2995 (N_2995,N_1869,N_1867);
or U2996 (N_2996,N_1719,N_1003);
or U2997 (N_2997,N_1562,N_1927);
or U2998 (N_2998,N_1773,N_1362);
xnor U2999 (N_2999,N_1019,N_1058);
nor U3000 (N_3000,N_2383,N_2813);
nand U3001 (N_3001,N_2764,N_2074);
or U3002 (N_3002,N_2785,N_2807);
and U3003 (N_3003,N_2523,N_2876);
nand U3004 (N_3004,N_2771,N_2806);
nand U3005 (N_3005,N_2061,N_2366);
and U3006 (N_3006,N_2069,N_2880);
and U3007 (N_3007,N_2335,N_2798);
and U3008 (N_3008,N_2904,N_2437);
and U3009 (N_3009,N_2739,N_2305);
or U3010 (N_3010,N_2923,N_2791);
nand U3011 (N_3011,N_2019,N_2992);
nor U3012 (N_3012,N_2847,N_2509);
nor U3013 (N_3013,N_2706,N_2021);
or U3014 (N_3014,N_2979,N_2529);
and U3015 (N_3015,N_2609,N_2583);
or U3016 (N_3016,N_2946,N_2499);
or U3017 (N_3017,N_2590,N_2298);
and U3018 (N_3018,N_2781,N_2647);
nand U3019 (N_3019,N_2471,N_2023);
or U3020 (N_3020,N_2972,N_2150);
and U3021 (N_3021,N_2873,N_2489);
nand U3022 (N_3022,N_2816,N_2456);
or U3023 (N_3023,N_2025,N_2115);
and U3024 (N_3024,N_2451,N_2263);
nor U3025 (N_3025,N_2886,N_2088);
or U3026 (N_3026,N_2430,N_2296);
and U3027 (N_3027,N_2967,N_2525);
and U3028 (N_3028,N_2405,N_2825);
xnor U3029 (N_3029,N_2618,N_2965);
and U3030 (N_3030,N_2854,N_2086);
nor U3031 (N_3031,N_2768,N_2137);
nand U3032 (N_3032,N_2547,N_2410);
and U3033 (N_3033,N_2146,N_2264);
nand U3034 (N_3034,N_2976,N_2777);
or U3035 (N_3035,N_2443,N_2311);
nor U3036 (N_3036,N_2013,N_2942);
nand U3037 (N_3037,N_2077,N_2314);
xor U3038 (N_3038,N_2063,N_2017);
xnor U3039 (N_3039,N_2655,N_2984);
or U3040 (N_3040,N_2789,N_2468);
nand U3041 (N_3041,N_2882,N_2543);
or U3042 (N_3042,N_2776,N_2527);
nand U3043 (N_3043,N_2670,N_2148);
or U3044 (N_3044,N_2246,N_2426);
nand U3045 (N_3045,N_2010,N_2810);
nor U3046 (N_3046,N_2557,N_2855);
nor U3047 (N_3047,N_2753,N_2496);
and U3048 (N_3048,N_2613,N_2531);
and U3049 (N_3049,N_2428,N_2308);
and U3050 (N_3050,N_2368,N_2695);
or U3051 (N_3051,N_2289,N_2015);
and U3052 (N_3052,N_2247,N_2605);
nand U3053 (N_3053,N_2804,N_2604);
nor U3054 (N_3054,N_2657,N_2945);
and U3055 (N_3055,N_2936,N_2567);
nand U3056 (N_3056,N_2755,N_2549);
nand U3057 (N_3057,N_2836,N_2584);
and U3058 (N_3058,N_2377,N_2352);
nand U3059 (N_3059,N_2351,N_2986);
or U3060 (N_3060,N_2414,N_2708);
and U3061 (N_3061,N_2217,N_2006);
nand U3062 (N_3062,N_2864,N_2096);
nand U3063 (N_3063,N_2388,N_2259);
nand U3064 (N_3064,N_2491,N_2920);
nor U3065 (N_3065,N_2282,N_2929);
and U3066 (N_3066,N_2078,N_2162);
nor U3067 (N_3067,N_2667,N_2126);
nor U3068 (N_3068,N_2733,N_2042);
and U3069 (N_3069,N_2619,N_2674);
nor U3070 (N_3070,N_2747,N_2062);
or U3071 (N_3071,N_2576,N_2101);
nor U3072 (N_3072,N_2363,N_2258);
and U3073 (N_3073,N_2169,N_2469);
or U3074 (N_3074,N_2828,N_2559);
nor U3075 (N_3075,N_2081,N_2602);
nor U3076 (N_3076,N_2441,N_2280);
and U3077 (N_3077,N_2159,N_2193);
and U3078 (N_3078,N_2370,N_2853);
nor U3079 (N_3079,N_2757,N_2401);
nand U3080 (N_3080,N_2980,N_2450);
nor U3081 (N_3081,N_2249,N_2534);
and U3082 (N_3082,N_2809,N_2540);
nor U3083 (N_3083,N_2808,N_2415);
nor U3084 (N_3084,N_2355,N_2843);
and U3085 (N_3085,N_2234,N_2286);
or U3086 (N_3086,N_2612,N_2925);
nor U3087 (N_3087,N_2216,N_2516);
and U3088 (N_3088,N_2849,N_2347);
nand U3089 (N_3089,N_2519,N_2682);
or U3090 (N_3090,N_2365,N_2959);
or U3091 (N_3091,N_2822,N_2707);
nor U3092 (N_3092,N_2453,N_2274);
nand U3093 (N_3093,N_2526,N_2236);
nand U3094 (N_3094,N_2727,N_2676);
nand U3095 (N_3095,N_2681,N_2575);
and U3096 (N_3096,N_2720,N_2799);
nor U3097 (N_3097,N_2710,N_2551);
or U3098 (N_3098,N_2654,N_2205);
or U3099 (N_3099,N_2743,N_2729);
nor U3100 (N_3100,N_2730,N_2037);
nor U3101 (N_3101,N_2599,N_2341);
and U3102 (N_3102,N_2046,N_2591);
and U3103 (N_3103,N_2458,N_2497);
and U3104 (N_3104,N_2664,N_2908);
nand U3105 (N_3105,N_2631,N_2932);
nand U3106 (N_3106,N_2470,N_2673);
and U3107 (N_3107,N_2878,N_2191);
or U3108 (N_3108,N_2542,N_2898);
nor U3109 (N_3109,N_2283,N_2750);
nand U3110 (N_3110,N_2724,N_2418);
and U3111 (N_3111,N_2248,N_2151);
xnor U3112 (N_3112,N_2866,N_2412);
nand U3113 (N_3113,N_2465,N_2054);
and U3114 (N_3114,N_2649,N_2581);
xor U3115 (N_3115,N_2722,N_2323);
and U3116 (N_3116,N_2887,N_2330);
or U3117 (N_3117,N_2120,N_2691);
or U3118 (N_3118,N_2702,N_2677);
or U3119 (N_3119,N_2005,N_2901);
xnor U3120 (N_3120,N_2011,N_2685);
nand U3121 (N_3121,N_2815,N_2772);
or U3122 (N_3122,N_2760,N_2281);
and U3123 (N_3123,N_2302,N_2686);
and U3124 (N_3124,N_2716,N_2990);
nand U3125 (N_3125,N_2462,N_2635);
nand U3126 (N_3126,N_2869,N_2475);
or U3127 (N_3127,N_2800,N_2284);
nand U3128 (N_3128,N_2883,N_2224);
nor U3129 (N_3129,N_2104,N_2279);
nand U3130 (N_3130,N_2830,N_2239);
and U3131 (N_3131,N_2593,N_2317);
nor U3132 (N_3132,N_2709,N_2937);
or U3133 (N_3133,N_2328,N_2407);
or U3134 (N_3134,N_2472,N_2732);
and U3135 (N_3135,N_2058,N_2877);
nand U3136 (N_3136,N_2174,N_2291);
nand U3137 (N_3137,N_2867,N_2027);
or U3138 (N_3138,N_2968,N_2031);
or U3139 (N_3139,N_2145,N_2287);
nand U3140 (N_3140,N_2072,N_2416);
xnor U3141 (N_3141,N_2127,N_2577);
or U3142 (N_3142,N_2009,N_2087);
nand U3143 (N_3143,N_2518,N_2422);
or U3144 (N_3144,N_2999,N_2406);
and U3145 (N_3145,N_2556,N_2859);
nand U3146 (N_3146,N_2502,N_2973);
nand U3147 (N_3147,N_2767,N_2500);
xor U3148 (N_3148,N_2628,N_2641);
nand U3149 (N_3149,N_2425,N_2554);
nor U3150 (N_3150,N_2638,N_2303);
and U3151 (N_3151,N_2048,N_2243);
and U3152 (N_3152,N_2211,N_2261);
nand U3153 (N_3153,N_2774,N_2988);
nor U3154 (N_3154,N_2269,N_2506);
or U3155 (N_3155,N_2343,N_2218);
nand U3156 (N_3156,N_2910,N_2693);
nor U3157 (N_3157,N_2299,N_2663);
nor U3158 (N_3158,N_2879,N_2884);
nor U3159 (N_3159,N_2260,N_2586);
nand U3160 (N_3160,N_2589,N_2580);
xnor U3161 (N_3161,N_2463,N_2212);
or U3162 (N_3162,N_2252,N_2913);
or U3163 (N_3163,N_2626,N_2158);
nor U3164 (N_3164,N_2226,N_2117);
and U3165 (N_3165,N_2488,N_2440);
nand U3166 (N_3166,N_2833,N_2672);
or U3167 (N_3167,N_2752,N_2424);
or U3168 (N_3168,N_2659,N_2636);
or U3169 (N_3169,N_2036,N_2943);
and U3170 (N_3170,N_2838,N_2241);
nor U3171 (N_3171,N_2178,N_2235);
nand U3172 (N_3172,N_2041,N_2438);
or U3173 (N_3173,N_2204,N_2503);
or U3174 (N_3174,N_2307,N_2487);
nor U3175 (N_3175,N_2220,N_2210);
or U3176 (N_3176,N_2356,N_2982);
and U3177 (N_3177,N_2138,N_2118);
and U3178 (N_3178,N_2257,N_2092);
or U3179 (N_3179,N_2924,N_2601);
nor U3180 (N_3180,N_2400,N_2136);
nand U3181 (N_3181,N_2060,N_2773);
nand U3182 (N_3182,N_2940,N_2206);
nand U3183 (N_3183,N_2070,N_2071);
or U3184 (N_3184,N_2826,N_2595);
or U3185 (N_3185,N_2790,N_2894);
and U3186 (N_3186,N_2219,N_2043);
and U3187 (N_3187,N_2630,N_2265);
or U3188 (N_3188,N_2934,N_2271);
or U3189 (N_3189,N_2566,N_2026);
nor U3190 (N_3190,N_2678,N_2033);
or U3191 (N_3191,N_2012,N_2433);
xor U3192 (N_3192,N_2020,N_2268);
or U3193 (N_3193,N_2508,N_2780);
nand U3194 (N_3194,N_2983,N_2787);
or U3195 (N_3195,N_2285,N_2395);
nand U3196 (N_3196,N_2978,N_2899);
nor U3197 (N_3197,N_2614,N_2479);
nor U3198 (N_3198,N_2277,N_2266);
and U3199 (N_3199,N_2004,N_2478);
or U3200 (N_3200,N_2000,N_2985);
nor U3201 (N_3201,N_2961,N_2511);
and U3202 (N_3202,N_2294,N_2018);
or U3203 (N_3203,N_2200,N_2570);
nand U3204 (N_3204,N_2652,N_2373);
nor U3205 (N_3205,N_2208,N_2524);
nand U3206 (N_3206,N_2522,N_2907);
nor U3207 (N_3207,N_2132,N_2571);
nand U3208 (N_3208,N_2893,N_2436);
or U3209 (N_3209,N_2477,N_2515);
nand U3210 (N_3210,N_2918,N_2858);
and U3211 (N_3211,N_2759,N_2155);
or U3212 (N_3212,N_2326,N_2817);
nand U3213 (N_3213,N_2568,N_2625);
nand U3214 (N_3214,N_2357,N_2761);
and U3215 (N_3215,N_2541,N_2738);
or U3216 (N_3216,N_2332,N_2981);
nor U3217 (N_3217,N_2250,N_2333);
nor U3218 (N_3218,N_2544,N_2318);
nor U3219 (N_3219,N_2313,N_2863);
or U3220 (N_3220,N_2569,N_2089);
and U3221 (N_3221,N_2109,N_2007);
nor U3222 (N_3222,N_2713,N_2545);
or U3223 (N_3223,N_2669,N_2270);
or U3224 (N_3224,N_2254,N_2349);
nand U3225 (N_3225,N_2537,N_2404);
nor U3226 (N_3226,N_2608,N_2044);
nor U3227 (N_3227,N_2172,N_2930);
nand U3228 (N_3228,N_2449,N_2827);
and U3229 (N_3229,N_2692,N_2059);
and U3230 (N_3230,N_2742,N_2834);
nand U3231 (N_3231,N_2675,N_2186);
nor U3232 (N_3232,N_2066,N_2788);
nand U3233 (N_3233,N_2413,N_2085);
nand U3234 (N_3234,N_2835,N_2875);
or U3235 (N_3235,N_2679,N_2080);
and U3236 (N_3236,N_2344,N_2874);
and U3237 (N_3237,N_2550,N_2871);
nor U3238 (N_3238,N_2035,N_2242);
nor U3239 (N_3239,N_2272,N_2001);
nor U3240 (N_3240,N_2480,N_2995);
and U3241 (N_3241,N_2331,N_2510);
nor U3242 (N_3242,N_2606,N_2689);
nor U3243 (N_3243,N_2624,N_2848);
nor U3244 (N_3244,N_2548,N_2369);
or U3245 (N_3245,N_2213,N_2306);
and U3246 (N_3246,N_2949,N_2735);
nor U3247 (N_3247,N_2900,N_2704);
nor U3248 (N_3248,N_2991,N_2596);
nor U3249 (N_3249,N_2233,N_2315);
nand U3250 (N_3250,N_2327,N_2513);
nand U3251 (N_3251,N_2448,N_2814);
nand U3252 (N_3252,N_2103,N_2494);
nand U3253 (N_3253,N_2338,N_2795);
nor U3254 (N_3254,N_2779,N_2643);
nor U3255 (N_3255,N_2350,N_2935);
and U3256 (N_3256,N_2737,N_2161);
nand U3257 (N_3257,N_2094,N_2435);
nand U3258 (N_3258,N_2954,N_2521);
nand U3259 (N_3259,N_2536,N_2564);
nand U3260 (N_3260,N_2758,N_2288);
nor U3261 (N_3261,N_2769,N_2546);
nand U3262 (N_3262,N_2446,N_2486);
and U3263 (N_3263,N_2616,N_2952);
or U3264 (N_3264,N_2135,N_2987);
nand U3265 (N_3265,N_2180,N_2354);
and U3266 (N_3266,N_2914,N_2736);
nand U3267 (N_3267,N_2290,N_2485);
and U3268 (N_3268,N_2749,N_2971);
nand U3269 (N_3269,N_2765,N_2931);
nor U3270 (N_3270,N_2533,N_2267);
nand U3271 (N_3271,N_2429,N_2579);
nor U3272 (N_3272,N_2455,N_2573);
nand U3273 (N_3273,N_2142,N_2361);
xnor U3274 (N_3274,N_2794,N_2922);
nand U3275 (N_3275,N_2228,N_2740);
nor U3276 (N_3276,N_2611,N_2770);
nor U3277 (N_3277,N_2839,N_2454);
nand U3278 (N_3278,N_2700,N_2562);
or U3279 (N_3279,N_2199,N_2711);
or U3280 (N_3280,N_2047,N_2008);
nand U3281 (N_3281,N_2963,N_2585);
or U3282 (N_3282,N_2292,N_2637);
and U3283 (N_3283,N_2627,N_2014);
and U3284 (N_3284,N_2998,N_2394);
or U3285 (N_3285,N_2157,N_2457);
nor U3286 (N_3286,N_2238,N_2346);
nand U3287 (N_3287,N_2181,N_2851);
or U3288 (N_3288,N_2818,N_2530);
nor U3289 (N_3289,N_2336,N_2371);
nor U3290 (N_3290,N_2053,N_2951);
and U3291 (N_3291,N_2055,N_2030);
or U3292 (N_3292,N_2131,N_2671);
or U3293 (N_3293,N_2597,N_2050);
or U3294 (N_3294,N_2362,N_2310);
nor U3295 (N_3295,N_2841,N_2688);
nand U3296 (N_3296,N_2507,N_2928);
nor U3297 (N_3297,N_2068,N_2461);
xnor U3298 (N_3298,N_2844,N_2187);
nand U3299 (N_3299,N_2316,N_2466);
nand U3300 (N_3300,N_2705,N_2119);
or U3301 (N_3301,N_2802,N_2143);
or U3302 (N_3302,N_2558,N_2411);
nor U3303 (N_3303,N_2334,N_2656);
and U3304 (N_3304,N_2147,N_2969);
or U3305 (N_3305,N_2796,N_2870);
or U3306 (N_3306,N_2116,N_2989);
xnor U3307 (N_3307,N_2762,N_2382);
nor U3308 (N_3308,N_2002,N_2417);
nor U3309 (N_3309,N_2182,N_2782);
or U3310 (N_3310,N_2057,N_2402);
nand U3311 (N_3311,N_2032,N_2783);
nor U3312 (N_3312,N_2823,N_2831);
xnor U3313 (N_3313,N_2490,N_2786);
or U3314 (N_3314,N_2237,N_2731);
nand U3315 (N_3315,N_2091,N_2578);
or U3316 (N_3316,N_2634,N_2372);
and U3317 (N_3317,N_2301,N_2065);
nand U3318 (N_3318,N_2207,N_2393);
nor U3319 (N_3319,N_2939,N_2051);
nor U3320 (N_3320,N_2251,N_2917);
xnor U3321 (N_3321,N_2231,N_2906);
or U3322 (N_3322,N_2728,N_2520);
nand U3323 (N_3323,N_2197,N_2964);
xor U3324 (N_3324,N_2803,N_2095);
nand U3325 (N_3325,N_2846,N_2275);
nand U3326 (N_3326,N_2431,N_2861);
and U3327 (N_3327,N_2842,N_2766);
and U3328 (N_3328,N_2793,N_2209);
xnor U3329 (N_3329,N_2916,N_2725);
or U3330 (N_3330,N_2167,N_2084);
nor U3331 (N_3331,N_2962,N_2572);
or U3332 (N_3332,N_2442,N_2482);
and U3333 (N_3333,N_2045,N_2493);
nor U3334 (N_3334,N_2113,N_2278);
or U3335 (N_3335,N_2840,N_2322);
nand U3336 (N_3336,N_2633,N_2295);
nand U3337 (N_3337,N_2797,N_2075);
nand U3338 (N_3338,N_2223,N_2171);
or U3339 (N_3339,N_2603,N_2476);
and U3340 (N_3340,N_2812,N_2152);
nand U3341 (N_3341,N_2367,N_2256);
or U3342 (N_3342,N_2194,N_2215);
nor U3343 (N_3343,N_2819,N_2121);
and U3344 (N_3344,N_2856,N_2105);
nand U3345 (N_3345,N_2865,N_2885);
nor U3346 (N_3346,N_2110,N_2746);
nand U3347 (N_3347,N_2646,N_2911);
nor U3348 (N_3348,N_2644,N_2409);
and U3349 (N_3349,N_2185,N_2598);
and U3350 (N_3350,N_2950,N_2312);
or U3351 (N_3351,N_2993,N_2651);
nand U3352 (N_3352,N_2850,N_2064);
nor U3353 (N_3353,N_2304,N_2067);
nand U3354 (N_3354,N_2229,N_2715);
or U3355 (N_3355,N_2378,N_2505);
and U3356 (N_3356,N_2621,N_2481);
nor U3357 (N_3357,N_2039,N_2666);
and U3358 (N_3358,N_2082,N_2380);
xor U3359 (N_3359,N_2240,N_2300);
or U3360 (N_3360,N_2112,N_2723);
and U3361 (N_3361,N_2535,N_2385);
nor U3362 (N_3362,N_2340,N_2909);
nand U3363 (N_3363,N_2915,N_2574);
and U3364 (N_3364,N_2653,N_2166);
and U3365 (N_3365,N_2560,N_2384);
and U3366 (N_3366,N_2040,N_2123);
and U3367 (N_3367,N_2245,N_2163);
and U3368 (N_3368,N_2358,N_2748);
and U3369 (N_3369,N_2763,N_2726);
or U3370 (N_3370,N_2498,N_2703);
or U3371 (N_3371,N_2845,N_2665);
nand U3372 (N_3372,N_2386,N_2829);
nor U3373 (N_3373,N_2563,N_2321);
nor U3374 (N_3374,N_2360,N_2403);
or U3375 (N_3375,N_2179,N_2617);
nor U3376 (N_3376,N_2375,N_2514);
nor U3377 (N_3377,N_2073,N_2690);
and U3378 (N_3378,N_2512,N_2203);
and U3379 (N_3379,N_2820,N_2111);
or U3380 (N_3380,N_2701,N_2214);
nor U3381 (N_3381,N_2588,N_2320);
nor U3382 (N_3382,N_2144,N_2532);
nor U3383 (N_3383,N_2387,N_2694);
and U3384 (N_3384,N_2891,N_2141);
nand U3385 (N_3385,N_2177,N_2620);
and U3386 (N_3386,N_2941,N_2889);
and U3387 (N_3387,N_2996,N_2160);
and U3388 (N_3388,N_2955,N_2140);
and U3389 (N_3389,N_2896,N_2607);
or U3390 (N_3390,N_2099,N_2460);
or U3391 (N_3391,N_2565,N_2473);
nor U3392 (N_3392,N_2658,N_2183);
xnor U3393 (N_3393,N_2697,N_2337);
nor U3394 (N_3394,N_2447,N_2339);
nor U3395 (N_3395,N_2439,N_2801);
and U3396 (N_3396,N_2421,N_2202);
nand U3397 (N_3397,N_2528,N_2124);
nand U3398 (N_3398,N_2090,N_2379);
nor U3399 (N_3399,N_2022,N_2432);
nor U3400 (N_3400,N_2504,N_2957);
or U3401 (N_3401,N_2668,N_2919);
and U3402 (N_3402,N_2190,N_2003);
and U3403 (N_3403,N_2642,N_2434);
nor U3404 (N_3404,N_2153,N_2134);
and U3405 (N_3405,N_2714,N_2038);
or U3406 (N_3406,N_2225,N_2221);
xor U3407 (N_3407,N_2698,N_2100);
nand U3408 (N_3408,N_2198,N_2696);
nand U3409 (N_3409,N_2125,N_2744);
or U3410 (N_3410,N_2538,N_2353);
nor U3411 (N_3411,N_2276,N_2852);
nand U3412 (N_3412,N_2881,N_2128);
nand U3413 (N_3413,N_2175,N_2149);
xnor U3414 (N_3414,N_2297,N_2227);
and U3415 (N_3415,N_2805,N_2398);
or U3416 (N_3416,N_2106,N_2684);
nor U3417 (N_3417,N_2645,N_2745);
or U3418 (N_3418,N_2821,N_2399);
or U3419 (N_3419,N_2364,N_2122);
nand U3420 (N_3420,N_2824,N_2872);
or U3421 (N_3421,N_2994,N_2639);
or U3422 (N_3422,N_2632,N_2097);
nand U3423 (N_3423,N_2927,N_2857);
nand U3424 (N_3424,N_2699,N_2107);
nand U3425 (N_3425,N_2419,N_2056);
nand U3426 (N_3426,N_2444,N_2622);
nor U3427 (N_3427,N_2130,N_2230);
nor U3428 (N_3428,N_2324,N_2255);
or U3429 (N_3429,N_2552,N_2467);
nor U3430 (N_3430,N_2102,N_2837);
and U3431 (N_3431,N_2662,N_2374);
xor U3432 (N_3432,N_2173,N_2028);
or U3433 (N_3433,N_2376,N_2342);
or U3434 (N_3434,N_2902,N_2648);
and U3435 (N_3435,N_2778,N_2164);
nand U3436 (N_3436,N_2517,N_2661);
or U3437 (N_3437,N_2495,N_2719);
and U3438 (N_3438,N_2660,N_2201);
and U3439 (N_3439,N_2629,N_2390);
nor U3440 (N_3440,N_2977,N_2391);
or U3441 (N_3441,N_2926,N_2445);
nor U3442 (N_3442,N_2396,N_2610);
nand U3443 (N_3443,N_2974,N_2483);
nor U3444 (N_3444,N_2960,N_2683);
nor U3445 (N_3445,N_2170,N_2975);
or U3446 (N_3446,N_2222,N_2492);
or U3447 (N_3447,N_2811,N_2024);
or U3448 (N_3448,N_2325,N_2751);
nand U3449 (N_3449,N_2687,N_2832);
and U3450 (N_3450,N_2903,N_2888);
and U3451 (N_3451,N_2273,N_2897);
or U3452 (N_3452,N_2615,N_2154);
and U3453 (N_3453,N_2262,N_2555);
nor U3454 (N_3454,N_2553,N_2156);
and U3455 (N_3455,N_2792,N_2452);
nand U3456 (N_3456,N_2966,N_2034);
nand U3457 (N_3457,N_2717,N_2195);
or U3458 (N_3458,N_2129,N_2862);
and U3459 (N_3459,N_2712,N_2944);
or U3460 (N_3460,N_2484,N_2345);
nand U3461 (N_3461,N_2189,N_2397);
or U3462 (N_3462,N_2079,N_2093);
nand U3463 (N_3463,N_2423,N_2892);
or U3464 (N_3464,N_2947,N_2905);
or U3465 (N_3465,N_2948,N_2895);
or U3466 (N_3466,N_2464,N_2938);
nand U3467 (N_3467,N_2293,N_2868);
and U3468 (N_3468,N_2775,N_2420);
nand U3469 (N_3469,N_2582,N_2168);
or U3470 (N_3470,N_2640,N_2592);
or U3471 (N_3471,N_2392,N_2427);
nor U3472 (N_3472,N_2958,N_2359);
and U3473 (N_3473,N_2329,N_2718);
and U3474 (N_3474,N_2196,N_2921);
nand U3475 (N_3475,N_2997,N_2052);
nor U3476 (N_3476,N_2348,N_2133);
nand U3477 (N_3477,N_2561,N_2188);
nand U3478 (N_3478,N_2912,N_2389);
nor U3479 (N_3479,N_2108,N_2319);
nor U3480 (N_3480,N_2192,N_2734);
nand U3481 (N_3481,N_2721,N_2309);
and U3482 (N_3482,N_2594,N_2890);
nor U3483 (N_3483,N_2381,N_2501);
nand U3484 (N_3484,N_2784,N_2165);
nand U3485 (N_3485,N_2244,N_2083);
and U3486 (N_3486,N_2459,N_2016);
nand U3487 (N_3487,N_2184,N_2623);
and U3488 (N_3488,N_2029,N_2860);
or U3489 (N_3489,N_2970,N_2933);
and U3490 (N_3490,N_2754,N_2176);
nor U3491 (N_3491,N_2741,N_2076);
or U3492 (N_3492,N_2956,N_2587);
nand U3493 (N_3493,N_2139,N_2650);
and U3494 (N_3494,N_2098,N_2680);
or U3495 (N_3495,N_2049,N_2408);
nor U3496 (N_3496,N_2114,N_2474);
nor U3497 (N_3497,N_2600,N_2253);
or U3498 (N_3498,N_2756,N_2232);
and U3499 (N_3499,N_2539,N_2953);
and U3500 (N_3500,N_2003,N_2913);
nor U3501 (N_3501,N_2159,N_2836);
and U3502 (N_3502,N_2709,N_2804);
and U3503 (N_3503,N_2319,N_2846);
nor U3504 (N_3504,N_2869,N_2874);
and U3505 (N_3505,N_2734,N_2003);
xor U3506 (N_3506,N_2520,N_2187);
or U3507 (N_3507,N_2106,N_2395);
and U3508 (N_3508,N_2278,N_2801);
nand U3509 (N_3509,N_2818,N_2205);
and U3510 (N_3510,N_2897,N_2113);
and U3511 (N_3511,N_2095,N_2840);
or U3512 (N_3512,N_2489,N_2663);
nand U3513 (N_3513,N_2399,N_2383);
nand U3514 (N_3514,N_2731,N_2181);
nor U3515 (N_3515,N_2673,N_2289);
nor U3516 (N_3516,N_2548,N_2672);
and U3517 (N_3517,N_2171,N_2846);
nor U3518 (N_3518,N_2318,N_2158);
nor U3519 (N_3519,N_2748,N_2832);
or U3520 (N_3520,N_2831,N_2446);
and U3521 (N_3521,N_2638,N_2958);
or U3522 (N_3522,N_2406,N_2289);
xor U3523 (N_3523,N_2534,N_2880);
nand U3524 (N_3524,N_2144,N_2202);
nand U3525 (N_3525,N_2450,N_2202);
nor U3526 (N_3526,N_2048,N_2426);
or U3527 (N_3527,N_2601,N_2358);
and U3528 (N_3528,N_2253,N_2554);
nor U3529 (N_3529,N_2853,N_2909);
and U3530 (N_3530,N_2503,N_2117);
and U3531 (N_3531,N_2621,N_2349);
and U3532 (N_3532,N_2425,N_2732);
nand U3533 (N_3533,N_2479,N_2795);
nand U3534 (N_3534,N_2930,N_2711);
or U3535 (N_3535,N_2803,N_2456);
and U3536 (N_3536,N_2326,N_2007);
and U3537 (N_3537,N_2413,N_2804);
and U3538 (N_3538,N_2683,N_2665);
and U3539 (N_3539,N_2505,N_2434);
and U3540 (N_3540,N_2265,N_2611);
and U3541 (N_3541,N_2112,N_2015);
and U3542 (N_3542,N_2013,N_2821);
nand U3543 (N_3543,N_2174,N_2643);
nor U3544 (N_3544,N_2704,N_2581);
xor U3545 (N_3545,N_2560,N_2568);
or U3546 (N_3546,N_2709,N_2998);
or U3547 (N_3547,N_2656,N_2370);
or U3548 (N_3548,N_2063,N_2220);
or U3549 (N_3549,N_2698,N_2965);
or U3550 (N_3550,N_2082,N_2907);
nor U3551 (N_3551,N_2518,N_2111);
nand U3552 (N_3552,N_2480,N_2062);
nor U3553 (N_3553,N_2539,N_2287);
nor U3554 (N_3554,N_2621,N_2119);
nand U3555 (N_3555,N_2008,N_2568);
nor U3556 (N_3556,N_2509,N_2201);
nor U3557 (N_3557,N_2437,N_2526);
or U3558 (N_3558,N_2316,N_2641);
nand U3559 (N_3559,N_2196,N_2543);
nor U3560 (N_3560,N_2472,N_2320);
or U3561 (N_3561,N_2773,N_2754);
or U3562 (N_3562,N_2666,N_2122);
and U3563 (N_3563,N_2279,N_2249);
and U3564 (N_3564,N_2010,N_2359);
or U3565 (N_3565,N_2020,N_2926);
or U3566 (N_3566,N_2732,N_2093);
or U3567 (N_3567,N_2093,N_2358);
nor U3568 (N_3568,N_2085,N_2394);
nand U3569 (N_3569,N_2452,N_2545);
nor U3570 (N_3570,N_2402,N_2483);
nand U3571 (N_3571,N_2227,N_2774);
or U3572 (N_3572,N_2227,N_2546);
or U3573 (N_3573,N_2722,N_2322);
xor U3574 (N_3574,N_2270,N_2407);
or U3575 (N_3575,N_2920,N_2108);
nand U3576 (N_3576,N_2666,N_2815);
or U3577 (N_3577,N_2224,N_2931);
nand U3578 (N_3578,N_2228,N_2611);
nand U3579 (N_3579,N_2747,N_2320);
or U3580 (N_3580,N_2843,N_2667);
nand U3581 (N_3581,N_2567,N_2991);
nor U3582 (N_3582,N_2666,N_2695);
nor U3583 (N_3583,N_2247,N_2914);
nor U3584 (N_3584,N_2077,N_2896);
nor U3585 (N_3585,N_2541,N_2780);
and U3586 (N_3586,N_2829,N_2106);
and U3587 (N_3587,N_2520,N_2826);
nand U3588 (N_3588,N_2362,N_2791);
nor U3589 (N_3589,N_2353,N_2475);
xor U3590 (N_3590,N_2926,N_2496);
nand U3591 (N_3591,N_2009,N_2183);
nand U3592 (N_3592,N_2374,N_2656);
or U3593 (N_3593,N_2137,N_2916);
nor U3594 (N_3594,N_2822,N_2884);
nor U3595 (N_3595,N_2731,N_2932);
and U3596 (N_3596,N_2727,N_2502);
nand U3597 (N_3597,N_2685,N_2909);
and U3598 (N_3598,N_2270,N_2662);
or U3599 (N_3599,N_2659,N_2645);
nor U3600 (N_3600,N_2506,N_2652);
or U3601 (N_3601,N_2070,N_2505);
nand U3602 (N_3602,N_2735,N_2397);
nor U3603 (N_3603,N_2583,N_2266);
and U3604 (N_3604,N_2518,N_2978);
nand U3605 (N_3605,N_2028,N_2265);
nor U3606 (N_3606,N_2405,N_2070);
and U3607 (N_3607,N_2791,N_2771);
xnor U3608 (N_3608,N_2042,N_2582);
and U3609 (N_3609,N_2835,N_2589);
nor U3610 (N_3610,N_2103,N_2751);
nor U3611 (N_3611,N_2617,N_2615);
nor U3612 (N_3612,N_2984,N_2029);
or U3613 (N_3613,N_2957,N_2686);
and U3614 (N_3614,N_2075,N_2769);
and U3615 (N_3615,N_2365,N_2195);
nor U3616 (N_3616,N_2466,N_2111);
nand U3617 (N_3617,N_2177,N_2687);
nand U3618 (N_3618,N_2706,N_2212);
nor U3619 (N_3619,N_2445,N_2332);
or U3620 (N_3620,N_2517,N_2062);
nand U3621 (N_3621,N_2352,N_2170);
nor U3622 (N_3622,N_2651,N_2900);
and U3623 (N_3623,N_2553,N_2308);
or U3624 (N_3624,N_2380,N_2761);
or U3625 (N_3625,N_2626,N_2043);
and U3626 (N_3626,N_2028,N_2494);
and U3627 (N_3627,N_2463,N_2116);
or U3628 (N_3628,N_2998,N_2205);
nor U3629 (N_3629,N_2114,N_2745);
or U3630 (N_3630,N_2777,N_2107);
and U3631 (N_3631,N_2166,N_2156);
and U3632 (N_3632,N_2480,N_2735);
or U3633 (N_3633,N_2416,N_2180);
nand U3634 (N_3634,N_2554,N_2732);
nor U3635 (N_3635,N_2873,N_2006);
nand U3636 (N_3636,N_2151,N_2704);
and U3637 (N_3637,N_2208,N_2935);
and U3638 (N_3638,N_2008,N_2217);
and U3639 (N_3639,N_2974,N_2485);
nand U3640 (N_3640,N_2350,N_2578);
nand U3641 (N_3641,N_2250,N_2493);
nand U3642 (N_3642,N_2919,N_2621);
nor U3643 (N_3643,N_2834,N_2149);
and U3644 (N_3644,N_2709,N_2470);
or U3645 (N_3645,N_2667,N_2106);
and U3646 (N_3646,N_2734,N_2903);
and U3647 (N_3647,N_2725,N_2450);
nor U3648 (N_3648,N_2658,N_2152);
nand U3649 (N_3649,N_2246,N_2415);
or U3650 (N_3650,N_2931,N_2646);
nor U3651 (N_3651,N_2094,N_2184);
and U3652 (N_3652,N_2921,N_2659);
or U3653 (N_3653,N_2070,N_2689);
and U3654 (N_3654,N_2737,N_2321);
nor U3655 (N_3655,N_2627,N_2940);
nand U3656 (N_3656,N_2414,N_2031);
and U3657 (N_3657,N_2453,N_2367);
and U3658 (N_3658,N_2053,N_2405);
nand U3659 (N_3659,N_2518,N_2532);
nand U3660 (N_3660,N_2318,N_2682);
or U3661 (N_3661,N_2962,N_2496);
nand U3662 (N_3662,N_2364,N_2225);
nor U3663 (N_3663,N_2877,N_2593);
nor U3664 (N_3664,N_2868,N_2006);
nand U3665 (N_3665,N_2533,N_2956);
nor U3666 (N_3666,N_2799,N_2401);
nand U3667 (N_3667,N_2507,N_2247);
nand U3668 (N_3668,N_2083,N_2265);
and U3669 (N_3669,N_2950,N_2527);
nand U3670 (N_3670,N_2841,N_2580);
nor U3671 (N_3671,N_2546,N_2526);
nand U3672 (N_3672,N_2443,N_2133);
and U3673 (N_3673,N_2802,N_2264);
nor U3674 (N_3674,N_2127,N_2156);
or U3675 (N_3675,N_2509,N_2967);
or U3676 (N_3676,N_2244,N_2901);
nand U3677 (N_3677,N_2049,N_2882);
and U3678 (N_3678,N_2481,N_2696);
nand U3679 (N_3679,N_2558,N_2580);
nor U3680 (N_3680,N_2434,N_2194);
nand U3681 (N_3681,N_2275,N_2427);
and U3682 (N_3682,N_2678,N_2902);
nor U3683 (N_3683,N_2712,N_2848);
nor U3684 (N_3684,N_2243,N_2189);
nand U3685 (N_3685,N_2726,N_2676);
or U3686 (N_3686,N_2507,N_2543);
nand U3687 (N_3687,N_2952,N_2180);
or U3688 (N_3688,N_2210,N_2665);
and U3689 (N_3689,N_2582,N_2052);
or U3690 (N_3690,N_2738,N_2753);
or U3691 (N_3691,N_2744,N_2668);
nor U3692 (N_3692,N_2166,N_2925);
nor U3693 (N_3693,N_2172,N_2837);
or U3694 (N_3694,N_2250,N_2147);
or U3695 (N_3695,N_2576,N_2116);
nand U3696 (N_3696,N_2998,N_2244);
nor U3697 (N_3697,N_2487,N_2235);
nand U3698 (N_3698,N_2590,N_2693);
nor U3699 (N_3699,N_2147,N_2646);
or U3700 (N_3700,N_2639,N_2356);
nor U3701 (N_3701,N_2893,N_2265);
nor U3702 (N_3702,N_2980,N_2923);
nand U3703 (N_3703,N_2960,N_2283);
nand U3704 (N_3704,N_2166,N_2124);
and U3705 (N_3705,N_2858,N_2681);
nand U3706 (N_3706,N_2450,N_2459);
and U3707 (N_3707,N_2014,N_2117);
nand U3708 (N_3708,N_2205,N_2200);
nand U3709 (N_3709,N_2865,N_2550);
nor U3710 (N_3710,N_2229,N_2786);
and U3711 (N_3711,N_2078,N_2229);
nand U3712 (N_3712,N_2990,N_2311);
and U3713 (N_3713,N_2067,N_2301);
and U3714 (N_3714,N_2163,N_2561);
and U3715 (N_3715,N_2924,N_2586);
xnor U3716 (N_3716,N_2024,N_2860);
nor U3717 (N_3717,N_2571,N_2669);
nand U3718 (N_3718,N_2566,N_2803);
nand U3719 (N_3719,N_2797,N_2825);
and U3720 (N_3720,N_2555,N_2335);
nor U3721 (N_3721,N_2286,N_2179);
nor U3722 (N_3722,N_2024,N_2632);
nand U3723 (N_3723,N_2439,N_2238);
and U3724 (N_3724,N_2038,N_2854);
and U3725 (N_3725,N_2011,N_2137);
or U3726 (N_3726,N_2996,N_2409);
or U3727 (N_3727,N_2397,N_2469);
nand U3728 (N_3728,N_2202,N_2998);
nand U3729 (N_3729,N_2544,N_2977);
and U3730 (N_3730,N_2419,N_2152);
nor U3731 (N_3731,N_2424,N_2520);
or U3732 (N_3732,N_2359,N_2341);
or U3733 (N_3733,N_2516,N_2012);
or U3734 (N_3734,N_2712,N_2531);
nand U3735 (N_3735,N_2768,N_2125);
nor U3736 (N_3736,N_2553,N_2938);
and U3737 (N_3737,N_2369,N_2897);
nor U3738 (N_3738,N_2590,N_2724);
nand U3739 (N_3739,N_2060,N_2599);
nand U3740 (N_3740,N_2416,N_2418);
and U3741 (N_3741,N_2758,N_2732);
nand U3742 (N_3742,N_2110,N_2671);
nor U3743 (N_3743,N_2918,N_2428);
nand U3744 (N_3744,N_2666,N_2583);
or U3745 (N_3745,N_2672,N_2742);
or U3746 (N_3746,N_2607,N_2352);
and U3747 (N_3747,N_2909,N_2308);
nor U3748 (N_3748,N_2943,N_2322);
nand U3749 (N_3749,N_2356,N_2440);
and U3750 (N_3750,N_2026,N_2445);
and U3751 (N_3751,N_2961,N_2036);
or U3752 (N_3752,N_2324,N_2386);
or U3753 (N_3753,N_2181,N_2745);
nor U3754 (N_3754,N_2415,N_2576);
or U3755 (N_3755,N_2209,N_2840);
or U3756 (N_3756,N_2798,N_2606);
nand U3757 (N_3757,N_2909,N_2302);
and U3758 (N_3758,N_2730,N_2489);
nand U3759 (N_3759,N_2752,N_2345);
nand U3760 (N_3760,N_2520,N_2253);
nor U3761 (N_3761,N_2158,N_2836);
nor U3762 (N_3762,N_2727,N_2369);
nand U3763 (N_3763,N_2208,N_2335);
or U3764 (N_3764,N_2245,N_2526);
and U3765 (N_3765,N_2546,N_2371);
nand U3766 (N_3766,N_2906,N_2169);
nor U3767 (N_3767,N_2659,N_2330);
nor U3768 (N_3768,N_2162,N_2051);
nand U3769 (N_3769,N_2801,N_2732);
nor U3770 (N_3770,N_2011,N_2537);
or U3771 (N_3771,N_2150,N_2447);
and U3772 (N_3772,N_2684,N_2876);
nand U3773 (N_3773,N_2574,N_2220);
or U3774 (N_3774,N_2222,N_2309);
or U3775 (N_3775,N_2201,N_2505);
nand U3776 (N_3776,N_2693,N_2638);
and U3777 (N_3777,N_2143,N_2150);
or U3778 (N_3778,N_2608,N_2353);
nand U3779 (N_3779,N_2047,N_2244);
nand U3780 (N_3780,N_2981,N_2428);
nand U3781 (N_3781,N_2724,N_2788);
or U3782 (N_3782,N_2578,N_2551);
and U3783 (N_3783,N_2303,N_2309);
and U3784 (N_3784,N_2429,N_2774);
or U3785 (N_3785,N_2764,N_2206);
or U3786 (N_3786,N_2185,N_2002);
nor U3787 (N_3787,N_2064,N_2876);
nand U3788 (N_3788,N_2502,N_2121);
nand U3789 (N_3789,N_2242,N_2284);
and U3790 (N_3790,N_2053,N_2872);
or U3791 (N_3791,N_2822,N_2984);
and U3792 (N_3792,N_2909,N_2737);
or U3793 (N_3793,N_2127,N_2616);
and U3794 (N_3794,N_2897,N_2323);
nand U3795 (N_3795,N_2607,N_2242);
and U3796 (N_3796,N_2218,N_2719);
nor U3797 (N_3797,N_2134,N_2701);
and U3798 (N_3798,N_2302,N_2369);
nor U3799 (N_3799,N_2482,N_2588);
nor U3800 (N_3800,N_2510,N_2266);
and U3801 (N_3801,N_2380,N_2008);
and U3802 (N_3802,N_2951,N_2910);
nor U3803 (N_3803,N_2865,N_2559);
and U3804 (N_3804,N_2704,N_2867);
or U3805 (N_3805,N_2285,N_2996);
nand U3806 (N_3806,N_2376,N_2908);
and U3807 (N_3807,N_2106,N_2170);
and U3808 (N_3808,N_2017,N_2970);
nand U3809 (N_3809,N_2454,N_2072);
nor U3810 (N_3810,N_2493,N_2520);
or U3811 (N_3811,N_2955,N_2968);
xnor U3812 (N_3812,N_2393,N_2347);
nor U3813 (N_3813,N_2763,N_2246);
nand U3814 (N_3814,N_2317,N_2967);
and U3815 (N_3815,N_2438,N_2673);
nand U3816 (N_3816,N_2559,N_2799);
nor U3817 (N_3817,N_2966,N_2491);
and U3818 (N_3818,N_2932,N_2995);
nor U3819 (N_3819,N_2946,N_2428);
nand U3820 (N_3820,N_2622,N_2534);
and U3821 (N_3821,N_2067,N_2906);
or U3822 (N_3822,N_2836,N_2563);
or U3823 (N_3823,N_2980,N_2394);
and U3824 (N_3824,N_2979,N_2361);
or U3825 (N_3825,N_2409,N_2238);
nor U3826 (N_3826,N_2388,N_2164);
or U3827 (N_3827,N_2913,N_2350);
or U3828 (N_3828,N_2180,N_2426);
or U3829 (N_3829,N_2915,N_2730);
nand U3830 (N_3830,N_2791,N_2163);
and U3831 (N_3831,N_2602,N_2711);
nor U3832 (N_3832,N_2975,N_2251);
or U3833 (N_3833,N_2394,N_2808);
nor U3834 (N_3834,N_2139,N_2007);
and U3835 (N_3835,N_2046,N_2656);
nand U3836 (N_3836,N_2759,N_2523);
and U3837 (N_3837,N_2166,N_2741);
xor U3838 (N_3838,N_2754,N_2524);
nor U3839 (N_3839,N_2222,N_2818);
nor U3840 (N_3840,N_2569,N_2977);
nand U3841 (N_3841,N_2655,N_2916);
xnor U3842 (N_3842,N_2430,N_2501);
nor U3843 (N_3843,N_2922,N_2130);
nand U3844 (N_3844,N_2427,N_2438);
nor U3845 (N_3845,N_2722,N_2706);
xnor U3846 (N_3846,N_2819,N_2205);
nand U3847 (N_3847,N_2892,N_2810);
nor U3848 (N_3848,N_2052,N_2148);
xor U3849 (N_3849,N_2456,N_2328);
nor U3850 (N_3850,N_2387,N_2438);
nor U3851 (N_3851,N_2865,N_2848);
xor U3852 (N_3852,N_2359,N_2526);
and U3853 (N_3853,N_2537,N_2840);
nor U3854 (N_3854,N_2383,N_2465);
nand U3855 (N_3855,N_2685,N_2108);
or U3856 (N_3856,N_2137,N_2109);
or U3857 (N_3857,N_2178,N_2663);
nand U3858 (N_3858,N_2634,N_2051);
nor U3859 (N_3859,N_2437,N_2300);
nand U3860 (N_3860,N_2086,N_2757);
nor U3861 (N_3861,N_2779,N_2950);
nand U3862 (N_3862,N_2528,N_2389);
and U3863 (N_3863,N_2951,N_2362);
nor U3864 (N_3864,N_2348,N_2326);
nand U3865 (N_3865,N_2578,N_2120);
xor U3866 (N_3866,N_2744,N_2216);
and U3867 (N_3867,N_2444,N_2976);
nand U3868 (N_3868,N_2362,N_2706);
and U3869 (N_3869,N_2117,N_2639);
or U3870 (N_3870,N_2732,N_2978);
or U3871 (N_3871,N_2928,N_2913);
and U3872 (N_3872,N_2382,N_2604);
nand U3873 (N_3873,N_2976,N_2133);
nor U3874 (N_3874,N_2056,N_2589);
xnor U3875 (N_3875,N_2094,N_2390);
or U3876 (N_3876,N_2482,N_2028);
nand U3877 (N_3877,N_2458,N_2369);
and U3878 (N_3878,N_2145,N_2295);
or U3879 (N_3879,N_2936,N_2222);
nand U3880 (N_3880,N_2599,N_2769);
nand U3881 (N_3881,N_2976,N_2366);
or U3882 (N_3882,N_2842,N_2931);
nand U3883 (N_3883,N_2038,N_2392);
xnor U3884 (N_3884,N_2138,N_2742);
and U3885 (N_3885,N_2296,N_2796);
xnor U3886 (N_3886,N_2890,N_2661);
and U3887 (N_3887,N_2873,N_2718);
nor U3888 (N_3888,N_2903,N_2257);
nand U3889 (N_3889,N_2158,N_2153);
nor U3890 (N_3890,N_2245,N_2921);
nand U3891 (N_3891,N_2834,N_2617);
and U3892 (N_3892,N_2670,N_2872);
nor U3893 (N_3893,N_2513,N_2010);
nor U3894 (N_3894,N_2321,N_2088);
nor U3895 (N_3895,N_2067,N_2810);
or U3896 (N_3896,N_2403,N_2262);
and U3897 (N_3897,N_2435,N_2305);
nor U3898 (N_3898,N_2348,N_2995);
or U3899 (N_3899,N_2658,N_2656);
and U3900 (N_3900,N_2853,N_2292);
nor U3901 (N_3901,N_2471,N_2087);
and U3902 (N_3902,N_2948,N_2040);
and U3903 (N_3903,N_2626,N_2907);
nand U3904 (N_3904,N_2146,N_2018);
and U3905 (N_3905,N_2842,N_2162);
nand U3906 (N_3906,N_2303,N_2137);
or U3907 (N_3907,N_2162,N_2342);
nor U3908 (N_3908,N_2173,N_2258);
or U3909 (N_3909,N_2624,N_2143);
and U3910 (N_3910,N_2201,N_2074);
xor U3911 (N_3911,N_2090,N_2992);
and U3912 (N_3912,N_2951,N_2493);
nor U3913 (N_3913,N_2284,N_2596);
or U3914 (N_3914,N_2057,N_2887);
and U3915 (N_3915,N_2583,N_2015);
nor U3916 (N_3916,N_2024,N_2981);
and U3917 (N_3917,N_2843,N_2862);
nand U3918 (N_3918,N_2798,N_2207);
nand U3919 (N_3919,N_2374,N_2626);
nand U3920 (N_3920,N_2747,N_2021);
and U3921 (N_3921,N_2993,N_2680);
nor U3922 (N_3922,N_2866,N_2719);
and U3923 (N_3923,N_2183,N_2435);
nand U3924 (N_3924,N_2635,N_2393);
nor U3925 (N_3925,N_2108,N_2752);
and U3926 (N_3926,N_2605,N_2578);
nor U3927 (N_3927,N_2116,N_2892);
nor U3928 (N_3928,N_2862,N_2653);
or U3929 (N_3929,N_2026,N_2990);
or U3930 (N_3930,N_2061,N_2822);
nand U3931 (N_3931,N_2400,N_2673);
nor U3932 (N_3932,N_2013,N_2440);
or U3933 (N_3933,N_2953,N_2796);
nor U3934 (N_3934,N_2953,N_2053);
nor U3935 (N_3935,N_2415,N_2525);
or U3936 (N_3936,N_2301,N_2263);
nand U3937 (N_3937,N_2471,N_2252);
nand U3938 (N_3938,N_2365,N_2995);
or U3939 (N_3939,N_2839,N_2104);
or U3940 (N_3940,N_2845,N_2336);
and U3941 (N_3941,N_2202,N_2453);
nor U3942 (N_3942,N_2772,N_2082);
or U3943 (N_3943,N_2731,N_2727);
nand U3944 (N_3944,N_2921,N_2376);
nor U3945 (N_3945,N_2823,N_2695);
and U3946 (N_3946,N_2077,N_2059);
nor U3947 (N_3947,N_2881,N_2811);
nor U3948 (N_3948,N_2386,N_2735);
nand U3949 (N_3949,N_2698,N_2109);
or U3950 (N_3950,N_2911,N_2323);
or U3951 (N_3951,N_2148,N_2783);
and U3952 (N_3952,N_2377,N_2394);
and U3953 (N_3953,N_2883,N_2750);
nand U3954 (N_3954,N_2567,N_2215);
or U3955 (N_3955,N_2700,N_2679);
nand U3956 (N_3956,N_2681,N_2544);
nor U3957 (N_3957,N_2550,N_2630);
and U3958 (N_3958,N_2003,N_2654);
nand U3959 (N_3959,N_2618,N_2787);
and U3960 (N_3960,N_2093,N_2466);
nand U3961 (N_3961,N_2176,N_2945);
nor U3962 (N_3962,N_2590,N_2061);
or U3963 (N_3963,N_2236,N_2245);
or U3964 (N_3964,N_2698,N_2763);
nor U3965 (N_3965,N_2467,N_2838);
and U3966 (N_3966,N_2191,N_2872);
or U3967 (N_3967,N_2945,N_2044);
or U3968 (N_3968,N_2309,N_2324);
or U3969 (N_3969,N_2771,N_2758);
and U3970 (N_3970,N_2877,N_2808);
and U3971 (N_3971,N_2792,N_2020);
or U3972 (N_3972,N_2289,N_2567);
nand U3973 (N_3973,N_2539,N_2442);
nand U3974 (N_3974,N_2441,N_2381);
nand U3975 (N_3975,N_2026,N_2838);
or U3976 (N_3976,N_2190,N_2136);
or U3977 (N_3977,N_2954,N_2378);
and U3978 (N_3978,N_2209,N_2077);
xnor U3979 (N_3979,N_2136,N_2277);
nand U3980 (N_3980,N_2817,N_2641);
and U3981 (N_3981,N_2042,N_2298);
or U3982 (N_3982,N_2614,N_2394);
and U3983 (N_3983,N_2285,N_2693);
or U3984 (N_3984,N_2027,N_2739);
or U3985 (N_3985,N_2733,N_2054);
nor U3986 (N_3986,N_2384,N_2421);
nor U3987 (N_3987,N_2998,N_2130);
nand U3988 (N_3988,N_2140,N_2980);
nand U3989 (N_3989,N_2515,N_2465);
and U3990 (N_3990,N_2559,N_2341);
nand U3991 (N_3991,N_2818,N_2920);
nand U3992 (N_3992,N_2754,N_2864);
nor U3993 (N_3993,N_2389,N_2873);
nand U3994 (N_3994,N_2494,N_2409);
nand U3995 (N_3995,N_2816,N_2183);
or U3996 (N_3996,N_2328,N_2973);
nor U3997 (N_3997,N_2333,N_2519);
or U3998 (N_3998,N_2938,N_2954);
nand U3999 (N_3999,N_2109,N_2841);
or U4000 (N_4000,N_3639,N_3960);
or U4001 (N_4001,N_3452,N_3297);
nand U4002 (N_4002,N_3380,N_3594);
nor U4003 (N_4003,N_3079,N_3977);
nand U4004 (N_4004,N_3888,N_3061);
nor U4005 (N_4005,N_3617,N_3915);
xor U4006 (N_4006,N_3476,N_3273);
nand U4007 (N_4007,N_3326,N_3455);
nand U4008 (N_4008,N_3771,N_3746);
nor U4009 (N_4009,N_3116,N_3574);
or U4010 (N_4010,N_3294,N_3472);
and U4011 (N_4011,N_3602,N_3481);
nand U4012 (N_4012,N_3364,N_3780);
nand U4013 (N_4013,N_3862,N_3194);
nor U4014 (N_4014,N_3291,N_3348);
and U4015 (N_4015,N_3508,N_3825);
nor U4016 (N_4016,N_3582,N_3456);
nand U4017 (N_4017,N_3665,N_3424);
or U4018 (N_4018,N_3994,N_3562);
nand U4019 (N_4019,N_3886,N_3894);
or U4020 (N_4020,N_3739,N_3725);
and U4021 (N_4021,N_3680,N_3317);
and U4022 (N_4022,N_3564,N_3839);
nand U4023 (N_4023,N_3415,N_3794);
nor U4024 (N_4024,N_3538,N_3512);
and U4025 (N_4025,N_3936,N_3851);
and U4026 (N_4026,N_3158,N_3596);
nor U4027 (N_4027,N_3514,N_3343);
nor U4028 (N_4028,N_3276,N_3443);
xor U4029 (N_4029,N_3671,N_3316);
xnor U4030 (N_4030,N_3949,N_3482);
nand U4031 (N_4031,N_3840,N_3879);
and U4032 (N_4032,N_3592,N_3823);
or U4033 (N_4033,N_3332,N_3664);
and U4034 (N_4034,N_3855,N_3820);
or U4035 (N_4035,N_3392,N_3454);
nand U4036 (N_4036,N_3585,N_3609);
nand U4037 (N_4037,N_3278,N_3515);
or U4038 (N_4038,N_3333,N_3480);
and U4039 (N_4039,N_3486,N_3106);
and U4040 (N_4040,N_3148,N_3487);
or U4041 (N_4041,N_3162,N_3988);
nor U4042 (N_4042,N_3433,N_3868);
and U4043 (N_4043,N_3793,N_3070);
nor U4044 (N_4044,N_3255,N_3293);
and U4045 (N_4045,N_3553,N_3361);
nand U4046 (N_4046,N_3812,N_3999);
or U4047 (N_4047,N_3922,N_3969);
or U4048 (N_4048,N_3686,N_3701);
nor U4049 (N_4049,N_3288,N_3075);
or U4050 (N_4050,N_3329,N_3144);
and U4051 (N_4051,N_3654,N_3952);
or U4052 (N_4052,N_3381,N_3765);
nor U4053 (N_4053,N_3890,N_3055);
nand U4054 (N_4054,N_3410,N_3253);
nand U4055 (N_4055,N_3753,N_3631);
or U4056 (N_4056,N_3178,N_3159);
or U4057 (N_4057,N_3434,N_3774);
nor U4058 (N_4058,N_3307,N_3470);
xnor U4059 (N_4059,N_3184,N_3981);
nor U4060 (N_4060,N_3087,N_3146);
or U4061 (N_4061,N_3575,N_3499);
and U4062 (N_4062,N_3968,N_3941);
xor U4063 (N_4063,N_3391,N_3783);
nand U4064 (N_4064,N_3718,N_3013);
nor U4065 (N_4065,N_3372,N_3349);
nand U4066 (N_4066,N_3599,N_3036);
nor U4067 (N_4067,N_3525,N_3659);
nand U4068 (N_4068,N_3996,N_3373);
nor U4069 (N_4069,N_3930,N_3787);
and U4070 (N_4070,N_3931,N_3719);
and U4071 (N_4071,N_3109,N_3691);
nor U4072 (N_4072,N_3681,N_3432);
and U4073 (N_4073,N_3034,N_3807);
nand U4074 (N_4074,N_3428,N_3099);
nand U4075 (N_4075,N_3679,N_3359);
and U4076 (N_4076,N_3479,N_3339);
or U4077 (N_4077,N_3046,N_3863);
or U4078 (N_4078,N_3925,N_3600);
or U4079 (N_4079,N_3243,N_3340);
nand U4080 (N_4080,N_3073,N_3260);
nand U4081 (N_4081,N_3658,N_3177);
nand U4082 (N_4082,N_3044,N_3323);
and U4083 (N_4083,N_3669,N_3636);
nor U4084 (N_4084,N_3401,N_3063);
nand U4085 (N_4085,N_3904,N_3453);
or U4086 (N_4086,N_3909,N_3503);
or U4087 (N_4087,N_3738,N_3675);
nor U4088 (N_4088,N_3580,N_3143);
nor U4089 (N_4089,N_3557,N_3924);
and U4090 (N_4090,N_3149,N_3744);
xnor U4091 (N_4091,N_3389,N_3634);
nor U4092 (N_4092,N_3704,N_3399);
or U4093 (N_4093,N_3165,N_3971);
or U4094 (N_4094,N_3475,N_3973);
and U4095 (N_4095,N_3218,N_3382);
or U4096 (N_4096,N_3684,N_3207);
and U4097 (N_4097,N_3590,N_3010);
nand U4098 (N_4098,N_3958,N_3069);
nor U4099 (N_4099,N_3641,N_3450);
nor U4100 (N_4100,N_3972,N_3570);
and U4101 (N_4101,N_3517,N_3773);
nor U4102 (N_4102,N_3319,N_3604);
nand U4103 (N_4103,N_3587,N_3191);
or U4104 (N_4104,N_3489,N_3029);
nand U4105 (N_4105,N_3713,N_3005);
nor U4106 (N_4106,N_3951,N_3056);
or U4107 (N_4107,N_3491,N_3175);
nor U4108 (N_4108,N_3770,N_3356);
nand U4109 (N_4109,N_3568,N_3174);
or U4110 (N_4110,N_3465,N_3237);
and U4111 (N_4111,N_3740,N_3039);
nand U4112 (N_4112,N_3384,N_3934);
xnor U4113 (N_4113,N_3712,N_3195);
or U4114 (N_4114,N_3483,N_3418);
nor U4115 (N_4115,N_3150,N_3190);
and U4116 (N_4116,N_3688,N_3231);
nor U4117 (N_4117,N_3663,N_3141);
nand U4118 (N_4118,N_3513,N_3901);
nand U4119 (N_4119,N_3806,N_3523);
or U4120 (N_4120,N_3019,N_3745);
or U4121 (N_4121,N_3074,N_3167);
nand U4122 (N_4122,N_3001,N_3090);
nor U4123 (N_4123,N_3752,N_3614);
nand U4124 (N_4124,N_3920,N_3731);
or U4125 (N_4125,N_3027,N_3749);
nand U4126 (N_4126,N_3270,N_3711);
and U4127 (N_4127,N_3308,N_3721);
or U4128 (N_4128,N_3921,N_3945);
nor U4129 (N_4129,N_3358,N_3495);
nand U4130 (N_4130,N_3086,N_3128);
nor U4131 (N_4131,N_3957,N_3347);
or U4132 (N_4132,N_3366,N_3067);
nor U4133 (N_4133,N_3605,N_3474);
nor U4134 (N_4134,N_3698,N_3155);
and U4135 (N_4135,N_3694,N_3420);
or U4136 (N_4136,N_3526,N_3633);
and U4137 (N_4137,N_3268,N_3064);
or U4138 (N_4138,N_3618,N_3181);
nor U4139 (N_4139,N_3997,N_3045);
nand U4140 (N_4140,N_3054,N_3315);
or U4141 (N_4141,N_3157,N_3431);
nand U4142 (N_4142,N_3735,N_3473);
or U4143 (N_4143,N_3959,N_3441);
nand U4144 (N_4144,N_3222,N_3186);
and U4145 (N_4145,N_3089,N_3369);
and U4146 (N_4146,N_3309,N_3018);
or U4147 (N_4147,N_3785,N_3354);
nand U4148 (N_4148,N_3285,N_3346);
or U4149 (N_4149,N_3710,N_3110);
or U4150 (N_4150,N_3892,N_3135);
and U4151 (N_4151,N_3648,N_3558);
nor U4152 (N_4152,N_3834,N_3142);
nor U4153 (N_4153,N_3066,N_3324);
nor U4154 (N_4154,N_3242,N_3581);
nor U4155 (N_4155,N_3012,N_3769);
and U4156 (N_4156,N_3060,N_3327);
nand U4157 (N_4157,N_3626,N_3986);
and U4158 (N_4158,N_3964,N_3091);
nand U4159 (N_4159,N_3795,N_3467);
nor U4160 (N_4160,N_3561,N_3030);
nand U4161 (N_4161,N_3955,N_3662);
or U4162 (N_4162,N_3504,N_3122);
nor U4163 (N_4163,N_3385,N_3727);
and U4164 (N_4164,N_3057,N_3038);
nand U4165 (N_4165,N_3935,N_3272);
and U4166 (N_4166,N_3383,N_3304);
nand U4167 (N_4167,N_3325,N_3397);
nor U4168 (N_4168,N_3543,N_3544);
nand U4169 (N_4169,N_3427,N_3943);
nand U4170 (N_4170,N_3559,N_3779);
nor U4171 (N_4171,N_3154,N_3040);
nand U4172 (N_4172,N_3918,N_3048);
nor U4173 (N_4173,N_3404,N_3937);
and U4174 (N_4174,N_3873,N_3406);
nand U4175 (N_4175,N_3928,N_3541);
or U4176 (N_4176,N_3192,N_3234);
or U4177 (N_4177,N_3932,N_3650);
or U4178 (N_4178,N_3976,N_3828);
or U4179 (N_4179,N_3613,N_3248);
nor U4180 (N_4180,N_3758,N_3117);
and U4181 (N_4181,N_3302,N_3676);
or U4182 (N_4182,N_3638,N_3031);
nand U4183 (N_4183,N_3775,N_3763);
or U4184 (N_4184,N_3173,N_3287);
or U4185 (N_4185,N_3419,N_3516);
or U4186 (N_4186,N_3011,N_3405);
and U4187 (N_4187,N_3303,N_3831);
nor U4188 (N_4188,N_3651,N_3071);
nor U4189 (N_4189,N_3202,N_3125);
nor U4190 (N_4190,N_3584,N_3096);
nor U4191 (N_4191,N_3520,N_3341);
nor U4192 (N_4192,N_3647,N_3777);
xor U4193 (N_4193,N_3172,N_3995);
or U4194 (N_4194,N_3942,N_3227);
nand U4195 (N_4195,N_3657,N_3209);
nand U4196 (N_4196,N_3728,N_3978);
nand U4197 (N_4197,N_3111,N_3497);
nor U4198 (N_4198,N_3300,N_3265);
or U4199 (N_4199,N_3801,N_3847);
nor U4200 (N_4200,N_3510,N_3789);
or U4201 (N_4201,N_3950,N_3910);
nor U4202 (N_4202,N_3351,N_3956);
nand U4203 (N_4203,N_3809,N_3982);
nand U4204 (N_4204,N_3593,N_3764);
and U4205 (N_4205,N_3621,N_3350);
or U4206 (N_4206,N_3630,N_3947);
or U4207 (N_4207,N_3717,N_3606);
and U4208 (N_4208,N_3707,N_3367);
nand U4209 (N_4209,N_3466,N_3571);
nor U4210 (N_4210,N_3238,N_3368);
nor U4211 (N_4211,N_3756,N_3786);
nand U4212 (N_4212,N_3266,N_3871);
nor U4213 (N_4213,N_3887,N_3980);
or U4214 (N_4214,N_3077,N_3199);
or U4215 (N_4215,N_3371,N_3610);
xor U4216 (N_4216,N_3896,N_3989);
nand U4217 (N_4217,N_3579,N_3761);
and U4218 (N_4218,N_3814,N_3741);
nor U4219 (N_4219,N_3414,N_3987);
nor U4220 (N_4220,N_3629,N_3138);
nand U4221 (N_4221,N_3660,N_3422);
nand U4222 (N_4222,N_3458,N_3500);
nor U4223 (N_4223,N_3459,N_3531);
nand U4224 (N_4224,N_3298,N_3824);
nor U4225 (N_4225,N_3290,N_3985);
nand U4226 (N_4226,N_3259,N_3137);
and U4227 (N_4227,N_3435,N_3673);
xor U4228 (N_4228,N_3672,N_3080);
nand U4229 (N_4229,N_3281,N_3878);
nor U4230 (N_4230,N_3519,N_3246);
nand U4231 (N_4231,N_3299,N_3292);
or U4232 (N_4232,N_3860,N_3693);
or U4233 (N_4233,N_3140,N_3189);
nand U4234 (N_4234,N_3378,N_3754);
and U4235 (N_4235,N_3295,N_3008);
nand U4236 (N_4236,N_3848,N_3180);
xnor U4237 (N_4237,N_3940,N_3284);
nand U4238 (N_4238,N_3169,N_3037);
or U4239 (N_4239,N_3521,N_3961);
or U4240 (N_4240,N_3661,N_3355);
and U4241 (N_4241,N_3226,N_3236);
nor U4242 (N_4242,N_3464,N_3869);
nand U4243 (N_4243,N_3042,N_3423);
xor U4244 (N_4244,N_3365,N_3205);
and U4245 (N_4245,N_3468,N_3667);
nor U4246 (N_4246,N_3889,N_3540);
nor U4247 (N_4247,N_3444,N_3993);
nand U4248 (N_4248,N_3724,N_3870);
and U4249 (N_4249,N_3534,N_3927);
or U4250 (N_4250,N_3767,N_3911);
and U4251 (N_4251,N_3898,N_3524);
nand U4252 (N_4252,N_3357,N_3656);
and U4253 (N_4253,N_3588,N_3800);
nor U4254 (N_4254,N_3328,N_3126);
nor U4255 (N_4255,N_3440,N_3463);
or U4256 (N_4256,N_3098,N_3261);
and U4257 (N_4257,N_3885,N_3121);
and U4258 (N_4258,N_3421,N_3219);
or U4259 (N_4259,N_3022,N_3829);
xnor U4260 (N_4260,N_3076,N_3509);
or U4261 (N_4261,N_3762,N_3100);
and U4262 (N_4262,N_3398,N_3637);
and U4263 (N_4263,N_3274,N_3002);
and U4264 (N_4264,N_3866,N_3803);
nand U4265 (N_4265,N_3345,N_3778);
nand U4266 (N_4266,N_3166,N_3914);
nor U4267 (N_4267,N_3546,N_3262);
and U4268 (N_4268,N_3645,N_3050);
and U4269 (N_4269,N_3845,N_3706);
and U4270 (N_4270,N_3537,N_3244);
nand U4271 (N_4271,N_3729,N_3640);
or U4272 (N_4272,N_3810,N_3591);
xor U4273 (N_4273,N_3245,N_3668);
nor U4274 (N_4274,N_3230,N_3084);
xnor U4275 (N_4275,N_3139,N_3204);
and U4276 (N_4276,N_3249,N_3395);
xnor U4277 (N_4277,N_3147,N_3179);
nor U4278 (N_4278,N_3817,N_3229);
nor U4279 (N_4279,N_3518,N_3269);
and U4280 (N_4280,N_3905,N_3788);
nand U4281 (N_4281,N_3289,N_3646);
and U4282 (N_4282,N_3842,N_3239);
and U4283 (N_4283,N_3830,N_3153);
and U4284 (N_4284,N_3696,N_3257);
nor U4285 (N_4285,N_3429,N_3446);
or U4286 (N_4286,N_3742,N_3835);
nor U4287 (N_4287,N_3695,N_3802);
or U4288 (N_4288,N_3277,N_3818);
or U4289 (N_4289,N_3565,N_3412);
nand U4290 (N_4290,N_3095,N_3374);
nor U4291 (N_4291,N_3737,N_3252);
nand U4292 (N_4292,N_3902,N_3020);
nor U4293 (N_4293,N_3082,N_3893);
and U4294 (N_4294,N_3113,N_3258);
nand U4295 (N_4295,N_3822,N_3335);
or U4296 (N_4296,N_3906,N_3849);
or U4297 (N_4297,N_3217,N_3403);
and U4298 (N_4298,N_3447,N_3185);
and U4299 (N_4299,N_3196,N_3628);
xor U4300 (N_4300,N_3460,N_3188);
or U4301 (N_4301,N_3880,N_3726);
or U4302 (N_4302,N_3296,N_3360);
and U4303 (N_4303,N_3334,N_3899);
or U4304 (N_4304,N_3306,N_3213);
or U4305 (N_4305,N_3053,N_3187);
nand U4306 (N_4306,N_3912,N_3305);
and U4307 (N_4307,N_3700,N_3097);
nand U4308 (N_4308,N_3838,N_3352);
or U4309 (N_4309,N_3131,N_3903);
nand U4310 (N_4310,N_3247,N_3677);
nor U4311 (N_4311,N_3983,N_3542);
nand U4312 (N_4312,N_3322,N_3438);
nand U4313 (N_4313,N_3750,N_3781);
or U4314 (N_4314,N_3279,N_3821);
xnor U4315 (N_4315,N_3891,N_3907);
nor U4316 (N_4316,N_3716,N_3757);
nor U4317 (N_4317,N_3413,N_3708);
and U4318 (N_4318,N_3612,N_3578);
nand U4319 (N_4319,N_3755,N_3923);
nand U4320 (N_4320,N_3161,N_3445);
nor U4321 (N_4321,N_3790,N_3678);
or U4322 (N_4322,N_3283,N_3990);
nor U4323 (N_4323,N_3967,N_3966);
and U4324 (N_4324,N_3088,N_3772);
and U4325 (N_4325,N_3023,N_3881);
nor U4326 (N_4326,N_3917,N_3732);
or U4327 (N_4327,N_3093,N_3709);
and U4328 (N_4328,N_3841,N_3362);
and U4329 (N_4329,N_3211,N_3595);
or U4330 (N_4330,N_3563,N_3589);
and U4331 (N_4331,N_3666,N_3390);
or U4332 (N_4332,N_3577,N_3548);
and U4333 (N_4333,N_3282,N_3759);
nor U4334 (N_4334,N_3017,N_3006);
or U4335 (N_4335,N_3566,N_3827);
or U4336 (N_4336,N_3511,N_3505);
nor U4337 (N_4337,N_3649,N_3919);
or U4338 (N_4338,N_3799,N_3624);
nand U4339 (N_4339,N_3114,N_3733);
nand U4340 (N_4340,N_3200,N_3151);
and U4341 (N_4341,N_3338,N_3461);
nor U4342 (N_4342,N_3102,N_3784);
or U4343 (N_4343,N_3974,N_3670);
nand U4344 (N_4344,N_3021,N_3336);
nand U4345 (N_4345,N_3622,N_3212);
nand U4346 (N_4346,N_3815,N_3522);
or U4347 (N_4347,N_3286,N_3094);
and U4348 (N_4348,N_3342,N_3393);
or U4349 (N_4349,N_3016,N_3689);
and U4350 (N_4350,N_3488,N_3556);
nand U4351 (N_4351,N_3233,N_3471);
and U4352 (N_4352,N_3895,N_3416);
nor U4353 (N_4353,N_3939,N_3442);
or U4354 (N_4354,N_3705,N_3051);
nand U4355 (N_4355,N_3083,N_3690);
nand U4356 (N_4356,N_3133,N_3998);
and U4357 (N_4357,N_3451,N_3597);
and U4358 (N_4358,N_3549,N_3394);
nor U4359 (N_4359,N_3882,N_3375);
nor U4360 (N_4360,N_3496,N_3176);
or U4361 (N_4361,N_3583,N_3948);
nor U4362 (N_4362,N_3032,N_3702);
or U4363 (N_4363,N_3620,N_3275);
nor U4364 (N_4364,N_3396,N_3736);
and U4365 (N_4365,N_3119,N_3944);
nor U4366 (N_4366,N_3850,N_3214);
and U4367 (N_4367,N_3506,N_3953);
nor U4368 (N_4368,N_3197,N_3208);
nand U4369 (N_4369,N_3081,N_3232);
nand U4370 (N_4370,N_3946,N_3337);
nor U4371 (N_4371,N_3545,N_3616);
nor U4372 (N_4372,N_3363,N_3766);
and U4373 (N_4373,N_3608,N_3530);
or U4374 (N_4374,N_3687,N_3417);
and U4375 (N_4375,N_3254,N_3832);
and U4376 (N_4376,N_3134,N_3816);
or U4377 (N_4377,N_3623,N_3062);
nor U4378 (N_4378,N_3550,N_3198);
and U4379 (N_4379,N_3223,N_3152);
and U4380 (N_4380,N_3182,N_3457);
nor U4381 (N_4381,N_3857,N_3007);
nor U4382 (N_4382,N_3250,N_3854);
nand U4383 (N_4383,N_3047,N_3224);
nand U4384 (N_4384,N_3168,N_3573);
nor U4385 (N_4385,N_3068,N_3035);
nand U4386 (N_4386,N_3430,N_3533);
or U4387 (N_4387,N_3101,N_3183);
and U4388 (N_4388,N_3791,N_3072);
nor U4389 (N_4389,N_3938,N_3536);
and U4390 (N_4390,N_3436,N_3256);
nand U4391 (N_4391,N_3843,N_3388);
or U4392 (N_4392,N_3136,N_3015);
nor U4393 (N_4393,N_3318,N_3808);
nor U4394 (N_4394,N_3092,N_3743);
nand U4395 (N_4395,N_3963,N_3933);
nand U4396 (N_4396,N_3164,N_3991);
nand U4397 (N_4397,N_3547,N_3852);
and U4398 (N_4398,N_3193,N_3897);
or U4399 (N_4399,N_3498,N_3979);
nand U4400 (N_4400,N_3024,N_3123);
or U4401 (N_4401,N_3201,N_3059);
nand U4402 (N_4402,N_3025,N_3876);
and U4403 (N_4403,N_3760,N_3104);
or U4404 (N_4404,N_3859,N_3798);
or U4405 (N_4405,N_3225,N_3856);
nand U4406 (N_4406,N_3883,N_3267);
or U4407 (N_4407,N_3813,N_3603);
nor U4408 (N_4408,N_3685,N_3108);
nand U4409 (N_4409,N_3567,N_3331);
nor U4410 (N_4410,N_3216,N_3844);
or U4411 (N_4411,N_3400,N_3026);
and U4412 (N_4412,N_3715,N_3635);
and U4413 (N_4413,N_3748,N_3954);
nor U4414 (N_4414,N_3120,N_3402);
or U4415 (N_4415,N_3052,N_3655);
nand U4416 (N_4416,N_3797,N_3449);
or U4417 (N_4417,N_3642,N_3112);
nand U4418 (N_4418,N_3720,N_3280);
nor U4419 (N_4419,N_3344,N_3043);
and U4420 (N_4420,N_3576,N_3379);
nand U4421 (N_4421,N_3532,N_3697);
nand U4422 (N_4422,N_3353,N_3408);
or U4423 (N_4423,N_3145,N_3539);
and U4424 (N_4424,N_3699,N_3041);
nand U4425 (N_4425,N_3643,N_3652);
and U4426 (N_4426,N_3529,N_3853);
or U4427 (N_4427,N_3220,N_3105);
and U4428 (N_4428,N_3858,N_3301);
nand U4429 (N_4429,N_3722,N_3235);
nand U4430 (N_4430,N_3560,N_3241);
nand U4431 (N_4431,N_3409,N_3776);
nand U4432 (N_4432,N_3163,N_3065);
nor U4433 (N_4433,N_3127,N_3751);
nand U4434 (N_4434,N_3425,N_3929);
and U4435 (N_4435,N_3913,N_3314);
nor U4436 (N_4436,N_3926,N_3377);
and U4437 (N_4437,N_3555,N_3884);
nand U4438 (N_4438,N_3313,N_3312);
nand U4439 (N_4439,N_3387,N_3692);
or U4440 (N_4440,N_3049,N_3311);
and U4441 (N_4441,N_3683,N_3796);
nor U4442 (N_4442,N_3569,N_3130);
nor U4443 (N_4443,N_3984,N_3484);
or U4444 (N_4444,N_3836,N_3107);
nor U4445 (N_4445,N_3846,N_3203);
or U4446 (N_4446,N_3619,N_3085);
or U4447 (N_4447,N_3228,N_3507);
nand U4448 (N_4448,N_3528,N_3310);
nand U4449 (N_4449,N_3674,N_3551);
and U4450 (N_4450,N_3864,N_3535);
nor U4451 (N_4451,N_3714,N_3552);
nor U4452 (N_4452,N_3867,N_3411);
nand U4453 (N_4453,N_3118,N_3826);
or U4454 (N_4454,N_3965,N_3819);
nor U4455 (N_4455,N_3320,N_3833);
and U4456 (N_4456,N_3448,N_3861);
and U4457 (N_4457,N_3407,N_3321);
nor U4458 (N_4458,N_3865,N_3601);
nand U4459 (N_4459,N_3462,N_3962);
and U4460 (N_4460,N_3734,N_3490);
nand U4461 (N_4461,N_3485,N_3625);
nor U4462 (N_4462,N_3330,N_3370);
nor U4463 (N_4463,N_3129,N_3527);
nand U4464 (N_4464,N_3682,N_3240);
nor U4465 (N_4465,N_3975,N_3386);
nor U4466 (N_4466,N_3494,N_3215);
and U4467 (N_4467,N_3837,N_3271);
and U4468 (N_4468,N_3703,N_3554);
nor U4469 (N_4469,N_3493,N_3908);
nor U4470 (N_4470,N_3768,N_3210);
or U4471 (N_4471,N_3028,N_3376);
and U4472 (N_4472,N_3426,N_3058);
and U4473 (N_4473,N_3078,N_3730);
or U4474 (N_4474,N_3874,N_3572);
nor U4475 (N_4475,N_3009,N_3170);
nand U4476 (N_4476,N_3805,N_3811);
nand U4477 (N_4477,N_3586,N_3004);
or U4478 (N_4478,N_3970,N_3598);
and U4479 (N_4479,N_3171,N_3003);
nand U4480 (N_4480,N_3723,N_3782);
and U4481 (N_4481,N_3206,N_3115);
or U4482 (N_4482,N_3156,N_3477);
and U4483 (N_4483,N_3653,N_3439);
nand U4484 (N_4484,N_3264,N_3103);
nor U4485 (N_4485,N_3900,N_3627);
nand U4486 (N_4486,N_3992,N_3124);
and U4487 (N_4487,N_3263,N_3501);
and U4488 (N_4488,N_3607,N_3632);
nor U4489 (N_4489,N_3000,N_3492);
nand U4490 (N_4490,N_3877,N_3469);
nand U4491 (N_4491,N_3502,N_3611);
or U4492 (N_4492,N_3916,N_3615);
nor U4493 (N_4493,N_3437,N_3132);
nand U4494 (N_4494,N_3251,N_3644);
or U4495 (N_4495,N_3875,N_3014);
nor U4496 (N_4496,N_3747,N_3033);
or U4497 (N_4497,N_3792,N_3804);
nand U4498 (N_4498,N_3478,N_3872);
and U4499 (N_4499,N_3160,N_3221);
and U4500 (N_4500,N_3308,N_3979);
nor U4501 (N_4501,N_3043,N_3903);
nor U4502 (N_4502,N_3011,N_3752);
nand U4503 (N_4503,N_3118,N_3624);
nand U4504 (N_4504,N_3184,N_3127);
and U4505 (N_4505,N_3296,N_3944);
nor U4506 (N_4506,N_3197,N_3563);
or U4507 (N_4507,N_3545,N_3933);
nor U4508 (N_4508,N_3572,N_3043);
nand U4509 (N_4509,N_3209,N_3204);
nand U4510 (N_4510,N_3777,N_3542);
nor U4511 (N_4511,N_3100,N_3373);
nand U4512 (N_4512,N_3580,N_3563);
nor U4513 (N_4513,N_3593,N_3295);
nand U4514 (N_4514,N_3339,N_3067);
nand U4515 (N_4515,N_3632,N_3535);
nor U4516 (N_4516,N_3733,N_3903);
and U4517 (N_4517,N_3225,N_3179);
or U4518 (N_4518,N_3007,N_3872);
or U4519 (N_4519,N_3441,N_3843);
and U4520 (N_4520,N_3738,N_3808);
nand U4521 (N_4521,N_3143,N_3528);
and U4522 (N_4522,N_3452,N_3078);
and U4523 (N_4523,N_3794,N_3697);
or U4524 (N_4524,N_3753,N_3427);
or U4525 (N_4525,N_3900,N_3100);
nor U4526 (N_4526,N_3768,N_3994);
or U4527 (N_4527,N_3225,N_3568);
or U4528 (N_4528,N_3037,N_3385);
or U4529 (N_4529,N_3240,N_3072);
or U4530 (N_4530,N_3518,N_3243);
nand U4531 (N_4531,N_3086,N_3046);
nor U4532 (N_4532,N_3234,N_3812);
nor U4533 (N_4533,N_3052,N_3960);
or U4534 (N_4534,N_3287,N_3779);
nand U4535 (N_4535,N_3629,N_3690);
nor U4536 (N_4536,N_3189,N_3149);
nor U4537 (N_4537,N_3733,N_3730);
or U4538 (N_4538,N_3867,N_3737);
or U4539 (N_4539,N_3503,N_3820);
or U4540 (N_4540,N_3307,N_3998);
and U4541 (N_4541,N_3675,N_3255);
and U4542 (N_4542,N_3905,N_3814);
xnor U4543 (N_4543,N_3011,N_3258);
nor U4544 (N_4544,N_3121,N_3623);
or U4545 (N_4545,N_3936,N_3865);
and U4546 (N_4546,N_3380,N_3006);
or U4547 (N_4547,N_3818,N_3305);
or U4548 (N_4548,N_3037,N_3831);
and U4549 (N_4549,N_3083,N_3798);
nor U4550 (N_4550,N_3556,N_3518);
nand U4551 (N_4551,N_3746,N_3821);
xnor U4552 (N_4552,N_3124,N_3229);
and U4553 (N_4553,N_3058,N_3446);
xor U4554 (N_4554,N_3402,N_3307);
nor U4555 (N_4555,N_3070,N_3698);
nor U4556 (N_4556,N_3326,N_3705);
nor U4557 (N_4557,N_3424,N_3658);
nor U4558 (N_4558,N_3149,N_3749);
nand U4559 (N_4559,N_3556,N_3210);
or U4560 (N_4560,N_3819,N_3015);
nand U4561 (N_4561,N_3553,N_3208);
nand U4562 (N_4562,N_3389,N_3538);
or U4563 (N_4563,N_3899,N_3662);
and U4564 (N_4564,N_3316,N_3232);
nor U4565 (N_4565,N_3161,N_3328);
nor U4566 (N_4566,N_3983,N_3760);
nand U4567 (N_4567,N_3300,N_3228);
or U4568 (N_4568,N_3183,N_3281);
and U4569 (N_4569,N_3143,N_3808);
or U4570 (N_4570,N_3758,N_3911);
nand U4571 (N_4571,N_3896,N_3537);
and U4572 (N_4572,N_3941,N_3628);
and U4573 (N_4573,N_3381,N_3016);
nor U4574 (N_4574,N_3687,N_3815);
nand U4575 (N_4575,N_3018,N_3941);
nand U4576 (N_4576,N_3594,N_3802);
or U4577 (N_4577,N_3846,N_3125);
or U4578 (N_4578,N_3040,N_3572);
and U4579 (N_4579,N_3164,N_3539);
nand U4580 (N_4580,N_3143,N_3740);
or U4581 (N_4581,N_3324,N_3607);
nand U4582 (N_4582,N_3209,N_3847);
or U4583 (N_4583,N_3898,N_3462);
or U4584 (N_4584,N_3621,N_3306);
nand U4585 (N_4585,N_3132,N_3047);
nand U4586 (N_4586,N_3322,N_3090);
and U4587 (N_4587,N_3653,N_3588);
nand U4588 (N_4588,N_3502,N_3316);
nand U4589 (N_4589,N_3999,N_3006);
nand U4590 (N_4590,N_3266,N_3465);
nand U4591 (N_4591,N_3714,N_3871);
nand U4592 (N_4592,N_3061,N_3248);
nor U4593 (N_4593,N_3129,N_3183);
and U4594 (N_4594,N_3304,N_3796);
nand U4595 (N_4595,N_3843,N_3757);
nor U4596 (N_4596,N_3410,N_3757);
nor U4597 (N_4597,N_3038,N_3478);
nand U4598 (N_4598,N_3095,N_3494);
or U4599 (N_4599,N_3513,N_3236);
and U4600 (N_4600,N_3056,N_3498);
or U4601 (N_4601,N_3753,N_3929);
xor U4602 (N_4602,N_3062,N_3578);
nor U4603 (N_4603,N_3581,N_3855);
nor U4604 (N_4604,N_3313,N_3435);
nand U4605 (N_4605,N_3389,N_3472);
and U4606 (N_4606,N_3747,N_3553);
or U4607 (N_4607,N_3314,N_3839);
nor U4608 (N_4608,N_3483,N_3370);
and U4609 (N_4609,N_3869,N_3527);
nand U4610 (N_4610,N_3258,N_3303);
nor U4611 (N_4611,N_3938,N_3047);
or U4612 (N_4612,N_3446,N_3288);
and U4613 (N_4613,N_3403,N_3629);
or U4614 (N_4614,N_3133,N_3842);
nand U4615 (N_4615,N_3777,N_3562);
and U4616 (N_4616,N_3489,N_3552);
xnor U4617 (N_4617,N_3355,N_3487);
nor U4618 (N_4618,N_3878,N_3232);
nor U4619 (N_4619,N_3251,N_3459);
and U4620 (N_4620,N_3440,N_3057);
or U4621 (N_4621,N_3227,N_3047);
and U4622 (N_4622,N_3112,N_3594);
or U4623 (N_4623,N_3872,N_3277);
nor U4624 (N_4624,N_3072,N_3794);
or U4625 (N_4625,N_3363,N_3622);
or U4626 (N_4626,N_3252,N_3832);
and U4627 (N_4627,N_3556,N_3199);
and U4628 (N_4628,N_3497,N_3555);
or U4629 (N_4629,N_3123,N_3104);
nor U4630 (N_4630,N_3165,N_3336);
nand U4631 (N_4631,N_3072,N_3526);
nand U4632 (N_4632,N_3183,N_3816);
and U4633 (N_4633,N_3340,N_3241);
nand U4634 (N_4634,N_3131,N_3375);
or U4635 (N_4635,N_3275,N_3712);
nor U4636 (N_4636,N_3680,N_3372);
nor U4637 (N_4637,N_3095,N_3650);
nor U4638 (N_4638,N_3034,N_3885);
nand U4639 (N_4639,N_3077,N_3690);
nor U4640 (N_4640,N_3882,N_3422);
nor U4641 (N_4641,N_3892,N_3153);
and U4642 (N_4642,N_3562,N_3585);
nand U4643 (N_4643,N_3423,N_3260);
nand U4644 (N_4644,N_3136,N_3108);
and U4645 (N_4645,N_3933,N_3016);
nand U4646 (N_4646,N_3674,N_3736);
nor U4647 (N_4647,N_3492,N_3041);
nand U4648 (N_4648,N_3122,N_3130);
nand U4649 (N_4649,N_3546,N_3825);
nand U4650 (N_4650,N_3820,N_3421);
or U4651 (N_4651,N_3454,N_3691);
and U4652 (N_4652,N_3343,N_3261);
and U4653 (N_4653,N_3782,N_3971);
and U4654 (N_4654,N_3867,N_3477);
nand U4655 (N_4655,N_3394,N_3270);
nand U4656 (N_4656,N_3868,N_3907);
or U4657 (N_4657,N_3473,N_3049);
and U4658 (N_4658,N_3078,N_3544);
and U4659 (N_4659,N_3284,N_3587);
nand U4660 (N_4660,N_3778,N_3295);
nor U4661 (N_4661,N_3380,N_3463);
nor U4662 (N_4662,N_3377,N_3468);
and U4663 (N_4663,N_3796,N_3953);
and U4664 (N_4664,N_3968,N_3797);
nand U4665 (N_4665,N_3604,N_3819);
nor U4666 (N_4666,N_3347,N_3825);
or U4667 (N_4667,N_3805,N_3586);
and U4668 (N_4668,N_3368,N_3703);
and U4669 (N_4669,N_3704,N_3662);
and U4670 (N_4670,N_3474,N_3801);
xnor U4671 (N_4671,N_3195,N_3232);
or U4672 (N_4672,N_3417,N_3592);
or U4673 (N_4673,N_3173,N_3290);
nand U4674 (N_4674,N_3248,N_3359);
and U4675 (N_4675,N_3077,N_3874);
or U4676 (N_4676,N_3829,N_3472);
nand U4677 (N_4677,N_3771,N_3656);
xor U4678 (N_4678,N_3970,N_3666);
nor U4679 (N_4679,N_3934,N_3557);
and U4680 (N_4680,N_3781,N_3964);
nor U4681 (N_4681,N_3319,N_3621);
and U4682 (N_4682,N_3269,N_3522);
and U4683 (N_4683,N_3175,N_3996);
nand U4684 (N_4684,N_3372,N_3292);
nor U4685 (N_4685,N_3055,N_3811);
nor U4686 (N_4686,N_3815,N_3952);
and U4687 (N_4687,N_3946,N_3485);
nand U4688 (N_4688,N_3211,N_3431);
and U4689 (N_4689,N_3095,N_3521);
nor U4690 (N_4690,N_3049,N_3991);
nand U4691 (N_4691,N_3914,N_3574);
and U4692 (N_4692,N_3432,N_3528);
nor U4693 (N_4693,N_3807,N_3371);
nand U4694 (N_4694,N_3827,N_3593);
nand U4695 (N_4695,N_3666,N_3605);
nor U4696 (N_4696,N_3916,N_3707);
nand U4697 (N_4697,N_3650,N_3195);
or U4698 (N_4698,N_3337,N_3458);
or U4699 (N_4699,N_3355,N_3287);
and U4700 (N_4700,N_3890,N_3122);
nand U4701 (N_4701,N_3248,N_3189);
or U4702 (N_4702,N_3216,N_3808);
and U4703 (N_4703,N_3037,N_3953);
nand U4704 (N_4704,N_3970,N_3463);
nor U4705 (N_4705,N_3704,N_3018);
nand U4706 (N_4706,N_3258,N_3328);
nor U4707 (N_4707,N_3594,N_3433);
and U4708 (N_4708,N_3244,N_3081);
xor U4709 (N_4709,N_3658,N_3155);
and U4710 (N_4710,N_3853,N_3041);
nand U4711 (N_4711,N_3823,N_3739);
nand U4712 (N_4712,N_3010,N_3160);
and U4713 (N_4713,N_3371,N_3629);
nand U4714 (N_4714,N_3018,N_3127);
or U4715 (N_4715,N_3380,N_3805);
or U4716 (N_4716,N_3670,N_3503);
and U4717 (N_4717,N_3454,N_3391);
and U4718 (N_4718,N_3599,N_3931);
nand U4719 (N_4719,N_3215,N_3112);
and U4720 (N_4720,N_3083,N_3610);
or U4721 (N_4721,N_3993,N_3371);
or U4722 (N_4722,N_3671,N_3971);
or U4723 (N_4723,N_3077,N_3391);
nor U4724 (N_4724,N_3358,N_3802);
nor U4725 (N_4725,N_3381,N_3100);
or U4726 (N_4726,N_3089,N_3374);
and U4727 (N_4727,N_3464,N_3200);
or U4728 (N_4728,N_3412,N_3868);
nor U4729 (N_4729,N_3683,N_3384);
and U4730 (N_4730,N_3763,N_3472);
or U4731 (N_4731,N_3069,N_3798);
or U4732 (N_4732,N_3801,N_3527);
nand U4733 (N_4733,N_3862,N_3669);
nand U4734 (N_4734,N_3906,N_3450);
nand U4735 (N_4735,N_3117,N_3795);
or U4736 (N_4736,N_3496,N_3361);
and U4737 (N_4737,N_3982,N_3534);
nor U4738 (N_4738,N_3854,N_3619);
or U4739 (N_4739,N_3940,N_3224);
or U4740 (N_4740,N_3240,N_3592);
xor U4741 (N_4741,N_3549,N_3644);
nand U4742 (N_4742,N_3356,N_3426);
and U4743 (N_4743,N_3947,N_3473);
or U4744 (N_4744,N_3286,N_3722);
or U4745 (N_4745,N_3119,N_3067);
nor U4746 (N_4746,N_3217,N_3053);
nand U4747 (N_4747,N_3594,N_3058);
or U4748 (N_4748,N_3958,N_3358);
or U4749 (N_4749,N_3724,N_3663);
nand U4750 (N_4750,N_3605,N_3221);
or U4751 (N_4751,N_3425,N_3409);
or U4752 (N_4752,N_3006,N_3793);
and U4753 (N_4753,N_3881,N_3024);
nand U4754 (N_4754,N_3230,N_3292);
or U4755 (N_4755,N_3529,N_3557);
nand U4756 (N_4756,N_3521,N_3566);
and U4757 (N_4757,N_3732,N_3592);
nor U4758 (N_4758,N_3634,N_3423);
and U4759 (N_4759,N_3824,N_3045);
and U4760 (N_4760,N_3416,N_3561);
and U4761 (N_4761,N_3979,N_3743);
nor U4762 (N_4762,N_3800,N_3307);
or U4763 (N_4763,N_3383,N_3397);
and U4764 (N_4764,N_3900,N_3846);
or U4765 (N_4765,N_3243,N_3784);
nand U4766 (N_4766,N_3859,N_3195);
nand U4767 (N_4767,N_3794,N_3103);
or U4768 (N_4768,N_3737,N_3273);
nor U4769 (N_4769,N_3642,N_3171);
nand U4770 (N_4770,N_3695,N_3214);
nor U4771 (N_4771,N_3216,N_3352);
nand U4772 (N_4772,N_3672,N_3466);
nor U4773 (N_4773,N_3897,N_3665);
or U4774 (N_4774,N_3752,N_3051);
and U4775 (N_4775,N_3254,N_3464);
or U4776 (N_4776,N_3910,N_3204);
nand U4777 (N_4777,N_3697,N_3493);
or U4778 (N_4778,N_3586,N_3704);
or U4779 (N_4779,N_3785,N_3071);
or U4780 (N_4780,N_3202,N_3631);
and U4781 (N_4781,N_3138,N_3183);
nand U4782 (N_4782,N_3725,N_3169);
nand U4783 (N_4783,N_3876,N_3952);
nor U4784 (N_4784,N_3047,N_3987);
or U4785 (N_4785,N_3074,N_3115);
and U4786 (N_4786,N_3911,N_3252);
xor U4787 (N_4787,N_3609,N_3476);
nand U4788 (N_4788,N_3378,N_3517);
nor U4789 (N_4789,N_3164,N_3955);
and U4790 (N_4790,N_3461,N_3964);
and U4791 (N_4791,N_3194,N_3036);
and U4792 (N_4792,N_3740,N_3392);
xor U4793 (N_4793,N_3818,N_3416);
and U4794 (N_4794,N_3358,N_3426);
nor U4795 (N_4795,N_3781,N_3475);
or U4796 (N_4796,N_3052,N_3346);
or U4797 (N_4797,N_3712,N_3833);
nand U4798 (N_4798,N_3328,N_3367);
nand U4799 (N_4799,N_3997,N_3111);
nand U4800 (N_4800,N_3257,N_3565);
and U4801 (N_4801,N_3920,N_3528);
nand U4802 (N_4802,N_3750,N_3470);
and U4803 (N_4803,N_3237,N_3374);
nand U4804 (N_4804,N_3091,N_3707);
nand U4805 (N_4805,N_3070,N_3044);
nand U4806 (N_4806,N_3640,N_3258);
and U4807 (N_4807,N_3507,N_3746);
nor U4808 (N_4808,N_3460,N_3040);
nor U4809 (N_4809,N_3180,N_3978);
nand U4810 (N_4810,N_3791,N_3959);
and U4811 (N_4811,N_3709,N_3588);
or U4812 (N_4812,N_3226,N_3487);
nand U4813 (N_4813,N_3734,N_3924);
or U4814 (N_4814,N_3766,N_3195);
nand U4815 (N_4815,N_3856,N_3152);
nand U4816 (N_4816,N_3467,N_3592);
or U4817 (N_4817,N_3092,N_3675);
or U4818 (N_4818,N_3743,N_3215);
nor U4819 (N_4819,N_3400,N_3555);
xor U4820 (N_4820,N_3550,N_3061);
nor U4821 (N_4821,N_3555,N_3885);
or U4822 (N_4822,N_3935,N_3516);
nor U4823 (N_4823,N_3895,N_3647);
and U4824 (N_4824,N_3645,N_3302);
nand U4825 (N_4825,N_3077,N_3554);
nand U4826 (N_4826,N_3369,N_3080);
or U4827 (N_4827,N_3813,N_3639);
nor U4828 (N_4828,N_3089,N_3623);
and U4829 (N_4829,N_3886,N_3726);
and U4830 (N_4830,N_3303,N_3976);
or U4831 (N_4831,N_3140,N_3175);
xnor U4832 (N_4832,N_3405,N_3971);
or U4833 (N_4833,N_3490,N_3601);
nand U4834 (N_4834,N_3622,N_3371);
or U4835 (N_4835,N_3052,N_3067);
or U4836 (N_4836,N_3768,N_3098);
and U4837 (N_4837,N_3240,N_3886);
or U4838 (N_4838,N_3857,N_3390);
or U4839 (N_4839,N_3444,N_3966);
nand U4840 (N_4840,N_3850,N_3711);
and U4841 (N_4841,N_3745,N_3936);
nor U4842 (N_4842,N_3684,N_3698);
and U4843 (N_4843,N_3323,N_3433);
nand U4844 (N_4844,N_3984,N_3380);
or U4845 (N_4845,N_3667,N_3184);
or U4846 (N_4846,N_3461,N_3325);
nand U4847 (N_4847,N_3467,N_3393);
and U4848 (N_4848,N_3434,N_3933);
or U4849 (N_4849,N_3757,N_3972);
and U4850 (N_4850,N_3280,N_3830);
nand U4851 (N_4851,N_3834,N_3586);
xnor U4852 (N_4852,N_3261,N_3235);
or U4853 (N_4853,N_3025,N_3653);
and U4854 (N_4854,N_3699,N_3580);
or U4855 (N_4855,N_3089,N_3429);
xor U4856 (N_4856,N_3392,N_3413);
or U4857 (N_4857,N_3964,N_3332);
or U4858 (N_4858,N_3000,N_3038);
nor U4859 (N_4859,N_3478,N_3540);
and U4860 (N_4860,N_3247,N_3047);
nand U4861 (N_4861,N_3926,N_3201);
nor U4862 (N_4862,N_3411,N_3623);
and U4863 (N_4863,N_3920,N_3727);
and U4864 (N_4864,N_3473,N_3115);
and U4865 (N_4865,N_3226,N_3349);
or U4866 (N_4866,N_3034,N_3471);
nand U4867 (N_4867,N_3869,N_3707);
or U4868 (N_4868,N_3414,N_3977);
nor U4869 (N_4869,N_3742,N_3079);
nor U4870 (N_4870,N_3809,N_3377);
or U4871 (N_4871,N_3884,N_3428);
or U4872 (N_4872,N_3195,N_3917);
and U4873 (N_4873,N_3749,N_3271);
or U4874 (N_4874,N_3733,N_3520);
or U4875 (N_4875,N_3364,N_3351);
or U4876 (N_4876,N_3988,N_3063);
and U4877 (N_4877,N_3847,N_3483);
nor U4878 (N_4878,N_3840,N_3154);
and U4879 (N_4879,N_3270,N_3460);
or U4880 (N_4880,N_3492,N_3413);
nand U4881 (N_4881,N_3442,N_3773);
or U4882 (N_4882,N_3868,N_3416);
or U4883 (N_4883,N_3141,N_3394);
nor U4884 (N_4884,N_3895,N_3659);
or U4885 (N_4885,N_3302,N_3316);
and U4886 (N_4886,N_3885,N_3426);
nand U4887 (N_4887,N_3467,N_3362);
nor U4888 (N_4888,N_3310,N_3157);
and U4889 (N_4889,N_3382,N_3469);
xor U4890 (N_4890,N_3814,N_3054);
nor U4891 (N_4891,N_3153,N_3136);
or U4892 (N_4892,N_3237,N_3820);
nand U4893 (N_4893,N_3081,N_3055);
or U4894 (N_4894,N_3945,N_3166);
and U4895 (N_4895,N_3364,N_3654);
nor U4896 (N_4896,N_3365,N_3284);
nand U4897 (N_4897,N_3009,N_3930);
nor U4898 (N_4898,N_3119,N_3676);
nor U4899 (N_4899,N_3729,N_3699);
or U4900 (N_4900,N_3127,N_3623);
nand U4901 (N_4901,N_3746,N_3074);
nand U4902 (N_4902,N_3010,N_3775);
xor U4903 (N_4903,N_3145,N_3580);
nor U4904 (N_4904,N_3087,N_3930);
and U4905 (N_4905,N_3168,N_3551);
nor U4906 (N_4906,N_3651,N_3072);
nand U4907 (N_4907,N_3640,N_3766);
nor U4908 (N_4908,N_3003,N_3446);
or U4909 (N_4909,N_3526,N_3547);
and U4910 (N_4910,N_3464,N_3126);
or U4911 (N_4911,N_3002,N_3787);
or U4912 (N_4912,N_3501,N_3016);
and U4913 (N_4913,N_3775,N_3850);
nand U4914 (N_4914,N_3210,N_3036);
xor U4915 (N_4915,N_3910,N_3573);
nand U4916 (N_4916,N_3314,N_3565);
or U4917 (N_4917,N_3067,N_3136);
nand U4918 (N_4918,N_3286,N_3944);
nand U4919 (N_4919,N_3598,N_3811);
and U4920 (N_4920,N_3042,N_3869);
nor U4921 (N_4921,N_3176,N_3343);
and U4922 (N_4922,N_3762,N_3978);
and U4923 (N_4923,N_3119,N_3972);
and U4924 (N_4924,N_3224,N_3550);
or U4925 (N_4925,N_3210,N_3743);
and U4926 (N_4926,N_3786,N_3180);
or U4927 (N_4927,N_3303,N_3923);
and U4928 (N_4928,N_3709,N_3642);
nand U4929 (N_4929,N_3092,N_3468);
nand U4930 (N_4930,N_3393,N_3825);
and U4931 (N_4931,N_3947,N_3719);
or U4932 (N_4932,N_3296,N_3667);
xor U4933 (N_4933,N_3468,N_3786);
or U4934 (N_4934,N_3751,N_3708);
or U4935 (N_4935,N_3953,N_3239);
nor U4936 (N_4936,N_3021,N_3853);
or U4937 (N_4937,N_3233,N_3328);
nand U4938 (N_4938,N_3730,N_3484);
nand U4939 (N_4939,N_3047,N_3559);
or U4940 (N_4940,N_3573,N_3095);
nand U4941 (N_4941,N_3150,N_3775);
or U4942 (N_4942,N_3593,N_3778);
or U4943 (N_4943,N_3628,N_3340);
nor U4944 (N_4944,N_3022,N_3474);
nand U4945 (N_4945,N_3956,N_3120);
or U4946 (N_4946,N_3687,N_3341);
and U4947 (N_4947,N_3323,N_3764);
or U4948 (N_4948,N_3327,N_3034);
and U4949 (N_4949,N_3625,N_3814);
nand U4950 (N_4950,N_3591,N_3331);
or U4951 (N_4951,N_3248,N_3662);
or U4952 (N_4952,N_3287,N_3413);
and U4953 (N_4953,N_3024,N_3457);
nand U4954 (N_4954,N_3023,N_3983);
nor U4955 (N_4955,N_3800,N_3763);
and U4956 (N_4956,N_3419,N_3823);
nor U4957 (N_4957,N_3774,N_3663);
nand U4958 (N_4958,N_3579,N_3551);
or U4959 (N_4959,N_3921,N_3843);
nand U4960 (N_4960,N_3557,N_3390);
or U4961 (N_4961,N_3812,N_3957);
nor U4962 (N_4962,N_3305,N_3703);
and U4963 (N_4963,N_3955,N_3925);
nand U4964 (N_4964,N_3396,N_3880);
or U4965 (N_4965,N_3352,N_3088);
and U4966 (N_4966,N_3901,N_3887);
and U4967 (N_4967,N_3749,N_3649);
or U4968 (N_4968,N_3927,N_3376);
nand U4969 (N_4969,N_3291,N_3669);
nand U4970 (N_4970,N_3168,N_3748);
nor U4971 (N_4971,N_3284,N_3240);
or U4972 (N_4972,N_3255,N_3188);
nand U4973 (N_4973,N_3793,N_3369);
and U4974 (N_4974,N_3071,N_3035);
nand U4975 (N_4975,N_3118,N_3377);
and U4976 (N_4976,N_3941,N_3370);
nand U4977 (N_4977,N_3144,N_3933);
nand U4978 (N_4978,N_3415,N_3442);
nand U4979 (N_4979,N_3594,N_3413);
nand U4980 (N_4980,N_3534,N_3119);
xor U4981 (N_4981,N_3547,N_3501);
or U4982 (N_4982,N_3540,N_3789);
or U4983 (N_4983,N_3090,N_3251);
nand U4984 (N_4984,N_3414,N_3964);
and U4985 (N_4985,N_3296,N_3153);
nor U4986 (N_4986,N_3849,N_3154);
nand U4987 (N_4987,N_3127,N_3428);
nand U4988 (N_4988,N_3528,N_3871);
nand U4989 (N_4989,N_3426,N_3309);
or U4990 (N_4990,N_3337,N_3188);
and U4991 (N_4991,N_3314,N_3074);
and U4992 (N_4992,N_3121,N_3312);
and U4993 (N_4993,N_3301,N_3700);
nand U4994 (N_4994,N_3209,N_3189);
or U4995 (N_4995,N_3787,N_3329);
nor U4996 (N_4996,N_3573,N_3915);
nand U4997 (N_4997,N_3791,N_3569);
nand U4998 (N_4998,N_3185,N_3253);
and U4999 (N_4999,N_3695,N_3094);
nor U5000 (N_5000,N_4997,N_4722);
nor U5001 (N_5001,N_4984,N_4256);
nand U5002 (N_5002,N_4601,N_4313);
nand U5003 (N_5003,N_4198,N_4671);
and U5004 (N_5004,N_4065,N_4149);
or U5005 (N_5005,N_4236,N_4834);
and U5006 (N_5006,N_4818,N_4152);
or U5007 (N_5007,N_4320,N_4993);
nand U5008 (N_5008,N_4892,N_4417);
nor U5009 (N_5009,N_4400,N_4630);
and U5010 (N_5010,N_4060,N_4334);
nand U5011 (N_5011,N_4962,N_4861);
nand U5012 (N_5012,N_4484,N_4944);
nor U5013 (N_5013,N_4987,N_4946);
nand U5014 (N_5014,N_4702,N_4415);
or U5015 (N_5015,N_4479,N_4387);
and U5016 (N_5016,N_4240,N_4838);
or U5017 (N_5017,N_4816,N_4524);
nand U5018 (N_5018,N_4475,N_4136);
and U5019 (N_5019,N_4683,N_4881);
or U5020 (N_5020,N_4604,N_4914);
nor U5021 (N_5021,N_4158,N_4583);
and U5022 (N_5022,N_4287,N_4961);
nor U5023 (N_5023,N_4602,N_4481);
or U5024 (N_5024,N_4598,N_4275);
nor U5025 (N_5025,N_4751,N_4628);
nor U5026 (N_5026,N_4770,N_4178);
nand U5027 (N_5027,N_4510,N_4373);
nand U5028 (N_5028,N_4954,N_4804);
nand U5029 (N_5029,N_4703,N_4335);
or U5030 (N_5030,N_4821,N_4966);
and U5031 (N_5031,N_4412,N_4805);
and U5032 (N_5032,N_4979,N_4483);
nor U5033 (N_5033,N_4221,N_4402);
and U5034 (N_5034,N_4740,N_4000);
nor U5035 (N_5035,N_4778,N_4720);
or U5036 (N_5036,N_4064,N_4612);
nor U5037 (N_5037,N_4904,N_4390);
or U5038 (N_5038,N_4348,N_4406);
nand U5039 (N_5039,N_4124,N_4786);
and U5040 (N_5040,N_4358,N_4186);
nand U5041 (N_5041,N_4204,N_4874);
or U5042 (N_5042,N_4854,N_4977);
or U5043 (N_5043,N_4968,N_4935);
and U5044 (N_5044,N_4055,N_4949);
nor U5045 (N_5045,N_4888,N_4127);
and U5046 (N_5046,N_4418,N_4921);
and U5047 (N_5047,N_4643,N_4650);
nor U5048 (N_5048,N_4285,N_4337);
nand U5049 (N_5049,N_4440,N_4659);
nand U5050 (N_5050,N_4085,N_4355);
nor U5051 (N_5051,N_4254,N_4880);
and U5052 (N_5052,N_4123,N_4163);
and U5053 (N_5053,N_4265,N_4772);
nor U5054 (N_5054,N_4174,N_4010);
xnor U5055 (N_5055,N_4663,N_4242);
nand U5056 (N_5056,N_4948,N_4468);
and U5057 (N_5057,N_4815,N_4326);
and U5058 (N_5058,N_4655,N_4088);
and U5059 (N_5059,N_4782,N_4523);
and U5060 (N_5060,N_4514,N_4747);
nor U5061 (N_5061,N_4025,N_4437);
nand U5062 (N_5062,N_4268,N_4789);
or U5063 (N_5063,N_4809,N_4687);
nor U5064 (N_5064,N_4783,N_4021);
nand U5065 (N_5065,N_4392,N_4905);
nor U5066 (N_5066,N_4425,N_4623);
nand U5067 (N_5067,N_4258,N_4332);
or U5068 (N_5068,N_4657,N_4513);
and U5069 (N_5069,N_4231,N_4384);
nand U5070 (N_5070,N_4173,N_4336);
nor U5071 (N_5071,N_4714,N_4252);
nor U5072 (N_5072,N_4379,N_4781);
nand U5073 (N_5073,N_4865,N_4758);
and U5074 (N_5074,N_4063,N_4721);
or U5075 (N_5075,N_4385,N_4718);
or U5076 (N_5076,N_4274,N_4677);
or U5077 (N_5077,N_4129,N_4044);
and U5078 (N_5078,N_4591,N_4796);
or U5079 (N_5079,N_4398,N_4201);
nor U5080 (N_5080,N_4419,N_4244);
nor U5081 (N_5081,N_4450,N_4199);
and U5082 (N_5082,N_4900,N_4713);
or U5083 (N_5083,N_4383,N_4208);
and U5084 (N_5084,N_4295,N_4726);
nor U5085 (N_5085,N_4491,N_4451);
nor U5086 (N_5086,N_4704,N_4863);
or U5087 (N_5087,N_4787,N_4641);
or U5088 (N_5088,N_4067,N_4100);
or U5089 (N_5089,N_4853,N_4835);
nand U5090 (N_5090,N_4742,N_4631);
nand U5091 (N_5091,N_4812,N_4730);
and U5092 (N_5092,N_4422,N_4975);
nor U5093 (N_5093,N_4446,N_4108);
nand U5094 (N_5094,N_4517,N_4745);
nand U5095 (N_5095,N_4988,N_4616);
nor U5096 (N_5096,N_4386,N_4648);
nand U5097 (N_5097,N_4506,N_4822);
nand U5098 (N_5098,N_4859,N_4994);
nand U5099 (N_5099,N_4073,N_4070);
nor U5100 (N_5100,N_4211,N_4288);
nand U5101 (N_5101,N_4773,N_4985);
and U5102 (N_5102,N_4875,N_4139);
nand U5103 (N_5103,N_4530,N_4543);
nor U5104 (N_5104,N_4272,N_4986);
and U5105 (N_5105,N_4008,N_4699);
nand U5106 (N_5106,N_4195,N_4637);
nor U5107 (N_5107,N_4515,N_4184);
nand U5108 (N_5108,N_4339,N_4982);
nand U5109 (N_5109,N_4978,N_4028);
and U5110 (N_5110,N_4929,N_4856);
or U5111 (N_5111,N_4364,N_4825);
and U5112 (N_5112,N_4462,N_4370);
nand U5113 (N_5113,N_4308,N_4014);
nor U5114 (N_5114,N_4595,N_4545);
or U5115 (N_5115,N_4790,N_4216);
nor U5116 (N_5116,N_4556,N_4585);
nand U5117 (N_5117,N_4849,N_4711);
and U5118 (N_5118,N_4759,N_4573);
or U5119 (N_5119,N_4052,N_4891);
nand U5120 (N_5120,N_4306,N_4951);
nand U5121 (N_5121,N_4066,N_4867);
nor U5122 (N_5122,N_4463,N_4666);
nand U5123 (N_5123,N_4305,N_4338);
and U5124 (N_5124,N_4138,N_4460);
nor U5125 (N_5125,N_4518,N_4056);
xnor U5126 (N_5126,N_4668,N_4624);
nor U5127 (N_5127,N_4762,N_4920);
nand U5128 (N_5128,N_4323,N_4399);
or U5129 (N_5129,N_4145,N_4860);
nor U5130 (N_5130,N_4899,N_4942);
nor U5131 (N_5131,N_4030,N_4766);
nand U5132 (N_5132,N_4095,N_4439);
nand U5133 (N_5133,N_4238,N_4661);
or U5134 (N_5134,N_4841,N_4527);
nor U5135 (N_5135,N_4317,N_4411);
nand U5136 (N_5136,N_4377,N_4808);
nand U5137 (N_5137,N_4688,N_4043);
and U5138 (N_5138,N_4345,N_4910);
nor U5139 (N_5139,N_4423,N_4858);
or U5140 (N_5140,N_4269,N_4576);
and U5141 (N_5141,N_4126,N_4069);
nor U5142 (N_5142,N_4474,N_4396);
and U5143 (N_5143,N_4803,N_4632);
nand U5144 (N_5144,N_4852,N_4130);
and U5145 (N_5145,N_4473,N_4389);
xnor U5146 (N_5146,N_4205,N_4071);
nor U5147 (N_5147,N_4405,N_4375);
or U5148 (N_5148,N_4015,N_4685);
nand U5149 (N_5149,N_4554,N_4734);
and U5150 (N_5150,N_4047,N_4083);
nor U5151 (N_5151,N_4270,N_4072);
nand U5152 (N_5152,N_4998,N_4404);
and U5153 (N_5153,N_4729,N_4110);
or U5154 (N_5154,N_4652,N_4087);
nand U5155 (N_5155,N_4525,N_4090);
or U5156 (N_5156,N_4393,N_4099);
nand U5157 (N_5157,N_4035,N_4864);
or U5158 (N_5158,N_4033,N_4538);
nand U5159 (N_5159,N_4784,N_4459);
or U5160 (N_5160,N_4774,N_4349);
and U5161 (N_5161,N_4619,N_4395);
nor U5162 (N_5162,N_4112,N_4508);
and U5163 (N_5163,N_4266,N_4048);
or U5164 (N_5164,N_4298,N_4885);
and U5165 (N_5165,N_4469,N_4731);
and U5166 (N_5166,N_4182,N_4420);
or U5167 (N_5167,N_4519,N_4464);
and U5168 (N_5168,N_4259,N_4520);
nor U5169 (N_5169,N_4571,N_4817);
or U5170 (N_5170,N_4811,N_4019);
nand U5171 (N_5171,N_4026,N_4561);
and U5172 (N_5172,N_4613,N_4441);
nand U5173 (N_5173,N_4160,N_4369);
or U5174 (N_5174,N_4599,N_4147);
nand U5175 (N_5175,N_4009,N_4889);
and U5176 (N_5176,N_4144,N_4780);
nand U5177 (N_5177,N_4156,N_4116);
and U5178 (N_5178,N_4995,N_4558);
nand U5179 (N_5179,N_4228,N_4103);
and U5180 (N_5180,N_4465,N_4963);
nand U5181 (N_5181,N_4159,N_4569);
or U5182 (N_5182,N_4357,N_4024);
and U5183 (N_5183,N_4365,N_4246);
or U5184 (N_5184,N_4600,N_4448);
or U5185 (N_5185,N_4798,N_4454);
or U5186 (N_5186,N_4102,N_4477);
xor U5187 (N_5187,N_4091,N_4115);
or U5188 (N_5188,N_4260,N_4820);
and U5189 (N_5189,N_4939,N_4727);
or U5190 (N_5190,N_4344,N_4132);
nor U5191 (N_5191,N_4027,N_4432);
nor U5192 (N_5192,N_4267,N_4225);
or U5193 (N_5193,N_4907,N_4281);
and U5194 (N_5194,N_4895,N_4372);
and U5195 (N_5195,N_4764,N_4074);
xor U5196 (N_5196,N_4621,N_4763);
or U5197 (N_5197,N_4190,N_4125);
and U5198 (N_5198,N_4273,N_4879);
nand U5199 (N_5199,N_4597,N_4844);
nor U5200 (N_5200,N_4094,N_4707);
and U5201 (N_5201,N_4593,N_4857);
and U5202 (N_5202,N_4941,N_4117);
nand U5203 (N_5203,N_4709,N_4622);
or U5204 (N_5204,N_4614,N_4098);
xor U5205 (N_5205,N_4578,N_4376);
nand U5206 (N_5206,N_4674,N_4931);
and U5207 (N_5207,N_4807,N_4059);
or U5208 (N_5208,N_4194,N_4492);
or U5209 (N_5209,N_4222,N_4006);
nor U5210 (N_5210,N_4493,N_4936);
and U5211 (N_5211,N_4113,N_4916);
nand U5212 (N_5212,N_4855,N_4947);
nor U5213 (N_5213,N_4728,N_4560);
nor U5214 (N_5214,N_4470,N_4366);
nand U5215 (N_5215,N_4733,N_4592);
and U5216 (N_5216,N_4175,N_4413);
or U5217 (N_5217,N_4062,N_4906);
or U5218 (N_5218,N_4280,N_4594);
and U5219 (N_5219,N_4361,N_4924);
or U5220 (N_5220,N_4188,N_4029);
or U5221 (N_5221,N_4325,N_4176);
and U5222 (N_5222,N_4548,N_4893);
nor U5223 (N_5223,N_4118,N_4151);
nand U5224 (N_5224,N_4953,N_4401);
nand U5225 (N_5225,N_4536,N_4250);
nand U5226 (N_5226,N_4956,N_4495);
and U5227 (N_5227,N_4509,N_4832);
nor U5228 (N_5228,N_4223,N_4967);
nand U5229 (N_5229,N_4570,N_4629);
and U5230 (N_5230,N_4237,N_4664);
and U5231 (N_5231,N_4847,N_4665);
nor U5232 (N_5232,N_4209,N_4011);
and U5233 (N_5233,N_4767,N_4206);
nor U5234 (N_5234,N_4533,N_4625);
and U5235 (N_5235,N_4938,N_4397);
nor U5236 (N_5236,N_4603,N_4486);
and U5237 (N_5237,N_4283,N_4974);
or U5238 (N_5238,N_4753,N_4324);
or U5239 (N_5239,N_4980,N_4981);
nand U5240 (N_5240,N_4693,N_4913);
and U5241 (N_5241,N_4076,N_4568);
nor U5242 (N_5242,N_4467,N_4292);
nand U5243 (N_5243,N_4732,N_4449);
and U5244 (N_5244,N_4848,N_4590);
or U5245 (N_5245,N_4919,N_4219);
nand U5246 (N_5246,N_4549,N_4925);
xnor U5247 (N_5247,N_4368,N_4589);
and U5248 (N_5248,N_4989,N_4452);
nor U5249 (N_5249,N_4694,N_4887);
nand U5250 (N_5250,N_4667,N_4302);
and U5251 (N_5251,N_4937,N_4884);
and U5252 (N_5252,N_4696,N_4607);
or U5253 (N_5253,N_4551,N_4512);
or U5254 (N_5254,N_4750,N_4894);
and U5255 (N_5255,N_4850,N_4608);
or U5256 (N_5256,N_4172,N_4971);
nand U5257 (N_5257,N_4669,N_4171);
or U5258 (N_5258,N_4952,N_4414);
nor U5259 (N_5259,N_4846,N_4797);
nor U5260 (N_5260,N_4553,N_4743);
or U5261 (N_5261,N_4391,N_4289);
and U5262 (N_5262,N_4075,N_4166);
nor U5263 (N_5263,N_4251,N_4433);
and U5264 (N_5264,N_4869,N_4672);
nor U5265 (N_5265,N_4564,N_4444);
nand U5266 (N_5266,N_4654,N_4224);
or U5267 (N_5267,N_4660,N_4723);
nand U5268 (N_5268,N_4586,N_4501);
and U5269 (N_5269,N_4878,N_4819);
nand U5270 (N_5270,N_4185,N_4823);
or U5271 (N_5271,N_4534,N_4263);
nand U5272 (N_5272,N_4068,N_4934);
or U5273 (N_5273,N_4430,N_4649);
nand U5274 (N_5274,N_4542,N_4351);
or U5275 (N_5275,N_4013,N_4284);
nand U5276 (N_5276,N_4957,N_4022);
and U5277 (N_5277,N_4084,N_4505);
or U5278 (N_5278,N_4701,N_4249);
or U5279 (N_5279,N_4296,N_4036);
nand U5280 (N_5280,N_4271,N_4016);
and U5281 (N_5281,N_4243,N_4378);
nor U5282 (N_5282,N_4077,N_4795);
nand U5283 (N_5283,N_4577,N_4086);
and U5284 (N_5284,N_4828,N_4636);
or U5285 (N_5285,N_4203,N_4557);
nor U5286 (N_5286,N_4079,N_4207);
and U5287 (N_5287,N_4646,N_4927);
or U5288 (N_5288,N_4682,N_4901);
or U5289 (N_5289,N_4005,N_4291);
or U5290 (N_5290,N_4196,N_4407);
nand U5291 (N_5291,N_4232,N_4466);
nand U5292 (N_5292,N_4041,N_4057);
nor U5293 (N_5293,N_4329,N_4507);
nor U5294 (N_5294,N_4990,N_4996);
or U5295 (N_5295,N_4686,N_4426);
and U5296 (N_5296,N_4058,N_4427);
and U5297 (N_5297,N_4245,N_4511);
and U5298 (N_5298,N_4278,N_4054);
nand U5299 (N_5299,N_4107,N_4403);
and U5300 (N_5300,N_4976,N_4300);
or U5301 (N_5301,N_4353,N_4488);
and U5302 (N_5302,N_4541,N_4180);
nand U5303 (N_5303,N_4294,N_4114);
or U5304 (N_5304,N_4168,N_4810);
or U5305 (N_5305,N_4955,N_4354);
nor U5306 (N_5306,N_4328,N_4200);
nand U5307 (N_5307,N_4213,N_4606);
or U5308 (N_5308,N_4690,N_4241);
or U5309 (N_5309,N_4537,N_4169);
nor U5310 (N_5310,N_4735,N_4179);
nand U5311 (N_5311,N_4550,N_4050);
nand U5312 (N_5312,N_4276,N_4775);
nand U5313 (N_5313,N_4922,N_4215);
or U5314 (N_5314,N_4814,N_4779);
and U5315 (N_5315,N_4316,N_4162);
or U5316 (N_5316,N_4579,N_4157);
nor U5317 (N_5317,N_4155,N_4676);
nor U5318 (N_5318,N_4141,N_4872);
nand U5319 (N_5319,N_4771,N_4247);
nor U5320 (N_5320,N_4004,N_4746);
or U5321 (N_5321,N_4757,N_4642);
or U5322 (N_5322,N_4480,N_4261);
nand U5323 (N_5323,N_4926,N_4165);
and U5324 (N_5324,N_4371,N_4193);
or U5325 (N_5325,N_4119,N_4902);
nand U5326 (N_5326,N_4045,N_4715);
and U5327 (N_5327,N_4627,N_4562);
nand U5328 (N_5328,N_4458,N_4826);
nor U5329 (N_5329,N_4264,N_4691);
or U5330 (N_5330,N_4455,N_4584);
or U5331 (N_5331,N_4609,N_4675);
nor U5332 (N_5332,N_4749,N_4792);
nor U5333 (N_5333,N_4321,N_4431);
or U5334 (N_5334,N_4133,N_4034);
and U5335 (N_5335,N_4343,N_4499);
or U5336 (N_5336,N_4496,N_4409);
and U5337 (N_5337,N_4279,N_4521);
or U5338 (N_5338,N_4574,N_4876);
nand U5339 (N_5339,N_4565,N_4487);
nand U5340 (N_5340,N_4333,N_4765);
and U5341 (N_5341,N_4806,N_4135);
or U5342 (N_5342,N_4662,N_4002);
nor U5343 (N_5343,N_4670,N_4716);
nor U5344 (N_5344,N_4327,N_4886);
or U5345 (N_5345,N_4837,N_4235);
or U5346 (N_5346,N_4105,N_4485);
or U5347 (N_5347,N_4472,N_4991);
and U5348 (N_5348,N_4843,N_4453);
and U5349 (N_5349,N_4134,N_4297);
nand U5350 (N_5350,N_4698,N_4421);
or U5351 (N_5351,N_4620,N_4410);
or U5352 (N_5352,N_4618,N_4255);
or U5353 (N_5353,N_4824,N_4429);
nand U5354 (N_5354,N_4424,N_4078);
nand U5355 (N_5355,N_4965,N_4871);
nor U5356 (N_5356,N_4873,N_4799);
and U5357 (N_5357,N_4360,N_4282);
or U5358 (N_5358,N_4725,N_4903);
and U5359 (N_5359,N_4791,N_4183);
nor U5360 (N_5360,N_4898,N_4374);
and U5361 (N_5361,N_4516,N_4862);
and U5362 (N_5362,N_4330,N_4830);
or U5363 (N_5363,N_4842,N_4457);
and U5364 (N_5364,N_4307,N_4739);
nand U5365 (N_5365,N_4311,N_4572);
nor U5366 (N_5366,N_4756,N_4089);
nand U5367 (N_5367,N_4752,N_4656);
nor U5368 (N_5368,N_4490,N_4104);
nand U5369 (N_5369,N_4580,N_4143);
or U5370 (N_5370,N_4970,N_4003);
and U5371 (N_5371,N_4061,N_4645);
xnor U5372 (N_5372,N_4737,N_4638);
nand U5373 (N_5373,N_4040,N_4992);
or U5374 (N_5374,N_4020,N_4303);
nor U5375 (N_5375,N_4833,N_4605);
and U5376 (N_5376,N_4708,N_4286);
nor U5377 (N_5377,N_4882,N_4918);
nand U5378 (N_5378,N_4122,N_4301);
or U5379 (N_5379,N_4964,N_4318);
nor U5380 (N_5380,N_4644,N_4299);
nand U5381 (N_5381,N_4528,N_4212);
nand U5382 (N_5382,N_4340,N_4131);
nor U5383 (N_5383,N_4785,N_4436);
nand U5384 (N_5384,N_4230,N_4960);
or U5385 (N_5385,N_4741,N_4322);
nand U5386 (N_5386,N_4314,N_4170);
nand U5387 (N_5387,N_4640,N_4476);
or U5388 (N_5388,N_4651,N_4788);
xnor U5389 (N_5389,N_4760,N_4587);
nor U5390 (N_5390,N_4503,N_4868);
and U5391 (N_5391,N_4234,N_4137);
nor U5392 (N_5392,N_4007,N_4018);
nand U5393 (N_5393,N_4497,N_4154);
or U5394 (N_5394,N_4109,N_4081);
nor U5395 (N_5395,N_4800,N_4500);
and U5396 (N_5396,N_4653,N_4181);
nor U5397 (N_5397,N_4001,N_4038);
nand U5398 (N_5398,N_4724,N_4983);
xnor U5399 (N_5399,N_4635,N_4319);
or U5400 (N_5400,N_4658,N_4754);
nand U5401 (N_5401,N_4972,N_4680);
nor U5402 (N_5402,N_4233,N_4673);
and U5403 (N_5403,N_4827,N_4046);
nand U5404 (N_5404,N_4121,N_4153);
or U5405 (N_5405,N_4191,N_4950);
and U5406 (N_5406,N_4262,N_4367);
nand U5407 (N_5407,N_4794,N_4214);
nor U5408 (N_5408,N_4229,N_4831);
nor U5409 (N_5409,N_4684,N_4836);
and U5410 (N_5410,N_4540,N_4610);
or U5411 (N_5411,N_4447,N_4217);
nand U5412 (N_5412,N_4761,N_4870);
and U5413 (N_5413,N_4080,N_4547);
and U5414 (N_5414,N_4164,N_4755);
nor U5415 (N_5415,N_4471,N_4310);
or U5416 (N_5416,N_4777,N_4456);
nor U5417 (N_5417,N_4227,N_4290);
or U5418 (N_5418,N_4712,N_4555);
nor U5419 (N_5419,N_4769,N_4482);
and U5420 (N_5420,N_4408,N_4930);
and U5421 (N_5421,N_4896,N_4544);
or U5422 (N_5422,N_4959,N_4695);
or U5423 (N_5423,N_4082,N_4639);
nor U5424 (N_5424,N_4973,N_4177);
or U5425 (N_5425,N_4945,N_4416);
nor U5426 (N_5426,N_4049,N_4142);
and U5427 (N_5427,N_4692,N_4350);
nand U5428 (N_5428,N_4908,N_4940);
or U5429 (N_5429,N_4443,N_4559);
and U5430 (N_5430,N_4346,N_4802);
nand U5431 (N_5431,N_4438,N_4093);
xnor U5432 (N_5432,N_4388,N_4567);
nand U5433 (N_5433,N_4167,N_4689);
nand U5434 (N_5434,N_4092,N_4829);
and U5435 (N_5435,N_4461,N_4969);
or U5436 (N_5436,N_4588,N_4192);
xnor U5437 (N_5437,N_4526,N_4257);
and U5438 (N_5438,N_4032,N_4435);
nor U5439 (N_5439,N_4813,N_4341);
nand U5440 (N_5440,N_4226,N_4210);
or U5441 (N_5441,N_4678,N_4037);
nand U5442 (N_5442,N_4220,N_4626);
nand U5443 (N_5443,N_4315,N_4096);
and U5444 (N_5444,N_4890,N_4738);
nand U5445 (N_5445,N_4529,N_4031);
and U5446 (N_5446,N_4552,N_4877);
nand U5447 (N_5447,N_4380,N_4647);
or U5448 (N_5448,N_4776,N_4359);
nand U5449 (N_5449,N_4793,N_4999);
and U5450 (N_5450,N_4611,N_4719);
and U5451 (N_5451,N_4017,N_4478);
nor U5452 (N_5452,N_4356,N_4498);
and U5453 (N_5453,N_4909,N_4504);
nor U5454 (N_5454,N_4042,N_4531);
and U5455 (N_5455,N_4148,N_4851);
nand U5456 (N_5456,N_4039,N_4958);
nand U5457 (N_5457,N_4111,N_4539);
nand U5458 (N_5458,N_4917,N_4146);
and U5459 (N_5459,N_4347,N_4362);
nand U5460 (N_5460,N_4866,N_4744);
nand U5461 (N_5461,N_4522,N_4012);
or U5462 (N_5462,N_4161,N_4928);
and U5463 (N_5463,N_4710,N_4897);
and U5464 (N_5464,N_4933,N_4445);
and U5465 (N_5465,N_4706,N_4845);
nand U5466 (N_5466,N_4202,N_4615);
xnor U5467 (N_5467,N_4331,N_4197);
nand U5468 (N_5468,N_4634,N_4150);
or U5469 (N_5469,N_4532,N_4700);
and U5470 (N_5470,N_4442,N_4494);
and U5471 (N_5471,N_4633,N_4434);
or U5472 (N_5472,N_4575,N_4382);
or U5473 (N_5473,N_4617,N_4106);
nand U5474 (N_5474,N_4023,N_4736);
nor U5475 (N_5475,N_4051,N_4932);
nand U5476 (N_5476,N_4582,N_4394);
or U5477 (N_5477,N_4428,N_4239);
nor U5478 (N_5478,N_4304,N_4546);
nor U5479 (N_5479,N_4312,N_4681);
and U5480 (N_5480,N_4705,N_4253);
or U5481 (N_5481,N_4679,N_4801);
nand U5482 (N_5482,N_4189,N_4489);
nor U5483 (N_5483,N_4277,N_4768);
xnor U5484 (N_5484,N_4697,N_4101);
and U5485 (N_5485,N_4502,N_4911);
or U5486 (N_5486,N_4915,N_4363);
or U5487 (N_5487,N_4563,N_4566);
or U5488 (N_5488,N_4839,N_4293);
and U5489 (N_5489,N_4748,N_4248);
nor U5490 (N_5490,N_4596,N_4717);
and U5491 (N_5491,N_4840,N_4128);
or U5492 (N_5492,N_4923,N_4535);
and U5493 (N_5493,N_4218,N_4140);
and U5494 (N_5494,N_4342,N_4053);
or U5495 (N_5495,N_4883,N_4581);
or U5496 (N_5496,N_4120,N_4943);
nand U5497 (N_5497,N_4309,N_4187);
nand U5498 (N_5498,N_4381,N_4352);
nor U5499 (N_5499,N_4097,N_4912);
or U5500 (N_5500,N_4498,N_4159);
or U5501 (N_5501,N_4603,N_4634);
xor U5502 (N_5502,N_4503,N_4246);
nand U5503 (N_5503,N_4694,N_4400);
nor U5504 (N_5504,N_4517,N_4003);
nor U5505 (N_5505,N_4015,N_4187);
or U5506 (N_5506,N_4433,N_4976);
or U5507 (N_5507,N_4445,N_4179);
nor U5508 (N_5508,N_4248,N_4909);
and U5509 (N_5509,N_4215,N_4053);
xor U5510 (N_5510,N_4197,N_4940);
nor U5511 (N_5511,N_4031,N_4647);
and U5512 (N_5512,N_4594,N_4157);
nor U5513 (N_5513,N_4443,N_4037);
or U5514 (N_5514,N_4044,N_4315);
nor U5515 (N_5515,N_4113,N_4025);
and U5516 (N_5516,N_4889,N_4879);
and U5517 (N_5517,N_4433,N_4113);
or U5518 (N_5518,N_4825,N_4914);
nor U5519 (N_5519,N_4793,N_4534);
and U5520 (N_5520,N_4452,N_4328);
or U5521 (N_5521,N_4922,N_4266);
and U5522 (N_5522,N_4158,N_4325);
and U5523 (N_5523,N_4405,N_4820);
nor U5524 (N_5524,N_4072,N_4597);
nand U5525 (N_5525,N_4969,N_4884);
or U5526 (N_5526,N_4938,N_4011);
and U5527 (N_5527,N_4961,N_4736);
or U5528 (N_5528,N_4986,N_4925);
and U5529 (N_5529,N_4225,N_4148);
nor U5530 (N_5530,N_4470,N_4428);
or U5531 (N_5531,N_4568,N_4034);
and U5532 (N_5532,N_4700,N_4585);
or U5533 (N_5533,N_4072,N_4162);
and U5534 (N_5534,N_4107,N_4427);
or U5535 (N_5535,N_4283,N_4791);
and U5536 (N_5536,N_4828,N_4434);
or U5537 (N_5537,N_4540,N_4565);
or U5538 (N_5538,N_4153,N_4358);
and U5539 (N_5539,N_4651,N_4144);
and U5540 (N_5540,N_4230,N_4912);
and U5541 (N_5541,N_4510,N_4223);
and U5542 (N_5542,N_4214,N_4451);
and U5543 (N_5543,N_4999,N_4557);
and U5544 (N_5544,N_4733,N_4118);
xor U5545 (N_5545,N_4605,N_4546);
or U5546 (N_5546,N_4568,N_4438);
nor U5547 (N_5547,N_4035,N_4471);
and U5548 (N_5548,N_4437,N_4538);
nor U5549 (N_5549,N_4578,N_4573);
nor U5550 (N_5550,N_4686,N_4728);
nand U5551 (N_5551,N_4219,N_4250);
nor U5552 (N_5552,N_4003,N_4734);
nor U5553 (N_5553,N_4842,N_4325);
nor U5554 (N_5554,N_4998,N_4099);
xnor U5555 (N_5555,N_4506,N_4585);
and U5556 (N_5556,N_4120,N_4359);
and U5557 (N_5557,N_4432,N_4276);
nor U5558 (N_5558,N_4879,N_4521);
nand U5559 (N_5559,N_4791,N_4641);
and U5560 (N_5560,N_4556,N_4721);
nor U5561 (N_5561,N_4963,N_4424);
or U5562 (N_5562,N_4413,N_4900);
nor U5563 (N_5563,N_4727,N_4429);
or U5564 (N_5564,N_4928,N_4955);
and U5565 (N_5565,N_4139,N_4855);
or U5566 (N_5566,N_4936,N_4959);
nor U5567 (N_5567,N_4268,N_4658);
nor U5568 (N_5568,N_4921,N_4313);
and U5569 (N_5569,N_4687,N_4947);
or U5570 (N_5570,N_4747,N_4889);
nand U5571 (N_5571,N_4665,N_4072);
and U5572 (N_5572,N_4002,N_4100);
nand U5573 (N_5573,N_4372,N_4270);
or U5574 (N_5574,N_4098,N_4353);
nor U5575 (N_5575,N_4653,N_4871);
or U5576 (N_5576,N_4948,N_4421);
nand U5577 (N_5577,N_4707,N_4820);
nand U5578 (N_5578,N_4664,N_4749);
and U5579 (N_5579,N_4245,N_4614);
and U5580 (N_5580,N_4428,N_4533);
nand U5581 (N_5581,N_4155,N_4737);
or U5582 (N_5582,N_4351,N_4023);
nor U5583 (N_5583,N_4172,N_4788);
nand U5584 (N_5584,N_4102,N_4373);
nand U5585 (N_5585,N_4338,N_4723);
or U5586 (N_5586,N_4544,N_4204);
or U5587 (N_5587,N_4361,N_4754);
nor U5588 (N_5588,N_4266,N_4217);
or U5589 (N_5589,N_4682,N_4783);
nand U5590 (N_5590,N_4282,N_4213);
nor U5591 (N_5591,N_4923,N_4470);
and U5592 (N_5592,N_4555,N_4287);
or U5593 (N_5593,N_4687,N_4568);
or U5594 (N_5594,N_4683,N_4346);
nand U5595 (N_5595,N_4216,N_4458);
xnor U5596 (N_5596,N_4551,N_4418);
and U5597 (N_5597,N_4541,N_4150);
nand U5598 (N_5598,N_4096,N_4612);
nand U5599 (N_5599,N_4238,N_4695);
nor U5600 (N_5600,N_4634,N_4775);
and U5601 (N_5601,N_4511,N_4175);
nor U5602 (N_5602,N_4865,N_4123);
and U5603 (N_5603,N_4269,N_4078);
nand U5604 (N_5604,N_4289,N_4636);
nand U5605 (N_5605,N_4527,N_4023);
and U5606 (N_5606,N_4108,N_4176);
nand U5607 (N_5607,N_4688,N_4601);
and U5608 (N_5608,N_4161,N_4254);
nand U5609 (N_5609,N_4175,N_4382);
nor U5610 (N_5610,N_4764,N_4466);
nand U5611 (N_5611,N_4380,N_4290);
or U5612 (N_5612,N_4907,N_4077);
or U5613 (N_5613,N_4968,N_4144);
nand U5614 (N_5614,N_4172,N_4026);
or U5615 (N_5615,N_4645,N_4012);
and U5616 (N_5616,N_4450,N_4328);
xnor U5617 (N_5617,N_4166,N_4779);
or U5618 (N_5618,N_4829,N_4517);
xor U5619 (N_5619,N_4011,N_4773);
and U5620 (N_5620,N_4329,N_4805);
nor U5621 (N_5621,N_4554,N_4670);
nor U5622 (N_5622,N_4164,N_4636);
and U5623 (N_5623,N_4471,N_4615);
and U5624 (N_5624,N_4373,N_4696);
nor U5625 (N_5625,N_4697,N_4292);
and U5626 (N_5626,N_4052,N_4921);
and U5627 (N_5627,N_4525,N_4067);
and U5628 (N_5628,N_4692,N_4954);
nand U5629 (N_5629,N_4390,N_4090);
or U5630 (N_5630,N_4648,N_4175);
and U5631 (N_5631,N_4699,N_4845);
and U5632 (N_5632,N_4814,N_4749);
nor U5633 (N_5633,N_4307,N_4959);
nor U5634 (N_5634,N_4415,N_4163);
nor U5635 (N_5635,N_4596,N_4834);
or U5636 (N_5636,N_4883,N_4035);
xnor U5637 (N_5637,N_4873,N_4896);
or U5638 (N_5638,N_4393,N_4628);
nor U5639 (N_5639,N_4988,N_4022);
nor U5640 (N_5640,N_4782,N_4884);
or U5641 (N_5641,N_4082,N_4449);
nor U5642 (N_5642,N_4000,N_4012);
and U5643 (N_5643,N_4337,N_4868);
nor U5644 (N_5644,N_4639,N_4409);
or U5645 (N_5645,N_4088,N_4261);
nand U5646 (N_5646,N_4373,N_4610);
or U5647 (N_5647,N_4217,N_4602);
nor U5648 (N_5648,N_4546,N_4329);
nand U5649 (N_5649,N_4677,N_4767);
and U5650 (N_5650,N_4559,N_4040);
or U5651 (N_5651,N_4231,N_4271);
and U5652 (N_5652,N_4901,N_4681);
and U5653 (N_5653,N_4505,N_4441);
and U5654 (N_5654,N_4129,N_4396);
nand U5655 (N_5655,N_4451,N_4572);
nor U5656 (N_5656,N_4837,N_4532);
and U5657 (N_5657,N_4069,N_4930);
or U5658 (N_5658,N_4854,N_4629);
or U5659 (N_5659,N_4743,N_4646);
nor U5660 (N_5660,N_4917,N_4038);
or U5661 (N_5661,N_4401,N_4799);
and U5662 (N_5662,N_4978,N_4535);
nor U5663 (N_5663,N_4528,N_4844);
nor U5664 (N_5664,N_4925,N_4387);
nand U5665 (N_5665,N_4870,N_4612);
and U5666 (N_5666,N_4840,N_4467);
nor U5667 (N_5667,N_4773,N_4742);
nor U5668 (N_5668,N_4045,N_4031);
nor U5669 (N_5669,N_4776,N_4452);
and U5670 (N_5670,N_4035,N_4876);
and U5671 (N_5671,N_4668,N_4449);
nor U5672 (N_5672,N_4587,N_4917);
nor U5673 (N_5673,N_4490,N_4940);
nand U5674 (N_5674,N_4233,N_4632);
or U5675 (N_5675,N_4002,N_4311);
nor U5676 (N_5676,N_4855,N_4530);
and U5677 (N_5677,N_4974,N_4342);
and U5678 (N_5678,N_4567,N_4551);
nand U5679 (N_5679,N_4334,N_4682);
or U5680 (N_5680,N_4187,N_4522);
or U5681 (N_5681,N_4134,N_4856);
nor U5682 (N_5682,N_4335,N_4522);
nand U5683 (N_5683,N_4494,N_4041);
or U5684 (N_5684,N_4584,N_4283);
and U5685 (N_5685,N_4601,N_4528);
or U5686 (N_5686,N_4537,N_4038);
nand U5687 (N_5687,N_4216,N_4220);
xor U5688 (N_5688,N_4320,N_4414);
xor U5689 (N_5689,N_4652,N_4628);
or U5690 (N_5690,N_4608,N_4282);
or U5691 (N_5691,N_4728,N_4743);
xnor U5692 (N_5692,N_4393,N_4678);
nor U5693 (N_5693,N_4556,N_4608);
and U5694 (N_5694,N_4056,N_4442);
nor U5695 (N_5695,N_4218,N_4437);
or U5696 (N_5696,N_4477,N_4991);
nor U5697 (N_5697,N_4632,N_4391);
and U5698 (N_5698,N_4236,N_4860);
and U5699 (N_5699,N_4536,N_4907);
nor U5700 (N_5700,N_4712,N_4051);
nor U5701 (N_5701,N_4377,N_4865);
and U5702 (N_5702,N_4859,N_4011);
nand U5703 (N_5703,N_4067,N_4029);
and U5704 (N_5704,N_4370,N_4650);
and U5705 (N_5705,N_4573,N_4292);
or U5706 (N_5706,N_4678,N_4961);
or U5707 (N_5707,N_4528,N_4862);
nand U5708 (N_5708,N_4544,N_4426);
nand U5709 (N_5709,N_4700,N_4993);
or U5710 (N_5710,N_4832,N_4376);
and U5711 (N_5711,N_4782,N_4881);
and U5712 (N_5712,N_4445,N_4125);
and U5713 (N_5713,N_4805,N_4350);
nor U5714 (N_5714,N_4713,N_4482);
nand U5715 (N_5715,N_4304,N_4623);
nand U5716 (N_5716,N_4420,N_4689);
nand U5717 (N_5717,N_4521,N_4462);
and U5718 (N_5718,N_4289,N_4320);
nand U5719 (N_5719,N_4795,N_4238);
nand U5720 (N_5720,N_4098,N_4810);
nand U5721 (N_5721,N_4038,N_4766);
or U5722 (N_5722,N_4810,N_4620);
nand U5723 (N_5723,N_4874,N_4248);
or U5724 (N_5724,N_4557,N_4130);
or U5725 (N_5725,N_4025,N_4715);
or U5726 (N_5726,N_4812,N_4778);
nor U5727 (N_5727,N_4813,N_4597);
nand U5728 (N_5728,N_4727,N_4135);
or U5729 (N_5729,N_4641,N_4760);
nand U5730 (N_5730,N_4139,N_4107);
and U5731 (N_5731,N_4294,N_4559);
nor U5732 (N_5732,N_4865,N_4011);
or U5733 (N_5733,N_4784,N_4475);
nand U5734 (N_5734,N_4484,N_4754);
nor U5735 (N_5735,N_4069,N_4961);
nor U5736 (N_5736,N_4134,N_4032);
nor U5737 (N_5737,N_4200,N_4446);
nor U5738 (N_5738,N_4278,N_4829);
and U5739 (N_5739,N_4654,N_4470);
xnor U5740 (N_5740,N_4517,N_4669);
nor U5741 (N_5741,N_4462,N_4467);
and U5742 (N_5742,N_4035,N_4283);
and U5743 (N_5743,N_4929,N_4585);
nand U5744 (N_5744,N_4341,N_4798);
and U5745 (N_5745,N_4270,N_4106);
or U5746 (N_5746,N_4298,N_4613);
nor U5747 (N_5747,N_4055,N_4921);
xnor U5748 (N_5748,N_4922,N_4439);
xor U5749 (N_5749,N_4944,N_4168);
nor U5750 (N_5750,N_4232,N_4182);
nand U5751 (N_5751,N_4383,N_4414);
nor U5752 (N_5752,N_4239,N_4219);
or U5753 (N_5753,N_4377,N_4640);
or U5754 (N_5754,N_4125,N_4428);
and U5755 (N_5755,N_4570,N_4396);
nand U5756 (N_5756,N_4984,N_4319);
and U5757 (N_5757,N_4059,N_4128);
and U5758 (N_5758,N_4590,N_4860);
and U5759 (N_5759,N_4916,N_4343);
or U5760 (N_5760,N_4505,N_4117);
nor U5761 (N_5761,N_4499,N_4134);
or U5762 (N_5762,N_4176,N_4968);
or U5763 (N_5763,N_4636,N_4980);
and U5764 (N_5764,N_4626,N_4355);
nand U5765 (N_5765,N_4630,N_4500);
nor U5766 (N_5766,N_4102,N_4306);
and U5767 (N_5767,N_4395,N_4890);
nor U5768 (N_5768,N_4114,N_4160);
or U5769 (N_5769,N_4178,N_4787);
and U5770 (N_5770,N_4122,N_4813);
and U5771 (N_5771,N_4372,N_4519);
nor U5772 (N_5772,N_4997,N_4076);
nor U5773 (N_5773,N_4123,N_4817);
nor U5774 (N_5774,N_4843,N_4919);
and U5775 (N_5775,N_4616,N_4093);
nor U5776 (N_5776,N_4617,N_4328);
or U5777 (N_5777,N_4406,N_4080);
and U5778 (N_5778,N_4860,N_4152);
nor U5779 (N_5779,N_4399,N_4673);
nor U5780 (N_5780,N_4203,N_4062);
nor U5781 (N_5781,N_4332,N_4853);
or U5782 (N_5782,N_4628,N_4523);
nand U5783 (N_5783,N_4863,N_4697);
or U5784 (N_5784,N_4967,N_4999);
or U5785 (N_5785,N_4050,N_4016);
nor U5786 (N_5786,N_4893,N_4947);
or U5787 (N_5787,N_4566,N_4733);
or U5788 (N_5788,N_4986,N_4466);
nor U5789 (N_5789,N_4550,N_4506);
or U5790 (N_5790,N_4504,N_4766);
or U5791 (N_5791,N_4811,N_4756);
and U5792 (N_5792,N_4132,N_4486);
or U5793 (N_5793,N_4215,N_4577);
or U5794 (N_5794,N_4683,N_4819);
nand U5795 (N_5795,N_4353,N_4432);
or U5796 (N_5796,N_4801,N_4876);
nor U5797 (N_5797,N_4321,N_4868);
nor U5798 (N_5798,N_4678,N_4895);
and U5799 (N_5799,N_4637,N_4098);
and U5800 (N_5800,N_4043,N_4494);
nor U5801 (N_5801,N_4693,N_4727);
nand U5802 (N_5802,N_4022,N_4417);
or U5803 (N_5803,N_4746,N_4043);
or U5804 (N_5804,N_4807,N_4625);
or U5805 (N_5805,N_4228,N_4794);
or U5806 (N_5806,N_4083,N_4474);
or U5807 (N_5807,N_4371,N_4155);
nor U5808 (N_5808,N_4989,N_4117);
and U5809 (N_5809,N_4119,N_4245);
or U5810 (N_5810,N_4878,N_4921);
and U5811 (N_5811,N_4229,N_4767);
nand U5812 (N_5812,N_4898,N_4446);
nor U5813 (N_5813,N_4922,N_4320);
and U5814 (N_5814,N_4894,N_4769);
and U5815 (N_5815,N_4798,N_4827);
or U5816 (N_5816,N_4799,N_4669);
nand U5817 (N_5817,N_4540,N_4852);
or U5818 (N_5818,N_4508,N_4434);
nand U5819 (N_5819,N_4368,N_4955);
and U5820 (N_5820,N_4492,N_4016);
nand U5821 (N_5821,N_4911,N_4699);
nor U5822 (N_5822,N_4873,N_4489);
or U5823 (N_5823,N_4658,N_4069);
and U5824 (N_5824,N_4777,N_4341);
nand U5825 (N_5825,N_4688,N_4981);
or U5826 (N_5826,N_4213,N_4752);
and U5827 (N_5827,N_4130,N_4874);
or U5828 (N_5828,N_4583,N_4999);
nand U5829 (N_5829,N_4637,N_4244);
and U5830 (N_5830,N_4858,N_4857);
nor U5831 (N_5831,N_4218,N_4248);
nor U5832 (N_5832,N_4008,N_4533);
or U5833 (N_5833,N_4874,N_4950);
or U5834 (N_5834,N_4526,N_4020);
or U5835 (N_5835,N_4590,N_4080);
nor U5836 (N_5836,N_4235,N_4377);
and U5837 (N_5837,N_4422,N_4505);
nor U5838 (N_5838,N_4966,N_4912);
or U5839 (N_5839,N_4143,N_4387);
nor U5840 (N_5840,N_4735,N_4877);
and U5841 (N_5841,N_4954,N_4947);
nand U5842 (N_5842,N_4443,N_4645);
and U5843 (N_5843,N_4216,N_4034);
nor U5844 (N_5844,N_4135,N_4570);
nand U5845 (N_5845,N_4858,N_4388);
or U5846 (N_5846,N_4615,N_4791);
nor U5847 (N_5847,N_4856,N_4043);
nor U5848 (N_5848,N_4922,N_4788);
nor U5849 (N_5849,N_4620,N_4668);
and U5850 (N_5850,N_4530,N_4175);
nor U5851 (N_5851,N_4845,N_4884);
or U5852 (N_5852,N_4453,N_4245);
nor U5853 (N_5853,N_4703,N_4638);
nor U5854 (N_5854,N_4221,N_4157);
or U5855 (N_5855,N_4226,N_4660);
or U5856 (N_5856,N_4207,N_4269);
nand U5857 (N_5857,N_4077,N_4123);
xnor U5858 (N_5858,N_4245,N_4464);
xor U5859 (N_5859,N_4183,N_4210);
xnor U5860 (N_5860,N_4833,N_4157);
nand U5861 (N_5861,N_4421,N_4614);
and U5862 (N_5862,N_4218,N_4885);
or U5863 (N_5863,N_4949,N_4955);
nor U5864 (N_5864,N_4999,N_4691);
and U5865 (N_5865,N_4436,N_4864);
nand U5866 (N_5866,N_4853,N_4367);
nand U5867 (N_5867,N_4414,N_4944);
and U5868 (N_5868,N_4557,N_4147);
nor U5869 (N_5869,N_4952,N_4428);
nor U5870 (N_5870,N_4867,N_4794);
nand U5871 (N_5871,N_4662,N_4838);
nand U5872 (N_5872,N_4298,N_4108);
or U5873 (N_5873,N_4040,N_4317);
nor U5874 (N_5874,N_4576,N_4614);
nor U5875 (N_5875,N_4575,N_4105);
nor U5876 (N_5876,N_4230,N_4721);
or U5877 (N_5877,N_4524,N_4987);
and U5878 (N_5878,N_4819,N_4524);
and U5879 (N_5879,N_4732,N_4658);
and U5880 (N_5880,N_4257,N_4480);
or U5881 (N_5881,N_4068,N_4119);
or U5882 (N_5882,N_4046,N_4248);
and U5883 (N_5883,N_4616,N_4243);
and U5884 (N_5884,N_4329,N_4263);
or U5885 (N_5885,N_4097,N_4388);
nand U5886 (N_5886,N_4446,N_4308);
nand U5887 (N_5887,N_4124,N_4416);
nand U5888 (N_5888,N_4088,N_4276);
nor U5889 (N_5889,N_4627,N_4303);
and U5890 (N_5890,N_4250,N_4906);
nand U5891 (N_5891,N_4853,N_4874);
or U5892 (N_5892,N_4628,N_4363);
and U5893 (N_5893,N_4335,N_4795);
or U5894 (N_5894,N_4802,N_4176);
nor U5895 (N_5895,N_4279,N_4857);
and U5896 (N_5896,N_4156,N_4783);
nand U5897 (N_5897,N_4967,N_4213);
nor U5898 (N_5898,N_4120,N_4729);
and U5899 (N_5899,N_4569,N_4936);
and U5900 (N_5900,N_4363,N_4439);
and U5901 (N_5901,N_4762,N_4203);
nor U5902 (N_5902,N_4525,N_4566);
nor U5903 (N_5903,N_4424,N_4088);
xnor U5904 (N_5904,N_4541,N_4046);
and U5905 (N_5905,N_4563,N_4083);
and U5906 (N_5906,N_4326,N_4104);
nor U5907 (N_5907,N_4167,N_4439);
and U5908 (N_5908,N_4547,N_4577);
nand U5909 (N_5909,N_4993,N_4622);
nor U5910 (N_5910,N_4505,N_4172);
nand U5911 (N_5911,N_4940,N_4977);
nand U5912 (N_5912,N_4941,N_4679);
and U5913 (N_5913,N_4209,N_4294);
or U5914 (N_5914,N_4619,N_4035);
nand U5915 (N_5915,N_4210,N_4859);
and U5916 (N_5916,N_4147,N_4958);
nor U5917 (N_5917,N_4305,N_4053);
and U5918 (N_5918,N_4078,N_4468);
and U5919 (N_5919,N_4322,N_4318);
nand U5920 (N_5920,N_4116,N_4939);
or U5921 (N_5921,N_4022,N_4461);
and U5922 (N_5922,N_4860,N_4782);
nor U5923 (N_5923,N_4576,N_4167);
nor U5924 (N_5924,N_4040,N_4329);
or U5925 (N_5925,N_4819,N_4456);
nand U5926 (N_5926,N_4706,N_4200);
xor U5927 (N_5927,N_4118,N_4261);
or U5928 (N_5928,N_4053,N_4183);
nand U5929 (N_5929,N_4084,N_4216);
and U5930 (N_5930,N_4910,N_4117);
nor U5931 (N_5931,N_4566,N_4797);
and U5932 (N_5932,N_4216,N_4338);
nand U5933 (N_5933,N_4304,N_4282);
and U5934 (N_5934,N_4601,N_4391);
and U5935 (N_5935,N_4384,N_4225);
nor U5936 (N_5936,N_4915,N_4357);
nand U5937 (N_5937,N_4838,N_4698);
xor U5938 (N_5938,N_4661,N_4165);
and U5939 (N_5939,N_4316,N_4273);
nor U5940 (N_5940,N_4799,N_4853);
and U5941 (N_5941,N_4619,N_4050);
nand U5942 (N_5942,N_4227,N_4094);
or U5943 (N_5943,N_4669,N_4140);
nand U5944 (N_5944,N_4780,N_4612);
and U5945 (N_5945,N_4702,N_4707);
xnor U5946 (N_5946,N_4612,N_4664);
nor U5947 (N_5947,N_4605,N_4692);
nand U5948 (N_5948,N_4311,N_4735);
and U5949 (N_5949,N_4942,N_4281);
and U5950 (N_5950,N_4594,N_4407);
or U5951 (N_5951,N_4238,N_4506);
and U5952 (N_5952,N_4258,N_4677);
and U5953 (N_5953,N_4192,N_4808);
and U5954 (N_5954,N_4575,N_4322);
nand U5955 (N_5955,N_4558,N_4742);
nand U5956 (N_5956,N_4699,N_4338);
nor U5957 (N_5957,N_4317,N_4986);
nand U5958 (N_5958,N_4500,N_4072);
nor U5959 (N_5959,N_4351,N_4585);
or U5960 (N_5960,N_4432,N_4070);
and U5961 (N_5961,N_4067,N_4824);
and U5962 (N_5962,N_4524,N_4018);
nor U5963 (N_5963,N_4073,N_4383);
and U5964 (N_5964,N_4019,N_4517);
nand U5965 (N_5965,N_4229,N_4373);
or U5966 (N_5966,N_4995,N_4044);
nor U5967 (N_5967,N_4665,N_4389);
nor U5968 (N_5968,N_4676,N_4478);
nand U5969 (N_5969,N_4581,N_4512);
xor U5970 (N_5970,N_4813,N_4018);
or U5971 (N_5971,N_4010,N_4457);
and U5972 (N_5972,N_4202,N_4606);
nor U5973 (N_5973,N_4973,N_4260);
and U5974 (N_5974,N_4280,N_4245);
and U5975 (N_5975,N_4310,N_4828);
xnor U5976 (N_5976,N_4557,N_4264);
or U5977 (N_5977,N_4599,N_4504);
nand U5978 (N_5978,N_4968,N_4876);
or U5979 (N_5979,N_4616,N_4771);
and U5980 (N_5980,N_4355,N_4124);
nor U5981 (N_5981,N_4038,N_4210);
nand U5982 (N_5982,N_4885,N_4486);
and U5983 (N_5983,N_4915,N_4632);
or U5984 (N_5984,N_4306,N_4428);
nor U5985 (N_5985,N_4619,N_4029);
nand U5986 (N_5986,N_4929,N_4265);
and U5987 (N_5987,N_4808,N_4649);
and U5988 (N_5988,N_4223,N_4449);
or U5989 (N_5989,N_4062,N_4467);
nand U5990 (N_5990,N_4416,N_4914);
nand U5991 (N_5991,N_4125,N_4704);
and U5992 (N_5992,N_4581,N_4922);
nand U5993 (N_5993,N_4673,N_4900);
or U5994 (N_5994,N_4204,N_4446);
xor U5995 (N_5995,N_4813,N_4164);
nand U5996 (N_5996,N_4789,N_4436);
and U5997 (N_5997,N_4371,N_4659);
nor U5998 (N_5998,N_4063,N_4927);
or U5999 (N_5999,N_4063,N_4809);
or U6000 (N_6000,N_5150,N_5435);
nand U6001 (N_6001,N_5142,N_5730);
or U6002 (N_6002,N_5058,N_5503);
or U6003 (N_6003,N_5995,N_5452);
or U6004 (N_6004,N_5663,N_5595);
nand U6005 (N_6005,N_5866,N_5565);
or U6006 (N_6006,N_5741,N_5299);
nor U6007 (N_6007,N_5370,N_5852);
or U6008 (N_6008,N_5260,N_5722);
or U6009 (N_6009,N_5786,N_5317);
and U6010 (N_6010,N_5512,N_5707);
nor U6011 (N_6011,N_5526,N_5388);
nor U6012 (N_6012,N_5720,N_5048);
or U6013 (N_6013,N_5180,N_5661);
nand U6014 (N_6014,N_5839,N_5132);
nand U6015 (N_6015,N_5110,N_5236);
nor U6016 (N_6016,N_5891,N_5557);
or U6017 (N_6017,N_5901,N_5264);
or U6018 (N_6018,N_5220,N_5499);
nor U6019 (N_6019,N_5815,N_5134);
and U6020 (N_6020,N_5588,N_5097);
or U6021 (N_6021,N_5768,N_5149);
and U6022 (N_6022,N_5255,N_5762);
and U6023 (N_6023,N_5480,N_5884);
and U6024 (N_6024,N_5396,N_5166);
nand U6025 (N_6025,N_5961,N_5310);
nand U6026 (N_6026,N_5051,N_5298);
nand U6027 (N_6027,N_5693,N_5071);
nor U6028 (N_6028,N_5656,N_5322);
or U6029 (N_6029,N_5613,N_5848);
and U6030 (N_6030,N_5361,N_5307);
or U6031 (N_6031,N_5266,N_5683);
and U6032 (N_6032,N_5511,N_5675);
nand U6033 (N_6033,N_5849,N_5198);
nand U6034 (N_6034,N_5125,N_5811);
nor U6035 (N_6035,N_5484,N_5842);
nand U6036 (N_6036,N_5203,N_5380);
and U6037 (N_6037,N_5709,N_5278);
nand U6038 (N_6038,N_5053,N_5382);
or U6039 (N_6039,N_5128,N_5805);
and U6040 (N_6040,N_5070,N_5778);
nand U6041 (N_6041,N_5272,N_5056);
and U6042 (N_6042,N_5518,N_5776);
or U6043 (N_6043,N_5340,N_5457);
or U6044 (N_6044,N_5104,N_5543);
or U6045 (N_6045,N_5772,N_5444);
nor U6046 (N_6046,N_5823,N_5785);
and U6047 (N_6047,N_5812,N_5034);
or U6048 (N_6048,N_5344,N_5471);
and U6049 (N_6049,N_5250,N_5515);
nand U6050 (N_6050,N_5075,N_5280);
and U6051 (N_6051,N_5064,N_5157);
and U6052 (N_6052,N_5969,N_5599);
nor U6053 (N_6053,N_5603,N_5323);
and U6054 (N_6054,N_5978,N_5558);
nand U6055 (N_6055,N_5637,N_5294);
or U6056 (N_6056,N_5485,N_5477);
and U6057 (N_6057,N_5464,N_5951);
nor U6058 (N_6058,N_5694,N_5226);
and U6059 (N_6059,N_5688,N_5508);
or U6060 (N_6060,N_5659,N_5871);
nand U6061 (N_6061,N_5817,N_5907);
nor U6062 (N_6062,N_5872,N_5647);
xnor U6063 (N_6063,N_5315,N_5006);
nand U6064 (N_6064,N_5689,N_5769);
or U6065 (N_6065,N_5943,N_5268);
and U6066 (N_6066,N_5212,N_5389);
or U6067 (N_6067,N_5617,N_5883);
nand U6068 (N_6068,N_5224,N_5256);
or U6069 (N_6069,N_5274,N_5265);
or U6070 (N_6070,N_5208,N_5218);
and U6071 (N_6071,N_5790,N_5390);
and U6072 (N_6072,N_5551,N_5939);
or U6073 (N_6073,N_5810,N_5442);
and U6074 (N_6074,N_5835,N_5467);
and U6075 (N_6075,N_5509,N_5343);
or U6076 (N_6076,N_5592,N_5845);
or U6077 (N_6077,N_5314,N_5788);
and U6078 (N_6078,N_5779,N_5590);
or U6079 (N_6079,N_5487,N_5710);
or U6080 (N_6080,N_5522,N_5743);
nand U6081 (N_6081,N_5666,N_5279);
nor U6082 (N_6082,N_5600,N_5738);
nor U6083 (N_6083,N_5712,N_5705);
nor U6084 (N_6084,N_5018,N_5654);
or U6085 (N_6085,N_5628,N_5148);
and U6086 (N_6086,N_5465,N_5041);
and U6087 (N_6087,N_5809,N_5765);
or U6088 (N_6088,N_5251,N_5195);
nor U6089 (N_6089,N_5427,N_5039);
nand U6090 (N_6090,N_5245,N_5986);
nand U6091 (N_6091,N_5934,N_5228);
nand U6092 (N_6092,N_5665,N_5035);
and U6093 (N_6093,N_5874,N_5231);
or U6094 (N_6094,N_5106,N_5135);
nor U6095 (N_6095,N_5119,N_5297);
nor U6096 (N_6096,N_5283,N_5843);
nor U6097 (N_6097,N_5957,N_5481);
or U6098 (N_6098,N_5140,N_5353);
nand U6099 (N_6099,N_5129,N_5649);
nor U6100 (N_6100,N_5660,N_5933);
and U6101 (N_6101,N_5523,N_5942);
and U6102 (N_6102,N_5821,N_5702);
and U6103 (N_6103,N_5998,N_5253);
nand U6104 (N_6104,N_5020,N_5413);
or U6105 (N_6105,N_5893,N_5873);
or U6106 (N_6106,N_5882,N_5763);
or U6107 (N_6107,N_5830,N_5540);
nor U6108 (N_6108,N_5581,N_5093);
nand U6109 (N_6109,N_5729,N_5336);
nor U6110 (N_6110,N_5202,N_5291);
nand U6111 (N_6111,N_5910,N_5597);
and U6112 (N_6112,N_5136,N_5755);
nor U6113 (N_6113,N_5716,N_5420);
and U6114 (N_6114,N_5573,N_5248);
nor U6115 (N_6115,N_5807,N_5384);
or U6116 (N_6116,N_5171,N_5703);
nor U6117 (N_6117,N_5400,N_5520);
and U6118 (N_6118,N_5112,N_5841);
xor U6119 (N_6119,N_5327,N_5434);
nand U6120 (N_6120,N_5914,N_5774);
nand U6121 (N_6121,N_5197,N_5909);
nand U6122 (N_6122,N_5867,N_5346);
nor U6123 (N_6123,N_5332,N_5455);
or U6124 (N_6124,N_5967,N_5182);
nand U6125 (N_6125,N_5429,N_5887);
or U6126 (N_6126,N_5886,N_5822);
or U6127 (N_6127,N_5145,N_5975);
or U6128 (N_6128,N_5046,N_5553);
nand U6129 (N_6129,N_5662,N_5284);
xor U6130 (N_6130,N_5672,N_5486);
nand U6131 (N_6131,N_5479,N_5431);
or U6132 (N_6132,N_5108,N_5160);
or U6133 (N_6133,N_5804,N_5366);
and U6134 (N_6134,N_5837,N_5917);
nor U6135 (N_6135,N_5582,N_5989);
nor U6136 (N_6136,N_5927,N_5773);
and U6137 (N_6137,N_5950,N_5879);
xor U6138 (N_6138,N_5211,N_5184);
nor U6139 (N_6139,N_5958,N_5838);
or U6140 (N_6140,N_5397,N_5889);
or U6141 (N_6141,N_5448,N_5881);
nand U6142 (N_6142,N_5156,N_5584);
nor U6143 (N_6143,N_5632,N_5983);
nand U6144 (N_6144,N_5271,N_5941);
or U6145 (N_6145,N_5766,N_5153);
or U6146 (N_6146,N_5623,N_5407);
and U6147 (N_6147,N_5191,N_5924);
nor U6148 (N_6148,N_5754,N_5609);
nand U6149 (N_6149,N_5894,N_5850);
nand U6150 (N_6150,N_5510,N_5036);
and U6151 (N_6151,N_5239,N_5799);
and U6152 (N_6152,N_5144,N_5364);
nor U6153 (N_6153,N_5542,N_5193);
and U6154 (N_6154,N_5579,N_5865);
xnor U6155 (N_6155,N_5190,N_5918);
nor U6156 (N_6156,N_5054,N_5759);
nor U6157 (N_6157,N_5357,N_5519);
nor U6158 (N_6158,N_5531,N_5834);
and U6159 (N_6159,N_5621,N_5101);
or U6160 (N_6160,N_5263,N_5399);
or U6161 (N_6161,N_5725,N_5025);
nor U6162 (N_6162,N_5751,N_5932);
nor U6163 (N_6163,N_5099,N_5846);
nand U6164 (N_6164,N_5922,N_5602);
nor U6165 (N_6165,N_5610,N_5066);
or U6166 (N_6166,N_5708,N_5063);
nand U6167 (N_6167,N_5005,N_5091);
nor U6168 (N_6168,N_5947,N_5270);
nand U6169 (N_6169,N_5437,N_5468);
nor U6170 (N_6170,N_5616,N_5719);
nand U6171 (N_6171,N_5973,N_5421);
or U6172 (N_6172,N_5282,N_5877);
xnor U6173 (N_6173,N_5223,N_5742);
nor U6174 (N_6174,N_5959,N_5147);
and U6175 (N_6175,N_5072,N_5217);
nor U6176 (N_6176,N_5293,N_5111);
or U6177 (N_6177,N_5169,N_5836);
nor U6178 (N_6178,N_5229,N_5764);
nand U6179 (N_6179,N_5533,N_5622);
nand U6180 (N_6180,N_5318,N_5612);
and U6181 (N_6181,N_5876,N_5492);
nor U6182 (N_6182,N_5858,N_5015);
nand U6183 (N_6183,N_5037,N_5436);
or U6184 (N_6184,N_5699,N_5210);
and U6185 (N_6185,N_5189,N_5962);
nor U6186 (N_6186,N_5721,N_5463);
or U6187 (N_6187,N_5999,N_5207);
or U6188 (N_6188,N_5690,N_5473);
and U6189 (N_6189,N_5563,N_5090);
nand U6190 (N_6190,N_5545,N_5371);
nor U6191 (N_6191,N_5033,N_5673);
and U6192 (N_6192,N_5349,N_5761);
nand U6193 (N_6193,N_5092,N_5938);
nor U6194 (N_6194,N_5777,N_5021);
nor U6195 (N_6195,N_5668,N_5124);
and U6196 (N_6196,N_5024,N_5117);
nand U6197 (N_6197,N_5158,N_5984);
nor U6198 (N_6198,N_5737,N_5974);
or U6199 (N_6199,N_5016,N_5929);
or U6200 (N_6200,N_5657,N_5564);
and U6201 (N_6201,N_5570,N_5476);
or U6202 (N_6202,N_5393,N_5440);
and U6203 (N_6203,N_5026,N_5546);
or U6204 (N_6204,N_5928,N_5856);
or U6205 (N_6205,N_5516,N_5395);
nand U6206 (N_6206,N_5908,N_5970);
nor U6207 (N_6207,N_5404,N_5601);
nand U6208 (N_6208,N_5781,N_5559);
or U6209 (N_6209,N_5347,N_5784);
or U6210 (N_6210,N_5915,N_5305);
and U6211 (N_6211,N_5254,N_5232);
nor U6212 (N_6212,N_5635,N_5269);
and U6213 (N_6213,N_5062,N_5782);
xor U6214 (N_6214,N_5328,N_5238);
nor U6215 (N_6215,N_5138,N_5733);
or U6216 (N_6216,N_5081,N_5855);
or U6217 (N_6217,N_5979,N_5824);
and U6218 (N_6218,N_5697,N_5611);
nand U6219 (N_6219,N_5030,N_5355);
and U6220 (N_6220,N_5281,N_5362);
and U6221 (N_6221,N_5406,N_5038);
or U6222 (N_6222,N_5205,N_5003);
nor U6223 (N_6223,N_5740,N_5443);
and U6224 (N_6224,N_5116,N_5461);
or U6225 (N_6225,N_5667,N_5744);
or U6226 (N_6226,N_5857,N_5820);
and U6227 (N_6227,N_5749,N_5985);
and U6228 (N_6228,N_5170,N_5639);
nand U6229 (N_6229,N_5560,N_5113);
nor U6230 (N_6230,N_5968,N_5055);
nor U6231 (N_6231,N_5794,N_5550);
nand U6232 (N_6232,N_5735,N_5895);
nor U6233 (N_6233,N_5528,N_5770);
and U6234 (N_6234,N_5105,N_5368);
nand U6235 (N_6235,N_5747,N_5296);
or U6236 (N_6236,N_5574,N_5188);
and U6237 (N_6237,N_5453,N_5791);
and U6238 (N_6238,N_5561,N_5500);
nor U6239 (N_6239,N_5593,N_5757);
and U6240 (N_6240,N_5944,N_5916);
and U6241 (N_6241,N_5981,N_5109);
or U6242 (N_6242,N_5329,N_5173);
and U6243 (N_6243,N_5162,N_5795);
or U6244 (N_6244,N_5724,N_5243);
nor U6245 (N_6245,N_5365,N_5651);
nand U6246 (N_6246,N_5402,N_5086);
and U6247 (N_6247,N_5900,N_5524);
and U6248 (N_6248,N_5752,N_5200);
nand U6249 (N_6249,N_5990,N_5050);
or U6250 (N_6250,N_5475,N_5289);
or U6251 (N_6251,N_5739,N_5789);
or U6252 (N_6252,N_5687,N_5460);
nor U6253 (N_6253,N_5320,N_5840);
or U6254 (N_6254,N_5861,N_5373);
or U6255 (N_6255,N_5258,N_5802);
and U6256 (N_6256,N_5504,N_5447);
xor U6257 (N_6257,N_5077,N_5215);
and U6258 (N_6258,N_5449,N_5972);
nor U6259 (N_6259,N_5060,N_5419);
or U6260 (N_6260,N_5607,N_5186);
and U6261 (N_6261,N_5598,N_5309);
nand U6262 (N_6262,N_5803,N_5439);
or U6263 (N_6263,N_5532,N_5178);
nor U6264 (N_6264,N_5065,N_5816);
nand U6265 (N_6265,N_5619,N_5267);
nor U6266 (N_6266,N_5342,N_5230);
xnor U6267 (N_6267,N_5426,N_5905);
or U6268 (N_6268,N_5566,N_5682);
and U6269 (N_6269,N_5870,N_5143);
nor U6270 (N_6270,N_5620,N_5017);
or U6271 (N_6271,N_5920,N_5605);
nor U6272 (N_6272,N_5625,N_5827);
nor U6273 (N_6273,N_5009,N_5808);
nand U6274 (N_6274,N_5031,N_5495);
nor U6275 (N_6275,N_5760,N_5120);
nand U6276 (N_6276,N_5521,N_5948);
and U6277 (N_6277,N_5316,N_5745);
nor U6278 (N_6278,N_5604,N_5892);
nor U6279 (N_6279,N_5261,N_5023);
xnor U6280 (N_6280,N_5146,N_5123);
nor U6281 (N_6281,N_5591,N_5089);
nand U6282 (N_6282,N_5411,N_5634);
nor U6283 (N_6283,N_5107,N_5864);
nor U6284 (N_6284,N_5335,N_5514);
xor U6285 (N_6285,N_5302,N_5825);
nand U6286 (N_6286,N_5646,N_5691);
or U6287 (N_6287,N_5676,N_5454);
and U6288 (N_6288,N_5414,N_5898);
or U6289 (N_6289,N_5409,N_5496);
nor U6290 (N_6290,N_5633,N_5432);
nand U6291 (N_6291,N_5771,N_5630);
and U6292 (N_6292,N_5043,N_5417);
nor U6293 (N_6293,N_5530,N_5982);
or U6294 (N_6294,N_5240,N_5288);
nand U6295 (N_6295,N_5076,N_5953);
nand U6296 (N_6296,N_5027,N_5010);
and U6297 (N_6297,N_5636,N_5201);
and U6298 (N_6298,N_5727,N_5832);
or U6299 (N_6299,N_5012,N_5706);
or U6300 (N_6300,N_5956,N_5736);
nand U6301 (N_6301,N_5438,N_5082);
and U6302 (N_6302,N_5234,N_5301);
or U6303 (N_6303,N_5833,N_5723);
nor U6304 (N_6304,N_5133,N_5539);
and U6305 (N_6305,N_5911,N_5606);
nand U6306 (N_6306,N_5244,N_5358);
or U6307 (N_6307,N_5470,N_5952);
nor U6308 (N_6308,N_5555,N_5235);
and U6309 (N_6309,N_5345,N_5576);
nor U6310 (N_6310,N_5356,N_5954);
and U6311 (N_6311,N_5088,N_5921);
and U6312 (N_6312,N_5185,N_5474);
nand U6313 (N_6313,N_5505,N_5919);
and U6314 (N_6314,N_5482,N_5937);
nor U6315 (N_6315,N_5330,N_5127);
nand U6316 (N_6316,N_5614,N_5159);
nor U6317 (N_6317,N_5897,N_5095);
nand U6318 (N_6318,N_5002,N_5130);
nor U6319 (N_6319,N_5341,N_5674);
nand U6320 (N_6320,N_5797,N_5433);
nor U6321 (N_6321,N_5529,N_5885);
nand U6322 (N_6322,N_5172,N_5194);
or U6323 (N_6323,N_5945,N_5678);
or U6324 (N_6324,N_5019,N_5940);
nor U6325 (N_6325,N_5387,N_5213);
or U6326 (N_6326,N_5013,N_5711);
and U6327 (N_6327,N_5534,N_5381);
or U6328 (N_6328,N_5174,N_5996);
and U6329 (N_6329,N_5949,N_5445);
or U6330 (N_6330,N_5748,N_5425);
nand U6331 (N_6331,N_5732,N_5306);
xor U6332 (N_6332,N_5446,N_5069);
or U6333 (N_6333,N_5352,N_5686);
and U6334 (N_6334,N_5624,N_5863);
or U6335 (N_6335,N_5237,N_5538);
nor U6336 (N_6336,N_5692,N_5494);
nor U6337 (N_6337,N_5233,N_5300);
or U6338 (N_6338,N_5204,N_5214);
or U6339 (N_6339,N_5008,N_5629);
nor U6340 (N_6340,N_5154,N_5793);
and U6341 (N_6341,N_5080,N_5700);
nor U6342 (N_6342,N_5287,N_5644);
nand U6343 (N_6343,N_5403,N_5746);
and U6344 (N_6344,N_5083,N_5627);
and U6345 (N_6345,N_5862,N_5798);
nand U6346 (N_6346,N_5466,N_5052);
nand U6347 (N_6347,N_5645,N_5507);
nand U6348 (N_6348,N_5715,N_5337);
and U6349 (N_6349,N_5567,N_5525);
and U6350 (N_6350,N_5257,N_5377);
and U6351 (N_6351,N_5199,N_5372);
and U6352 (N_6352,N_5502,N_5814);
nand U6353 (N_6353,N_5139,N_5728);
nor U6354 (N_6354,N_5562,N_5685);
or U6355 (N_6355,N_5497,N_5308);
nor U6356 (N_6356,N_5638,N_5118);
nand U6357 (N_6357,N_5734,N_5079);
nand U6358 (N_6358,N_5577,N_5926);
or U6359 (N_6359,N_5653,N_5714);
nand U6360 (N_6360,N_5196,N_5047);
and U6361 (N_6361,N_5087,N_5094);
nor U6362 (N_6362,N_5575,N_5626);
nor U6363 (N_6363,N_5913,N_5430);
nand U6364 (N_6364,N_5994,N_5100);
or U6365 (N_6365,N_5681,N_5275);
or U6366 (N_6366,N_5506,N_5696);
and U6367 (N_6367,N_5594,N_5787);
nor U6368 (N_6368,N_5114,N_5935);
and U6369 (N_6369,N_5115,N_5078);
nor U6370 (N_6370,N_5780,N_5664);
and U6371 (N_6371,N_5326,N_5312);
or U6372 (N_6372,N_5398,N_5875);
nand U6373 (N_6373,N_5163,N_5459);
and U6374 (N_6374,N_5792,N_5818);
or U6375 (N_6375,N_5483,N_5311);
nor U6376 (N_6376,N_5348,N_5585);
nor U6377 (N_6377,N_5963,N_5596);
or U6378 (N_6378,N_5868,N_5325);
nand U6379 (N_6379,N_5175,N_5339);
or U6380 (N_6380,N_5187,N_5847);
or U6381 (N_6381,N_5331,N_5209);
xnor U6382 (N_6382,N_5775,N_5014);
nor U6383 (N_6383,N_5354,N_5084);
or U6384 (N_6384,N_5273,N_5044);
and U6385 (N_6385,N_5225,N_5640);
and U6386 (N_6386,N_5152,N_5408);
nor U6387 (N_6387,N_5537,N_5800);
and U6388 (N_6388,N_5045,N_5126);
or U6389 (N_6389,N_5412,N_5806);
nor U6390 (N_6390,N_5057,N_5569);
nand U6391 (N_6391,N_5303,N_5642);
or U6392 (N_6392,N_5394,N_5227);
and U6393 (N_6393,N_5102,N_5964);
and U6394 (N_6394,N_5880,N_5992);
nand U6395 (N_6395,N_5441,N_5164);
nand U6396 (N_6396,N_5277,N_5589);
nand U6397 (N_6397,N_5643,N_5378);
nor U6398 (N_6398,N_5501,N_5670);
and U6399 (N_6399,N_5096,N_5376);
nor U6400 (N_6400,N_5618,N_5796);
or U6401 (N_6401,N_5980,N_5878);
nor U6402 (N_6402,N_5383,N_5903);
nor U6403 (N_6403,N_5498,N_5583);
nand U6404 (N_6404,N_5717,N_5179);
nand U6405 (N_6405,N_5042,N_5819);
nand U6406 (N_6406,N_5375,N_5648);
nor U6407 (N_6407,N_5993,N_5758);
nand U6408 (N_6408,N_5801,N_5247);
or U6409 (N_6409,N_5718,N_5890);
or U6410 (N_6410,N_5535,N_5061);
or U6411 (N_6411,N_5987,N_5828);
nor U6412 (N_6412,N_5177,N_5386);
or U6413 (N_6413,N_5568,N_5321);
nand U6414 (N_6414,N_5141,N_5416);
and U6415 (N_6415,N_5290,N_5165);
nand U6416 (N_6416,N_5168,N_5369);
or U6417 (N_6417,N_5285,N_5965);
nor U6418 (N_6418,N_5292,N_5462);
or U6419 (N_6419,N_5068,N_5641);
nor U6420 (N_6420,N_5161,N_5698);
and U6421 (N_6421,N_5571,N_5029);
and U6422 (N_6422,N_5022,N_5181);
nor U6423 (N_6423,N_5671,N_5360);
nor U6424 (N_6424,N_5456,N_5242);
or U6425 (N_6425,N_5904,N_5669);
and U6426 (N_6426,N_5572,N_5826);
or U6427 (N_6427,N_5246,N_5726);
and U6428 (N_6428,N_5695,N_5392);
and U6429 (N_6429,N_5423,N_5955);
or U6430 (N_6430,N_5011,N_5677);
and U6431 (N_6431,N_5478,N_5586);
nor U6432 (N_6432,N_5991,N_5750);
nand U6433 (N_6433,N_5385,N_5912);
and U6434 (N_6434,N_5854,N_5259);
and U6435 (N_6435,N_5658,N_5363);
or U6436 (N_6436,N_5131,N_5338);
and U6437 (N_6437,N_5216,N_5631);
nor U6438 (N_6438,N_5073,N_5249);
and U6439 (N_6439,N_5121,N_5192);
nand U6440 (N_6440,N_5680,N_5701);
nand U6441 (N_6441,N_5415,N_5401);
or U6442 (N_6442,N_5704,N_5925);
and U6443 (N_6443,N_5085,N_5333);
nand U6444 (N_6444,N_5319,N_5960);
nand U6445 (N_6445,N_5527,N_5410);
or U6446 (N_6446,N_5513,N_5679);
or U6447 (N_6447,N_5966,N_5831);
xnor U6448 (N_6448,N_5608,N_5899);
and U6449 (N_6449,N_5536,N_5059);
nor U6450 (N_6450,N_5262,N_5151);
nand U6451 (N_6451,N_5853,N_5241);
nor U6452 (N_6452,N_5813,N_5578);
or U6453 (N_6453,N_5552,N_5753);
nand U6454 (N_6454,N_5829,N_5334);
or U6455 (N_6455,N_5451,N_5988);
nor U6456 (N_6456,N_5931,N_5547);
and U6457 (N_6457,N_5548,N_5103);
or U6458 (N_6458,N_5137,N_5450);
nor U6459 (N_6459,N_5324,N_5000);
and U6460 (N_6460,N_5040,N_5731);
or U6461 (N_6461,N_5860,N_5490);
nor U6462 (N_6462,N_5888,N_5049);
or U6463 (N_6463,N_5971,N_5488);
nor U6464 (N_6464,N_5428,N_5098);
or U6465 (N_6465,N_5756,N_5276);
nor U6466 (N_6466,N_5902,N_5374);
nand U6467 (N_6467,N_5554,N_5391);
nand U6468 (N_6468,N_5424,N_5004);
nor U6469 (N_6469,N_5517,N_5295);
or U6470 (N_6470,N_5028,N_5844);
or U6471 (N_6471,N_5544,N_5074);
nor U6472 (N_6472,N_5976,N_5155);
and U6473 (N_6473,N_5304,N_5351);
nor U6474 (N_6474,N_5997,N_5206);
nor U6475 (N_6475,N_5379,N_5923);
nand U6476 (N_6476,N_5859,N_5491);
or U6477 (N_6477,N_5767,N_5549);
nand U6478 (N_6478,N_5183,N_5219);
nand U6479 (N_6479,N_5122,N_5350);
nand U6480 (N_6480,N_5469,N_5977);
nor U6481 (N_6481,N_5252,N_5067);
nand U6482 (N_6482,N_5869,N_5652);
or U6483 (N_6483,N_5936,N_5587);
or U6484 (N_6484,N_5405,N_5930);
nor U6485 (N_6485,N_5851,N_5222);
and U6486 (N_6486,N_5615,N_5167);
or U6487 (N_6487,N_5946,N_5221);
and U6488 (N_6488,N_5286,N_5580);
nand U6489 (N_6489,N_5007,N_5472);
nor U6490 (N_6490,N_5367,N_5032);
and U6491 (N_6491,N_5359,N_5458);
nand U6492 (N_6492,N_5489,N_5493);
or U6493 (N_6493,N_5422,N_5906);
nor U6494 (N_6494,N_5713,N_5896);
xnor U6495 (N_6495,N_5001,N_5541);
nor U6496 (N_6496,N_5650,N_5556);
and U6497 (N_6497,N_5655,N_5176);
nand U6498 (N_6498,N_5418,N_5684);
or U6499 (N_6499,N_5783,N_5313);
nor U6500 (N_6500,N_5332,N_5579);
or U6501 (N_6501,N_5379,N_5431);
or U6502 (N_6502,N_5785,N_5816);
nand U6503 (N_6503,N_5996,N_5897);
nor U6504 (N_6504,N_5668,N_5673);
or U6505 (N_6505,N_5516,N_5738);
nor U6506 (N_6506,N_5599,N_5201);
nor U6507 (N_6507,N_5815,N_5840);
and U6508 (N_6508,N_5580,N_5318);
nor U6509 (N_6509,N_5401,N_5038);
nor U6510 (N_6510,N_5995,N_5084);
nor U6511 (N_6511,N_5603,N_5935);
nand U6512 (N_6512,N_5674,N_5104);
nand U6513 (N_6513,N_5746,N_5188);
nor U6514 (N_6514,N_5937,N_5678);
nand U6515 (N_6515,N_5202,N_5261);
xor U6516 (N_6516,N_5930,N_5803);
or U6517 (N_6517,N_5431,N_5095);
or U6518 (N_6518,N_5601,N_5032);
and U6519 (N_6519,N_5885,N_5659);
nor U6520 (N_6520,N_5888,N_5838);
nor U6521 (N_6521,N_5304,N_5428);
and U6522 (N_6522,N_5782,N_5275);
or U6523 (N_6523,N_5119,N_5358);
or U6524 (N_6524,N_5511,N_5166);
nor U6525 (N_6525,N_5479,N_5742);
nand U6526 (N_6526,N_5044,N_5253);
nand U6527 (N_6527,N_5140,N_5069);
nand U6528 (N_6528,N_5832,N_5619);
nand U6529 (N_6529,N_5169,N_5325);
and U6530 (N_6530,N_5720,N_5428);
nand U6531 (N_6531,N_5003,N_5509);
or U6532 (N_6532,N_5424,N_5193);
nor U6533 (N_6533,N_5766,N_5128);
nor U6534 (N_6534,N_5511,N_5803);
or U6535 (N_6535,N_5032,N_5496);
and U6536 (N_6536,N_5229,N_5392);
nor U6537 (N_6537,N_5471,N_5807);
and U6538 (N_6538,N_5640,N_5236);
xor U6539 (N_6539,N_5089,N_5793);
nor U6540 (N_6540,N_5929,N_5151);
nor U6541 (N_6541,N_5738,N_5866);
nor U6542 (N_6542,N_5536,N_5350);
nor U6543 (N_6543,N_5070,N_5040);
xnor U6544 (N_6544,N_5086,N_5409);
or U6545 (N_6545,N_5389,N_5581);
and U6546 (N_6546,N_5825,N_5733);
or U6547 (N_6547,N_5367,N_5735);
nand U6548 (N_6548,N_5635,N_5990);
nand U6549 (N_6549,N_5700,N_5213);
or U6550 (N_6550,N_5856,N_5989);
and U6551 (N_6551,N_5103,N_5832);
and U6552 (N_6552,N_5387,N_5644);
or U6553 (N_6553,N_5920,N_5088);
nor U6554 (N_6554,N_5601,N_5321);
and U6555 (N_6555,N_5339,N_5024);
or U6556 (N_6556,N_5992,N_5121);
xor U6557 (N_6557,N_5265,N_5959);
nor U6558 (N_6558,N_5830,N_5880);
nand U6559 (N_6559,N_5608,N_5876);
or U6560 (N_6560,N_5658,N_5021);
xnor U6561 (N_6561,N_5666,N_5132);
or U6562 (N_6562,N_5836,N_5899);
or U6563 (N_6563,N_5536,N_5906);
nand U6564 (N_6564,N_5835,N_5882);
xor U6565 (N_6565,N_5214,N_5058);
nor U6566 (N_6566,N_5637,N_5052);
and U6567 (N_6567,N_5155,N_5857);
nand U6568 (N_6568,N_5770,N_5226);
nand U6569 (N_6569,N_5241,N_5830);
nand U6570 (N_6570,N_5798,N_5928);
nor U6571 (N_6571,N_5562,N_5313);
and U6572 (N_6572,N_5883,N_5142);
or U6573 (N_6573,N_5158,N_5548);
xnor U6574 (N_6574,N_5279,N_5060);
and U6575 (N_6575,N_5324,N_5567);
nor U6576 (N_6576,N_5797,N_5063);
nand U6577 (N_6577,N_5166,N_5994);
or U6578 (N_6578,N_5340,N_5221);
and U6579 (N_6579,N_5474,N_5213);
or U6580 (N_6580,N_5431,N_5320);
nand U6581 (N_6581,N_5183,N_5128);
and U6582 (N_6582,N_5782,N_5918);
nand U6583 (N_6583,N_5676,N_5854);
nand U6584 (N_6584,N_5023,N_5448);
xor U6585 (N_6585,N_5337,N_5378);
nand U6586 (N_6586,N_5669,N_5256);
nor U6587 (N_6587,N_5825,N_5183);
or U6588 (N_6588,N_5458,N_5274);
nand U6589 (N_6589,N_5684,N_5930);
nor U6590 (N_6590,N_5720,N_5229);
nand U6591 (N_6591,N_5117,N_5492);
or U6592 (N_6592,N_5003,N_5355);
and U6593 (N_6593,N_5226,N_5689);
nand U6594 (N_6594,N_5736,N_5094);
or U6595 (N_6595,N_5682,N_5085);
and U6596 (N_6596,N_5661,N_5201);
nand U6597 (N_6597,N_5850,N_5099);
nor U6598 (N_6598,N_5145,N_5683);
and U6599 (N_6599,N_5550,N_5563);
and U6600 (N_6600,N_5183,N_5760);
and U6601 (N_6601,N_5528,N_5006);
or U6602 (N_6602,N_5047,N_5552);
or U6603 (N_6603,N_5962,N_5822);
nand U6604 (N_6604,N_5914,N_5180);
nor U6605 (N_6605,N_5088,N_5440);
or U6606 (N_6606,N_5123,N_5430);
or U6607 (N_6607,N_5913,N_5630);
nand U6608 (N_6608,N_5554,N_5094);
nand U6609 (N_6609,N_5566,N_5576);
nor U6610 (N_6610,N_5064,N_5562);
nor U6611 (N_6611,N_5952,N_5761);
nor U6612 (N_6612,N_5608,N_5049);
nor U6613 (N_6613,N_5561,N_5395);
nand U6614 (N_6614,N_5560,N_5955);
nand U6615 (N_6615,N_5290,N_5125);
nor U6616 (N_6616,N_5167,N_5685);
and U6617 (N_6617,N_5633,N_5863);
and U6618 (N_6618,N_5449,N_5632);
nand U6619 (N_6619,N_5233,N_5816);
xor U6620 (N_6620,N_5401,N_5681);
and U6621 (N_6621,N_5701,N_5835);
or U6622 (N_6622,N_5985,N_5732);
nor U6623 (N_6623,N_5940,N_5887);
or U6624 (N_6624,N_5300,N_5564);
nand U6625 (N_6625,N_5987,N_5959);
nor U6626 (N_6626,N_5585,N_5193);
nand U6627 (N_6627,N_5531,N_5753);
nand U6628 (N_6628,N_5299,N_5912);
xnor U6629 (N_6629,N_5968,N_5871);
or U6630 (N_6630,N_5504,N_5008);
xnor U6631 (N_6631,N_5436,N_5675);
or U6632 (N_6632,N_5302,N_5022);
nand U6633 (N_6633,N_5344,N_5364);
nand U6634 (N_6634,N_5586,N_5976);
and U6635 (N_6635,N_5976,N_5882);
xnor U6636 (N_6636,N_5406,N_5360);
and U6637 (N_6637,N_5382,N_5902);
nand U6638 (N_6638,N_5975,N_5408);
nand U6639 (N_6639,N_5128,N_5889);
xor U6640 (N_6640,N_5694,N_5863);
and U6641 (N_6641,N_5733,N_5427);
and U6642 (N_6642,N_5619,N_5796);
and U6643 (N_6643,N_5177,N_5309);
and U6644 (N_6644,N_5903,N_5910);
nor U6645 (N_6645,N_5332,N_5035);
or U6646 (N_6646,N_5533,N_5053);
nand U6647 (N_6647,N_5870,N_5892);
and U6648 (N_6648,N_5742,N_5990);
nor U6649 (N_6649,N_5675,N_5443);
nor U6650 (N_6650,N_5912,N_5633);
and U6651 (N_6651,N_5659,N_5790);
and U6652 (N_6652,N_5649,N_5588);
or U6653 (N_6653,N_5222,N_5921);
nand U6654 (N_6654,N_5477,N_5875);
nand U6655 (N_6655,N_5355,N_5635);
nand U6656 (N_6656,N_5396,N_5120);
nand U6657 (N_6657,N_5699,N_5827);
or U6658 (N_6658,N_5526,N_5733);
or U6659 (N_6659,N_5940,N_5353);
nor U6660 (N_6660,N_5453,N_5676);
nand U6661 (N_6661,N_5044,N_5004);
or U6662 (N_6662,N_5384,N_5816);
or U6663 (N_6663,N_5142,N_5379);
nor U6664 (N_6664,N_5561,N_5414);
nand U6665 (N_6665,N_5554,N_5448);
nand U6666 (N_6666,N_5533,N_5982);
nand U6667 (N_6667,N_5840,N_5856);
nand U6668 (N_6668,N_5955,N_5749);
or U6669 (N_6669,N_5200,N_5974);
and U6670 (N_6670,N_5918,N_5301);
nand U6671 (N_6671,N_5455,N_5746);
or U6672 (N_6672,N_5739,N_5722);
or U6673 (N_6673,N_5961,N_5456);
nor U6674 (N_6674,N_5862,N_5302);
or U6675 (N_6675,N_5608,N_5930);
or U6676 (N_6676,N_5849,N_5911);
or U6677 (N_6677,N_5338,N_5813);
nor U6678 (N_6678,N_5150,N_5718);
nand U6679 (N_6679,N_5827,N_5631);
or U6680 (N_6680,N_5741,N_5983);
and U6681 (N_6681,N_5430,N_5257);
and U6682 (N_6682,N_5423,N_5336);
and U6683 (N_6683,N_5863,N_5300);
nand U6684 (N_6684,N_5953,N_5657);
nor U6685 (N_6685,N_5424,N_5310);
and U6686 (N_6686,N_5232,N_5984);
or U6687 (N_6687,N_5657,N_5508);
and U6688 (N_6688,N_5711,N_5729);
and U6689 (N_6689,N_5666,N_5817);
and U6690 (N_6690,N_5736,N_5988);
and U6691 (N_6691,N_5216,N_5125);
nand U6692 (N_6692,N_5813,N_5663);
nand U6693 (N_6693,N_5739,N_5221);
nor U6694 (N_6694,N_5745,N_5499);
or U6695 (N_6695,N_5914,N_5728);
and U6696 (N_6696,N_5525,N_5248);
or U6697 (N_6697,N_5488,N_5491);
nor U6698 (N_6698,N_5469,N_5013);
and U6699 (N_6699,N_5944,N_5767);
and U6700 (N_6700,N_5099,N_5123);
and U6701 (N_6701,N_5068,N_5741);
and U6702 (N_6702,N_5461,N_5330);
and U6703 (N_6703,N_5872,N_5591);
nand U6704 (N_6704,N_5439,N_5705);
nor U6705 (N_6705,N_5647,N_5345);
nor U6706 (N_6706,N_5382,N_5250);
xnor U6707 (N_6707,N_5614,N_5938);
nor U6708 (N_6708,N_5477,N_5549);
nand U6709 (N_6709,N_5392,N_5294);
and U6710 (N_6710,N_5540,N_5859);
nand U6711 (N_6711,N_5247,N_5775);
nor U6712 (N_6712,N_5701,N_5139);
nor U6713 (N_6713,N_5265,N_5056);
nor U6714 (N_6714,N_5452,N_5417);
nand U6715 (N_6715,N_5764,N_5842);
or U6716 (N_6716,N_5134,N_5678);
nand U6717 (N_6717,N_5106,N_5982);
nand U6718 (N_6718,N_5196,N_5539);
nand U6719 (N_6719,N_5721,N_5780);
nand U6720 (N_6720,N_5626,N_5748);
nor U6721 (N_6721,N_5033,N_5053);
and U6722 (N_6722,N_5120,N_5389);
nor U6723 (N_6723,N_5513,N_5968);
or U6724 (N_6724,N_5629,N_5213);
nor U6725 (N_6725,N_5472,N_5036);
xor U6726 (N_6726,N_5213,N_5976);
and U6727 (N_6727,N_5365,N_5358);
and U6728 (N_6728,N_5304,N_5300);
nor U6729 (N_6729,N_5821,N_5450);
and U6730 (N_6730,N_5719,N_5811);
and U6731 (N_6731,N_5752,N_5956);
nor U6732 (N_6732,N_5805,N_5349);
nor U6733 (N_6733,N_5480,N_5113);
and U6734 (N_6734,N_5867,N_5555);
or U6735 (N_6735,N_5924,N_5346);
nor U6736 (N_6736,N_5400,N_5939);
and U6737 (N_6737,N_5613,N_5509);
and U6738 (N_6738,N_5922,N_5367);
nor U6739 (N_6739,N_5232,N_5502);
and U6740 (N_6740,N_5496,N_5072);
nand U6741 (N_6741,N_5595,N_5578);
nand U6742 (N_6742,N_5818,N_5270);
and U6743 (N_6743,N_5510,N_5973);
or U6744 (N_6744,N_5808,N_5341);
and U6745 (N_6745,N_5050,N_5295);
or U6746 (N_6746,N_5816,N_5501);
nand U6747 (N_6747,N_5148,N_5818);
and U6748 (N_6748,N_5142,N_5946);
or U6749 (N_6749,N_5337,N_5890);
nor U6750 (N_6750,N_5837,N_5029);
xor U6751 (N_6751,N_5119,N_5336);
or U6752 (N_6752,N_5321,N_5358);
or U6753 (N_6753,N_5468,N_5254);
nand U6754 (N_6754,N_5711,N_5681);
nand U6755 (N_6755,N_5016,N_5277);
and U6756 (N_6756,N_5434,N_5800);
or U6757 (N_6757,N_5752,N_5014);
or U6758 (N_6758,N_5811,N_5067);
nor U6759 (N_6759,N_5801,N_5370);
nand U6760 (N_6760,N_5882,N_5515);
or U6761 (N_6761,N_5871,N_5941);
and U6762 (N_6762,N_5526,N_5041);
or U6763 (N_6763,N_5470,N_5971);
nor U6764 (N_6764,N_5515,N_5382);
nor U6765 (N_6765,N_5251,N_5327);
xnor U6766 (N_6766,N_5225,N_5586);
nor U6767 (N_6767,N_5021,N_5172);
nand U6768 (N_6768,N_5715,N_5357);
nand U6769 (N_6769,N_5433,N_5706);
nand U6770 (N_6770,N_5497,N_5424);
and U6771 (N_6771,N_5349,N_5516);
or U6772 (N_6772,N_5633,N_5149);
nor U6773 (N_6773,N_5666,N_5638);
nand U6774 (N_6774,N_5381,N_5237);
nor U6775 (N_6775,N_5575,N_5239);
nor U6776 (N_6776,N_5609,N_5907);
or U6777 (N_6777,N_5534,N_5060);
or U6778 (N_6778,N_5146,N_5867);
or U6779 (N_6779,N_5220,N_5710);
and U6780 (N_6780,N_5960,N_5022);
or U6781 (N_6781,N_5873,N_5081);
nor U6782 (N_6782,N_5876,N_5154);
or U6783 (N_6783,N_5574,N_5859);
nand U6784 (N_6784,N_5144,N_5270);
or U6785 (N_6785,N_5812,N_5432);
or U6786 (N_6786,N_5255,N_5771);
or U6787 (N_6787,N_5145,N_5898);
nor U6788 (N_6788,N_5759,N_5929);
nor U6789 (N_6789,N_5693,N_5143);
and U6790 (N_6790,N_5250,N_5581);
xnor U6791 (N_6791,N_5142,N_5652);
nand U6792 (N_6792,N_5079,N_5645);
and U6793 (N_6793,N_5417,N_5018);
and U6794 (N_6794,N_5599,N_5182);
and U6795 (N_6795,N_5051,N_5226);
nand U6796 (N_6796,N_5897,N_5423);
or U6797 (N_6797,N_5469,N_5641);
nor U6798 (N_6798,N_5499,N_5736);
or U6799 (N_6799,N_5506,N_5967);
xor U6800 (N_6800,N_5420,N_5411);
and U6801 (N_6801,N_5136,N_5965);
and U6802 (N_6802,N_5914,N_5312);
and U6803 (N_6803,N_5709,N_5084);
or U6804 (N_6804,N_5912,N_5139);
nor U6805 (N_6805,N_5528,N_5364);
nand U6806 (N_6806,N_5432,N_5325);
or U6807 (N_6807,N_5440,N_5394);
nor U6808 (N_6808,N_5423,N_5941);
xnor U6809 (N_6809,N_5431,N_5418);
or U6810 (N_6810,N_5162,N_5294);
nor U6811 (N_6811,N_5394,N_5744);
or U6812 (N_6812,N_5917,N_5847);
or U6813 (N_6813,N_5889,N_5138);
nor U6814 (N_6814,N_5533,N_5364);
nor U6815 (N_6815,N_5051,N_5997);
xor U6816 (N_6816,N_5211,N_5154);
or U6817 (N_6817,N_5868,N_5244);
and U6818 (N_6818,N_5238,N_5932);
nor U6819 (N_6819,N_5340,N_5316);
and U6820 (N_6820,N_5415,N_5991);
and U6821 (N_6821,N_5406,N_5428);
nand U6822 (N_6822,N_5106,N_5944);
nand U6823 (N_6823,N_5559,N_5338);
or U6824 (N_6824,N_5327,N_5295);
and U6825 (N_6825,N_5264,N_5065);
and U6826 (N_6826,N_5009,N_5724);
nand U6827 (N_6827,N_5418,N_5053);
and U6828 (N_6828,N_5794,N_5365);
nand U6829 (N_6829,N_5152,N_5186);
nand U6830 (N_6830,N_5297,N_5620);
and U6831 (N_6831,N_5649,N_5943);
nand U6832 (N_6832,N_5003,N_5976);
and U6833 (N_6833,N_5273,N_5340);
nor U6834 (N_6834,N_5217,N_5905);
nand U6835 (N_6835,N_5557,N_5076);
nor U6836 (N_6836,N_5486,N_5124);
nor U6837 (N_6837,N_5409,N_5607);
nand U6838 (N_6838,N_5900,N_5777);
nand U6839 (N_6839,N_5130,N_5561);
nor U6840 (N_6840,N_5389,N_5635);
xor U6841 (N_6841,N_5006,N_5457);
nor U6842 (N_6842,N_5590,N_5036);
nand U6843 (N_6843,N_5759,N_5871);
and U6844 (N_6844,N_5069,N_5314);
xor U6845 (N_6845,N_5834,N_5044);
nor U6846 (N_6846,N_5331,N_5717);
nor U6847 (N_6847,N_5025,N_5858);
nand U6848 (N_6848,N_5803,N_5487);
and U6849 (N_6849,N_5692,N_5566);
nand U6850 (N_6850,N_5902,N_5878);
nor U6851 (N_6851,N_5571,N_5121);
and U6852 (N_6852,N_5817,N_5289);
nand U6853 (N_6853,N_5914,N_5620);
or U6854 (N_6854,N_5502,N_5892);
nand U6855 (N_6855,N_5767,N_5494);
nand U6856 (N_6856,N_5858,N_5070);
and U6857 (N_6857,N_5228,N_5007);
nand U6858 (N_6858,N_5572,N_5844);
nor U6859 (N_6859,N_5471,N_5827);
nor U6860 (N_6860,N_5126,N_5660);
nor U6861 (N_6861,N_5207,N_5323);
nor U6862 (N_6862,N_5230,N_5090);
nand U6863 (N_6863,N_5316,N_5540);
and U6864 (N_6864,N_5080,N_5252);
nand U6865 (N_6865,N_5311,N_5743);
and U6866 (N_6866,N_5466,N_5761);
or U6867 (N_6867,N_5973,N_5534);
nor U6868 (N_6868,N_5003,N_5892);
xor U6869 (N_6869,N_5570,N_5344);
nand U6870 (N_6870,N_5784,N_5767);
nand U6871 (N_6871,N_5944,N_5019);
or U6872 (N_6872,N_5836,N_5320);
and U6873 (N_6873,N_5632,N_5661);
nand U6874 (N_6874,N_5424,N_5818);
nand U6875 (N_6875,N_5891,N_5868);
and U6876 (N_6876,N_5575,N_5171);
nor U6877 (N_6877,N_5912,N_5609);
xnor U6878 (N_6878,N_5340,N_5219);
nand U6879 (N_6879,N_5104,N_5553);
xor U6880 (N_6880,N_5747,N_5184);
and U6881 (N_6881,N_5851,N_5502);
nand U6882 (N_6882,N_5800,N_5594);
and U6883 (N_6883,N_5837,N_5742);
and U6884 (N_6884,N_5598,N_5410);
nand U6885 (N_6885,N_5339,N_5859);
nor U6886 (N_6886,N_5321,N_5226);
nand U6887 (N_6887,N_5205,N_5956);
and U6888 (N_6888,N_5983,N_5946);
nor U6889 (N_6889,N_5054,N_5328);
nor U6890 (N_6890,N_5088,N_5796);
nor U6891 (N_6891,N_5870,N_5900);
nand U6892 (N_6892,N_5845,N_5790);
and U6893 (N_6893,N_5189,N_5125);
nor U6894 (N_6894,N_5679,N_5312);
or U6895 (N_6895,N_5464,N_5811);
xor U6896 (N_6896,N_5810,N_5818);
and U6897 (N_6897,N_5409,N_5689);
and U6898 (N_6898,N_5023,N_5964);
nor U6899 (N_6899,N_5781,N_5336);
nand U6900 (N_6900,N_5071,N_5421);
or U6901 (N_6901,N_5394,N_5027);
xnor U6902 (N_6902,N_5508,N_5080);
and U6903 (N_6903,N_5184,N_5204);
nand U6904 (N_6904,N_5631,N_5127);
nand U6905 (N_6905,N_5230,N_5148);
nand U6906 (N_6906,N_5536,N_5087);
and U6907 (N_6907,N_5558,N_5116);
and U6908 (N_6908,N_5826,N_5691);
or U6909 (N_6909,N_5456,N_5086);
or U6910 (N_6910,N_5798,N_5313);
nor U6911 (N_6911,N_5266,N_5248);
nor U6912 (N_6912,N_5009,N_5042);
nor U6913 (N_6913,N_5562,N_5945);
nand U6914 (N_6914,N_5205,N_5084);
nor U6915 (N_6915,N_5777,N_5945);
nor U6916 (N_6916,N_5454,N_5844);
or U6917 (N_6917,N_5409,N_5548);
and U6918 (N_6918,N_5790,N_5714);
or U6919 (N_6919,N_5025,N_5004);
and U6920 (N_6920,N_5590,N_5647);
or U6921 (N_6921,N_5136,N_5665);
nand U6922 (N_6922,N_5108,N_5710);
nand U6923 (N_6923,N_5967,N_5754);
or U6924 (N_6924,N_5223,N_5595);
nor U6925 (N_6925,N_5123,N_5356);
or U6926 (N_6926,N_5704,N_5319);
and U6927 (N_6927,N_5544,N_5423);
nor U6928 (N_6928,N_5605,N_5118);
or U6929 (N_6929,N_5997,N_5450);
nand U6930 (N_6930,N_5994,N_5860);
xor U6931 (N_6931,N_5995,N_5731);
nor U6932 (N_6932,N_5741,N_5416);
and U6933 (N_6933,N_5398,N_5907);
or U6934 (N_6934,N_5285,N_5455);
nor U6935 (N_6935,N_5671,N_5876);
nand U6936 (N_6936,N_5137,N_5964);
or U6937 (N_6937,N_5501,N_5564);
nor U6938 (N_6938,N_5649,N_5966);
and U6939 (N_6939,N_5631,N_5324);
or U6940 (N_6940,N_5845,N_5663);
xnor U6941 (N_6941,N_5983,N_5024);
and U6942 (N_6942,N_5760,N_5712);
and U6943 (N_6943,N_5327,N_5162);
nor U6944 (N_6944,N_5149,N_5835);
or U6945 (N_6945,N_5833,N_5534);
nand U6946 (N_6946,N_5993,N_5771);
or U6947 (N_6947,N_5925,N_5468);
or U6948 (N_6948,N_5543,N_5951);
nand U6949 (N_6949,N_5689,N_5704);
nor U6950 (N_6950,N_5934,N_5733);
nor U6951 (N_6951,N_5212,N_5497);
nor U6952 (N_6952,N_5560,N_5725);
nand U6953 (N_6953,N_5054,N_5958);
and U6954 (N_6954,N_5316,N_5334);
or U6955 (N_6955,N_5004,N_5988);
nor U6956 (N_6956,N_5476,N_5090);
nor U6957 (N_6957,N_5705,N_5629);
nor U6958 (N_6958,N_5229,N_5618);
nand U6959 (N_6959,N_5435,N_5935);
or U6960 (N_6960,N_5091,N_5094);
or U6961 (N_6961,N_5100,N_5754);
and U6962 (N_6962,N_5854,N_5779);
nor U6963 (N_6963,N_5922,N_5581);
nor U6964 (N_6964,N_5272,N_5294);
nand U6965 (N_6965,N_5667,N_5722);
and U6966 (N_6966,N_5269,N_5831);
nor U6967 (N_6967,N_5086,N_5561);
and U6968 (N_6968,N_5541,N_5300);
nand U6969 (N_6969,N_5639,N_5099);
or U6970 (N_6970,N_5973,N_5867);
and U6971 (N_6971,N_5443,N_5332);
or U6972 (N_6972,N_5603,N_5223);
xnor U6973 (N_6973,N_5242,N_5284);
nor U6974 (N_6974,N_5874,N_5076);
and U6975 (N_6975,N_5338,N_5253);
nand U6976 (N_6976,N_5347,N_5629);
or U6977 (N_6977,N_5655,N_5601);
nand U6978 (N_6978,N_5296,N_5033);
or U6979 (N_6979,N_5707,N_5678);
and U6980 (N_6980,N_5215,N_5268);
and U6981 (N_6981,N_5357,N_5025);
nor U6982 (N_6982,N_5701,N_5555);
and U6983 (N_6983,N_5824,N_5246);
and U6984 (N_6984,N_5874,N_5907);
nor U6985 (N_6985,N_5606,N_5779);
nand U6986 (N_6986,N_5515,N_5045);
nand U6987 (N_6987,N_5630,N_5446);
nor U6988 (N_6988,N_5279,N_5064);
nor U6989 (N_6989,N_5196,N_5913);
nand U6990 (N_6990,N_5972,N_5035);
or U6991 (N_6991,N_5035,N_5356);
and U6992 (N_6992,N_5860,N_5082);
nor U6993 (N_6993,N_5765,N_5531);
nor U6994 (N_6994,N_5403,N_5205);
and U6995 (N_6995,N_5532,N_5313);
or U6996 (N_6996,N_5643,N_5449);
nor U6997 (N_6997,N_5694,N_5130);
nor U6998 (N_6998,N_5743,N_5759);
and U6999 (N_6999,N_5685,N_5384);
and U7000 (N_7000,N_6546,N_6069);
nand U7001 (N_7001,N_6732,N_6346);
or U7002 (N_7002,N_6739,N_6345);
or U7003 (N_7003,N_6397,N_6671);
and U7004 (N_7004,N_6216,N_6073);
or U7005 (N_7005,N_6609,N_6390);
nand U7006 (N_7006,N_6202,N_6068);
nor U7007 (N_7007,N_6638,N_6142);
and U7008 (N_7008,N_6600,N_6511);
nor U7009 (N_7009,N_6398,N_6439);
nand U7010 (N_7010,N_6574,N_6150);
or U7011 (N_7011,N_6370,N_6348);
nand U7012 (N_7012,N_6233,N_6502);
and U7013 (N_7013,N_6626,N_6571);
or U7014 (N_7014,N_6604,N_6186);
nand U7015 (N_7015,N_6723,N_6116);
and U7016 (N_7016,N_6608,N_6055);
nand U7017 (N_7017,N_6673,N_6475);
nor U7018 (N_7018,N_6735,N_6736);
or U7019 (N_7019,N_6588,N_6261);
or U7020 (N_7020,N_6619,N_6708);
and U7021 (N_7021,N_6407,N_6665);
nand U7022 (N_7022,N_6957,N_6895);
nor U7023 (N_7023,N_6305,N_6770);
or U7024 (N_7024,N_6935,N_6288);
nand U7025 (N_7025,N_6196,N_6717);
and U7026 (N_7026,N_6046,N_6765);
nand U7027 (N_7027,N_6238,N_6806);
and U7028 (N_7028,N_6644,N_6500);
and U7029 (N_7029,N_6654,N_6155);
and U7030 (N_7030,N_6760,N_6563);
and U7031 (N_7031,N_6713,N_6968);
nor U7032 (N_7032,N_6321,N_6698);
or U7033 (N_7033,N_6816,N_6389);
nor U7034 (N_7034,N_6249,N_6940);
nand U7035 (N_7035,N_6701,N_6464);
and U7036 (N_7036,N_6415,N_6484);
nor U7037 (N_7037,N_6289,N_6519);
nor U7038 (N_7038,N_6236,N_6531);
and U7039 (N_7039,N_6996,N_6171);
or U7040 (N_7040,N_6999,N_6232);
and U7041 (N_7041,N_6871,N_6905);
xnor U7042 (N_7042,N_6700,N_6720);
nor U7043 (N_7043,N_6727,N_6878);
and U7044 (N_7044,N_6589,N_6498);
nor U7045 (N_7045,N_6024,N_6877);
and U7046 (N_7046,N_6991,N_6075);
nand U7047 (N_7047,N_6280,N_6093);
xnor U7048 (N_7048,N_6958,N_6941);
nor U7049 (N_7049,N_6801,N_6317);
and U7050 (N_7050,N_6344,N_6924);
nand U7051 (N_7051,N_6356,N_6256);
and U7052 (N_7052,N_6688,N_6219);
or U7053 (N_7053,N_6306,N_6932);
and U7054 (N_7054,N_6143,N_6065);
and U7055 (N_7055,N_6781,N_6018);
or U7056 (N_7056,N_6663,N_6284);
or U7057 (N_7057,N_6897,N_6821);
nand U7058 (N_7058,N_6025,N_6326);
nand U7059 (N_7059,N_6315,N_6586);
and U7060 (N_7060,N_6056,N_6121);
nor U7061 (N_7061,N_6004,N_6165);
and U7062 (N_7062,N_6386,N_6445);
and U7063 (N_7063,N_6336,N_6988);
nor U7064 (N_7064,N_6487,N_6054);
or U7065 (N_7065,N_6862,N_6809);
or U7066 (N_7066,N_6434,N_6516);
nor U7067 (N_7067,N_6329,N_6140);
nand U7068 (N_7068,N_6613,N_6000);
and U7069 (N_7069,N_6677,N_6578);
nor U7070 (N_7070,N_6339,N_6179);
nand U7071 (N_7071,N_6485,N_6423);
and U7072 (N_7072,N_6522,N_6377);
nand U7073 (N_7073,N_6402,N_6625);
or U7074 (N_7074,N_6614,N_6915);
nor U7075 (N_7075,N_6972,N_6109);
nor U7076 (N_7076,N_6570,N_6031);
xor U7077 (N_7077,N_6145,N_6430);
and U7078 (N_7078,N_6208,N_6680);
nand U7079 (N_7079,N_6412,N_6361);
and U7080 (N_7080,N_6246,N_6852);
nand U7081 (N_7081,N_6505,N_6265);
or U7082 (N_7082,N_6598,N_6101);
or U7083 (N_7083,N_6785,N_6019);
or U7084 (N_7084,N_6763,N_6063);
nor U7085 (N_7085,N_6038,N_6911);
xnor U7086 (N_7086,N_6307,N_6777);
xor U7087 (N_7087,N_6242,N_6603);
nand U7088 (N_7088,N_6002,N_6567);
nand U7089 (N_7089,N_6125,N_6363);
or U7090 (N_7090,N_6615,N_6824);
nand U7091 (N_7091,N_6864,N_6380);
nand U7092 (N_7092,N_6008,N_6553);
or U7093 (N_7093,N_6836,N_6089);
nand U7094 (N_7094,N_6297,N_6168);
nand U7095 (N_7095,N_6985,N_6354);
nor U7096 (N_7096,N_6561,N_6893);
xnor U7097 (N_7097,N_6646,N_6802);
and U7098 (N_7098,N_6198,N_6514);
nand U7099 (N_7099,N_6926,N_6631);
xor U7100 (N_7100,N_6313,N_6870);
nor U7101 (N_7101,N_6748,N_6855);
or U7102 (N_7102,N_6755,N_6225);
nand U7103 (N_7103,N_6081,N_6020);
and U7104 (N_7104,N_6993,N_6979);
or U7105 (N_7105,N_6764,N_6092);
nor U7106 (N_7106,N_6136,N_6391);
nand U7107 (N_7107,N_6704,N_6449);
or U7108 (N_7108,N_6630,N_6820);
nor U7109 (N_7109,N_6263,N_6368);
or U7110 (N_7110,N_6118,N_6367);
nand U7111 (N_7111,N_6767,N_6119);
and U7112 (N_7112,N_6648,N_6460);
nand U7113 (N_7113,N_6994,N_6072);
nand U7114 (N_7114,N_6797,N_6813);
nand U7115 (N_7115,N_6021,N_6602);
nor U7116 (N_7116,N_6956,N_6314);
nand U7117 (N_7117,N_6917,N_6210);
nand U7118 (N_7118,N_6651,N_6928);
or U7119 (N_7119,N_6844,N_6827);
nand U7120 (N_7120,N_6756,N_6164);
and U7121 (N_7121,N_6403,N_6879);
nand U7122 (N_7122,N_6009,N_6962);
nand U7123 (N_7123,N_6859,N_6703);
nand U7124 (N_7124,N_6632,N_6845);
or U7125 (N_7125,N_6973,N_6240);
xnor U7126 (N_7126,N_6294,N_6441);
nand U7127 (N_7127,N_6465,N_6450);
or U7128 (N_7128,N_6691,N_6983);
nand U7129 (N_7129,N_6520,N_6894);
xor U7130 (N_7130,N_6846,N_6309);
and U7131 (N_7131,N_6507,N_6287);
and U7132 (N_7132,N_6085,N_6424);
and U7133 (N_7133,N_6998,N_6098);
nand U7134 (N_7134,N_6359,N_6599);
or U7135 (N_7135,N_6550,N_6784);
nor U7136 (N_7136,N_6396,N_6624);
nand U7137 (N_7137,N_6523,N_6524);
and U7138 (N_7138,N_6906,N_6180);
or U7139 (N_7139,N_6178,N_6733);
nor U7140 (N_7140,N_6851,N_6264);
and U7141 (N_7141,N_6823,N_6016);
and U7142 (N_7142,N_6921,N_6947);
or U7143 (N_7143,N_6577,N_6141);
nand U7144 (N_7144,N_6655,N_6003);
nand U7145 (N_7145,N_6048,N_6527);
and U7146 (N_7146,N_6095,N_6759);
and U7147 (N_7147,N_6462,N_6248);
or U7148 (N_7148,N_6130,N_6686);
or U7149 (N_7149,N_6010,N_6869);
xor U7150 (N_7150,N_6788,N_6942);
nor U7151 (N_7151,N_6173,N_6187);
nor U7152 (N_7152,N_6742,N_6714);
and U7153 (N_7153,N_6904,N_6409);
and U7154 (N_7154,N_6255,N_6637);
nor U7155 (N_7155,N_6298,N_6436);
or U7156 (N_7156,N_6352,N_6585);
nor U7157 (N_7157,N_6378,N_6576);
nand U7158 (N_7158,N_6030,N_6506);
and U7159 (N_7159,N_6918,N_6273);
or U7160 (N_7160,N_6192,N_6448);
and U7161 (N_7161,N_6997,N_6042);
xnor U7162 (N_7162,N_6283,N_6419);
and U7163 (N_7163,N_6177,N_6960);
nor U7164 (N_7164,N_6129,N_6382);
and U7165 (N_7165,N_6153,N_6395);
nor U7166 (N_7166,N_6780,N_6606);
nor U7167 (N_7167,N_6982,N_6104);
nor U7168 (N_7168,N_6071,N_6687);
and U7169 (N_7169,N_6067,N_6090);
nand U7170 (N_7170,N_6226,N_6260);
nor U7171 (N_7171,N_6454,N_6682);
and U7172 (N_7172,N_6185,N_6676);
or U7173 (N_7173,N_6244,N_6819);
and U7174 (N_7174,N_6222,N_6959);
and U7175 (N_7175,N_6047,N_6479);
nand U7176 (N_7176,N_6693,N_6931);
xnor U7177 (N_7177,N_6715,N_6817);
nor U7178 (N_7178,N_6954,N_6981);
and U7179 (N_7179,N_6400,N_6868);
nand U7180 (N_7180,N_6721,N_6621);
or U7181 (N_7181,N_6909,N_6132);
and U7182 (N_7182,N_6992,N_6131);
nor U7183 (N_7183,N_6182,N_6882);
and U7184 (N_7184,N_6889,N_6169);
nand U7185 (N_7185,N_6944,N_6333);
nor U7186 (N_7186,N_6933,N_6310);
nand U7187 (N_7187,N_6989,N_6938);
nor U7188 (N_7188,N_6568,N_6672);
nor U7189 (N_7189,N_6271,N_6835);
nand U7190 (N_7190,N_6683,N_6383);
nor U7191 (N_7191,N_6228,N_6496);
nor U7192 (N_7192,N_6681,N_6761);
or U7193 (N_7193,N_6416,N_6480);
nor U7194 (N_7194,N_6768,N_6694);
or U7195 (N_7195,N_6901,N_6752);
nand U7196 (N_7196,N_6828,N_6467);
or U7197 (N_7197,N_6203,N_6541);
nand U7198 (N_7198,N_6443,N_6799);
and U7199 (N_7199,N_6984,N_6552);
xor U7200 (N_7200,N_6778,N_6290);
nor U7201 (N_7201,N_6393,N_6808);
xor U7202 (N_7202,N_6741,N_6937);
and U7203 (N_7203,N_6980,N_6079);
or U7204 (N_7204,N_6478,N_6867);
or U7205 (N_7205,N_6731,N_6342);
and U7206 (N_7206,N_6295,N_6340);
or U7207 (N_7207,N_6034,N_6587);
nand U7208 (N_7208,N_6229,N_6495);
or U7209 (N_7209,N_6471,N_6668);
nand U7210 (N_7210,N_6257,N_6839);
and U7211 (N_7211,N_6650,N_6557);
or U7212 (N_7212,N_6302,N_6209);
and U7213 (N_7213,N_6213,N_6537);
and U7214 (N_7214,N_6746,N_6803);
and U7215 (N_7215,N_6757,N_6188);
nand U7216 (N_7216,N_6880,N_6087);
or U7217 (N_7217,N_6438,N_6250);
and U7218 (N_7218,N_6887,N_6706);
nor U7219 (N_7219,N_6322,N_6888);
nand U7220 (N_7220,N_6365,N_6842);
or U7221 (N_7221,N_6292,N_6634);
and U7222 (N_7222,N_6532,N_6328);
nand U7223 (N_7223,N_6312,N_6167);
nand U7224 (N_7224,N_6435,N_6040);
nand U7225 (N_7225,N_6388,N_6617);
nor U7226 (N_7226,N_6530,N_6951);
xnor U7227 (N_7227,N_6679,N_6105);
or U7228 (N_7228,N_6610,N_6123);
and U7229 (N_7229,N_6512,N_6433);
nand U7230 (N_7230,N_6633,N_6440);
nand U7231 (N_7231,N_6151,N_6783);
or U7232 (N_7232,N_6592,N_6555);
nand U7233 (N_7233,N_6920,N_6647);
or U7234 (N_7234,N_6394,N_6724);
nand U7235 (N_7235,N_6320,N_6896);
and U7236 (N_7236,N_6899,N_6157);
nor U7237 (N_7237,N_6127,N_6582);
and U7238 (N_7238,N_6750,N_6028);
and U7239 (N_7239,N_6176,N_6884);
xnor U7240 (N_7240,N_6133,N_6270);
nor U7241 (N_7241,N_6364,N_6074);
nor U7242 (N_7242,N_6111,N_6032);
and U7243 (N_7243,N_6707,N_6482);
and U7244 (N_7244,N_6375,N_6840);
nand U7245 (N_7245,N_6719,N_6622);
nor U7246 (N_7246,N_6734,N_6952);
or U7247 (N_7247,N_6853,N_6499);
nand U7248 (N_7248,N_6866,N_6103);
and U7249 (N_7249,N_6268,N_6045);
nand U7250 (N_7250,N_6080,N_6830);
xor U7251 (N_7251,N_6709,N_6689);
nand U7252 (N_7252,N_6543,N_6276);
nor U7253 (N_7253,N_6515,N_6108);
or U7254 (N_7254,N_6754,N_6749);
or U7255 (N_7255,N_6262,N_6408);
and U7256 (N_7256,N_6885,N_6170);
nand U7257 (N_7257,N_6976,N_6371);
nand U7258 (N_7258,N_6296,N_6274);
and U7259 (N_7259,N_6832,N_6861);
nor U7260 (N_7260,N_6334,N_6607);
or U7261 (N_7261,N_6955,N_6873);
nor U7262 (N_7262,N_6453,N_6540);
or U7263 (N_7263,N_6725,N_6774);
and U7264 (N_7264,N_6062,N_6892);
and U7265 (N_7265,N_6327,N_6946);
xor U7266 (N_7266,N_6597,N_6649);
or U7267 (N_7267,N_6191,N_6446);
nor U7268 (N_7268,N_6456,N_6833);
and U7269 (N_7269,N_6653,N_6122);
or U7270 (N_7270,N_6324,N_6061);
nor U7271 (N_7271,N_6037,N_6301);
or U7272 (N_7272,N_6579,N_6805);
nor U7273 (N_7273,N_6929,N_6117);
or U7274 (N_7274,N_6426,N_6147);
or U7275 (N_7275,N_6559,N_6970);
or U7276 (N_7276,N_6569,N_6641);
or U7277 (N_7277,N_6086,N_6964);
or U7278 (N_7278,N_6158,N_6697);
or U7279 (N_7279,N_6975,N_6775);
and U7280 (N_7280,N_6907,N_6206);
or U7281 (N_7281,N_6199,N_6154);
or U7282 (N_7282,N_6227,N_6044);
and U7283 (N_7283,N_6536,N_6126);
nand U7284 (N_7284,N_6110,N_6627);
and U7285 (N_7285,N_6927,N_6146);
nor U7286 (N_7286,N_6945,N_6266);
or U7287 (N_7287,N_6429,N_6195);
or U7288 (N_7288,N_6469,N_6645);
and U7289 (N_7289,N_6277,N_6476);
or U7290 (N_7290,N_6481,N_6762);
or U7291 (N_7291,N_6591,N_6427);
nor U7292 (N_7292,N_6751,N_6282);
or U7293 (N_7293,N_6883,N_6362);
and U7294 (N_7294,N_6793,N_6323);
nand U7295 (N_7295,N_6399,N_6548);
nand U7296 (N_7296,N_6337,N_6161);
or U7297 (N_7297,N_6912,N_6181);
or U7298 (N_7298,N_6084,N_6099);
or U7299 (N_7299,N_6696,N_6890);
nor U7300 (N_7300,N_6966,N_6451);
nand U7301 (N_7301,N_6269,N_6057);
and U7302 (N_7302,N_6776,N_6134);
and U7303 (N_7303,N_6488,N_6690);
or U7304 (N_7304,N_6669,N_6163);
or U7305 (N_7305,N_6369,N_6950);
or U7306 (N_7306,N_6251,N_6508);
or U7307 (N_7307,N_6967,N_6335);
and U7308 (N_7308,N_6566,N_6818);
nor U7309 (N_7309,N_6461,N_6442);
nor U7310 (N_7310,N_6102,N_6194);
nor U7311 (N_7311,N_6376,N_6737);
and U7312 (N_7312,N_6043,N_6373);
nand U7313 (N_7313,N_6138,N_6064);
or U7314 (N_7314,N_6790,N_6695);
or U7315 (N_7315,N_6285,N_6425);
or U7316 (N_7316,N_6652,N_6316);
nand U7317 (N_7317,N_6712,N_6560);
nor U7318 (N_7318,N_6913,N_6898);
and U7319 (N_7319,N_6015,N_6472);
nor U7320 (N_7320,N_6971,N_6549);
nand U7321 (N_7321,N_6815,N_6189);
nand U7322 (N_7322,N_6916,N_6458);
nand U7323 (N_7323,N_6636,N_6293);
and U7324 (N_7324,N_6214,N_6410);
or U7325 (N_7325,N_6060,N_6078);
or U7326 (N_7326,N_6299,N_6662);
xnor U7327 (N_7327,N_6418,N_6212);
nand U7328 (N_7328,N_6207,N_6466);
or U7329 (N_7329,N_6643,N_6711);
nor U7330 (N_7330,N_6573,N_6013);
and U7331 (N_7331,N_6304,N_6554);
nor U7332 (N_7332,N_6743,N_6534);
nor U7333 (N_7333,N_6059,N_6773);
and U7334 (N_7334,N_6457,N_6058);
and U7335 (N_7335,N_6347,N_6023);
nor U7336 (N_7336,N_6923,N_6053);
nor U7337 (N_7337,N_6990,N_6355);
and U7338 (N_7338,N_6657,N_6166);
nor U7339 (N_7339,N_6925,N_6175);
or U7340 (N_7340,N_6077,N_6794);
nand U7341 (N_7341,N_6738,N_6834);
and U7342 (N_7342,N_6772,N_6413);
nand U7343 (N_7343,N_6360,N_6358);
and U7344 (N_7344,N_6857,N_6629);
and U7345 (N_7345,N_6281,N_6740);
nand U7346 (N_7346,N_6831,N_6542);
nand U7347 (N_7347,N_6049,N_6217);
nand U7348 (N_7348,N_6097,N_6247);
nor U7349 (N_7349,N_6455,N_6468);
and U7350 (N_7350,N_6100,N_6528);
and U7351 (N_7351,N_6486,N_6353);
nand U7352 (N_7352,N_6432,N_6533);
nand U7353 (N_7353,N_6319,N_6675);
nand U7354 (N_7354,N_6826,N_6995);
nand U7355 (N_7355,N_6969,N_6786);
nand U7356 (N_7356,N_6135,N_6474);
nor U7357 (N_7357,N_6200,N_6572);
nand U7358 (N_7358,N_6350,N_6120);
xor U7359 (N_7359,N_6728,N_6437);
or U7360 (N_7360,N_6385,N_6332);
nor U7361 (N_7361,N_6193,N_6939);
and U7362 (N_7362,N_6144,N_6492);
and U7363 (N_7363,N_6856,N_6753);
or U7364 (N_7364,N_6091,N_6804);
nor U7365 (N_7365,N_6218,N_6308);
nand U7366 (N_7366,N_6076,N_6036);
or U7367 (N_7367,N_6201,N_6444);
or U7368 (N_7368,N_6148,N_6027);
or U7369 (N_7369,N_6903,N_6539);
and U7370 (N_7370,N_6594,N_6275);
nor U7371 (N_7371,N_6220,N_6529);
and U7372 (N_7372,N_6575,N_6494);
nor U7373 (N_7373,N_6230,N_6252);
or U7374 (N_7374,N_6318,N_6565);
or U7375 (N_7375,N_6891,N_6279);
nor U7376 (N_7376,N_6798,N_6473);
or U7377 (N_7377,N_6769,N_6149);
or U7378 (N_7378,N_6452,N_6729);
or U7379 (N_7379,N_6658,N_6900);
nor U7380 (N_7380,N_6605,N_6812);
nor U7381 (N_7381,N_6745,N_6006);
xor U7382 (N_7382,N_6544,N_6744);
nor U7383 (N_7383,N_6374,N_6387);
and U7384 (N_7384,N_6272,N_6493);
nor U7385 (N_7385,N_6595,N_6051);
xnor U7386 (N_7386,N_6183,N_6664);
or U7387 (N_7387,N_6501,N_6420);
or U7388 (N_7388,N_6303,N_6822);
nand U7389 (N_7389,N_6007,N_6463);
nor U7390 (N_7390,N_6267,N_6381);
nor U7391 (N_7391,N_6628,N_6779);
nand U7392 (N_7392,N_6112,N_6033);
nand U7393 (N_7393,N_6211,N_6291);
and U7394 (N_7394,N_6841,N_6243);
or U7395 (N_7395,N_6863,N_6716);
nor U7396 (N_7396,N_6223,N_6829);
nand U7397 (N_7397,N_6325,N_6490);
and U7398 (N_7398,N_6300,N_6612);
and U7399 (N_7399,N_6771,N_6551);
nor U7400 (N_7400,N_6949,N_6022);
or U7401 (N_7401,N_6810,N_6459);
and U7402 (N_7402,N_6963,N_6787);
nor U7403 (N_7403,N_6039,N_6160);
and U7404 (N_7404,N_6351,N_6562);
nand U7405 (N_7405,N_6096,N_6792);
nor U7406 (N_7406,N_6491,N_6366);
nand U7407 (N_7407,N_6766,N_6215);
nor U7408 (N_7408,N_6124,N_6384);
nand U7409 (N_7409,N_6847,N_6837);
or U7410 (N_7410,N_6881,N_6710);
and U7411 (N_7411,N_6667,N_6477);
xor U7412 (N_7412,N_6017,N_6666);
or U7413 (N_7413,N_6526,N_6747);
nand U7414 (N_7414,N_6235,N_6489);
or U7415 (N_7415,N_6417,N_6029);
and U7416 (N_7416,N_6796,N_6872);
nand U7417 (N_7417,N_6011,N_6580);
or U7418 (N_7418,N_6692,N_6874);
or U7419 (N_7419,N_6902,N_6807);
nor U7420 (N_7420,N_6876,N_6684);
and U7421 (N_7421,N_6886,N_6128);
nor U7422 (N_7422,N_6421,N_6838);
nand U7423 (N_7423,N_6858,N_6428);
nor U7424 (N_7424,N_6848,N_6914);
nor U7425 (N_7425,N_6854,N_6184);
nand U7426 (N_7426,N_6865,N_6259);
and U7427 (N_7427,N_6343,N_6814);
nor U7428 (N_7428,N_6330,N_6190);
or U7429 (N_7429,N_6618,N_6311);
or U7430 (N_7430,N_6699,N_6137);
nand U7431 (N_7431,N_6115,N_6593);
nor U7432 (N_7432,N_6372,N_6088);
nor U7433 (N_7433,N_6224,N_6558);
xor U7434 (N_7434,N_6504,N_6642);
nand U7435 (N_7435,N_6221,N_6050);
nand U7436 (N_7436,N_6258,N_6510);
nand U7437 (N_7437,N_6234,N_6422);
or U7438 (N_7438,N_6411,N_6497);
nand U7439 (N_7439,N_6965,N_6811);
xor U7440 (N_7440,N_6789,N_6556);
nand U7441 (N_7441,N_6782,N_6922);
nor U7442 (N_7442,N_6503,N_6107);
or U7443 (N_7443,N_6930,N_6678);
or U7444 (N_7444,N_6114,N_6919);
nor U7445 (N_7445,N_6843,N_6231);
nand U7446 (N_7446,N_6106,N_6616);
or U7447 (N_7447,N_6401,N_6656);
nor U7448 (N_7448,N_6948,N_6205);
and U7449 (N_7449,N_6583,N_6414);
or U7450 (N_7450,N_6910,N_6404);
nor U7451 (N_7451,N_6953,N_6082);
or U7452 (N_7452,N_6012,N_6239);
or U7453 (N_7453,N_6978,N_6518);
nand U7454 (N_7454,N_6718,N_6685);
xor U7455 (N_7455,N_6943,N_6172);
or U7456 (N_7456,N_6961,N_6525);
or U7457 (N_7457,N_6596,N_6509);
nor U7458 (N_7458,N_6139,N_6241);
or U7459 (N_7459,N_6670,N_6547);
nor U7460 (N_7460,N_6908,N_6405);
nand U7461 (N_7461,N_6156,N_6379);
nor U7462 (N_7462,N_6517,N_6825);
and U7463 (N_7463,N_6521,N_6850);
and U7464 (N_7464,N_6800,N_6623);
nor U7465 (N_7465,N_6174,N_6674);
and U7466 (N_7466,N_6791,N_6005);
nor U7467 (N_7467,N_6041,N_6035);
nand U7468 (N_7468,N_6849,N_6001);
and U7469 (N_7469,N_6639,N_6705);
and U7470 (N_7470,N_6661,N_6254);
nor U7471 (N_7471,N_6722,N_6795);
and U7472 (N_7472,N_6447,N_6584);
and U7473 (N_7473,N_6535,N_6513);
nor U7474 (N_7474,N_6094,N_6986);
or U7475 (N_7475,N_6357,N_6470);
nor U7476 (N_7476,N_6113,N_6014);
nor U7477 (N_7477,N_6083,N_6278);
and U7478 (N_7478,N_6162,N_6875);
or U7479 (N_7479,N_6204,N_6253);
and U7480 (N_7480,N_6331,N_6581);
nor U7481 (N_7481,N_6601,N_6730);
nor U7482 (N_7482,N_6758,N_6286);
or U7483 (N_7483,N_6934,N_6052);
nor U7484 (N_7484,N_6159,N_6860);
and U7485 (N_7485,N_6483,N_6564);
or U7486 (N_7486,N_6977,N_6066);
nand U7487 (N_7487,N_6070,N_6726);
nand U7488 (N_7488,N_6406,N_6392);
nand U7489 (N_7489,N_6538,N_6341);
xor U7490 (N_7490,N_6987,N_6431);
nand U7491 (N_7491,N_6640,N_6620);
or U7492 (N_7492,N_6026,N_6590);
nor U7493 (N_7493,N_6660,N_6545);
nand U7494 (N_7494,N_6611,N_6338);
nor U7495 (N_7495,N_6635,N_6702);
xor U7496 (N_7496,N_6197,N_6152);
nand U7497 (N_7497,N_6936,N_6237);
nand U7498 (N_7498,N_6974,N_6349);
nand U7499 (N_7499,N_6245,N_6659);
and U7500 (N_7500,N_6015,N_6123);
or U7501 (N_7501,N_6876,N_6868);
and U7502 (N_7502,N_6760,N_6861);
and U7503 (N_7503,N_6437,N_6972);
nand U7504 (N_7504,N_6004,N_6877);
xnor U7505 (N_7505,N_6388,N_6304);
nand U7506 (N_7506,N_6109,N_6156);
nand U7507 (N_7507,N_6397,N_6665);
and U7508 (N_7508,N_6741,N_6161);
nor U7509 (N_7509,N_6098,N_6543);
nor U7510 (N_7510,N_6884,N_6414);
and U7511 (N_7511,N_6682,N_6040);
nor U7512 (N_7512,N_6819,N_6210);
nor U7513 (N_7513,N_6572,N_6429);
or U7514 (N_7514,N_6770,N_6490);
nand U7515 (N_7515,N_6388,N_6459);
or U7516 (N_7516,N_6570,N_6362);
or U7517 (N_7517,N_6440,N_6997);
or U7518 (N_7518,N_6271,N_6079);
nand U7519 (N_7519,N_6700,N_6105);
and U7520 (N_7520,N_6014,N_6789);
nor U7521 (N_7521,N_6965,N_6301);
and U7522 (N_7522,N_6417,N_6469);
and U7523 (N_7523,N_6704,N_6146);
nor U7524 (N_7524,N_6784,N_6782);
nand U7525 (N_7525,N_6372,N_6802);
nand U7526 (N_7526,N_6027,N_6777);
or U7527 (N_7527,N_6689,N_6918);
and U7528 (N_7528,N_6904,N_6899);
nor U7529 (N_7529,N_6730,N_6671);
nand U7530 (N_7530,N_6565,N_6451);
and U7531 (N_7531,N_6468,N_6851);
or U7532 (N_7532,N_6382,N_6335);
or U7533 (N_7533,N_6929,N_6860);
nor U7534 (N_7534,N_6166,N_6340);
and U7535 (N_7535,N_6980,N_6976);
or U7536 (N_7536,N_6247,N_6227);
or U7537 (N_7537,N_6127,N_6325);
nand U7538 (N_7538,N_6668,N_6498);
and U7539 (N_7539,N_6822,N_6078);
nand U7540 (N_7540,N_6915,N_6743);
and U7541 (N_7541,N_6556,N_6292);
nor U7542 (N_7542,N_6086,N_6703);
nor U7543 (N_7543,N_6643,N_6034);
nor U7544 (N_7544,N_6650,N_6821);
and U7545 (N_7545,N_6813,N_6072);
nor U7546 (N_7546,N_6170,N_6623);
nand U7547 (N_7547,N_6054,N_6151);
nor U7548 (N_7548,N_6826,N_6494);
and U7549 (N_7549,N_6630,N_6285);
or U7550 (N_7550,N_6842,N_6035);
nor U7551 (N_7551,N_6925,N_6859);
xnor U7552 (N_7552,N_6362,N_6858);
and U7553 (N_7553,N_6408,N_6515);
or U7554 (N_7554,N_6266,N_6767);
nor U7555 (N_7555,N_6368,N_6900);
and U7556 (N_7556,N_6726,N_6974);
and U7557 (N_7557,N_6072,N_6756);
nand U7558 (N_7558,N_6602,N_6831);
nand U7559 (N_7559,N_6660,N_6120);
and U7560 (N_7560,N_6398,N_6079);
nor U7561 (N_7561,N_6917,N_6954);
and U7562 (N_7562,N_6487,N_6998);
nand U7563 (N_7563,N_6800,N_6324);
or U7564 (N_7564,N_6421,N_6218);
nand U7565 (N_7565,N_6479,N_6171);
and U7566 (N_7566,N_6366,N_6160);
nor U7567 (N_7567,N_6264,N_6950);
and U7568 (N_7568,N_6822,N_6352);
nand U7569 (N_7569,N_6454,N_6859);
and U7570 (N_7570,N_6325,N_6788);
and U7571 (N_7571,N_6118,N_6695);
nand U7572 (N_7572,N_6415,N_6298);
and U7573 (N_7573,N_6133,N_6125);
nor U7574 (N_7574,N_6094,N_6922);
and U7575 (N_7575,N_6075,N_6941);
or U7576 (N_7576,N_6582,N_6474);
or U7577 (N_7577,N_6832,N_6785);
nand U7578 (N_7578,N_6048,N_6059);
or U7579 (N_7579,N_6003,N_6673);
nor U7580 (N_7580,N_6483,N_6665);
or U7581 (N_7581,N_6381,N_6795);
xor U7582 (N_7582,N_6860,N_6934);
nand U7583 (N_7583,N_6367,N_6607);
nand U7584 (N_7584,N_6751,N_6859);
nor U7585 (N_7585,N_6194,N_6892);
nand U7586 (N_7586,N_6229,N_6621);
and U7587 (N_7587,N_6604,N_6372);
or U7588 (N_7588,N_6431,N_6380);
and U7589 (N_7589,N_6475,N_6608);
and U7590 (N_7590,N_6598,N_6162);
and U7591 (N_7591,N_6010,N_6603);
nand U7592 (N_7592,N_6563,N_6316);
nand U7593 (N_7593,N_6270,N_6623);
or U7594 (N_7594,N_6905,N_6821);
or U7595 (N_7595,N_6225,N_6182);
or U7596 (N_7596,N_6506,N_6286);
xnor U7597 (N_7597,N_6145,N_6070);
or U7598 (N_7598,N_6488,N_6197);
and U7599 (N_7599,N_6965,N_6869);
and U7600 (N_7600,N_6630,N_6200);
nand U7601 (N_7601,N_6366,N_6721);
or U7602 (N_7602,N_6023,N_6727);
nand U7603 (N_7603,N_6090,N_6647);
nor U7604 (N_7604,N_6206,N_6431);
and U7605 (N_7605,N_6152,N_6817);
or U7606 (N_7606,N_6612,N_6708);
nand U7607 (N_7607,N_6506,N_6343);
nand U7608 (N_7608,N_6412,N_6372);
nand U7609 (N_7609,N_6612,N_6992);
nor U7610 (N_7610,N_6440,N_6625);
nand U7611 (N_7611,N_6304,N_6717);
and U7612 (N_7612,N_6152,N_6169);
and U7613 (N_7613,N_6501,N_6965);
nand U7614 (N_7614,N_6766,N_6822);
nor U7615 (N_7615,N_6810,N_6771);
nand U7616 (N_7616,N_6878,N_6902);
nand U7617 (N_7617,N_6506,N_6479);
and U7618 (N_7618,N_6297,N_6088);
nand U7619 (N_7619,N_6668,N_6556);
nor U7620 (N_7620,N_6720,N_6287);
nand U7621 (N_7621,N_6107,N_6300);
xor U7622 (N_7622,N_6876,N_6765);
and U7623 (N_7623,N_6727,N_6789);
nor U7624 (N_7624,N_6668,N_6549);
nand U7625 (N_7625,N_6741,N_6627);
and U7626 (N_7626,N_6616,N_6864);
nor U7627 (N_7627,N_6833,N_6617);
or U7628 (N_7628,N_6893,N_6642);
nand U7629 (N_7629,N_6269,N_6155);
and U7630 (N_7630,N_6949,N_6213);
and U7631 (N_7631,N_6389,N_6904);
or U7632 (N_7632,N_6792,N_6819);
and U7633 (N_7633,N_6457,N_6439);
and U7634 (N_7634,N_6671,N_6639);
nor U7635 (N_7635,N_6372,N_6934);
or U7636 (N_7636,N_6839,N_6236);
and U7637 (N_7637,N_6820,N_6654);
nor U7638 (N_7638,N_6035,N_6141);
nand U7639 (N_7639,N_6082,N_6513);
or U7640 (N_7640,N_6931,N_6738);
nor U7641 (N_7641,N_6439,N_6281);
nand U7642 (N_7642,N_6028,N_6590);
xor U7643 (N_7643,N_6820,N_6050);
or U7644 (N_7644,N_6750,N_6200);
nand U7645 (N_7645,N_6384,N_6670);
nand U7646 (N_7646,N_6491,N_6435);
and U7647 (N_7647,N_6906,N_6347);
and U7648 (N_7648,N_6106,N_6173);
or U7649 (N_7649,N_6937,N_6774);
and U7650 (N_7650,N_6460,N_6828);
and U7651 (N_7651,N_6049,N_6635);
and U7652 (N_7652,N_6580,N_6582);
and U7653 (N_7653,N_6854,N_6145);
and U7654 (N_7654,N_6576,N_6514);
or U7655 (N_7655,N_6029,N_6667);
or U7656 (N_7656,N_6681,N_6180);
nand U7657 (N_7657,N_6480,N_6939);
and U7658 (N_7658,N_6930,N_6955);
nand U7659 (N_7659,N_6047,N_6391);
nor U7660 (N_7660,N_6166,N_6854);
and U7661 (N_7661,N_6051,N_6974);
or U7662 (N_7662,N_6374,N_6558);
nand U7663 (N_7663,N_6908,N_6622);
or U7664 (N_7664,N_6463,N_6716);
nor U7665 (N_7665,N_6292,N_6989);
nand U7666 (N_7666,N_6862,N_6167);
or U7667 (N_7667,N_6719,N_6781);
nor U7668 (N_7668,N_6628,N_6451);
xor U7669 (N_7669,N_6589,N_6905);
nor U7670 (N_7670,N_6139,N_6574);
and U7671 (N_7671,N_6088,N_6374);
or U7672 (N_7672,N_6244,N_6895);
or U7673 (N_7673,N_6551,N_6501);
and U7674 (N_7674,N_6683,N_6785);
nor U7675 (N_7675,N_6536,N_6133);
or U7676 (N_7676,N_6089,N_6218);
and U7677 (N_7677,N_6687,N_6286);
or U7678 (N_7678,N_6308,N_6570);
nor U7679 (N_7679,N_6289,N_6570);
and U7680 (N_7680,N_6636,N_6590);
and U7681 (N_7681,N_6556,N_6023);
or U7682 (N_7682,N_6783,N_6120);
nand U7683 (N_7683,N_6672,N_6460);
and U7684 (N_7684,N_6536,N_6128);
or U7685 (N_7685,N_6995,N_6686);
or U7686 (N_7686,N_6829,N_6660);
or U7687 (N_7687,N_6872,N_6999);
or U7688 (N_7688,N_6638,N_6677);
nor U7689 (N_7689,N_6859,N_6020);
xnor U7690 (N_7690,N_6269,N_6708);
or U7691 (N_7691,N_6121,N_6851);
or U7692 (N_7692,N_6399,N_6740);
nor U7693 (N_7693,N_6269,N_6399);
or U7694 (N_7694,N_6430,N_6985);
and U7695 (N_7695,N_6624,N_6809);
or U7696 (N_7696,N_6745,N_6154);
and U7697 (N_7697,N_6869,N_6853);
or U7698 (N_7698,N_6219,N_6889);
or U7699 (N_7699,N_6056,N_6893);
and U7700 (N_7700,N_6956,N_6577);
nor U7701 (N_7701,N_6928,N_6180);
or U7702 (N_7702,N_6703,N_6369);
nand U7703 (N_7703,N_6253,N_6258);
nor U7704 (N_7704,N_6658,N_6097);
nor U7705 (N_7705,N_6898,N_6882);
and U7706 (N_7706,N_6702,N_6790);
and U7707 (N_7707,N_6024,N_6909);
and U7708 (N_7708,N_6845,N_6269);
or U7709 (N_7709,N_6433,N_6545);
and U7710 (N_7710,N_6066,N_6590);
nand U7711 (N_7711,N_6127,N_6200);
and U7712 (N_7712,N_6640,N_6012);
and U7713 (N_7713,N_6140,N_6373);
nand U7714 (N_7714,N_6217,N_6577);
nor U7715 (N_7715,N_6154,N_6015);
nand U7716 (N_7716,N_6151,N_6897);
or U7717 (N_7717,N_6833,N_6487);
nand U7718 (N_7718,N_6914,N_6143);
nand U7719 (N_7719,N_6541,N_6755);
or U7720 (N_7720,N_6014,N_6111);
xor U7721 (N_7721,N_6749,N_6997);
or U7722 (N_7722,N_6381,N_6873);
or U7723 (N_7723,N_6091,N_6801);
nand U7724 (N_7724,N_6503,N_6728);
nor U7725 (N_7725,N_6757,N_6804);
nand U7726 (N_7726,N_6805,N_6918);
nor U7727 (N_7727,N_6082,N_6695);
and U7728 (N_7728,N_6995,N_6343);
and U7729 (N_7729,N_6917,N_6433);
nor U7730 (N_7730,N_6037,N_6546);
nor U7731 (N_7731,N_6423,N_6833);
or U7732 (N_7732,N_6038,N_6883);
nand U7733 (N_7733,N_6015,N_6803);
nor U7734 (N_7734,N_6199,N_6191);
and U7735 (N_7735,N_6712,N_6188);
and U7736 (N_7736,N_6341,N_6687);
and U7737 (N_7737,N_6162,N_6621);
and U7738 (N_7738,N_6911,N_6527);
or U7739 (N_7739,N_6238,N_6913);
nor U7740 (N_7740,N_6169,N_6575);
nor U7741 (N_7741,N_6308,N_6507);
and U7742 (N_7742,N_6832,N_6181);
nand U7743 (N_7743,N_6648,N_6660);
and U7744 (N_7744,N_6390,N_6727);
nor U7745 (N_7745,N_6191,N_6616);
and U7746 (N_7746,N_6904,N_6844);
or U7747 (N_7747,N_6249,N_6212);
nand U7748 (N_7748,N_6041,N_6165);
and U7749 (N_7749,N_6667,N_6884);
nor U7750 (N_7750,N_6111,N_6952);
nor U7751 (N_7751,N_6217,N_6392);
nor U7752 (N_7752,N_6646,N_6004);
nand U7753 (N_7753,N_6214,N_6601);
or U7754 (N_7754,N_6323,N_6408);
nor U7755 (N_7755,N_6018,N_6832);
or U7756 (N_7756,N_6221,N_6376);
nand U7757 (N_7757,N_6137,N_6787);
and U7758 (N_7758,N_6798,N_6764);
or U7759 (N_7759,N_6330,N_6808);
nor U7760 (N_7760,N_6947,N_6263);
or U7761 (N_7761,N_6465,N_6413);
and U7762 (N_7762,N_6643,N_6061);
and U7763 (N_7763,N_6318,N_6062);
or U7764 (N_7764,N_6662,N_6486);
nand U7765 (N_7765,N_6331,N_6808);
and U7766 (N_7766,N_6406,N_6814);
nand U7767 (N_7767,N_6101,N_6652);
and U7768 (N_7768,N_6788,N_6407);
and U7769 (N_7769,N_6115,N_6615);
and U7770 (N_7770,N_6634,N_6766);
nand U7771 (N_7771,N_6179,N_6056);
or U7772 (N_7772,N_6135,N_6946);
xnor U7773 (N_7773,N_6075,N_6304);
and U7774 (N_7774,N_6493,N_6386);
or U7775 (N_7775,N_6932,N_6599);
or U7776 (N_7776,N_6677,N_6078);
and U7777 (N_7777,N_6449,N_6216);
nand U7778 (N_7778,N_6486,N_6122);
nor U7779 (N_7779,N_6165,N_6986);
nand U7780 (N_7780,N_6595,N_6804);
or U7781 (N_7781,N_6548,N_6139);
nand U7782 (N_7782,N_6269,N_6350);
or U7783 (N_7783,N_6265,N_6723);
nand U7784 (N_7784,N_6583,N_6653);
or U7785 (N_7785,N_6577,N_6711);
nor U7786 (N_7786,N_6571,N_6059);
and U7787 (N_7787,N_6833,N_6524);
or U7788 (N_7788,N_6651,N_6646);
nor U7789 (N_7789,N_6092,N_6157);
xnor U7790 (N_7790,N_6406,N_6381);
and U7791 (N_7791,N_6769,N_6279);
nand U7792 (N_7792,N_6170,N_6611);
nand U7793 (N_7793,N_6673,N_6689);
or U7794 (N_7794,N_6219,N_6875);
nor U7795 (N_7795,N_6576,N_6030);
and U7796 (N_7796,N_6249,N_6855);
nand U7797 (N_7797,N_6456,N_6445);
and U7798 (N_7798,N_6920,N_6675);
or U7799 (N_7799,N_6371,N_6255);
and U7800 (N_7800,N_6471,N_6060);
and U7801 (N_7801,N_6745,N_6372);
and U7802 (N_7802,N_6660,N_6220);
nor U7803 (N_7803,N_6847,N_6785);
or U7804 (N_7804,N_6880,N_6758);
or U7805 (N_7805,N_6415,N_6493);
or U7806 (N_7806,N_6182,N_6679);
nand U7807 (N_7807,N_6738,N_6138);
and U7808 (N_7808,N_6983,N_6686);
nand U7809 (N_7809,N_6525,N_6902);
nand U7810 (N_7810,N_6337,N_6940);
nand U7811 (N_7811,N_6411,N_6197);
xnor U7812 (N_7812,N_6307,N_6584);
or U7813 (N_7813,N_6551,N_6882);
nor U7814 (N_7814,N_6290,N_6237);
or U7815 (N_7815,N_6425,N_6776);
nand U7816 (N_7816,N_6693,N_6812);
or U7817 (N_7817,N_6571,N_6511);
nand U7818 (N_7818,N_6461,N_6488);
and U7819 (N_7819,N_6376,N_6749);
nand U7820 (N_7820,N_6477,N_6114);
and U7821 (N_7821,N_6391,N_6779);
or U7822 (N_7822,N_6661,N_6167);
nor U7823 (N_7823,N_6728,N_6436);
and U7824 (N_7824,N_6310,N_6509);
nor U7825 (N_7825,N_6278,N_6862);
nor U7826 (N_7826,N_6404,N_6682);
nand U7827 (N_7827,N_6241,N_6938);
nor U7828 (N_7828,N_6018,N_6176);
nand U7829 (N_7829,N_6235,N_6290);
or U7830 (N_7830,N_6646,N_6437);
or U7831 (N_7831,N_6779,N_6974);
nand U7832 (N_7832,N_6796,N_6301);
nand U7833 (N_7833,N_6421,N_6323);
and U7834 (N_7834,N_6905,N_6226);
or U7835 (N_7835,N_6548,N_6146);
xnor U7836 (N_7836,N_6185,N_6807);
nor U7837 (N_7837,N_6585,N_6266);
and U7838 (N_7838,N_6148,N_6093);
and U7839 (N_7839,N_6802,N_6590);
or U7840 (N_7840,N_6113,N_6159);
nor U7841 (N_7841,N_6145,N_6835);
nand U7842 (N_7842,N_6028,N_6079);
and U7843 (N_7843,N_6155,N_6771);
or U7844 (N_7844,N_6606,N_6239);
nor U7845 (N_7845,N_6530,N_6254);
xnor U7846 (N_7846,N_6877,N_6083);
nor U7847 (N_7847,N_6600,N_6605);
nand U7848 (N_7848,N_6734,N_6610);
and U7849 (N_7849,N_6367,N_6708);
and U7850 (N_7850,N_6281,N_6605);
nor U7851 (N_7851,N_6498,N_6377);
nor U7852 (N_7852,N_6138,N_6397);
nor U7853 (N_7853,N_6456,N_6724);
nand U7854 (N_7854,N_6384,N_6457);
nor U7855 (N_7855,N_6869,N_6944);
and U7856 (N_7856,N_6698,N_6614);
nor U7857 (N_7857,N_6747,N_6220);
and U7858 (N_7858,N_6486,N_6181);
and U7859 (N_7859,N_6881,N_6363);
nand U7860 (N_7860,N_6419,N_6117);
nand U7861 (N_7861,N_6233,N_6918);
and U7862 (N_7862,N_6368,N_6794);
nand U7863 (N_7863,N_6092,N_6889);
nor U7864 (N_7864,N_6010,N_6651);
and U7865 (N_7865,N_6993,N_6115);
nor U7866 (N_7866,N_6108,N_6809);
and U7867 (N_7867,N_6634,N_6536);
xnor U7868 (N_7868,N_6293,N_6403);
nand U7869 (N_7869,N_6094,N_6144);
or U7870 (N_7870,N_6246,N_6508);
and U7871 (N_7871,N_6850,N_6591);
and U7872 (N_7872,N_6682,N_6634);
and U7873 (N_7873,N_6443,N_6172);
nand U7874 (N_7874,N_6718,N_6181);
or U7875 (N_7875,N_6590,N_6035);
and U7876 (N_7876,N_6336,N_6858);
nand U7877 (N_7877,N_6651,N_6179);
nand U7878 (N_7878,N_6790,N_6533);
nand U7879 (N_7879,N_6137,N_6942);
and U7880 (N_7880,N_6180,N_6517);
and U7881 (N_7881,N_6526,N_6146);
and U7882 (N_7882,N_6965,N_6215);
or U7883 (N_7883,N_6103,N_6001);
nand U7884 (N_7884,N_6004,N_6154);
and U7885 (N_7885,N_6376,N_6414);
nand U7886 (N_7886,N_6922,N_6133);
and U7887 (N_7887,N_6004,N_6207);
nor U7888 (N_7888,N_6404,N_6551);
nand U7889 (N_7889,N_6410,N_6781);
nor U7890 (N_7890,N_6418,N_6142);
or U7891 (N_7891,N_6309,N_6816);
nor U7892 (N_7892,N_6802,N_6709);
nor U7893 (N_7893,N_6588,N_6388);
or U7894 (N_7894,N_6466,N_6048);
nor U7895 (N_7895,N_6215,N_6615);
and U7896 (N_7896,N_6909,N_6348);
nand U7897 (N_7897,N_6580,N_6370);
nor U7898 (N_7898,N_6129,N_6709);
nor U7899 (N_7899,N_6920,N_6607);
nand U7900 (N_7900,N_6738,N_6395);
nand U7901 (N_7901,N_6702,N_6131);
or U7902 (N_7902,N_6564,N_6401);
and U7903 (N_7903,N_6839,N_6800);
nand U7904 (N_7904,N_6366,N_6889);
and U7905 (N_7905,N_6169,N_6736);
and U7906 (N_7906,N_6980,N_6516);
or U7907 (N_7907,N_6901,N_6285);
nor U7908 (N_7908,N_6466,N_6843);
nand U7909 (N_7909,N_6449,N_6808);
and U7910 (N_7910,N_6957,N_6484);
nand U7911 (N_7911,N_6249,N_6142);
nor U7912 (N_7912,N_6342,N_6841);
nor U7913 (N_7913,N_6130,N_6540);
and U7914 (N_7914,N_6126,N_6321);
xnor U7915 (N_7915,N_6849,N_6666);
or U7916 (N_7916,N_6846,N_6345);
nand U7917 (N_7917,N_6537,N_6777);
and U7918 (N_7918,N_6768,N_6550);
nand U7919 (N_7919,N_6565,N_6406);
and U7920 (N_7920,N_6580,N_6033);
nor U7921 (N_7921,N_6021,N_6141);
or U7922 (N_7922,N_6578,N_6562);
or U7923 (N_7923,N_6646,N_6973);
nor U7924 (N_7924,N_6953,N_6529);
or U7925 (N_7925,N_6727,N_6307);
nor U7926 (N_7926,N_6361,N_6639);
nand U7927 (N_7927,N_6277,N_6164);
nand U7928 (N_7928,N_6210,N_6664);
nor U7929 (N_7929,N_6595,N_6628);
nand U7930 (N_7930,N_6660,N_6215);
or U7931 (N_7931,N_6799,N_6894);
and U7932 (N_7932,N_6436,N_6312);
or U7933 (N_7933,N_6825,N_6577);
or U7934 (N_7934,N_6675,N_6179);
or U7935 (N_7935,N_6369,N_6530);
nand U7936 (N_7936,N_6970,N_6082);
nand U7937 (N_7937,N_6818,N_6830);
nor U7938 (N_7938,N_6477,N_6134);
and U7939 (N_7939,N_6999,N_6551);
or U7940 (N_7940,N_6432,N_6895);
nor U7941 (N_7941,N_6179,N_6934);
and U7942 (N_7942,N_6108,N_6597);
nand U7943 (N_7943,N_6005,N_6102);
or U7944 (N_7944,N_6778,N_6832);
nand U7945 (N_7945,N_6277,N_6279);
or U7946 (N_7946,N_6628,N_6224);
and U7947 (N_7947,N_6132,N_6933);
xor U7948 (N_7948,N_6872,N_6750);
and U7949 (N_7949,N_6157,N_6196);
or U7950 (N_7950,N_6420,N_6361);
nand U7951 (N_7951,N_6713,N_6256);
or U7952 (N_7952,N_6403,N_6348);
nand U7953 (N_7953,N_6027,N_6457);
and U7954 (N_7954,N_6813,N_6058);
and U7955 (N_7955,N_6756,N_6941);
nand U7956 (N_7956,N_6940,N_6528);
nor U7957 (N_7957,N_6410,N_6599);
nor U7958 (N_7958,N_6011,N_6021);
and U7959 (N_7959,N_6533,N_6361);
nand U7960 (N_7960,N_6535,N_6066);
and U7961 (N_7961,N_6168,N_6863);
nand U7962 (N_7962,N_6173,N_6930);
nand U7963 (N_7963,N_6644,N_6517);
nor U7964 (N_7964,N_6568,N_6736);
nor U7965 (N_7965,N_6580,N_6170);
or U7966 (N_7966,N_6205,N_6195);
xor U7967 (N_7967,N_6410,N_6334);
nand U7968 (N_7968,N_6577,N_6753);
nand U7969 (N_7969,N_6998,N_6024);
and U7970 (N_7970,N_6529,N_6413);
and U7971 (N_7971,N_6851,N_6651);
nor U7972 (N_7972,N_6734,N_6137);
nor U7973 (N_7973,N_6841,N_6873);
or U7974 (N_7974,N_6715,N_6208);
nor U7975 (N_7975,N_6428,N_6108);
or U7976 (N_7976,N_6637,N_6936);
xnor U7977 (N_7977,N_6874,N_6190);
and U7978 (N_7978,N_6343,N_6201);
and U7979 (N_7979,N_6085,N_6065);
nand U7980 (N_7980,N_6077,N_6753);
nand U7981 (N_7981,N_6927,N_6266);
nor U7982 (N_7982,N_6820,N_6699);
nor U7983 (N_7983,N_6363,N_6441);
or U7984 (N_7984,N_6494,N_6383);
nand U7985 (N_7985,N_6633,N_6796);
nor U7986 (N_7986,N_6374,N_6470);
or U7987 (N_7987,N_6296,N_6038);
nand U7988 (N_7988,N_6700,N_6190);
and U7989 (N_7989,N_6777,N_6261);
nand U7990 (N_7990,N_6658,N_6682);
and U7991 (N_7991,N_6325,N_6965);
xnor U7992 (N_7992,N_6191,N_6749);
nor U7993 (N_7993,N_6920,N_6159);
and U7994 (N_7994,N_6349,N_6158);
or U7995 (N_7995,N_6068,N_6332);
nor U7996 (N_7996,N_6410,N_6791);
nor U7997 (N_7997,N_6761,N_6830);
nor U7998 (N_7998,N_6059,N_6292);
and U7999 (N_7999,N_6457,N_6935);
nor U8000 (N_8000,N_7621,N_7216);
nand U8001 (N_8001,N_7335,N_7030);
and U8002 (N_8002,N_7154,N_7541);
nor U8003 (N_8003,N_7495,N_7913);
or U8004 (N_8004,N_7288,N_7822);
nor U8005 (N_8005,N_7098,N_7857);
and U8006 (N_8006,N_7411,N_7380);
nand U8007 (N_8007,N_7117,N_7743);
or U8008 (N_8008,N_7974,N_7150);
nand U8009 (N_8009,N_7929,N_7761);
or U8010 (N_8010,N_7844,N_7052);
nand U8011 (N_8011,N_7053,N_7181);
xnor U8012 (N_8012,N_7206,N_7125);
and U8013 (N_8013,N_7609,N_7666);
or U8014 (N_8014,N_7491,N_7373);
or U8015 (N_8015,N_7207,N_7866);
nand U8016 (N_8016,N_7975,N_7047);
nor U8017 (N_8017,N_7337,N_7029);
nor U8018 (N_8018,N_7391,N_7210);
and U8019 (N_8019,N_7062,N_7064);
nor U8020 (N_8020,N_7983,N_7296);
nor U8021 (N_8021,N_7916,N_7838);
nor U8022 (N_8022,N_7370,N_7235);
nand U8023 (N_8023,N_7338,N_7504);
nor U8024 (N_8024,N_7189,N_7744);
nor U8025 (N_8025,N_7539,N_7617);
or U8026 (N_8026,N_7396,N_7148);
nand U8027 (N_8027,N_7453,N_7478);
and U8028 (N_8028,N_7114,N_7177);
or U8029 (N_8029,N_7323,N_7341);
nor U8030 (N_8030,N_7737,N_7771);
nor U8031 (N_8031,N_7674,N_7871);
and U8032 (N_8032,N_7054,N_7729);
xnor U8033 (N_8033,N_7951,N_7861);
nand U8034 (N_8034,N_7694,N_7420);
xor U8035 (N_8035,N_7646,N_7108);
nor U8036 (N_8036,N_7863,N_7889);
nand U8037 (N_8037,N_7229,N_7718);
and U8038 (N_8038,N_7026,N_7332);
nor U8039 (N_8039,N_7434,N_7078);
nor U8040 (N_8040,N_7712,N_7074);
or U8041 (N_8041,N_7497,N_7309);
and U8042 (N_8042,N_7225,N_7215);
or U8043 (N_8043,N_7707,N_7877);
nand U8044 (N_8044,N_7019,N_7873);
and U8045 (N_8045,N_7874,N_7915);
nand U8046 (N_8046,N_7232,N_7616);
nor U8047 (N_8047,N_7456,N_7855);
or U8048 (N_8048,N_7615,N_7265);
and U8049 (N_8049,N_7261,N_7551);
nor U8050 (N_8050,N_7101,N_7727);
or U8051 (N_8051,N_7113,N_7318);
or U8052 (N_8052,N_7233,N_7825);
nor U8053 (N_8053,N_7776,N_7998);
and U8054 (N_8054,N_7398,N_7284);
or U8055 (N_8055,N_7024,N_7275);
nor U8056 (N_8056,N_7255,N_7662);
nor U8057 (N_8057,N_7685,N_7700);
and U8058 (N_8058,N_7957,N_7543);
xor U8059 (N_8059,N_7953,N_7118);
and U8060 (N_8060,N_7741,N_7775);
and U8061 (N_8061,N_7642,N_7413);
nand U8062 (N_8062,N_7433,N_7440);
nand U8063 (N_8063,N_7553,N_7564);
nor U8064 (N_8064,N_7194,N_7003);
and U8065 (N_8065,N_7509,N_7481);
nor U8066 (N_8066,N_7529,N_7138);
and U8067 (N_8067,N_7698,N_7010);
or U8068 (N_8068,N_7182,N_7750);
nor U8069 (N_8069,N_7578,N_7445);
nor U8070 (N_8070,N_7406,N_7800);
nand U8071 (N_8071,N_7720,N_7832);
or U8072 (N_8072,N_7381,N_7186);
nor U8073 (N_8073,N_7902,N_7333);
nand U8074 (N_8074,N_7152,N_7277);
nand U8075 (N_8075,N_7936,N_7937);
nand U8076 (N_8076,N_7886,N_7670);
nand U8077 (N_8077,N_7093,N_7124);
and U8078 (N_8078,N_7013,N_7912);
or U8079 (N_8079,N_7887,N_7172);
or U8080 (N_8080,N_7379,N_7076);
and U8081 (N_8081,N_7583,N_7753);
nor U8082 (N_8082,N_7585,N_7828);
nor U8083 (N_8083,N_7127,N_7544);
nand U8084 (N_8084,N_7486,N_7352);
or U8085 (N_8085,N_7414,N_7268);
xnor U8086 (N_8086,N_7867,N_7677);
or U8087 (N_8087,N_7831,N_7371);
nor U8088 (N_8088,N_7151,N_7608);
and U8089 (N_8089,N_7409,N_7360);
nor U8090 (N_8090,N_7970,N_7365);
and U8091 (N_8091,N_7952,N_7386);
xor U8092 (N_8092,N_7724,N_7930);
or U8093 (N_8093,N_7244,N_7258);
nand U8094 (N_8094,N_7789,N_7967);
nand U8095 (N_8095,N_7826,N_7900);
nor U8096 (N_8096,N_7623,N_7682);
and U8097 (N_8097,N_7584,N_7131);
and U8098 (N_8098,N_7656,N_7441);
or U8099 (N_8099,N_7343,N_7159);
or U8100 (N_8100,N_7068,N_7103);
nand U8101 (N_8101,N_7102,N_7267);
nand U8102 (N_8102,N_7175,N_7600);
nor U8103 (N_8103,N_7959,N_7762);
nor U8104 (N_8104,N_7071,N_7725);
and U8105 (N_8105,N_7756,N_7701);
nor U8106 (N_8106,N_7419,N_7683);
nand U8107 (N_8107,N_7565,N_7249);
nor U8108 (N_8108,N_7031,N_7870);
nand U8109 (N_8109,N_7574,N_7279);
nor U8110 (N_8110,N_7452,N_7395);
or U8111 (N_8111,N_7226,N_7895);
or U8112 (N_8112,N_7596,N_7254);
or U8113 (N_8113,N_7001,N_7634);
and U8114 (N_8114,N_7465,N_7447);
nor U8115 (N_8115,N_7763,N_7805);
and U8116 (N_8116,N_7639,N_7483);
or U8117 (N_8117,N_7179,N_7988);
and U8118 (N_8118,N_7307,N_7095);
or U8119 (N_8119,N_7143,N_7963);
nand U8120 (N_8120,N_7271,N_7176);
nor U8121 (N_8121,N_7824,N_7620);
nor U8122 (N_8122,N_7752,N_7555);
nand U8123 (N_8123,N_7270,N_7035);
and U8124 (N_8124,N_7853,N_7740);
nor U8125 (N_8125,N_7810,N_7348);
and U8126 (N_8126,N_7790,N_7573);
xor U8127 (N_8127,N_7430,N_7164);
and U8128 (N_8128,N_7330,N_7292);
and U8129 (N_8129,N_7291,N_7947);
nand U8130 (N_8130,N_7846,N_7556);
nor U8131 (N_8131,N_7462,N_7550);
nand U8132 (N_8132,N_7667,N_7697);
and U8133 (N_8133,N_7022,N_7444);
nor U8134 (N_8134,N_7868,N_7845);
nor U8135 (N_8135,N_7392,N_7474);
nand U8136 (N_8136,N_7663,N_7829);
or U8137 (N_8137,N_7911,N_7436);
and U8138 (N_8138,N_7507,N_7067);
and U8139 (N_8139,N_7702,N_7094);
or U8140 (N_8140,N_7965,N_7402);
or U8141 (N_8141,N_7416,N_7467);
and U8142 (N_8142,N_7384,N_7817);
nor U8143 (N_8143,N_7922,N_7709);
nand U8144 (N_8144,N_7269,N_7532);
and U8145 (N_8145,N_7180,N_7032);
or U8146 (N_8146,N_7298,N_7213);
or U8147 (N_8147,N_7178,N_7905);
and U8148 (N_8148,N_7304,N_7714);
nand U8149 (N_8149,N_7759,N_7320);
nand U8150 (N_8150,N_7498,N_7185);
or U8151 (N_8151,N_7121,N_7948);
nand U8152 (N_8152,N_7859,N_7297);
nand U8153 (N_8153,N_7579,N_7387);
or U8154 (N_8154,N_7356,N_7769);
and U8155 (N_8155,N_7144,N_7107);
or U8156 (N_8156,N_7605,N_7891);
and U8157 (N_8157,N_7517,N_7624);
xor U8158 (N_8158,N_7722,N_7588);
nor U8159 (N_8159,N_7376,N_7918);
nand U8160 (N_8160,N_7766,N_7306);
and U8161 (N_8161,N_7319,N_7253);
and U8162 (N_8162,N_7777,N_7042);
or U8163 (N_8163,N_7116,N_7212);
nand U8164 (N_8164,N_7571,N_7612);
nor U8165 (N_8165,N_7650,N_7316);
nand U8166 (N_8166,N_7326,N_7548);
or U8167 (N_8167,N_7183,N_7807);
nand U8168 (N_8168,N_7500,N_7536);
and U8169 (N_8169,N_7699,N_7665);
or U8170 (N_8170,N_7086,N_7986);
nor U8171 (N_8171,N_7346,N_7136);
and U8172 (N_8172,N_7184,N_7781);
and U8173 (N_8173,N_7835,N_7765);
and U8174 (N_8174,N_7515,N_7328);
nand U8175 (N_8175,N_7793,N_7243);
and U8176 (N_8176,N_7405,N_7601);
and U8177 (N_8177,N_7802,N_7490);
nand U8178 (N_8178,N_7485,N_7821);
nand U8179 (N_8179,N_7115,N_7366);
or U8180 (N_8180,N_7072,N_7980);
or U8181 (N_8181,N_7191,N_7954);
nor U8182 (N_8182,N_7083,N_7520);
and U8183 (N_8183,N_7657,N_7885);
nand U8184 (N_8184,N_7518,N_7009);
and U8185 (N_8185,N_7850,N_7484);
and U8186 (N_8186,N_7836,N_7494);
xnor U8187 (N_8187,N_7973,N_7170);
nor U8188 (N_8188,N_7208,N_7716);
nor U8189 (N_8189,N_7531,N_7157);
and U8190 (N_8190,N_7214,N_7008);
nor U8191 (N_8191,N_7197,N_7303);
or U8192 (N_8192,N_7492,N_7424);
nor U8193 (N_8193,N_7129,N_7378);
nor U8194 (N_8194,N_7349,N_7968);
nand U8195 (N_8195,N_7946,N_7259);
nor U8196 (N_8196,N_7519,N_7188);
or U8197 (N_8197,N_7941,N_7917);
and U8198 (N_8198,N_7751,N_7687);
nor U8199 (N_8199,N_7914,N_7849);
and U8200 (N_8200,N_7016,N_7659);
nand U8201 (N_8201,N_7603,N_7069);
or U8202 (N_8202,N_7399,N_7390);
and U8203 (N_8203,N_7950,N_7311);
or U8204 (N_8204,N_7691,N_7407);
or U8205 (N_8205,N_7192,N_7437);
and U8206 (N_8206,N_7927,N_7971);
nand U8207 (N_8207,N_7881,N_7949);
and U8208 (N_8208,N_7245,N_7460);
nor U8209 (N_8209,N_7506,N_7535);
or U8210 (N_8210,N_7020,N_7589);
and U8211 (N_8211,N_7527,N_7339);
nand U8212 (N_8212,N_7449,N_7542);
nand U8213 (N_8213,N_7158,N_7290);
nor U8214 (N_8214,N_7894,N_7732);
and U8215 (N_8215,N_7048,N_7163);
and U8216 (N_8216,N_7648,N_7742);
or U8217 (N_8217,N_7593,N_7363);
nor U8218 (N_8218,N_7372,N_7595);
or U8219 (N_8219,N_7782,N_7477);
nand U8220 (N_8220,N_7223,N_7066);
nor U8221 (N_8221,N_7109,N_7679);
nor U8222 (N_8222,N_7241,N_7140);
or U8223 (N_8223,N_7325,N_7770);
and U8224 (N_8224,N_7631,N_7045);
and U8225 (N_8225,N_7193,N_7299);
nand U8226 (N_8226,N_7160,N_7547);
or U8227 (N_8227,N_7510,N_7077);
and U8228 (N_8228,N_7196,N_7156);
or U8229 (N_8229,N_7100,N_7302);
or U8230 (N_8230,N_7021,N_7023);
or U8231 (N_8231,N_7374,N_7499);
or U8232 (N_8232,N_7669,N_7979);
or U8233 (N_8233,N_7658,N_7684);
nor U8234 (N_8234,N_7635,N_7926);
nor U8235 (N_8235,N_7856,N_7622);
nand U8236 (N_8236,N_7592,N_7317);
and U8237 (N_8237,N_7190,N_7931);
and U8238 (N_8238,N_7237,N_7672);
or U8239 (N_8239,N_7962,N_7221);
and U8240 (N_8240,N_7784,N_7070);
and U8241 (N_8241,N_7613,N_7295);
nor U8242 (N_8242,N_7723,N_7678);
nand U8243 (N_8243,N_7576,N_7961);
nor U8244 (N_8244,N_7025,N_7393);
nand U8245 (N_8245,N_7928,N_7418);
nand U8246 (N_8246,N_7017,N_7038);
and U8247 (N_8247,N_7198,N_7883);
nor U8248 (N_8248,N_7664,N_7110);
nand U8249 (N_8249,N_7511,N_7065);
and U8250 (N_8250,N_7218,N_7713);
nor U8251 (N_8251,N_7690,N_7755);
and U8252 (N_8252,N_7878,N_7502);
nand U8253 (N_8253,N_7004,N_7458);
nand U8254 (N_8254,N_7734,N_7758);
or U8255 (N_8255,N_7530,N_7869);
nand U8256 (N_8256,N_7731,N_7899);
nand U8257 (N_8257,N_7220,N_7310);
nand U8258 (N_8258,N_7106,N_7400);
or U8259 (N_8259,N_7155,N_7661);
or U8260 (N_8260,N_7966,N_7351);
nor U8261 (N_8261,N_7660,N_7939);
and U8262 (N_8262,N_7813,N_7359);
and U8263 (N_8263,N_7227,N_7513);
or U8264 (N_8264,N_7272,N_7626);
nor U8265 (N_8265,N_7875,N_7142);
nand U8266 (N_8266,N_7767,N_7860);
or U8267 (N_8267,N_7369,N_7091);
nor U8268 (N_8268,N_7431,N_7280);
nor U8269 (N_8269,N_7976,N_7528);
nor U8270 (N_8270,N_7276,N_7768);
nor U8271 (N_8271,N_7327,N_7563);
and U8272 (N_8272,N_7858,N_7429);
nor U8273 (N_8273,N_7345,N_7787);
or U8274 (N_8274,N_7778,N_7897);
nand U8275 (N_8275,N_7786,N_7834);
nor U8276 (N_8276,N_7710,N_7049);
and U8277 (N_8277,N_7128,N_7161);
and U8278 (N_8278,N_7361,N_7099);
nor U8279 (N_8279,N_7063,N_7201);
nand U8280 (N_8280,N_7808,N_7839);
nor U8281 (N_8281,N_7818,N_7422);
nor U8282 (N_8282,N_7676,N_7582);
and U8283 (N_8283,N_7638,N_7993);
nand U8284 (N_8284,N_7126,N_7693);
and U8285 (N_8285,N_7559,N_7643);
nor U8286 (N_8286,N_7721,N_7872);
nor U8287 (N_8287,N_7036,N_7096);
and U8288 (N_8288,N_7473,N_7843);
or U8289 (N_8289,N_7920,N_7283);
and U8290 (N_8290,N_7815,N_7014);
nand U8291 (N_8291,N_7606,N_7996);
nor U8292 (N_8292,N_7910,N_7903);
nor U8293 (N_8293,N_7746,N_7814);
or U8294 (N_8294,N_7503,N_7239);
nand U8295 (N_8295,N_7219,N_7749);
nor U8296 (N_8296,N_7262,N_7308);
or U8297 (N_8297,N_7516,N_7525);
or U8298 (N_8298,N_7594,N_7353);
and U8299 (N_8299,N_7681,N_7907);
xnor U8300 (N_8300,N_7133,N_7137);
nor U8301 (N_8301,N_7882,N_7044);
nor U8302 (N_8302,N_7586,N_7628);
nor U8303 (N_8303,N_7404,N_7377);
nand U8304 (N_8304,N_7222,N_7342);
nand U8305 (N_8305,N_7446,N_7251);
or U8306 (N_8306,N_7480,N_7978);
nor U8307 (N_8307,N_7908,N_7240);
nor U8308 (N_8308,N_7075,N_7748);
and U8309 (N_8309,N_7415,N_7892);
nor U8310 (N_8310,N_7566,N_7006);
or U8311 (N_8311,N_7149,N_7043);
or U8312 (N_8312,N_7165,N_7087);
or U8313 (N_8313,N_7058,N_7122);
and U8314 (N_8314,N_7614,N_7324);
nor U8315 (N_8315,N_7408,N_7388);
nor U8316 (N_8316,N_7994,N_7512);
nor U8317 (N_8317,N_7134,N_7633);
or U8318 (N_8318,N_7364,N_7848);
and U8319 (N_8319,N_7773,N_7037);
or U8320 (N_8320,N_7797,N_7427);
nand U8321 (N_8321,N_7457,N_7187);
nor U8322 (N_8322,N_7533,N_7321);
nand U8323 (N_8323,N_7654,N_7514);
nor U8324 (N_8324,N_7285,N_7455);
or U8325 (N_8325,N_7217,N_7286);
and U8326 (N_8326,N_7056,N_7312);
or U8327 (N_8327,N_7082,N_7464);
nand U8328 (N_8328,N_7730,N_7708);
nor U8329 (N_8329,N_7266,N_7675);
and U8330 (N_8330,N_7088,N_7935);
and U8331 (N_8331,N_7476,N_7479);
and U8332 (N_8332,N_7552,N_7774);
nand U8333 (N_8333,N_7619,N_7123);
or U8334 (N_8334,N_7211,N_7294);
nand U8335 (N_8335,N_7092,N_7879);
nor U8336 (N_8336,N_7987,N_7046);
nand U8337 (N_8337,N_7819,N_7538);
and U8338 (N_8338,N_7247,N_7119);
and U8339 (N_8339,N_7367,N_7577);
nand U8340 (N_8340,N_7314,N_7686);
and U8341 (N_8341,N_7558,N_7015);
nor U8342 (N_8342,N_7598,N_7000);
and U8343 (N_8343,N_7997,N_7554);
or U8344 (N_8344,N_7717,N_7924);
or U8345 (N_8345,N_7153,N_7442);
and U8346 (N_8346,N_7898,N_7146);
nand U8347 (N_8347,N_7322,N_7050);
nor U8348 (N_8348,N_7166,N_7147);
nor U8349 (N_8349,N_7696,N_7545);
nand U8350 (N_8350,N_7120,N_7085);
nor U8351 (N_8351,N_7745,N_7385);
nor U8352 (N_8352,N_7097,N_7073);
nor U8353 (N_8353,N_7162,N_7715);
and U8354 (N_8354,N_7537,N_7027);
and U8355 (N_8355,N_7599,N_7990);
nor U8356 (N_8356,N_7804,N_7890);
or U8357 (N_8357,N_7468,N_7007);
xor U8358 (N_8358,N_7984,N_7847);
nand U8359 (N_8359,N_7135,N_7471);
or U8360 (N_8360,N_7852,N_7803);
nand U8361 (N_8361,N_7199,N_7354);
or U8362 (N_8362,N_7355,N_7827);
and U8363 (N_8363,N_7801,N_7488);
nand U8364 (N_8364,N_7340,N_7806);
nor U8365 (N_8365,N_7647,N_7470);
or U8366 (N_8366,N_7637,N_7055);
and U8367 (N_8367,N_7991,N_7412);
or U8368 (N_8368,N_7602,N_7816);
nand U8369 (N_8369,N_7689,N_7876);
or U8370 (N_8370,N_7726,N_7234);
nor U8371 (N_8371,N_7489,N_7278);
nand U8372 (N_8372,N_7250,N_7644);
and U8373 (N_8373,N_7611,N_7228);
nand U8374 (N_8374,N_7522,N_7534);
and U8375 (N_8375,N_7041,N_7651);
nor U8376 (N_8376,N_7028,N_7587);
nand U8377 (N_8377,N_7747,N_7493);
xnor U8378 (N_8378,N_7933,N_7591);
or U8379 (N_8379,N_7671,N_7736);
or U8380 (N_8380,N_7200,N_7130);
nand U8381 (N_8381,N_7443,N_7012);
and U8382 (N_8382,N_7812,N_7925);
nor U8383 (N_8383,N_7132,N_7809);
and U8384 (N_8384,N_7772,N_7604);
nor U8385 (N_8385,N_7383,N_7864);
nand U8386 (N_8386,N_7139,N_7540);
nor U8387 (N_8387,N_7079,N_7051);
or U8388 (N_8388,N_7273,N_7459);
and U8389 (N_8389,N_7688,N_7842);
and U8390 (N_8390,N_7059,N_7425);
and U8391 (N_8391,N_7173,N_7830);
xnor U8392 (N_8392,N_7618,N_7331);
nand U8393 (N_8393,N_7673,N_7081);
nand U8394 (N_8394,N_7263,N_7854);
and U8395 (N_8395,N_7796,N_7033);
or U8396 (N_8396,N_7719,N_7649);
and U8397 (N_8397,N_7305,N_7002);
and U8398 (N_8398,N_7989,N_7630);
xor U8399 (N_8399,N_7347,N_7627);
nand U8400 (N_8400,N_7111,N_7487);
nand U8401 (N_8401,N_7865,N_7590);
or U8402 (N_8402,N_7260,N_7706);
or U8403 (N_8403,N_7421,N_7287);
xnor U8404 (N_8404,N_7840,N_7168);
nand U8405 (N_8405,N_7203,N_7981);
and U8406 (N_8406,N_7549,N_7389);
and U8407 (N_8407,N_7329,N_7692);
or U8408 (N_8408,N_7909,N_7906);
nand U8409 (N_8409,N_7641,N_7569);
nand U8410 (N_8410,N_7851,N_7655);
and U8411 (N_8411,N_7972,N_7705);
nand U8412 (N_8412,N_7760,N_7735);
nor U8413 (N_8413,N_7368,N_7791);
and U8414 (N_8414,N_7257,N_7080);
or U8415 (N_8415,N_7224,N_7728);
or U8416 (N_8416,N_7944,N_7580);
xor U8417 (N_8417,N_7739,N_7607);
nand U8418 (N_8418,N_7202,N_7561);
nand U8419 (N_8419,N_7293,N_7382);
and U8420 (N_8420,N_7252,N_7652);
or U8421 (N_8421,N_7209,N_7426);
nor U8422 (N_8422,N_7089,N_7238);
and U8423 (N_8423,N_7896,N_7526);
or U8424 (N_8424,N_7466,N_7105);
nand U8425 (N_8425,N_7837,N_7754);
and U8426 (N_8426,N_7375,N_7454);
and U8427 (N_8427,N_7904,N_7938);
nor U8428 (N_8428,N_7779,N_7448);
nor U8429 (N_8429,N_7572,N_7785);
and U8430 (N_8430,N_7357,N_7942);
and U8431 (N_8431,N_7482,N_7820);
and U8432 (N_8432,N_7982,N_7956);
and U8433 (N_8433,N_7282,N_7546);
nor U8434 (N_8434,N_7171,N_7940);
or U8435 (N_8435,N_7174,N_7955);
and U8436 (N_8436,N_7632,N_7496);
nor U8437 (N_8437,N_7403,N_7438);
nand U8438 (N_8438,N_7417,N_7246);
or U8439 (N_8439,N_7501,N_7281);
nor U8440 (N_8440,N_7823,N_7841);
nand U8441 (N_8441,N_7195,N_7084);
and U8442 (N_8442,N_7923,N_7472);
and U8443 (N_8443,N_7733,N_7039);
nand U8444 (N_8444,N_7231,N_7977);
or U8445 (N_8445,N_7862,N_7428);
and U8446 (N_8446,N_7248,N_7521);
or U8447 (N_8447,N_7524,N_7040);
nand U8448 (N_8448,N_7090,N_7230);
nor U8449 (N_8449,N_7005,N_7833);
or U8450 (N_8450,N_7167,N_7798);
or U8451 (N_8451,N_7523,N_7934);
or U8452 (N_8452,N_7236,N_7011);
or U8453 (N_8453,N_7680,N_7653);
nor U8454 (N_8454,N_7636,N_7792);
nand U8455 (N_8455,N_7141,N_7711);
nor U8456 (N_8456,N_7795,N_7640);
or U8457 (N_8457,N_7562,N_7919);
or U8458 (N_8458,N_7570,N_7557);
or U8459 (N_8459,N_7992,N_7567);
and U8460 (N_8460,N_7313,N_7738);
or U8461 (N_8461,N_7610,N_7884);
nor U8462 (N_8462,N_7783,N_7880);
nand U8463 (N_8463,N_7289,N_7960);
nor U8464 (N_8464,N_7794,N_7450);
and U8465 (N_8465,N_7061,N_7018);
nor U8466 (N_8466,N_7242,N_7435);
and U8467 (N_8467,N_7475,N_7629);
and U8468 (N_8468,N_7204,N_7703);
or U8469 (N_8469,N_7799,N_7764);
nor U8470 (N_8470,N_7757,N_7505);
or U8471 (N_8471,N_7999,N_7461);
nor U8472 (N_8472,N_7893,N_7145);
or U8473 (N_8473,N_7439,N_7410);
and U8474 (N_8474,N_7256,N_7336);
nand U8475 (N_8475,N_7625,N_7104);
nor U8476 (N_8476,N_7394,N_7315);
nor U8477 (N_8477,N_7397,N_7034);
nor U8478 (N_8478,N_7780,N_7958);
nand U8479 (N_8479,N_7463,N_7597);
xnor U8480 (N_8480,N_7788,N_7943);
nor U8481 (N_8481,N_7451,N_7264);
and U8482 (N_8482,N_7057,N_7362);
nor U8483 (N_8483,N_7344,N_7888);
and U8484 (N_8484,N_7358,N_7901);
nor U8485 (N_8485,N_7169,N_7423);
and U8486 (N_8486,N_7969,N_7668);
xor U8487 (N_8487,N_7508,N_7432);
and U8488 (N_8488,N_7274,N_7581);
nor U8489 (N_8489,N_7568,N_7645);
and U8490 (N_8490,N_7995,N_7964);
nand U8491 (N_8491,N_7350,N_7334);
and U8492 (N_8492,N_7060,N_7560);
and U8493 (N_8493,N_7811,N_7945);
and U8494 (N_8494,N_7112,N_7921);
nor U8495 (N_8495,N_7932,N_7575);
or U8496 (N_8496,N_7985,N_7695);
and U8497 (N_8497,N_7205,N_7469);
and U8498 (N_8498,N_7301,N_7401);
nor U8499 (N_8499,N_7300,N_7704);
nor U8500 (N_8500,N_7971,N_7966);
nor U8501 (N_8501,N_7457,N_7919);
or U8502 (N_8502,N_7549,N_7442);
and U8503 (N_8503,N_7582,N_7863);
and U8504 (N_8504,N_7998,N_7487);
or U8505 (N_8505,N_7064,N_7861);
nor U8506 (N_8506,N_7103,N_7088);
nand U8507 (N_8507,N_7862,N_7684);
nor U8508 (N_8508,N_7781,N_7081);
nor U8509 (N_8509,N_7139,N_7247);
or U8510 (N_8510,N_7736,N_7853);
nor U8511 (N_8511,N_7052,N_7806);
or U8512 (N_8512,N_7382,N_7779);
or U8513 (N_8513,N_7000,N_7917);
nor U8514 (N_8514,N_7228,N_7589);
nand U8515 (N_8515,N_7965,N_7452);
nor U8516 (N_8516,N_7000,N_7080);
nor U8517 (N_8517,N_7362,N_7899);
nand U8518 (N_8518,N_7103,N_7309);
and U8519 (N_8519,N_7238,N_7144);
and U8520 (N_8520,N_7165,N_7105);
and U8521 (N_8521,N_7273,N_7605);
nand U8522 (N_8522,N_7238,N_7167);
nand U8523 (N_8523,N_7969,N_7680);
nand U8524 (N_8524,N_7202,N_7710);
nor U8525 (N_8525,N_7288,N_7682);
nor U8526 (N_8526,N_7927,N_7030);
nor U8527 (N_8527,N_7998,N_7379);
nand U8528 (N_8528,N_7590,N_7837);
and U8529 (N_8529,N_7434,N_7605);
and U8530 (N_8530,N_7278,N_7186);
or U8531 (N_8531,N_7178,N_7412);
nand U8532 (N_8532,N_7997,N_7259);
or U8533 (N_8533,N_7691,N_7223);
or U8534 (N_8534,N_7580,N_7801);
or U8535 (N_8535,N_7100,N_7386);
nor U8536 (N_8536,N_7790,N_7291);
nand U8537 (N_8537,N_7140,N_7229);
and U8538 (N_8538,N_7270,N_7829);
and U8539 (N_8539,N_7948,N_7375);
or U8540 (N_8540,N_7621,N_7949);
nor U8541 (N_8541,N_7576,N_7306);
or U8542 (N_8542,N_7008,N_7613);
or U8543 (N_8543,N_7010,N_7835);
nor U8544 (N_8544,N_7384,N_7866);
or U8545 (N_8545,N_7769,N_7879);
or U8546 (N_8546,N_7155,N_7545);
nand U8547 (N_8547,N_7074,N_7512);
and U8548 (N_8548,N_7746,N_7543);
and U8549 (N_8549,N_7376,N_7827);
nor U8550 (N_8550,N_7538,N_7209);
nand U8551 (N_8551,N_7290,N_7004);
nand U8552 (N_8552,N_7938,N_7547);
and U8553 (N_8553,N_7114,N_7656);
and U8554 (N_8554,N_7188,N_7027);
and U8555 (N_8555,N_7041,N_7969);
or U8556 (N_8556,N_7530,N_7600);
nor U8557 (N_8557,N_7923,N_7556);
and U8558 (N_8558,N_7233,N_7393);
nor U8559 (N_8559,N_7882,N_7220);
and U8560 (N_8560,N_7676,N_7196);
and U8561 (N_8561,N_7835,N_7883);
nand U8562 (N_8562,N_7980,N_7386);
or U8563 (N_8563,N_7118,N_7942);
and U8564 (N_8564,N_7262,N_7340);
nand U8565 (N_8565,N_7449,N_7636);
nand U8566 (N_8566,N_7571,N_7044);
nor U8567 (N_8567,N_7317,N_7243);
and U8568 (N_8568,N_7976,N_7030);
and U8569 (N_8569,N_7855,N_7434);
and U8570 (N_8570,N_7850,N_7110);
nor U8571 (N_8571,N_7968,N_7728);
or U8572 (N_8572,N_7324,N_7942);
xnor U8573 (N_8573,N_7907,N_7759);
or U8574 (N_8574,N_7528,N_7045);
nand U8575 (N_8575,N_7846,N_7721);
nand U8576 (N_8576,N_7231,N_7778);
and U8577 (N_8577,N_7959,N_7704);
nor U8578 (N_8578,N_7871,N_7716);
or U8579 (N_8579,N_7339,N_7750);
nand U8580 (N_8580,N_7099,N_7407);
and U8581 (N_8581,N_7191,N_7254);
and U8582 (N_8582,N_7530,N_7806);
nand U8583 (N_8583,N_7535,N_7255);
nand U8584 (N_8584,N_7083,N_7613);
or U8585 (N_8585,N_7973,N_7377);
or U8586 (N_8586,N_7922,N_7500);
and U8587 (N_8587,N_7141,N_7938);
nor U8588 (N_8588,N_7409,N_7758);
nand U8589 (N_8589,N_7335,N_7227);
and U8590 (N_8590,N_7006,N_7539);
nor U8591 (N_8591,N_7825,N_7945);
and U8592 (N_8592,N_7641,N_7013);
or U8593 (N_8593,N_7355,N_7042);
nand U8594 (N_8594,N_7820,N_7463);
or U8595 (N_8595,N_7743,N_7146);
and U8596 (N_8596,N_7365,N_7667);
or U8597 (N_8597,N_7229,N_7642);
and U8598 (N_8598,N_7025,N_7870);
nand U8599 (N_8599,N_7674,N_7328);
and U8600 (N_8600,N_7297,N_7457);
and U8601 (N_8601,N_7690,N_7051);
nand U8602 (N_8602,N_7983,N_7508);
and U8603 (N_8603,N_7952,N_7755);
nand U8604 (N_8604,N_7229,N_7698);
and U8605 (N_8605,N_7859,N_7510);
nor U8606 (N_8606,N_7812,N_7207);
nand U8607 (N_8607,N_7574,N_7622);
xnor U8608 (N_8608,N_7314,N_7037);
nand U8609 (N_8609,N_7749,N_7934);
or U8610 (N_8610,N_7396,N_7473);
or U8611 (N_8611,N_7150,N_7628);
nand U8612 (N_8612,N_7977,N_7012);
and U8613 (N_8613,N_7711,N_7951);
nand U8614 (N_8614,N_7963,N_7261);
and U8615 (N_8615,N_7291,N_7822);
nand U8616 (N_8616,N_7037,N_7513);
or U8617 (N_8617,N_7721,N_7899);
nor U8618 (N_8618,N_7675,N_7487);
nand U8619 (N_8619,N_7864,N_7577);
or U8620 (N_8620,N_7412,N_7117);
nand U8621 (N_8621,N_7776,N_7365);
nand U8622 (N_8622,N_7218,N_7437);
or U8623 (N_8623,N_7546,N_7668);
or U8624 (N_8624,N_7936,N_7221);
and U8625 (N_8625,N_7881,N_7913);
nor U8626 (N_8626,N_7956,N_7162);
nor U8627 (N_8627,N_7268,N_7401);
nor U8628 (N_8628,N_7856,N_7244);
or U8629 (N_8629,N_7269,N_7419);
nor U8630 (N_8630,N_7014,N_7847);
and U8631 (N_8631,N_7512,N_7986);
nor U8632 (N_8632,N_7343,N_7747);
xnor U8633 (N_8633,N_7557,N_7228);
xnor U8634 (N_8634,N_7189,N_7227);
nand U8635 (N_8635,N_7313,N_7386);
nor U8636 (N_8636,N_7198,N_7913);
nand U8637 (N_8637,N_7665,N_7392);
nand U8638 (N_8638,N_7098,N_7112);
or U8639 (N_8639,N_7675,N_7431);
and U8640 (N_8640,N_7930,N_7806);
nand U8641 (N_8641,N_7765,N_7592);
nor U8642 (N_8642,N_7197,N_7210);
and U8643 (N_8643,N_7050,N_7013);
or U8644 (N_8644,N_7059,N_7396);
and U8645 (N_8645,N_7411,N_7039);
and U8646 (N_8646,N_7303,N_7872);
nand U8647 (N_8647,N_7231,N_7317);
nor U8648 (N_8648,N_7776,N_7682);
or U8649 (N_8649,N_7025,N_7521);
and U8650 (N_8650,N_7594,N_7060);
and U8651 (N_8651,N_7785,N_7910);
or U8652 (N_8652,N_7127,N_7616);
nand U8653 (N_8653,N_7785,N_7537);
or U8654 (N_8654,N_7972,N_7066);
nor U8655 (N_8655,N_7798,N_7951);
or U8656 (N_8656,N_7336,N_7813);
and U8657 (N_8657,N_7959,N_7821);
nand U8658 (N_8658,N_7392,N_7108);
or U8659 (N_8659,N_7553,N_7849);
and U8660 (N_8660,N_7804,N_7135);
nor U8661 (N_8661,N_7645,N_7572);
nand U8662 (N_8662,N_7158,N_7786);
or U8663 (N_8663,N_7642,N_7178);
and U8664 (N_8664,N_7330,N_7662);
nor U8665 (N_8665,N_7821,N_7681);
and U8666 (N_8666,N_7584,N_7788);
nor U8667 (N_8667,N_7766,N_7140);
nand U8668 (N_8668,N_7802,N_7771);
nand U8669 (N_8669,N_7251,N_7304);
or U8670 (N_8670,N_7288,N_7512);
or U8671 (N_8671,N_7020,N_7092);
nor U8672 (N_8672,N_7614,N_7229);
and U8673 (N_8673,N_7754,N_7174);
nor U8674 (N_8674,N_7612,N_7607);
nand U8675 (N_8675,N_7199,N_7182);
nand U8676 (N_8676,N_7395,N_7408);
and U8677 (N_8677,N_7049,N_7659);
or U8678 (N_8678,N_7349,N_7732);
and U8679 (N_8679,N_7312,N_7150);
or U8680 (N_8680,N_7688,N_7327);
or U8681 (N_8681,N_7497,N_7921);
nor U8682 (N_8682,N_7314,N_7997);
nor U8683 (N_8683,N_7924,N_7658);
nand U8684 (N_8684,N_7564,N_7651);
nor U8685 (N_8685,N_7126,N_7814);
and U8686 (N_8686,N_7253,N_7580);
or U8687 (N_8687,N_7423,N_7076);
nand U8688 (N_8688,N_7394,N_7787);
nor U8689 (N_8689,N_7197,N_7203);
and U8690 (N_8690,N_7265,N_7470);
nand U8691 (N_8691,N_7282,N_7238);
or U8692 (N_8692,N_7409,N_7512);
or U8693 (N_8693,N_7631,N_7872);
and U8694 (N_8694,N_7244,N_7110);
or U8695 (N_8695,N_7061,N_7476);
nor U8696 (N_8696,N_7562,N_7705);
or U8697 (N_8697,N_7077,N_7817);
nor U8698 (N_8698,N_7792,N_7921);
and U8699 (N_8699,N_7132,N_7876);
or U8700 (N_8700,N_7295,N_7993);
or U8701 (N_8701,N_7506,N_7648);
or U8702 (N_8702,N_7929,N_7196);
nand U8703 (N_8703,N_7113,N_7002);
or U8704 (N_8704,N_7671,N_7954);
and U8705 (N_8705,N_7493,N_7128);
nor U8706 (N_8706,N_7080,N_7044);
nor U8707 (N_8707,N_7714,N_7189);
and U8708 (N_8708,N_7316,N_7996);
nand U8709 (N_8709,N_7993,N_7281);
nand U8710 (N_8710,N_7819,N_7754);
or U8711 (N_8711,N_7123,N_7583);
or U8712 (N_8712,N_7014,N_7655);
xor U8713 (N_8713,N_7972,N_7460);
nor U8714 (N_8714,N_7922,N_7330);
or U8715 (N_8715,N_7371,N_7065);
and U8716 (N_8716,N_7316,N_7308);
nand U8717 (N_8717,N_7153,N_7103);
and U8718 (N_8718,N_7527,N_7770);
nor U8719 (N_8719,N_7977,N_7043);
and U8720 (N_8720,N_7920,N_7397);
or U8721 (N_8721,N_7555,N_7235);
nor U8722 (N_8722,N_7949,N_7555);
and U8723 (N_8723,N_7643,N_7635);
and U8724 (N_8724,N_7031,N_7353);
and U8725 (N_8725,N_7995,N_7815);
nand U8726 (N_8726,N_7826,N_7329);
nor U8727 (N_8727,N_7915,N_7637);
nand U8728 (N_8728,N_7177,N_7965);
xnor U8729 (N_8729,N_7272,N_7113);
and U8730 (N_8730,N_7370,N_7573);
nor U8731 (N_8731,N_7233,N_7650);
or U8732 (N_8732,N_7119,N_7913);
or U8733 (N_8733,N_7434,N_7974);
and U8734 (N_8734,N_7568,N_7818);
nor U8735 (N_8735,N_7554,N_7474);
and U8736 (N_8736,N_7160,N_7874);
nand U8737 (N_8737,N_7885,N_7084);
nand U8738 (N_8738,N_7884,N_7808);
and U8739 (N_8739,N_7618,N_7876);
or U8740 (N_8740,N_7975,N_7203);
or U8741 (N_8741,N_7957,N_7904);
nand U8742 (N_8742,N_7135,N_7676);
or U8743 (N_8743,N_7124,N_7089);
xnor U8744 (N_8744,N_7188,N_7451);
or U8745 (N_8745,N_7413,N_7913);
nor U8746 (N_8746,N_7180,N_7246);
and U8747 (N_8747,N_7105,N_7581);
nand U8748 (N_8748,N_7778,N_7868);
nand U8749 (N_8749,N_7704,N_7712);
nand U8750 (N_8750,N_7592,N_7835);
and U8751 (N_8751,N_7291,N_7611);
nor U8752 (N_8752,N_7677,N_7240);
nand U8753 (N_8753,N_7138,N_7168);
or U8754 (N_8754,N_7939,N_7969);
or U8755 (N_8755,N_7712,N_7474);
or U8756 (N_8756,N_7501,N_7901);
nor U8757 (N_8757,N_7928,N_7364);
nor U8758 (N_8758,N_7316,N_7351);
or U8759 (N_8759,N_7130,N_7415);
nand U8760 (N_8760,N_7140,N_7332);
nor U8761 (N_8761,N_7289,N_7931);
and U8762 (N_8762,N_7094,N_7621);
and U8763 (N_8763,N_7695,N_7226);
or U8764 (N_8764,N_7236,N_7791);
and U8765 (N_8765,N_7432,N_7879);
nor U8766 (N_8766,N_7002,N_7631);
nand U8767 (N_8767,N_7286,N_7648);
and U8768 (N_8768,N_7192,N_7117);
nand U8769 (N_8769,N_7143,N_7783);
nor U8770 (N_8770,N_7212,N_7616);
or U8771 (N_8771,N_7822,N_7330);
nand U8772 (N_8772,N_7915,N_7494);
or U8773 (N_8773,N_7658,N_7920);
or U8774 (N_8774,N_7080,N_7751);
nor U8775 (N_8775,N_7762,N_7167);
and U8776 (N_8776,N_7222,N_7701);
nand U8777 (N_8777,N_7403,N_7166);
and U8778 (N_8778,N_7558,N_7543);
and U8779 (N_8779,N_7134,N_7202);
nand U8780 (N_8780,N_7314,N_7038);
nor U8781 (N_8781,N_7325,N_7255);
or U8782 (N_8782,N_7038,N_7368);
and U8783 (N_8783,N_7287,N_7172);
nand U8784 (N_8784,N_7578,N_7680);
or U8785 (N_8785,N_7059,N_7882);
and U8786 (N_8786,N_7093,N_7331);
and U8787 (N_8787,N_7821,N_7854);
or U8788 (N_8788,N_7867,N_7009);
nor U8789 (N_8789,N_7617,N_7422);
nor U8790 (N_8790,N_7351,N_7806);
nand U8791 (N_8791,N_7723,N_7903);
or U8792 (N_8792,N_7279,N_7981);
nor U8793 (N_8793,N_7054,N_7224);
xnor U8794 (N_8794,N_7618,N_7598);
or U8795 (N_8795,N_7581,N_7564);
and U8796 (N_8796,N_7544,N_7343);
nand U8797 (N_8797,N_7481,N_7050);
nor U8798 (N_8798,N_7197,N_7663);
nand U8799 (N_8799,N_7089,N_7067);
nand U8800 (N_8800,N_7415,N_7264);
or U8801 (N_8801,N_7273,N_7776);
or U8802 (N_8802,N_7369,N_7912);
or U8803 (N_8803,N_7199,N_7492);
nor U8804 (N_8804,N_7100,N_7398);
nand U8805 (N_8805,N_7390,N_7431);
nand U8806 (N_8806,N_7279,N_7145);
or U8807 (N_8807,N_7813,N_7826);
or U8808 (N_8808,N_7487,N_7158);
nor U8809 (N_8809,N_7583,N_7044);
and U8810 (N_8810,N_7637,N_7694);
and U8811 (N_8811,N_7970,N_7699);
nor U8812 (N_8812,N_7402,N_7321);
nor U8813 (N_8813,N_7995,N_7457);
and U8814 (N_8814,N_7378,N_7666);
nor U8815 (N_8815,N_7345,N_7509);
nand U8816 (N_8816,N_7846,N_7455);
or U8817 (N_8817,N_7597,N_7370);
and U8818 (N_8818,N_7093,N_7181);
or U8819 (N_8819,N_7583,N_7949);
nor U8820 (N_8820,N_7857,N_7554);
or U8821 (N_8821,N_7987,N_7722);
and U8822 (N_8822,N_7553,N_7685);
nand U8823 (N_8823,N_7714,N_7664);
nor U8824 (N_8824,N_7451,N_7967);
xor U8825 (N_8825,N_7264,N_7832);
and U8826 (N_8826,N_7940,N_7371);
or U8827 (N_8827,N_7197,N_7813);
or U8828 (N_8828,N_7970,N_7270);
and U8829 (N_8829,N_7482,N_7154);
or U8830 (N_8830,N_7805,N_7601);
nand U8831 (N_8831,N_7850,N_7830);
nand U8832 (N_8832,N_7349,N_7191);
nor U8833 (N_8833,N_7576,N_7529);
and U8834 (N_8834,N_7702,N_7324);
or U8835 (N_8835,N_7344,N_7545);
and U8836 (N_8836,N_7867,N_7702);
nand U8837 (N_8837,N_7590,N_7118);
and U8838 (N_8838,N_7038,N_7160);
or U8839 (N_8839,N_7044,N_7688);
nand U8840 (N_8840,N_7521,N_7741);
nor U8841 (N_8841,N_7198,N_7964);
nor U8842 (N_8842,N_7969,N_7910);
nand U8843 (N_8843,N_7886,N_7373);
or U8844 (N_8844,N_7078,N_7774);
or U8845 (N_8845,N_7959,N_7022);
nor U8846 (N_8846,N_7640,N_7190);
nand U8847 (N_8847,N_7749,N_7855);
and U8848 (N_8848,N_7521,N_7763);
nor U8849 (N_8849,N_7332,N_7358);
nor U8850 (N_8850,N_7271,N_7015);
xnor U8851 (N_8851,N_7112,N_7848);
or U8852 (N_8852,N_7357,N_7921);
nor U8853 (N_8853,N_7081,N_7699);
or U8854 (N_8854,N_7086,N_7570);
and U8855 (N_8855,N_7525,N_7680);
and U8856 (N_8856,N_7686,N_7678);
and U8857 (N_8857,N_7134,N_7980);
xnor U8858 (N_8858,N_7834,N_7315);
or U8859 (N_8859,N_7938,N_7777);
nand U8860 (N_8860,N_7108,N_7349);
or U8861 (N_8861,N_7288,N_7911);
or U8862 (N_8862,N_7912,N_7354);
nand U8863 (N_8863,N_7305,N_7564);
or U8864 (N_8864,N_7954,N_7331);
or U8865 (N_8865,N_7330,N_7985);
nand U8866 (N_8866,N_7829,N_7170);
and U8867 (N_8867,N_7613,N_7232);
nor U8868 (N_8868,N_7541,N_7773);
or U8869 (N_8869,N_7730,N_7480);
nand U8870 (N_8870,N_7114,N_7412);
nor U8871 (N_8871,N_7286,N_7791);
or U8872 (N_8872,N_7868,N_7237);
nand U8873 (N_8873,N_7264,N_7444);
nand U8874 (N_8874,N_7193,N_7667);
or U8875 (N_8875,N_7232,N_7373);
and U8876 (N_8876,N_7266,N_7367);
and U8877 (N_8877,N_7485,N_7607);
and U8878 (N_8878,N_7077,N_7382);
nand U8879 (N_8879,N_7367,N_7347);
nand U8880 (N_8880,N_7841,N_7396);
or U8881 (N_8881,N_7749,N_7113);
nor U8882 (N_8882,N_7216,N_7108);
or U8883 (N_8883,N_7905,N_7114);
nor U8884 (N_8884,N_7303,N_7279);
nor U8885 (N_8885,N_7040,N_7355);
nor U8886 (N_8886,N_7546,N_7626);
nand U8887 (N_8887,N_7751,N_7809);
nand U8888 (N_8888,N_7053,N_7174);
or U8889 (N_8889,N_7624,N_7456);
nor U8890 (N_8890,N_7798,N_7858);
nor U8891 (N_8891,N_7263,N_7911);
and U8892 (N_8892,N_7580,N_7507);
nand U8893 (N_8893,N_7922,N_7784);
nor U8894 (N_8894,N_7892,N_7410);
and U8895 (N_8895,N_7670,N_7232);
or U8896 (N_8896,N_7584,N_7137);
nand U8897 (N_8897,N_7003,N_7046);
nor U8898 (N_8898,N_7819,N_7336);
xor U8899 (N_8899,N_7257,N_7501);
nor U8900 (N_8900,N_7253,N_7115);
nand U8901 (N_8901,N_7354,N_7943);
xnor U8902 (N_8902,N_7735,N_7042);
nor U8903 (N_8903,N_7411,N_7281);
and U8904 (N_8904,N_7655,N_7888);
or U8905 (N_8905,N_7584,N_7128);
nor U8906 (N_8906,N_7548,N_7336);
or U8907 (N_8907,N_7374,N_7296);
or U8908 (N_8908,N_7174,N_7871);
nor U8909 (N_8909,N_7748,N_7605);
and U8910 (N_8910,N_7640,N_7177);
and U8911 (N_8911,N_7280,N_7048);
nand U8912 (N_8912,N_7885,N_7163);
nor U8913 (N_8913,N_7726,N_7818);
or U8914 (N_8914,N_7978,N_7638);
or U8915 (N_8915,N_7433,N_7687);
and U8916 (N_8916,N_7102,N_7336);
and U8917 (N_8917,N_7146,N_7235);
and U8918 (N_8918,N_7075,N_7582);
nand U8919 (N_8919,N_7317,N_7373);
nor U8920 (N_8920,N_7566,N_7946);
and U8921 (N_8921,N_7859,N_7546);
or U8922 (N_8922,N_7767,N_7562);
nor U8923 (N_8923,N_7866,N_7905);
nand U8924 (N_8924,N_7283,N_7666);
or U8925 (N_8925,N_7334,N_7605);
and U8926 (N_8926,N_7388,N_7981);
or U8927 (N_8927,N_7764,N_7379);
or U8928 (N_8928,N_7778,N_7796);
xnor U8929 (N_8929,N_7400,N_7055);
nor U8930 (N_8930,N_7423,N_7080);
or U8931 (N_8931,N_7472,N_7619);
or U8932 (N_8932,N_7417,N_7153);
nand U8933 (N_8933,N_7157,N_7017);
nand U8934 (N_8934,N_7706,N_7100);
or U8935 (N_8935,N_7516,N_7963);
or U8936 (N_8936,N_7690,N_7273);
and U8937 (N_8937,N_7684,N_7922);
and U8938 (N_8938,N_7885,N_7805);
nor U8939 (N_8939,N_7928,N_7403);
or U8940 (N_8940,N_7810,N_7373);
and U8941 (N_8941,N_7258,N_7955);
or U8942 (N_8942,N_7469,N_7214);
nor U8943 (N_8943,N_7965,N_7693);
or U8944 (N_8944,N_7307,N_7367);
and U8945 (N_8945,N_7383,N_7017);
nand U8946 (N_8946,N_7908,N_7958);
nand U8947 (N_8947,N_7059,N_7219);
nand U8948 (N_8948,N_7367,N_7331);
nor U8949 (N_8949,N_7200,N_7461);
nand U8950 (N_8950,N_7451,N_7062);
and U8951 (N_8951,N_7427,N_7636);
or U8952 (N_8952,N_7653,N_7598);
nand U8953 (N_8953,N_7596,N_7461);
nor U8954 (N_8954,N_7878,N_7814);
nor U8955 (N_8955,N_7838,N_7971);
nor U8956 (N_8956,N_7494,N_7175);
xnor U8957 (N_8957,N_7495,N_7225);
and U8958 (N_8958,N_7265,N_7624);
and U8959 (N_8959,N_7548,N_7304);
nor U8960 (N_8960,N_7983,N_7621);
nor U8961 (N_8961,N_7718,N_7224);
and U8962 (N_8962,N_7446,N_7827);
or U8963 (N_8963,N_7284,N_7773);
and U8964 (N_8964,N_7750,N_7500);
xor U8965 (N_8965,N_7127,N_7838);
and U8966 (N_8966,N_7761,N_7738);
and U8967 (N_8967,N_7780,N_7256);
or U8968 (N_8968,N_7447,N_7336);
or U8969 (N_8969,N_7379,N_7495);
or U8970 (N_8970,N_7002,N_7961);
and U8971 (N_8971,N_7335,N_7608);
or U8972 (N_8972,N_7789,N_7008);
nor U8973 (N_8973,N_7838,N_7143);
or U8974 (N_8974,N_7539,N_7051);
xnor U8975 (N_8975,N_7369,N_7772);
nor U8976 (N_8976,N_7094,N_7609);
nand U8977 (N_8977,N_7879,N_7716);
or U8978 (N_8978,N_7996,N_7353);
or U8979 (N_8979,N_7026,N_7996);
nand U8980 (N_8980,N_7185,N_7092);
xor U8981 (N_8981,N_7654,N_7646);
and U8982 (N_8982,N_7372,N_7040);
nand U8983 (N_8983,N_7317,N_7052);
nor U8984 (N_8984,N_7014,N_7981);
or U8985 (N_8985,N_7371,N_7536);
nor U8986 (N_8986,N_7009,N_7664);
nand U8987 (N_8987,N_7297,N_7022);
or U8988 (N_8988,N_7791,N_7128);
and U8989 (N_8989,N_7630,N_7599);
and U8990 (N_8990,N_7079,N_7829);
nand U8991 (N_8991,N_7372,N_7892);
nor U8992 (N_8992,N_7904,N_7016);
nor U8993 (N_8993,N_7790,N_7452);
and U8994 (N_8994,N_7777,N_7264);
or U8995 (N_8995,N_7053,N_7712);
and U8996 (N_8996,N_7628,N_7000);
nor U8997 (N_8997,N_7064,N_7928);
nor U8998 (N_8998,N_7610,N_7675);
nor U8999 (N_8999,N_7996,N_7076);
or U9000 (N_9000,N_8622,N_8729);
and U9001 (N_9001,N_8690,N_8509);
and U9002 (N_9002,N_8401,N_8546);
nor U9003 (N_9003,N_8040,N_8723);
nor U9004 (N_9004,N_8349,N_8032);
nor U9005 (N_9005,N_8335,N_8074);
and U9006 (N_9006,N_8190,N_8938);
and U9007 (N_9007,N_8293,N_8997);
and U9008 (N_9008,N_8779,N_8771);
or U9009 (N_9009,N_8925,N_8072);
nor U9010 (N_9010,N_8863,N_8718);
xor U9011 (N_9011,N_8353,N_8113);
and U9012 (N_9012,N_8213,N_8902);
nand U9013 (N_9013,N_8035,N_8466);
nand U9014 (N_9014,N_8034,N_8756);
nand U9015 (N_9015,N_8002,N_8308);
and U9016 (N_9016,N_8602,N_8890);
or U9017 (N_9017,N_8667,N_8581);
nand U9018 (N_9018,N_8585,N_8411);
and U9019 (N_9019,N_8115,N_8854);
and U9020 (N_9020,N_8681,N_8506);
or U9021 (N_9021,N_8793,N_8721);
and U9022 (N_9022,N_8226,N_8534);
nand U9023 (N_9023,N_8805,N_8028);
and U9024 (N_9024,N_8281,N_8832);
and U9025 (N_9025,N_8322,N_8788);
nor U9026 (N_9026,N_8419,N_8862);
xor U9027 (N_9027,N_8640,N_8043);
nor U9028 (N_9028,N_8164,N_8892);
nor U9029 (N_9029,N_8387,N_8962);
nand U9030 (N_9030,N_8780,N_8031);
and U9031 (N_9031,N_8971,N_8166);
nor U9032 (N_9032,N_8237,N_8184);
and U9033 (N_9033,N_8926,N_8508);
nor U9034 (N_9034,N_8198,N_8671);
nor U9035 (N_9035,N_8445,N_8374);
nor U9036 (N_9036,N_8498,N_8452);
or U9037 (N_9037,N_8242,N_8417);
nand U9038 (N_9038,N_8936,N_8619);
or U9039 (N_9039,N_8144,N_8751);
or U9040 (N_9040,N_8029,N_8464);
nand U9041 (N_9041,N_8183,N_8995);
or U9042 (N_9042,N_8104,N_8341);
and U9043 (N_9043,N_8727,N_8342);
or U9044 (N_9044,N_8017,N_8261);
nor U9045 (N_9045,N_8803,N_8696);
nand U9046 (N_9046,N_8057,N_8064);
nand U9047 (N_9047,N_8864,N_8548);
nor U9048 (N_9048,N_8639,N_8837);
nand U9049 (N_9049,N_8791,N_8649);
and U9050 (N_9050,N_8071,N_8122);
and U9051 (N_9051,N_8354,N_8310);
and U9052 (N_9052,N_8384,N_8872);
and U9053 (N_9053,N_8940,N_8535);
or U9054 (N_9054,N_8066,N_8078);
or U9055 (N_9055,N_8448,N_8421);
or U9056 (N_9056,N_8594,N_8959);
nor U9057 (N_9057,N_8928,N_8303);
or U9058 (N_9058,N_8097,N_8912);
nor U9059 (N_9059,N_8138,N_8263);
and U9060 (N_9060,N_8063,N_8519);
and U9061 (N_9061,N_8675,N_8547);
nand U9062 (N_9062,N_8019,N_8740);
and U9063 (N_9063,N_8558,N_8825);
nand U9064 (N_9064,N_8259,N_8277);
and U9065 (N_9065,N_8255,N_8895);
nand U9066 (N_9066,N_8362,N_8116);
and U9067 (N_9067,N_8752,N_8893);
nor U9068 (N_9068,N_8045,N_8023);
nand U9069 (N_9069,N_8973,N_8518);
and U9070 (N_9070,N_8403,N_8267);
xnor U9071 (N_9071,N_8933,N_8566);
and U9072 (N_9072,N_8471,N_8501);
or U9073 (N_9073,N_8919,N_8150);
and U9074 (N_9074,N_8260,N_8358);
or U9075 (N_9075,N_8312,N_8024);
and U9076 (N_9076,N_8393,N_8661);
and U9077 (N_9077,N_8006,N_8219);
and U9078 (N_9078,N_8402,N_8268);
nand U9079 (N_9079,N_8824,N_8207);
nand U9080 (N_9080,N_8212,N_8795);
nand U9081 (N_9081,N_8099,N_8380);
and U9082 (N_9082,N_8388,N_8443);
nor U9083 (N_9083,N_8953,N_8192);
and U9084 (N_9084,N_8887,N_8672);
nor U9085 (N_9085,N_8470,N_8790);
nand U9086 (N_9086,N_8369,N_8128);
nand U9087 (N_9087,N_8822,N_8852);
and U9088 (N_9088,N_8203,N_8797);
xor U9089 (N_9089,N_8942,N_8450);
and U9090 (N_9090,N_8903,N_8200);
and U9091 (N_9091,N_8248,N_8980);
or U9092 (N_9092,N_8278,N_8230);
and U9093 (N_9093,N_8706,N_8974);
nor U9094 (N_9094,N_8279,N_8440);
nand U9095 (N_9095,N_8944,N_8699);
nor U9096 (N_9096,N_8305,N_8773);
or U9097 (N_9097,N_8073,N_8117);
nor U9098 (N_9098,N_8542,N_8720);
nor U9099 (N_9099,N_8961,N_8911);
xor U9100 (N_9100,N_8420,N_8205);
nor U9101 (N_9101,N_8968,N_8896);
or U9102 (N_9102,N_8127,N_8722);
or U9103 (N_9103,N_8931,N_8301);
or U9104 (N_9104,N_8060,N_8414);
and U9105 (N_9105,N_8357,N_8298);
and U9106 (N_9106,N_8586,N_8172);
and U9107 (N_9107,N_8486,N_8970);
nand U9108 (N_9108,N_8934,N_8886);
nor U9109 (N_9109,N_8676,N_8058);
or U9110 (N_9110,N_8784,N_8673);
nor U9111 (N_9111,N_8817,N_8476);
nor U9112 (N_9112,N_8449,N_8037);
or U9113 (N_9113,N_8777,N_8763);
and U9114 (N_9114,N_8734,N_8831);
or U9115 (N_9115,N_8713,N_8992);
or U9116 (N_9116,N_8601,N_8810);
nor U9117 (N_9117,N_8576,N_8525);
nand U9118 (N_9118,N_8493,N_8569);
and U9119 (N_9119,N_8759,N_8544);
nor U9120 (N_9120,N_8376,N_8819);
or U9121 (N_9121,N_8422,N_8733);
nand U9122 (N_9122,N_8287,N_8062);
nor U9123 (N_9123,N_8208,N_8774);
and U9124 (N_9124,N_8868,N_8846);
nand U9125 (N_9125,N_8372,N_8103);
and U9126 (N_9126,N_8584,N_8976);
nor U9127 (N_9127,N_8030,N_8725);
xor U9128 (N_9128,N_8536,N_8206);
nand U9129 (N_9129,N_8829,N_8054);
and U9130 (N_9130,N_8314,N_8254);
nand U9131 (N_9131,N_8964,N_8592);
xnor U9132 (N_9132,N_8177,N_8702);
nand U9133 (N_9133,N_8156,N_8036);
and U9134 (N_9134,N_8100,N_8361);
nor U9135 (N_9135,N_8528,N_8408);
and U9136 (N_9136,N_8583,N_8485);
and U9137 (N_9137,N_8913,N_8830);
nand U9138 (N_9138,N_8674,N_8530);
and U9139 (N_9139,N_8302,N_8628);
or U9140 (N_9140,N_8227,N_8855);
nor U9141 (N_9141,N_8008,N_8350);
and U9142 (N_9142,N_8404,N_8717);
and U9143 (N_9143,N_8806,N_8328);
or U9144 (N_9144,N_8869,N_8038);
nand U9145 (N_9145,N_8575,N_8923);
and U9146 (N_9146,N_8510,N_8413);
or U9147 (N_9147,N_8845,N_8056);
and U9148 (N_9148,N_8551,N_8977);
nand U9149 (N_9149,N_8613,N_8851);
and U9150 (N_9150,N_8772,N_8441);
and U9151 (N_9151,N_8552,N_8716);
nand U9152 (N_9152,N_8798,N_8426);
and U9153 (N_9153,N_8459,N_8764);
nor U9154 (N_9154,N_8669,N_8949);
nand U9155 (N_9155,N_8815,N_8630);
and U9156 (N_9156,N_8888,N_8329);
nand U9157 (N_9157,N_8410,N_8710);
and U9158 (N_9158,N_8231,N_8965);
and U9159 (N_9159,N_8339,N_8559);
or U9160 (N_9160,N_8707,N_8625);
nor U9161 (N_9161,N_8935,N_8407);
nor U9162 (N_9162,N_8048,N_8574);
nor U9163 (N_9163,N_8655,N_8635);
nor U9164 (N_9164,N_8238,N_8069);
nor U9165 (N_9165,N_8957,N_8685);
nand U9166 (N_9166,N_8873,N_8749);
xnor U9167 (N_9167,N_8521,N_8125);
or U9168 (N_9168,N_8275,N_8106);
nand U9169 (N_9169,N_8007,N_8646);
or U9170 (N_9170,N_8143,N_8334);
and U9171 (N_9171,N_8126,N_8804);
nor U9172 (N_9172,N_8665,N_8579);
or U9173 (N_9173,N_8446,N_8516);
nand U9174 (N_9174,N_8682,N_8611);
or U9175 (N_9175,N_8243,N_8090);
and U9176 (N_9176,N_8504,N_8637);
or U9177 (N_9177,N_8644,N_8969);
or U9178 (N_9178,N_8187,N_8194);
and U9179 (N_9179,N_8105,N_8463);
nor U9180 (N_9180,N_8306,N_8657);
or U9181 (N_9181,N_8119,N_8599);
nor U9182 (N_9182,N_8381,N_8332);
xnor U9183 (N_9183,N_8162,N_8220);
or U9184 (N_9184,N_8047,N_8891);
and U9185 (N_9185,N_8709,N_8222);
or U9186 (N_9186,N_8904,N_8169);
or U9187 (N_9187,N_8778,N_8315);
and U9188 (N_9188,N_8561,N_8745);
nand U9189 (N_9189,N_8295,N_8430);
nand U9190 (N_9190,N_8170,N_8762);
nor U9191 (N_9191,N_8171,N_8431);
nand U9192 (N_9192,N_8724,N_8787);
and U9193 (N_9193,N_8251,N_8311);
nand U9194 (N_9194,N_8000,N_8785);
and U9195 (N_9195,N_8370,N_8618);
nand U9196 (N_9196,N_8916,N_8726);
or U9197 (N_9197,N_8983,N_8768);
nand U9198 (N_9198,N_8889,N_8783);
nor U9199 (N_9199,N_8929,N_8433);
and U9200 (N_9200,N_8760,N_8405);
nand U9201 (N_9201,N_8866,N_8324);
nand U9202 (N_9202,N_8225,N_8526);
or U9203 (N_9203,N_8648,N_8879);
and U9204 (N_9204,N_8013,N_8397);
or U9205 (N_9205,N_8645,N_8683);
and U9206 (N_9206,N_8009,N_8826);
nor U9207 (N_9207,N_8967,N_8375);
nor U9208 (N_9208,N_8221,N_8107);
nor U9209 (N_9209,N_8603,N_8775);
nand U9210 (N_9210,N_8336,N_8309);
nor U9211 (N_9211,N_8877,N_8136);
and U9212 (N_9212,N_8499,N_8185);
xor U9213 (N_9213,N_8694,N_8130);
nand U9214 (N_9214,N_8598,N_8562);
nand U9215 (N_9215,N_8077,N_8697);
or U9216 (N_9216,N_8870,N_8587);
nand U9217 (N_9217,N_8214,N_8391);
nor U9218 (N_9218,N_8428,N_8621);
nor U9219 (N_9219,N_8321,N_8153);
and U9220 (N_9220,N_8055,N_8823);
or U9221 (N_9221,N_8642,N_8294);
and U9222 (N_9222,N_8157,N_8347);
nor U9223 (N_9223,N_8394,N_8480);
nand U9224 (N_9224,N_8897,N_8865);
or U9225 (N_9225,N_8258,N_8218);
nand U9226 (N_9226,N_8202,N_8998);
nor U9227 (N_9227,N_8507,N_8022);
nor U9228 (N_9228,N_8155,N_8059);
nor U9229 (N_9229,N_8615,N_8836);
nor U9230 (N_9230,N_8075,N_8741);
nor U9231 (N_9231,N_8092,N_8271);
nand U9232 (N_9232,N_8839,N_8432);
or U9233 (N_9233,N_8299,N_8182);
or U9234 (N_9234,N_8487,N_8545);
or U9235 (N_9235,N_8094,N_8366);
nand U9236 (N_9236,N_8849,N_8769);
nor U9237 (N_9237,N_8132,N_8371);
nand U9238 (N_9238,N_8827,N_8500);
nor U9239 (N_9239,N_8910,N_8666);
nor U9240 (N_9240,N_8605,N_8564);
nand U9241 (N_9241,N_8313,N_8765);
or U9242 (N_9242,N_8282,N_8999);
nor U9243 (N_9243,N_8927,N_8898);
and U9244 (N_9244,N_8816,N_8137);
nand U9245 (N_9245,N_8050,N_8027);
and U9246 (N_9246,N_8490,N_8560);
nand U9247 (N_9247,N_8684,N_8146);
and U9248 (N_9248,N_8447,N_8654);
and U9249 (N_9249,N_8712,N_8604);
nand U9250 (N_9250,N_8847,N_8531);
and U9251 (N_9251,N_8262,N_8240);
or U9252 (N_9252,N_8856,N_8761);
nand U9253 (N_9253,N_8320,N_8894);
nand U9254 (N_9254,N_8860,N_8624);
and U9255 (N_9255,N_8689,N_8241);
xnor U9256 (N_9256,N_8838,N_8285);
nor U9257 (N_9257,N_8818,N_8399);
nand U9258 (N_9258,N_8932,N_8789);
or U9259 (N_9259,N_8568,N_8101);
nor U9260 (N_9260,N_8691,N_8900);
nor U9261 (N_9261,N_8861,N_8664);
nor U9262 (N_9262,N_8921,N_8539);
nor U9263 (N_9263,N_8327,N_8236);
and U9264 (N_9264,N_8738,N_8120);
and U9265 (N_9265,N_8821,N_8478);
nand U9266 (N_9266,N_8437,N_8468);
nor U9267 (N_9267,N_8735,N_8616);
nor U9268 (N_9268,N_8754,N_8700);
or U9269 (N_9269,N_8042,N_8475);
and U9270 (N_9270,N_8416,N_8705);
nand U9271 (N_9271,N_8692,N_8981);
nand U9272 (N_9272,N_8833,N_8907);
or U9273 (N_9273,N_8757,N_8307);
or U9274 (N_9274,N_8245,N_8946);
nor U9275 (N_9275,N_8139,N_8522);
xor U9276 (N_9276,N_8800,N_8317);
nand U9277 (N_9277,N_8828,N_8383);
nand U9278 (N_9278,N_8079,N_8010);
xnor U9279 (N_9279,N_8858,N_8356);
or U9280 (N_9280,N_8363,N_8770);
nand U9281 (N_9281,N_8917,N_8954);
nand U9282 (N_9282,N_8193,N_8112);
or U9283 (N_9283,N_8265,N_8914);
nor U9284 (N_9284,N_8151,N_8496);
nand U9285 (N_9285,N_8148,N_8958);
nor U9286 (N_9286,N_8986,N_8427);
nand U9287 (N_9287,N_8052,N_8367);
nand U9288 (N_9288,N_8633,N_8623);
nand U9289 (N_9289,N_8109,N_8606);
or U9290 (N_9290,N_8880,N_8386);
nand U9291 (N_9291,N_8001,N_8435);
or U9292 (N_9292,N_8085,N_8316);
xnor U9293 (N_9293,N_8110,N_8807);
or U9294 (N_9294,N_8458,N_8631);
nand U9295 (N_9295,N_8044,N_8456);
or U9296 (N_9296,N_8406,N_8686);
and U9297 (N_9297,N_8515,N_8679);
and U9298 (N_9298,N_8211,N_8163);
nor U9299 (N_9299,N_8159,N_8972);
or U9300 (N_9300,N_8960,N_8479);
nor U9301 (N_9301,N_8589,N_8084);
nand U9302 (N_9302,N_8878,N_8520);
nor U9303 (N_9303,N_8739,N_8351);
nand U9304 (N_9304,N_8451,N_8750);
and U9305 (N_9305,N_8532,N_8502);
or U9306 (N_9306,N_8874,N_8434);
nor U9307 (N_9307,N_8199,N_8698);
or U9308 (N_9308,N_8483,N_8111);
and U9309 (N_9309,N_8996,N_8990);
xor U9310 (N_9310,N_8453,N_8053);
nor U9311 (N_9311,N_8677,N_8252);
nand U9312 (N_9312,N_8550,N_8337);
or U9313 (N_9313,N_8292,N_8175);
or U9314 (N_9314,N_8802,N_8688);
nand U9315 (N_9315,N_8840,N_8930);
nand U9316 (N_9316,N_8093,N_8647);
nand U9317 (N_9317,N_8472,N_8975);
nor U9318 (N_9318,N_8368,N_8429);
xor U9319 (N_9319,N_8235,N_8348);
nand U9320 (N_9320,N_8273,N_8484);
nand U9321 (N_9321,N_8003,N_8796);
or U9322 (N_9322,N_8881,N_8557);
and U9323 (N_9323,N_8956,N_8168);
nand U9324 (N_9324,N_8607,N_8680);
or U9325 (N_9325,N_8901,N_8549);
and U9326 (N_9326,N_8442,N_8591);
or U9327 (N_9327,N_8588,N_8494);
xnor U9328 (N_9328,N_8991,N_8253);
or U9329 (N_9329,N_8985,N_8488);
and U9330 (N_9330,N_8814,N_8668);
or U9331 (N_9331,N_8951,N_8149);
nor U9332 (N_9332,N_8952,N_8651);
nor U9333 (N_9333,N_8670,N_8323);
or U9334 (N_9334,N_8989,N_8269);
and U9335 (N_9335,N_8517,N_8196);
nor U9336 (N_9336,N_8409,N_8915);
nand U9337 (N_9337,N_8284,N_8834);
nand U9338 (N_9338,N_8482,N_8514);
nor U9339 (N_9339,N_8563,N_8161);
nor U9340 (N_9340,N_8994,N_8270);
nand U9341 (N_9341,N_8004,N_8714);
nor U9342 (N_9342,N_8141,N_8905);
and U9343 (N_9343,N_8179,N_8979);
nand U9344 (N_9344,N_8246,N_8108);
and U9345 (N_9345,N_8233,N_8018);
and U9346 (N_9346,N_8663,N_8918);
xnor U9347 (N_9347,N_8652,N_8636);
nor U9348 (N_9348,N_8118,N_8039);
or U9349 (N_9349,N_8133,N_8080);
or U9350 (N_9350,N_8656,N_8065);
nor U9351 (N_9351,N_8614,N_8180);
nor U9352 (N_9352,N_8481,N_8014);
nor U9353 (N_9353,N_8626,N_8088);
nand U9354 (N_9354,N_8215,N_8596);
nor U9355 (N_9355,N_8378,N_8853);
nor U9356 (N_9356,N_8844,N_8966);
and U9357 (N_9357,N_8529,N_8081);
or U9358 (N_9358,N_8091,N_8503);
and U9359 (N_9359,N_8608,N_8266);
xnor U9360 (N_9360,N_8082,N_8781);
nor U9361 (N_9361,N_8939,N_8609);
nor U9362 (N_9362,N_8385,N_8473);
and U9363 (N_9363,N_8859,N_8540);
nor U9364 (N_9364,N_8753,N_8121);
nor U9365 (N_9365,N_8289,N_8181);
nand U9366 (N_9366,N_8595,N_8297);
and U9367 (N_9367,N_8573,N_8033);
xor U9368 (N_9368,N_8474,N_8909);
nand U9369 (N_9369,N_8590,N_8597);
xnor U9370 (N_9370,N_8687,N_8343);
nor U9371 (N_9371,N_8283,N_8167);
nor U9372 (N_9372,N_8249,N_8813);
and U9373 (N_9373,N_8497,N_8556);
and U9374 (N_9374,N_8732,N_8742);
and U9375 (N_9375,N_8577,N_8578);
xor U9376 (N_9376,N_8715,N_8477);
and U9377 (N_9377,N_8178,N_8489);
nand U9378 (N_9378,N_8580,N_8012);
nor U9379 (N_9379,N_8086,N_8145);
and U9380 (N_9380,N_8461,N_8244);
nor U9381 (N_9381,N_8454,N_8899);
nor U9382 (N_9382,N_8982,N_8610);
and U9383 (N_9383,N_8331,N_8660);
and U9384 (N_9384,N_8061,N_8993);
nor U9385 (N_9385,N_8746,N_8462);
and U9386 (N_9386,N_8216,N_8924);
and U9387 (N_9387,N_8300,N_8377);
nor U9388 (N_9388,N_8129,N_8436);
and U9389 (N_9389,N_8988,N_8189);
nor U9390 (N_9390,N_8955,N_8850);
nand U9391 (N_9391,N_8650,N_8703);
and U9392 (N_9392,N_8820,N_8280);
nor U9393 (N_9393,N_8567,N_8812);
nand U9394 (N_9394,N_8809,N_8906);
xnor U9395 (N_9395,N_8304,N_8201);
or U9396 (N_9396,N_8748,N_8076);
and U9397 (N_9397,N_8617,N_8782);
and U9398 (N_9398,N_8704,N_8843);
nand U9399 (N_9399,N_8412,N_8658);
or U9400 (N_9400,N_8398,N_8444);
or U9401 (N_9401,N_8743,N_8465);
nor U9402 (N_9402,N_8209,N_8087);
or U9403 (N_9403,N_8016,N_8659);
nor U9404 (N_9404,N_8011,N_8555);
nor U9405 (N_9405,N_8389,N_8695);
or U9406 (N_9406,N_8867,N_8641);
and U9407 (N_9407,N_8360,N_8786);
and U9408 (N_9408,N_8392,N_8799);
or U9409 (N_9409,N_8922,N_8067);
nor U9410 (N_9410,N_8296,N_8096);
and U9411 (N_9411,N_8600,N_8191);
and U9412 (N_9412,N_8176,N_8025);
or U9413 (N_9413,N_8257,N_8662);
and U9414 (N_9414,N_8920,N_8882);
and U9415 (N_9415,N_8538,N_8693);
nand U9416 (N_9416,N_8134,N_8424);
or U9417 (N_9417,N_8095,N_8131);
or U9418 (N_9418,N_8264,N_8083);
nand U9419 (N_9419,N_8020,N_8512);
nand U9420 (N_9420,N_8229,N_8570);
or U9421 (N_9421,N_8731,N_8565);
or U9422 (N_9422,N_8359,N_8767);
or U9423 (N_9423,N_8719,N_8533);
nor U9424 (N_9424,N_8553,N_8541);
nor U9425 (N_9425,N_8188,N_8195);
nand U9426 (N_9426,N_8758,N_8158);
or U9427 (N_9427,N_8286,N_8423);
or U9428 (N_9428,N_8744,N_8152);
or U9429 (N_9429,N_8792,N_8593);
nand U9430 (N_9430,N_8345,N_8492);
or U9431 (N_9431,N_8395,N_8841);
nand U9432 (N_9432,N_8455,N_8276);
or U9433 (N_9433,N_8288,N_8875);
and U9434 (N_9434,N_8711,N_8883);
nor U9435 (N_9435,N_8495,N_8941);
and U9436 (N_9436,N_8114,N_8848);
and U9437 (N_9437,N_8232,N_8140);
or U9438 (N_9438,N_8643,N_8963);
nand U9439 (N_9439,N_8250,N_8174);
and U9440 (N_9440,N_8333,N_8505);
and U9441 (N_9441,N_8467,N_8124);
or U9442 (N_9442,N_8021,N_8382);
nor U9443 (N_9443,N_8885,N_8554);
or U9444 (N_9444,N_8186,N_8364);
nor U9445 (N_9445,N_8123,N_8290);
nor U9446 (N_9446,N_8701,N_8572);
and U9447 (N_9447,N_8318,N_8801);
or U9448 (N_9448,N_8046,N_8835);
and U9449 (N_9449,N_8272,N_8415);
or U9450 (N_9450,N_8620,N_8365);
nand U9451 (N_9451,N_8638,N_8811);
nor U9452 (N_9452,N_8256,N_8527);
or U9453 (N_9453,N_8747,N_8418);
nor U9454 (N_9454,N_8766,N_8049);
nand U9455 (N_9455,N_8755,N_8632);
and U9456 (N_9456,N_8239,N_8987);
nand U9457 (N_9457,N_8326,N_8026);
or U9458 (N_9458,N_8173,N_8224);
and U9459 (N_9459,N_8160,N_8228);
and U9460 (N_9460,N_8340,N_8247);
and U9461 (N_9461,N_8943,N_8438);
or U9462 (N_9462,N_8884,N_8460);
and U9463 (N_9463,N_8776,N_8102);
and U9464 (N_9464,N_8947,N_8338);
nand U9465 (N_9465,N_8937,N_8612);
nand U9466 (N_9466,N_8400,N_8736);
xnor U9467 (N_9467,N_8015,N_8876);
or U9468 (N_9468,N_8325,N_8330);
or U9469 (N_9469,N_8948,N_8197);
or U9470 (N_9470,N_8469,N_8629);
nor U9471 (N_9471,N_8978,N_8728);
nor U9472 (N_9472,N_8147,N_8154);
and U9473 (N_9473,N_8005,N_8165);
nor U9474 (N_9474,N_8439,N_8135);
and U9475 (N_9475,N_8204,N_8217);
nor U9476 (N_9476,N_8511,N_8210);
nand U9477 (N_9477,N_8070,N_8041);
or U9478 (N_9478,N_8950,N_8571);
or U9479 (N_9479,N_8627,N_8730);
or U9480 (N_9480,N_8373,N_8379);
and U9481 (N_9481,N_8513,N_8537);
or U9482 (N_9482,N_8523,N_8842);
and U9483 (N_9483,N_8794,N_8396);
or U9484 (N_9484,N_8984,N_8274);
nor U9485 (N_9485,N_8634,N_8346);
and U9486 (N_9486,N_8708,N_8223);
nand U9487 (N_9487,N_8808,N_8355);
nand U9488 (N_9488,N_8425,N_8582);
nand U9489 (N_9489,N_8857,N_8871);
or U9490 (N_9490,N_8098,N_8068);
and U9491 (N_9491,N_8945,N_8653);
and U9492 (N_9492,N_8543,N_8319);
xor U9493 (N_9493,N_8524,N_8234);
nor U9494 (N_9494,N_8908,N_8344);
nor U9495 (N_9495,N_8089,N_8142);
or U9496 (N_9496,N_8491,N_8390);
nand U9497 (N_9497,N_8678,N_8291);
nor U9498 (N_9498,N_8457,N_8352);
xnor U9499 (N_9499,N_8737,N_8051);
nor U9500 (N_9500,N_8736,N_8127);
and U9501 (N_9501,N_8470,N_8945);
nor U9502 (N_9502,N_8192,N_8873);
nand U9503 (N_9503,N_8502,N_8827);
and U9504 (N_9504,N_8726,N_8753);
or U9505 (N_9505,N_8175,N_8925);
or U9506 (N_9506,N_8174,N_8878);
or U9507 (N_9507,N_8144,N_8071);
or U9508 (N_9508,N_8393,N_8564);
nor U9509 (N_9509,N_8566,N_8711);
xnor U9510 (N_9510,N_8621,N_8110);
or U9511 (N_9511,N_8728,N_8380);
nor U9512 (N_9512,N_8636,N_8572);
and U9513 (N_9513,N_8275,N_8119);
and U9514 (N_9514,N_8074,N_8588);
nor U9515 (N_9515,N_8721,N_8622);
or U9516 (N_9516,N_8948,N_8360);
and U9517 (N_9517,N_8994,N_8047);
and U9518 (N_9518,N_8668,N_8499);
xor U9519 (N_9519,N_8769,N_8630);
xor U9520 (N_9520,N_8629,N_8987);
nor U9521 (N_9521,N_8940,N_8805);
nor U9522 (N_9522,N_8468,N_8118);
or U9523 (N_9523,N_8896,N_8970);
or U9524 (N_9524,N_8751,N_8603);
nor U9525 (N_9525,N_8460,N_8575);
and U9526 (N_9526,N_8493,N_8974);
xnor U9527 (N_9527,N_8308,N_8071);
nor U9528 (N_9528,N_8012,N_8472);
nor U9529 (N_9529,N_8383,N_8267);
nand U9530 (N_9530,N_8398,N_8990);
nand U9531 (N_9531,N_8893,N_8681);
or U9532 (N_9532,N_8918,N_8037);
nand U9533 (N_9533,N_8656,N_8326);
and U9534 (N_9534,N_8846,N_8238);
and U9535 (N_9535,N_8362,N_8779);
and U9536 (N_9536,N_8996,N_8521);
or U9537 (N_9537,N_8094,N_8768);
or U9538 (N_9538,N_8561,N_8398);
and U9539 (N_9539,N_8245,N_8587);
nor U9540 (N_9540,N_8012,N_8058);
nand U9541 (N_9541,N_8420,N_8965);
nor U9542 (N_9542,N_8487,N_8282);
nand U9543 (N_9543,N_8097,N_8119);
nor U9544 (N_9544,N_8128,N_8633);
nor U9545 (N_9545,N_8352,N_8824);
xnor U9546 (N_9546,N_8888,N_8491);
nor U9547 (N_9547,N_8857,N_8793);
nand U9548 (N_9548,N_8650,N_8066);
nand U9549 (N_9549,N_8437,N_8411);
nand U9550 (N_9550,N_8536,N_8779);
nor U9551 (N_9551,N_8548,N_8831);
nand U9552 (N_9552,N_8709,N_8919);
or U9553 (N_9553,N_8615,N_8324);
or U9554 (N_9554,N_8097,N_8245);
nand U9555 (N_9555,N_8094,N_8142);
nor U9556 (N_9556,N_8978,N_8533);
nand U9557 (N_9557,N_8592,N_8665);
nor U9558 (N_9558,N_8205,N_8229);
nor U9559 (N_9559,N_8825,N_8413);
and U9560 (N_9560,N_8716,N_8183);
and U9561 (N_9561,N_8401,N_8689);
and U9562 (N_9562,N_8214,N_8752);
nor U9563 (N_9563,N_8749,N_8699);
xor U9564 (N_9564,N_8188,N_8113);
nand U9565 (N_9565,N_8723,N_8957);
nor U9566 (N_9566,N_8180,N_8345);
nand U9567 (N_9567,N_8017,N_8149);
nand U9568 (N_9568,N_8765,N_8745);
nor U9569 (N_9569,N_8420,N_8120);
nor U9570 (N_9570,N_8657,N_8111);
and U9571 (N_9571,N_8610,N_8410);
or U9572 (N_9572,N_8338,N_8086);
and U9573 (N_9573,N_8123,N_8307);
or U9574 (N_9574,N_8287,N_8274);
and U9575 (N_9575,N_8488,N_8973);
and U9576 (N_9576,N_8485,N_8033);
or U9577 (N_9577,N_8964,N_8343);
nor U9578 (N_9578,N_8076,N_8378);
nor U9579 (N_9579,N_8272,N_8630);
nand U9580 (N_9580,N_8813,N_8161);
nand U9581 (N_9581,N_8568,N_8489);
nor U9582 (N_9582,N_8946,N_8502);
nand U9583 (N_9583,N_8851,N_8084);
nand U9584 (N_9584,N_8995,N_8596);
nand U9585 (N_9585,N_8829,N_8421);
or U9586 (N_9586,N_8615,N_8716);
nor U9587 (N_9587,N_8493,N_8867);
nand U9588 (N_9588,N_8542,N_8476);
nand U9589 (N_9589,N_8668,N_8055);
nand U9590 (N_9590,N_8234,N_8555);
nor U9591 (N_9591,N_8208,N_8023);
or U9592 (N_9592,N_8938,N_8897);
nor U9593 (N_9593,N_8502,N_8495);
and U9594 (N_9594,N_8655,N_8183);
nor U9595 (N_9595,N_8870,N_8881);
and U9596 (N_9596,N_8015,N_8607);
nor U9597 (N_9597,N_8966,N_8383);
and U9598 (N_9598,N_8455,N_8072);
nand U9599 (N_9599,N_8148,N_8585);
and U9600 (N_9600,N_8641,N_8374);
nand U9601 (N_9601,N_8588,N_8844);
and U9602 (N_9602,N_8583,N_8349);
or U9603 (N_9603,N_8780,N_8716);
and U9604 (N_9604,N_8513,N_8794);
and U9605 (N_9605,N_8632,N_8789);
and U9606 (N_9606,N_8769,N_8959);
or U9607 (N_9607,N_8839,N_8952);
or U9608 (N_9608,N_8361,N_8969);
nand U9609 (N_9609,N_8048,N_8655);
or U9610 (N_9610,N_8960,N_8186);
nor U9611 (N_9611,N_8708,N_8477);
and U9612 (N_9612,N_8785,N_8929);
nor U9613 (N_9613,N_8852,N_8554);
nor U9614 (N_9614,N_8142,N_8672);
nor U9615 (N_9615,N_8740,N_8897);
nand U9616 (N_9616,N_8381,N_8524);
nand U9617 (N_9617,N_8423,N_8906);
nor U9618 (N_9618,N_8183,N_8844);
nor U9619 (N_9619,N_8056,N_8627);
and U9620 (N_9620,N_8733,N_8706);
or U9621 (N_9621,N_8953,N_8712);
nand U9622 (N_9622,N_8603,N_8962);
and U9623 (N_9623,N_8959,N_8173);
nand U9624 (N_9624,N_8879,N_8928);
nor U9625 (N_9625,N_8169,N_8120);
or U9626 (N_9626,N_8336,N_8504);
or U9627 (N_9627,N_8050,N_8885);
or U9628 (N_9628,N_8896,N_8649);
or U9629 (N_9629,N_8827,N_8580);
or U9630 (N_9630,N_8499,N_8465);
or U9631 (N_9631,N_8846,N_8694);
nand U9632 (N_9632,N_8374,N_8950);
nor U9633 (N_9633,N_8291,N_8848);
xnor U9634 (N_9634,N_8941,N_8803);
nand U9635 (N_9635,N_8048,N_8252);
and U9636 (N_9636,N_8666,N_8083);
or U9637 (N_9637,N_8049,N_8513);
nand U9638 (N_9638,N_8985,N_8360);
nor U9639 (N_9639,N_8773,N_8390);
nand U9640 (N_9640,N_8418,N_8532);
or U9641 (N_9641,N_8365,N_8289);
nor U9642 (N_9642,N_8789,N_8620);
nand U9643 (N_9643,N_8105,N_8440);
nor U9644 (N_9644,N_8032,N_8661);
nand U9645 (N_9645,N_8306,N_8976);
or U9646 (N_9646,N_8416,N_8963);
nor U9647 (N_9647,N_8274,N_8515);
and U9648 (N_9648,N_8768,N_8177);
nand U9649 (N_9649,N_8522,N_8825);
or U9650 (N_9650,N_8349,N_8953);
nor U9651 (N_9651,N_8850,N_8294);
or U9652 (N_9652,N_8883,N_8770);
or U9653 (N_9653,N_8447,N_8411);
nand U9654 (N_9654,N_8546,N_8353);
or U9655 (N_9655,N_8201,N_8440);
nand U9656 (N_9656,N_8884,N_8107);
nor U9657 (N_9657,N_8140,N_8632);
and U9658 (N_9658,N_8404,N_8852);
nor U9659 (N_9659,N_8256,N_8222);
nand U9660 (N_9660,N_8526,N_8577);
nor U9661 (N_9661,N_8085,N_8272);
nor U9662 (N_9662,N_8974,N_8368);
or U9663 (N_9663,N_8414,N_8003);
nor U9664 (N_9664,N_8976,N_8926);
and U9665 (N_9665,N_8640,N_8850);
or U9666 (N_9666,N_8736,N_8092);
nand U9667 (N_9667,N_8440,N_8303);
nor U9668 (N_9668,N_8828,N_8446);
nand U9669 (N_9669,N_8380,N_8570);
or U9670 (N_9670,N_8667,N_8384);
and U9671 (N_9671,N_8247,N_8586);
nand U9672 (N_9672,N_8392,N_8130);
nand U9673 (N_9673,N_8854,N_8132);
and U9674 (N_9674,N_8010,N_8188);
nor U9675 (N_9675,N_8295,N_8641);
nand U9676 (N_9676,N_8647,N_8277);
nand U9677 (N_9677,N_8230,N_8522);
nand U9678 (N_9678,N_8756,N_8280);
nor U9679 (N_9679,N_8681,N_8583);
and U9680 (N_9680,N_8092,N_8974);
and U9681 (N_9681,N_8393,N_8095);
and U9682 (N_9682,N_8612,N_8924);
xnor U9683 (N_9683,N_8267,N_8621);
or U9684 (N_9684,N_8511,N_8674);
nand U9685 (N_9685,N_8154,N_8180);
and U9686 (N_9686,N_8108,N_8139);
or U9687 (N_9687,N_8867,N_8008);
nand U9688 (N_9688,N_8345,N_8516);
and U9689 (N_9689,N_8548,N_8238);
and U9690 (N_9690,N_8433,N_8299);
nor U9691 (N_9691,N_8122,N_8837);
nor U9692 (N_9692,N_8166,N_8872);
and U9693 (N_9693,N_8855,N_8818);
nand U9694 (N_9694,N_8292,N_8128);
and U9695 (N_9695,N_8262,N_8518);
nor U9696 (N_9696,N_8947,N_8653);
nand U9697 (N_9697,N_8438,N_8755);
nand U9698 (N_9698,N_8344,N_8464);
nor U9699 (N_9699,N_8397,N_8136);
or U9700 (N_9700,N_8081,N_8200);
or U9701 (N_9701,N_8561,N_8986);
and U9702 (N_9702,N_8814,N_8524);
nor U9703 (N_9703,N_8245,N_8885);
nand U9704 (N_9704,N_8634,N_8643);
or U9705 (N_9705,N_8503,N_8337);
xnor U9706 (N_9706,N_8852,N_8553);
nand U9707 (N_9707,N_8366,N_8722);
nand U9708 (N_9708,N_8824,N_8585);
or U9709 (N_9709,N_8764,N_8800);
nand U9710 (N_9710,N_8335,N_8652);
and U9711 (N_9711,N_8394,N_8308);
and U9712 (N_9712,N_8320,N_8637);
nor U9713 (N_9713,N_8901,N_8855);
nor U9714 (N_9714,N_8828,N_8907);
or U9715 (N_9715,N_8842,N_8787);
and U9716 (N_9716,N_8865,N_8636);
and U9717 (N_9717,N_8925,N_8886);
nor U9718 (N_9718,N_8071,N_8674);
nand U9719 (N_9719,N_8866,N_8705);
and U9720 (N_9720,N_8009,N_8143);
nand U9721 (N_9721,N_8462,N_8345);
and U9722 (N_9722,N_8694,N_8780);
and U9723 (N_9723,N_8956,N_8776);
or U9724 (N_9724,N_8718,N_8751);
xnor U9725 (N_9725,N_8393,N_8699);
nand U9726 (N_9726,N_8836,N_8157);
and U9727 (N_9727,N_8045,N_8083);
nand U9728 (N_9728,N_8402,N_8995);
nand U9729 (N_9729,N_8289,N_8126);
and U9730 (N_9730,N_8886,N_8219);
and U9731 (N_9731,N_8745,N_8600);
nand U9732 (N_9732,N_8100,N_8946);
xor U9733 (N_9733,N_8358,N_8230);
and U9734 (N_9734,N_8862,N_8159);
nor U9735 (N_9735,N_8854,N_8606);
nand U9736 (N_9736,N_8014,N_8976);
and U9737 (N_9737,N_8765,N_8994);
or U9738 (N_9738,N_8337,N_8564);
nor U9739 (N_9739,N_8539,N_8659);
nand U9740 (N_9740,N_8910,N_8825);
and U9741 (N_9741,N_8337,N_8704);
or U9742 (N_9742,N_8313,N_8971);
and U9743 (N_9743,N_8457,N_8026);
and U9744 (N_9744,N_8894,N_8953);
and U9745 (N_9745,N_8046,N_8450);
nand U9746 (N_9746,N_8572,N_8327);
nand U9747 (N_9747,N_8845,N_8710);
nand U9748 (N_9748,N_8966,N_8363);
or U9749 (N_9749,N_8661,N_8585);
nand U9750 (N_9750,N_8487,N_8173);
and U9751 (N_9751,N_8482,N_8176);
nand U9752 (N_9752,N_8435,N_8371);
nor U9753 (N_9753,N_8435,N_8650);
or U9754 (N_9754,N_8573,N_8906);
and U9755 (N_9755,N_8837,N_8435);
and U9756 (N_9756,N_8203,N_8066);
nand U9757 (N_9757,N_8348,N_8543);
nor U9758 (N_9758,N_8339,N_8348);
or U9759 (N_9759,N_8559,N_8097);
xor U9760 (N_9760,N_8893,N_8062);
or U9761 (N_9761,N_8984,N_8690);
nand U9762 (N_9762,N_8018,N_8670);
nor U9763 (N_9763,N_8357,N_8378);
or U9764 (N_9764,N_8415,N_8169);
or U9765 (N_9765,N_8192,N_8421);
nand U9766 (N_9766,N_8847,N_8783);
xor U9767 (N_9767,N_8159,N_8531);
nand U9768 (N_9768,N_8679,N_8851);
or U9769 (N_9769,N_8297,N_8612);
and U9770 (N_9770,N_8299,N_8117);
nand U9771 (N_9771,N_8774,N_8380);
or U9772 (N_9772,N_8476,N_8123);
nor U9773 (N_9773,N_8948,N_8240);
and U9774 (N_9774,N_8807,N_8060);
nor U9775 (N_9775,N_8991,N_8578);
xnor U9776 (N_9776,N_8347,N_8376);
and U9777 (N_9777,N_8956,N_8907);
and U9778 (N_9778,N_8625,N_8682);
xnor U9779 (N_9779,N_8003,N_8726);
xnor U9780 (N_9780,N_8646,N_8744);
nor U9781 (N_9781,N_8449,N_8248);
nor U9782 (N_9782,N_8888,N_8245);
xnor U9783 (N_9783,N_8330,N_8434);
nand U9784 (N_9784,N_8091,N_8743);
or U9785 (N_9785,N_8859,N_8900);
nand U9786 (N_9786,N_8010,N_8411);
and U9787 (N_9787,N_8629,N_8498);
nand U9788 (N_9788,N_8876,N_8333);
or U9789 (N_9789,N_8670,N_8039);
nand U9790 (N_9790,N_8023,N_8617);
nand U9791 (N_9791,N_8350,N_8039);
nand U9792 (N_9792,N_8821,N_8029);
and U9793 (N_9793,N_8194,N_8344);
nor U9794 (N_9794,N_8987,N_8466);
nand U9795 (N_9795,N_8212,N_8871);
nand U9796 (N_9796,N_8161,N_8405);
or U9797 (N_9797,N_8665,N_8145);
and U9798 (N_9798,N_8998,N_8112);
nor U9799 (N_9799,N_8154,N_8252);
or U9800 (N_9800,N_8988,N_8468);
and U9801 (N_9801,N_8794,N_8484);
nor U9802 (N_9802,N_8884,N_8052);
xnor U9803 (N_9803,N_8524,N_8536);
or U9804 (N_9804,N_8875,N_8401);
nor U9805 (N_9805,N_8344,N_8988);
and U9806 (N_9806,N_8671,N_8944);
or U9807 (N_9807,N_8364,N_8363);
or U9808 (N_9808,N_8878,N_8166);
nor U9809 (N_9809,N_8863,N_8829);
and U9810 (N_9810,N_8691,N_8005);
or U9811 (N_9811,N_8241,N_8982);
nor U9812 (N_9812,N_8815,N_8928);
nand U9813 (N_9813,N_8953,N_8331);
and U9814 (N_9814,N_8237,N_8650);
and U9815 (N_9815,N_8959,N_8390);
nor U9816 (N_9816,N_8863,N_8445);
and U9817 (N_9817,N_8158,N_8737);
and U9818 (N_9818,N_8421,N_8395);
and U9819 (N_9819,N_8796,N_8428);
and U9820 (N_9820,N_8564,N_8835);
nor U9821 (N_9821,N_8947,N_8641);
nand U9822 (N_9822,N_8676,N_8900);
or U9823 (N_9823,N_8090,N_8309);
or U9824 (N_9824,N_8753,N_8007);
nand U9825 (N_9825,N_8957,N_8979);
nand U9826 (N_9826,N_8009,N_8520);
or U9827 (N_9827,N_8340,N_8912);
nor U9828 (N_9828,N_8202,N_8891);
and U9829 (N_9829,N_8817,N_8933);
and U9830 (N_9830,N_8524,N_8661);
or U9831 (N_9831,N_8228,N_8964);
and U9832 (N_9832,N_8717,N_8368);
nand U9833 (N_9833,N_8403,N_8815);
or U9834 (N_9834,N_8234,N_8142);
and U9835 (N_9835,N_8011,N_8524);
nor U9836 (N_9836,N_8966,N_8253);
nand U9837 (N_9837,N_8104,N_8726);
nand U9838 (N_9838,N_8630,N_8703);
and U9839 (N_9839,N_8536,N_8118);
nor U9840 (N_9840,N_8691,N_8017);
or U9841 (N_9841,N_8395,N_8281);
and U9842 (N_9842,N_8846,N_8864);
or U9843 (N_9843,N_8529,N_8104);
or U9844 (N_9844,N_8389,N_8319);
and U9845 (N_9845,N_8522,N_8685);
and U9846 (N_9846,N_8293,N_8025);
or U9847 (N_9847,N_8551,N_8318);
nand U9848 (N_9848,N_8598,N_8430);
and U9849 (N_9849,N_8677,N_8381);
and U9850 (N_9850,N_8027,N_8564);
and U9851 (N_9851,N_8638,N_8957);
or U9852 (N_9852,N_8319,N_8253);
xnor U9853 (N_9853,N_8667,N_8281);
nor U9854 (N_9854,N_8827,N_8900);
nand U9855 (N_9855,N_8196,N_8947);
nand U9856 (N_9856,N_8639,N_8386);
or U9857 (N_9857,N_8862,N_8511);
nand U9858 (N_9858,N_8603,N_8351);
and U9859 (N_9859,N_8131,N_8331);
nor U9860 (N_9860,N_8412,N_8999);
and U9861 (N_9861,N_8639,N_8388);
nand U9862 (N_9862,N_8276,N_8230);
nand U9863 (N_9863,N_8338,N_8578);
xor U9864 (N_9864,N_8977,N_8361);
nor U9865 (N_9865,N_8765,N_8099);
nor U9866 (N_9866,N_8802,N_8400);
or U9867 (N_9867,N_8004,N_8568);
and U9868 (N_9868,N_8264,N_8043);
or U9869 (N_9869,N_8256,N_8064);
nand U9870 (N_9870,N_8663,N_8228);
and U9871 (N_9871,N_8549,N_8751);
nand U9872 (N_9872,N_8545,N_8156);
and U9873 (N_9873,N_8025,N_8831);
or U9874 (N_9874,N_8701,N_8002);
xnor U9875 (N_9875,N_8502,N_8655);
and U9876 (N_9876,N_8796,N_8669);
or U9877 (N_9877,N_8711,N_8171);
and U9878 (N_9878,N_8640,N_8106);
and U9879 (N_9879,N_8247,N_8245);
nor U9880 (N_9880,N_8755,N_8963);
nand U9881 (N_9881,N_8926,N_8792);
or U9882 (N_9882,N_8393,N_8836);
or U9883 (N_9883,N_8921,N_8786);
nand U9884 (N_9884,N_8808,N_8227);
nor U9885 (N_9885,N_8378,N_8627);
and U9886 (N_9886,N_8188,N_8790);
or U9887 (N_9887,N_8235,N_8452);
nor U9888 (N_9888,N_8187,N_8327);
nand U9889 (N_9889,N_8574,N_8947);
nand U9890 (N_9890,N_8332,N_8143);
and U9891 (N_9891,N_8038,N_8842);
or U9892 (N_9892,N_8625,N_8363);
or U9893 (N_9893,N_8834,N_8020);
and U9894 (N_9894,N_8188,N_8354);
nor U9895 (N_9895,N_8206,N_8984);
nor U9896 (N_9896,N_8813,N_8433);
or U9897 (N_9897,N_8479,N_8345);
or U9898 (N_9898,N_8409,N_8073);
nor U9899 (N_9899,N_8798,N_8519);
nand U9900 (N_9900,N_8621,N_8200);
or U9901 (N_9901,N_8792,N_8509);
and U9902 (N_9902,N_8242,N_8031);
and U9903 (N_9903,N_8756,N_8426);
or U9904 (N_9904,N_8628,N_8886);
nand U9905 (N_9905,N_8944,N_8307);
nor U9906 (N_9906,N_8339,N_8916);
and U9907 (N_9907,N_8802,N_8219);
nor U9908 (N_9908,N_8503,N_8776);
nand U9909 (N_9909,N_8698,N_8934);
and U9910 (N_9910,N_8674,N_8750);
and U9911 (N_9911,N_8081,N_8524);
nor U9912 (N_9912,N_8851,N_8258);
nor U9913 (N_9913,N_8732,N_8095);
and U9914 (N_9914,N_8621,N_8551);
or U9915 (N_9915,N_8482,N_8220);
nand U9916 (N_9916,N_8211,N_8901);
nand U9917 (N_9917,N_8205,N_8970);
nor U9918 (N_9918,N_8713,N_8273);
xor U9919 (N_9919,N_8614,N_8549);
and U9920 (N_9920,N_8776,N_8668);
nor U9921 (N_9921,N_8030,N_8864);
and U9922 (N_9922,N_8873,N_8322);
nor U9923 (N_9923,N_8091,N_8000);
nand U9924 (N_9924,N_8621,N_8458);
nand U9925 (N_9925,N_8038,N_8763);
nor U9926 (N_9926,N_8941,N_8304);
nand U9927 (N_9927,N_8461,N_8375);
and U9928 (N_9928,N_8999,N_8869);
nor U9929 (N_9929,N_8191,N_8594);
and U9930 (N_9930,N_8666,N_8515);
or U9931 (N_9931,N_8099,N_8723);
and U9932 (N_9932,N_8609,N_8729);
or U9933 (N_9933,N_8297,N_8726);
nand U9934 (N_9934,N_8078,N_8230);
nand U9935 (N_9935,N_8486,N_8067);
nor U9936 (N_9936,N_8072,N_8786);
and U9937 (N_9937,N_8512,N_8910);
and U9938 (N_9938,N_8534,N_8600);
or U9939 (N_9939,N_8963,N_8354);
and U9940 (N_9940,N_8198,N_8800);
nand U9941 (N_9941,N_8142,N_8438);
nor U9942 (N_9942,N_8920,N_8664);
nor U9943 (N_9943,N_8052,N_8681);
nand U9944 (N_9944,N_8324,N_8483);
and U9945 (N_9945,N_8721,N_8975);
nand U9946 (N_9946,N_8534,N_8299);
and U9947 (N_9947,N_8341,N_8077);
nor U9948 (N_9948,N_8418,N_8676);
and U9949 (N_9949,N_8942,N_8608);
and U9950 (N_9950,N_8815,N_8615);
nor U9951 (N_9951,N_8820,N_8545);
nor U9952 (N_9952,N_8046,N_8738);
and U9953 (N_9953,N_8676,N_8242);
nor U9954 (N_9954,N_8008,N_8358);
nor U9955 (N_9955,N_8258,N_8454);
nand U9956 (N_9956,N_8280,N_8420);
and U9957 (N_9957,N_8193,N_8175);
xnor U9958 (N_9958,N_8131,N_8655);
or U9959 (N_9959,N_8411,N_8374);
nand U9960 (N_9960,N_8662,N_8538);
nor U9961 (N_9961,N_8115,N_8763);
xnor U9962 (N_9962,N_8375,N_8565);
or U9963 (N_9963,N_8020,N_8646);
nand U9964 (N_9964,N_8443,N_8819);
and U9965 (N_9965,N_8307,N_8806);
or U9966 (N_9966,N_8508,N_8216);
nor U9967 (N_9967,N_8227,N_8740);
nor U9968 (N_9968,N_8008,N_8364);
or U9969 (N_9969,N_8802,N_8741);
and U9970 (N_9970,N_8516,N_8555);
or U9971 (N_9971,N_8580,N_8383);
and U9972 (N_9972,N_8683,N_8893);
or U9973 (N_9973,N_8253,N_8218);
and U9974 (N_9974,N_8625,N_8694);
nor U9975 (N_9975,N_8124,N_8103);
nand U9976 (N_9976,N_8076,N_8394);
nand U9977 (N_9977,N_8749,N_8310);
nand U9978 (N_9978,N_8574,N_8524);
and U9979 (N_9979,N_8158,N_8810);
or U9980 (N_9980,N_8997,N_8209);
or U9981 (N_9981,N_8174,N_8551);
or U9982 (N_9982,N_8078,N_8171);
nor U9983 (N_9983,N_8100,N_8200);
nor U9984 (N_9984,N_8807,N_8030);
nand U9985 (N_9985,N_8720,N_8621);
nand U9986 (N_9986,N_8320,N_8974);
nor U9987 (N_9987,N_8555,N_8628);
nor U9988 (N_9988,N_8192,N_8163);
or U9989 (N_9989,N_8079,N_8734);
and U9990 (N_9990,N_8762,N_8537);
and U9991 (N_9991,N_8988,N_8305);
or U9992 (N_9992,N_8581,N_8573);
or U9993 (N_9993,N_8860,N_8171);
nor U9994 (N_9994,N_8662,N_8856);
nor U9995 (N_9995,N_8335,N_8409);
nand U9996 (N_9996,N_8178,N_8244);
nand U9997 (N_9997,N_8259,N_8144);
nor U9998 (N_9998,N_8973,N_8866);
nor U9999 (N_9999,N_8825,N_8728);
and UO_0 (O_0,N_9023,N_9344);
or UO_1 (O_1,N_9405,N_9500);
or UO_2 (O_2,N_9640,N_9190);
nand UO_3 (O_3,N_9379,N_9106);
nand UO_4 (O_4,N_9246,N_9769);
and UO_5 (O_5,N_9997,N_9943);
nand UO_6 (O_6,N_9755,N_9192);
or UO_7 (O_7,N_9313,N_9412);
and UO_8 (O_8,N_9267,N_9275);
or UO_9 (O_9,N_9522,N_9837);
nor UO_10 (O_10,N_9309,N_9579);
and UO_11 (O_11,N_9422,N_9633);
nor UO_12 (O_12,N_9988,N_9416);
nand UO_13 (O_13,N_9550,N_9558);
nand UO_14 (O_14,N_9661,N_9217);
nor UO_15 (O_15,N_9025,N_9229);
and UO_16 (O_16,N_9816,N_9084);
nand UO_17 (O_17,N_9095,N_9950);
nand UO_18 (O_18,N_9101,N_9610);
and UO_19 (O_19,N_9375,N_9711);
and UO_20 (O_20,N_9506,N_9480);
nand UO_21 (O_21,N_9647,N_9776);
nor UO_22 (O_22,N_9089,N_9280);
and UO_23 (O_23,N_9790,N_9669);
and UO_24 (O_24,N_9105,N_9597);
xnor UO_25 (O_25,N_9334,N_9922);
nor UO_26 (O_26,N_9858,N_9665);
nor UO_27 (O_27,N_9678,N_9593);
and UO_28 (O_28,N_9842,N_9866);
and UO_29 (O_29,N_9384,N_9469);
nor UO_30 (O_30,N_9450,N_9975);
and UO_31 (O_31,N_9195,N_9814);
and UO_32 (O_32,N_9960,N_9463);
nor UO_33 (O_33,N_9607,N_9944);
and UO_34 (O_34,N_9555,N_9887);
and UO_35 (O_35,N_9478,N_9079);
nor UO_36 (O_36,N_9525,N_9492);
and UO_37 (O_37,N_9371,N_9205);
nand UO_38 (O_38,N_9342,N_9382);
nand UO_39 (O_39,N_9533,N_9928);
and UO_40 (O_40,N_9904,N_9452);
nand UO_41 (O_41,N_9426,N_9763);
nor UO_42 (O_42,N_9850,N_9263);
or UO_43 (O_43,N_9973,N_9630);
and UO_44 (O_44,N_9157,N_9886);
and UO_45 (O_45,N_9148,N_9113);
nor UO_46 (O_46,N_9750,N_9815);
nor UO_47 (O_47,N_9176,N_9325);
nor UO_48 (O_48,N_9540,N_9649);
or UO_49 (O_49,N_9241,N_9038);
or UO_50 (O_50,N_9707,N_9938);
and UO_51 (O_51,N_9662,N_9874);
or UO_52 (O_52,N_9486,N_9511);
nand UO_53 (O_53,N_9543,N_9393);
nand UO_54 (O_54,N_9715,N_9727);
nand UO_55 (O_55,N_9618,N_9413);
or UO_56 (O_56,N_9085,N_9681);
xnor UO_57 (O_57,N_9799,N_9590);
or UO_58 (O_58,N_9078,N_9933);
or UO_59 (O_59,N_9531,N_9884);
nand UO_60 (O_60,N_9166,N_9392);
nor UO_61 (O_61,N_9920,N_9692);
nand UO_62 (O_62,N_9901,N_9453);
or UO_63 (O_63,N_9722,N_9602);
nand UO_64 (O_64,N_9057,N_9521);
nand UO_65 (O_65,N_9729,N_9349);
nand UO_66 (O_66,N_9826,N_9179);
or UO_67 (O_67,N_9357,N_9910);
nor UO_68 (O_68,N_9080,N_9804);
and UO_69 (O_69,N_9774,N_9093);
nor UO_70 (O_70,N_9249,N_9970);
nor UO_71 (O_71,N_9472,N_9096);
nor UO_72 (O_72,N_9073,N_9706);
or UO_73 (O_73,N_9206,N_9447);
nor UO_74 (O_74,N_9359,N_9165);
nor UO_75 (O_75,N_9367,N_9738);
or UO_76 (O_76,N_9351,N_9830);
and UO_77 (O_77,N_9848,N_9098);
and UO_78 (O_78,N_9471,N_9339);
nand UO_79 (O_79,N_9264,N_9028);
and UO_80 (O_80,N_9926,N_9369);
and UO_81 (O_81,N_9908,N_9578);
nand UO_82 (O_82,N_9230,N_9104);
or UO_83 (O_83,N_9658,N_9575);
nor UO_84 (O_84,N_9406,N_9968);
or UO_85 (O_85,N_9680,N_9508);
nor UO_86 (O_86,N_9451,N_9321);
or UO_87 (O_87,N_9236,N_9697);
or UO_88 (O_88,N_9861,N_9324);
nor UO_89 (O_89,N_9732,N_9783);
nand UO_90 (O_90,N_9231,N_9601);
or UO_91 (O_91,N_9168,N_9978);
nand UO_92 (O_92,N_9801,N_9062);
and UO_93 (O_93,N_9636,N_9880);
nor UO_94 (O_94,N_9121,N_9298);
nand UO_95 (O_95,N_9833,N_9855);
xnor UO_96 (O_96,N_9477,N_9110);
nand UO_97 (O_97,N_9704,N_9523);
nand UO_98 (O_98,N_9122,N_9891);
and UO_99 (O_99,N_9224,N_9254);
nor UO_100 (O_100,N_9075,N_9137);
nand UO_101 (O_101,N_9401,N_9262);
and UO_102 (O_102,N_9112,N_9840);
or UO_103 (O_103,N_9204,N_9541);
nand UO_104 (O_104,N_9355,N_9823);
nand UO_105 (O_105,N_9900,N_9788);
xor UO_106 (O_106,N_9552,N_9741);
nor UO_107 (O_107,N_9791,N_9146);
nor UO_108 (O_108,N_9239,N_9169);
nand UO_109 (O_109,N_9036,N_9035);
nand UO_110 (O_110,N_9197,N_9644);
nand UO_111 (O_111,N_9818,N_9949);
nor UO_112 (O_112,N_9210,N_9460);
or UO_113 (O_113,N_9536,N_9825);
and UO_114 (O_114,N_9553,N_9809);
or UO_115 (O_115,N_9088,N_9177);
and UO_116 (O_116,N_9772,N_9445);
and UO_117 (O_117,N_9048,N_9620);
or UO_118 (O_118,N_9466,N_9753);
nand UO_119 (O_119,N_9985,N_9131);
nand UO_120 (O_120,N_9304,N_9526);
nand UO_121 (O_121,N_9333,N_9650);
nor UO_122 (O_122,N_9399,N_9227);
and UO_123 (O_123,N_9097,N_9864);
nor UO_124 (O_124,N_9293,N_9296);
nand UO_125 (O_125,N_9652,N_9058);
and UO_126 (O_126,N_9017,N_9063);
xnor UO_127 (O_127,N_9198,N_9588);
or UO_128 (O_128,N_9468,N_9042);
nand UO_129 (O_129,N_9921,N_9076);
and UO_130 (O_130,N_9128,N_9568);
xnor UO_131 (O_131,N_9797,N_9530);
or UO_132 (O_132,N_9504,N_9292);
and UO_133 (O_133,N_9002,N_9178);
or UO_134 (O_134,N_9667,N_9152);
and UO_135 (O_135,N_9449,N_9418);
or UO_136 (O_136,N_9821,N_9118);
and UO_137 (O_137,N_9643,N_9311);
or UO_138 (O_138,N_9872,N_9346);
nand UO_139 (O_139,N_9135,N_9976);
and UO_140 (O_140,N_9429,N_9488);
and UO_141 (O_141,N_9679,N_9686);
and UO_142 (O_142,N_9415,N_9362);
nor UO_143 (O_143,N_9951,N_9109);
and UO_144 (O_144,N_9745,N_9690);
and UO_145 (O_145,N_9688,N_9993);
nand UO_146 (O_146,N_9796,N_9187);
nor UO_147 (O_147,N_9592,N_9102);
nand UO_148 (O_148,N_9059,N_9759);
and UO_149 (O_149,N_9441,N_9605);
or UO_150 (O_150,N_9044,N_9744);
or UO_151 (O_151,N_9201,N_9594);
nor UO_152 (O_152,N_9424,N_9077);
xnor UO_153 (O_153,N_9845,N_9743);
nand UO_154 (O_154,N_9243,N_9974);
and UO_155 (O_155,N_9302,N_9386);
and UO_156 (O_156,N_9829,N_9794);
or UO_157 (O_157,N_9972,N_9461);
nand UO_158 (O_158,N_9454,N_9871);
and UO_159 (O_159,N_9383,N_9895);
or UO_160 (O_160,N_9655,N_9014);
nor UO_161 (O_161,N_9162,N_9233);
or UO_162 (O_162,N_9863,N_9639);
nor UO_163 (O_163,N_9223,N_9024);
or UO_164 (O_164,N_9033,N_9070);
nand UO_165 (O_165,N_9853,N_9475);
and UO_166 (O_166,N_9585,N_9115);
nor UO_167 (O_167,N_9225,N_9251);
and UO_168 (O_168,N_9403,N_9586);
or UO_169 (O_169,N_9410,N_9494);
nand UO_170 (O_170,N_9072,N_9006);
nor UO_171 (O_171,N_9474,N_9003);
and UO_172 (O_172,N_9625,N_9203);
nand UO_173 (O_173,N_9981,N_9685);
nor UO_174 (O_174,N_9544,N_9503);
nor UO_175 (O_175,N_9828,N_9687);
or UO_176 (O_176,N_9125,N_9498);
nand UO_177 (O_177,N_9491,N_9221);
nand UO_178 (O_178,N_9222,N_9709);
nand UO_179 (O_179,N_9979,N_9465);
nand UO_180 (O_180,N_9473,N_9082);
or UO_181 (O_181,N_9385,N_9303);
nor UO_182 (O_182,N_9623,N_9752);
or UO_183 (O_183,N_9443,N_9932);
xnor UO_184 (O_184,N_9562,N_9305);
nor UO_185 (O_185,N_9020,N_9720);
or UO_186 (O_186,N_9153,N_9893);
nand UO_187 (O_187,N_9778,N_9701);
nor UO_188 (O_188,N_9318,N_9297);
or UO_189 (O_189,N_9582,N_9402);
or UO_190 (O_190,N_9785,N_9260);
or UO_191 (O_191,N_9616,N_9635);
nand UO_192 (O_192,N_9631,N_9634);
nor UO_193 (O_193,N_9434,N_9328);
nand UO_194 (O_194,N_9323,N_9497);
nor UO_195 (O_195,N_9992,N_9677);
nand UO_196 (O_196,N_9695,N_9749);
nor UO_197 (O_197,N_9945,N_9648);
or UO_198 (O_198,N_9326,N_9322);
nand UO_199 (O_199,N_9138,N_9409);
or UO_200 (O_200,N_9708,N_9388);
nor UO_201 (O_201,N_9606,N_9805);
and UO_202 (O_202,N_9617,N_9366);
xnor UO_203 (O_203,N_9865,N_9438);
nand UO_204 (O_204,N_9567,N_9545);
nand UO_205 (O_205,N_9282,N_9551);
nand UO_206 (O_206,N_9219,N_9032);
nor UO_207 (O_207,N_9923,N_9261);
and UO_208 (O_208,N_9614,N_9611);
and UO_209 (O_209,N_9030,N_9045);
nand UO_210 (O_210,N_9247,N_9040);
or UO_211 (O_211,N_9969,N_9966);
and UO_212 (O_212,N_9439,N_9398);
nand UO_213 (O_213,N_9564,N_9760);
or UO_214 (O_214,N_9358,N_9250);
nor UO_215 (O_215,N_9719,N_9565);
or UO_216 (O_216,N_9561,N_9228);
nor UO_217 (O_217,N_9820,N_9627);
nand UO_218 (O_218,N_9052,N_9394);
and UO_219 (O_219,N_9535,N_9289);
nor UO_220 (O_220,N_9589,N_9888);
nand UO_221 (O_221,N_9184,N_9598);
or UO_222 (O_222,N_9761,N_9869);
or UO_223 (O_223,N_9400,N_9381);
nor UO_224 (O_224,N_9834,N_9780);
or UO_225 (O_225,N_9812,N_9638);
or UO_226 (O_226,N_9983,N_9090);
nand UO_227 (O_227,N_9717,N_9411);
nor UO_228 (O_228,N_9004,N_9144);
nand UO_229 (O_229,N_9907,N_9516);
or UO_230 (O_230,N_9257,N_9918);
nand UO_231 (O_231,N_9576,N_9307);
nor UO_232 (O_232,N_9877,N_9034);
and UO_233 (O_233,N_9064,N_9986);
or UO_234 (O_234,N_9609,N_9518);
nand UO_235 (O_235,N_9114,N_9671);
nand UO_236 (O_236,N_9885,N_9327);
nor UO_237 (O_237,N_9245,N_9906);
or UO_238 (O_238,N_9710,N_9193);
nand UO_239 (O_239,N_9811,N_9622);
or UO_240 (O_240,N_9031,N_9237);
nor UO_241 (O_241,N_9124,N_9255);
or UO_242 (O_242,N_9786,N_9879);
or UO_243 (O_243,N_9947,N_9273);
and UO_244 (O_244,N_9501,N_9599);
nor UO_245 (O_245,N_9442,N_9682);
nand UO_246 (O_246,N_9942,N_9314);
and UO_247 (O_247,N_9462,N_9141);
nand UO_248 (O_248,N_9768,N_9207);
or UO_249 (O_249,N_9621,N_9499);
nor UO_250 (O_250,N_9773,N_9538);
and UO_251 (O_251,N_9813,N_9420);
nor UO_252 (O_252,N_9554,N_9889);
nand UO_253 (O_253,N_9764,N_9962);
nor UO_254 (O_254,N_9862,N_9702);
nor UO_255 (O_255,N_9288,N_9946);
nor UO_256 (O_256,N_9642,N_9963);
nor UO_257 (O_257,N_9183,N_9977);
and UO_258 (O_258,N_9742,N_9464);
nor UO_259 (O_259,N_9345,N_9703);
nor UO_260 (O_260,N_9698,N_9924);
nor UO_261 (O_261,N_9276,N_9580);
or UO_262 (O_262,N_9931,N_9330);
nand UO_263 (O_263,N_9007,N_9286);
and UO_264 (O_264,N_9151,N_9196);
nand UO_265 (O_265,N_9091,N_9363);
and UO_266 (O_266,N_9479,N_9507);
and UO_267 (O_267,N_9374,N_9641);
and UO_268 (O_268,N_9242,N_9542);
nor UO_269 (O_269,N_9068,N_9739);
and UO_270 (O_270,N_9147,N_9890);
or UO_271 (O_271,N_9191,N_9170);
nand UO_272 (O_272,N_9336,N_9365);
and UO_273 (O_273,N_9684,N_9515);
or UO_274 (O_274,N_9039,N_9046);
or UO_275 (O_275,N_9290,N_9514);
and UO_276 (O_276,N_9612,N_9537);
xor UO_277 (O_277,N_9991,N_9127);
and UO_278 (O_278,N_9637,N_9407);
and UO_279 (O_279,N_9019,N_9512);
nand UO_280 (O_280,N_9496,N_9390);
nand UO_281 (O_281,N_9347,N_9935);
nor UO_282 (O_282,N_9746,N_9911);
or UO_283 (O_283,N_9111,N_9934);
or UO_284 (O_284,N_9283,N_9689);
nand UO_285 (O_285,N_9481,N_9332);
nand UO_286 (O_286,N_9832,N_9150);
or UO_287 (O_287,N_9457,N_9356);
and UO_288 (O_288,N_9967,N_9748);
and UO_289 (O_289,N_9489,N_9524);
and UO_290 (O_290,N_9186,N_9806);
nand UO_291 (O_291,N_9999,N_9431);
and UO_292 (O_292,N_9574,N_9490);
or UO_293 (O_293,N_9435,N_9939);
and UO_294 (O_294,N_9802,N_9675);
or UO_295 (O_295,N_9725,N_9259);
and UO_296 (O_296,N_9808,N_9256);
or UO_297 (O_297,N_9757,N_9714);
nor UO_298 (O_298,N_9881,N_9027);
or UO_299 (O_299,N_9726,N_9800);
nand UO_300 (O_300,N_9632,N_9716);
nor UO_301 (O_301,N_9265,N_9335);
nor UO_302 (O_302,N_9244,N_9312);
and UO_303 (O_303,N_9069,N_9484);
nand UO_304 (O_304,N_9957,N_9149);
or UO_305 (O_305,N_9787,N_9408);
and UO_306 (O_306,N_9958,N_9291);
nor UO_307 (O_307,N_9056,N_9160);
xnor UO_308 (O_308,N_9470,N_9629);
or UO_309 (O_309,N_9456,N_9839);
nand UO_310 (O_310,N_9458,N_9646);
and UO_311 (O_311,N_9734,N_9827);
nor UO_312 (O_312,N_9654,N_9546);
and UO_313 (O_313,N_9316,N_9132);
and UO_314 (O_314,N_9389,N_9860);
or UO_315 (O_315,N_9691,N_9026);
nor UO_316 (O_316,N_9437,N_9446);
and UO_317 (O_317,N_9560,N_9831);
nor UO_318 (O_318,N_9696,N_9964);
xnor UO_319 (O_319,N_9735,N_9119);
nand UO_320 (O_320,N_9436,N_9174);
nor UO_321 (O_321,N_9754,N_9216);
nand UO_322 (O_322,N_9199,N_9041);
xnor UO_323 (O_323,N_9455,N_9817);
and UO_324 (O_324,N_9919,N_9235);
nand UO_325 (O_325,N_9844,N_9664);
and UO_326 (O_326,N_9182,N_9253);
and UO_327 (O_327,N_9859,N_9914);
nand UO_328 (O_328,N_9737,N_9306);
nand UO_329 (O_329,N_9171,N_9836);
nor UO_330 (O_330,N_9854,N_9092);
nor UO_331 (O_331,N_9232,N_9099);
nor UO_332 (O_332,N_9329,N_9194);
nor UO_333 (O_333,N_9271,N_9378);
xor UO_334 (O_334,N_9857,N_9338);
nor UO_335 (O_335,N_9867,N_9021);
nor UO_336 (O_336,N_9941,N_9397);
nor UO_337 (O_337,N_9838,N_9081);
and UO_338 (O_338,N_9142,N_9573);
or UO_339 (O_339,N_9459,N_9188);
nor UO_340 (O_340,N_9534,N_9651);
or UO_341 (O_341,N_9736,N_9810);
or UO_342 (O_342,N_9668,N_9584);
and UO_343 (O_343,N_9718,N_9209);
or UO_344 (O_344,N_9427,N_9930);
nor UO_345 (O_345,N_9730,N_9071);
or UO_346 (O_346,N_9348,N_9285);
nand UO_347 (O_347,N_9485,N_9495);
nor UO_348 (O_348,N_9909,N_9894);
nor UO_349 (O_349,N_9164,N_9172);
or UO_350 (O_350,N_9672,N_9956);
nor UO_351 (O_351,N_9547,N_9372);
nor UO_352 (O_352,N_9238,N_9912);
and UO_353 (O_353,N_9361,N_9699);
and UO_354 (O_354,N_9126,N_9683);
and UO_355 (O_355,N_9782,N_9936);
and UO_356 (O_356,N_9843,N_9980);
nor UO_357 (O_357,N_9117,N_9915);
and UO_358 (O_358,N_9012,N_9892);
and UO_359 (O_359,N_9493,N_9143);
nand UO_360 (O_360,N_9566,N_9583);
and UO_361 (O_361,N_9154,N_9903);
nand UO_362 (O_362,N_9331,N_9156);
xor UO_363 (O_363,N_9781,N_9532);
nor UO_364 (O_364,N_9758,N_9295);
and UO_365 (O_365,N_9234,N_9954);
nand UO_366 (O_366,N_9299,N_9433);
or UO_367 (O_367,N_9878,N_9281);
and UO_368 (O_368,N_9569,N_9423);
or UO_369 (O_369,N_9873,N_9368);
or UO_370 (O_370,N_9220,N_9161);
nor UO_371 (O_371,N_9315,N_9279);
or UO_372 (O_372,N_9103,N_9659);
or UO_373 (O_373,N_9807,N_9548);
nand UO_374 (O_374,N_9929,N_9376);
nor UO_375 (O_375,N_9100,N_9430);
nor UO_376 (O_376,N_9123,N_9882);
or UO_377 (O_377,N_9483,N_9337);
or UO_378 (O_378,N_9913,N_9795);
or UO_379 (O_379,N_9563,N_9428);
nor UO_380 (O_380,N_9784,N_9916);
nand UO_381 (O_381,N_9268,N_9513);
and UO_382 (O_382,N_9301,N_9693);
and UO_383 (O_383,N_9824,N_9868);
and UO_384 (O_384,N_9343,N_9953);
nor UO_385 (O_385,N_9107,N_9883);
or UO_386 (O_386,N_9529,N_9215);
nor UO_387 (O_387,N_9572,N_9159);
nor UO_388 (O_388,N_9937,N_9364);
nand UO_389 (O_389,N_9779,N_9340);
nor UO_390 (O_390,N_9984,N_9419);
and UO_391 (O_391,N_9517,N_9798);
or UO_392 (O_392,N_9440,N_9140);
xnor UO_393 (O_393,N_9060,N_9875);
or UO_394 (O_394,N_9663,N_9694);
xor UO_395 (O_395,N_9009,N_9425);
xor UO_396 (O_396,N_9700,N_9214);
and UO_397 (O_397,N_9835,N_9065);
xnor UO_398 (O_398,N_9766,N_9284);
nand UO_399 (O_399,N_9723,N_9628);
nor UO_400 (O_400,N_9982,N_9948);
xor UO_401 (O_401,N_9917,N_9448);
or UO_402 (O_402,N_9341,N_9008);
and UO_403 (O_403,N_9061,N_9352);
and UO_404 (O_404,N_9851,N_9721);
nand UO_405 (O_405,N_9300,N_9167);
or UO_406 (O_406,N_9899,N_9670);
nor UO_407 (O_407,N_9136,N_9556);
nor UO_408 (O_408,N_9660,N_9175);
nor UO_409 (O_409,N_9226,N_9591);
nor UO_410 (O_410,N_9849,N_9527);
nand UO_411 (O_411,N_9971,N_9756);
and UO_412 (O_412,N_9876,N_9615);
nor UO_413 (O_413,N_9989,N_9116);
xor UO_414 (O_414,N_9898,N_9391);
nor UO_415 (O_415,N_9212,N_9319);
and UO_416 (O_416,N_9505,N_9603);
nand UO_417 (O_417,N_9240,N_9596);
or UO_418 (O_418,N_9277,N_9108);
nor UO_419 (O_419,N_9417,N_9010);
or UO_420 (O_420,N_9404,N_9139);
nor UO_421 (O_421,N_9130,N_9770);
and UO_422 (O_422,N_9444,N_9018);
or UO_423 (O_423,N_9539,N_9927);
and UO_424 (O_424,N_9145,N_9278);
and UO_425 (O_425,N_9666,N_9673);
or UO_426 (O_426,N_9751,N_9998);
nand UO_427 (O_427,N_9803,N_9896);
nand UO_428 (O_428,N_9731,N_9747);
and UO_429 (O_429,N_9373,N_9120);
xnor UO_430 (O_430,N_9414,N_9952);
nor UO_431 (O_431,N_9158,N_9762);
and UO_432 (O_432,N_9476,N_9252);
and UO_433 (O_433,N_9266,N_9509);
nand UO_434 (O_434,N_9767,N_9467);
nand UO_435 (O_435,N_9287,N_9377);
and UO_436 (O_436,N_9571,N_9789);
nand UO_437 (O_437,N_9841,N_9847);
nand UO_438 (O_438,N_9487,N_9990);
and UO_439 (O_439,N_9705,N_9185);
nand UO_440 (O_440,N_9712,N_9624);
or UO_441 (O_441,N_9370,N_9846);
xor UO_442 (O_442,N_9856,N_9902);
or UO_443 (O_443,N_9519,N_9765);
or UO_444 (O_444,N_9005,N_9029);
nand UO_445 (O_445,N_9066,N_9000);
or UO_446 (O_446,N_9897,N_9054);
and UO_447 (O_447,N_9218,N_9955);
nand UO_448 (O_448,N_9520,N_9961);
or UO_449 (O_449,N_9353,N_9987);
and UO_450 (O_450,N_9208,N_9996);
nor UO_451 (O_451,N_9270,N_9350);
xor UO_452 (O_452,N_9055,N_9053);
nor UO_453 (O_453,N_9482,N_9549);
nand UO_454 (O_454,N_9294,N_9272);
and UO_455 (O_455,N_9308,N_9994);
nand UO_456 (O_456,N_9380,N_9676);
and UO_457 (O_457,N_9733,N_9587);
or UO_458 (O_458,N_9310,N_9740);
nor UO_459 (O_459,N_9870,N_9015);
or UO_460 (O_460,N_9129,N_9777);
nand UO_461 (O_461,N_9793,N_9570);
or UO_462 (O_462,N_9094,N_9395);
or UO_463 (O_463,N_9925,N_9771);
and UO_464 (O_464,N_9248,N_9134);
and UO_465 (O_465,N_9626,N_9940);
and UO_466 (O_466,N_9087,N_9905);
nand UO_467 (O_467,N_9724,N_9822);
or UO_468 (O_468,N_9581,N_9200);
nor UO_469 (O_469,N_9074,N_9595);
nor UO_470 (O_470,N_9713,N_9163);
and UO_471 (O_471,N_9421,N_9317);
nand UO_472 (O_472,N_9645,N_9001);
nand UO_473 (O_473,N_9396,N_9959);
nand UO_474 (O_474,N_9360,N_9155);
nand UO_475 (O_475,N_9604,N_9037);
or UO_476 (O_476,N_9067,N_9728);
nor UO_477 (O_477,N_9173,N_9354);
and UO_478 (O_478,N_9608,N_9653);
or UO_479 (O_479,N_9502,N_9011);
nand UO_480 (O_480,N_9202,N_9852);
nand UO_481 (O_481,N_9387,N_9613);
or UO_482 (O_482,N_9086,N_9320);
or UO_483 (O_483,N_9189,N_9049);
nor UO_484 (O_484,N_9269,N_9657);
nor UO_485 (O_485,N_9559,N_9016);
and UO_486 (O_486,N_9181,N_9022);
nor UO_487 (O_487,N_9432,N_9180);
nand UO_488 (O_488,N_9528,N_9274);
nor UO_489 (O_489,N_9043,N_9213);
nor UO_490 (O_490,N_9258,N_9577);
and UO_491 (O_491,N_9819,N_9995);
nand UO_492 (O_492,N_9775,N_9965);
and UO_493 (O_493,N_9013,N_9557);
nand UO_494 (O_494,N_9083,N_9656);
and UO_495 (O_495,N_9600,N_9674);
nand UO_496 (O_496,N_9133,N_9792);
nand UO_497 (O_497,N_9510,N_9050);
and UO_498 (O_498,N_9619,N_9051);
nand UO_499 (O_499,N_9047,N_9211);
and UO_500 (O_500,N_9297,N_9423);
or UO_501 (O_501,N_9165,N_9953);
or UO_502 (O_502,N_9703,N_9182);
and UO_503 (O_503,N_9485,N_9152);
nand UO_504 (O_504,N_9860,N_9844);
nor UO_505 (O_505,N_9034,N_9398);
nor UO_506 (O_506,N_9216,N_9303);
and UO_507 (O_507,N_9430,N_9095);
or UO_508 (O_508,N_9877,N_9591);
nand UO_509 (O_509,N_9647,N_9385);
nor UO_510 (O_510,N_9184,N_9692);
nor UO_511 (O_511,N_9990,N_9371);
xor UO_512 (O_512,N_9734,N_9934);
nor UO_513 (O_513,N_9412,N_9638);
nor UO_514 (O_514,N_9357,N_9034);
nor UO_515 (O_515,N_9577,N_9802);
xor UO_516 (O_516,N_9629,N_9344);
nand UO_517 (O_517,N_9789,N_9046);
and UO_518 (O_518,N_9824,N_9755);
or UO_519 (O_519,N_9167,N_9596);
nand UO_520 (O_520,N_9074,N_9265);
or UO_521 (O_521,N_9209,N_9482);
or UO_522 (O_522,N_9671,N_9092);
nand UO_523 (O_523,N_9144,N_9708);
nor UO_524 (O_524,N_9884,N_9061);
and UO_525 (O_525,N_9646,N_9703);
and UO_526 (O_526,N_9597,N_9886);
nor UO_527 (O_527,N_9773,N_9625);
and UO_528 (O_528,N_9745,N_9116);
and UO_529 (O_529,N_9533,N_9024);
or UO_530 (O_530,N_9311,N_9107);
nand UO_531 (O_531,N_9699,N_9431);
and UO_532 (O_532,N_9209,N_9197);
and UO_533 (O_533,N_9997,N_9412);
xor UO_534 (O_534,N_9666,N_9745);
nor UO_535 (O_535,N_9649,N_9570);
or UO_536 (O_536,N_9660,N_9105);
nand UO_537 (O_537,N_9102,N_9316);
xor UO_538 (O_538,N_9126,N_9047);
or UO_539 (O_539,N_9796,N_9870);
nor UO_540 (O_540,N_9293,N_9331);
and UO_541 (O_541,N_9018,N_9546);
or UO_542 (O_542,N_9660,N_9983);
nand UO_543 (O_543,N_9487,N_9371);
nand UO_544 (O_544,N_9213,N_9230);
nor UO_545 (O_545,N_9385,N_9648);
and UO_546 (O_546,N_9868,N_9559);
and UO_547 (O_547,N_9972,N_9106);
or UO_548 (O_548,N_9949,N_9914);
nand UO_549 (O_549,N_9721,N_9577);
nand UO_550 (O_550,N_9531,N_9297);
or UO_551 (O_551,N_9019,N_9834);
nor UO_552 (O_552,N_9228,N_9287);
or UO_553 (O_553,N_9491,N_9040);
and UO_554 (O_554,N_9492,N_9550);
nand UO_555 (O_555,N_9528,N_9663);
nor UO_556 (O_556,N_9887,N_9955);
xor UO_557 (O_557,N_9934,N_9340);
and UO_558 (O_558,N_9945,N_9303);
nand UO_559 (O_559,N_9868,N_9969);
nor UO_560 (O_560,N_9916,N_9747);
nand UO_561 (O_561,N_9842,N_9181);
and UO_562 (O_562,N_9938,N_9918);
nor UO_563 (O_563,N_9018,N_9280);
nand UO_564 (O_564,N_9064,N_9615);
and UO_565 (O_565,N_9739,N_9696);
or UO_566 (O_566,N_9645,N_9902);
or UO_567 (O_567,N_9349,N_9314);
nand UO_568 (O_568,N_9242,N_9194);
nor UO_569 (O_569,N_9051,N_9694);
nand UO_570 (O_570,N_9237,N_9185);
nand UO_571 (O_571,N_9136,N_9502);
and UO_572 (O_572,N_9927,N_9482);
and UO_573 (O_573,N_9103,N_9733);
nand UO_574 (O_574,N_9292,N_9497);
and UO_575 (O_575,N_9156,N_9581);
or UO_576 (O_576,N_9781,N_9645);
nand UO_577 (O_577,N_9036,N_9874);
nand UO_578 (O_578,N_9329,N_9916);
nor UO_579 (O_579,N_9147,N_9103);
nand UO_580 (O_580,N_9898,N_9229);
and UO_581 (O_581,N_9858,N_9467);
or UO_582 (O_582,N_9337,N_9354);
and UO_583 (O_583,N_9679,N_9715);
and UO_584 (O_584,N_9574,N_9831);
nor UO_585 (O_585,N_9127,N_9295);
and UO_586 (O_586,N_9704,N_9586);
nor UO_587 (O_587,N_9983,N_9361);
nand UO_588 (O_588,N_9143,N_9184);
nand UO_589 (O_589,N_9571,N_9007);
nand UO_590 (O_590,N_9065,N_9920);
nor UO_591 (O_591,N_9532,N_9543);
nor UO_592 (O_592,N_9522,N_9888);
or UO_593 (O_593,N_9365,N_9632);
and UO_594 (O_594,N_9361,N_9090);
nor UO_595 (O_595,N_9805,N_9078);
nor UO_596 (O_596,N_9319,N_9895);
nand UO_597 (O_597,N_9606,N_9372);
or UO_598 (O_598,N_9923,N_9496);
nor UO_599 (O_599,N_9685,N_9912);
nor UO_600 (O_600,N_9977,N_9519);
nand UO_601 (O_601,N_9674,N_9143);
and UO_602 (O_602,N_9223,N_9157);
or UO_603 (O_603,N_9028,N_9001);
nand UO_604 (O_604,N_9405,N_9079);
and UO_605 (O_605,N_9807,N_9413);
and UO_606 (O_606,N_9975,N_9510);
or UO_607 (O_607,N_9466,N_9427);
nor UO_608 (O_608,N_9728,N_9917);
nand UO_609 (O_609,N_9462,N_9741);
and UO_610 (O_610,N_9529,N_9895);
and UO_611 (O_611,N_9515,N_9189);
and UO_612 (O_612,N_9983,N_9574);
and UO_613 (O_613,N_9830,N_9375);
nand UO_614 (O_614,N_9816,N_9434);
nand UO_615 (O_615,N_9689,N_9330);
or UO_616 (O_616,N_9650,N_9812);
or UO_617 (O_617,N_9553,N_9276);
and UO_618 (O_618,N_9410,N_9880);
and UO_619 (O_619,N_9524,N_9243);
and UO_620 (O_620,N_9500,N_9301);
and UO_621 (O_621,N_9301,N_9042);
and UO_622 (O_622,N_9323,N_9037);
nand UO_623 (O_623,N_9288,N_9277);
and UO_624 (O_624,N_9591,N_9193);
nand UO_625 (O_625,N_9997,N_9337);
or UO_626 (O_626,N_9305,N_9496);
or UO_627 (O_627,N_9874,N_9524);
nand UO_628 (O_628,N_9530,N_9811);
or UO_629 (O_629,N_9757,N_9862);
nand UO_630 (O_630,N_9240,N_9907);
nand UO_631 (O_631,N_9123,N_9730);
nor UO_632 (O_632,N_9308,N_9449);
nand UO_633 (O_633,N_9471,N_9564);
and UO_634 (O_634,N_9741,N_9652);
nand UO_635 (O_635,N_9604,N_9227);
or UO_636 (O_636,N_9211,N_9637);
nand UO_637 (O_637,N_9562,N_9377);
and UO_638 (O_638,N_9133,N_9257);
and UO_639 (O_639,N_9995,N_9005);
and UO_640 (O_640,N_9486,N_9802);
nor UO_641 (O_641,N_9788,N_9422);
nand UO_642 (O_642,N_9712,N_9218);
nor UO_643 (O_643,N_9214,N_9835);
nand UO_644 (O_644,N_9090,N_9367);
or UO_645 (O_645,N_9334,N_9272);
nand UO_646 (O_646,N_9061,N_9631);
and UO_647 (O_647,N_9383,N_9177);
and UO_648 (O_648,N_9174,N_9775);
nand UO_649 (O_649,N_9152,N_9980);
nand UO_650 (O_650,N_9258,N_9696);
or UO_651 (O_651,N_9153,N_9827);
and UO_652 (O_652,N_9106,N_9512);
and UO_653 (O_653,N_9047,N_9604);
or UO_654 (O_654,N_9775,N_9370);
nor UO_655 (O_655,N_9935,N_9817);
nand UO_656 (O_656,N_9956,N_9382);
nor UO_657 (O_657,N_9748,N_9889);
or UO_658 (O_658,N_9550,N_9447);
nand UO_659 (O_659,N_9967,N_9925);
and UO_660 (O_660,N_9859,N_9586);
nor UO_661 (O_661,N_9589,N_9228);
or UO_662 (O_662,N_9356,N_9140);
and UO_663 (O_663,N_9698,N_9353);
nor UO_664 (O_664,N_9366,N_9345);
nor UO_665 (O_665,N_9072,N_9546);
and UO_666 (O_666,N_9125,N_9932);
nand UO_667 (O_667,N_9828,N_9007);
or UO_668 (O_668,N_9272,N_9619);
nand UO_669 (O_669,N_9504,N_9287);
and UO_670 (O_670,N_9882,N_9574);
nor UO_671 (O_671,N_9486,N_9038);
nand UO_672 (O_672,N_9368,N_9598);
or UO_673 (O_673,N_9073,N_9055);
or UO_674 (O_674,N_9655,N_9427);
or UO_675 (O_675,N_9158,N_9070);
nor UO_676 (O_676,N_9832,N_9851);
and UO_677 (O_677,N_9946,N_9375);
nor UO_678 (O_678,N_9284,N_9712);
nor UO_679 (O_679,N_9677,N_9695);
xnor UO_680 (O_680,N_9826,N_9918);
and UO_681 (O_681,N_9599,N_9742);
or UO_682 (O_682,N_9143,N_9416);
nand UO_683 (O_683,N_9361,N_9866);
and UO_684 (O_684,N_9689,N_9149);
nand UO_685 (O_685,N_9997,N_9994);
or UO_686 (O_686,N_9524,N_9041);
or UO_687 (O_687,N_9110,N_9074);
nor UO_688 (O_688,N_9846,N_9243);
and UO_689 (O_689,N_9387,N_9732);
nor UO_690 (O_690,N_9113,N_9306);
nand UO_691 (O_691,N_9702,N_9228);
nor UO_692 (O_692,N_9317,N_9524);
and UO_693 (O_693,N_9884,N_9611);
xor UO_694 (O_694,N_9703,N_9606);
nor UO_695 (O_695,N_9316,N_9940);
nor UO_696 (O_696,N_9820,N_9243);
and UO_697 (O_697,N_9215,N_9331);
and UO_698 (O_698,N_9341,N_9335);
and UO_699 (O_699,N_9781,N_9992);
or UO_700 (O_700,N_9758,N_9893);
and UO_701 (O_701,N_9382,N_9365);
or UO_702 (O_702,N_9089,N_9557);
and UO_703 (O_703,N_9449,N_9568);
or UO_704 (O_704,N_9524,N_9996);
nor UO_705 (O_705,N_9861,N_9521);
nor UO_706 (O_706,N_9456,N_9757);
and UO_707 (O_707,N_9525,N_9072);
nand UO_708 (O_708,N_9377,N_9731);
and UO_709 (O_709,N_9539,N_9016);
nand UO_710 (O_710,N_9574,N_9872);
nand UO_711 (O_711,N_9991,N_9521);
nand UO_712 (O_712,N_9190,N_9011);
or UO_713 (O_713,N_9067,N_9853);
and UO_714 (O_714,N_9792,N_9014);
nor UO_715 (O_715,N_9423,N_9063);
nand UO_716 (O_716,N_9692,N_9749);
and UO_717 (O_717,N_9043,N_9989);
xor UO_718 (O_718,N_9615,N_9228);
or UO_719 (O_719,N_9873,N_9298);
and UO_720 (O_720,N_9765,N_9381);
nand UO_721 (O_721,N_9200,N_9293);
and UO_722 (O_722,N_9253,N_9486);
or UO_723 (O_723,N_9931,N_9213);
nor UO_724 (O_724,N_9474,N_9933);
or UO_725 (O_725,N_9990,N_9120);
nand UO_726 (O_726,N_9948,N_9298);
nand UO_727 (O_727,N_9598,N_9107);
and UO_728 (O_728,N_9840,N_9490);
nor UO_729 (O_729,N_9097,N_9858);
nand UO_730 (O_730,N_9018,N_9554);
or UO_731 (O_731,N_9519,N_9060);
nor UO_732 (O_732,N_9112,N_9979);
nor UO_733 (O_733,N_9007,N_9193);
or UO_734 (O_734,N_9731,N_9787);
nand UO_735 (O_735,N_9490,N_9836);
nor UO_736 (O_736,N_9079,N_9638);
nor UO_737 (O_737,N_9931,N_9654);
or UO_738 (O_738,N_9557,N_9541);
nand UO_739 (O_739,N_9216,N_9708);
nand UO_740 (O_740,N_9192,N_9438);
and UO_741 (O_741,N_9397,N_9897);
xnor UO_742 (O_742,N_9534,N_9887);
nor UO_743 (O_743,N_9661,N_9488);
and UO_744 (O_744,N_9721,N_9816);
and UO_745 (O_745,N_9333,N_9613);
nor UO_746 (O_746,N_9470,N_9872);
nand UO_747 (O_747,N_9689,N_9093);
nor UO_748 (O_748,N_9354,N_9765);
nand UO_749 (O_749,N_9892,N_9828);
or UO_750 (O_750,N_9451,N_9177);
and UO_751 (O_751,N_9939,N_9436);
nand UO_752 (O_752,N_9504,N_9634);
and UO_753 (O_753,N_9766,N_9367);
and UO_754 (O_754,N_9584,N_9464);
or UO_755 (O_755,N_9468,N_9237);
nand UO_756 (O_756,N_9197,N_9314);
and UO_757 (O_757,N_9044,N_9625);
nor UO_758 (O_758,N_9342,N_9957);
or UO_759 (O_759,N_9083,N_9534);
and UO_760 (O_760,N_9860,N_9461);
or UO_761 (O_761,N_9135,N_9631);
and UO_762 (O_762,N_9573,N_9956);
nor UO_763 (O_763,N_9229,N_9490);
nor UO_764 (O_764,N_9772,N_9530);
and UO_765 (O_765,N_9163,N_9699);
xnor UO_766 (O_766,N_9044,N_9048);
and UO_767 (O_767,N_9636,N_9586);
and UO_768 (O_768,N_9212,N_9051);
or UO_769 (O_769,N_9593,N_9545);
or UO_770 (O_770,N_9635,N_9435);
or UO_771 (O_771,N_9481,N_9559);
and UO_772 (O_772,N_9782,N_9615);
or UO_773 (O_773,N_9970,N_9618);
or UO_774 (O_774,N_9417,N_9481);
and UO_775 (O_775,N_9992,N_9785);
and UO_776 (O_776,N_9385,N_9157);
xor UO_777 (O_777,N_9269,N_9069);
or UO_778 (O_778,N_9468,N_9306);
nor UO_779 (O_779,N_9885,N_9333);
and UO_780 (O_780,N_9881,N_9821);
xnor UO_781 (O_781,N_9308,N_9009);
nand UO_782 (O_782,N_9994,N_9155);
nand UO_783 (O_783,N_9116,N_9477);
or UO_784 (O_784,N_9881,N_9273);
nor UO_785 (O_785,N_9411,N_9401);
and UO_786 (O_786,N_9762,N_9003);
nand UO_787 (O_787,N_9157,N_9098);
nor UO_788 (O_788,N_9256,N_9691);
xor UO_789 (O_789,N_9691,N_9212);
xor UO_790 (O_790,N_9326,N_9293);
nor UO_791 (O_791,N_9213,N_9405);
nand UO_792 (O_792,N_9824,N_9546);
nand UO_793 (O_793,N_9859,N_9736);
and UO_794 (O_794,N_9457,N_9526);
and UO_795 (O_795,N_9476,N_9037);
nor UO_796 (O_796,N_9174,N_9207);
and UO_797 (O_797,N_9221,N_9259);
or UO_798 (O_798,N_9789,N_9269);
and UO_799 (O_799,N_9597,N_9464);
and UO_800 (O_800,N_9955,N_9319);
nand UO_801 (O_801,N_9190,N_9256);
nor UO_802 (O_802,N_9556,N_9119);
and UO_803 (O_803,N_9015,N_9930);
nor UO_804 (O_804,N_9260,N_9761);
nor UO_805 (O_805,N_9560,N_9996);
nor UO_806 (O_806,N_9216,N_9566);
nand UO_807 (O_807,N_9244,N_9458);
nor UO_808 (O_808,N_9455,N_9513);
and UO_809 (O_809,N_9091,N_9073);
nor UO_810 (O_810,N_9860,N_9124);
nor UO_811 (O_811,N_9165,N_9497);
and UO_812 (O_812,N_9206,N_9471);
or UO_813 (O_813,N_9025,N_9186);
nor UO_814 (O_814,N_9451,N_9115);
nand UO_815 (O_815,N_9000,N_9935);
or UO_816 (O_816,N_9146,N_9324);
nor UO_817 (O_817,N_9913,N_9835);
or UO_818 (O_818,N_9595,N_9602);
nor UO_819 (O_819,N_9747,N_9403);
or UO_820 (O_820,N_9205,N_9586);
nand UO_821 (O_821,N_9736,N_9716);
and UO_822 (O_822,N_9845,N_9081);
nor UO_823 (O_823,N_9273,N_9251);
and UO_824 (O_824,N_9101,N_9728);
xnor UO_825 (O_825,N_9939,N_9005);
or UO_826 (O_826,N_9913,N_9121);
nand UO_827 (O_827,N_9772,N_9062);
nor UO_828 (O_828,N_9792,N_9708);
nand UO_829 (O_829,N_9765,N_9865);
nand UO_830 (O_830,N_9064,N_9161);
and UO_831 (O_831,N_9296,N_9247);
nand UO_832 (O_832,N_9599,N_9426);
or UO_833 (O_833,N_9331,N_9888);
and UO_834 (O_834,N_9781,N_9810);
and UO_835 (O_835,N_9731,N_9748);
nor UO_836 (O_836,N_9234,N_9740);
nand UO_837 (O_837,N_9885,N_9918);
nand UO_838 (O_838,N_9757,N_9290);
nand UO_839 (O_839,N_9699,N_9884);
nand UO_840 (O_840,N_9870,N_9489);
nor UO_841 (O_841,N_9522,N_9109);
and UO_842 (O_842,N_9336,N_9003);
and UO_843 (O_843,N_9361,N_9214);
nand UO_844 (O_844,N_9477,N_9445);
nand UO_845 (O_845,N_9934,N_9652);
nor UO_846 (O_846,N_9426,N_9840);
and UO_847 (O_847,N_9951,N_9537);
and UO_848 (O_848,N_9401,N_9836);
or UO_849 (O_849,N_9884,N_9646);
nor UO_850 (O_850,N_9306,N_9634);
xnor UO_851 (O_851,N_9641,N_9823);
or UO_852 (O_852,N_9493,N_9969);
nor UO_853 (O_853,N_9526,N_9868);
and UO_854 (O_854,N_9198,N_9613);
or UO_855 (O_855,N_9415,N_9381);
and UO_856 (O_856,N_9086,N_9175);
nand UO_857 (O_857,N_9717,N_9347);
or UO_858 (O_858,N_9539,N_9229);
nand UO_859 (O_859,N_9752,N_9786);
nor UO_860 (O_860,N_9455,N_9374);
or UO_861 (O_861,N_9945,N_9992);
nor UO_862 (O_862,N_9733,N_9866);
nor UO_863 (O_863,N_9146,N_9779);
nor UO_864 (O_864,N_9302,N_9260);
nor UO_865 (O_865,N_9756,N_9123);
nand UO_866 (O_866,N_9988,N_9283);
nor UO_867 (O_867,N_9645,N_9701);
or UO_868 (O_868,N_9448,N_9949);
nor UO_869 (O_869,N_9771,N_9430);
and UO_870 (O_870,N_9678,N_9788);
nor UO_871 (O_871,N_9017,N_9177);
nand UO_872 (O_872,N_9152,N_9538);
or UO_873 (O_873,N_9928,N_9026);
nor UO_874 (O_874,N_9622,N_9201);
nand UO_875 (O_875,N_9696,N_9378);
nor UO_876 (O_876,N_9776,N_9910);
nor UO_877 (O_877,N_9284,N_9135);
nor UO_878 (O_878,N_9678,N_9631);
or UO_879 (O_879,N_9000,N_9695);
or UO_880 (O_880,N_9593,N_9976);
and UO_881 (O_881,N_9523,N_9292);
nor UO_882 (O_882,N_9512,N_9617);
nor UO_883 (O_883,N_9631,N_9540);
or UO_884 (O_884,N_9136,N_9348);
and UO_885 (O_885,N_9666,N_9514);
nor UO_886 (O_886,N_9138,N_9984);
or UO_887 (O_887,N_9296,N_9022);
nor UO_888 (O_888,N_9907,N_9824);
or UO_889 (O_889,N_9454,N_9333);
or UO_890 (O_890,N_9229,N_9807);
nor UO_891 (O_891,N_9495,N_9782);
and UO_892 (O_892,N_9761,N_9824);
nand UO_893 (O_893,N_9819,N_9330);
and UO_894 (O_894,N_9719,N_9563);
and UO_895 (O_895,N_9685,N_9733);
nand UO_896 (O_896,N_9726,N_9283);
and UO_897 (O_897,N_9672,N_9919);
or UO_898 (O_898,N_9654,N_9156);
nor UO_899 (O_899,N_9622,N_9979);
nand UO_900 (O_900,N_9599,N_9471);
and UO_901 (O_901,N_9246,N_9337);
or UO_902 (O_902,N_9237,N_9343);
xnor UO_903 (O_903,N_9078,N_9560);
or UO_904 (O_904,N_9686,N_9645);
nor UO_905 (O_905,N_9901,N_9635);
nor UO_906 (O_906,N_9203,N_9463);
nor UO_907 (O_907,N_9822,N_9274);
nor UO_908 (O_908,N_9133,N_9040);
nand UO_909 (O_909,N_9226,N_9023);
or UO_910 (O_910,N_9825,N_9453);
nand UO_911 (O_911,N_9151,N_9023);
and UO_912 (O_912,N_9830,N_9755);
and UO_913 (O_913,N_9845,N_9339);
nor UO_914 (O_914,N_9951,N_9692);
nand UO_915 (O_915,N_9868,N_9896);
nor UO_916 (O_916,N_9142,N_9528);
nor UO_917 (O_917,N_9272,N_9482);
and UO_918 (O_918,N_9803,N_9053);
and UO_919 (O_919,N_9269,N_9517);
nand UO_920 (O_920,N_9000,N_9191);
and UO_921 (O_921,N_9126,N_9665);
or UO_922 (O_922,N_9996,N_9637);
nor UO_923 (O_923,N_9935,N_9008);
and UO_924 (O_924,N_9919,N_9428);
nand UO_925 (O_925,N_9814,N_9145);
or UO_926 (O_926,N_9555,N_9425);
nand UO_927 (O_927,N_9495,N_9719);
or UO_928 (O_928,N_9277,N_9674);
nand UO_929 (O_929,N_9463,N_9638);
nor UO_930 (O_930,N_9370,N_9467);
nor UO_931 (O_931,N_9448,N_9467);
or UO_932 (O_932,N_9192,N_9688);
or UO_933 (O_933,N_9912,N_9678);
nand UO_934 (O_934,N_9713,N_9650);
nor UO_935 (O_935,N_9211,N_9050);
nand UO_936 (O_936,N_9149,N_9321);
and UO_937 (O_937,N_9777,N_9511);
nor UO_938 (O_938,N_9196,N_9602);
and UO_939 (O_939,N_9011,N_9098);
or UO_940 (O_940,N_9137,N_9874);
nand UO_941 (O_941,N_9926,N_9295);
nand UO_942 (O_942,N_9844,N_9182);
or UO_943 (O_943,N_9937,N_9935);
xnor UO_944 (O_944,N_9256,N_9503);
nor UO_945 (O_945,N_9100,N_9039);
or UO_946 (O_946,N_9661,N_9118);
nor UO_947 (O_947,N_9942,N_9733);
and UO_948 (O_948,N_9810,N_9573);
xor UO_949 (O_949,N_9944,N_9631);
nand UO_950 (O_950,N_9638,N_9713);
nor UO_951 (O_951,N_9448,N_9559);
or UO_952 (O_952,N_9180,N_9146);
xor UO_953 (O_953,N_9594,N_9778);
nor UO_954 (O_954,N_9711,N_9114);
xnor UO_955 (O_955,N_9820,N_9045);
nand UO_956 (O_956,N_9731,N_9040);
nor UO_957 (O_957,N_9273,N_9575);
and UO_958 (O_958,N_9693,N_9252);
nor UO_959 (O_959,N_9529,N_9410);
or UO_960 (O_960,N_9927,N_9006);
and UO_961 (O_961,N_9905,N_9419);
nor UO_962 (O_962,N_9563,N_9630);
and UO_963 (O_963,N_9807,N_9606);
or UO_964 (O_964,N_9170,N_9766);
nand UO_965 (O_965,N_9638,N_9587);
and UO_966 (O_966,N_9137,N_9963);
or UO_967 (O_967,N_9238,N_9345);
and UO_968 (O_968,N_9395,N_9534);
or UO_969 (O_969,N_9075,N_9051);
and UO_970 (O_970,N_9791,N_9099);
or UO_971 (O_971,N_9290,N_9770);
nand UO_972 (O_972,N_9259,N_9774);
or UO_973 (O_973,N_9668,N_9168);
or UO_974 (O_974,N_9064,N_9079);
nand UO_975 (O_975,N_9575,N_9029);
and UO_976 (O_976,N_9396,N_9106);
and UO_977 (O_977,N_9568,N_9223);
or UO_978 (O_978,N_9412,N_9541);
nor UO_979 (O_979,N_9028,N_9275);
and UO_980 (O_980,N_9983,N_9713);
nand UO_981 (O_981,N_9473,N_9605);
nor UO_982 (O_982,N_9826,N_9556);
nand UO_983 (O_983,N_9246,N_9095);
and UO_984 (O_984,N_9434,N_9984);
nor UO_985 (O_985,N_9190,N_9161);
nor UO_986 (O_986,N_9492,N_9287);
nand UO_987 (O_987,N_9697,N_9405);
nor UO_988 (O_988,N_9833,N_9898);
or UO_989 (O_989,N_9697,N_9852);
nor UO_990 (O_990,N_9877,N_9991);
and UO_991 (O_991,N_9343,N_9294);
or UO_992 (O_992,N_9854,N_9882);
and UO_993 (O_993,N_9161,N_9367);
or UO_994 (O_994,N_9322,N_9263);
or UO_995 (O_995,N_9801,N_9308);
or UO_996 (O_996,N_9286,N_9532);
or UO_997 (O_997,N_9509,N_9749);
or UO_998 (O_998,N_9688,N_9212);
nand UO_999 (O_999,N_9404,N_9923);
nand UO_1000 (O_1000,N_9852,N_9468);
or UO_1001 (O_1001,N_9203,N_9392);
and UO_1002 (O_1002,N_9248,N_9955);
nand UO_1003 (O_1003,N_9123,N_9125);
nand UO_1004 (O_1004,N_9487,N_9207);
or UO_1005 (O_1005,N_9034,N_9649);
or UO_1006 (O_1006,N_9994,N_9719);
and UO_1007 (O_1007,N_9411,N_9017);
or UO_1008 (O_1008,N_9870,N_9021);
and UO_1009 (O_1009,N_9308,N_9180);
nor UO_1010 (O_1010,N_9360,N_9378);
nor UO_1011 (O_1011,N_9775,N_9077);
or UO_1012 (O_1012,N_9503,N_9537);
and UO_1013 (O_1013,N_9569,N_9640);
nor UO_1014 (O_1014,N_9600,N_9841);
nand UO_1015 (O_1015,N_9084,N_9563);
nand UO_1016 (O_1016,N_9375,N_9708);
nor UO_1017 (O_1017,N_9807,N_9944);
nand UO_1018 (O_1018,N_9984,N_9630);
or UO_1019 (O_1019,N_9829,N_9770);
xnor UO_1020 (O_1020,N_9056,N_9997);
and UO_1021 (O_1021,N_9399,N_9804);
and UO_1022 (O_1022,N_9262,N_9587);
nand UO_1023 (O_1023,N_9982,N_9030);
nor UO_1024 (O_1024,N_9272,N_9315);
nand UO_1025 (O_1025,N_9518,N_9047);
nand UO_1026 (O_1026,N_9112,N_9608);
or UO_1027 (O_1027,N_9085,N_9972);
nand UO_1028 (O_1028,N_9288,N_9172);
nand UO_1029 (O_1029,N_9972,N_9133);
nand UO_1030 (O_1030,N_9141,N_9781);
nand UO_1031 (O_1031,N_9852,N_9578);
nor UO_1032 (O_1032,N_9931,N_9522);
nor UO_1033 (O_1033,N_9057,N_9535);
and UO_1034 (O_1034,N_9580,N_9361);
nand UO_1035 (O_1035,N_9158,N_9208);
nor UO_1036 (O_1036,N_9309,N_9383);
and UO_1037 (O_1037,N_9912,N_9661);
xnor UO_1038 (O_1038,N_9105,N_9271);
and UO_1039 (O_1039,N_9408,N_9784);
nand UO_1040 (O_1040,N_9206,N_9325);
and UO_1041 (O_1041,N_9538,N_9036);
and UO_1042 (O_1042,N_9534,N_9864);
or UO_1043 (O_1043,N_9593,N_9389);
or UO_1044 (O_1044,N_9729,N_9028);
nand UO_1045 (O_1045,N_9583,N_9652);
nor UO_1046 (O_1046,N_9455,N_9720);
or UO_1047 (O_1047,N_9870,N_9027);
or UO_1048 (O_1048,N_9080,N_9087);
and UO_1049 (O_1049,N_9984,N_9074);
xor UO_1050 (O_1050,N_9588,N_9942);
and UO_1051 (O_1051,N_9684,N_9424);
nor UO_1052 (O_1052,N_9321,N_9057);
and UO_1053 (O_1053,N_9768,N_9433);
or UO_1054 (O_1054,N_9411,N_9630);
nor UO_1055 (O_1055,N_9675,N_9517);
or UO_1056 (O_1056,N_9763,N_9850);
nand UO_1057 (O_1057,N_9598,N_9618);
and UO_1058 (O_1058,N_9626,N_9232);
nand UO_1059 (O_1059,N_9226,N_9929);
nand UO_1060 (O_1060,N_9109,N_9436);
or UO_1061 (O_1061,N_9373,N_9925);
and UO_1062 (O_1062,N_9569,N_9867);
and UO_1063 (O_1063,N_9032,N_9740);
xor UO_1064 (O_1064,N_9717,N_9190);
and UO_1065 (O_1065,N_9222,N_9525);
and UO_1066 (O_1066,N_9949,N_9854);
nand UO_1067 (O_1067,N_9605,N_9674);
nor UO_1068 (O_1068,N_9128,N_9324);
nand UO_1069 (O_1069,N_9515,N_9269);
nor UO_1070 (O_1070,N_9995,N_9685);
nand UO_1071 (O_1071,N_9495,N_9763);
and UO_1072 (O_1072,N_9530,N_9821);
nand UO_1073 (O_1073,N_9399,N_9016);
nand UO_1074 (O_1074,N_9330,N_9564);
nor UO_1075 (O_1075,N_9915,N_9152);
nand UO_1076 (O_1076,N_9899,N_9667);
and UO_1077 (O_1077,N_9472,N_9476);
or UO_1078 (O_1078,N_9481,N_9828);
and UO_1079 (O_1079,N_9492,N_9935);
and UO_1080 (O_1080,N_9781,N_9140);
or UO_1081 (O_1081,N_9499,N_9121);
or UO_1082 (O_1082,N_9433,N_9064);
and UO_1083 (O_1083,N_9386,N_9001);
nand UO_1084 (O_1084,N_9876,N_9203);
and UO_1085 (O_1085,N_9205,N_9848);
nand UO_1086 (O_1086,N_9875,N_9135);
and UO_1087 (O_1087,N_9585,N_9080);
nor UO_1088 (O_1088,N_9636,N_9607);
and UO_1089 (O_1089,N_9054,N_9131);
or UO_1090 (O_1090,N_9419,N_9575);
or UO_1091 (O_1091,N_9130,N_9897);
or UO_1092 (O_1092,N_9682,N_9760);
nand UO_1093 (O_1093,N_9364,N_9094);
or UO_1094 (O_1094,N_9789,N_9192);
nand UO_1095 (O_1095,N_9655,N_9398);
nand UO_1096 (O_1096,N_9234,N_9261);
and UO_1097 (O_1097,N_9147,N_9680);
nor UO_1098 (O_1098,N_9805,N_9959);
nor UO_1099 (O_1099,N_9741,N_9276);
or UO_1100 (O_1100,N_9236,N_9288);
nand UO_1101 (O_1101,N_9491,N_9861);
nand UO_1102 (O_1102,N_9140,N_9999);
nand UO_1103 (O_1103,N_9078,N_9626);
and UO_1104 (O_1104,N_9438,N_9809);
nor UO_1105 (O_1105,N_9746,N_9102);
or UO_1106 (O_1106,N_9204,N_9822);
nand UO_1107 (O_1107,N_9920,N_9888);
and UO_1108 (O_1108,N_9257,N_9103);
nand UO_1109 (O_1109,N_9090,N_9644);
and UO_1110 (O_1110,N_9577,N_9461);
or UO_1111 (O_1111,N_9841,N_9363);
nand UO_1112 (O_1112,N_9611,N_9142);
nand UO_1113 (O_1113,N_9430,N_9949);
nor UO_1114 (O_1114,N_9457,N_9144);
and UO_1115 (O_1115,N_9361,N_9513);
or UO_1116 (O_1116,N_9318,N_9581);
and UO_1117 (O_1117,N_9074,N_9381);
or UO_1118 (O_1118,N_9666,N_9888);
and UO_1119 (O_1119,N_9013,N_9479);
or UO_1120 (O_1120,N_9135,N_9099);
or UO_1121 (O_1121,N_9450,N_9063);
or UO_1122 (O_1122,N_9828,N_9998);
nand UO_1123 (O_1123,N_9101,N_9048);
or UO_1124 (O_1124,N_9009,N_9956);
nand UO_1125 (O_1125,N_9620,N_9195);
or UO_1126 (O_1126,N_9093,N_9844);
nand UO_1127 (O_1127,N_9020,N_9087);
or UO_1128 (O_1128,N_9873,N_9131);
or UO_1129 (O_1129,N_9995,N_9135);
or UO_1130 (O_1130,N_9187,N_9953);
and UO_1131 (O_1131,N_9511,N_9725);
and UO_1132 (O_1132,N_9899,N_9837);
or UO_1133 (O_1133,N_9618,N_9222);
and UO_1134 (O_1134,N_9720,N_9841);
nor UO_1135 (O_1135,N_9867,N_9625);
xor UO_1136 (O_1136,N_9350,N_9333);
nand UO_1137 (O_1137,N_9741,N_9327);
nor UO_1138 (O_1138,N_9390,N_9863);
or UO_1139 (O_1139,N_9384,N_9314);
and UO_1140 (O_1140,N_9251,N_9168);
nor UO_1141 (O_1141,N_9223,N_9818);
or UO_1142 (O_1142,N_9042,N_9115);
and UO_1143 (O_1143,N_9023,N_9934);
and UO_1144 (O_1144,N_9006,N_9783);
nand UO_1145 (O_1145,N_9363,N_9276);
nor UO_1146 (O_1146,N_9935,N_9883);
nor UO_1147 (O_1147,N_9249,N_9624);
nand UO_1148 (O_1148,N_9334,N_9655);
nor UO_1149 (O_1149,N_9774,N_9700);
nor UO_1150 (O_1150,N_9386,N_9781);
and UO_1151 (O_1151,N_9382,N_9549);
and UO_1152 (O_1152,N_9173,N_9930);
xor UO_1153 (O_1153,N_9405,N_9185);
nor UO_1154 (O_1154,N_9802,N_9394);
nor UO_1155 (O_1155,N_9699,N_9651);
nand UO_1156 (O_1156,N_9626,N_9578);
nand UO_1157 (O_1157,N_9716,N_9411);
nor UO_1158 (O_1158,N_9207,N_9589);
or UO_1159 (O_1159,N_9207,N_9782);
or UO_1160 (O_1160,N_9340,N_9182);
nand UO_1161 (O_1161,N_9408,N_9491);
and UO_1162 (O_1162,N_9593,N_9365);
nand UO_1163 (O_1163,N_9551,N_9203);
nor UO_1164 (O_1164,N_9053,N_9200);
nand UO_1165 (O_1165,N_9958,N_9123);
and UO_1166 (O_1166,N_9939,N_9043);
nand UO_1167 (O_1167,N_9057,N_9350);
or UO_1168 (O_1168,N_9269,N_9590);
nor UO_1169 (O_1169,N_9300,N_9270);
nand UO_1170 (O_1170,N_9660,N_9848);
and UO_1171 (O_1171,N_9258,N_9202);
and UO_1172 (O_1172,N_9824,N_9517);
nand UO_1173 (O_1173,N_9506,N_9776);
and UO_1174 (O_1174,N_9290,N_9584);
and UO_1175 (O_1175,N_9688,N_9209);
nand UO_1176 (O_1176,N_9052,N_9855);
or UO_1177 (O_1177,N_9519,N_9459);
or UO_1178 (O_1178,N_9267,N_9370);
or UO_1179 (O_1179,N_9121,N_9016);
nand UO_1180 (O_1180,N_9091,N_9795);
and UO_1181 (O_1181,N_9669,N_9428);
or UO_1182 (O_1182,N_9084,N_9719);
or UO_1183 (O_1183,N_9858,N_9153);
and UO_1184 (O_1184,N_9565,N_9811);
or UO_1185 (O_1185,N_9747,N_9527);
or UO_1186 (O_1186,N_9607,N_9031);
and UO_1187 (O_1187,N_9105,N_9407);
nand UO_1188 (O_1188,N_9736,N_9516);
nor UO_1189 (O_1189,N_9526,N_9052);
nor UO_1190 (O_1190,N_9758,N_9015);
and UO_1191 (O_1191,N_9695,N_9390);
or UO_1192 (O_1192,N_9440,N_9340);
or UO_1193 (O_1193,N_9660,N_9369);
nand UO_1194 (O_1194,N_9867,N_9777);
nand UO_1195 (O_1195,N_9393,N_9181);
or UO_1196 (O_1196,N_9841,N_9905);
nor UO_1197 (O_1197,N_9821,N_9042);
nor UO_1198 (O_1198,N_9116,N_9743);
nand UO_1199 (O_1199,N_9855,N_9514);
nor UO_1200 (O_1200,N_9210,N_9941);
and UO_1201 (O_1201,N_9515,N_9251);
nand UO_1202 (O_1202,N_9967,N_9905);
or UO_1203 (O_1203,N_9575,N_9700);
nand UO_1204 (O_1204,N_9320,N_9491);
and UO_1205 (O_1205,N_9083,N_9616);
nor UO_1206 (O_1206,N_9976,N_9751);
nor UO_1207 (O_1207,N_9472,N_9178);
nor UO_1208 (O_1208,N_9013,N_9794);
nand UO_1209 (O_1209,N_9059,N_9006);
nor UO_1210 (O_1210,N_9427,N_9784);
nor UO_1211 (O_1211,N_9334,N_9942);
or UO_1212 (O_1212,N_9050,N_9379);
or UO_1213 (O_1213,N_9261,N_9347);
or UO_1214 (O_1214,N_9884,N_9920);
nand UO_1215 (O_1215,N_9193,N_9809);
or UO_1216 (O_1216,N_9040,N_9830);
and UO_1217 (O_1217,N_9361,N_9982);
or UO_1218 (O_1218,N_9848,N_9832);
or UO_1219 (O_1219,N_9920,N_9846);
nand UO_1220 (O_1220,N_9251,N_9025);
or UO_1221 (O_1221,N_9703,N_9458);
nor UO_1222 (O_1222,N_9137,N_9066);
nor UO_1223 (O_1223,N_9666,N_9581);
nor UO_1224 (O_1224,N_9830,N_9449);
and UO_1225 (O_1225,N_9236,N_9495);
or UO_1226 (O_1226,N_9385,N_9037);
and UO_1227 (O_1227,N_9400,N_9453);
and UO_1228 (O_1228,N_9998,N_9537);
and UO_1229 (O_1229,N_9287,N_9112);
nand UO_1230 (O_1230,N_9678,N_9179);
nand UO_1231 (O_1231,N_9487,N_9366);
and UO_1232 (O_1232,N_9774,N_9379);
nand UO_1233 (O_1233,N_9352,N_9853);
nand UO_1234 (O_1234,N_9726,N_9551);
and UO_1235 (O_1235,N_9626,N_9561);
or UO_1236 (O_1236,N_9690,N_9249);
or UO_1237 (O_1237,N_9505,N_9141);
or UO_1238 (O_1238,N_9710,N_9383);
and UO_1239 (O_1239,N_9929,N_9577);
nand UO_1240 (O_1240,N_9357,N_9151);
and UO_1241 (O_1241,N_9848,N_9281);
or UO_1242 (O_1242,N_9595,N_9523);
nor UO_1243 (O_1243,N_9255,N_9172);
and UO_1244 (O_1244,N_9580,N_9749);
xnor UO_1245 (O_1245,N_9493,N_9973);
nor UO_1246 (O_1246,N_9257,N_9811);
or UO_1247 (O_1247,N_9693,N_9144);
or UO_1248 (O_1248,N_9236,N_9883);
nand UO_1249 (O_1249,N_9969,N_9228);
nand UO_1250 (O_1250,N_9520,N_9602);
nor UO_1251 (O_1251,N_9288,N_9391);
or UO_1252 (O_1252,N_9916,N_9462);
and UO_1253 (O_1253,N_9989,N_9118);
nand UO_1254 (O_1254,N_9877,N_9460);
nand UO_1255 (O_1255,N_9159,N_9114);
nand UO_1256 (O_1256,N_9287,N_9376);
nand UO_1257 (O_1257,N_9635,N_9452);
nand UO_1258 (O_1258,N_9422,N_9035);
nor UO_1259 (O_1259,N_9281,N_9810);
nand UO_1260 (O_1260,N_9782,N_9494);
nand UO_1261 (O_1261,N_9039,N_9000);
and UO_1262 (O_1262,N_9979,N_9293);
and UO_1263 (O_1263,N_9878,N_9913);
or UO_1264 (O_1264,N_9582,N_9462);
or UO_1265 (O_1265,N_9843,N_9942);
or UO_1266 (O_1266,N_9685,N_9911);
or UO_1267 (O_1267,N_9438,N_9415);
nor UO_1268 (O_1268,N_9957,N_9728);
and UO_1269 (O_1269,N_9785,N_9641);
and UO_1270 (O_1270,N_9796,N_9846);
or UO_1271 (O_1271,N_9560,N_9694);
nand UO_1272 (O_1272,N_9940,N_9318);
nor UO_1273 (O_1273,N_9481,N_9521);
or UO_1274 (O_1274,N_9166,N_9517);
or UO_1275 (O_1275,N_9195,N_9091);
nand UO_1276 (O_1276,N_9669,N_9417);
or UO_1277 (O_1277,N_9995,N_9515);
and UO_1278 (O_1278,N_9951,N_9120);
and UO_1279 (O_1279,N_9265,N_9911);
and UO_1280 (O_1280,N_9266,N_9101);
nor UO_1281 (O_1281,N_9256,N_9411);
and UO_1282 (O_1282,N_9608,N_9008);
nor UO_1283 (O_1283,N_9669,N_9699);
nand UO_1284 (O_1284,N_9667,N_9558);
xnor UO_1285 (O_1285,N_9324,N_9638);
and UO_1286 (O_1286,N_9528,N_9968);
or UO_1287 (O_1287,N_9413,N_9354);
nand UO_1288 (O_1288,N_9859,N_9283);
and UO_1289 (O_1289,N_9153,N_9295);
nor UO_1290 (O_1290,N_9645,N_9339);
or UO_1291 (O_1291,N_9106,N_9645);
nand UO_1292 (O_1292,N_9513,N_9681);
nand UO_1293 (O_1293,N_9888,N_9186);
or UO_1294 (O_1294,N_9339,N_9989);
nand UO_1295 (O_1295,N_9920,N_9396);
or UO_1296 (O_1296,N_9983,N_9801);
nor UO_1297 (O_1297,N_9107,N_9559);
or UO_1298 (O_1298,N_9619,N_9875);
and UO_1299 (O_1299,N_9611,N_9570);
and UO_1300 (O_1300,N_9050,N_9834);
xnor UO_1301 (O_1301,N_9892,N_9453);
nand UO_1302 (O_1302,N_9147,N_9608);
nor UO_1303 (O_1303,N_9368,N_9595);
or UO_1304 (O_1304,N_9804,N_9970);
xnor UO_1305 (O_1305,N_9017,N_9247);
nor UO_1306 (O_1306,N_9045,N_9126);
nand UO_1307 (O_1307,N_9808,N_9296);
xnor UO_1308 (O_1308,N_9221,N_9700);
or UO_1309 (O_1309,N_9215,N_9738);
or UO_1310 (O_1310,N_9848,N_9680);
and UO_1311 (O_1311,N_9092,N_9592);
and UO_1312 (O_1312,N_9537,N_9638);
nor UO_1313 (O_1313,N_9455,N_9484);
nand UO_1314 (O_1314,N_9683,N_9181);
or UO_1315 (O_1315,N_9066,N_9642);
xor UO_1316 (O_1316,N_9542,N_9707);
nor UO_1317 (O_1317,N_9737,N_9233);
nand UO_1318 (O_1318,N_9266,N_9124);
nand UO_1319 (O_1319,N_9509,N_9143);
or UO_1320 (O_1320,N_9349,N_9165);
or UO_1321 (O_1321,N_9406,N_9142);
and UO_1322 (O_1322,N_9705,N_9153);
nand UO_1323 (O_1323,N_9072,N_9846);
nand UO_1324 (O_1324,N_9955,N_9680);
and UO_1325 (O_1325,N_9256,N_9345);
nor UO_1326 (O_1326,N_9459,N_9632);
nor UO_1327 (O_1327,N_9850,N_9677);
nand UO_1328 (O_1328,N_9339,N_9987);
nand UO_1329 (O_1329,N_9709,N_9033);
nand UO_1330 (O_1330,N_9895,N_9626);
nand UO_1331 (O_1331,N_9172,N_9352);
and UO_1332 (O_1332,N_9435,N_9972);
nor UO_1333 (O_1333,N_9747,N_9994);
or UO_1334 (O_1334,N_9654,N_9544);
nand UO_1335 (O_1335,N_9592,N_9850);
and UO_1336 (O_1336,N_9474,N_9964);
nor UO_1337 (O_1337,N_9813,N_9800);
and UO_1338 (O_1338,N_9981,N_9381);
and UO_1339 (O_1339,N_9139,N_9015);
nand UO_1340 (O_1340,N_9742,N_9094);
or UO_1341 (O_1341,N_9656,N_9484);
and UO_1342 (O_1342,N_9397,N_9876);
xnor UO_1343 (O_1343,N_9809,N_9424);
nand UO_1344 (O_1344,N_9063,N_9445);
and UO_1345 (O_1345,N_9689,N_9331);
nand UO_1346 (O_1346,N_9763,N_9237);
nand UO_1347 (O_1347,N_9631,N_9320);
or UO_1348 (O_1348,N_9487,N_9856);
nor UO_1349 (O_1349,N_9740,N_9551);
nor UO_1350 (O_1350,N_9483,N_9486);
and UO_1351 (O_1351,N_9033,N_9921);
or UO_1352 (O_1352,N_9863,N_9951);
and UO_1353 (O_1353,N_9826,N_9387);
and UO_1354 (O_1354,N_9889,N_9898);
nor UO_1355 (O_1355,N_9570,N_9726);
nor UO_1356 (O_1356,N_9041,N_9145);
or UO_1357 (O_1357,N_9169,N_9455);
or UO_1358 (O_1358,N_9433,N_9966);
and UO_1359 (O_1359,N_9137,N_9591);
nor UO_1360 (O_1360,N_9980,N_9854);
nand UO_1361 (O_1361,N_9534,N_9568);
or UO_1362 (O_1362,N_9427,N_9367);
nor UO_1363 (O_1363,N_9747,N_9478);
nor UO_1364 (O_1364,N_9509,N_9037);
and UO_1365 (O_1365,N_9564,N_9600);
xor UO_1366 (O_1366,N_9268,N_9500);
nor UO_1367 (O_1367,N_9080,N_9773);
and UO_1368 (O_1368,N_9090,N_9521);
nor UO_1369 (O_1369,N_9701,N_9042);
nand UO_1370 (O_1370,N_9932,N_9751);
nand UO_1371 (O_1371,N_9263,N_9422);
and UO_1372 (O_1372,N_9267,N_9990);
and UO_1373 (O_1373,N_9151,N_9597);
nand UO_1374 (O_1374,N_9917,N_9370);
and UO_1375 (O_1375,N_9281,N_9307);
nand UO_1376 (O_1376,N_9041,N_9341);
nand UO_1377 (O_1377,N_9641,N_9181);
nand UO_1378 (O_1378,N_9365,N_9500);
nor UO_1379 (O_1379,N_9434,N_9848);
nand UO_1380 (O_1380,N_9719,N_9369);
nand UO_1381 (O_1381,N_9220,N_9698);
and UO_1382 (O_1382,N_9153,N_9038);
nor UO_1383 (O_1383,N_9000,N_9276);
nor UO_1384 (O_1384,N_9957,N_9159);
nand UO_1385 (O_1385,N_9940,N_9234);
or UO_1386 (O_1386,N_9499,N_9457);
nand UO_1387 (O_1387,N_9368,N_9304);
nor UO_1388 (O_1388,N_9097,N_9320);
and UO_1389 (O_1389,N_9839,N_9539);
or UO_1390 (O_1390,N_9582,N_9645);
or UO_1391 (O_1391,N_9357,N_9329);
and UO_1392 (O_1392,N_9516,N_9680);
xor UO_1393 (O_1393,N_9613,N_9479);
and UO_1394 (O_1394,N_9861,N_9703);
nor UO_1395 (O_1395,N_9951,N_9272);
nor UO_1396 (O_1396,N_9899,N_9223);
nor UO_1397 (O_1397,N_9731,N_9366);
or UO_1398 (O_1398,N_9023,N_9606);
nor UO_1399 (O_1399,N_9741,N_9370);
nor UO_1400 (O_1400,N_9375,N_9967);
nor UO_1401 (O_1401,N_9574,N_9485);
nor UO_1402 (O_1402,N_9235,N_9036);
nand UO_1403 (O_1403,N_9844,N_9250);
nand UO_1404 (O_1404,N_9049,N_9511);
nor UO_1405 (O_1405,N_9148,N_9865);
nor UO_1406 (O_1406,N_9411,N_9768);
nor UO_1407 (O_1407,N_9154,N_9956);
and UO_1408 (O_1408,N_9402,N_9016);
and UO_1409 (O_1409,N_9015,N_9354);
and UO_1410 (O_1410,N_9065,N_9885);
nand UO_1411 (O_1411,N_9273,N_9192);
and UO_1412 (O_1412,N_9424,N_9384);
or UO_1413 (O_1413,N_9914,N_9915);
or UO_1414 (O_1414,N_9426,N_9052);
and UO_1415 (O_1415,N_9453,N_9597);
nand UO_1416 (O_1416,N_9872,N_9389);
nor UO_1417 (O_1417,N_9618,N_9367);
nand UO_1418 (O_1418,N_9852,N_9964);
nand UO_1419 (O_1419,N_9937,N_9563);
nor UO_1420 (O_1420,N_9130,N_9973);
nand UO_1421 (O_1421,N_9129,N_9078);
or UO_1422 (O_1422,N_9517,N_9551);
nor UO_1423 (O_1423,N_9015,N_9370);
nor UO_1424 (O_1424,N_9350,N_9232);
xor UO_1425 (O_1425,N_9043,N_9321);
or UO_1426 (O_1426,N_9949,N_9621);
nand UO_1427 (O_1427,N_9764,N_9268);
and UO_1428 (O_1428,N_9309,N_9187);
nand UO_1429 (O_1429,N_9907,N_9704);
and UO_1430 (O_1430,N_9490,N_9930);
and UO_1431 (O_1431,N_9532,N_9136);
xnor UO_1432 (O_1432,N_9461,N_9788);
and UO_1433 (O_1433,N_9833,N_9778);
or UO_1434 (O_1434,N_9389,N_9637);
and UO_1435 (O_1435,N_9237,N_9909);
and UO_1436 (O_1436,N_9772,N_9460);
and UO_1437 (O_1437,N_9045,N_9454);
and UO_1438 (O_1438,N_9570,N_9346);
and UO_1439 (O_1439,N_9082,N_9261);
nand UO_1440 (O_1440,N_9368,N_9453);
nor UO_1441 (O_1441,N_9904,N_9400);
nand UO_1442 (O_1442,N_9638,N_9397);
and UO_1443 (O_1443,N_9187,N_9274);
nand UO_1444 (O_1444,N_9376,N_9255);
nor UO_1445 (O_1445,N_9798,N_9645);
nand UO_1446 (O_1446,N_9695,N_9544);
or UO_1447 (O_1447,N_9927,N_9958);
or UO_1448 (O_1448,N_9872,N_9509);
nand UO_1449 (O_1449,N_9560,N_9538);
nand UO_1450 (O_1450,N_9462,N_9515);
nand UO_1451 (O_1451,N_9257,N_9163);
or UO_1452 (O_1452,N_9104,N_9605);
and UO_1453 (O_1453,N_9863,N_9897);
nor UO_1454 (O_1454,N_9969,N_9502);
nor UO_1455 (O_1455,N_9249,N_9762);
nand UO_1456 (O_1456,N_9367,N_9764);
and UO_1457 (O_1457,N_9417,N_9507);
nand UO_1458 (O_1458,N_9233,N_9757);
nor UO_1459 (O_1459,N_9775,N_9578);
nand UO_1460 (O_1460,N_9202,N_9068);
nor UO_1461 (O_1461,N_9523,N_9869);
and UO_1462 (O_1462,N_9578,N_9606);
xor UO_1463 (O_1463,N_9929,N_9337);
and UO_1464 (O_1464,N_9051,N_9834);
nand UO_1465 (O_1465,N_9468,N_9650);
or UO_1466 (O_1466,N_9236,N_9384);
nor UO_1467 (O_1467,N_9837,N_9942);
or UO_1468 (O_1468,N_9490,N_9137);
and UO_1469 (O_1469,N_9597,N_9026);
nor UO_1470 (O_1470,N_9253,N_9701);
and UO_1471 (O_1471,N_9896,N_9736);
nand UO_1472 (O_1472,N_9754,N_9876);
nor UO_1473 (O_1473,N_9532,N_9013);
nand UO_1474 (O_1474,N_9061,N_9522);
nor UO_1475 (O_1475,N_9787,N_9955);
nand UO_1476 (O_1476,N_9586,N_9895);
nor UO_1477 (O_1477,N_9211,N_9603);
and UO_1478 (O_1478,N_9064,N_9676);
and UO_1479 (O_1479,N_9497,N_9606);
xnor UO_1480 (O_1480,N_9579,N_9999);
nand UO_1481 (O_1481,N_9725,N_9962);
nand UO_1482 (O_1482,N_9070,N_9230);
or UO_1483 (O_1483,N_9254,N_9169);
nand UO_1484 (O_1484,N_9592,N_9579);
and UO_1485 (O_1485,N_9755,N_9612);
or UO_1486 (O_1486,N_9717,N_9072);
nand UO_1487 (O_1487,N_9378,N_9867);
nand UO_1488 (O_1488,N_9348,N_9945);
nor UO_1489 (O_1489,N_9249,N_9460);
nor UO_1490 (O_1490,N_9438,N_9351);
and UO_1491 (O_1491,N_9421,N_9634);
nor UO_1492 (O_1492,N_9585,N_9702);
nand UO_1493 (O_1493,N_9687,N_9329);
nand UO_1494 (O_1494,N_9748,N_9849);
nand UO_1495 (O_1495,N_9711,N_9210);
nor UO_1496 (O_1496,N_9430,N_9434);
nand UO_1497 (O_1497,N_9124,N_9450);
and UO_1498 (O_1498,N_9901,N_9506);
and UO_1499 (O_1499,N_9627,N_9546);
endmodule