module basic_500_3000_500_40_levels_2xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_236,In_402);
nand U1 (N_1,In_281,In_7);
nand U2 (N_2,In_432,In_112);
nand U3 (N_3,In_439,In_472);
or U4 (N_4,In_337,In_444);
and U5 (N_5,In_296,In_206);
nor U6 (N_6,In_125,In_97);
or U7 (N_7,In_393,In_204);
nand U8 (N_8,In_146,In_47);
and U9 (N_9,In_480,In_376);
nor U10 (N_10,In_63,In_134);
and U11 (N_11,In_258,In_95);
or U12 (N_12,In_40,In_308);
nand U13 (N_13,In_162,In_357);
nand U14 (N_14,In_88,In_365);
nand U15 (N_15,In_27,In_271);
and U16 (N_16,In_441,In_447);
and U17 (N_17,In_413,In_44);
or U18 (N_18,In_317,In_153);
nor U19 (N_19,In_187,In_228);
or U20 (N_20,In_494,In_222);
or U21 (N_21,In_461,In_75);
nand U22 (N_22,In_121,In_157);
nor U23 (N_23,In_349,In_0);
nor U24 (N_24,In_60,In_225);
nor U25 (N_25,In_417,In_195);
or U26 (N_26,In_249,In_465);
nor U27 (N_27,In_318,In_16);
nand U28 (N_28,In_129,In_245);
or U29 (N_29,In_17,In_102);
nand U30 (N_30,In_115,In_110);
nor U31 (N_31,In_107,In_471);
or U32 (N_32,In_20,In_213);
nor U33 (N_33,In_197,In_426);
nor U34 (N_34,In_468,In_34);
or U35 (N_35,In_404,In_360);
and U36 (N_36,In_248,In_114);
or U37 (N_37,In_184,In_333);
nor U38 (N_38,In_78,In_205);
nand U39 (N_39,In_10,In_268);
and U40 (N_40,In_384,In_92);
nand U41 (N_41,In_454,In_85);
nand U42 (N_42,In_239,In_288);
nand U43 (N_43,In_346,In_409);
nor U44 (N_44,In_351,In_411);
nand U45 (N_45,In_499,In_490);
nor U46 (N_46,In_183,In_263);
nand U47 (N_47,In_304,In_159);
nor U48 (N_48,In_152,In_434);
and U49 (N_49,In_270,In_166);
nor U50 (N_50,In_292,In_389);
nand U51 (N_51,In_366,In_113);
nand U52 (N_52,In_164,In_279);
or U53 (N_53,In_335,In_273);
and U54 (N_54,In_93,In_190);
and U55 (N_55,In_23,In_182);
nor U56 (N_56,In_329,In_32);
nor U57 (N_57,In_66,In_94);
nand U58 (N_58,In_74,In_52);
nor U59 (N_59,In_22,In_13);
and U60 (N_60,In_478,In_386);
or U61 (N_61,In_62,In_381);
and U62 (N_62,In_429,In_254);
or U63 (N_63,In_283,In_211);
nor U64 (N_64,In_12,In_436);
or U65 (N_65,In_262,In_364);
nor U66 (N_66,In_358,In_124);
or U67 (N_67,In_339,In_145);
or U68 (N_68,In_420,In_498);
or U69 (N_69,In_477,In_325);
nor U70 (N_70,In_445,In_57);
or U71 (N_71,In_255,In_280);
nor U72 (N_72,In_485,In_31);
or U73 (N_73,In_135,In_352);
nand U74 (N_74,In_370,In_488);
nor U75 (N_75,In_3,N_48);
xnor U76 (N_76,In_49,In_24);
nor U77 (N_77,In_141,In_421);
or U78 (N_78,N_29,In_104);
nor U79 (N_79,In_403,In_448);
and U80 (N_80,In_290,In_398);
or U81 (N_81,In_54,In_437);
nand U82 (N_82,In_315,In_122);
or U83 (N_83,N_59,In_450);
and U84 (N_84,N_30,In_231);
and U85 (N_85,N_46,In_43);
or U86 (N_86,In_19,In_176);
nor U87 (N_87,In_451,In_497);
nand U88 (N_88,In_342,In_482);
nand U89 (N_89,In_87,In_408);
or U90 (N_90,In_362,In_274);
nor U91 (N_91,In_460,In_181);
nand U92 (N_92,In_167,In_82);
and U93 (N_93,N_16,In_394);
and U94 (N_94,In_210,N_41);
and U95 (N_95,N_33,In_138);
nor U96 (N_96,In_15,In_470);
or U97 (N_97,In_56,In_269);
nand U98 (N_98,In_155,In_265);
nor U99 (N_99,In_350,In_128);
or U100 (N_100,In_380,In_440);
or U101 (N_101,N_15,In_185);
nand U102 (N_102,In_142,In_233);
nand U103 (N_103,In_143,N_51);
and U104 (N_104,In_61,In_243);
nand U105 (N_105,In_286,In_492);
nor U106 (N_106,In_226,In_382);
nand U107 (N_107,In_35,N_68);
and U108 (N_108,In_202,In_18);
nand U109 (N_109,In_84,In_449);
and U110 (N_110,In_310,In_193);
nand U111 (N_111,In_46,N_63);
nor U112 (N_112,In_400,In_45);
nor U113 (N_113,In_169,In_319);
nand U114 (N_114,In_117,In_201);
and U115 (N_115,In_285,In_36);
nand U116 (N_116,N_5,In_67);
or U117 (N_117,N_18,In_373);
nand U118 (N_118,N_17,In_305);
and U119 (N_119,In_89,In_455);
and U120 (N_120,N_6,In_474);
and U121 (N_121,In_363,In_453);
nand U122 (N_122,In_313,In_396);
and U123 (N_123,In_29,In_163);
or U124 (N_124,In_147,In_495);
xor U125 (N_125,In_8,In_230);
and U126 (N_126,In_234,In_422);
and U127 (N_127,In_433,In_221);
nor U128 (N_128,In_321,In_341);
or U129 (N_129,In_70,In_322);
and U130 (N_130,N_49,In_377);
nand U131 (N_131,N_26,In_241);
or U132 (N_132,In_303,In_173);
nor U133 (N_133,In_459,In_106);
nor U134 (N_134,In_469,In_212);
and U135 (N_135,N_67,N_7);
nand U136 (N_136,In_108,In_224);
or U137 (N_137,In_232,In_48);
and U138 (N_138,In_332,In_264);
nand U139 (N_139,In_372,In_30);
xnor U140 (N_140,In_257,In_475);
nand U141 (N_141,In_144,In_25);
and U142 (N_142,In_50,In_424);
and U143 (N_143,In_493,In_479);
or U144 (N_144,In_237,In_276);
nor U145 (N_145,In_253,In_150);
nand U146 (N_146,In_180,In_220);
nand U147 (N_147,N_44,In_189);
and U148 (N_148,In_385,In_473);
nand U149 (N_149,In_359,In_399);
or U150 (N_150,In_390,N_12);
nand U151 (N_151,In_291,N_20);
nand U152 (N_152,N_101,In_136);
and U153 (N_153,In_328,N_113);
and U154 (N_154,N_138,In_81);
or U155 (N_155,In_59,In_240);
or U156 (N_156,N_50,N_39);
nand U157 (N_157,In_26,N_121);
or U158 (N_158,N_24,In_37);
nor U159 (N_159,N_42,N_95);
nand U160 (N_160,N_132,N_4);
nand U161 (N_161,In_246,In_1);
and U162 (N_162,In_284,In_344);
nor U163 (N_163,In_149,N_57);
or U164 (N_164,N_100,N_10);
or U165 (N_165,N_82,In_484);
or U166 (N_166,In_306,N_27);
nand U167 (N_167,In_235,In_367);
and U168 (N_168,N_108,In_397);
or U169 (N_169,In_238,N_34);
or U170 (N_170,N_89,N_143);
and U171 (N_171,N_90,In_229);
nand U172 (N_172,In_481,N_13);
and U173 (N_173,N_102,In_98);
nand U174 (N_174,In_215,In_406);
nand U175 (N_175,In_130,In_309);
and U176 (N_176,N_96,In_353);
and U177 (N_177,N_62,N_71);
and U178 (N_178,N_21,In_42);
and U179 (N_179,In_68,In_307);
or U180 (N_180,In_218,In_83);
and U181 (N_181,In_378,In_4);
or U182 (N_182,In_6,N_111);
or U183 (N_183,In_250,N_125);
or U184 (N_184,N_22,In_428);
and U185 (N_185,N_87,In_331);
nor U186 (N_186,N_149,N_119);
or U187 (N_187,In_247,N_127);
or U188 (N_188,In_69,N_77);
or U189 (N_189,N_123,In_298);
nor U190 (N_190,In_435,In_77);
or U191 (N_191,In_133,In_132);
xnor U192 (N_192,N_86,In_371);
or U193 (N_193,In_21,In_316);
and U194 (N_194,In_178,N_136);
and U195 (N_195,In_415,In_355);
and U196 (N_196,In_334,N_19);
xnor U197 (N_197,In_175,In_369);
or U198 (N_198,N_84,N_25);
or U199 (N_199,N_115,In_356);
nand U200 (N_200,In_491,N_8);
or U201 (N_201,N_99,N_40);
nand U202 (N_202,In_295,In_137);
or U203 (N_203,In_423,In_338);
or U204 (N_204,In_158,N_116);
or U205 (N_205,N_61,In_261);
or U206 (N_206,In_196,In_266);
nand U207 (N_207,In_2,N_97);
nand U208 (N_208,N_112,In_139);
and U209 (N_209,N_75,In_214);
nor U210 (N_210,In_76,In_466);
and U211 (N_211,In_242,In_96);
nor U212 (N_212,N_43,N_147);
nor U213 (N_213,N_85,N_122);
nor U214 (N_214,N_2,In_414);
and U215 (N_215,In_343,N_94);
nor U216 (N_216,N_74,N_31);
or U217 (N_217,In_151,N_66);
and U218 (N_218,N_35,In_320);
or U219 (N_219,N_134,In_156);
nand U220 (N_220,In_347,In_442);
nor U221 (N_221,In_90,N_107);
or U222 (N_222,N_109,In_383);
or U223 (N_223,In_251,In_39);
and U224 (N_224,In_278,N_60);
and U225 (N_225,N_199,In_28);
or U226 (N_226,In_191,N_154);
nand U227 (N_227,N_177,In_119);
nand U228 (N_228,N_174,N_130);
and U229 (N_229,N_171,In_198);
and U230 (N_230,In_171,N_222);
nor U231 (N_231,In_219,N_78);
or U232 (N_232,N_203,In_314);
and U233 (N_233,N_129,N_223);
and U234 (N_234,In_330,In_170);
nor U235 (N_235,In_203,N_165);
nor U236 (N_236,In_487,In_186);
and U237 (N_237,In_11,N_164);
nor U238 (N_238,N_209,In_327);
and U239 (N_239,N_32,In_361);
or U240 (N_240,N_224,N_37);
or U241 (N_241,N_219,In_99);
nand U242 (N_242,In_324,In_174);
nor U243 (N_243,In_5,N_1);
or U244 (N_244,In_188,In_419);
or U245 (N_245,In_9,In_73);
and U246 (N_246,N_126,N_152);
and U247 (N_247,In_438,N_167);
and U248 (N_248,In_208,N_220);
nand U249 (N_249,N_56,N_215);
or U250 (N_250,N_105,In_462);
nand U251 (N_251,N_187,In_486);
nor U252 (N_252,In_489,N_173);
nor U253 (N_253,N_162,In_51);
or U254 (N_254,In_148,N_218);
nand U255 (N_255,In_443,In_412);
or U256 (N_256,N_64,N_169);
or U257 (N_257,In_80,N_180);
nand U258 (N_258,In_282,In_275);
nand U259 (N_259,N_212,N_178);
or U260 (N_260,In_407,In_53);
nor U261 (N_261,In_55,In_91);
or U262 (N_262,N_201,N_70);
or U263 (N_263,N_93,In_375);
or U264 (N_264,N_150,N_0);
or U265 (N_265,N_137,In_345);
nand U266 (N_266,N_36,N_146);
and U267 (N_267,N_208,In_312);
nor U268 (N_268,N_140,N_114);
or U269 (N_269,N_185,In_14);
nand U270 (N_270,In_118,N_76);
nand U271 (N_271,N_128,In_38);
nor U272 (N_272,In_294,In_354);
and U273 (N_273,N_157,In_109);
and U274 (N_274,In_348,N_52);
or U275 (N_275,N_91,In_177);
nor U276 (N_276,N_186,In_392);
nand U277 (N_277,N_205,N_179);
nand U278 (N_278,In_405,In_311);
nor U279 (N_279,N_182,N_88);
nor U280 (N_280,N_210,N_65);
and U281 (N_281,N_188,In_259);
or U282 (N_282,In_131,N_14);
or U283 (N_283,In_199,In_100);
and U284 (N_284,In_127,In_299);
or U285 (N_285,N_166,In_297);
nand U286 (N_286,N_217,N_211);
and U287 (N_287,N_221,N_9);
and U288 (N_288,N_124,In_368);
or U289 (N_289,N_189,N_117);
nand U290 (N_290,In_272,N_38);
or U291 (N_291,In_165,In_223);
and U292 (N_292,N_131,N_206);
nor U293 (N_293,N_197,In_410);
nand U294 (N_294,In_431,N_214);
or U295 (N_295,In_172,In_123);
and U296 (N_296,In_58,N_191);
and U297 (N_297,In_425,In_179);
nand U298 (N_298,In_287,N_183);
or U299 (N_299,In_452,In_302);
nand U300 (N_300,N_58,In_244);
nand U301 (N_301,N_273,In_105);
nor U302 (N_302,N_251,In_256);
nand U303 (N_303,N_278,N_159);
nor U304 (N_304,In_71,N_172);
or U305 (N_305,In_217,N_257);
or U306 (N_306,In_374,N_283);
and U307 (N_307,N_237,N_246);
nor U308 (N_308,In_41,N_106);
nor U309 (N_309,In_401,N_243);
and U310 (N_310,In_379,In_64);
and U311 (N_311,In_154,N_247);
or U312 (N_312,N_103,In_340);
or U313 (N_313,In_326,In_252);
and U314 (N_314,N_288,N_190);
nor U315 (N_315,N_153,In_457);
xnor U316 (N_316,N_272,In_289);
nor U317 (N_317,N_294,In_458);
nor U318 (N_318,N_47,In_140);
and U319 (N_319,In_79,N_244);
nor U320 (N_320,N_264,N_250);
nand U321 (N_321,N_192,In_209);
nand U322 (N_322,N_282,N_110);
nor U323 (N_323,N_281,In_456);
or U324 (N_324,N_181,N_231);
nand U325 (N_325,In_194,In_200);
or U326 (N_326,N_69,N_226);
nand U327 (N_327,N_53,N_3);
or U328 (N_328,N_163,N_239);
and U329 (N_329,N_298,N_170);
and U330 (N_330,N_228,N_259);
and U331 (N_331,N_213,In_260);
nand U332 (N_332,In_336,N_253);
nand U333 (N_333,N_263,N_240);
nand U334 (N_334,N_284,In_207);
and U335 (N_335,N_254,N_289);
nor U336 (N_336,In_168,N_45);
nand U337 (N_337,In_33,N_160);
or U338 (N_338,In_86,In_388);
nand U339 (N_339,N_11,In_120);
nor U340 (N_340,N_242,In_464);
or U341 (N_341,N_194,N_156);
or U342 (N_342,In_395,N_295);
and U343 (N_343,N_23,N_293);
and U344 (N_344,N_248,In_277);
nand U345 (N_345,N_290,N_269);
or U346 (N_346,N_80,N_265);
and U347 (N_347,N_241,N_286);
nand U348 (N_348,N_275,In_116);
and U349 (N_349,N_271,In_416);
or U350 (N_350,In_300,N_216);
nand U351 (N_351,N_285,In_103);
or U352 (N_352,N_292,N_236);
nor U353 (N_353,N_232,N_133);
nand U354 (N_354,N_291,N_144);
nand U355 (N_355,N_249,N_135);
and U356 (N_356,In_267,N_276);
and U357 (N_357,N_72,N_176);
nor U358 (N_358,In_227,N_277);
nor U359 (N_359,In_323,N_195);
nor U360 (N_360,N_256,In_111);
nor U361 (N_361,N_193,In_446);
nand U362 (N_362,N_202,N_297);
and U363 (N_363,In_467,In_216);
nand U364 (N_364,N_270,N_238);
and U365 (N_365,N_235,N_118);
nand U366 (N_366,In_418,In_65);
or U367 (N_367,N_79,N_28);
and U368 (N_368,In_293,N_258);
nor U369 (N_369,N_279,N_161);
or U370 (N_370,N_155,In_161);
nor U371 (N_371,N_287,N_196);
or U372 (N_372,In_391,N_296);
nor U373 (N_373,In_496,N_198);
and U374 (N_374,In_430,N_145);
nand U375 (N_375,N_148,N_92);
or U376 (N_376,N_54,N_204);
or U377 (N_377,N_313,N_280);
nand U378 (N_378,N_83,N_261);
nand U379 (N_379,N_299,N_369);
and U380 (N_380,N_300,N_274);
or U381 (N_381,N_349,N_342);
or U382 (N_382,N_353,N_345);
and U383 (N_383,N_371,N_104);
or U384 (N_384,N_306,N_81);
nor U385 (N_385,In_126,N_341);
or U386 (N_386,In_160,N_304);
and U387 (N_387,N_338,N_55);
nor U388 (N_388,N_139,N_302);
or U389 (N_389,N_233,N_348);
or U390 (N_390,N_312,N_309);
nor U391 (N_391,N_303,N_255);
and U392 (N_392,N_307,In_483);
nor U393 (N_393,N_252,N_364);
nand U394 (N_394,N_360,N_230);
or U395 (N_395,N_336,N_354);
or U396 (N_396,N_310,N_200);
or U397 (N_397,N_324,N_318);
xnor U398 (N_398,N_356,N_339);
and U399 (N_399,N_344,N_325);
or U400 (N_400,N_322,N_120);
nand U401 (N_401,N_373,N_229);
and U402 (N_402,In_301,N_268);
and U403 (N_403,N_374,N_366);
or U404 (N_404,N_73,N_335);
nand U405 (N_405,N_321,N_346);
nand U406 (N_406,N_207,N_350);
or U407 (N_407,N_370,N_361);
nor U408 (N_408,N_184,N_332);
and U409 (N_409,N_319,N_355);
and U410 (N_410,In_72,N_267);
nor U411 (N_411,N_225,N_359);
nor U412 (N_412,N_333,N_352);
nand U413 (N_413,N_351,N_317);
or U414 (N_414,N_368,N_175);
and U415 (N_415,N_260,N_151);
xnor U416 (N_416,N_308,N_329);
nor U417 (N_417,N_357,N_347);
or U418 (N_418,In_192,N_358);
nand U419 (N_419,N_141,N_234);
or U420 (N_420,N_315,N_331);
nor U421 (N_421,N_372,N_98);
nor U422 (N_422,N_328,In_427);
nand U423 (N_423,N_158,N_316);
or U424 (N_424,N_367,N_262);
or U425 (N_425,N_326,N_343);
and U426 (N_426,N_320,N_227);
nand U427 (N_427,N_142,In_463);
nor U428 (N_428,N_363,N_311);
or U429 (N_429,N_340,N_266);
nand U430 (N_430,In_476,In_101);
or U431 (N_431,N_168,N_337);
nand U432 (N_432,N_245,N_314);
and U433 (N_433,N_327,N_334);
or U434 (N_434,N_330,N_365);
or U435 (N_435,In_387,N_362);
and U436 (N_436,N_301,N_305);
and U437 (N_437,N_323,N_168);
nor U438 (N_438,N_266,N_333);
or U439 (N_439,N_120,In_160);
and U440 (N_440,N_54,N_252);
or U441 (N_441,N_252,N_354);
nand U442 (N_442,N_268,N_339);
nor U443 (N_443,N_200,N_354);
nand U444 (N_444,N_362,N_333);
nand U445 (N_445,N_299,N_262);
and U446 (N_446,N_274,N_318);
and U447 (N_447,N_299,N_331);
and U448 (N_448,In_72,N_365);
nand U449 (N_449,N_142,N_314);
or U450 (N_450,N_382,N_442);
and U451 (N_451,N_400,N_404);
nand U452 (N_452,N_383,N_424);
nand U453 (N_453,N_402,N_419);
and U454 (N_454,N_433,N_435);
nor U455 (N_455,N_445,N_378);
and U456 (N_456,N_390,N_449);
nor U457 (N_457,N_375,N_394);
nor U458 (N_458,N_410,N_408);
or U459 (N_459,N_417,N_411);
and U460 (N_460,N_413,N_444);
and U461 (N_461,N_396,N_414);
or U462 (N_462,N_381,N_427);
or U463 (N_463,N_376,N_407);
nor U464 (N_464,N_380,N_392);
or U465 (N_465,N_398,N_399);
and U466 (N_466,N_391,N_416);
and U467 (N_467,N_393,N_423);
xnor U468 (N_468,N_425,N_415);
nor U469 (N_469,N_447,N_428);
nand U470 (N_470,N_420,N_441);
or U471 (N_471,N_439,N_388);
nand U472 (N_472,N_426,N_379);
nand U473 (N_473,N_384,N_448);
nand U474 (N_474,N_432,N_409);
or U475 (N_475,N_436,N_387);
xor U476 (N_476,N_434,N_430);
nor U477 (N_477,N_437,N_446);
and U478 (N_478,N_395,N_406);
or U479 (N_479,N_431,N_421);
and U480 (N_480,N_412,N_440);
nor U481 (N_481,N_443,N_438);
or U482 (N_482,N_422,N_389);
and U483 (N_483,N_405,N_397);
and U484 (N_484,N_385,N_386);
nor U485 (N_485,N_418,N_401);
and U486 (N_486,N_377,N_429);
and U487 (N_487,N_403,N_383);
or U488 (N_488,N_419,N_435);
or U489 (N_489,N_424,N_407);
and U490 (N_490,N_392,N_385);
xor U491 (N_491,N_447,N_375);
and U492 (N_492,N_426,N_435);
or U493 (N_493,N_443,N_383);
or U494 (N_494,N_393,N_427);
and U495 (N_495,N_399,N_384);
nand U496 (N_496,N_401,N_383);
nor U497 (N_497,N_385,N_449);
xnor U498 (N_498,N_378,N_447);
nand U499 (N_499,N_399,N_395);
and U500 (N_500,N_395,N_438);
nor U501 (N_501,N_401,N_429);
nor U502 (N_502,N_408,N_403);
and U503 (N_503,N_441,N_401);
nand U504 (N_504,N_377,N_437);
nand U505 (N_505,N_393,N_413);
nand U506 (N_506,N_417,N_405);
or U507 (N_507,N_431,N_379);
nor U508 (N_508,N_383,N_427);
nor U509 (N_509,N_387,N_400);
nor U510 (N_510,N_429,N_427);
and U511 (N_511,N_415,N_416);
and U512 (N_512,N_400,N_418);
nand U513 (N_513,N_443,N_378);
nor U514 (N_514,N_429,N_380);
nand U515 (N_515,N_411,N_402);
nand U516 (N_516,N_418,N_416);
and U517 (N_517,N_383,N_444);
and U518 (N_518,N_415,N_418);
or U519 (N_519,N_420,N_390);
or U520 (N_520,N_440,N_436);
xor U521 (N_521,N_448,N_415);
and U522 (N_522,N_407,N_440);
nor U523 (N_523,N_448,N_376);
and U524 (N_524,N_416,N_446);
or U525 (N_525,N_472,N_506);
nor U526 (N_526,N_518,N_524);
or U527 (N_527,N_520,N_467);
nand U528 (N_528,N_499,N_502);
and U529 (N_529,N_458,N_523);
nor U530 (N_530,N_509,N_461);
and U531 (N_531,N_513,N_479);
or U532 (N_532,N_460,N_488);
nand U533 (N_533,N_473,N_489);
nor U534 (N_534,N_452,N_454);
nor U535 (N_535,N_503,N_517);
nand U536 (N_536,N_490,N_486);
or U537 (N_537,N_451,N_464);
nor U538 (N_538,N_521,N_470);
nand U539 (N_539,N_507,N_515);
and U540 (N_540,N_456,N_455);
and U541 (N_541,N_481,N_505);
nand U542 (N_542,N_450,N_497);
or U543 (N_543,N_477,N_469);
nand U544 (N_544,N_463,N_457);
and U545 (N_545,N_483,N_514);
nor U546 (N_546,N_508,N_504);
nand U547 (N_547,N_485,N_495);
nor U548 (N_548,N_476,N_475);
or U549 (N_549,N_462,N_491);
and U550 (N_550,N_496,N_494);
and U551 (N_551,N_482,N_487);
and U552 (N_552,N_471,N_522);
and U553 (N_553,N_501,N_511);
nor U554 (N_554,N_459,N_510);
or U555 (N_555,N_493,N_492);
or U556 (N_556,N_466,N_500);
and U557 (N_557,N_468,N_480);
and U558 (N_558,N_512,N_478);
nor U559 (N_559,N_474,N_484);
nor U560 (N_560,N_453,N_516);
nor U561 (N_561,N_465,N_498);
and U562 (N_562,N_519,N_520);
or U563 (N_563,N_465,N_485);
nor U564 (N_564,N_515,N_496);
nor U565 (N_565,N_489,N_466);
and U566 (N_566,N_499,N_453);
nand U567 (N_567,N_477,N_486);
nor U568 (N_568,N_451,N_472);
nand U569 (N_569,N_484,N_499);
nand U570 (N_570,N_516,N_463);
or U571 (N_571,N_464,N_463);
nor U572 (N_572,N_463,N_487);
nor U573 (N_573,N_451,N_476);
or U574 (N_574,N_497,N_512);
nand U575 (N_575,N_481,N_460);
nand U576 (N_576,N_468,N_515);
and U577 (N_577,N_464,N_458);
and U578 (N_578,N_501,N_484);
and U579 (N_579,N_469,N_493);
or U580 (N_580,N_464,N_489);
and U581 (N_581,N_486,N_499);
or U582 (N_582,N_475,N_522);
nor U583 (N_583,N_505,N_509);
nor U584 (N_584,N_454,N_480);
nand U585 (N_585,N_520,N_493);
nor U586 (N_586,N_462,N_458);
or U587 (N_587,N_495,N_513);
and U588 (N_588,N_480,N_517);
xor U589 (N_589,N_503,N_482);
or U590 (N_590,N_494,N_475);
nor U591 (N_591,N_506,N_456);
and U592 (N_592,N_515,N_522);
or U593 (N_593,N_489,N_509);
nand U594 (N_594,N_481,N_502);
nor U595 (N_595,N_492,N_503);
nand U596 (N_596,N_513,N_507);
nor U597 (N_597,N_462,N_494);
nor U598 (N_598,N_476,N_466);
or U599 (N_599,N_504,N_486);
and U600 (N_600,N_536,N_530);
nor U601 (N_601,N_566,N_570);
nor U602 (N_602,N_575,N_564);
nand U603 (N_603,N_574,N_589);
nand U604 (N_604,N_550,N_549);
nand U605 (N_605,N_599,N_563);
nor U606 (N_606,N_572,N_558);
xnor U607 (N_607,N_571,N_576);
nand U608 (N_608,N_593,N_587);
or U609 (N_609,N_534,N_596);
and U610 (N_610,N_545,N_557);
and U611 (N_611,N_547,N_527);
or U612 (N_612,N_561,N_567);
nor U613 (N_613,N_541,N_538);
and U614 (N_614,N_569,N_594);
and U615 (N_615,N_585,N_588);
nor U616 (N_616,N_540,N_542);
nor U617 (N_617,N_552,N_560);
or U618 (N_618,N_543,N_531);
nand U619 (N_619,N_586,N_548);
nor U620 (N_620,N_581,N_535);
and U621 (N_621,N_562,N_590);
or U622 (N_622,N_528,N_592);
or U623 (N_623,N_553,N_577);
and U624 (N_624,N_573,N_597);
or U625 (N_625,N_546,N_565);
nor U626 (N_626,N_578,N_555);
nand U627 (N_627,N_556,N_539);
and U628 (N_628,N_584,N_526);
or U629 (N_629,N_580,N_537);
nor U630 (N_630,N_568,N_532);
and U631 (N_631,N_544,N_554);
xor U632 (N_632,N_533,N_529);
and U633 (N_633,N_583,N_559);
nor U634 (N_634,N_579,N_591);
nand U635 (N_635,N_595,N_525);
nor U636 (N_636,N_551,N_598);
and U637 (N_637,N_582,N_591);
nand U638 (N_638,N_542,N_567);
nor U639 (N_639,N_527,N_535);
or U640 (N_640,N_577,N_546);
nor U641 (N_641,N_568,N_581);
and U642 (N_642,N_555,N_572);
nor U643 (N_643,N_535,N_541);
nor U644 (N_644,N_599,N_554);
nor U645 (N_645,N_583,N_560);
nor U646 (N_646,N_558,N_582);
nor U647 (N_647,N_537,N_529);
nor U648 (N_648,N_539,N_534);
or U649 (N_649,N_596,N_544);
and U650 (N_650,N_564,N_568);
and U651 (N_651,N_536,N_577);
or U652 (N_652,N_561,N_532);
nor U653 (N_653,N_582,N_526);
nor U654 (N_654,N_599,N_561);
and U655 (N_655,N_526,N_532);
or U656 (N_656,N_581,N_584);
nor U657 (N_657,N_577,N_598);
or U658 (N_658,N_564,N_537);
or U659 (N_659,N_528,N_578);
and U660 (N_660,N_567,N_571);
or U661 (N_661,N_585,N_552);
and U662 (N_662,N_562,N_527);
nand U663 (N_663,N_569,N_541);
nand U664 (N_664,N_544,N_599);
or U665 (N_665,N_584,N_588);
nand U666 (N_666,N_597,N_592);
or U667 (N_667,N_551,N_529);
nand U668 (N_668,N_582,N_559);
and U669 (N_669,N_594,N_576);
or U670 (N_670,N_569,N_562);
or U671 (N_671,N_592,N_569);
nor U672 (N_672,N_594,N_547);
and U673 (N_673,N_574,N_554);
or U674 (N_674,N_556,N_596);
and U675 (N_675,N_645,N_672);
nor U676 (N_676,N_644,N_605);
or U677 (N_677,N_628,N_611);
nor U678 (N_678,N_602,N_646);
nand U679 (N_679,N_653,N_608);
nor U680 (N_680,N_649,N_606);
or U681 (N_681,N_638,N_663);
and U682 (N_682,N_661,N_667);
nand U683 (N_683,N_627,N_636);
nand U684 (N_684,N_673,N_601);
xnor U685 (N_685,N_671,N_634);
nand U686 (N_686,N_631,N_619);
nor U687 (N_687,N_633,N_656);
nor U688 (N_688,N_629,N_652);
nand U689 (N_689,N_648,N_642);
or U690 (N_690,N_660,N_639);
nor U691 (N_691,N_641,N_659);
nor U692 (N_692,N_612,N_658);
nor U693 (N_693,N_637,N_600);
nor U694 (N_694,N_668,N_674);
nor U695 (N_695,N_643,N_607);
and U696 (N_696,N_650,N_662);
and U697 (N_697,N_620,N_621);
nand U698 (N_698,N_610,N_622);
xor U699 (N_699,N_615,N_630);
or U700 (N_700,N_609,N_617);
or U701 (N_701,N_635,N_625);
nor U702 (N_702,N_604,N_654);
or U703 (N_703,N_651,N_670);
nand U704 (N_704,N_666,N_623);
nor U705 (N_705,N_640,N_613);
nor U706 (N_706,N_603,N_655);
nand U707 (N_707,N_632,N_624);
or U708 (N_708,N_626,N_657);
and U709 (N_709,N_614,N_618);
or U710 (N_710,N_664,N_616);
or U711 (N_711,N_669,N_647);
nand U712 (N_712,N_665,N_634);
or U713 (N_713,N_610,N_643);
nand U714 (N_714,N_649,N_612);
or U715 (N_715,N_628,N_670);
or U716 (N_716,N_606,N_648);
and U717 (N_717,N_641,N_615);
nand U718 (N_718,N_674,N_671);
or U719 (N_719,N_610,N_667);
xor U720 (N_720,N_614,N_674);
nor U721 (N_721,N_604,N_659);
or U722 (N_722,N_625,N_605);
nor U723 (N_723,N_642,N_619);
or U724 (N_724,N_663,N_614);
nand U725 (N_725,N_659,N_654);
nor U726 (N_726,N_640,N_630);
and U727 (N_727,N_634,N_636);
nand U728 (N_728,N_622,N_617);
nand U729 (N_729,N_623,N_600);
and U730 (N_730,N_655,N_601);
nor U731 (N_731,N_669,N_670);
or U732 (N_732,N_650,N_619);
nand U733 (N_733,N_624,N_644);
nand U734 (N_734,N_646,N_611);
xor U735 (N_735,N_646,N_668);
or U736 (N_736,N_636,N_602);
nand U737 (N_737,N_629,N_661);
nand U738 (N_738,N_646,N_653);
or U739 (N_739,N_631,N_636);
and U740 (N_740,N_659,N_610);
or U741 (N_741,N_667,N_653);
nand U742 (N_742,N_635,N_673);
nor U743 (N_743,N_625,N_629);
and U744 (N_744,N_668,N_613);
or U745 (N_745,N_630,N_603);
and U746 (N_746,N_635,N_668);
or U747 (N_747,N_632,N_612);
or U748 (N_748,N_674,N_636);
nor U749 (N_749,N_629,N_674);
nand U750 (N_750,N_692,N_683);
or U751 (N_751,N_679,N_713);
and U752 (N_752,N_704,N_747);
and U753 (N_753,N_744,N_748);
and U754 (N_754,N_728,N_711);
or U755 (N_755,N_705,N_732);
or U756 (N_756,N_706,N_709);
nand U757 (N_757,N_703,N_690);
xnor U758 (N_758,N_720,N_694);
nand U759 (N_759,N_714,N_727);
nand U760 (N_760,N_701,N_726);
nor U761 (N_761,N_700,N_696);
and U762 (N_762,N_723,N_695);
nand U763 (N_763,N_729,N_689);
nor U764 (N_764,N_739,N_678);
nand U765 (N_765,N_735,N_715);
nand U766 (N_766,N_740,N_697);
and U767 (N_767,N_737,N_738);
or U768 (N_768,N_693,N_725);
nand U769 (N_769,N_686,N_681);
nor U770 (N_770,N_724,N_699);
nand U771 (N_771,N_736,N_710);
or U772 (N_772,N_688,N_718);
nor U773 (N_773,N_745,N_676);
nand U774 (N_774,N_708,N_702);
or U775 (N_775,N_698,N_675);
nor U776 (N_776,N_743,N_717);
nand U777 (N_777,N_733,N_742);
nand U778 (N_778,N_734,N_677);
nand U779 (N_779,N_707,N_716);
nand U780 (N_780,N_721,N_680);
nand U781 (N_781,N_685,N_746);
nor U782 (N_782,N_731,N_741);
nor U783 (N_783,N_682,N_749);
nor U784 (N_784,N_687,N_730);
nor U785 (N_785,N_722,N_719);
nor U786 (N_786,N_684,N_712);
or U787 (N_787,N_691,N_700);
nor U788 (N_788,N_697,N_748);
or U789 (N_789,N_675,N_730);
and U790 (N_790,N_684,N_747);
and U791 (N_791,N_684,N_724);
and U792 (N_792,N_679,N_719);
nor U793 (N_793,N_737,N_747);
or U794 (N_794,N_708,N_744);
nand U795 (N_795,N_749,N_748);
or U796 (N_796,N_741,N_689);
nor U797 (N_797,N_702,N_736);
nand U798 (N_798,N_710,N_678);
and U799 (N_799,N_676,N_721);
nor U800 (N_800,N_688,N_697);
nand U801 (N_801,N_690,N_679);
nand U802 (N_802,N_735,N_709);
or U803 (N_803,N_715,N_714);
and U804 (N_804,N_749,N_708);
nor U805 (N_805,N_727,N_716);
or U806 (N_806,N_731,N_748);
or U807 (N_807,N_714,N_737);
nor U808 (N_808,N_724,N_682);
or U809 (N_809,N_676,N_736);
nor U810 (N_810,N_734,N_737);
or U811 (N_811,N_688,N_701);
or U812 (N_812,N_725,N_717);
nor U813 (N_813,N_690,N_675);
nor U814 (N_814,N_676,N_681);
nand U815 (N_815,N_700,N_684);
nor U816 (N_816,N_687,N_690);
and U817 (N_817,N_684,N_687);
nand U818 (N_818,N_714,N_698);
or U819 (N_819,N_744,N_747);
nand U820 (N_820,N_693,N_696);
nand U821 (N_821,N_731,N_723);
nor U822 (N_822,N_688,N_691);
xnor U823 (N_823,N_681,N_718);
and U824 (N_824,N_705,N_678);
nand U825 (N_825,N_771,N_776);
or U826 (N_826,N_790,N_808);
and U827 (N_827,N_789,N_802);
and U828 (N_828,N_805,N_756);
nand U829 (N_829,N_755,N_784);
nand U830 (N_830,N_820,N_786);
or U831 (N_831,N_796,N_770);
nor U832 (N_832,N_797,N_806);
or U833 (N_833,N_754,N_781);
nand U834 (N_834,N_814,N_765);
or U835 (N_835,N_807,N_751);
nor U836 (N_836,N_768,N_759);
or U837 (N_837,N_794,N_795);
nand U838 (N_838,N_758,N_763);
nor U839 (N_839,N_817,N_774);
and U840 (N_840,N_804,N_782);
and U841 (N_841,N_766,N_769);
or U842 (N_842,N_780,N_762);
or U843 (N_843,N_793,N_801);
and U844 (N_844,N_799,N_812);
and U845 (N_845,N_761,N_777);
and U846 (N_846,N_773,N_811);
nor U847 (N_847,N_824,N_787);
nor U848 (N_848,N_753,N_752);
nor U849 (N_849,N_778,N_822);
nor U850 (N_850,N_783,N_785);
and U851 (N_851,N_760,N_816);
nor U852 (N_852,N_750,N_800);
nand U853 (N_853,N_809,N_791);
or U854 (N_854,N_775,N_798);
nand U855 (N_855,N_813,N_772);
xnor U856 (N_856,N_803,N_788);
nor U857 (N_857,N_819,N_764);
nor U858 (N_858,N_767,N_823);
and U859 (N_859,N_821,N_815);
nand U860 (N_860,N_792,N_810);
nand U861 (N_861,N_779,N_757);
nand U862 (N_862,N_818,N_789);
nor U863 (N_863,N_813,N_783);
xor U864 (N_864,N_786,N_811);
nor U865 (N_865,N_816,N_765);
nor U866 (N_866,N_756,N_786);
or U867 (N_867,N_789,N_804);
and U868 (N_868,N_758,N_760);
nor U869 (N_869,N_806,N_783);
nor U870 (N_870,N_790,N_757);
or U871 (N_871,N_760,N_802);
xnor U872 (N_872,N_781,N_757);
or U873 (N_873,N_818,N_788);
xor U874 (N_874,N_756,N_759);
nor U875 (N_875,N_808,N_824);
nand U876 (N_876,N_788,N_769);
and U877 (N_877,N_759,N_754);
nand U878 (N_878,N_775,N_805);
nand U879 (N_879,N_792,N_778);
or U880 (N_880,N_781,N_756);
xor U881 (N_881,N_816,N_807);
nand U882 (N_882,N_765,N_756);
or U883 (N_883,N_779,N_793);
and U884 (N_884,N_821,N_810);
nand U885 (N_885,N_753,N_805);
nand U886 (N_886,N_789,N_795);
nand U887 (N_887,N_811,N_775);
and U888 (N_888,N_750,N_754);
and U889 (N_889,N_754,N_797);
nand U890 (N_890,N_777,N_812);
and U891 (N_891,N_794,N_813);
or U892 (N_892,N_819,N_768);
and U893 (N_893,N_765,N_809);
nor U894 (N_894,N_798,N_795);
or U895 (N_895,N_762,N_768);
nor U896 (N_896,N_770,N_792);
nand U897 (N_897,N_765,N_817);
nor U898 (N_898,N_793,N_822);
nand U899 (N_899,N_810,N_761);
nand U900 (N_900,N_868,N_834);
nand U901 (N_901,N_874,N_842);
and U902 (N_902,N_898,N_867);
nor U903 (N_903,N_876,N_830);
and U904 (N_904,N_854,N_863);
and U905 (N_905,N_850,N_853);
nand U906 (N_906,N_884,N_878);
or U907 (N_907,N_858,N_846);
nand U908 (N_908,N_861,N_895);
nand U909 (N_909,N_827,N_882);
nand U910 (N_910,N_890,N_886);
and U911 (N_911,N_845,N_881);
nor U912 (N_912,N_828,N_894);
and U913 (N_913,N_844,N_856);
nand U914 (N_914,N_899,N_832);
and U915 (N_915,N_838,N_839);
nand U916 (N_916,N_826,N_829);
nor U917 (N_917,N_883,N_851);
and U918 (N_918,N_862,N_877);
nor U919 (N_919,N_860,N_825);
nor U920 (N_920,N_891,N_896);
and U921 (N_921,N_885,N_837);
and U922 (N_922,N_892,N_889);
and U923 (N_923,N_880,N_869);
and U924 (N_924,N_893,N_859);
nor U925 (N_925,N_831,N_887);
xnor U926 (N_926,N_897,N_840);
nor U927 (N_927,N_871,N_852);
or U928 (N_928,N_879,N_873);
nor U929 (N_929,N_875,N_866);
and U930 (N_930,N_870,N_847);
xnor U931 (N_931,N_857,N_836);
nor U932 (N_932,N_888,N_848);
nand U933 (N_933,N_835,N_849);
nand U934 (N_934,N_864,N_855);
and U935 (N_935,N_843,N_872);
or U936 (N_936,N_865,N_841);
nand U937 (N_937,N_833,N_873);
and U938 (N_938,N_894,N_836);
nand U939 (N_939,N_831,N_861);
nor U940 (N_940,N_827,N_893);
nand U941 (N_941,N_860,N_840);
nor U942 (N_942,N_829,N_847);
and U943 (N_943,N_843,N_899);
or U944 (N_944,N_898,N_889);
nand U945 (N_945,N_825,N_885);
xnor U946 (N_946,N_847,N_871);
or U947 (N_947,N_833,N_842);
nand U948 (N_948,N_841,N_894);
nand U949 (N_949,N_843,N_884);
nor U950 (N_950,N_858,N_876);
nor U951 (N_951,N_865,N_875);
nor U952 (N_952,N_876,N_857);
nor U953 (N_953,N_868,N_874);
or U954 (N_954,N_856,N_861);
or U955 (N_955,N_869,N_866);
and U956 (N_956,N_863,N_850);
and U957 (N_957,N_837,N_881);
nor U958 (N_958,N_826,N_871);
nor U959 (N_959,N_859,N_837);
nor U960 (N_960,N_852,N_847);
or U961 (N_961,N_828,N_873);
and U962 (N_962,N_888,N_855);
nand U963 (N_963,N_834,N_883);
and U964 (N_964,N_869,N_859);
nor U965 (N_965,N_882,N_894);
and U966 (N_966,N_879,N_883);
and U967 (N_967,N_850,N_848);
nand U968 (N_968,N_895,N_872);
and U969 (N_969,N_862,N_870);
nand U970 (N_970,N_885,N_867);
nand U971 (N_971,N_846,N_848);
nand U972 (N_972,N_885,N_898);
or U973 (N_973,N_874,N_854);
and U974 (N_974,N_876,N_863);
nand U975 (N_975,N_934,N_942);
and U976 (N_976,N_927,N_916);
nand U977 (N_977,N_943,N_974);
nor U978 (N_978,N_907,N_933);
and U979 (N_979,N_970,N_941);
and U980 (N_980,N_918,N_900);
or U981 (N_981,N_958,N_956);
nor U982 (N_982,N_950,N_953);
nand U983 (N_983,N_961,N_903);
nand U984 (N_984,N_968,N_919);
and U985 (N_985,N_931,N_922);
nand U986 (N_986,N_930,N_901);
or U987 (N_987,N_928,N_947);
or U988 (N_988,N_920,N_912);
nand U989 (N_989,N_910,N_905);
and U990 (N_990,N_967,N_938);
and U991 (N_991,N_973,N_929);
xnor U992 (N_992,N_906,N_969);
nand U993 (N_993,N_964,N_935);
nand U994 (N_994,N_957,N_923);
and U995 (N_995,N_904,N_914);
xnor U996 (N_996,N_925,N_959);
nand U997 (N_997,N_960,N_951);
xor U998 (N_998,N_908,N_966);
xnor U999 (N_999,N_936,N_902);
nor U1000 (N_1000,N_944,N_948);
nor U1001 (N_1001,N_924,N_909);
nor U1002 (N_1002,N_954,N_915);
or U1003 (N_1003,N_972,N_952);
or U1004 (N_1004,N_963,N_932);
nand U1005 (N_1005,N_971,N_939);
and U1006 (N_1006,N_962,N_926);
or U1007 (N_1007,N_946,N_937);
and U1008 (N_1008,N_965,N_917);
and U1009 (N_1009,N_921,N_955);
nor U1010 (N_1010,N_940,N_949);
nand U1011 (N_1011,N_913,N_945);
nor U1012 (N_1012,N_911,N_938);
or U1013 (N_1013,N_952,N_928);
or U1014 (N_1014,N_927,N_924);
and U1015 (N_1015,N_961,N_966);
nand U1016 (N_1016,N_946,N_913);
nand U1017 (N_1017,N_942,N_932);
nand U1018 (N_1018,N_974,N_937);
and U1019 (N_1019,N_906,N_955);
or U1020 (N_1020,N_902,N_926);
or U1021 (N_1021,N_956,N_954);
nor U1022 (N_1022,N_932,N_928);
and U1023 (N_1023,N_964,N_969);
nand U1024 (N_1024,N_932,N_935);
and U1025 (N_1025,N_910,N_933);
nor U1026 (N_1026,N_934,N_914);
or U1027 (N_1027,N_944,N_953);
or U1028 (N_1028,N_921,N_914);
and U1029 (N_1029,N_902,N_965);
xor U1030 (N_1030,N_901,N_966);
nor U1031 (N_1031,N_933,N_974);
or U1032 (N_1032,N_965,N_946);
nand U1033 (N_1033,N_932,N_944);
nor U1034 (N_1034,N_905,N_915);
and U1035 (N_1035,N_926,N_954);
nand U1036 (N_1036,N_951,N_956);
and U1037 (N_1037,N_906,N_901);
or U1038 (N_1038,N_939,N_958);
and U1039 (N_1039,N_907,N_971);
nand U1040 (N_1040,N_939,N_938);
or U1041 (N_1041,N_920,N_900);
nand U1042 (N_1042,N_924,N_973);
or U1043 (N_1043,N_969,N_952);
or U1044 (N_1044,N_961,N_956);
and U1045 (N_1045,N_932,N_957);
and U1046 (N_1046,N_910,N_925);
and U1047 (N_1047,N_910,N_917);
or U1048 (N_1048,N_910,N_935);
xnor U1049 (N_1049,N_956,N_974);
nor U1050 (N_1050,N_1048,N_1005);
or U1051 (N_1051,N_1047,N_977);
xor U1052 (N_1052,N_1002,N_1042);
xor U1053 (N_1053,N_978,N_1027);
and U1054 (N_1054,N_999,N_1024);
nor U1055 (N_1055,N_1017,N_1032);
and U1056 (N_1056,N_1014,N_1045);
and U1057 (N_1057,N_986,N_1011);
or U1058 (N_1058,N_1019,N_1033);
and U1059 (N_1059,N_1030,N_989);
nand U1060 (N_1060,N_997,N_981);
or U1061 (N_1061,N_993,N_1035);
or U1062 (N_1062,N_1001,N_992);
and U1063 (N_1063,N_1041,N_988);
and U1064 (N_1064,N_1007,N_983);
and U1065 (N_1065,N_1000,N_1029);
nand U1066 (N_1066,N_1049,N_1031);
nand U1067 (N_1067,N_1013,N_982);
nand U1068 (N_1068,N_1020,N_998);
nor U1069 (N_1069,N_980,N_1015);
and U1070 (N_1070,N_990,N_1038);
nor U1071 (N_1071,N_1025,N_1003);
or U1072 (N_1072,N_984,N_1016);
nand U1073 (N_1073,N_1004,N_1006);
nor U1074 (N_1074,N_1009,N_1028);
or U1075 (N_1075,N_1008,N_976);
and U1076 (N_1076,N_985,N_1036);
nand U1077 (N_1077,N_979,N_1026);
nor U1078 (N_1078,N_1046,N_1021);
nand U1079 (N_1079,N_1043,N_1018);
or U1080 (N_1080,N_1023,N_1039);
nor U1081 (N_1081,N_1037,N_1044);
or U1082 (N_1082,N_1010,N_994);
nand U1083 (N_1083,N_987,N_1040);
and U1084 (N_1084,N_991,N_996);
nor U1085 (N_1085,N_975,N_995);
or U1086 (N_1086,N_1034,N_1012);
nor U1087 (N_1087,N_1022,N_1009);
nor U1088 (N_1088,N_1031,N_1028);
or U1089 (N_1089,N_1003,N_994);
nand U1090 (N_1090,N_1001,N_1028);
or U1091 (N_1091,N_1035,N_985);
or U1092 (N_1092,N_1042,N_1038);
nor U1093 (N_1093,N_1042,N_1008);
nor U1094 (N_1094,N_1009,N_1033);
nor U1095 (N_1095,N_1008,N_985);
nand U1096 (N_1096,N_1043,N_1007);
xnor U1097 (N_1097,N_978,N_992);
and U1098 (N_1098,N_1011,N_984);
nand U1099 (N_1099,N_1012,N_1032);
nor U1100 (N_1100,N_1033,N_1022);
xor U1101 (N_1101,N_1003,N_977);
or U1102 (N_1102,N_1035,N_996);
nor U1103 (N_1103,N_983,N_992);
or U1104 (N_1104,N_1005,N_1002);
nand U1105 (N_1105,N_1026,N_984);
nor U1106 (N_1106,N_1032,N_1027);
nor U1107 (N_1107,N_1005,N_1012);
or U1108 (N_1108,N_1020,N_984);
or U1109 (N_1109,N_992,N_1032);
and U1110 (N_1110,N_978,N_1028);
or U1111 (N_1111,N_990,N_1020);
and U1112 (N_1112,N_979,N_1002);
nand U1113 (N_1113,N_992,N_999);
and U1114 (N_1114,N_1046,N_1027);
nand U1115 (N_1115,N_1018,N_1023);
or U1116 (N_1116,N_1001,N_990);
nand U1117 (N_1117,N_1019,N_989);
and U1118 (N_1118,N_1031,N_1033);
nand U1119 (N_1119,N_991,N_1029);
or U1120 (N_1120,N_1046,N_1000);
xnor U1121 (N_1121,N_1039,N_1005);
nand U1122 (N_1122,N_989,N_999);
nand U1123 (N_1123,N_995,N_1048);
and U1124 (N_1124,N_1014,N_1022);
nor U1125 (N_1125,N_1087,N_1063);
or U1126 (N_1126,N_1121,N_1067);
and U1127 (N_1127,N_1081,N_1077);
nor U1128 (N_1128,N_1113,N_1120);
nand U1129 (N_1129,N_1057,N_1096);
nor U1130 (N_1130,N_1099,N_1101);
nand U1131 (N_1131,N_1088,N_1051);
nor U1132 (N_1132,N_1050,N_1094);
nor U1133 (N_1133,N_1085,N_1107);
or U1134 (N_1134,N_1054,N_1102);
or U1135 (N_1135,N_1072,N_1083);
nor U1136 (N_1136,N_1103,N_1084);
nor U1137 (N_1137,N_1119,N_1068);
and U1138 (N_1138,N_1073,N_1055);
and U1139 (N_1139,N_1086,N_1082);
and U1140 (N_1140,N_1109,N_1114);
nand U1141 (N_1141,N_1065,N_1052);
nand U1142 (N_1142,N_1122,N_1069);
nand U1143 (N_1143,N_1108,N_1123);
nor U1144 (N_1144,N_1059,N_1116);
nor U1145 (N_1145,N_1091,N_1076);
or U1146 (N_1146,N_1062,N_1053);
and U1147 (N_1147,N_1070,N_1100);
and U1148 (N_1148,N_1080,N_1093);
and U1149 (N_1149,N_1056,N_1089);
and U1150 (N_1150,N_1118,N_1075);
or U1151 (N_1151,N_1124,N_1090);
xnor U1152 (N_1152,N_1066,N_1097);
and U1153 (N_1153,N_1098,N_1115);
or U1154 (N_1154,N_1117,N_1078);
or U1155 (N_1155,N_1106,N_1064);
and U1156 (N_1156,N_1061,N_1111);
and U1157 (N_1157,N_1079,N_1105);
and U1158 (N_1158,N_1092,N_1071);
nand U1159 (N_1159,N_1095,N_1060);
nor U1160 (N_1160,N_1110,N_1104);
nand U1161 (N_1161,N_1074,N_1058);
nand U1162 (N_1162,N_1112,N_1074);
and U1163 (N_1163,N_1062,N_1104);
nand U1164 (N_1164,N_1075,N_1078);
and U1165 (N_1165,N_1102,N_1058);
xor U1166 (N_1166,N_1124,N_1057);
nor U1167 (N_1167,N_1065,N_1123);
nand U1168 (N_1168,N_1053,N_1105);
nand U1169 (N_1169,N_1053,N_1107);
or U1170 (N_1170,N_1077,N_1108);
xor U1171 (N_1171,N_1091,N_1092);
nor U1172 (N_1172,N_1072,N_1090);
nor U1173 (N_1173,N_1098,N_1083);
nor U1174 (N_1174,N_1099,N_1092);
nor U1175 (N_1175,N_1124,N_1097);
nand U1176 (N_1176,N_1084,N_1069);
nand U1177 (N_1177,N_1087,N_1097);
nor U1178 (N_1178,N_1098,N_1101);
or U1179 (N_1179,N_1106,N_1059);
nor U1180 (N_1180,N_1060,N_1104);
or U1181 (N_1181,N_1082,N_1053);
or U1182 (N_1182,N_1073,N_1100);
nand U1183 (N_1183,N_1051,N_1099);
nand U1184 (N_1184,N_1050,N_1089);
and U1185 (N_1185,N_1100,N_1075);
and U1186 (N_1186,N_1104,N_1090);
nor U1187 (N_1187,N_1099,N_1055);
xnor U1188 (N_1188,N_1067,N_1095);
nor U1189 (N_1189,N_1103,N_1051);
and U1190 (N_1190,N_1104,N_1100);
nor U1191 (N_1191,N_1092,N_1064);
nor U1192 (N_1192,N_1065,N_1107);
or U1193 (N_1193,N_1121,N_1071);
nor U1194 (N_1194,N_1084,N_1061);
nor U1195 (N_1195,N_1092,N_1119);
and U1196 (N_1196,N_1063,N_1050);
and U1197 (N_1197,N_1074,N_1091);
and U1198 (N_1198,N_1106,N_1078);
and U1199 (N_1199,N_1105,N_1123);
and U1200 (N_1200,N_1195,N_1139);
nand U1201 (N_1201,N_1162,N_1175);
and U1202 (N_1202,N_1199,N_1165);
nand U1203 (N_1203,N_1152,N_1130);
or U1204 (N_1204,N_1154,N_1166);
and U1205 (N_1205,N_1172,N_1183);
and U1206 (N_1206,N_1136,N_1191);
nor U1207 (N_1207,N_1147,N_1168);
nor U1208 (N_1208,N_1131,N_1197);
nand U1209 (N_1209,N_1148,N_1198);
nand U1210 (N_1210,N_1170,N_1143);
and U1211 (N_1211,N_1138,N_1187);
nor U1212 (N_1212,N_1126,N_1179);
nor U1213 (N_1213,N_1185,N_1164);
nor U1214 (N_1214,N_1156,N_1159);
and U1215 (N_1215,N_1176,N_1137);
or U1216 (N_1216,N_1140,N_1142);
nor U1217 (N_1217,N_1155,N_1173);
or U1218 (N_1218,N_1149,N_1153);
nor U1219 (N_1219,N_1145,N_1134);
and U1220 (N_1220,N_1186,N_1188);
nor U1221 (N_1221,N_1163,N_1141);
nand U1222 (N_1222,N_1160,N_1157);
or U1223 (N_1223,N_1150,N_1190);
nor U1224 (N_1224,N_1167,N_1161);
nand U1225 (N_1225,N_1184,N_1192);
nand U1226 (N_1226,N_1125,N_1193);
nor U1227 (N_1227,N_1133,N_1144);
or U1228 (N_1228,N_1135,N_1174);
or U1229 (N_1229,N_1189,N_1171);
and U1230 (N_1230,N_1182,N_1127);
or U1231 (N_1231,N_1177,N_1146);
nand U1232 (N_1232,N_1178,N_1158);
nand U1233 (N_1233,N_1132,N_1169);
nand U1234 (N_1234,N_1180,N_1196);
or U1235 (N_1235,N_1129,N_1194);
and U1236 (N_1236,N_1128,N_1181);
nand U1237 (N_1237,N_1151,N_1150);
or U1238 (N_1238,N_1171,N_1129);
nor U1239 (N_1239,N_1184,N_1172);
and U1240 (N_1240,N_1158,N_1164);
and U1241 (N_1241,N_1159,N_1190);
or U1242 (N_1242,N_1138,N_1192);
nand U1243 (N_1243,N_1198,N_1169);
or U1244 (N_1244,N_1163,N_1164);
and U1245 (N_1245,N_1170,N_1129);
and U1246 (N_1246,N_1172,N_1186);
nand U1247 (N_1247,N_1133,N_1148);
and U1248 (N_1248,N_1127,N_1179);
nand U1249 (N_1249,N_1184,N_1127);
or U1250 (N_1250,N_1157,N_1168);
and U1251 (N_1251,N_1182,N_1191);
nor U1252 (N_1252,N_1145,N_1176);
nor U1253 (N_1253,N_1146,N_1133);
nor U1254 (N_1254,N_1145,N_1198);
nand U1255 (N_1255,N_1148,N_1135);
nor U1256 (N_1256,N_1194,N_1133);
nor U1257 (N_1257,N_1142,N_1130);
and U1258 (N_1258,N_1170,N_1158);
or U1259 (N_1259,N_1151,N_1127);
nor U1260 (N_1260,N_1133,N_1127);
nor U1261 (N_1261,N_1166,N_1195);
nand U1262 (N_1262,N_1143,N_1145);
or U1263 (N_1263,N_1189,N_1137);
or U1264 (N_1264,N_1158,N_1141);
nor U1265 (N_1265,N_1140,N_1181);
nor U1266 (N_1266,N_1177,N_1149);
or U1267 (N_1267,N_1171,N_1141);
nor U1268 (N_1268,N_1177,N_1162);
or U1269 (N_1269,N_1188,N_1139);
nand U1270 (N_1270,N_1166,N_1172);
and U1271 (N_1271,N_1136,N_1190);
or U1272 (N_1272,N_1170,N_1180);
or U1273 (N_1273,N_1178,N_1140);
nand U1274 (N_1274,N_1151,N_1168);
and U1275 (N_1275,N_1223,N_1271);
and U1276 (N_1276,N_1211,N_1261);
nor U1277 (N_1277,N_1274,N_1204);
or U1278 (N_1278,N_1265,N_1267);
or U1279 (N_1279,N_1221,N_1243);
nand U1280 (N_1280,N_1231,N_1242);
nand U1281 (N_1281,N_1232,N_1252);
nand U1282 (N_1282,N_1255,N_1247);
nor U1283 (N_1283,N_1260,N_1227);
and U1284 (N_1284,N_1233,N_1206);
or U1285 (N_1285,N_1215,N_1225);
and U1286 (N_1286,N_1264,N_1210);
and U1287 (N_1287,N_1237,N_1262);
nand U1288 (N_1288,N_1244,N_1205);
nand U1289 (N_1289,N_1250,N_1218);
and U1290 (N_1290,N_1251,N_1238);
nor U1291 (N_1291,N_1272,N_1202);
and U1292 (N_1292,N_1209,N_1201);
nand U1293 (N_1293,N_1222,N_1236);
and U1294 (N_1294,N_1200,N_1203);
nand U1295 (N_1295,N_1273,N_1214);
nand U1296 (N_1296,N_1256,N_1220);
and U1297 (N_1297,N_1213,N_1240);
or U1298 (N_1298,N_1245,N_1259);
or U1299 (N_1299,N_1266,N_1254);
nor U1300 (N_1300,N_1268,N_1253);
nand U1301 (N_1301,N_1217,N_1224);
nand U1302 (N_1302,N_1235,N_1263);
nand U1303 (N_1303,N_1212,N_1207);
or U1304 (N_1304,N_1219,N_1246);
and U1305 (N_1305,N_1229,N_1241);
nor U1306 (N_1306,N_1270,N_1248);
xor U1307 (N_1307,N_1249,N_1230);
nand U1308 (N_1308,N_1226,N_1257);
or U1309 (N_1309,N_1228,N_1208);
or U1310 (N_1310,N_1269,N_1239);
and U1311 (N_1311,N_1234,N_1216);
and U1312 (N_1312,N_1258,N_1209);
and U1313 (N_1313,N_1262,N_1252);
or U1314 (N_1314,N_1220,N_1236);
nor U1315 (N_1315,N_1233,N_1240);
or U1316 (N_1316,N_1227,N_1206);
and U1317 (N_1317,N_1232,N_1205);
nor U1318 (N_1318,N_1268,N_1228);
or U1319 (N_1319,N_1240,N_1261);
nand U1320 (N_1320,N_1215,N_1235);
or U1321 (N_1321,N_1232,N_1234);
or U1322 (N_1322,N_1244,N_1271);
nor U1323 (N_1323,N_1213,N_1208);
and U1324 (N_1324,N_1233,N_1230);
and U1325 (N_1325,N_1201,N_1214);
nand U1326 (N_1326,N_1216,N_1245);
nand U1327 (N_1327,N_1224,N_1254);
and U1328 (N_1328,N_1224,N_1236);
or U1329 (N_1329,N_1256,N_1259);
nor U1330 (N_1330,N_1204,N_1219);
or U1331 (N_1331,N_1256,N_1232);
nand U1332 (N_1332,N_1256,N_1248);
and U1333 (N_1333,N_1263,N_1224);
nor U1334 (N_1334,N_1235,N_1202);
xor U1335 (N_1335,N_1272,N_1214);
or U1336 (N_1336,N_1263,N_1208);
nand U1337 (N_1337,N_1200,N_1224);
and U1338 (N_1338,N_1209,N_1271);
nand U1339 (N_1339,N_1212,N_1256);
or U1340 (N_1340,N_1211,N_1238);
nand U1341 (N_1341,N_1231,N_1221);
or U1342 (N_1342,N_1225,N_1211);
nor U1343 (N_1343,N_1215,N_1236);
or U1344 (N_1344,N_1215,N_1248);
and U1345 (N_1345,N_1203,N_1255);
nand U1346 (N_1346,N_1230,N_1231);
or U1347 (N_1347,N_1273,N_1253);
nor U1348 (N_1348,N_1210,N_1266);
nand U1349 (N_1349,N_1245,N_1243);
or U1350 (N_1350,N_1278,N_1276);
and U1351 (N_1351,N_1321,N_1304);
or U1352 (N_1352,N_1338,N_1337);
nand U1353 (N_1353,N_1290,N_1309);
and U1354 (N_1354,N_1296,N_1341);
or U1355 (N_1355,N_1311,N_1326);
nor U1356 (N_1356,N_1319,N_1318);
nand U1357 (N_1357,N_1335,N_1306);
nor U1358 (N_1358,N_1283,N_1284);
nand U1359 (N_1359,N_1330,N_1313);
nor U1360 (N_1360,N_1292,N_1339);
nor U1361 (N_1361,N_1316,N_1343);
nand U1362 (N_1362,N_1295,N_1324);
nand U1363 (N_1363,N_1345,N_1346);
or U1364 (N_1364,N_1302,N_1323);
nor U1365 (N_1365,N_1314,N_1308);
or U1366 (N_1366,N_1320,N_1348);
nand U1367 (N_1367,N_1277,N_1327);
nor U1368 (N_1368,N_1286,N_1289);
xnor U1369 (N_1369,N_1300,N_1344);
or U1370 (N_1370,N_1303,N_1333);
and U1371 (N_1371,N_1294,N_1331);
and U1372 (N_1372,N_1297,N_1310);
or U1373 (N_1373,N_1293,N_1279);
nand U1374 (N_1374,N_1305,N_1325);
and U1375 (N_1375,N_1332,N_1288);
nand U1376 (N_1376,N_1280,N_1301);
nand U1377 (N_1377,N_1281,N_1299);
nor U1378 (N_1378,N_1342,N_1329);
nand U1379 (N_1379,N_1322,N_1336);
nor U1380 (N_1380,N_1282,N_1315);
nor U1381 (N_1381,N_1287,N_1312);
or U1382 (N_1382,N_1291,N_1349);
nand U1383 (N_1383,N_1317,N_1307);
nand U1384 (N_1384,N_1275,N_1328);
nand U1385 (N_1385,N_1285,N_1347);
nor U1386 (N_1386,N_1340,N_1298);
nor U1387 (N_1387,N_1334,N_1284);
nor U1388 (N_1388,N_1308,N_1341);
nand U1389 (N_1389,N_1316,N_1327);
or U1390 (N_1390,N_1324,N_1345);
and U1391 (N_1391,N_1285,N_1310);
nand U1392 (N_1392,N_1276,N_1338);
or U1393 (N_1393,N_1280,N_1345);
and U1394 (N_1394,N_1317,N_1325);
and U1395 (N_1395,N_1328,N_1289);
and U1396 (N_1396,N_1349,N_1298);
nand U1397 (N_1397,N_1294,N_1317);
nor U1398 (N_1398,N_1310,N_1293);
xnor U1399 (N_1399,N_1308,N_1332);
nand U1400 (N_1400,N_1319,N_1294);
or U1401 (N_1401,N_1332,N_1328);
and U1402 (N_1402,N_1287,N_1296);
and U1403 (N_1403,N_1309,N_1324);
or U1404 (N_1404,N_1326,N_1300);
nand U1405 (N_1405,N_1344,N_1309);
xnor U1406 (N_1406,N_1314,N_1290);
nor U1407 (N_1407,N_1279,N_1277);
or U1408 (N_1408,N_1343,N_1310);
nand U1409 (N_1409,N_1299,N_1332);
nand U1410 (N_1410,N_1312,N_1315);
xnor U1411 (N_1411,N_1299,N_1326);
nor U1412 (N_1412,N_1310,N_1282);
or U1413 (N_1413,N_1315,N_1287);
or U1414 (N_1414,N_1338,N_1327);
or U1415 (N_1415,N_1295,N_1299);
nor U1416 (N_1416,N_1293,N_1289);
and U1417 (N_1417,N_1306,N_1307);
nor U1418 (N_1418,N_1347,N_1303);
nor U1419 (N_1419,N_1301,N_1345);
nand U1420 (N_1420,N_1321,N_1296);
nand U1421 (N_1421,N_1318,N_1333);
or U1422 (N_1422,N_1311,N_1279);
nor U1423 (N_1423,N_1335,N_1329);
nor U1424 (N_1424,N_1344,N_1329);
nor U1425 (N_1425,N_1363,N_1359);
xnor U1426 (N_1426,N_1378,N_1423);
or U1427 (N_1427,N_1418,N_1389);
nand U1428 (N_1428,N_1395,N_1362);
nor U1429 (N_1429,N_1394,N_1376);
or U1430 (N_1430,N_1406,N_1367);
nor U1431 (N_1431,N_1401,N_1390);
and U1432 (N_1432,N_1407,N_1360);
nor U1433 (N_1433,N_1405,N_1409);
nor U1434 (N_1434,N_1420,N_1412);
or U1435 (N_1435,N_1366,N_1396);
and U1436 (N_1436,N_1402,N_1357);
nand U1437 (N_1437,N_1391,N_1419);
and U1438 (N_1438,N_1421,N_1384);
nand U1439 (N_1439,N_1404,N_1424);
and U1440 (N_1440,N_1386,N_1369);
nand U1441 (N_1441,N_1356,N_1358);
and U1442 (N_1442,N_1416,N_1375);
nor U1443 (N_1443,N_1414,N_1364);
nand U1444 (N_1444,N_1399,N_1388);
nand U1445 (N_1445,N_1377,N_1361);
nand U1446 (N_1446,N_1400,N_1372);
and U1447 (N_1447,N_1380,N_1371);
or U1448 (N_1448,N_1422,N_1411);
nor U1449 (N_1449,N_1374,N_1393);
or U1450 (N_1450,N_1354,N_1351);
or U1451 (N_1451,N_1392,N_1413);
nor U1452 (N_1452,N_1382,N_1385);
nor U1453 (N_1453,N_1410,N_1373);
or U1454 (N_1454,N_1403,N_1381);
and U1455 (N_1455,N_1387,N_1352);
and U1456 (N_1456,N_1408,N_1350);
nand U1457 (N_1457,N_1370,N_1417);
or U1458 (N_1458,N_1368,N_1383);
nand U1459 (N_1459,N_1353,N_1398);
nor U1460 (N_1460,N_1397,N_1365);
nand U1461 (N_1461,N_1355,N_1415);
and U1462 (N_1462,N_1379,N_1406);
nor U1463 (N_1463,N_1363,N_1352);
nor U1464 (N_1464,N_1399,N_1401);
or U1465 (N_1465,N_1424,N_1400);
nand U1466 (N_1466,N_1371,N_1373);
nor U1467 (N_1467,N_1363,N_1382);
and U1468 (N_1468,N_1414,N_1354);
or U1469 (N_1469,N_1416,N_1419);
nor U1470 (N_1470,N_1418,N_1386);
nand U1471 (N_1471,N_1369,N_1400);
nor U1472 (N_1472,N_1416,N_1393);
or U1473 (N_1473,N_1380,N_1386);
nand U1474 (N_1474,N_1365,N_1357);
and U1475 (N_1475,N_1385,N_1403);
and U1476 (N_1476,N_1356,N_1367);
and U1477 (N_1477,N_1422,N_1393);
nand U1478 (N_1478,N_1360,N_1370);
nand U1479 (N_1479,N_1419,N_1396);
or U1480 (N_1480,N_1363,N_1413);
or U1481 (N_1481,N_1402,N_1387);
and U1482 (N_1482,N_1410,N_1419);
and U1483 (N_1483,N_1410,N_1358);
and U1484 (N_1484,N_1366,N_1376);
or U1485 (N_1485,N_1351,N_1353);
or U1486 (N_1486,N_1374,N_1421);
or U1487 (N_1487,N_1374,N_1405);
and U1488 (N_1488,N_1359,N_1388);
nand U1489 (N_1489,N_1409,N_1424);
and U1490 (N_1490,N_1424,N_1389);
and U1491 (N_1491,N_1423,N_1399);
or U1492 (N_1492,N_1400,N_1380);
nor U1493 (N_1493,N_1358,N_1424);
nor U1494 (N_1494,N_1364,N_1408);
nand U1495 (N_1495,N_1418,N_1402);
nor U1496 (N_1496,N_1402,N_1361);
or U1497 (N_1497,N_1385,N_1365);
and U1498 (N_1498,N_1408,N_1399);
or U1499 (N_1499,N_1382,N_1395);
nor U1500 (N_1500,N_1435,N_1455);
nand U1501 (N_1501,N_1428,N_1453);
nor U1502 (N_1502,N_1440,N_1499);
nor U1503 (N_1503,N_1490,N_1438);
nor U1504 (N_1504,N_1464,N_1469);
and U1505 (N_1505,N_1462,N_1492);
nor U1506 (N_1506,N_1463,N_1447);
nor U1507 (N_1507,N_1479,N_1432);
or U1508 (N_1508,N_1445,N_1461);
nand U1509 (N_1509,N_1480,N_1484);
or U1510 (N_1510,N_1457,N_1491);
nor U1511 (N_1511,N_1497,N_1446);
or U1512 (N_1512,N_1474,N_1486);
nand U1513 (N_1513,N_1460,N_1430);
or U1514 (N_1514,N_1441,N_1465);
nand U1515 (N_1515,N_1431,N_1475);
and U1516 (N_1516,N_1470,N_1448);
or U1517 (N_1517,N_1483,N_1487);
or U1518 (N_1518,N_1485,N_1496);
nor U1519 (N_1519,N_1452,N_1425);
or U1520 (N_1520,N_1439,N_1459);
nand U1521 (N_1521,N_1426,N_1493);
and U1522 (N_1522,N_1488,N_1449);
nor U1523 (N_1523,N_1442,N_1456);
nor U1524 (N_1524,N_1471,N_1466);
and U1525 (N_1525,N_1444,N_1436);
and U1526 (N_1526,N_1450,N_1489);
and U1527 (N_1527,N_1458,N_1472);
or U1528 (N_1528,N_1434,N_1498);
and U1529 (N_1529,N_1451,N_1473);
or U1530 (N_1530,N_1427,N_1477);
or U1531 (N_1531,N_1433,N_1443);
nor U1532 (N_1532,N_1468,N_1495);
nor U1533 (N_1533,N_1494,N_1478);
nand U1534 (N_1534,N_1437,N_1467);
or U1535 (N_1535,N_1454,N_1429);
nand U1536 (N_1536,N_1481,N_1482);
and U1537 (N_1537,N_1476,N_1441);
nand U1538 (N_1538,N_1470,N_1468);
nand U1539 (N_1539,N_1487,N_1481);
nor U1540 (N_1540,N_1471,N_1483);
and U1541 (N_1541,N_1470,N_1478);
nand U1542 (N_1542,N_1484,N_1491);
or U1543 (N_1543,N_1480,N_1478);
nand U1544 (N_1544,N_1427,N_1481);
nand U1545 (N_1545,N_1490,N_1442);
and U1546 (N_1546,N_1428,N_1465);
and U1547 (N_1547,N_1485,N_1466);
nor U1548 (N_1548,N_1430,N_1488);
nor U1549 (N_1549,N_1497,N_1447);
or U1550 (N_1550,N_1427,N_1464);
nor U1551 (N_1551,N_1492,N_1490);
xor U1552 (N_1552,N_1465,N_1457);
nand U1553 (N_1553,N_1468,N_1444);
or U1554 (N_1554,N_1437,N_1497);
or U1555 (N_1555,N_1436,N_1498);
nor U1556 (N_1556,N_1443,N_1435);
xnor U1557 (N_1557,N_1469,N_1496);
and U1558 (N_1558,N_1461,N_1467);
nand U1559 (N_1559,N_1426,N_1491);
and U1560 (N_1560,N_1479,N_1456);
and U1561 (N_1561,N_1471,N_1448);
nand U1562 (N_1562,N_1426,N_1425);
or U1563 (N_1563,N_1481,N_1429);
nand U1564 (N_1564,N_1440,N_1448);
or U1565 (N_1565,N_1499,N_1484);
or U1566 (N_1566,N_1445,N_1438);
xnor U1567 (N_1567,N_1464,N_1442);
nor U1568 (N_1568,N_1457,N_1469);
or U1569 (N_1569,N_1459,N_1474);
and U1570 (N_1570,N_1427,N_1487);
nor U1571 (N_1571,N_1486,N_1494);
or U1572 (N_1572,N_1442,N_1438);
nor U1573 (N_1573,N_1463,N_1480);
or U1574 (N_1574,N_1433,N_1471);
xnor U1575 (N_1575,N_1555,N_1531);
and U1576 (N_1576,N_1556,N_1518);
and U1577 (N_1577,N_1539,N_1560);
nand U1578 (N_1578,N_1500,N_1559);
nand U1579 (N_1579,N_1512,N_1508);
nor U1580 (N_1580,N_1525,N_1543);
nand U1581 (N_1581,N_1538,N_1545);
and U1582 (N_1582,N_1557,N_1529);
nand U1583 (N_1583,N_1553,N_1507);
and U1584 (N_1584,N_1527,N_1572);
xnor U1585 (N_1585,N_1547,N_1533);
and U1586 (N_1586,N_1510,N_1534);
or U1587 (N_1587,N_1532,N_1528);
nand U1588 (N_1588,N_1546,N_1561);
or U1589 (N_1589,N_1536,N_1535);
and U1590 (N_1590,N_1554,N_1570);
and U1591 (N_1591,N_1564,N_1573);
or U1592 (N_1592,N_1523,N_1511);
nor U1593 (N_1593,N_1524,N_1503);
or U1594 (N_1594,N_1541,N_1537);
nor U1595 (N_1595,N_1549,N_1544);
or U1596 (N_1596,N_1521,N_1522);
and U1597 (N_1597,N_1552,N_1520);
nand U1598 (N_1598,N_1501,N_1516);
and U1599 (N_1599,N_1574,N_1567);
and U1600 (N_1600,N_1569,N_1526);
and U1601 (N_1601,N_1565,N_1513);
xnor U1602 (N_1602,N_1509,N_1542);
nor U1603 (N_1603,N_1551,N_1568);
or U1604 (N_1604,N_1530,N_1504);
nor U1605 (N_1605,N_1558,N_1514);
and U1606 (N_1606,N_1517,N_1562);
nor U1607 (N_1607,N_1506,N_1548);
or U1608 (N_1608,N_1571,N_1515);
nand U1609 (N_1609,N_1505,N_1540);
and U1610 (N_1610,N_1563,N_1519);
and U1611 (N_1611,N_1502,N_1566);
nor U1612 (N_1612,N_1550,N_1555);
xnor U1613 (N_1613,N_1510,N_1550);
nor U1614 (N_1614,N_1528,N_1565);
or U1615 (N_1615,N_1555,N_1534);
and U1616 (N_1616,N_1557,N_1545);
nand U1617 (N_1617,N_1560,N_1557);
or U1618 (N_1618,N_1537,N_1553);
xnor U1619 (N_1619,N_1549,N_1535);
and U1620 (N_1620,N_1540,N_1572);
or U1621 (N_1621,N_1532,N_1504);
or U1622 (N_1622,N_1523,N_1573);
or U1623 (N_1623,N_1549,N_1533);
and U1624 (N_1624,N_1536,N_1514);
nand U1625 (N_1625,N_1569,N_1572);
or U1626 (N_1626,N_1507,N_1512);
and U1627 (N_1627,N_1545,N_1558);
nor U1628 (N_1628,N_1529,N_1502);
and U1629 (N_1629,N_1549,N_1537);
nand U1630 (N_1630,N_1552,N_1571);
and U1631 (N_1631,N_1506,N_1510);
or U1632 (N_1632,N_1565,N_1506);
and U1633 (N_1633,N_1568,N_1512);
or U1634 (N_1634,N_1532,N_1505);
nor U1635 (N_1635,N_1520,N_1504);
xor U1636 (N_1636,N_1537,N_1500);
nand U1637 (N_1637,N_1559,N_1561);
and U1638 (N_1638,N_1555,N_1508);
nand U1639 (N_1639,N_1501,N_1543);
nand U1640 (N_1640,N_1530,N_1510);
nor U1641 (N_1641,N_1518,N_1563);
and U1642 (N_1642,N_1507,N_1554);
nor U1643 (N_1643,N_1534,N_1537);
nand U1644 (N_1644,N_1530,N_1508);
nor U1645 (N_1645,N_1553,N_1503);
and U1646 (N_1646,N_1501,N_1510);
nor U1647 (N_1647,N_1537,N_1556);
xnor U1648 (N_1648,N_1505,N_1515);
nand U1649 (N_1649,N_1526,N_1571);
and U1650 (N_1650,N_1632,N_1640);
xor U1651 (N_1651,N_1630,N_1596);
or U1652 (N_1652,N_1631,N_1614);
and U1653 (N_1653,N_1599,N_1633);
or U1654 (N_1654,N_1635,N_1604);
or U1655 (N_1655,N_1605,N_1585);
or U1656 (N_1656,N_1649,N_1611);
xnor U1657 (N_1657,N_1638,N_1641);
or U1658 (N_1658,N_1646,N_1592);
nor U1659 (N_1659,N_1634,N_1576);
nor U1660 (N_1660,N_1577,N_1647);
or U1661 (N_1661,N_1618,N_1582);
nand U1662 (N_1662,N_1627,N_1623);
nor U1663 (N_1663,N_1579,N_1642);
or U1664 (N_1664,N_1603,N_1602);
xor U1665 (N_1665,N_1607,N_1598);
nand U1666 (N_1666,N_1593,N_1619);
or U1667 (N_1667,N_1586,N_1588);
nor U1668 (N_1668,N_1626,N_1628);
and U1669 (N_1669,N_1648,N_1591);
nand U1670 (N_1670,N_1644,N_1590);
and U1671 (N_1671,N_1600,N_1615);
or U1672 (N_1672,N_1620,N_1637);
and U1673 (N_1673,N_1621,N_1580);
nor U1674 (N_1674,N_1597,N_1581);
nor U1675 (N_1675,N_1622,N_1583);
nand U1676 (N_1676,N_1629,N_1643);
nor U1677 (N_1677,N_1625,N_1636);
nand U1678 (N_1678,N_1616,N_1595);
nand U1679 (N_1679,N_1624,N_1612);
nand U1680 (N_1680,N_1587,N_1639);
nor U1681 (N_1681,N_1610,N_1609);
or U1682 (N_1682,N_1584,N_1645);
and U1683 (N_1683,N_1613,N_1606);
nand U1684 (N_1684,N_1589,N_1601);
nor U1685 (N_1685,N_1575,N_1617);
and U1686 (N_1686,N_1594,N_1608);
or U1687 (N_1687,N_1578,N_1583);
and U1688 (N_1688,N_1604,N_1578);
nand U1689 (N_1689,N_1593,N_1627);
xnor U1690 (N_1690,N_1593,N_1583);
nor U1691 (N_1691,N_1599,N_1594);
nor U1692 (N_1692,N_1629,N_1611);
nor U1693 (N_1693,N_1597,N_1623);
and U1694 (N_1694,N_1637,N_1590);
nor U1695 (N_1695,N_1639,N_1634);
or U1696 (N_1696,N_1598,N_1575);
nand U1697 (N_1697,N_1614,N_1642);
or U1698 (N_1698,N_1586,N_1621);
nor U1699 (N_1699,N_1587,N_1622);
nor U1700 (N_1700,N_1587,N_1582);
or U1701 (N_1701,N_1606,N_1615);
and U1702 (N_1702,N_1576,N_1583);
xnor U1703 (N_1703,N_1630,N_1609);
nand U1704 (N_1704,N_1633,N_1631);
and U1705 (N_1705,N_1583,N_1628);
or U1706 (N_1706,N_1588,N_1644);
or U1707 (N_1707,N_1578,N_1595);
nor U1708 (N_1708,N_1575,N_1590);
nand U1709 (N_1709,N_1608,N_1591);
nand U1710 (N_1710,N_1577,N_1636);
and U1711 (N_1711,N_1622,N_1591);
nand U1712 (N_1712,N_1609,N_1582);
and U1713 (N_1713,N_1636,N_1588);
and U1714 (N_1714,N_1600,N_1605);
nor U1715 (N_1715,N_1580,N_1581);
or U1716 (N_1716,N_1648,N_1617);
or U1717 (N_1717,N_1591,N_1632);
nor U1718 (N_1718,N_1594,N_1579);
nor U1719 (N_1719,N_1627,N_1602);
or U1720 (N_1720,N_1629,N_1631);
and U1721 (N_1721,N_1647,N_1607);
nor U1722 (N_1722,N_1603,N_1611);
nor U1723 (N_1723,N_1575,N_1616);
nor U1724 (N_1724,N_1633,N_1596);
nor U1725 (N_1725,N_1689,N_1711);
and U1726 (N_1726,N_1660,N_1668);
or U1727 (N_1727,N_1714,N_1656);
nor U1728 (N_1728,N_1699,N_1708);
and U1729 (N_1729,N_1710,N_1722);
nand U1730 (N_1730,N_1700,N_1667);
nand U1731 (N_1731,N_1674,N_1658);
nor U1732 (N_1732,N_1709,N_1653);
nor U1733 (N_1733,N_1695,N_1694);
nand U1734 (N_1734,N_1696,N_1665);
nor U1735 (N_1735,N_1664,N_1712);
nor U1736 (N_1736,N_1672,N_1661);
and U1737 (N_1737,N_1704,N_1703);
and U1738 (N_1738,N_1720,N_1680);
and U1739 (N_1739,N_1678,N_1702);
and U1740 (N_1740,N_1697,N_1651);
and U1741 (N_1741,N_1673,N_1721);
nand U1742 (N_1742,N_1671,N_1663);
nor U1743 (N_1743,N_1676,N_1655);
nand U1744 (N_1744,N_1690,N_1669);
and U1745 (N_1745,N_1705,N_1713);
nor U1746 (N_1746,N_1657,N_1715);
nand U1747 (N_1747,N_1723,N_1666);
xnor U1748 (N_1748,N_1686,N_1687);
or U1749 (N_1749,N_1693,N_1677);
and U1750 (N_1750,N_1692,N_1650);
and U1751 (N_1751,N_1652,N_1716);
or U1752 (N_1752,N_1684,N_1724);
nor U1753 (N_1753,N_1682,N_1701);
or U1754 (N_1754,N_1681,N_1679);
xnor U1755 (N_1755,N_1662,N_1719);
and U1756 (N_1756,N_1654,N_1683);
nor U1757 (N_1757,N_1691,N_1698);
and U1758 (N_1758,N_1675,N_1707);
and U1759 (N_1759,N_1717,N_1685);
or U1760 (N_1760,N_1659,N_1688);
nor U1761 (N_1761,N_1670,N_1718);
or U1762 (N_1762,N_1706,N_1719);
nand U1763 (N_1763,N_1690,N_1660);
or U1764 (N_1764,N_1667,N_1664);
or U1765 (N_1765,N_1720,N_1682);
nor U1766 (N_1766,N_1656,N_1701);
and U1767 (N_1767,N_1713,N_1699);
or U1768 (N_1768,N_1664,N_1658);
or U1769 (N_1769,N_1650,N_1707);
and U1770 (N_1770,N_1684,N_1677);
and U1771 (N_1771,N_1660,N_1692);
or U1772 (N_1772,N_1708,N_1706);
and U1773 (N_1773,N_1689,N_1697);
nor U1774 (N_1774,N_1677,N_1706);
nand U1775 (N_1775,N_1652,N_1664);
nand U1776 (N_1776,N_1695,N_1653);
nor U1777 (N_1777,N_1687,N_1679);
nor U1778 (N_1778,N_1699,N_1663);
and U1779 (N_1779,N_1671,N_1701);
or U1780 (N_1780,N_1722,N_1719);
and U1781 (N_1781,N_1680,N_1678);
or U1782 (N_1782,N_1686,N_1672);
and U1783 (N_1783,N_1651,N_1722);
or U1784 (N_1784,N_1721,N_1662);
nor U1785 (N_1785,N_1655,N_1704);
nand U1786 (N_1786,N_1702,N_1655);
nor U1787 (N_1787,N_1724,N_1699);
and U1788 (N_1788,N_1704,N_1687);
or U1789 (N_1789,N_1670,N_1711);
and U1790 (N_1790,N_1696,N_1662);
and U1791 (N_1791,N_1660,N_1705);
nand U1792 (N_1792,N_1720,N_1666);
nand U1793 (N_1793,N_1700,N_1680);
nand U1794 (N_1794,N_1666,N_1679);
and U1795 (N_1795,N_1684,N_1710);
nor U1796 (N_1796,N_1687,N_1673);
or U1797 (N_1797,N_1714,N_1703);
nor U1798 (N_1798,N_1673,N_1688);
and U1799 (N_1799,N_1650,N_1721);
or U1800 (N_1800,N_1743,N_1732);
or U1801 (N_1801,N_1791,N_1786);
nor U1802 (N_1802,N_1756,N_1751);
nand U1803 (N_1803,N_1747,N_1725);
and U1804 (N_1804,N_1745,N_1788);
nor U1805 (N_1805,N_1738,N_1730);
nand U1806 (N_1806,N_1768,N_1727);
nor U1807 (N_1807,N_1729,N_1737);
xnor U1808 (N_1808,N_1749,N_1746);
and U1809 (N_1809,N_1752,N_1757);
nor U1810 (N_1810,N_1779,N_1799);
and U1811 (N_1811,N_1796,N_1754);
nor U1812 (N_1812,N_1778,N_1735);
nor U1813 (N_1813,N_1731,N_1794);
nor U1814 (N_1814,N_1793,N_1726);
nor U1815 (N_1815,N_1797,N_1758);
or U1816 (N_1816,N_1741,N_1772);
and U1817 (N_1817,N_1770,N_1789);
and U1818 (N_1818,N_1748,N_1781);
and U1819 (N_1819,N_1785,N_1766);
or U1820 (N_1820,N_1763,N_1742);
nor U1821 (N_1821,N_1771,N_1753);
or U1822 (N_1822,N_1774,N_1769);
nor U1823 (N_1823,N_1744,N_1777);
and U1824 (N_1824,N_1783,N_1784);
nor U1825 (N_1825,N_1790,N_1787);
nor U1826 (N_1826,N_1759,N_1736);
and U1827 (N_1827,N_1728,N_1762);
or U1828 (N_1828,N_1750,N_1767);
nor U1829 (N_1829,N_1740,N_1733);
nand U1830 (N_1830,N_1764,N_1773);
and U1831 (N_1831,N_1798,N_1782);
or U1832 (N_1832,N_1755,N_1776);
and U1833 (N_1833,N_1761,N_1775);
nand U1834 (N_1834,N_1760,N_1734);
nor U1835 (N_1835,N_1739,N_1792);
nor U1836 (N_1836,N_1780,N_1765);
and U1837 (N_1837,N_1795,N_1731);
and U1838 (N_1838,N_1741,N_1780);
nand U1839 (N_1839,N_1745,N_1757);
and U1840 (N_1840,N_1763,N_1773);
and U1841 (N_1841,N_1752,N_1749);
nor U1842 (N_1842,N_1795,N_1772);
or U1843 (N_1843,N_1777,N_1748);
nor U1844 (N_1844,N_1798,N_1763);
nand U1845 (N_1845,N_1772,N_1763);
nor U1846 (N_1846,N_1735,N_1749);
or U1847 (N_1847,N_1775,N_1757);
xnor U1848 (N_1848,N_1775,N_1763);
and U1849 (N_1849,N_1762,N_1742);
nor U1850 (N_1850,N_1785,N_1757);
and U1851 (N_1851,N_1738,N_1755);
and U1852 (N_1852,N_1739,N_1756);
or U1853 (N_1853,N_1781,N_1790);
nand U1854 (N_1854,N_1730,N_1753);
or U1855 (N_1855,N_1739,N_1766);
and U1856 (N_1856,N_1778,N_1757);
nand U1857 (N_1857,N_1777,N_1784);
and U1858 (N_1858,N_1747,N_1761);
or U1859 (N_1859,N_1779,N_1752);
nor U1860 (N_1860,N_1782,N_1796);
and U1861 (N_1861,N_1737,N_1751);
or U1862 (N_1862,N_1771,N_1734);
and U1863 (N_1863,N_1777,N_1786);
or U1864 (N_1864,N_1736,N_1791);
nor U1865 (N_1865,N_1733,N_1746);
nor U1866 (N_1866,N_1767,N_1765);
and U1867 (N_1867,N_1796,N_1780);
nor U1868 (N_1868,N_1752,N_1799);
or U1869 (N_1869,N_1756,N_1730);
nor U1870 (N_1870,N_1759,N_1728);
nand U1871 (N_1871,N_1755,N_1748);
nand U1872 (N_1872,N_1794,N_1747);
or U1873 (N_1873,N_1740,N_1760);
nand U1874 (N_1874,N_1753,N_1770);
nand U1875 (N_1875,N_1815,N_1857);
nand U1876 (N_1876,N_1824,N_1816);
and U1877 (N_1877,N_1828,N_1805);
or U1878 (N_1878,N_1870,N_1819);
nor U1879 (N_1879,N_1846,N_1839);
or U1880 (N_1880,N_1849,N_1861);
nor U1881 (N_1881,N_1813,N_1837);
nor U1882 (N_1882,N_1860,N_1872);
nor U1883 (N_1883,N_1865,N_1871);
nand U1884 (N_1884,N_1818,N_1866);
and U1885 (N_1885,N_1801,N_1842);
nor U1886 (N_1886,N_1800,N_1829);
or U1887 (N_1887,N_1855,N_1845);
nand U1888 (N_1888,N_1862,N_1804);
nand U1889 (N_1889,N_1832,N_1847);
nor U1890 (N_1890,N_1843,N_1874);
nor U1891 (N_1891,N_1841,N_1833);
nor U1892 (N_1892,N_1812,N_1811);
or U1893 (N_1893,N_1869,N_1807);
nor U1894 (N_1894,N_1859,N_1814);
or U1895 (N_1895,N_1873,N_1858);
xnor U1896 (N_1896,N_1825,N_1836);
and U1897 (N_1897,N_1822,N_1827);
xor U1898 (N_1898,N_1854,N_1867);
nand U1899 (N_1899,N_1809,N_1852);
and U1900 (N_1900,N_1823,N_1806);
and U1901 (N_1901,N_1844,N_1856);
or U1902 (N_1902,N_1863,N_1810);
nor U1903 (N_1903,N_1830,N_1808);
or U1904 (N_1904,N_1831,N_1802);
nand U1905 (N_1905,N_1834,N_1803);
nand U1906 (N_1906,N_1838,N_1864);
and U1907 (N_1907,N_1853,N_1835);
or U1908 (N_1908,N_1820,N_1851);
nor U1909 (N_1909,N_1850,N_1868);
nand U1910 (N_1910,N_1848,N_1821);
nand U1911 (N_1911,N_1826,N_1817);
and U1912 (N_1912,N_1840,N_1820);
and U1913 (N_1913,N_1819,N_1844);
nand U1914 (N_1914,N_1813,N_1809);
nor U1915 (N_1915,N_1873,N_1841);
nand U1916 (N_1916,N_1828,N_1868);
nor U1917 (N_1917,N_1803,N_1845);
nand U1918 (N_1918,N_1843,N_1822);
nor U1919 (N_1919,N_1842,N_1822);
nor U1920 (N_1920,N_1841,N_1807);
or U1921 (N_1921,N_1841,N_1824);
or U1922 (N_1922,N_1811,N_1837);
nor U1923 (N_1923,N_1822,N_1848);
or U1924 (N_1924,N_1830,N_1869);
nand U1925 (N_1925,N_1843,N_1802);
nor U1926 (N_1926,N_1842,N_1841);
or U1927 (N_1927,N_1807,N_1856);
or U1928 (N_1928,N_1832,N_1822);
xnor U1929 (N_1929,N_1805,N_1863);
or U1930 (N_1930,N_1819,N_1855);
nor U1931 (N_1931,N_1801,N_1854);
and U1932 (N_1932,N_1821,N_1862);
and U1933 (N_1933,N_1818,N_1874);
and U1934 (N_1934,N_1836,N_1814);
nor U1935 (N_1935,N_1834,N_1861);
nor U1936 (N_1936,N_1804,N_1859);
nand U1937 (N_1937,N_1855,N_1844);
nand U1938 (N_1938,N_1829,N_1812);
nor U1939 (N_1939,N_1827,N_1865);
and U1940 (N_1940,N_1855,N_1812);
and U1941 (N_1941,N_1834,N_1806);
and U1942 (N_1942,N_1830,N_1820);
or U1943 (N_1943,N_1844,N_1832);
nand U1944 (N_1944,N_1852,N_1854);
and U1945 (N_1945,N_1834,N_1811);
nand U1946 (N_1946,N_1800,N_1824);
nand U1947 (N_1947,N_1844,N_1822);
nand U1948 (N_1948,N_1802,N_1846);
nor U1949 (N_1949,N_1816,N_1821);
nand U1950 (N_1950,N_1892,N_1928);
and U1951 (N_1951,N_1916,N_1885);
and U1952 (N_1952,N_1935,N_1888);
nand U1953 (N_1953,N_1907,N_1921);
or U1954 (N_1954,N_1941,N_1936);
or U1955 (N_1955,N_1917,N_1881);
and U1956 (N_1956,N_1937,N_1879);
nand U1957 (N_1957,N_1882,N_1939);
nor U1958 (N_1958,N_1895,N_1923);
nand U1959 (N_1959,N_1887,N_1945);
nand U1960 (N_1960,N_1927,N_1932);
and U1961 (N_1961,N_1883,N_1925);
nor U1962 (N_1962,N_1946,N_1899);
or U1963 (N_1963,N_1908,N_1912);
and U1964 (N_1964,N_1944,N_1929);
nor U1965 (N_1965,N_1889,N_1884);
nand U1966 (N_1966,N_1918,N_1905);
or U1967 (N_1967,N_1911,N_1901);
and U1968 (N_1968,N_1893,N_1934);
nor U1969 (N_1969,N_1896,N_1909);
nand U1970 (N_1970,N_1915,N_1890);
or U1971 (N_1971,N_1875,N_1914);
nand U1972 (N_1972,N_1940,N_1933);
nand U1973 (N_1973,N_1910,N_1880);
nand U1974 (N_1974,N_1920,N_1949);
nor U1975 (N_1975,N_1886,N_1926);
nand U1976 (N_1976,N_1938,N_1924);
and U1977 (N_1977,N_1913,N_1898);
nor U1978 (N_1978,N_1943,N_1897);
and U1979 (N_1979,N_1894,N_1891);
nand U1980 (N_1980,N_1931,N_1900);
nand U1981 (N_1981,N_1948,N_1919);
nor U1982 (N_1982,N_1902,N_1877);
nor U1983 (N_1983,N_1878,N_1903);
nand U1984 (N_1984,N_1922,N_1942);
or U1985 (N_1985,N_1906,N_1947);
xor U1986 (N_1986,N_1876,N_1930);
nor U1987 (N_1987,N_1904,N_1885);
and U1988 (N_1988,N_1943,N_1892);
xnor U1989 (N_1989,N_1918,N_1937);
or U1990 (N_1990,N_1933,N_1892);
nand U1991 (N_1991,N_1928,N_1936);
nand U1992 (N_1992,N_1937,N_1911);
nor U1993 (N_1993,N_1882,N_1908);
nor U1994 (N_1994,N_1943,N_1949);
nor U1995 (N_1995,N_1933,N_1908);
nand U1996 (N_1996,N_1882,N_1933);
nor U1997 (N_1997,N_1892,N_1900);
or U1998 (N_1998,N_1918,N_1876);
and U1999 (N_1999,N_1928,N_1942);
xor U2000 (N_2000,N_1901,N_1943);
nand U2001 (N_2001,N_1883,N_1900);
nand U2002 (N_2002,N_1885,N_1897);
nor U2003 (N_2003,N_1932,N_1889);
nand U2004 (N_2004,N_1884,N_1913);
nor U2005 (N_2005,N_1900,N_1901);
nor U2006 (N_2006,N_1892,N_1912);
and U2007 (N_2007,N_1892,N_1895);
nand U2008 (N_2008,N_1905,N_1900);
or U2009 (N_2009,N_1943,N_1944);
or U2010 (N_2010,N_1899,N_1942);
or U2011 (N_2011,N_1908,N_1949);
nor U2012 (N_2012,N_1928,N_1890);
nand U2013 (N_2013,N_1890,N_1917);
nand U2014 (N_2014,N_1903,N_1945);
nand U2015 (N_2015,N_1882,N_1941);
nor U2016 (N_2016,N_1881,N_1912);
nor U2017 (N_2017,N_1886,N_1876);
nor U2018 (N_2018,N_1938,N_1886);
and U2019 (N_2019,N_1876,N_1927);
or U2020 (N_2020,N_1921,N_1949);
nor U2021 (N_2021,N_1932,N_1894);
xnor U2022 (N_2022,N_1940,N_1902);
or U2023 (N_2023,N_1883,N_1879);
nor U2024 (N_2024,N_1909,N_1884);
or U2025 (N_2025,N_1953,N_1959);
or U2026 (N_2026,N_2006,N_2002);
nor U2027 (N_2027,N_2010,N_1966);
nor U2028 (N_2028,N_2024,N_1977);
nor U2029 (N_2029,N_1956,N_2012);
nand U2030 (N_2030,N_2021,N_1983);
xor U2031 (N_2031,N_1994,N_1967);
and U2032 (N_2032,N_2004,N_1961);
or U2033 (N_2033,N_2007,N_1989);
nor U2034 (N_2034,N_2018,N_2023);
and U2035 (N_2035,N_2016,N_1981);
or U2036 (N_2036,N_1978,N_1995);
nand U2037 (N_2037,N_1960,N_1958);
and U2038 (N_2038,N_2011,N_2009);
nor U2039 (N_2039,N_1997,N_1999);
xor U2040 (N_2040,N_1965,N_1950);
xnor U2041 (N_2041,N_1957,N_1954);
nor U2042 (N_2042,N_2008,N_1988);
nor U2043 (N_2043,N_1971,N_2014);
and U2044 (N_2044,N_1973,N_1968);
or U2045 (N_2045,N_2020,N_1951);
and U2046 (N_2046,N_1987,N_1979);
or U2047 (N_2047,N_2003,N_1972);
nor U2048 (N_2048,N_1976,N_1992);
and U2049 (N_2049,N_2005,N_2001);
and U2050 (N_2050,N_1952,N_1984);
nand U2051 (N_2051,N_1964,N_1996);
nand U2052 (N_2052,N_1991,N_1980);
or U2053 (N_2053,N_2019,N_2000);
and U2054 (N_2054,N_2022,N_2017);
and U2055 (N_2055,N_1975,N_1969);
and U2056 (N_2056,N_1962,N_2013);
or U2057 (N_2057,N_1993,N_1970);
or U2058 (N_2058,N_1955,N_1990);
nor U2059 (N_2059,N_1974,N_2015);
nor U2060 (N_2060,N_1982,N_1986);
or U2061 (N_2061,N_1963,N_1985);
nor U2062 (N_2062,N_1998,N_1956);
nor U2063 (N_2063,N_1975,N_2010);
or U2064 (N_2064,N_2009,N_1975);
or U2065 (N_2065,N_1990,N_1976);
or U2066 (N_2066,N_1976,N_2022);
or U2067 (N_2067,N_2019,N_2002);
nand U2068 (N_2068,N_1953,N_1972);
xor U2069 (N_2069,N_2008,N_1979);
nand U2070 (N_2070,N_1957,N_1979);
nand U2071 (N_2071,N_1997,N_1958);
nand U2072 (N_2072,N_1957,N_1999);
nand U2073 (N_2073,N_1970,N_1965);
and U2074 (N_2074,N_1987,N_2023);
or U2075 (N_2075,N_2017,N_1991);
and U2076 (N_2076,N_2018,N_1973);
and U2077 (N_2077,N_2020,N_2016);
nand U2078 (N_2078,N_1974,N_1972);
or U2079 (N_2079,N_2013,N_1956);
or U2080 (N_2080,N_1969,N_2003);
and U2081 (N_2081,N_1955,N_1956);
nand U2082 (N_2082,N_1999,N_1996);
nand U2083 (N_2083,N_1980,N_2009);
nor U2084 (N_2084,N_1984,N_2022);
or U2085 (N_2085,N_1966,N_1953);
xnor U2086 (N_2086,N_1982,N_2018);
xnor U2087 (N_2087,N_1989,N_1974);
or U2088 (N_2088,N_2015,N_2011);
or U2089 (N_2089,N_2011,N_2013);
nand U2090 (N_2090,N_1985,N_1986);
or U2091 (N_2091,N_2000,N_1992);
or U2092 (N_2092,N_1957,N_1992);
and U2093 (N_2093,N_1972,N_1969);
xor U2094 (N_2094,N_2006,N_1997);
nand U2095 (N_2095,N_1984,N_2012);
and U2096 (N_2096,N_1990,N_1961);
or U2097 (N_2097,N_1965,N_1967);
and U2098 (N_2098,N_1976,N_1977);
or U2099 (N_2099,N_1950,N_2018);
or U2100 (N_2100,N_2043,N_2047);
and U2101 (N_2101,N_2053,N_2051);
nand U2102 (N_2102,N_2063,N_2086);
and U2103 (N_2103,N_2026,N_2083);
or U2104 (N_2104,N_2084,N_2027);
nor U2105 (N_2105,N_2092,N_2095);
nor U2106 (N_2106,N_2078,N_2034);
nand U2107 (N_2107,N_2025,N_2069);
nand U2108 (N_2108,N_2073,N_2074);
or U2109 (N_2109,N_2055,N_2079);
nor U2110 (N_2110,N_2097,N_2090);
nand U2111 (N_2111,N_2061,N_2099);
and U2112 (N_2112,N_2065,N_2085);
and U2113 (N_2113,N_2075,N_2089);
or U2114 (N_2114,N_2030,N_2057);
and U2115 (N_2115,N_2036,N_2035);
or U2116 (N_2116,N_2062,N_2088);
nor U2117 (N_2117,N_2041,N_2042);
or U2118 (N_2118,N_2052,N_2081);
and U2119 (N_2119,N_2044,N_2072);
nand U2120 (N_2120,N_2029,N_2048);
nand U2121 (N_2121,N_2039,N_2059);
and U2122 (N_2122,N_2049,N_2093);
or U2123 (N_2123,N_2087,N_2066);
and U2124 (N_2124,N_2050,N_2094);
and U2125 (N_2125,N_2046,N_2091);
nand U2126 (N_2126,N_2033,N_2038);
and U2127 (N_2127,N_2032,N_2058);
nor U2128 (N_2128,N_2064,N_2070);
and U2129 (N_2129,N_2031,N_2071);
nor U2130 (N_2130,N_2060,N_2082);
nor U2131 (N_2131,N_2028,N_2054);
nor U2132 (N_2132,N_2056,N_2076);
or U2133 (N_2133,N_2068,N_2098);
nor U2134 (N_2134,N_2045,N_2040);
nor U2135 (N_2135,N_2096,N_2080);
nor U2136 (N_2136,N_2067,N_2037);
nand U2137 (N_2137,N_2077,N_2037);
or U2138 (N_2138,N_2043,N_2087);
or U2139 (N_2139,N_2055,N_2085);
nand U2140 (N_2140,N_2042,N_2044);
nand U2141 (N_2141,N_2080,N_2028);
or U2142 (N_2142,N_2069,N_2071);
nor U2143 (N_2143,N_2093,N_2080);
or U2144 (N_2144,N_2071,N_2027);
or U2145 (N_2145,N_2066,N_2094);
nor U2146 (N_2146,N_2026,N_2042);
nor U2147 (N_2147,N_2060,N_2033);
or U2148 (N_2148,N_2049,N_2081);
nor U2149 (N_2149,N_2087,N_2051);
and U2150 (N_2150,N_2077,N_2038);
nor U2151 (N_2151,N_2061,N_2058);
nor U2152 (N_2152,N_2088,N_2077);
xnor U2153 (N_2153,N_2050,N_2038);
and U2154 (N_2154,N_2045,N_2084);
and U2155 (N_2155,N_2033,N_2077);
nand U2156 (N_2156,N_2070,N_2097);
nor U2157 (N_2157,N_2052,N_2034);
nand U2158 (N_2158,N_2030,N_2090);
xor U2159 (N_2159,N_2038,N_2034);
nor U2160 (N_2160,N_2089,N_2031);
or U2161 (N_2161,N_2069,N_2077);
nor U2162 (N_2162,N_2039,N_2074);
nand U2163 (N_2163,N_2045,N_2044);
and U2164 (N_2164,N_2079,N_2068);
nor U2165 (N_2165,N_2050,N_2078);
nor U2166 (N_2166,N_2056,N_2091);
and U2167 (N_2167,N_2062,N_2028);
nand U2168 (N_2168,N_2095,N_2072);
or U2169 (N_2169,N_2033,N_2037);
nand U2170 (N_2170,N_2097,N_2060);
or U2171 (N_2171,N_2060,N_2087);
nor U2172 (N_2172,N_2062,N_2047);
nand U2173 (N_2173,N_2045,N_2037);
nor U2174 (N_2174,N_2027,N_2079);
nor U2175 (N_2175,N_2124,N_2131);
and U2176 (N_2176,N_2101,N_2119);
and U2177 (N_2177,N_2142,N_2122);
nor U2178 (N_2178,N_2144,N_2164);
or U2179 (N_2179,N_2155,N_2126);
nor U2180 (N_2180,N_2149,N_2139);
and U2181 (N_2181,N_2115,N_2129);
nor U2182 (N_2182,N_2100,N_2153);
nand U2183 (N_2183,N_2109,N_2163);
nor U2184 (N_2184,N_2111,N_2116);
xnor U2185 (N_2185,N_2156,N_2125);
or U2186 (N_2186,N_2140,N_2166);
nand U2187 (N_2187,N_2154,N_2143);
or U2188 (N_2188,N_2169,N_2132);
and U2189 (N_2189,N_2104,N_2145);
or U2190 (N_2190,N_2150,N_2123);
and U2191 (N_2191,N_2137,N_2121);
nor U2192 (N_2192,N_2141,N_2117);
and U2193 (N_2193,N_2128,N_2162);
or U2194 (N_2194,N_2135,N_2161);
or U2195 (N_2195,N_2106,N_2105);
nor U2196 (N_2196,N_2170,N_2102);
or U2197 (N_2197,N_2173,N_2147);
or U2198 (N_2198,N_2103,N_2152);
nand U2199 (N_2199,N_2148,N_2172);
nor U2200 (N_2200,N_2171,N_2114);
xnor U2201 (N_2201,N_2108,N_2146);
and U2202 (N_2202,N_2157,N_2127);
and U2203 (N_2203,N_2160,N_2138);
nor U2204 (N_2204,N_2167,N_2159);
or U2205 (N_2205,N_2133,N_2158);
nand U2206 (N_2206,N_2110,N_2118);
or U2207 (N_2207,N_2151,N_2165);
and U2208 (N_2208,N_2130,N_2120);
or U2209 (N_2209,N_2168,N_2174);
or U2210 (N_2210,N_2113,N_2136);
or U2211 (N_2211,N_2134,N_2112);
nor U2212 (N_2212,N_2107,N_2129);
and U2213 (N_2213,N_2127,N_2147);
and U2214 (N_2214,N_2136,N_2120);
or U2215 (N_2215,N_2151,N_2164);
and U2216 (N_2216,N_2119,N_2169);
nor U2217 (N_2217,N_2129,N_2116);
and U2218 (N_2218,N_2139,N_2124);
or U2219 (N_2219,N_2112,N_2123);
and U2220 (N_2220,N_2160,N_2107);
nor U2221 (N_2221,N_2135,N_2111);
or U2222 (N_2222,N_2172,N_2153);
nand U2223 (N_2223,N_2107,N_2115);
nand U2224 (N_2224,N_2108,N_2143);
nor U2225 (N_2225,N_2152,N_2133);
or U2226 (N_2226,N_2146,N_2117);
and U2227 (N_2227,N_2158,N_2160);
nand U2228 (N_2228,N_2151,N_2146);
and U2229 (N_2229,N_2141,N_2119);
and U2230 (N_2230,N_2172,N_2123);
nand U2231 (N_2231,N_2130,N_2127);
nand U2232 (N_2232,N_2144,N_2160);
xor U2233 (N_2233,N_2119,N_2111);
or U2234 (N_2234,N_2100,N_2130);
xor U2235 (N_2235,N_2125,N_2164);
nand U2236 (N_2236,N_2117,N_2125);
and U2237 (N_2237,N_2134,N_2133);
and U2238 (N_2238,N_2152,N_2154);
and U2239 (N_2239,N_2171,N_2107);
and U2240 (N_2240,N_2111,N_2151);
or U2241 (N_2241,N_2150,N_2116);
nor U2242 (N_2242,N_2112,N_2111);
nor U2243 (N_2243,N_2162,N_2151);
and U2244 (N_2244,N_2134,N_2113);
nand U2245 (N_2245,N_2111,N_2136);
nor U2246 (N_2246,N_2104,N_2131);
and U2247 (N_2247,N_2135,N_2145);
nand U2248 (N_2248,N_2136,N_2164);
and U2249 (N_2249,N_2167,N_2145);
or U2250 (N_2250,N_2211,N_2178);
or U2251 (N_2251,N_2223,N_2205);
nand U2252 (N_2252,N_2196,N_2214);
nor U2253 (N_2253,N_2182,N_2228);
or U2254 (N_2254,N_2232,N_2230);
and U2255 (N_2255,N_2179,N_2225);
nand U2256 (N_2256,N_2247,N_2197);
nand U2257 (N_2257,N_2212,N_2209);
nand U2258 (N_2258,N_2176,N_2222);
nand U2259 (N_2259,N_2183,N_2215);
and U2260 (N_2260,N_2233,N_2201);
xor U2261 (N_2261,N_2243,N_2193);
nor U2262 (N_2262,N_2192,N_2231);
nor U2263 (N_2263,N_2188,N_2219);
xnor U2264 (N_2264,N_2202,N_2185);
and U2265 (N_2265,N_2246,N_2175);
and U2266 (N_2266,N_2220,N_2206);
and U2267 (N_2267,N_2218,N_2236);
and U2268 (N_2268,N_2189,N_2217);
nor U2269 (N_2269,N_2242,N_2234);
and U2270 (N_2270,N_2241,N_2187);
nand U2271 (N_2271,N_2191,N_2177);
nand U2272 (N_2272,N_2203,N_2208);
or U2273 (N_2273,N_2181,N_2207);
xnor U2274 (N_2274,N_2210,N_2184);
or U2275 (N_2275,N_2180,N_2238);
or U2276 (N_2276,N_2245,N_2200);
and U2277 (N_2277,N_2199,N_2186);
or U2278 (N_2278,N_2213,N_2240);
nand U2279 (N_2279,N_2226,N_2229);
nand U2280 (N_2280,N_2194,N_2235);
and U2281 (N_2281,N_2244,N_2221);
nor U2282 (N_2282,N_2239,N_2248);
or U2283 (N_2283,N_2195,N_2237);
nor U2284 (N_2284,N_2204,N_2190);
nand U2285 (N_2285,N_2227,N_2216);
nand U2286 (N_2286,N_2198,N_2249);
nand U2287 (N_2287,N_2224,N_2246);
xnor U2288 (N_2288,N_2237,N_2184);
nor U2289 (N_2289,N_2243,N_2192);
or U2290 (N_2290,N_2233,N_2208);
and U2291 (N_2291,N_2239,N_2180);
nand U2292 (N_2292,N_2241,N_2178);
nand U2293 (N_2293,N_2203,N_2228);
nor U2294 (N_2294,N_2242,N_2248);
nand U2295 (N_2295,N_2195,N_2225);
xor U2296 (N_2296,N_2221,N_2240);
nand U2297 (N_2297,N_2219,N_2182);
and U2298 (N_2298,N_2241,N_2227);
nor U2299 (N_2299,N_2213,N_2200);
or U2300 (N_2300,N_2215,N_2191);
nor U2301 (N_2301,N_2198,N_2197);
or U2302 (N_2302,N_2226,N_2244);
nand U2303 (N_2303,N_2177,N_2235);
nor U2304 (N_2304,N_2227,N_2226);
and U2305 (N_2305,N_2228,N_2184);
and U2306 (N_2306,N_2204,N_2211);
or U2307 (N_2307,N_2215,N_2248);
nor U2308 (N_2308,N_2248,N_2202);
nand U2309 (N_2309,N_2213,N_2220);
nor U2310 (N_2310,N_2218,N_2237);
or U2311 (N_2311,N_2205,N_2182);
nand U2312 (N_2312,N_2206,N_2179);
xnor U2313 (N_2313,N_2209,N_2178);
nor U2314 (N_2314,N_2197,N_2202);
or U2315 (N_2315,N_2182,N_2226);
or U2316 (N_2316,N_2209,N_2191);
nand U2317 (N_2317,N_2190,N_2188);
and U2318 (N_2318,N_2188,N_2239);
or U2319 (N_2319,N_2191,N_2214);
or U2320 (N_2320,N_2181,N_2205);
or U2321 (N_2321,N_2182,N_2187);
nand U2322 (N_2322,N_2201,N_2202);
nand U2323 (N_2323,N_2176,N_2241);
nand U2324 (N_2324,N_2218,N_2195);
nor U2325 (N_2325,N_2299,N_2251);
nand U2326 (N_2326,N_2271,N_2264);
or U2327 (N_2327,N_2272,N_2318);
nor U2328 (N_2328,N_2316,N_2295);
nand U2329 (N_2329,N_2265,N_2268);
and U2330 (N_2330,N_2273,N_2288);
and U2331 (N_2331,N_2308,N_2303);
nand U2332 (N_2332,N_2291,N_2312);
nand U2333 (N_2333,N_2257,N_2292);
or U2334 (N_2334,N_2262,N_2275);
or U2335 (N_2335,N_2321,N_2267);
or U2336 (N_2336,N_2261,N_2269);
or U2337 (N_2337,N_2277,N_2315);
nor U2338 (N_2338,N_2278,N_2280);
or U2339 (N_2339,N_2270,N_2281);
or U2340 (N_2340,N_2282,N_2279);
nor U2341 (N_2341,N_2255,N_2258);
xnor U2342 (N_2342,N_2309,N_2300);
nor U2343 (N_2343,N_2302,N_2256);
or U2344 (N_2344,N_2293,N_2322);
nand U2345 (N_2345,N_2298,N_2290);
or U2346 (N_2346,N_2296,N_2252);
nand U2347 (N_2347,N_2297,N_2306);
nand U2348 (N_2348,N_2285,N_2274);
nor U2349 (N_2349,N_2254,N_2317);
nand U2350 (N_2350,N_2287,N_2250);
nor U2351 (N_2351,N_2304,N_2289);
or U2352 (N_2352,N_2286,N_2307);
nor U2353 (N_2353,N_2320,N_2301);
and U2354 (N_2354,N_2263,N_2323);
and U2355 (N_2355,N_2266,N_2314);
xnor U2356 (N_2356,N_2253,N_2324);
or U2357 (N_2357,N_2310,N_2276);
nor U2358 (N_2358,N_2305,N_2319);
or U2359 (N_2359,N_2313,N_2284);
nor U2360 (N_2360,N_2294,N_2283);
nor U2361 (N_2361,N_2259,N_2260);
xnor U2362 (N_2362,N_2311,N_2322);
nand U2363 (N_2363,N_2286,N_2255);
nor U2364 (N_2364,N_2322,N_2292);
and U2365 (N_2365,N_2302,N_2280);
and U2366 (N_2366,N_2296,N_2253);
or U2367 (N_2367,N_2280,N_2272);
or U2368 (N_2368,N_2260,N_2314);
xor U2369 (N_2369,N_2305,N_2299);
and U2370 (N_2370,N_2302,N_2266);
or U2371 (N_2371,N_2320,N_2252);
nor U2372 (N_2372,N_2278,N_2289);
and U2373 (N_2373,N_2294,N_2298);
nor U2374 (N_2374,N_2306,N_2293);
or U2375 (N_2375,N_2274,N_2289);
or U2376 (N_2376,N_2251,N_2268);
nor U2377 (N_2377,N_2299,N_2297);
nand U2378 (N_2378,N_2283,N_2274);
or U2379 (N_2379,N_2264,N_2270);
nor U2380 (N_2380,N_2284,N_2319);
nand U2381 (N_2381,N_2298,N_2251);
or U2382 (N_2382,N_2250,N_2322);
nor U2383 (N_2383,N_2258,N_2305);
xor U2384 (N_2384,N_2284,N_2308);
nand U2385 (N_2385,N_2274,N_2271);
nor U2386 (N_2386,N_2269,N_2313);
nor U2387 (N_2387,N_2304,N_2277);
nand U2388 (N_2388,N_2298,N_2300);
and U2389 (N_2389,N_2304,N_2254);
or U2390 (N_2390,N_2262,N_2305);
or U2391 (N_2391,N_2278,N_2317);
and U2392 (N_2392,N_2285,N_2298);
or U2393 (N_2393,N_2310,N_2320);
or U2394 (N_2394,N_2264,N_2300);
and U2395 (N_2395,N_2251,N_2285);
and U2396 (N_2396,N_2293,N_2268);
nand U2397 (N_2397,N_2301,N_2310);
and U2398 (N_2398,N_2304,N_2282);
nand U2399 (N_2399,N_2257,N_2255);
or U2400 (N_2400,N_2334,N_2388);
nand U2401 (N_2401,N_2333,N_2352);
nor U2402 (N_2402,N_2355,N_2339);
or U2403 (N_2403,N_2383,N_2330);
nand U2404 (N_2404,N_2349,N_2326);
and U2405 (N_2405,N_2369,N_2373);
and U2406 (N_2406,N_2393,N_2399);
and U2407 (N_2407,N_2382,N_2378);
or U2408 (N_2408,N_2395,N_2377);
nand U2409 (N_2409,N_2357,N_2364);
nor U2410 (N_2410,N_2375,N_2380);
nor U2411 (N_2411,N_2372,N_2345);
or U2412 (N_2412,N_2394,N_2386);
nor U2413 (N_2413,N_2387,N_2391);
nor U2414 (N_2414,N_2389,N_2351);
nor U2415 (N_2415,N_2379,N_2359);
or U2416 (N_2416,N_2366,N_2350);
nand U2417 (N_2417,N_2325,N_2398);
or U2418 (N_2418,N_2341,N_2368);
or U2419 (N_2419,N_2353,N_2367);
and U2420 (N_2420,N_2329,N_2384);
or U2421 (N_2421,N_2332,N_2385);
xor U2422 (N_2422,N_2336,N_2363);
or U2423 (N_2423,N_2348,N_2371);
nand U2424 (N_2424,N_2338,N_2356);
nor U2425 (N_2425,N_2354,N_2370);
nor U2426 (N_2426,N_2392,N_2327);
and U2427 (N_2427,N_2397,N_2360);
nor U2428 (N_2428,N_2343,N_2358);
and U2429 (N_2429,N_2337,N_2346);
and U2430 (N_2430,N_2344,N_2381);
and U2431 (N_2431,N_2331,N_2374);
or U2432 (N_2432,N_2335,N_2362);
and U2433 (N_2433,N_2365,N_2328);
nor U2434 (N_2434,N_2340,N_2396);
xnor U2435 (N_2435,N_2361,N_2347);
nand U2436 (N_2436,N_2342,N_2390);
nand U2437 (N_2437,N_2376,N_2330);
nor U2438 (N_2438,N_2384,N_2341);
and U2439 (N_2439,N_2336,N_2373);
nor U2440 (N_2440,N_2353,N_2383);
or U2441 (N_2441,N_2344,N_2375);
and U2442 (N_2442,N_2359,N_2337);
nand U2443 (N_2443,N_2330,N_2333);
and U2444 (N_2444,N_2365,N_2325);
nor U2445 (N_2445,N_2332,N_2374);
and U2446 (N_2446,N_2375,N_2355);
or U2447 (N_2447,N_2360,N_2330);
and U2448 (N_2448,N_2340,N_2334);
nor U2449 (N_2449,N_2387,N_2379);
xor U2450 (N_2450,N_2385,N_2399);
nor U2451 (N_2451,N_2347,N_2383);
and U2452 (N_2452,N_2341,N_2357);
nand U2453 (N_2453,N_2325,N_2332);
nand U2454 (N_2454,N_2382,N_2384);
nor U2455 (N_2455,N_2395,N_2338);
nor U2456 (N_2456,N_2349,N_2371);
nor U2457 (N_2457,N_2339,N_2368);
or U2458 (N_2458,N_2364,N_2393);
nand U2459 (N_2459,N_2396,N_2390);
nor U2460 (N_2460,N_2343,N_2327);
nor U2461 (N_2461,N_2366,N_2395);
nor U2462 (N_2462,N_2343,N_2373);
and U2463 (N_2463,N_2364,N_2384);
nand U2464 (N_2464,N_2375,N_2399);
nand U2465 (N_2465,N_2369,N_2389);
or U2466 (N_2466,N_2373,N_2348);
nand U2467 (N_2467,N_2372,N_2342);
nor U2468 (N_2468,N_2333,N_2396);
nand U2469 (N_2469,N_2367,N_2398);
or U2470 (N_2470,N_2358,N_2372);
nand U2471 (N_2471,N_2355,N_2347);
or U2472 (N_2472,N_2370,N_2364);
nor U2473 (N_2473,N_2343,N_2353);
nand U2474 (N_2474,N_2352,N_2368);
or U2475 (N_2475,N_2459,N_2464);
nor U2476 (N_2476,N_2452,N_2432);
or U2477 (N_2477,N_2405,N_2440);
nand U2478 (N_2478,N_2402,N_2437);
and U2479 (N_2479,N_2429,N_2434);
nand U2480 (N_2480,N_2466,N_2410);
and U2481 (N_2481,N_2424,N_2414);
nor U2482 (N_2482,N_2474,N_2461);
and U2483 (N_2483,N_2430,N_2409);
and U2484 (N_2484,N_2448,N_2454);
and U2485 (N_2485,N_2455,N_2403);
nor U2486 (N_2486,N_2427,N_2425);
nor U2487 (N_2487,N_2400,N_2444);
and U2488 (N_2488,N_2413,N_2447);
nand U2489 (N_2489,N_2438,N_2418);
xnor U2490 (N_2490,N_2453,N_2433);
nand U2491 (N_2491,N_2422,N_2407);
or U2492 (N_2492,N_2406,N_2401);
nand U2493 (N_2493,N_2416,N_2408);
nor U2494 (N_2494,N_2421,N_2473);
nand U2495 (N_2495,N_2456,N_2445);
nor U2496 (N_2496,N_2436,N_2441);
nand U2497 (N_2497,N_2428,N_2467);
nor U2498 (N_2498,N_2468,N_2460);
nor U2499 (N_2499,N_2419,N_2462);
nor U2500 (N_2500,N_2449,N_2439);
nor U2501 (N_2501,N_2443,N_2471);
nand U2502 (N_2502,N_2451,N_2435);
nor U2503 (N_2503,N_2469,N_2423);
nand U2504 (N_2504,N_2465,N_2458);
and U2505 (N_2505,N_2420,N_2412);
or U2506 (N_2506,N_2446,N_2457);
and U2507 (N_2507,N_2442,N_2426);
xnor U2508 (N_2508,N_2470,N_2411);
nor U2509 (N_2509,N_2472,N_2415);
nor U2510 (N_2510,N_2463,N_2417);
and U2511 (N_2511,N_2404,N_2450);
nor U2512 (N_2512,N_2431,N_2446);
or U2513 (N_2513,N_2424,N_2412);
nor U2514 (N_2514,N_2457,N_2407);
nor U2515 (N_2515,N_2464,N_2442);
nand U2516 (N_2516,N_2472,N_2435);
or U2517 (N_2517,N_2403,N_2421);
or U2518 (N_2518,N_2400,N_2470);
nor U2519 (N_2519,N_2463,N_2441);
and U2520 (N_2520,N_2439,N_2417);
xnor U2521 (N_2521,N_2420,N_2400);
and U2522 (N_2522,N_2408,N_2465);
and U2523 (N_2523,N_2402,N_2466);
and U2524 (N_2524,N_2428,N_2409);
nor U2525 (N_2525,N_2400,N_2438);
and U2526 (N_2526,N_2423,N_2410);
nand U2527 (N_2527,N_2462,N_2452);
nor U2528 (N_2528,N_2438,N_2456);
or U2529 (N_2529,N_2417,N_2409);
nor U2530 (N_2530,N_2442,N_2437);
or U2531 (N_2531,N_2439,N_2441);
or U2532 (N_2532,N_2450,N_2462);
nand U2533 (N_2533,N_2437,N_2431);
nor U2534 (N_2534,N_2433,N_2421);
nand U2535 (N_2535,N_2457,N_2410);
nand U2536 (N_2536,N_2453,N_2412);
nand U2537 (N_2537,N_2402,N_2432);
nand U2538 (N_2538,N_2403,N_2453);
or U2539 (N_2539,N_2416,N_2451);
and U2540 (N_2540,N_2463,N_2472);
and U2541 (N_2541,N_2420,N_2416);
and U2542 (N_2542,N_2413,N_2405);
xor U2543 (N_2543,N_2445,N_2449);
nor U2544 (N_2544,N_2408,N_2411);
nor U2545 (N_2545,N_2474,N_2453);
nor U2546 (N_2546,N_2406,N_2456);
nor U2547 (N_2547,N_2463,N_2401);
nand U2548 (N_2548,N_2444,N_2467);
or U2549 (N_2549,N_2419,N_2472);
and U2550 (N_2550,N_2516,N_2533);
or U2551 (N_2551,N_2487,N_2532);
nand U2552 (N_2552,N_2536,N_2511);
or U2553 (N_2553,N_2549,N_2480);
or U2554 (N_2554,N_2504,N_2538);
nor U2555 (N_2555,N_2489,N_2479);
nand U2556 (N_2556,N_2535,N_2527);
and U2557 (N_2557,N_2541,N_2512);
nor U2558 (N_2558,N_2523,N_2503);
nand U2559 (N_2559,N_2542,N_2495);
and U2560 (N_2560,N_2492,N_2507);
xor U2561 (N_2561,N_2546,N_2505);
and U2562 (N_2562,N_2486,N_2501);
nor U2563 (N_2563,N_2484,N_2528);
and U2564 (N_2564,N_2478,N_2510);
nor U2565 (N_2565,N_2509,N_2498);
and U2566 (N_2566,N_2494,N_2513);
nand U2567 (N_2567,N_2502,N_2529);
or U2568 (N_2568,N_2485,N_2517);
or U2569 (N_2569,N_2481,N_2482);
and U2570 (N_2570,N_2518,N_2539);
and U2571 (N_2571,N_2525,N_2496);
nand U2572 (N_2572,N_2475,N_2477);
or U2573 (N_2573,N_2497,N_2514);
nand U2574 (N_2574,N_2520,N_2534);
nor U2575 (N_2575,N_2524,N_2548);
and U2576 (N_2576,N_2547,N_2515);
nand U2577 (N_2577,N_2521,N_2519);
nor U2578 (N_2578,N_2522,N_2490);
nor U2579 (N_2579,N_2500,N_2537);
nand U2580 (N_2580,N_2493,N_2491);
or U2581 (N_2581,N_2543,N_2476);
nand U2582 (N_2582,N_2488,N_2508);
nor U2583 (N_2583,N_2540,N_2483);
nand U2584 (N_2584,N_2506,N_2499);
or U2585 (N_2585,N_2544,N_2526);
nand U2586 (N_2586,N_2531,N_2545);
nand U2587 (N_2587,N_2530,N_2525);
or U2588 (N_2588,N_2534,N_2481);
nand U2589 (N_2589,N_2476,N_2502);
nand U2590 (N_2590,N_2519,N_2502);
and U2591 (N_2591,N_2494,N_2476);
or U2592 (N_2592,N_2543,N_2530);
or U2593 (N_2593,N_2533,N_2506);
nand U2594 (N_2594,N_2506,N_2515);
and U2595 (N_2595,N_2496,N_2506);
xor U2596 (N_2596,N_2483,N_2517);
or U2597 (N_2597,N_2508,N_2539);
or U2598 (N_2598,N_2548,N_2493);
and U2599 (N_2599,N_2520,N_2481);
nor U2600 (N_2600,N_2530,N_2494);
or U2601 (N_2601,N_2491,N_2506);
nand U2602 (N_2602,N_2510,N_2519);
nand U2603 (N_2603,N_2534,N_2477);
nand U2604 (N_2604,N_2548,N_2538);
or U2605 (N_2605,N_2503,N_2495);
or U2606 (N_2606,N_2483,N_2488);
nand U2607 (N_2607,N_2489,N_2514);
nand U2608 (N_2608,N_2478,N_2502);
nand U2609 (N_2609,N_2502,N_2515);
nand U2610 (N_2610,N_2481,N_2486);
and U2611 (N_2611,N_2531,N_2490);
nor U2612 (N_2612,N_2491,N_2526);
and U2613 (N_2613,N_2500,N_2518);
nand U2614 (N_2614,N_2527,N_2489);
nand U2615 (N_2615,N_2496,N_2527);
nor U2616 (N_2616,N_2489,N_2529);
nor U2617 (N_2617,N_2504,N_2490);
and U2618 (N_2618,N_2510,N_2477);
or U2619 (N_2619,N_2539,N_2492);
nor U2620 (N_2620,N_2516,N_2510);
nand U2621 (N_2621,N_2494,N_2503);
xnor U2622 (N_2622,N_2527,N_2477);
and U2623 (N_2623,N_2478,N_2519);
nor U2624 (N_2624,N_2533,N_2484);
or U2625 (N_2625,N_2553,N_2555);
or U2626 (N_2626,N_2585,N_2573);
and U2627 (N_2627,N_2557,N_2579);
nor U2628 (N_2628,N_2615,N_2578);
or U2629 (N_2629,N_2570,N_2592);
and U2630 (N_2630,N_2582,N_2564);
nand U2631 (N_2631,N_2551,N_2594);
nor U2632 (N_2632,N_2565,N_2608);
nor U2633 (N_2633,N_2589,N_2561);
nand U2634 (N_2634,N_2568,N_2558);
nand U2635 (N_2635,N_2621,N_2622);
xnor U2636 (N_2636,N_2550,N_2617);
or U2637 (N_2637,N_2599,N_2614);
or U2638 (N_2638,N_2588,N_2576);
nand U2639 (N_2639,N_2566,N_2597);
and U2640 (N_2640,N_2569,N_2612);
or U2641 (N_2641,N_2580,N_2616);
nor U2642 (N_2642,N_2602,N_2562);
and U2643 (N_2643,N_2611,N_2577);
nand U2644 (N_2644,N_2607,N_2604);
nor U2645 (N_2645,N_2563,N_2600);
nand U2646 (N_2646,N_2575,N_2590);
nor U2647 (N_2647,N_2587,N_2581);
and U2648 (N_2648,N_2552,N_2620);
nand U2649 (N_2649,N_2609,N_2583);
nand U2650 (N_2650,N_2574,N_2572);
nand U2651 (N_2651,N_2605,N_2598);
nor U2652 (N_2652,N_2567,N_2596);
xnor U2653 (N_2653,N_2619,N_2624);
nand U2654 (N_2654,N_2584,N_2591);
or U2655 (N_2655,N_2603,N_2571);
and U2656 (N_2656,N_2560,N_2554);
nor U2657 (N_2657,N_2559,N_2623);
xor U2658 (N_2658,N_2556,N_2610);
and U2659 (N_2659,N_2613,N_2586);
or U2660 (N_2660,N_2593,N_2606);
nor U2661 (N_2661,N_2601,N_2595);
or U2662 (N_2662,N_2618,N_2610);
and U2663 (N_2663,N_2609,N_2559);
and U2664 (N_2664,N_2579,N_2611);
or U2665 (N_2665,N_2550,N_2579);
nand U2666 (N_2666,N_2571,N_2588);
nor U2667 (N_2667,N_2572,N_2605);
or U2668 (N_2668,N_2580,N_2556);
xor U2669 (N_2669,N_2589,N_2554);
or U2670 (N_2670,N_2610,N_2595);
nor U2671 (N_2671,N_2583,N_2608);
or U2672 (N_2672,N_2600,N_2568);
nor U2673 (N_2673,N_2623,N_2620);
nand U2674 (N_2674,N_2603,N_2598);
xor U2675 (N_2675,N_2565,N_2593);
nor U2676 (N_2676,N_2616,N_2554);
nand U2677 (N_2677,N_2582,N_2614);
and U2678 (N_2678,N_2613,N_2603);
nor U2679 (N_2679,N_2624,N_2616);
and U2680 (N_2680,N_2575,N_2593);
nor U2681 (N_2681,N_2624,N_2603);
or U2682 (N_2682,N_2552,N_2615);
nand U2683 (N_2683,N_2573,N_2584);
nand U2684 (N_2684,N_2550,N_2563);
and U2685 (N_2685,N_2558,N_2581);
and U2686 (N_2686,N_2613,N_2623);
nand U2687 (N_2687,N_2585,N_2570);
or U2688 (N_2688,N_2570,N_2556);
or U2689 (N_2689,N_2563,N_2603);
or U2690 (N_2690,N_2595,N_2556);
or U2691 (N_2691,N_2578,N_2601);
nor U2692 (N_2692,N_2596,N_2564);
nand U2693 (N_2693,N_2561,N_2569);
nand U2694 (N_2694,N_2613,N_2606);
nand U2695 (N_2695,N_2577,N_2564);
nor U2696 (N_2696,N_2561,N_2592);
and U2697 (N_2697,N_2597,N_2556);
and U2698 (N_2698,N_2592,N_2581);
nand U2699 (N_2699,N_2563,N_2591);
and U2700 (N_2700,N_2631,N_2630);
nand U2701 (N_2701,N_2652,N_2679);
and U2702 (N_2702,N_2666,N_2625);
nand U2703 (N_2703,N_2648,N_2654);
xnor U2704 (N_2704,N_2682,N_2669);
and U2705 (N_2705,N_2650,N_2696);
or U2706 (N_2706,N_2626,N_2659);
nor U2707 (N_2707,N_2646,N_2628);
and U2708 (N_2708,N_2661,N_2668);
nor U2709 (N_2709,N_2698,N_2673);
nor U2710 (N_2710,N_2687,N_2664);
nor U2711 (N_2711,N_2642,N_2694);
nor U2712 (N_2712,N_2627,N_2685);
and U2713 (N_2713,N_2655,N_2690);
or U2714 (N_2714,N_2644,N_2662);
nand U2715 (N_2715,N_2635,N_2643);
nand U2716 (N_2716,N_2653,N_2640);
xnor U2717 (N_2717,N_2693,N_2672);
nand U2718 (N_2718,N_2692,N_2637);
nor U2719 (N_2719,N_2632,N_2629);
nor U2720 (N_2720,N_2667,N_2651);
or U2721 (N_2721,N_2678,N_2645);
xor U2722 (N_2722,N_2681,N_2674);
nand U2723 (N_2723,N_2647,N_2689);
nor U2724 (N_2724,N_2649,N_2665);
or U2725 (N_2725,N_2660,N_2697);
nand U2726 (N_2726,N_2691,N_2677);
and U2727 (N_2727,N_2684,N_2641);
and U2728 (N_2728,N_2683,N_2658);
nor U2729 (N_2729,N_2680,N_2688);
nor U2730 (N_2730,N_2676,N_2695);
nand U2731 (N_2731,N_2675,N_2670);
nor U2732 (N_2732,N_2639,N_2671);
nor U2733 (N_2733,N_2657,N_2699);
and U2734 (N_2734,N_2634,N_2633);
nor U2735 (N_2735,N_2663,N_2638);
nand U2736 (N_2736,N_2636,N_2656);
nor U2737 (N_2737,N_2686,N_2648);
or U2738 (N_2738,N_2631,N_2629);
and U2739 (N_2739,N_2647,N_2694);
and U2740 (N_2740,N_2693,N_2668);
nor U2741 (N_2741,N_2645,N_2668);
nor U2742 (N_2742,N_2651,N_2675);
and U2743 (N_2743,N_2697,N_2635);
nor U2744 (N_2744,N_2630,N_2657);
nand U2745 (N_2745,N_2677,N_2666);
or U2746 (N_2746,N_2667,N_2657);
nand U2747 (N_2747,N_2650,N_2645);
or U2748 (N_2748,N_2680,N_2647);
nor U2749 (N_2749,N_2660,N_2635);
xor U2750 (N_2750,N_2644,N_2656);
nand U2751 (N_2751,N_2670,N_2666);
nand U2752 (N_2752,N_2646,N_2681);
nor U2753 (N_2753,N_2670,N_2659);
and U2754 (N_2754,N_2667,N_2690);
nor U2755 (N_2755,N_2634,N_2692);
and U2756 (N_2756,N_2667,N_2638);
nand U2757 (N_2757,N_2648,N_2699);
nand U2758 (N_2758,N_2638,N_2680);
xnor U2759 (N_2759,N_2695,N_2698);
nand U2760 (N_2760,N_2668,N_2674);
nor U2761 (N_2761,N_2680,N_2650);
and U2762 (N_2762,N_2685,N_2691);
nor U2763 (N_2763,N_2656,N_2659);
or U2764 (N_2764,N_2679,N_2647);
and U2765 (N_2765,N_2659,N_2694);
and U2766 (N_2766,N_2672,N_2669);
or U2767 (N_2767,N_2679,N_2654);
or U2768 (N_2768,N_2634,N_2659);
nor U2769 (N_2769,N_2645,N_2633);
and U2770 (N_2770,N_2628,N_2684);
and U2771 (N_2771,N_2631,N_2668);
nand U2772 (N_2772,N_2654,N_2652);
nor U2773 (N_2773,N_2633,N_2631);
nor U2774 (N_2774,N_2666,N_2694);
or U2775 (N_2775,N_2749,N_2722);
and U2776 (N_2776,N_2743,N_2774);
xor U2777 (N_2777,N_2710,N_2754);
nand U2778 (N_2778,N_2700,N_2747);
and U2779 (N_2779,N_2746,N_2708);
nand U2780 (N_2780,N_2760,N_2733);
or U2781 (N_2781,N_2721,N_2735);
or U2782 (N_2782,N_2716,N_2758);
or U2783 (N_2783,N_2728,N_2729);
or U2784 (N_2784,N_2711,N_2740);
and U2785 (N_2785,N_2771,N_2709);
and U2786 (N_2786,N_2703,N_2772);
or U2787 (N_2787,N_2765,N_2744);
or U2788 (N_2788,N_2705,N_2713);
nand U2789 (N_2789,N_2764,N_2770);
nand U2790 (N_2790,N_2753,N_2755);
nand U2791 (N_2791,N_2720,N_2768);
or U2792 (N_2792,N_2773,N_2706);
nor U2793 (N_2793,N_2707,N_2714);
nor U2794 (N_2794,N_2741,N_2704);
or U2795 (N_2795,N_2701,N_2727);
and U2796 (N_2796,N_2732,N_2763);
nand U2797 (N_2797,N_2745,N_2750);
and U2798 (N_2798,N_2767,N_2756);
xor U2799 (N_2799,N_2725,N_2757);
or U2800 (N_2800,N_2712,N_2731);
and U2801 (N_2801,N_2736,N_2739);
or U2802 (N_2802,N_2702,N_2738);
nor U2803 (N_2803,N_2748,N_2742);
nand U2804 (N_2804,N_2759,N_2730);
and U2805 (N_2805,N_2734,N_2769);
nand U2806 (N_2806,N_2762,N_2724);
and U2807 (N_2807,N_2718,N_2726);
xor U2808 (N_2808,N_2717,N_2719);
and U2809 (N_2809,N_2737,N_2715);
nand U2810 (N_2810,N_2751,N_2761);
nand U2811 (N_2811,N_2752,N_2723);
nand U2812 (N_2812,N_2766,N_2768);
and U2813 (N_2813,N_2756,N_2753);
nor U2814 (N_2814,N_2722,N_2739);
and U2815 (N_2815,N_2718,N_2767);
nand U2816 (N_2816,N_2747,N_2711);
nand U2817 (N_2817,N_2755,N_2720);
nor U2818 (N_2818,N_2758,N_2763);
nand U2819 (N_2819,N_2768,N_2759);
or U2820 (N_2820,N_2763,N_2741);
nor U2821 (N_2821,N_2743,N_2770);
and U2822 (N_2822,N_2750,N_2709);
nor U2823 (N_2823,N_2735,N_2729);
nand U2824 (N_2824,N_2731,N_2729);
nor U2825 (N_2825,N_2745,N_2774);
nor U2826 (N_2826,N_2761,N_2733);
and U2827 (N_2827,N_2717,N_2705);
nand U2828 (N_2828,N_2756,N_2763);
nor U2829 (N_2829,N_2768,N_2755);
or U2830 (N_2830,N_2744,N_2758);
nand U2831 (N_2831,N_2772,N_2700);
nand U2832 (N_2832,N_2727,N_2753);
or U2833 (N_2833,N_2703,N_2764);
nor U2834 (N_2834,N_2737,N_2739);
nand U2835 (N_2835,N_2735,N_2762);
or U2836 (N_2836,N_2705,N_2757);
nor U2837 (N_2837,N_2772,N_2711);
nand U2838 (N_2838,N_2704,N_2751);
or U2839 (N_2839,N_2743,N_2771);
or U2840 (N_2840,N_2753,N_2716);
nand U2841 (N_2841,N_2751,N_2771);
nor U2842 (N_2842,N_2756,N_2713);
or U2843 (N_2843,N_2729,N_2770);
nand U2844 (N_2844,N_2735,N_2713);
nor U2845 (N_2845,N_2746,N_2756);
and U2846 (N_2846,N_2763,N_2707);
nor U2847 (N_2847,N_2706,N_2709);
nor U2848 (N_2848,N_2730,N_2712);
nor U2849 (N_2849,N_2766,N_2724);
or U2850 (N_2850,N_2847,N_2832);
and U2851 (N_2851,N_2809,N_2798);
or U2852 (N_2852,N_2831,N_2840);
nor U2853 (N_2853,N_2826,N_2801);
nand U2854 (N_2854,N_2796,N_2844);
nor U2855 (N_2855,N_2810,N_2775);
or U2856 (N_2856,N_2778,N_2811);
nor U2857 (N_2857,N_2817,N_2837);
and U2858 (N_2858,N_2833,N_2821);
nor U2859 (N_2859,N_2839,N_2792);
and U2860 (N_2860,N_2830,N_2827);
or U2861 (N_2861,N_2783,N_2802);
xnor U2862 (N_2862,N_2834,N_2784);
nor U2863 (N_2863,N_2838,N_2780);
nand U2864 (N_2864,N_2790,N_2806);
or U2865 (N_2865,N_2781,N_2814);
or U2866 (N_2866,N_2788,N_2828);
and U2867 (N_2867,N_2829,N_2787);
nor U2868 (N_2868,N_2800,N_2779);
nand U2869 (N_2869,N_2843,N_2799);
nor U2870 (N_2870,N_2794,N_2789);
xor U2871 (N_2871,N_2804,N_2808);
nand U2872 (N_2872,N_2824,N_2813);
xor U2873 (N_2873,N_2818,N_2777);
nor U2874 (N_2874,N_2807,N_2812);
nand U2875 (N_2875,N_2791,N_2819);
nor U2876 (N_2876,N_2825,N_2797);
nor U2877 (N_2877,N_2842,N_2782);
nor U2878 (N_2878,N_2793,N_2841);
nand U2879 (N_2879,N_2846,N_2835);
nand U2880 (N_2880,N_2836,N_2848);
or U2881 (N_2881,N_2822,N_2795);
and U2882 (N_2882,N_2845,N_2785);
or U2883 (N_2883,N_2776,N_2816);
or U2884 (N_2884,N_2803,N_2820);
or U2885 (N_2885,N_2805,N_2849);
and U2886 (N_2886,N_2815,N_2786);
nand U2887 (N_2887,N_2823,N_2797);
xor U2888 (N_2888,N_2825,N_2836);
nor U2889 (N_2889,N_2821,N_2832);
and U2890 (N_2890,N_2804,N_2844);
nor U2891 (N_2891,N_2775,N_2796);
nor U2892 (N_2892,N_2793,N_2780);
and U2893 (N_2893,N_2779,N_2795);
or U2894 (N_2894,N_2834,N_2799);
or U2895 (N_2895,N_2777,N_2847);
nor U2896 (N_2896,N_2788,N_2812);
or U2897 (N_2897,N_2815,N_2780);
nor U2898 (N_2898,N_2846,N_2787);
and U2899 (N_2899,N_2791,N_2820);
nor U2900 (N_2900,N_2839,N_2789);
or U2901 (N_2901,N_2819,N_2830);
or U2902 (N_2902,N_2795,N_2803);
xnor U2903 (N_2903,N_2782,N_2818);
or U2904 (N_2904,N_2784,N_2783);
and U2905 (N_2905,N_2833,N_2839);
or U2906 (N_2906,N_2787,N_2824);
and U2907 (N_2907,N_2793,N_2825);
and U2908 (N_2908,N_2789,N_2786);
nor U2909 (N_2909,N_2831,N_2813);
nand U2910 (N_2910,N_2823,N_2793);
nand U2911 (N_2911,N_2825,N_2801);
nand U2912 (N_2912,N_2821,N_2795);
nor U2913 (N_2913,N_2793,N_2797);
and U2914 (N_2914,N_2807,N_2814);
or U2915 (N_2915,N_2827,N_2817);
or U2916 (N_2916,N_2826,N_2829);
or U2917 (N_2917,N_2830,N_2792);
nor U2918 (N_2918,N_2822,N_2810);
and U2919 (N_2919,N_2800,N_2808);
nor U2920 (N_2920,N_2784,N_2809);
xnor U2921 (N_2921,N_2819,N_2794);
nor U2922 (N_2922,N_2811,N_2839);
and U2923 (N_2923,N_2779,N_2849);
or U2924 (N_2924,N_2775,N_2848);
and U2925 (N_2925,N_2899,N_2881);
or U2926 (N_2926,N_2870,N_2887);
and U2927 (N_2927,N_2894,N_2914);
or U2928 (N_2928,N_2867,N_2898);
nand U2929 (N_2929,N_2880,N_2916);
nor U2930 (N_2930,N_2893,N_2874);
or U2931 (N_2931,N_2920,N_2905);
nor U2932 (N_2932,N_2897,N_2908);
nand U2933 (N_2933,N_2918,N_2903);
nand U2934 (N_2934,N_2924,N_2858);
or U2935 (N_2935,N_2868,N_2892);
nor U2936 (N_2936,N_2857,N_2891);
nor U2937 (N_2937,N_2910,N_2878);
or U2938 (N_2938,N_2909,N_2882);
and U2939 (N_2939,N_2879,N_2862);
nor U2940 (N_2940,N_2919,N_2871);
and U2941 (N_2941,N_2866,N_2861);
or U2942 (N_2942,N_2923,N_2912);
or U2943 (N_2943,N_2900,N_2852);
and U2944 (N_2944,N_2855,N_2851);
nor U2945 (N_2945,N_2902,N_2883);
or U2946 (N_2946,N_2863,N_2917);
and U2947 (N_2947,N_2895,N_2854);
or U2948 (N_2948,N_2906,N_2850);
or U2949 (N_2949,N_2859,N_2904);
nor U2950 (N_2950,N_2921,N_2884);
or U2951 (N_2951,N_2888,N_2853);
nor U2952 (N_2952,N_2890,N_2915);
nand U2953 (N_2953,N_2877,N_2864);
xnor U2954 (N_2954,N_2913,N_2896);
nand U2955 (N_2955,N_2886,N_2911);
and U2956 (N_2956,N_2901,N_2885);
nor U2957 (N_2957,N_2876,N_2922);
and U2958 (N_2958,N_2872,N_2873);
or U2959 (N_2959,N_2875,N_2889);
and U2960 (N_2960,N_2865,N_2907);
or U2961 (N_2961,N_2860,N_2856);
or U2962 (N_2962,N_2869,N_2919);
nor U2963 (N_2963,N_2904,N_2896);
nand U2964 (N_2964,N_2890,N_2923);
nand U2965 (N_2965,N_2884,N_2899);
xor U2966 (N_2966,N_2894,N_2915);
nor U2967 (N_2967,N_2851,N_2863);
nor U2968 (N_2968,N_2866,N_2872);
or U2969 (N_2969,N_2881,N_2869);
nand U2970 (N_2970,N_2877,N_2862);
xor U2971 (N_2971,N_2881,N_2886);
nand U2972 (N_2972,N_2876,N_2907);
and U2973 (N_2973,N_2909,N_2858);
nor U2974 (N_2974,N_2901,N_2903);
nand U2975 (N_2975,N_2900,N_2879);
and U2976 (N_2976,N_2852,N_2909);
and U2977 (N_2977,N_2907,N_2872);
nand U2978 (N_2978,N_2859,N_2915);
nor U2979 (N_2979,N_2872,N_2881);
or U2980 (N_2980,N_2886,N_2888);
nor U2981 (N_2981,N_2897,N_2871);
nand U2982 (N_2982,N_2868,N_2885);
nor U2983 (N_2983,N_2873,N_2889);
and U2984 (N_2984,N_2850,N_2877);
nor U2985 (N_2985,N_2900,N_2904);
nor U2986 (N_2986,N_2856,N_2854);
and U2987 (N_2987,N_2881,N_2911);
or U2988 (N_2988,N_2924,N_2869);
nand U2989 (N_2989,N_2856,N_2908);
nor U2990 (N_2990,N_2922,N_2851);
xor U2991 (N_2991,N_2867,N_2861);
nand U2992 (N_2992,N_2882,N_2911);
and U2993 (N_2993,N_2863,N_2885);
nor U2994 (N_2994,N_2916,N_2893);
or U2995 (N_2995,N_2876,N_2883);
nor U2996 (N_2996,N_2907,N_2905);
or U2997 (N_2997,N_2855,N_2869);
nor U2998 (N_2998,N_2854,N_2878);
nor U2999 (N_2999,N_2851,N_2895);
and UO_0 (O_0,N_2926,N_2989);
nand UO_1 (O_1,N_2993,N_2961);
nor UO_2 (O_2,N_2974,N_2939);
and UO_3 (O_3,N_2930,N_2985);
nor UO_4 (O_4,N_2957,N_2978);
and UO_5 (O_5,N_2990,N_2959);
or UO_6 (O_6,N_2952,N_2969);
and UO_7 (O_7,N_2931,N_2938);
or UO_8 (O_8,N_2946,N_2945);
xor UO_9 (O_9,N_2970,N_2963);
nor UO_10 (O_10,N_2940,N_2951);
nor UO_11 (O_11,N_2972,N_2986);
nor UO_12 (O_12,N_2984,N_2953);
nor UO_13 (O_13,N_2997,N_2964);
and UO_14 (O_14,N_2928,N_2994);
or UO_15 (O_15,N_2991,N_2956);
nor UO_16 (O_16,N_2998,N_2979);
nor UO_17 (O_17,N_2935,N_2943);
nor UO_18 (O_18,N_2934,N_2947);
or UO_19 (O_19,N_2958,N_2929);
or UO_20 (O_20,N_2971,N_2982);
nor UO_21 (O_21,N_2933,N_2983);
nor UO_22 (O_22,N_2941,N_2949);
or UO_23 (O_23,N_2996,N_2932);
nand UO_24 (O_24,N_2925,N_2987);
nor UO_25 (O_25,N_2976,N_2936);
or UO_26 (O_26,N_2999,N_2968);
and UO_27 (O_27,N_2948,N_2955);
and UO_28 (O_28,N_2954,N_2960);
nand UO_29 (O_29,N_2950,N_2981);
or UO_30 (O_30,N_2966,N_2992);
nor UO_31 (O_31,N_2967,N_2962);
nand UO_32 (O_32,N_2927,N_2977);
nand UO_33 (O_33,N_2995,N_2942);
nor UO_34 (O_34,N_2965,N_2973);
and UO_35 (O_35,N_2980,N_2975);
nor UO_36 (O_36,N_2937,N_2988);
nor UO_37 (O_37,N_2944,N_2982);
nand UO_38 (O_38,N_2936,N_2927);
or UO_39 (O_39,N_2954,N_2981);
and UO_40 (O_40,N_2978,N_2991);
nand UO_41 (O_41,N_2989,N_2985);
nor UO_42 (O_42,N_2998,N_2969);
or UO_43 (O_43,N_2965,N_2948);
and UO_44 (O_44,N_2943,N_2995);
nor UO_45 (O_45,N_2966,N_2945);
xor UO_46 (O_46,N_2954,N_2996);
nor UO_47 (O_47,N_2984,N_2962);
nand UO_48 (O_48,N_2971,N_2994);
or UO_49 (O_49,N_2943,N_2994);
nand UO_50 (O_50,N_2951,N_2964);
nand UO_51 (O_51,N_2959,N_2967);
and UO_52 (O_52,N_2992,N_2993);
and UO_53 (O_53,N_2963,N_2955);
and UO_54 (O_54,N_2966,N_2939);
nand UO_55 (O_55,N_2987,N_2931);
nor UO_56 (O_56,N_2927,N_2998);
or UO_57 (O_57,N_2998,N_2984);
and UO_58 (O_58,N_2987,N_2970);
nor UO_59 (O_59,N_2931,N_2949);
nand UO_60 (O_60,N_2965,N_2988);
or UO_61 (O_61,N_2946,N_2953);
or UO_62 (O_62,N_2945,N_2982);
or UO_63 (O_63,N_2938,N_2955);
or UO_64 (O_64,N_2932,N_2962);
or UO_65 (O_65,N_2949,N_2989);
xnor UO_66 (O_66,N_2973,N_2980);
and UO_67 (O_67,N_2938,N_2932);
or UO_68 (O_68,N_2966,N_2930);
nor UO_69 (O_69,N_2967,N_2939);
or UO_70 (O_70,N_2962,N_2944);
or UO_71 (O_71,N_2998,N_2941);
nor UO_72 (O_72,N_2961,N_2945);
nor UO_73 (O_73,N_2936,N_2961);
and UO_74 (O_74,N_2961,N_2938);
xnor UO_75 (O_75,N_2982,N_2958);
nand UO_76 (O_76,N_2962,N_2933);
and UO_77 (O_77,N_2926,N_2971);
and UO_78 (O_78,N_2984,N_2929);
and UO_79 (O_79,N_2953,N_2932);
nand UO_80 (O_80,N_2972,N_2989);
and UO_81 (O_81,N_2982,N_2952);
nand UO_82 (O_82,N_2941,N_2981);
or UO_83 (O_83,N_2925,N_2926);
and UO_84 (O_84,N_2976,N_2996);
nor UO_85 (O_85,N_2940,N_2958);
nand UO_86 (O_86,N_2927,N_2946);
or UO_87 (O_87,N_2948,N_2970);
and UO_88 (O_88,N_2934,N_2940);
and UO_89 (O_89,N_2969,N_2974);
or UO_90 (O_90,N_2927,N_2976);
and UO_91 (O_91,N_2985,N_2993);
and UO_92 (O_92,N_2945,N_2952);
or UO_93 (O_93,N_2998,N_2966);
or UO_94 (O_94,N_2926,N_2961);
nand UO_95 (O_95,N_2942,N_2978);
and UO_96 (O_96,N_2941,N_2927);
nand UO_97 (O_97,N_2968,N_2948);
nand UO_98 (O_98,N_2945,N_2926);
nor UO_99 (O_99,N_2946,N_2952);
xnor UO_100 (O_100,N_2949,N_2973);
nor UO_101 (O_101,N_2986,N_2925);
nand UO_102 (O_102,N_2947,N_2941);
and UO_103 (O_103,N_2954,N_2958);
nor UO_104 (O_104,N_2935,N_2981);
nand UO_105 (O_105,N_2955,N_2964);
nand UO_106 (O_106,N_2999,N_2929);
nand UO_107 (O_107,N_2930,N_2999);
nor UO_108 (O_108,N_2934,N_2970);
nor UO_109 (O_109,N_2939,N_2965);
or UO_110 (O_110,N_2960,N_2955);
nand UO_111 (O_111,N_2938,N_2958);
nand UO_112 (O_112,N_2932,N_2965);
or UO_113 (O_113,N_2960,N_2975);
nor UO_114 (O_114,N_2994,N_2933);
and UO_115 (O_115,N_2948,N_2971);
or UO_116 (O_116,N_2986,N_2944);
and UO_117 (O_117,N_2968,N_2995);
nor UO_118 (O_118,N_2971,N_2961);
or UO_119 (O_119,N_2983,N_2964);
and UO_120 (O_120,N_2933,N_2969);
nor UO_121 (O_121,N_2976,N_2944);
nor UO_122 (O_122,N_2951,N_2965);
nor UO_123 (O_123,N_2988,N_2967);
nand UO_124 (O_124,N_2951,N_2968);
nor UO_125 (O_125,N_2927,N_2926);
or UO_126 (O_126,N_2955,N_2954);
and UO_127 (O_127,N_2973,N_2954);
and UO_128 (O_128,N_2999,N_2983);
nand UO_129 (O_129,N_2938,N_2936);
nand UO_130 (O_130,N_2964,N_2947);
or UO_131 (O_131,N_2989,N_2994);
nor UO_132 (O_132,N_2938,N_2953);
and UO_133 (O_133,N_2932,N_2972);
or UO_134 (O_134,N_2987,N_2941);
and UO_135 (O_135,N_2961,N_2944);
or UO_136 (O_136,N_2947,N_2986);
or UO_137 (O_137,N_2947,N_2987);
nor UO_138 (O_138,N_2991,N_2932);
nor UO_139 (O_139,N_2999,N_2928);
nand UO_140 (O_140,N_2965,N_2944);
nor UO_141 (O_141,N_2967,N_2972);
and UO_142 (O_142,N_2929,N_2942);
nor UO_143 (O_143,N_2949,N_2968);
xnor UO_144 (O_144,N_2986,N_2926);
nor UO_145 (O_145,N_2935,N_2985);
or UO_146 (O_146,N_2961,N_2982);
nand UO_147 (O_147,N_2953,N_2959);
or UO_148 (O_148,N_2991,N_2933);
nand UO_149 (O_149,N_2929,N_2959);
or UO_150 (O_150,N_2990,N_2952);
nand UO_151 (O_151,N_2935,N_2995);
or UO_152 (O_152,N_2934,N_2983);
nand UO_153 (O_153,N_2948,N_2973);
or UO_154 (O_154,N_2960,N_2988);
nand UO_155 (O_155,N_2955,N_2994);
and UO_156 (O_156,N_2979,N_2992);
nor UO_157 (O_157,N_2938,N_2935);
nand UO_158 (O_158,N_2989,N_2958);
and UO_159 (O_159,N_2979,N_2961);
or UO_160 (O_160,N_2930,N_2948);
nand UO_161 (O_161,N_2993,N_2928);
or UO_162 (O_162,N_2992,N_2949);
or UO_163 (O_163,N_2972,N_2975);
nor UO_164 (O_164,N_2973,N_2957);
xor UO_165 (O_165,N_2933,N_2930);
or UO_166 (O_166,N_2934,N_2950);
and UO_167 (O_167,N_2948,N_2962);
or UO_168 (O_168,N_2977,N_2950);
nor UO_169 (O_169,N_2944,N_2949);
and UO_170 (O_170,N_2963,N_2928);
or UO_171 (O_171,N_2978,N_2945);
or UO_172 (O_172,N_2969,N_2948);
nor UO_173 (O_173,N_2986,N_2960);
or UO_174 (O_174,N_2947,N_2926);
nand UO_175 (O_175,N_2972,N_2951);
nor UO_176 (O_176,N_2986,N_2998);
nand UO_177 (O_177,N_2961,N_2931);
nand UO_178 (O_178,N_2951,N_2950);
nor UO_179 (O_179,N_2984,N_2992);
or UO_180 (O_180,N_2984,N_2946);
nor UO_181 (O_181,N_2992,N_2925);
nand UO_182 (O_182,N_2978,N_2933);
or UO_183 (O_183,N_2998,N_2945);
nor UO_184 (O_184,N_2994,N_2978);
nand UO_185 (O_185,N_2973,N_2977);
or UO_186 (O_186,N_2941,N_2964);
and UO_187 (O_187,N_2940,N_2998);
or UO_188 (O_188,N_2967,N_2982);
nand UO_189 (O_189,N_2930,N_2971);
and UO_190 (O_190,N_2957,N_2968);
and UO_191 (O_191,N_2944,N_2977);
nand UO_192 (O_192,N_2939,N_2995);
and UO_193 (O_193,N_2951,N_2989);
and UO_194 (O_194,N_2975,N_2986);
nand UO_195 (O_195,N_2991,N_2985);
nor UO_196 (O_196,N_2943,N_2939);
or UO_197 (O_197,N_2931,N_2945);
nor UO_198 (O_198,N_2988,N_2946);
nand UO_199 (O_199,N_2980,N_2996);
nor UO_200 (O_200,N_2980,N_2937);
nor UO_201 (O_201,N_2941,N_2993);
or UO_202 (O_202,N_2955,N_2956);
and UO_203 (O_203,N_2965,N_2971);
nand UO_204 (O_204,N_2943,N_2930);
nor UO_205 (O_205,N_2972,N_2994);
nand UO_206 (O_206,N_2971,N_2950);
nor UO_207 (O_207,N_2974,N_2975);
and UO_208 (O_208,N_2931,N_2946);
or UO_209 (O_209,N_2947,N_2957);
nand UO_210 (O_210,N_2986,N_2932);
and UO_211 (O_211,N_2941,N_2978);
nand UO_212 (O_212,N_2992,N_2980);
nor UO_213 (O_213,N_2943,N_2951);
or UO_214 (O_214,N_2930,N_2975);
or UO_215 (O_215,N_2958,N_2978);
nor UO_216 (O_216,N_2942,N_2939);
nand UO_217 (O_217,N_2958,N_2977);
nor UO_218 (O_218,N_2938,N_2982);
nor UO_219 (O_219,N_2983,N_2952);
nor UO_220 (O_220,N_2948,N_2929);
nor UO_221 (O_221,N_2984,N_2975);
or UO_222 (O_222,N_2937,N_2968);
nor UO_223 (O_223,N_2987,N_2998);
nand UO_224 (O_224,N_2992,N_2998);
and UO_225 (O_225,N_2981,N_2926);
xor UO_226 (O_226,N_2945,N_2937);
and UO_227 (O_227,N_2937,N_2983);
nor UO_228 (O_228,N_2940,N_2969);
nand UO_229 (O_229,N_2977,N_2985);
nand UO_230 (O_230,N_2993,N_2929);
nor UO_231 (O_231,N_2996,N_2979);
or UO_232 (O_232,N_2990,N_2972);
or UO_233 (O_233,N_2959,N_2945);
nand UO_234 (O_234,N_2967,N_2978);
nor UO_235 (O_235,N_2927,N_2985);
and UO_236 (O_236,N_2944,N_2960);
and UO_237 (O_237,N_2995,N_2992);
and UO_238 (O_238,N_2996,N_2952);
nor UO_239 (O_239,N_2947,N_2943);
xnor UO_240 (O_240,N_2964,N_2970);
and UO_241 (O_241,N_2951,N_2971);
nor UO_242 (O_242,N_2929,N_2998);
or UO_243 (O_243,N_2969,N_2987);
and UO_244 (O_244,N_2960,N_2941);
nand UO_245 (O_245,N_2989,N_2971);
and UO_246 (O_246,N_2995,N_2960);
and UO_247 (O_247,N_2944,N_2970);
nor UO_248 (O_248,N_2996,N_2978);
nand UO_249 (O_249,N_2948,N_2956);
or UO_250 (O_250,N_2972,N_2983);
nor UO_251 (O_251,N_2997,N_2984);
nand UO_252 (O_252,N_2996,N_2974);
xnor UO_253 (O_253,N_2936,N_2986);
nand UO_254 (O_254,N_2996,N_2998);
nor UO_255 (O_255,N_2973,N_2962);
and UO_256 (O_256,N_2965,N_2999);
and UO_257 (O_257,N_2953,N_2954);
nor UO_258 (O_258,N_2961,N_2966);
or UO_259 (O_259,N_2979,N_2978);
or UO_260 (O_260,N_2996,N_2931);
nor UO_261 (O_261,N_2935,N_2940);
and UO_262 (O_262,N_2957,N_2966);
nand UO_263 (O_263,N_2969,N_2963);
xnor UO_264 (O_264,N_2965,N_2957);
nand UO_265 (O_265,N_2940,N_2941);
and UO_266 (O_266,N_2986,N_2970);
or UO_267 (O_267,N_2971,N_2940);
or UO_268 (O_268,N_2940,N_2930);
and UO_269 (O_269,N_2938,N_2934);
nor UO_270 (O_270,N_2949,N_2933);
nor UO_271 (O_271,N_2969,N_2936);
and UO_272 (O_272,N_2959,N_2932);
xnor UO_273 (O_273,N_2997,N_2976);
and UO_274 (O_274,N_2957,N_2974);
nand UO_275 (O_275,N_2973,N_2990);
nor UO_276 (O_276,N_2963,N_2999);
or UO_277 (O_277,N_2984,N_2949);
and UO_278 (O_278,N_2967,N_2947);
nor UO_279 (O_279,N_2962,N_2950);
nand UO_280 (O_280,N_2952,N_2948);
and UO_281 (O_281,N_2977,N_2953);
nor UO_282 (O_282,N_2971,N_2929);
nor UO_283 (O_283,N_2990,N_2991);
nor UO_284 (O_284,N_2977,N_2967);
nand UO_285 (O_285,N_2931,N_2986);
or UO_286 (O_286,N_2962,N_2931);
nor UO_287 (O_287,N_2935,N_2986);
nor UO_288 (O_288,N_2984,N_2972);
nand UO_289 (O_289,N_2941,N_2925);
nor UO_290 (O_290,N_2947,N_2969);
or UO_291 (O_291,N_2951,N_2998);
and UO_292 (O_292,N_2932,N_2971);
nor UO_293 (O_293,N_2991,N_2930);
nand UO_294 (O_294,N_2934,N_2956);
nand UO_295 (O_295,N_2954,N_2971);
and UO_296 (O_296,N_2990,N_2944);
and UO_297 (O_297,N_2981,N_2970);
nand UO_298 (O_298,N_2961,N_2968);
and UO_299 (O_299,N_2999,N_2979);
nor UO_300 (O_300,N_2965,N_2980);
or UO_301 (O_301,N_2976,N_2973);
or UO_302 (O_302,N_2949,N_2970);
xnor UO_303 (O_303,N_2951,N_2984);
nor UO_304 (O_304,N_2983,N_2968);
nor UO_305 (O_305,N_2938,N_2943);
nand UO_306 (O_306,N_2964,N_2948);
and UO_307 (O_307,N_2962,N_2929);
or UO_308 (O_308,N_2958,N_2987);
or UO_309 (O_309,N_2926,N_2964);
nor UO_310 (O_310,N_2988,N_2932);
and UO_311 (O_311,N_2950,N_2980);
and UO_312 (O_312,N_2993,N_2963);
nand UO_313 (O_313,N_2935,N_2973);
nand UO_314 (O_314,N_2988,N_2984);
and UO_315 (O_315,N_2947,N_2981);
nand UO_316 (O_316,N_2929,N_2936);
nor UO_317 (O_317,N_2963,N_2965);
or UO_318 (O_318,N_2930,N_2976);
nor UO_319 (O_319,N_2962,N_2978);
or UO_320 (O_320,N_2996,N_2970);
or UO_321 (O_321,N_2965,N_2987);
nor UO_322 (O_322,N_2945,N_2955);
or UO_323 (O_323,N_2953,N_2931);
nor UO_324 (O_324,N_2993,N_2980);
nor UO_325 (O_325,N_2967,N_2974);
nand UO_326 (O_326,N_2931,N_2940);
nand UO_327 (O_327,N_2926,N_2933);
nand UO_328 (O_328,N_2984,N_2933);
xnor UO_329 (O_329,N_2939,N_2977);
nand UO_330 (O_330,N_2993,N_2959);
nor UO_331 (O_331,N_2944,N_2984);
nand UO_332 (O_332,N_2989,N_2973);
nor UO_333 (O_333,N_2962,N_2925);
or UO_334 (O_334,N_2925,N_2928);
xor UO_335 (O_335,N_2948,N_2981);
and UO_336 (O_336,N_2968,N_2935);
nand UO_337 (O_337,N_2997,N_2940);
nand UO_338 (O_338,N_2983,N_2997);
and UO_339 (O_339,N_2925,N_2984);
or UO_340 (O_340,N_2931,N_2937);
and UO_341 (O_341,N_2939,N_2954);
and UO_342 (O_342,N_2997,N_2967);
nand UO_343 (O_343,N_2973,N_2930);
nor UO_344 (O_344,N_2961,N_2930);
or UO_345 (O_345,N_2948,N_2985);
nor UO_346 (O_346,N_2951,N_2973);
and UO_347 (O_347,N_2993,N_2994);
nand UO_348 (O_348,N_2977,N_2932);
and UO_349 (O_349,N_2965,N_2972);
nor UO_350 (O_350,N_2972,N_2943);
or UO_351 (O_351,N_2964,N_2929);
nor UO_352 (O_352,N_2972,N_2931);
and UO_353 (O_353,N_2974,N_2946);
nor UO_354 (O_354,N_2939,N_2952);
or UO_355 (O_355,N_2998,N_2958);
and UO_356 (O_356,N_2934,N_2971);
nor UO_357 (O_357,N_2998,N_2988);
and UO_358 (O_358,N_2941,N_2968);
nor UO_359 (O_359,N_2992,N_2991);
nand UO_360 (O_360,N_2940,N_2991);
nand UO_361 (O_361,N_2932,N_2952);
nand UO_362 (O_362,N_2968,N_2984);
xnor UO_363 (O_363,N_2978,N_2939);
and UO_364 (O_364,N_2977,N_2988);
nor UO_365 (O_365,N_2985,N_2957);
nand UO_366 (O_366,N_2961,N_2997);
nand UO_367 (O_367,N_2956,N_2926);
nor UO_368 (O_368,N_2999,N_2927);
and UO_369 (O_369,N_2994,N_2977);
and UO_370 (O_370,N_2967,N_2957);
and UO_371 (O_371,N_2955,N_2930);
and UO_372 (O_372,N_2970,N_2927);
and UO_373 (O_373,N_2996,N_2969);
nand UO_374 (O_374,N_2933,N_2928);
nor UO_375 (O_375,N_2961,N_2939);
or UO_376 (O_376,N_2974,N_2950);
and UO_377 (O_377,N_2937,N_2967);
or UO_378 (O_378,N_2979,N_2963);
nor UO_379 (O_379,N_2951,N_2997);
or UO_380 (O_380,N_2987,N_2994);
nor UO_381 (O_381,N_2926,N_2931);
or UO_382 (O_382,N_2957,N_2935);
and UO_383 (O_383,N_2960,N_2949);
nor UO_384 (O_384,N_2993,N_2972);
or UO_385 (O_385,N_2956,N_2946);
or UO_386 (O_386,N_2974,N_2984);
nor UO_387 (O_387,N_2929,N_2981);
nand UO_388 (O_388,N_2961,N_2940);
or UO_389 (O_389,N_2983,N_2932);
or UO_390 (O_390,N_2993,N_2944);
xnor UO_391 (O_391,N_2931,N_2998);
or UO_392 (O_392,N_2933,N_2941);
nor UO_393 (O_393,N_2927,N_2928);
or UO_394 (O_394,N_2991,N_2949);
and UO_395 (O_395,N_2929,N_2966);
or UO_396 (O_396,N_2939,N_2953);
nor UO_397 (O_397,N_2940,N_2984);
nor UO_398 (O_398,N_2945,N_2944);
and UO_399 (O_399,N_2985,N_2987);
and UO_400 (O_400,N_2991,N_2965);
nand UO_401 (O_401,N_2993,N_2953);
nand UO_402 (O_402,N_2938,N_2926);
nand UO_403 (O_403,N_2928,N_2938);
nor UO_404 (O_404,N_2931,N_2955);
nor UO_405 (O_405,N_2948,N_2983);
xor UO_406 (O_406,N_2943,N_2925);
and UO_407 (O_407,N_2926,N_2936);
nor UO_408 (O_408,N_2994,N_2931);
and UO_409 (O_409,N_2939,N_2989);
or UO_410 (O_410,N_2929,N_2977);
nand UO_411 (O_411,N_2980,N_2930);
xnor UO_412 (O_412,N_2987,N_2954);
or UO_413 (O_413,N_2985,N_2969);
and UO_414 (O_414,N_2960,N_2958);
and UO_415 (O_415,N_2928,N_2926);
or UO_416 (O_416,N_2927,N_2979);
nor UO_417 (O_417,N_2985,N_2971);
or UO_418 (O_418,N_2966,N_2934);
nor UO_419 (O_419,N_2965,N_2931);
or UO_420 (O_420,N_2971,N_2943);
or UO_421 (O_421,N_2936,N_2950);
nand UO_422 (O_422,N_2950,N_2940);
or UO_423 (O_423,N_2926,N_2991);
or UO_424 (O_424,N_2980,N_2935);
nor UO_425 (O_425,N_2997,N_2996);
or UO_426 (O_426,N_2925,N_2945);
nor UO_427 (O_427,N_2959,N_2995);
and UO_428 (O_428,N_2981,N_2966);
nand UO_429 (O_429,N_2994,N_2948);
nand UO_430 (O_430,N_2995,N_2958);
nand UO_431 (O_431,N_2987,N_2968);
nor UO_432 (O_432,N_2982,N_2941);
nand UO_433 (O_433,N_2946,N_2947);
and UO_434 (O_434,N_2951,N_2982);
nand UO_435 (O_435,N_2935,N_2972);
nand UO_436 (O_436,N_2991,N_2945);
nand UO_437 (O_437,N_2942,N_2985);
nor UO_438 (O_438,N_2944,N_2943);
or UO_439 (O_439,N_2973,N_2964);
nand UO_440 (O_440,N_2978,N_2988);
or UO_441 (O_441,N_2970,N_2974);
nand UO_442 (O_442,N_2952,N_2953);
and UO_443 (O_443,N_2977,N_2952);
or UO_444 (O_444,N_2972,N_2955);
nor UO_445 (O_445,N_2941,N_2937);
nor UO_446 (O_446,N_2959,N_2968);
nor UO_447 (O_447,N_2979,N_2926);
nand UO_448 (O_448,N_2946,N_2996);
nand UO_449 (O_449,N_2960,N_2977);
nor UO_450 (O_450,N_2990,N_2968);
or UO_451 (O_451,N_2964,N_2925);
or UO_452 (O_452,N_2959,N_2942);
nand UO_453 (O_453,N_2969,N_2977);
nor UO_454 (O_454,N_2942,N_2962);
nand UO_455 (O_455,N_2952,N_2967);
nand UO_456 (O_456,N_2995,N_2928);
or UO_457 (O_457,N_2946,N_2928);
and UO_458 (O_458,N_2989,N_2945);
or UO_459 (O_459,N_2929,N_2963);
nor UO_460 (O_460,N_2937,N_2994);
or UO_461 (O_461,N_2997,N_2995);
and UO_462 (O_462,N_2997,N_2929);
nor UO_463 (O_463,N_2943,N_2934);
nand UO_464 (O_464,N_2991,N_2976);
or UO_465 (O_465,N_2978,N_2936);
or UO_466 (O_466,N_2985,N_2953);
or UO_467 (O_467,N_2929,N_2947);
and UO_468 (O_468,N_2951,N_2978);
and UO_469 (O_469,N_2943,N_2964);
nor UO_470 (O_470,N_2934,N_2996);
or UO_471 (O_471,N_2938,N_2973);
nor UO_472 (O_472,N_2955,N_2977);
nor UO_473 (O_473,N_2965,N_2938);
nand UO_474 (O_474,N_2976,N_2999);
and UO_475 (O_475,N_2976,N_2945);
or UO_476 (O_476,N_2969,N_2984);
and UO_477 (O_477,N_2993,N_2988);
and UO_478 (O_478,N_2953,N_2967);
nand UO_479 (O_479,N_2965,N_2937);
and UO_480 (O_480,N_2993,N_2968);
and UO_481 (O_481,N_2994,N_2995);
or UO_482 (O_482,N_2933,N_2988);
nor UO_483 (O_483,N_2987,N_2960);
nand UO_484 (O_484,N_2926,N_2967);
nand UO_485 (O_485,N_2931,N_2976);
nand UO_486 (O_486,N_2932,N_2974);
nor UO_487 (O_487,N_2990,N_2981);
nand UO_488 (O_488,N_2962,N_2977);
and UO_489 (O_489,N_2987,N_2943);
or UO_490 (O_490,N_2988,N_2973);
nor UO_491 (O_491,N_2964,N_2996);
nor UO_492 (O_492,N_2976,N_2960);
nand UO_493 (O_493,N_2977,N_2990);
and UO_494 (O_494,N_2945,N_2957);
or UO_495 (O_495,N_2937,N_2982);
nor UO_496 (O_496,N_2988,N_2951);
or UO_497 (O_497,N_2962,N_2971);
nand UO_498 (O_498,N_2986,N_2954);
and UO_499 (O_499,N_2958,N_2985);
endmodule