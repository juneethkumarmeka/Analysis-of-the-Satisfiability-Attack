module basic_1000_10000_1500_2_levels_10xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5002,N_5006,N_5009,N_5010,N_5011,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5023,N_5024,N_5026,N_5027,N_5028,N_5029,N_5032,N_5033,N_5035,N_5036,N_5039,N_5040,N_5041,N_5042,N_5044,N_5046,N_5047,N_5048,N_5052,N_5053,N_5057,N_5060,N_5061,N_5063,N_5064,N_5065,N_5066,N_5068,N_5069,N_5070,N_5071,N_5072,N_5077,N_5078,N_5084,N_5086,N_5088,N_5091,N_5092,N_5094,N_5096,N_5100,N_5102,N_5104,N_5105,N_5106,N_5110,N_5111,N_5113,N_5115,N_5118,N_5119,N_5121,N_5122,N_5123,N_5124,N_5125,N_5131,N_5134,N_5136,N_5137,N_5140,N_5141,N_5142,N_5144,N_5145,N_5146,N_5148,N_5150,N_5151,N_5152,N_5153,N_5155,N_5157,N_5159,N_5160,N_5161,N_5163,N_5167,N_5171,N_5175,N_5176,N_5178,N_5179,N_5180,N_5181,N_5182,N_5186,N_5188,N_5189,N_5195,N_5196,N_5197,N_5200,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5213,N_5214,N_5215,N_5217,N_5218,N_5220,N_5224,N_5225,N_5227,N_5228,N_5230,N_5231,N_5232,N_5237,N_5238,N_5240,N_5242,N_5243,N_5244,N_5245,N_5248,N_5249,N_5250,N_5252,N_5254,N_5255,N_5258,N_5259,N_5260,N_5261,N_5263,N_5264,N_5265,N_5267,N_5270,N_5271,N_5272,N_5274,N_5281,N_5283,N_5286,N_5287,N_5288,N_5289,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5300,N_5304,N_5306,N_5310,N_5311,N_5315,N_5317,N_5318,N_5321,N_5322,N_5323,N_5325,N_5326,N_5327,N_5328,N_5330,N_5331,N_5333,N_5335,N_5336,N_5338,N_5340,N_5341,N_5342,N_5343,N_5345,N_5346,N_5347,N_5348,N_5352,N_5354,N_5355,N_5357,N_5358,N_5360,N_5361,N_5363,N_5364,N_5366,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5375,N_5376,N_5379,N_5380,N_5381,N_5383,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5400,N_5403,N_5406,N_5407,N_5408,N_5409,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5418,N_5419,N_5420,N_5423,N_5425,N_5426,N_5429,N_5432,N_5437,N_5440,N_5443,N_5446,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5456,N_5458,N_5459,N_5461,N_5464,N_5465,N_5466,N_5467,N_5470,N_5473,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5482,N_5483,N_5485,N_5487,N_5491,N_5492,N_5494,N_5495,N_5496,N_5498,N_5499,N_5500,N_5502,N_5505,N_5506,N_5509,N_5510,N_5511,N_5512,N_5515,N_5516,N_5517,N_5521,N_5522,N_5524,N_5528,N_5529,N_5531,N_5533,N_5534,N_5535,N_5540,N_5541,N_5542,N_5543,N_5544,N_5549,N_5551,N_5553,N_5555,N_5556,N_5558,N_5562,N_5564,N_5566,N_5567,N_5569,N_5570,N_5571,N_5572,N_5575,N_5576,N_5578,N_5580,N_5581,N_5582,N_5584,N_5587,N_5593,N_5594,N_5595,N_5596,N_5603,N_5605,N_5606,N_5607,N_5609,N_5612,N_5614,N_5615,N_5616,N_5617,N_5620,N_5621,N_5622,N_5623,N_5625,N_5626,N_5627,N_5629,N_5632,N_5635,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5645,N_5646,N_5648,N_5649,N_5650,N_5651,N_5653,N_5654,N_5655,N_5656,N_5658,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5668,N_5669,N_5671,N_5672,N_5673,N_5674,N_5675,N_5677,N_5678,N_5685,N_5686,N_5687,N_5688,N_5690,N_5691,N_5693,N_5694,N_5695,N_5696,N_5699,N_5701,N_5703,N_5706,N_5707,N_5708,N_5710,N_5715,N_5716,N_5720,N_5722,N_5725,N_5726,N_5727,N_5730,N_5733,N_5736,N_5737,N_5740,N_5742,N_5746,N_5748,N_5749,N_5750,N_5754,N_5758,N_5759,N_5760,N_5762,N_5765,N_5767,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5782,N_5783,N_5784,N_5786,N_5788,N_5791,N_5793,N_5795,N_5796,N_5797,N_5798,N_5800,N_5802,N_5804,N_5805,N_5807,N_5808,N_5809,N_5810,N_5812,N_5813,N_5814,N_5817,N_5819,N_5820,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5831,N_5832,N_5834,N_5835,N_5837,N_5838,N_5839,N_5840,N_5841,N_5844,N_5846,N_5848,N_5849,N_5850,N_5851,N_5852,N_5854,N_5855,N_5856,N_5857,N_5859,N_5862,N_5863,N_5865,N_5866,N_5868,N_5869,N_5870,N_5871,N_5872,N_5874,N_5875,N_5876,N_5877,N_5878,N_5883,N_5886,N_5887,N_5888,N_5889,N_5890,N_5892,N_5893,N_5899,N_5900,N_5903,N_5904,N_5906,N_5907,N_5910,N_5911,N_5912,N_5914,N_5915,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5926,N_5928,N_5932,N_5934,N_5935,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5946,N_5947,N_5950,N_5953,N_5954,N_5956,N_5958,N_5961,N_5963,N_5965,N_5966,N_5967,N_5969,N_5971,N_5972,N_5973,N_5976,N_5977,N_5978,N_5979,N_5980,N_5982,N_5985,N_5986,N_5990,N_5992,N_5993,N_5994,N_5995,N_5998,N_6000,N_6001,N_6002,N_6006,N_6007,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6017,N_6018,N_6019,N_6020,N_6021,N_6023,N_6024,N_6025,N_6028,N_6029,N_6030,N_6031,N_6032,N_6035,N_6036,N_6038,N_6040,N_6041,N_6042,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6072,N_6073,N_6074,N_6076,N_6078,N_6079,N_6081,N_6082,N_6084,N_6089,N_6090,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6103,N_6105,N_6108,N_6109,N_6112,N_6114,N_6116,N_6117,N_6118,N_6119,N_6122,N_6125,N_6126,N_6127,N_6130,N_6131,N_6133,N_6134,N_6136,N_6138,N_6139,N_6141,N_6142,N_6143,N_6144,N_6145,N_6147,N_6148,N_6149,N_6150,N_6153,N_6154,N_6159,N_6161,N_6162,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6176,N_6177,N_6178,N_6180,N_6182,N_6185,N_6187,N_6188,N_6189,N_6190,N_6191,N_6193,N_6194,N_6196,N_6197,N_6199,N_6200,N_6201,N_6202,N_6209,N_6210,N_6212,N_6213,N_6217,N_6218,N_6219,N_6220,N_6222,N_6224,N_6225,N_6226,N_6227,N_6229,N_6233,N_6235,N_6236,N_6239,N_6240,N_6241,N_6243,N_6248,N_6252,N_6255,N_6257,N_6258,N_6259,N_6261,N_6262,N_6263,N_6264,N_6265,N_6267,N_6270,N_6271,N_6272,N_6273,N_6274,N_6276,N_6277,N_6278,N_6281,N_6282,N_6284,N_6285,N_6286,N_6287,N_6288,N_6290,N_6291,N_6293,N_6296,N_6298,N_6299,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6311,N_6313,N_6314,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6325,N_6326,N_6328,N_6330,N_6331,N_6332,N_6333,N_6335,N_6336,N_6337,N_6340,N_6341,N_6343,N_6344,N_6347,N_6348,N_6349,N_6350,N_6351,N_6353,N_6354,N_6355,N_6357,N_6358,N_6360,N_6361,N_6366,N_6367,N_6369,N_6370,N_6371,N_6373,N_6375,N_6376,N_6378,N_6379,N_6380,N_6383,N_6384,N_6386,N_6387,N_6388,N_6389,N_6392,N_6395,N_6400,N_6401,N_6407,N_6409,N_6411,N_6412,N_6413,N_6414,N_6416,N_6418,N_6419,N_6423,N_6424,N_6425,N_6426,N_6427,N_6429,N_6430,N_6431,N_6435,N_6436,N_6438,N_6441,N_6442,N_6445,N_6446,N_6447,N_6449,N_6450,N_6451,N_6452,N_6453,N_6456,N_6458,N_6460,N_6461,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6470,N_6472,N_6474,N_6475,N_6476,N_6477,N_6480,N_6481,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6492,N_6494,N_6495,N_6497,N_6498,N_6500,N_6502,N_6505,N_6506,N_6510,N_6512,N_6517,N_6518,N_6520,N_6521,N_6522,N_6523,N_6524,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6537,N_6538,N_6539,N_6540,N_6541,N_6543,N_6546,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6557,N_6558,N_6559,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6573,N_6575,N_6577,N_6579,N_6584,N_6585,N_6586,N_6587,N_6588,N_6591,N_6592,N_6593,N_6599,N_6603,N_6604,N_6609,N_6610,N_6612,N_6613,N_6615,N_6616,N_6617,N_6618,N_6619,N_6621,N_6622,N_6623,N_6624,N_6625,N_6627,N_6628,N_6629,N_6632,N_6638,N_6639,N_6640,N_6642,N_6643,N_6644,N_6646,N_6647,N_6649,N_6653,N_6654,N_6655,N_6657,N_6658,N_6659,N_6661,N_6665,N_6667,N_6668,N_6669,N_6671,N_6672,N_6674,N_6675,N_6676,N_6677,N_6678,N_6680,N_6682,N_6683,N_6684,N_6685,N_6686,N_6688,N_6691,N_6693,N_6698,N_6701,N_6703,N_6705,N_6706,N_6711,N_6712,N_6714,N_6715,N_6717,N_6719,N_6720,N_6723,N_6727,N_6728,N_6729,N_6730,N_6731,N_6734,N_6737,N_6738,N_6739,N_6744,N_6745,N_6750,N_6751,N_6752,N_6754,N_6755,N_6756,N_6757,N_6759,N_6761,N_6763,N_6764,N_6765,N_6767,N_6769,N_6770,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6781,N_6782,N_6783,N_6785,N_6786,N_6788,N_6792,N_6793,N_6794,N_6795,N_6796,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6806,N_6808,N_6812,N_6813,N_6814,N_6815,N_6816,N_6819,N_6820,N_6821,N_6823,N_6824,N_6826,N_6827,N_6828,N_6829,N_6831,N_6833,N_6835,N_6836,N_6837,N_6838,N_6841,N_6842,N_6843,N_6847,N_6849,N_6850,N_6851,N_6855,N_6858,N_6859,N_6860,N_6862,N_6863,N_6865,N_6866,N_6867,N_6873,N_6874,N_6875,N_6876,N_6878,N_6879,N_6880,N_6881,N_6883,N_6885,N_6886,N_6888,N_6889,N_6890,N_6892,N_6893,N_6895,N_6901,N_6902,N_6904,N_6907,N_6909,N_6910,N_6912,N_6913,N_6915,N_6916,N_6918,N_6919,N_6920,N_6922,N_6923,N_6924,N_6927,N_6928,N_6931,N_6932,N_6933,N_6936,N_6937,N_6938,N_6941,N_6942,N_6945,N_6948,N_6949,N_6950,N_6952,N_6954,N_6955,N_6957,N_6958,N_6959,N_6960,N_6961,N_6963,N_6964,N_6968,N_6970,N_6971,N_6972,N_6973,N_6975,N_6976,N_6977,N_6980,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6995,N_6997,N_6999,N_7000,N_7002,N_7004,N_7005,N_7006,N_7007,N_7009,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7020,N_7021,N_7022,N_7025,N_7027,N_7028,N_7031,N_7033,N_7035,N_7036,N_7037,N_7038,N_7040,N_7044,N_7046,N_7048,N_7050,N_7051,N_7053,N_7054,N_7055,N_7056,N_7057,N_7059,N_7060,N_7062,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7091,N_7092,N_7094,N_7095,N_7098,N_7100,N_7101,N_7102,N_7103,N_7104,N_7106,N_7108,N_7109,N_7115,N_7117,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7132,N_7134,N_7135,N_7136,N_7138,N_7139,N_7140,N_7142,N_7143,N_7145,N_7146,N_7147,N_7148,N_7150,N_7151,N_7154,N_7156,N_7157,N_7158,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7168,N_7169,N_7171,N_7172,N_7176,N_7177,N_7178,N_7180,N_7181,N_7184,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7194,N_7195,N_7197,N_7203,N_7204,N_7205,N_7207,N_7209,N_7210,N_7213,N_7214,N_7215,N_7217,N_7218,N_7223,N_7225,N_7226,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7248,N_7250,N_7252,N_7253,N_7254,N_7255,N_7256,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7269,N_7270,N_7271,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7284,N_7285,N_7290,N_7291,N_7295,N_7296,N_7297,N_7300,N_7302,N_7304,N_7305,N_7307,N_7308,N_7309,N_7310,N_7314,N_7316,N_7318,N_7320,N_7321,N_7322,N_7323,N_7324,N_7327,N_7328,N_7335,N_7337,N_7338,N_7339,N_7341,N_7343,N_7345,N_7346,N_7347,N_7348,N_7350,N_7351,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7360,N_7361,N_7363,N_7367,N_7368,N_7370,N_7373,N_7374,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7385,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7398,N_7399,N_7400,N_7404,N_7408,N_7413,N_7414,N_7415,N_7416,N_7418,N_7419,N_7420,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7442,N_7443,N_7445,N_7446,N_7449,N_7451,N_7452,N_7454,N_7456,N_7457,N_7459,N_7460,N_7462,N_7464,N_7465,N_7470,N_7471,N_7474,N_7475,N_7481,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7491,N_7492,N_7494,N_7495,N_7496,N_7497,N_7500,N_7501,N_7502,N_7504,N_7505,N_7506,N_7507,N_7508,N_7510,N_7514,N_7515,N_7517,N_7518,N_7520,N_7522,N_7523,N_7524,N_7526,N_7528,N_7529,N_7530,N_7532,N_7533,N_7534,N_7535,N_7536,N_7538,N_7539,N_7540,N_7541,N_7543,N_7544,N_7545,N_7546,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7565,N_7567,N_7568,N_7573,N_7574,N_7575,N_7576,N_7578,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7587,N_7588,N_7592,N_7593,N_7595,N_7598,N_7600,N_7601,N_7602,N_7604,N_7605,N_7608,N_7609,N_7611,N_7615,N_7616,N_7618,N_7622,N_7625,N_7628,N_7631,N_7633,N_7634,N_7637,N_7639,N_7641,N_7642,N_7643,N_7644,N_7647,N_7649,N_7651,N_7652,N_7654,N_7655,N_7656,N_7657,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7671,N_7673,N_7674,N_7676,N_7677,N_7679,N_7680,N_7682,N_7684,N_7685,N_7686,N_7689,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7700,N_7703,N_7704,N_7705,N_7706,N_7707,N_7709,N_7710,N_7713,N_7714,N_7715,N_7716,N_7717,N_7720,N_7721,N_7722,N_7723,N_7725,N_7728,N_7729,N_7731,N_7732,N_7741,N_7743,N_7746,N_7748,N_7749,N_7750,N_7753,N_7755,N_7756,N_7757,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7772,N_7773,N_7774,N_7775,N_7777,N_7779,N_7780,N_7783,N_7784,N_7785,N_7787,N_7789,N_7790,N_7793,N_7795,N_7799,N_7800,N_7802,N_7804,N_7808,N_7809,N_7810,N_7811,N_7813,N_7814,N_7815,N_7817,N_7819,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7829,N_7831,N_7833,N_7834,N_7835,N_7837,N_7838,N_7839,N_7840,N_7843,N_7844,N_7849,N_7850,N_7853,N_7854,N_7855,N_7856,N_7858,N_7859,N_7861,N_7862,N_7864,N_7865,N_7871,N_7872,N_7876,N_7877,N_7878,N_7881,N_7882,N_7883,N_7885,N_7887,N_7889,N_7890,N_7892,N_7894,N_7897,N_7898,N_7899,N_7907,N_7908,N_7909,N_7913,N_7915,N_7917,N_7918,N_7919,N_7920,N_7922,N_7925,N_7928,N_7929,N_7930,N_7934,N_7935,N_7936,N_7938,N_7940,N_7941,N_7943,N_7944,N_7946,N_7950,N_7951,N_7952,N_7955,N_7958,N_7959,N_7961,N_7963,N_7966,N_7971,N_7975,N_7976,N_7978,N_7979,N_7981,N_7982,N_7983,N_7984,N_7985,N_7990,N_7991,N_7994,N_7995,N_7997,N_7998,N_8002,N_8005,N_8006,N_8007,N_8009,N_8010,N_8012,N_8013,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8025,N_8026,N_8027,N_8029,N_8030,N_8032,N_8036,N_8037,N_8038,N_8039,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8053,N_8054,N_8055,N_8057,N_8058,N_8059,N_8060,N_8062,N_8063,N_8064,N_8066,N_8068,N_8069,N_8070,N_8072,N_8074,N_8078,N_8082,N_8083,N_8085,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8096,N_8097,N_8099,N_8101,N_8102,N_8104,N_8106,N_8108,N_8111,N_8113,N_8115,N_8116,N_8117,N_8118,N_8119,N_8121,N_8122,N_8124,N_8125,N_8126,N_8128,N_8130,N_8131,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8145,N_8147,N_8149,N_8151,N_8152,N_8153,N_8156,N_8157,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8170,N_8171,N_8172,N_8173,N_8174,N_8177,N_8178,N_8181,N_8182,N_8183,N_8186,N_8187,N_8189,N_8192,N_8195,N_8198,N_8199,N_8200,N_8201,N_8203,N_8205,N_8209,N_8210,N_8218,N_8220,N_8222,N_8223,N_8224,N_8225,N_8227,N_8229,N_8231,N_8232,N_8233,N_8234,N_8235,N_8237,N_8239,N_8240,N_8242,N_8243,N_8244,N_8248,N_8249,N_8250,N_8251,N_8252,N_8254,N_8255,N_8257,N_8261,N_8264,N_8265,N_8266,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8275,N_8276,N_8278,N_8281,N_8283,N_8285,N_8287,N_8288,N_8291,N_8294,N_8297,N_8298,N_8300,N_8301,N_8302,N_8305,N_8306,N_8307,N_8309,N_8313,N_8315,N_8316,N_8318,N_8321,N_8323,N_8324,N_8325,N_8326,N_8328,N_8332,N_8333,N_8334,N_8335,N_8337,N_8338,N_8339,N_8340,N_8342,N_8344,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8353,N_8354,N_8355,N_8357,N_8358,N_8359,N_8363,N_8364,N_8365,N_8366,N_8368,N_8369,N_8370,N_8372,N_8373,N_8374,N_8376,N_8377,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8387,N_8389,N_8392,N_8395,N_8396,N_8397,N_8399,N_8402,N_8404,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8414,N_8415,N_8416,N_8419,N_8421,N_8425,N_8428,N_8429,N_8430,N_8431,N_8436,N_8439,N_8440,N_8441,N_8443,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8454,N_8456,N_8459,N_8460,N_8461,N_8462,N_8463,N_8465,N_8466,N_8467,N_8469,N_8470,N_8471,N_8472,N_8473,N_8475,N_8476,N_8477,N_8479,N_8480,N_8481,N_8482,N_8489,N_8490,N_8491,N_8492,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8502,N_8503,N_8504,N_8505,N_8507,N_8508,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8517,N_8518,N_8520,N_8522,N_8524,N_8526,N_8527,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8540,N_8541,N_8544,N_8546,N_8547,N_8548,N_8549,N_8551,N_8552,N_8553,N_8555,N_8556,N_8557,N_8558,N_8561,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8573,N_8575,N_8576,N_8578,N_8579,N_8581,N_8582,N_8583,N_8587,N_8588,N_8591,N_8592,N_8593,N_8596,N_8597,N_8599,N_8600,N_8601,N_8602,N_8604,N_8606,N_8607,N_8609,N_8611,N_8612,N_8613,N_8615,N_8619,N_8620,N_8621,N_8623,N_8625,N_8627,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8637,N_8640,N_8641,N_8643,N_8644,N_8645,N_8647,N_8648,N_8651,N_8653,N_8656,N_8658,N_8659,N_8660,N_8662,N_8663,N_8666,N_8668,N_8671,N_8672,N_8673,N_8674,N_8675,N_8678,N_8681,N_8683,N_8685,N_8686,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8702,N_8703,N_8705,N_8708,N_8709,N_8710,N_8711,N_8712,N_8714,N_8716,N_8718,N_8719,N_8721,N_8722,N_8723,N_8725,N_8726,N_8727,N_8729,N_8731,N_8732,N_8735,N_8736,N_8737,N_8742,N_8743,N_8745,N_8746,N_8749,N_8750,N_8751,N_8752,N_8753,N_8758,N_8759,N_8760,N_8762,N_8763,N_8764,N_8765,N_8766,N_8768,N_8770,N_8771,N_8772,N_8773,N_8775,N_8776,N_8777,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8788,N_8789,N_8791,N_8792,N_8794,N_8795,N_8797,N_8799,N_8803,N_8804,N_8806,N_8809,N_8810,N_8811,N_8813,N_8815,N_8817,N_8819,N_8821,N_8822,N_8823,N_8824,N_8826,N_8827,N_8828,N_8830,N_8831,N_8832,N_8836,N_8839,N_8842,N_8843,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8857,N_8858,N_8859,N_8861,N_8862,N_8863,N_8864,N_8865,N_8872,N_8873,N_8874,N_8876,N_8877,N_8879,N_8881,N_8883,N_8884,N_8887,N_8889,N_8890,N_8893,N_8896,N_8898,N_8899,N_8901,N_8903,N_8904,N_8907,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8925,N_8926,N_8928,N_8929,N_8930,N_8933,N_8941,N_8942,N_8944,N_8946,N_8947,N_8948,N_8949,N_8951,N_8953,N_8957,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8975,N_8976,N_8977,N_8979,N_8980,N_8981,N_8983,N_8984,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8998,N_8999,N_9000,N_9001,N_9002,N_9004,N_9005,N_9006,N_9008,N_9009,N_9010,N_9011,N_9012,N_9014,N_9015,N_9016,N_9022,N_9023,N_9024,N_9026,N_9027,N_9031,N_9032,N_9033,N_9034,N_9035,N_9038,N_9040,N_9041,N_9042,N_9043,N_9045,N_9046,N_9047,N_9050,N_9052,N_9053,N_9055,N_9056,N_9058,N_9060,N_9061,N_9062,N_9069,N_9070,N_9073,N_9075,N_9076,N_9077,N_9078,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9088,N_9090,N_9091,N_9092,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9105,N_9106,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9116,N_9117,N_9118,N_9119,N_9121,N_9122,N_9123,N_9124,N_9125,N_9127,N_9129,N_9130,N_9131,N_9135,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9144,N_9145,N_9146,N_9147,N_9148,N_9150,N_9152,N_9153,N_9154,N_9155,N_9157,N_9158,N_9160,N_9167,N_9168,N_9169,N_9170,N_9174,N_9176,N_9177,N_9178,N_9179,N_9181,N_9183,N_9184,N_9186,N_9187,N_9189,N_9190,N_9191,N_9192,N_9195,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9212,N_9216,N_9217,N_9219,N_9221,N_9222,N_9225,N_9226,N_9227,N_9229,N_9230,N_9231,N_9233,N_9234,N_9235,N_9236,N_9238,N_9240,N_9243,N_9244,N_9245,N_9247,N_9249,N_9253,N_9255,N_9256,N_9258,N_9260,N_9262,N_9264,N_9266,N_9268,N_9269,N_9270,N_9272,N_9273,N_9274,N_9275,N_9276,N_9278,N_9280,N_9281,N_9284,N_9285,N_9287,N_9288,N_9289,N_9290,N_9291,N_9293,N_9294,N_9295,N_9296,N_9299,N_9300,N_9301,N_9303,N_9304,N_9306,N_9309,N_9311,N_9312,N_9314,N_9316,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9331,N_9332,N_9334,N_9335,N_9336,N_9337,N_9340,N_9341,N_9342,N_9343,N_9345,N_9347,N_9349,N_9352,N_9355,N_9356,N_9357,N_9359,N_9360,N_9361,N_9362,N_9363,N_9365,N_9368,N_9369,N_9371,N_9372,N_9374,N_9375,N_9376,N_9378,N_9381,N_9382,N_9384,N_9385,N_9388,N_9392,N_9394,N_9396,N_9398,N_9399,N_9400,N_9401,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9411,N_9412,N_9415,N_9416,N_9418,N_9420,N_9421,N_9423,N_9425,N_9427,N_9429,N_9431,N_9432,N_9433,N_9434,N_9436,N_9437,N_9439,N_9445,N_9451,N_9452,N_9453,N_9454,N_9456,N_9458,N_9459,N_9460,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9474,N_9475,N_9477,N_9478,N_9481,N_9483,N_9484,N_9487,N_9488,N_9490,N_9493,N_9494,N_9495,N_9496,N_9497,N_9499,N_9500,N_9502,N_9504,N_9505,N_9506,N_9507,N_9509,N_9511,N_9512,N_9514,N_9515,N_9516,N_9518,N_9519,N_9523,N_9525,N_9527,N_9528,N_9529,N_9530,N_9533,N_9535,N_9536,N_9537,N_9538,N_9539,N_9547,N_9548,N_9549,N_9552,N_9554,N_9556,N_9560,N_9561,N_9565,N_9566,N_9569,N_9570,N_9573,N_9574,N_9575,N_9577,N_9578,N_9579,N_9580,N_9581,N_9583,N_9584,N_9585,N_9586,N_9587,N_9590,N_9591,N_9593,N_9596,N_9597,N_9598,N_9601,N_9602,N_9603,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9615,N_9617,N_9619,N_9623,N_9625,N_9626,N_9627,N_9628,N_9629,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9638,N_9639,N_9640,N_9641,N_9642,N_9647,N_9648,N_9649,N_9655,N_9656,N_9658,N_9659,N_9660,N_9665,N_9666,N_9667,N_9668,N_9669,N_9671,N_9673,N_9674,N_9675,N_9676,N_9678,N_9679,N_9681,N_9685,N_9686,N_9688,N_9689,N_9690,N_9691,N_9692,N_9695,N_9697,N_9698,N_9701,N_9702,N_9703,N_9704,N_9705,N_9707,N_9708,N_9710,N_9716,N_9719,N_9720,N_9724,N_9725,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9736,N_9739,N_9740,N_9741,N_9743,N_9745,N_9748,N_9749,N_9750,N_9753,N_9755,N_9757,N_9758,N_9760,N_9762,N_9763,N_9766,N_9769,N_9770,N_9775,N_9777,N_9781,N_9782,N_9786,N_9787,N_9788,N_9792,N_9793,N_9795,N_9796,N_9797,N_9798,N_9799,N_9802,N_9803,N_9805,N_9807,N_9810,N_9811,N_9814,N_9816,N_9817,N_9821,N_9824,N_9825,N_9827,N_9828,N_9832,N_9833,N_9834,N_9837,N_9840,N_9841,N_9844,N_9845,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9858,N_9859,N_9861,N_9866,N_9867,N_9868,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9879,N_9884,N_9885,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9895,N_9896,N_9897,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9907,N_9908,N_9910,N_9912,N_9915,N_9917,N_9919,N_9920,N_9922,N_9924,N_9926,N_9927,N_9928,N_9930,N_9931,N_9932,N_9934,N_9937,N_9938,N_9940,N_9945,N_9947,N_9949,N_9950,N_9951,N_9953,N_9959,N_9962,N_9963,N_9964,N_9966,N_9967,N_9970,N_9971,N_9974,N_9975,N_9976,N_9977,N_9978,N_9983,N_9984,N_9986,N_9989,N_9990,N_9991,N_9994,N_9995,N_9996,N_9998;
nand U0 (N_0,In_112,In_214);
or U1 (N_1,In_456,In_275);
xor U2 (N_2,In_607,In_406);
nor U3 (N_3,In_647,In_658);
nand U4 (N_4,In_762,In_369);
or U5 (N_5,In_128,In_978);
xor U6 (N_6,In_713,In_543);
nand U7 (N_7,In_17,In_56);
xor U8 (N_8,In_157,In_315);
or U9 (N_9,In_969,In_907);
and U10 (N_10,In_160,In_480);
nor U11 (N_11,In_866,In_2);
or U12 (N_12,In_858,In_224);
and U13 (N_13,In_876,In_131);
nand U14 (N_14,In_80,In_21);
or U15 (N_15,In_494,In_91);
nand U16 (N_16,In_405,In_190);
and U17 (N_17,In_634,In_878);
nor U18 (N_18,In_362,In_443);
xnor U19 (N_19,In_587,In_371);
nor U20 (N_20,In_152,In_423);
or U21 (N_21,In_95,In_759);
xnor U22 (N_22,In_243,In_548);
nor U23 (N_23,In_886,In_798);
nand U24 (N_24,In_918,In_835);
nor U25 (N_25,In_301,In_189);
and U26 (N_26,In_603,In_339);
and U27 (N_27,In_495,In_983);
nand U28 (N_28,In_779,In_106);
nand U29 (N_29,In_240,In_967);
nand U30 (N_30,In_428,In_807);
nand U31 (N_31,In_816,In_242);
nand U32 (N_32,In_879,In_192);
or U33 (N_33,In_533,In_864);
or U34 (N_34,In_414,In_757);
and U35 (N_35,In_552,In_20);
and U36 (N_36,In_280,In_733);
nor U37 (N_37,In_582,In_684);
and U38 (N_38,In_183,In_248);
nor U39 (N_39,In_953,In_149);
or U40 (N_40,In_86,In_295);
nor U41 (N_41,In_806,In_900);
xor U42 (N_42,In_588,In_792);
nand U43 (N_43,In_674,In_343);
xnor U44 (N_44,In_468,In_155);
xnor U45 (N_45,In_635,In_67);
xor U46 (N_46,In_83,In_44);
xnor U47 (N_47,In_450,In_624);
nor U48 (N_48,In_466,In_58);
nand U49 (N_49,In_230,In_204);
and U50 (N_50,In_659,In_167);
or U51 (N_51,In_312,In_935);
nand U52 (N_52,In_591,In_769);
nor U53 (N_53,In_293,In_620);
nor U54 (N_54,In_619,In_368);
or U55 (N_55,In_887,In_997);
nor U56 (N_56,In_42,In_531);
and U57 (N_57,In_170,In_814);
nand U58 (N_58,In_576,In_891);
nand U59 (N_59,In_114,In_228);
nor U60 (N_60,In_258,In_926);
nor U61 (N_61,In_453,In_309);
or U62 (N_62,In_393,In_968);
and U63 (N_63,In_925,In_89);
xnor U64 (N_64,In_458,In_193);
or U65 (N_65,In_986,In_874);
or U66 (N_66,In_827,In_566);
and U67 (N_67,In_246,In_344);
nand U68 (N_68,In_46,In_294);
nor U69 (N_69,In_300,In_679);
and U70 (N_70,In_132,In_52);
and U71 (N_71,In_562,In_783);
nor U72 (N_72,In_179,In_854);
nand U73 (N_73,In_174,In_14);
nor U74 (N_74,In_310,In_743);
or U75 (N_75,In_688,In_475);
nor U76 (N_76,In_868,In_387);
or U77 (N_77,In_751,In_556);
xor U78 (N_78,In_830,In_216);
nor U79 (N_79,In_436,In_119);
nor U80 (N_80,In_286,In_832);
and U81 (N_81,In_937,In_943);
and U82 (N_82,In_687,In_270);
or U83 (N_83,In_561,In_860);
nor U84 (N_84,In_485,In_66);
xnor U85 (N_85,In_975,In_580);
or U86 (N_86,In_991,In_723);
nand U87 (N_87,In_559,In_675);
or U88 (N_88,In_784,In_261);
nor U89 (N_89,In_927,In_319);
or U90 (N_90,In_626,In_734);
and U91 (N_91,In_715,In_172);
nand U92 (N_92,In_32,In_717);
or U93 (N_93,In_802,In_249);
nand U94 (N_94,In_316,In_471);
and U95 (N_95,In_856,In_19);
nand U96 (N_96,In_716,In_277);
nand U97 (N_97,In_867,In_841);
or U98 (N_98,In_245,In_694);
xnor U99 (N_99,In_60,In_585);
nor U100 (N_100,In_911,In_53);
nand U101 (N_101,In_262,In_373);
nor U102 (N_102,In_822,In_180);
nand U103 (N_103,In_442,In_460);
or U104 (N_104,In_98,In_434);
nor U105 (N_105,In_699,In_695);
nand U106 (N_106,In_944,In_411);
or U107 (N_107,In_643,In_993);
nor U108 (N_108,In_962,In_354);
or U109 (N_109,In_45,In_178);
nand U110 (N_110,In_903,In_211);
nand U111 (N_111,In_998,In_218);
nor U112 (N_112,In_209,In_398);
or U113 (N_113,In_296,In_483);
or U114 (N_114,In_74,In_308);
nor U115 (N_115,In_516,In_313);
and U116 (N_116,In_375,In_191);
nor U117 (N_117,In_614,In_124);
xnor U118 (N_118,In_642,In_645);
nand U119 (N_119,In_419,In_196);
nand U120 (N_120,In_959,In_142);
and U121 (N_121,In_578,In_696);
nand U122 (N_122,In_284,In_401);
nand U123 (N_123,In_96,In_622);
nand U124 (N_124,In_115,In_589);
and U125 (N_125,In_444,In_523);
xor U126 (N_126,In_996,In_438);
and U127 (N_127,In_956,In_256);
xnor U128 (N_128,In_502,In_794);
xnor U129 (N_129,In_730,In_655);
xnor U130 (N_130,In_71,In_150);
nor U131 (N_131,In_754,In_768);
xnor U132 (N_132,In_415,In_667);
or U133 (N_133,In_791,In_636);
nor U134 (N_134,In_666,In_109);
nand U135 (N_135,In_527,In_338);
and U136 (N_136,In_11,In_726);
or U137 (N_137,In_382,In_662);
nor U138 (N_138,In_464,In_36);
and U139 (N_139,In_676,In_951);
xnor U140 (N_140,In_708,In_611);
xnor U141 (N_141,In_113,In_568);
nor U142 (N_142,In_93,In_892);
or U143 (N_143,In_722,In_283);
or U144 (N_144,In_473,In_704);
and U145 (N_145,In_452,In_459);
nor U146 (N_146,In_62,In_197);
nor U147 (N_147,In_347,In_542);
or U148 (N_148,In_328,In_989);
xnor U149 (N_149,In_223,In_537);
or U150 (N_150,In_522,In_73);
xnor U151 (N_151,In_893,In_187);
nand U152 (N_152,In_805,In_839);
or U153 (N_153,In_593,In_381);
or U154 (N_154,In_644,In_970);
and U155 (N_155,In_532,In_517);
nand U156 (N_156,In_208,In_306);
xor U157 (N_157,In_597,In_365);
nand U158 (N_158,In_166,In_933);
or U159 (N_159,In_273,In_302);
xnor U160 (N_160,In_212,In_184);
nor U161 (N_161,In_916,In_432);
nor U162 (N_162,In_952,In_617);
nand U163 (N_163,In_749,In_333);
nand U164 (N_164,In_169,In_233);
nand U165 (N_165,In_311,In_815);
or U166 (N_166,In_318,In_143);
xnor U167 (N_167,In_549,In_28);
nor U168 (N_168,In_496,In_345);
nand U169 (N_169,In_427,In_917);
nor U170 (N_170,In_278,In_287);
xor U171 (N_171,In_263,In_595);
and U172 (N_172,In_239,In_380);
or U173 (N_173,In_984,In_747);
nor U174 (N_174,In_241,In_819);
and U175 (N_175,In_817,In_631);
xnor U176 (N_176,In_946,In_812);
and U177 (N_177,In_663,In_140);
xnor U178 (N_178,In_162,In_221);
nor U179 (N_179,In_325,In_99);
and U180 (N_180,In_481,In_253);
or U181 (N_181,In_870,In_513);
and U182 (N_182,In_244,In_22);
xnor U183 (N_183,In_748,In_857);
nor U184 (N_184,In_225,In_650);
and U185 (N_185,In_147,In_837);
nor U186 (N_186,In_350,In_890);
or U187 (N_187,In_669,In_487);
nand U188 (N_188,In_441,In_729);
or U189 (N_189,In_521,In_863);
nor U190 (N_190,In_340,In_418);
or U191 (N_191,In_520,In_236);
or U192 (N_192,In_711,In_201);
or U193 (N_193,In_950,In_3);
and U194 (N_194,In_331,In_888);
xnor U195 (N_195,In_508,In_506);
and U196 (N_196,In_269,In_709);
nor U197 (N_197,In_665,In_102);
nand U198 (N_198,In_596,In_755);
nand U199 (N_199,In_810,In_247);
and U200 (N_200,In_871,In_898);
nor U201 (N_201,In_629,In_175);
or U202 (N_202,In_202,In_292);
xnor U203 (N_203,In_281,In_107);
nor U204 (N_204,In_939,In_195);
or U205 (N_205,In_116,In_842);
xor U206 (N_206,In_721,In_500);
and U207 (N_207,In_601,In_237);
nor U208 (N_208,In_648,In_605);
or U209 (N_209,In_905,In_198);
or U210 (N_210,In_31,In_422);
nor U211 (N_211,In_100,In_425);
nand U212 (N_212,In_942,In_744);
nand U213 (N_213,In_793,In_484);
nand U214 (N_214,In_999,In_24);
nor U215 (N_215,In_901,In_367);
nand U216 (N_216,In_719,In_510);
and U217 (N_217,In_971,In_586);
nand U218 (N_218,In_811,In_206);
and U219 (N_219,In_376,In_266);
and U220 (N_220,In_320,In_440);
xor U221 (N_221,In_104,In_606);
nand U222 (N_222,In_564,In_35);
xnor U223 (N_223,In_923,In_492);
or U224 (N_224,In_451,In_932);
xor U225 (N_225,In_641,In_61);
nand U226 (N_226,In_122,In_739);
and U227 (N_227,In_68,In_335);
nor U228 (N_228,In_349,In_499);
nor U229 (N_229,In_465,In_985);
xor U230 (N_230,In_472,In_448);
nor U231 (N_231,In_288,In_795);
or U232 (N_232,In_33,In_539);
nand U233 (N_233,In_538,In_821);
nor U234 (N_234,In_251,In_904);
nor U235 (N_235,In_990,In_972);
xor U236 (N_236,In_234,In_291);
nor U237 (N_237,In_255,In_359);
xnor U238 (N_238,In_735,In_766);
nor U239 (N_239,In_76,In_540);
nor U240 (N_240,In_571,In_859);
and U241 (N_241,In_701,In_579);
nand U242 (N_242,In_621,In_988);
nor U243 (N_243,In_279,In_899);
xor U244 (N_244,In_470,In_765);
nor U245 (N_245,In_388,In_849);
nand U246 (N_246,In_455,In_829);
nand U247 (N_247,In_123,In_536);
and U248 (N_248,In_215,In_924);
or U249 (N_249,In_534,In_77);
nand U250 (N_250,In_491,In_47);
and U251 (N_251,In_976,In_718);
and U252 (N_252,In_360,In_163);
or U253 (N_253,In_673,In_81);
nor U254 (N_254,In_395,In_908);
nand U255 (N_255,In_809,In_139);
nor U256 (N_256,In_229,In_207);
or U257 (N_257,In_352,In_390);
xor U258 (N_258,In_10,In_897);
and U259 (N_259,In_745,In_630);
xor U260 (N_260,In_252,In_613);
nand U261 (N_261,In_355,In_238);
or U262 (N_262,In_69,In_929);
nand U263 (N_263,In_609,In_557);
nand U264 (N_264,In_703,In_803);
and U265 (N_265,In_125,In_181);
nor U266 (N_266,In_65,In_396);
and U267 (N_267,In_94,In_383);
and U268 (N_268,In_353,In_884);
or U269 (N_269,In_752,In_357);
xnor U270 (N_270,In_638,In_767);
and U271 (N_271,In_490,In_678);
nor U272 (N_272,In_25,In_111);
or U273 (N_273,In_590,In_672);
xnor U274 (N_274,In_154,In_332);
xor U275 (N_275,In_895,In_40);
and U276 (N_276,In_153,In_97);
nand U277 (N_277,In_205,In_546);
nor U278 (N_278,In_57,In_509);
or U279 (N_279,In_844,In_148);
and U280 (N_280,In_324,In_934);
nand U281 (N_281,In_63,In_88);
or U282 (N_282,In_572,In_652);
nand U283 (N_283,In_705,In_38);
or U284 (N_284,In_50,In_670);
xnor U285 (N_285,In_158,In_34);
nor U286 (N_286,In_714,In_285);
xnor U287 (N_287,In_321,In_210);
nand U288 (N_288,In_182,In_447);
nand U289 (N_289,In_775,In_746);
and U290 (N_290,In_526,In_764);
or U291 (N_291,In_341,In_250);
nor U292 (N_292,In_400,In_433);
or U293 (N_293,In_840,In_493);
xnor U294 (N_294,In_569,In_512);
or U295 (N_295,In_813,In_342);
or U296 (N_296,In_307,In_529);
and U297 (N_297,In_728,In_130);
nand U298 (N_298,In_727,In_482);
nand U299 (N_299,In_161,In_39);
and U300 (N_300,In_530,In_424);
or U301 (N_301,In_168,In_48);
nand U302 (N_302,In_497,In_873);
nor U303 (N_303,In_16,In_51);
and U304 (N_304,In_412,In_936);
nand U305 (N_305,In_173,In_958);
nand U306 (N_306,In_909,In_846);
or U307 (N_307,In_254,In_941);
and U308 (N_308,In_865,In_454);
nor U309 (N_309,In_786,In_782);
and U310 (N_310,In_87,In_27);
nor U311 (N_311,In_4,In_501);
and U312 (N_312,In_750,In_9);
or U313 (N_313,In_374,In_686);
nand U314 (N_314,In_789,In_79);
or U315 (N_315,In_217,In_915);
nor U316 (N_316,In_555,In_553);
and U317 (N_317,In_314,In_788);
nor U318 (N_318,In_511,In_610);
nor U319 (N_319,In_889,In_861);
or U320 (N_320,In_82,In_682);
or U321 (N_321,In_710,In_504);
nor U322 (N_322,In_156,In_394);
xnor U323 (N_323,In_877,In_303);
and U324 (N_324,In_760,In_677);
nand U325 (N_325,In_691,In_615);
xor U326 (N_326,In_731,In_668);
nor U327 (N_327,In_758,In_322);
or U328 (N_328,In_777,In_558);
nor U329 (N_329,In_737,In_41);
nor U330 (N_330,In_987,In_826);
or U331 (N_331,In_351,In_720);
and U332 (N_332,In_741,In_828);
or U333 (N_333,In_219,In_43);
nand U334 (N_334,In_289,In_298);
nor U335 (N_335,In_370,In_651);
xor U336 (N_336,In_426,In_922);
xor U337 (N_337,In_824,In_257);
and U338 (N_338,In_883,In_267);
nand U339 (N_339,In_276,In_72);
and U340 (N_340,In_358,In_573);
nor U341 (N_341,In_476,In_875);
nand U342 (N_342,In_583,In_171);
nand U343 (N_343,In_323,In_290);
and U344 (N_344,In_524,In_633);
nand U345 (N_345,In_541,In_92);
or U346 (N_346,In_577,In_271);
nand U347 (N_347,In_820,In_707);
or U348 (N_348,In_507,In_327);
nand U349 (N_349,In_75,In_656);
nor U350 (N_350,In_954,In_386);
xor U351 (N_351,In_421,In_384);
nand U352 (N_352,In_435,In_855);
or U353 (N_353,In_136,In_264);
and U354 (N_354,In_117,In_823);
and U355 (N_355,In_706,In_600);
and U356 (N_356,In_213,In_995);
or U357 (N_357,In_920,In_389);
and U358 (N_358,In_649,In_625);
and U359 (N_359,In_474,In_274);
nor U360 (N_360,In_957,In_780);
nor U361 (N_361,In_712,In_282);
nor U362 (N_362,In_90,In_403);
nand U363 (N_363,In_78,In_29);
xor U364 (N_364,In_439,In_979);
nand U365 (N_365,In_671,In_778);
or U366 (N_366,In_231,In_268);
xor U367 (N_367,In_544,In_612);
nand U368 (N_368,In_177,In_399);
nand U369 (N_369,In_49,In_964);
nor U370 (N_370,In_463,In_992);
or U371 (N_371,In_965,In_151);
nand U372 (N_372,In_519,In_602);
nand U373 (N_373,In_657,In_692);
nand U374 (N_374,In_551,In_337);
nand U375 (N_375,In_15,In_348);
and U376 (N_376,In_771,In_785);
nor U377 (N_377,In_317,In_449);
nor U378 (N_378,In_260,In_70);
nor U379 (N_379,In_948,In_220);
and U380 (N_380,In_200,In_584);
and U381 (N_381,In_894,In_397);
nand U382 (N_382,In_378,In_781);
and U383 (N_383,In_845,In_304);
xnor U384 (N_384,In_848,In_364);
nor U385 (N_385,In_489,In_413);
xnor U386 (N_386,In_850,In_392);
nand U387 (N_387,In_947,In_235);
nand U388 (N_388,In_346,In_818);
nor U389 (N_389,In_847,In_931);
or U390 (N_390,In_836,In_462);
nor U391 (N_391,In_134,In_693);
nor U392 (N_392,In_640,In_773);
nor U393 (N_393,In_330,In_660);
nand U394 (N_394,In_862,In_974);
xor U395 (N_395,In_599,In_632);
and U396 (N_396,In_402,In_445);
nand U397 (N_397,In_0,In_554);
xnor U398 (N_398,In_639,In_469);
or U399 (N_399,In_272,In_664);
or U400 (N_400,In_804,In_940);
xnor U401 (N_401,In_110,In_361);
nand U402 (N_402,In_627,In_408);
xor U403 (N_403,In_404,In_960);
or U404 (N_404,In_683,In_437);
and U405 (N_405,In_297,In_120);
nor U406 (N_406,In_146,In_431);
nand U407 (N_407,In_736,In_981);
nor U408 (N_408,In_882,In_770);
xnor U409 (N_409,In_938,In_186);
nor U410 (N_410,In_831,In_808);
or U411 (N_411,In_326,In_869);
and U412 (N_412,In_906,In_646);
or U413 (N_413,In_618,In_385);
nand U414 (N_414,In_429,In_680);
xor U415 (N_415,In_801,In_921);
and U416 (N_416,In_410,In_545);
xor U417 (N_417,In_738,In_653);
xor U418 (N_418,In_834,In_138);
xor U419 (N_419,In_772,In_616);
or U420 (N_420,In_790,In_30);
and U421 (N_421,In_912,In_567);
and U422 (N_422,In_977,In_881);
and U423 (N_423,In_26,In_188);
nor U424 (N_424,In_407,In_7);
xnor U425 (N_425,In_137,In_176);
nand U426 (N_426,In_159,In_853);
and U427 (N_427,In_838,In_259);
and U428 (N_428,In_843,In_604);
nor U429 (N_429,In_574,In_363);
and U430 (N_430,In_129,In_961);
xor U431 (N_431,In_661,In_689);
and U432 (N_432,In_880,In_467);
or U433 (N_433,In_199,In_515);
xor U434 (N_434,In_852,In_756);
xnor U435 (N_435,In_305,In_222);
and U436 (N_436,In_299,In_654);
xnor U437 (N_437,In_232,In_37);
xnor U438 (N_438,In_1,In_800);
nor U439 (N_439,In_690,In_896);
xnor U440 (N_440,In_949,In_776);
and U441 (N_441,In_575,In_64);
nand U442 (N_442,In_377,In_226);
xnor U443 (N_443,In_930,In_702);
and U444 (N_444,In_637,In_356);
nor U445 (N_445,In_477,In_851);
nand U446 (N_446,In_528,In_165);
nor U447 (N_447,In_144,In_334);
and U448 (N_448,In_565,In_141);
nand U449 (N_449,In_608,In_535);
and U450 (N_450,In_379,In_700);
nor U451 (N_451,In_963,In_724);
nand U452 (N_452,In_121,In_833);
and U453 (N_453,In_84,In_145);
nand U454 (N_454,In_914,In_461);
and U455 (N_455,In_118,In_416);
and U456 (N_456,In_763,In_753);
nor U457 (N_457,In_498,In_581);
nand U458 (N_458,In_265,In_488);
and U459 (N_459,In_955,In_913);
xor U460 (N_460,In_486,In_23);
xor U461 (N_461,In_761,In_503);
or U462 (N_462,In_18,In_525);
and U463 (N_463,In_628,In_945);
or U464 (N_464,In_366,In_885);
nand U465 (N_465,In_774,In_902);
or U466 (N_466,In_592,In_919);
nor U467 (N_467,In_547,In_973);
and U468 (N_468,In_797,In_164);
nand U469 (N_469,In_505,In_127);
xnor U470 (N_470,In_697,In_872);
or U471 (N_471,In_910,In_799);
and U472 (N_472,In_681,In_740);
xor U473 (N_473,In_994,In_5);
xnor U474 (N_474,In_550,In_329);
or U475 (N_475,In_194,In_514);
or U476 (N_476,In_13,In_12);
and U477 (N_477,In_928,In_135);
xnor U478 (N_478,In_563,In_185);
xnor U479 (N_479,In_732,In_623);
or U480 (N_480,In_203,In_980);
xnor U481 (N_481,In_133,In_796);
nor U482 (N_482,In_982,In_103);
nor U483 (N_483,In_594,In_966);
xor U484 (N_484,In_372,In_6);
nor U485 (N_485,In_59,In_457);
nor U486 (N_486,In_8,In_101);
xor U487 (N_487,In_391,In_54);
xor U488 (N_488,In_336,In_409);
nor U489 (N_489,In_108,In_685);
nor U490 (N_490,In_430,In_825);
nor U491 (N_491,In_227,In_725);
xor U492 (N_492,In_570,In_105);
and U493 (N_493,In_787,In_126);
or U494 (N_494,In_479,In_478);
nor U495 (N_495,In_417,In_598);
and U496 (N_496,In_85,In_698);
and U497 (N_497,In_420,In_446);
nand U498 (N_498,In_560,In_55);
nand U499 (N_499,In_742,In_518);
nor U500 (N_500,In_807,In_458);
or U501 (N_501,In_63,In_541);
xnor U502 (N_502,In_917,In_12);
nand U503 (N_503,In_425,In_213);
and U504 (N_504,In_245,In_269);
nand U505 (N_505,In_351,In_682);
nor U506 (N_506,In_989,In_969);
and U507 (N_507,In_812,In_426);
or U508 (N_508,In_17,In_825);
or U509 (N_509,In_707,In_64);
xor U510 (N_510,In_758,In_685);
nand U511 (N_511,In_508,In_223);
or U512 (N_512,In_142,In_751);
and U513 (N_513,In_405,In_415);
or U514 (N_514,In_48,In_855);
nor U515 (N_515,In_65,In_200);
and U516 (N_516,In_296,In_320);
nand U517 (N_517,In_100,In_950);
and U518 (N_518,In_784,In_889);
xor U519 (N_519,In_803,In_873);
and U520 (N_520,In_345,In_558);
nand U521 (N_521,In_810,In_521);
nand U522 (N_522,In_995,In_676);
nor U523 (N_523,In_179,In_648);
nand U524 (N_524,In_755,In_639);
and U525 (N_525,In_652,In_903);
nor U526 (N_526,In_445,In_678);
and U527 (N_527,In_228,In_662);
xnor U528 (N_528,In_513,In_340);
nand U529 (N_529,In_701,In_383);
nor U530 (N_530,In_546,In_450);
nor U531 (N_531,In_267,In_411);
nand U532 (N_532,In_587,In_773);
nand U533 (N_533,In_407,In_965);
xnor U534 (N_534,In_743,In_363);
or U535 (N_535,In_444,In_215);
nor U536 (N_536,In_558,In_322);
and U537 (N_537,In_113,In_73);
nand U538 (N_538,In_973,In_908);
nand U539 (N_539,In_837,In_777);
nor U540 (N_540,In_893,In_172);
nand U541 (N_541,In_541,In_479);
nand U542 (N_542,In_458,In_364);
nand U543 (N_543,In_23,In_274);
nand U544 (N_544,In_793,In_229);
nor U545 (N_545,In_334,In_572);
or U546 (N_546,In_711,In_422);
xnor U547 (N_547,In_411,In_966);
and U548 (N_548,In_77,In_576);
xor U549 (N_549,In_702,In_156);
nor U550 (N_550,In_984,In_744);
nand U551 (N_551,In_335,In_385);
nor U552 (N_552,In_481,In_563);
nor U553 (N_553,In_9,In_966);
or U554 (N_554,In_438,In_53);
nor U555 (N_555,In_401,In_56);
or U556 (N_556,In_834,In_379);
or U557 (N_557,In_997,In_576);
or U558 (N_558,In_733,In_736);
or U559 (N_559,In_548,In_305);
and U560 (N_560,In_79,In_431);
nand U561 (N_561,In_114,In_515);
or U562 (N_562,In_622,In_61);
nand U563 (N_563,In_49,In_27);
nand U564 (N_564,In_332,In_799);
nand U565 (N_565,In_119,In_435);
nor U566 (N_566,In_576,In_748);
nor U567 (N_567,In_4,In_305);
nand U568 (N_568,In_872,In_451);
nor U569 (N_569,In_160,In_593);
or U570 (N_570,In_146,In_859);
or U571 (N_571,In_531,In_614);
xor U572 (N_572,In_570,In_379);
nand U573 (N_573,In_480,In_369);
xnor U574 (N_574,In_626,In_78);
or U575 (N_575,In_403,In_426);
nand U576 (N_576,In_709,In_393);
or U577 (N_577,In_621,In_311);
xnor U578 (N_578,In_462,In_128);
nor U579 (N_579,In_19,In_970);
nor U580 (N_580,In_632,In_527);
nand U581 (N_581,In_261,In_525);
nor U582 (N_582,In_722,In_984);
xnor U583 (N_583,In_524,In_513);
nand U584 (N_584,In_782,In_973);
or U585 (N_585,In_689,In_608);
and U586 (N_586,In_389,In_673);
nand U587 (N_587,In_441,In_723);
nand U588 (N_588,In_33,In_807);
or U589 (N_589,In_679,In_390);
xor U590 (N_590,In_620,In_642);
nand U591 (N_591,In_940,In_926);
or U592 (N_592,In_968,In_717);
nor U593 (N_593,In_686,In_32);
or U594 (N_594,In_135,In_879);
xnor U595 (N_595,In_142,In_225);
nand U596 (N_596,In_177,In_496);
xnor U597 (N_597,In_701,In_445);
or U598 (N_598,In_144,In_282);
xor U599 (N_599,In_726,In_528);
and U600 (N_600,In_656,In_212);
nor U601 (N_601,In_230,In_998);
nor U602 (N_602,In_579,In_960);
nand U603 (N_603,In_890,In_610);
and U604 (N_604,In_282,In_400);
xor U605 (N_605,In_653,In_560);
nand U606 (N_606,In_556,In_8);
and U607 (N_607,In_486,In_100);
and U608 (N_608,In_92,In_955);
xnor U609 (N_609,In_725,In_724);
nand U610 (N_610,In_199,In_990);
and U611 (N_611,In_356,In_354);
or U612 (N_612,In_418,In_489);
xor U613 (N_613,In_38,In_233);
nand U614 (N_614,In_881,In_410);
xor U615 (N_615,In_278,In_962);
nand U616 (N_616,In_511,In_679);
or U617 (N_617,In_667,In_537);
xnor U618 (N_618,In_307,In_381);
xnor U619 (N_619,In_352,In_44);
nand U620 (N_620,In_962,In_86);
nand U621 (N_621,In_79,In_925);
xnor U622 (N_622,In_573,In_57);
or U623 (N_623,In_422,In_493);
nand U624 (N_624,In_180,In_539);
or U625 (N_625,In_972,In_108);
or U626 (N_626,In_27,In_190);
xnor U627 (N_627,In_913,In_613);
nand U628 (N_628,In_186,In_349);
and U629 (N_629,In_303,In_945);
nor U630 (N_630,In_246,In_562);
nor U631 (N_631,In_44,In_295);
nor U632 (N_632,In_403,In_551);
xor U633 (N_633,In_444,In_442);
or U634 (N_634,In_585,In_412);
xnor U635 (N_635,In_65,In_257);
nor U636 (N_636,In_263,In_890);
nand U637 (N_637,In_146,In_678);
nand U638 (N_638,In_558,In_456);
and U639 (N_639,In_903,In_129);
nor U640 (N_640,In_626,In_964);
and U641 (N_641,In_672,In_329);
nor U642 (N_642,In_379,In_676);
nand U643 (N_643,In_97,In_377);
nand U644 (N_644,In_967,In_343);
nor U645 (N_645,In_774,In_10);
xnor U646 (N_646,In_312,In_551);
nor U647 (N_647,In_411,In_136);
nor U648 (N_648,In_763,In_684);
and U649 (N_649,In_485,In_687);
or U650 (N_650,In_765,In_832);
and U651 (N_651,In_690,In_926);
xnor U652 (N_652,In_715,In_981);
nor U653 (N_653,In_728,In_633);
and U654 (N_654,In_624,In_424);
and U655 (N_655,In_469,In_624);
nor U656 (N_656,In_84,In_938);
nor U657 (N_657,In_403,In_888);
nand U658 (N_658,In_133,In_38);
xnor U659 (N_659,In_920,In_369);
or U660 (N_660,In_90,In_621);
xnor U661 (N_661,In_972,In_994);
nand U662 (N_662,In_98,In_269);
and U663 (N_663,In_124,In_224);
xnor U664 (N_664,In_739,In_925);
nand U665 (N_665,In_141,In_636);
and U666 (N_666,In_630,In_231);
or U667 (N_667,In_96,In_321);
xnor U668 (N_668,In_606,In_319);
xor U669 (N_669,In_232,In_136);
or U670 (N_670,In_589,In_902);
xnor U671 (N_671,In_349,In_18);
and U672 (N_672,In_896,In_230);
and U673 (N_673,In_730,In_843);
xnor U674 (N_674,In_503,In_917);
xor U675 (N_675,In_836,In_736);
nor U676 (N_676,In_816,In_547);
nor U677 (N_677,In_341,In_625);
nand U678 (N_678,In_745,In_522);
xnor U679 (N_679,In_83,In_474);
nand U680 (N_680,In_772,In_502);
and U681 (N_681,In_851,In_617);
nor U682 (N_682,In_138,In_41);
and U683 (N_683,In_30,In_377);
or U684 (N_684,In_347,In_333);
and U685 (N_685,In_581,In_981);
or U686 (N_686,In_139,In_285);
xnor U687 (N_687,In_675,In_252);
nor U688 (N_688,In_915,In_802);
xor U689 (N_689,In_956,In_932);
xnor U690 (N_690,In_81,In_621);
nor U691 (N_691,In_124,In_404);
nor U692 (N_692,In_364,In_652);
nand U693 (N_693,In_609,In_781);
nand U694 (N_694,In_780,In_87);
and U695 (N_695,In_102,In_733);
nor U696 (N_696,In_779,In_461);
or U697 (N_697,In_50,In_631);
or U698 (N_698,In_876,In_272);
nand U699 (N_699,In_644,In_82);
or U700 (N_700,In_578,In_185);
nand U701 (N_701,In_544,In_205);
xnor U702 (N_702,In_602,In_553);
nand U703 (N_703,In_289,In_718);
nor U704 (N_704,In_343,In_147);
xor U705 (N_705,In_573,In_375);
nand U706 (N_706,In_386,In_601);
and U707 (N_707,In_940,In_637);
and U708 (N_708,In_985,In_590);
or U709 (N_709,In_556,In_514);
nand U710 (N_710,In_6,In_986);
nor U711 (N_711,In_155,In_472);
nor U712 (N_712,In_918,In_867);
and U713 (N_713,In_831,In_441);
nor U714 (N_714,In_196,In_996);
xnor U715 (N_715,In_518,In_601);
nand U716 (N_716,In_919,In_940);
xnor U717 (N_717,In_897,In_929);
xor U718 (N_718,In_1,In_965);
nor U719 (N_719,In_573,In_183);
or U720 (N_720,In_346,In_709);
and U721 (N_721,In_436,In_786);
nor U722 (N_722,In_358,In_197);
and U723 (N_723,In_56,In_117);
or U724 (N_724,In_973,In_173);
or U725 (N_725,In_23,In_139);
nand U726 (N_726,In_768,In_286);
or U727 (N_727,In_297,In_138);
nor U728 (N_728,In_973,In_590);
or U729 (N_729,In_788,In_503);
xor U730 (N_730,In_448,In_828);
nand U731 (N_731,In_917,In_389);
nand U732 (N_732,In_497,In_605);
and U733 (N_733,In_38,In_997);
or U734 (N_734,In_208,In_227);
nor U735 (N_735,In_574,In_367);
nor U736 (N_736,In_651,In_926);
and U737 (N_737,In_146,In_410);
xnor U738 (N_738,In_390,In_316);
or U739 (N_739,In_482,In_207);
nor U740 (N_740,In_422,In_195);
and U741 (N_741,In_678,In_104);
nand U742 (N_742,In_152,In_698);
nor U743 (N_743,In_664,In_36);
nand U744 (N_744,In_382,In_918);
or U745 (N_745,In_605,In_253);
or U746 (N_746,In_712,In_916);
nand U747 (N_747,In_466,In_22);
or U748 (N_748,In_556,In_157);
xor U749 (N_749,In_402,In_326);
nand U750 (N_750,In_49,In_313);
or U751 (N_751,In_470,In_638);
nor U752 (N_752,In_283,In_208);
nor U753 (N_753,In_687,In_525);
nor U754 (N_754,In_483,In_847);
nand U755 (N_755,In_601,In_398);
nand U756 (N_756,In_946,In_318);
or U757 (N_757,In_578,In_724);
and U758 (N_758,In_665,In_542);
or U759 (N_759,In_960,In_291);
nor U760 (N_760,In_337,In_767);
and U761 (N_761,In_610,In_918);
nor U762 (N_762,In_333,In_779);
nor U763 (N_763,In_743,In_65);
nand U764 (N_764,In_198,In_297);
nor U765 (N_765,In_381,In_599);
xor U766 (N_766,In_734,In_576);
or U767 (N_767,In_748,In_194);
and U768 (N_768,In_613,In_812);
and U769 (N_769,In_551,In_703);
nor U770 (N_770,In_657,In_547);
xnor U771 (N_771,In_447,In_330);
nand U772 (N_772,In_72,In_773);
nand U773 (N_773,In_642,In_74);
or U774 (N_774,In_769,In_57);
xor U775 (N_775,In_116,In_209);
xnor U776 (N_776,In_399,In_9);
nor U777 (N_777,In_199,In_125);
and U778 (N_778,In_980,In_70);
nand U779 (N_779,In_855,In_470);
nor U780 (N_780,In_673,In_109);
nor U781 (N_781,In_153,In_198);
nand U782 (N_782,In_350,In_841);
or U783 (N_783,In_981,In_575);
nand U784 (N_784,In_10,In_302);
xnor U785 (N_785,In_817,In_478);
nor U786 (N_786,In_463,In_243);
xnor U787 (N_787,In_652,In_48);
or U788 (N_788,In_333,In_23);
nand U789 (N_789,In_174,In_82);
nand U790 (N_790,In_173,In_302);
nand U791 (N_791,In_271,In_525);
nor U792 (N_792,In_128,In_998);
nor U793 (N_793,In_120,In_870);
nand U794 (N_794,In_842,In_401);
or U795 (N_795,In_976,In_277);
nor U796 (N_796,In_538,In_285);
or U797 (N_797,In_470,In_285);
or U798 (N_798,In_311,In_558);
nand U799 (N_799,In_591,In_33);
xor U800 (N_800,In_577,In_942);
nand U801 (N_801,In_651,In_279);
nand U802 (N_802,In_804,In_781);
nor U803 (N_803,In_838,In_646);
nor U804 (N_804,In_328,In_869);
or U805 (N_805,In_34,In_400);
xnor U806 (N_806,In_681,In_957);
nor U807 (N_807,In_57,In_888);
nand U808 (N_808,In_906,In_568);
nand U809 (N_809,In_606,In_743);
and U810 (N_810,In_390,In_776);
xor U811 (N_811,In_628,In_724);
and U812 (N_812,In_372,In_790);
xnor U813 (N_813,In_716,In_85);
nand U814 (N_814,In_235,In_705);
and U815 (N_815,In_352,In_471);
nand U816 (N_816,In_187,In_814);
and U817 (N_817,In_885,In_784);
or U818 (N_818,In_332,In_251);
and U819 (N_819,In_521,In_707);
nor U820 (N_820,In_212,In_510);
nand U821 (N_821,In_685,In_188);
nand U822 (N_822,In_776,In_169);
nand U823 (N_823,In_825,In_725);
and U824 (N_824,In_415,In_130);
and U825 (N_825,In_616,In_924);
and U826 (N_826,In_681,In_585);
nand U827 (N_827,In_920,In_69);
or U828 (N_828,In_360,In_483);
nand U829 (N_829,In_450,In_88);
nor U830 (N_830,In_741,In_930);
nor U831 (N_831,In_627,In_232);
xor U832 (N_832,In_888,In_374);
nor U833 (N_833,In_71,In_817);
nor U834 (N_834,In_864,In_398);
nor U835 (N_835,In_921,In_246);
nand U836 (N_836,In_331,In_598);
nor U837 (N_837,In_731,In_526);
or U838 (N_838,In_625,In_828);
xnor U839 (N_839,In_815,In_87);
xnor U840 (N_840,In_459,In_250);
nand U841 (N_841,In_730,In_49);
xor U842 (N_842,In_512,In_143);
or U843 (N_843,In_823,In_92);
nand U844 (N_844,In_606,In_80);
nand U845 (N_845,In_365,In_592);
nand U846 (N_846,In_342,In_985);
nand U847 (N_847,In_765,In_286);
xor U848 (N_848,In_843,In_777);
nor U849 (N_849,In_304,In_532);
or U850 (N_850,In_775,In_256);
or U851 (N_851,In_99,In_482);
and U852 (N_852,In_162,In_23);
nor U853 (N_853,In_914,In_613);
xor U854 (N_854,In_230,In_840);
and U855 (N_855,In_95,In_241);
and U856 (N_856,In_510,In_957);
and U857 (N_857,In_199,In_217);
and U858 (N_858,In_316,In_105);
and U859 (N_859,In_504,In_838);
and U860 (N_860,In_97,In_235);
nand U861 (N_861,In_334,In_27);
nor U862 (N_862,In_565,In_161);
xnor U863 (N_863,In_765,In_30);
xnor U864 (N_864,In_874,In_980);
or U865 (N_865,In_855,In_611);
and U866 (N_866,In_373,In_195);
nor U867 (N_867,In_71,In_427);
nor U868 (N_868,In_222,In_431);
or U869 (N_869,In_907,In_86);
xor U870 (N_870,In_878,In_337);
nand U871 (N_871,In_547,In_834);
xor U872 (N_872,In_828,In_85);
nor U873 (N_873,In_481,In_143);
and U874 (N_874,In_794,In_851);
and U875 (N_875,In_530,In_338);
or U876 (N_876,In_124,In_211);
nor U877 (N_877,In_853,In_37);
xor U878 (N_878,In_478,In_512);
and U879 (N_879,In_321,In_940);
or U880 (N_880,In_916,In_777);
nand U881 (N_881,In_51,In_480);
or U882 (N_882,In_372,In_458);
xnor U883 (N_883,In_939,In_135);
or U884 (N_884,In_797,In_37);
xor U885 (N_885,In_32,In_75);
or U886 (N_886,In_157,In_214);
or U887 (N_887,In_866,In_164);
or U888 (N_888,In_221,In_213);
nor U889 (N_889,In_376,In_92);
nand U890 (N_890,In_573,In_419);
and U891 (N_891,In_45,In_606);
and U892 (N_892,In_616,In_303);
and U893 (N_893,In_495,In_340);
nand U894 (N_894,In_185,In_297);
nor U895 (N_895,In_607,In_740);
xor U896 (N_896,In_178,In_723);
nand U897 (N_897,In_470,In_146);
nand U898 (N_898,In_995,In_47);
and U899 (N_899,In_991,In_676);
nor U900 (N_900,In_650,In_416);
and U901 (N_901,In_819,In_392);
or U902 (N_902,In_691,In_556);
xor U903 (N_903,In_207,In_251);
or U904 (N_904,In_263,In_923);
xnor U905 (N_905,In_677,In_211);
nor U906 (N_906,In_26,In_905);
xor U907 (N_907,In_843,In_931);
and U908 (N_908,In_758,In_994);
or U909 (N_909,In_348,In_276);
and U910 (N_910,In_378,In_753);
nor U911 (N_911,In_533,In_459);
xor U912 (N_912,In_88,In_621);
nand U913 (N_913,In_914,In_655);
nor U914 (N_914,In_615,In_784);
xor U915 (N_915,In_91,In_634);
xnor U916 (N_916,In_773,In_627);
nand U917 (N_917,In_631,In_101);
nand U918 (N_918,In_665,In_973);
nand U919 (N_919,In_496,In_894);
and U920 (N_920,In_726,In_919);
or U921 (N_921,In_486,In_813);
xor U922 (N_922,In_841,In_650);
or U923 (N_923,In_58,In_314);
xnor U924 (N_924,In_671,In_720);
xor U925 (N_925,In_743,In_21);
nand U926 (N_926,In_814,In_284);
xnor U927 (N_927,In_983,In_965);
or U928 (N_928,In_646,In_488);
and U929 (N_929,In_794,In_338);
nand U930 (N_930,In_860,In_333);
nand U931 (N_931,In_122,In_842);
xor U932 (N_932,In_857,In_984);
nand U933 (N_933,In_697,In_978);
nor U934 (N_934,In_823,In_764);
and U935 (N_935,In_632,In_612);
nor U936 (N_936,In_861,In_40);
nor U937 (N_937,In_213,In_52);
or U938 (N_938,In_446,In_14);
or U939 (N_939,In_352,In_204);
and U940 (N_940,In_280,In_0);
and U941 (N_941,In_14,In_370);
nor U942 (N_942,In_178,In_971);
xnor U943 (N_943,In_275,In_192);
and U944 (N_944,In_885,In_380);
or U945 (N_945,In_395,In_961);
and U946 (N_946,In_757,In_63);
and U947 (N_947,In_579,In_559);
nand U948 (N_948,In_830,In_764);
or U949 (N_949,In_950,In_739);
and U950 (N_950,In_653,In_808);
and U951 (N_951,In_729,In_674);
nand U952 (N_952,In_211,In_329);
nor U953 (N_953,In_639,In_412);
nor U954 (N_954,In_457,In_474);
and U955 (N_955,In_622,In_15);
and U956 (N_956,In_785,In_157);
and U957 (N_957,In_289,In_767);
and U958 (N_958,In_57,In_54);
or U959 (N_959,In_777,In_338);
or U960 (N_960,In_483,In_357);
xnor U961 (N_961,In_500,In_530);
and U962 (N_962,In_685,In_501);
and U963 (N_963,In_857,In_633);
or U964 (N_964,In_612,In_555);
nand U965 (N_965,In_282,In_765);
xor U966 (N_966,In_755,In_620);
nor U967 (N_967,In_982,In_382);
nor U968 (N_968,In_955,In_594);
and U969 (N_969,In_563,In_872);
or U970 (N_970,In_967,In_477);
nand U971 (N_971,In_844,In_651);
and U972 (N_972,In_645,In_330);
xor U973 (N_973,In_724,In_486);
nor U974 (N_974,In_680,In_665);
nand U975 (N_975,In_145,In_601);
xnor U976 (N_976,In_429,In_709);
xnor U977 (N_977,In_982,In_378);
and U978 (N_978,In_670,In_322);
or U979 (N_979,In_775,In_833);
or U980 (N_980,In_557,In_348);
xnor U981 (N_981,In_167,In_999);
xor U982 (N_982,In_225,In_248);
xnor U983 (N_983,In_186,In_633);
and U984 (N_984,In_477,In_721);
nand U985 (N_985,In_659,In_43);
and U986 (N_986,In_678,In_9);
nor U987 (N_987,In_142,In_978);
nor U988 (N_988,In_580,In_802);
or U989 (N_989,In_400,In_365);
nor U990 (N_990,In_746,In_184);
xor U991 (N_991,In_395,In_645);
nand U992 (N_992,In_760,In_166);
or U993 (N_993,In_336,In_731);
or U994 (N_994,In_815,In_697);
and U995 (N_995,In_826,In_478);
and U996 (N_996,In_339,In_495);
nor U997 (N_997,In_27,In_444);
nor U998 (N_998,In_512,In_180);
xnor U999 (N_999,In_14,In_929);
xor U1000 (N_1000,In_435,In_374);
and U1001 (N_1001,In_584,In_724);
xnor U1002 (N_1002,In_796,In_485);
nand U1003 (N_1003,In_572,In_951);
and U1004 (N_1004,In_601,In_656);
or U1005 (N_1005,In_890,In_677);
or U1006 (N_1006,In_578,In_883);
or U1007 (N_1007,In_210,In_486);
nand U1008 (N_1008,In_626,In_612);
xnor U1009 (N_1009,In_229,In_471);
or U1010 (N_1010,In_303,In_257);
or U1011 (N_1011,In_952,In_258);
and U1012 (N_1012,In_906,In_577);
and U1013 (N_1013,In_366,In_568);
and U1014 (N_1014,In_507,In_873);
nor U1015 (N_1015,In_820,In_22);
nand U1016 (N_1016,In_64,In_439);
nand U1017 (N_1017,In_552,In_168);
nor U1018 (N_1018,In_651,In_277);
nor U1019 (N_1019,In_616,In_426);
or U1020 (N_1020,In_429,In_847);
nand U1021 (N_1021,In_461,In_173);
nand U1022 (N_1022,In_361,In_158);
and U1023 (N_1023,In_13,In_55);
or U1024 (N_1024,In_327,In_472);
or U1025 (N_1025,In_23,In_673);
xor U1026 (N_1026,In_577,In_951);
nand U1027 (N_1027,In_293,In_600);
nand U1028 (N_1028,In_181,In_130);
nand U1029 (N_1029,In_358,In_223);
xor U1030 (N_1030,In_797,In_732);
or U1031 (N_1031,In_245,In_658);
nand U1032 (N_1032,In_456,In_870);
xor U1033 (N_1033,In_119,In_477);
or U1034 (N_1034,In_850,In_298);
or U1035 (N_1035,In_981,In_149);
or U1036 (N_1036,In_400,In_653);
and U1037 (N_1037,In_786,In_89);
xor U1038 (N_1038,In_303,In_183);
and U1039 (N_1039,In_77,In_597);
or U1040 (N_1040,In_606,In_526);
nand U1041 (N_1041,In_182,In_88);
or U1042 (N_1042,In_329,In_564);
nor U1043 (N_1043,In_232,In_279);
nor U1044 (N_1044,In_710,In_586);
nor U1045 (N_1045,In_789,In_564);
and U1046 (N_1046,In_137,In_75);
and U1047 (N_1047,In_653,In_588);
nand U1048 (N_1048,In_877,In_6);
nand U1049 (N_1049,In_774,In_44);
or U1050 (N_1050,In_422,In_383);
nand U1051 (N_1051,In_691,In_896);
xor U1052 (N_1052,In_240,In_868);
and U1053 (N_1053,In_222,In_230);
nor U1054 (N_1054,In_100,In_857);
and U1055 (N_1055,In_837,In_462);
or U1056 (N_1056,In_810,In_563);
nor U1057 (N_1057,In_665,In_320);
xnor U1058 (N_1058,In_936,In_197);
xor U1059 (N_1059,In_681,In_205);
nand U1060 (N_1060,In_916,In_437);
nor U1061 (N_1061,In_660,In_261);
xor U1062 (N_1062,In_104,In_312);
xnor U1063 (N_1063,In_648,In_541);
nor U1064 (N_1064,In_305,In_491);
nand U1065 (N_1065,In_683,In_695);
nor U1066 (N_1066,In_291,In_414);
xnor U1067 (N_1067,In_384,In_805);
nand U1068 (N_1068,In_311,In_265);
xnor U1069 (N_1069,In_728,In_163);
and U1070 (N_1070,In_330,In_790);
nor U1071 (N_1071,In_323,In_497);
or U1072 (N_1072,In_156,In_454);
and U1073 (N_1073,In_582,In_236);
nand U1074 (N_1074,In_592,In_616);
and U1075 (N_1075,In_135,In_40);
nor U1076 (N_1076,In_137,In_973);
nand U1077 (N_1077,In_116,In_766);
nor U1078 (N_1078,In_527,In_558);
and U1079 (N_1079,In_48,In_258);
nor U1080 (N_1080,In_806,In_206);
xnor U1081 (N_1081,In_572,In_1);
nor U1082 (N_1082,In_200,In_171);
and U1083 (N_1083,In_241,In_871);
xnor U1084 (N_1084,In_177,In_516);
or U1085 (N_1085,In_155,In_360);
nor U1086 (N_1086,In_695,In_162);
nand U1087 (N_1087,In_973,In_643);
or U1088 (N_1088,In_882,In_339);
nor U1089 (N_1089,In_414,In_197);
xor U1090 (N_1090,In_791,In_433);
or U1091 (N_1091,In_31,In_105);
nor U1092 (N_1092,In_96,In_3);
and U1093 (N_1093,In_158,In_938);
nor U1094 (N_1094,In_172,In_497);
xnor U1095 (N_1095,In_782,In_851);
and U1096 (N_1096,In_35,In_518);
or U1097 (N_1097,In_741,In_719);
or U1098 (N_1098,In_369,In_319);
and U1099 (N_1099,In_649,In_673);
nor U1100 (N_1100,In_441,In_774);
nand U1101 (N_1101,In_924,In_640);
nand U1102 (N_1102,In_44,In_373);
nor U1103 (N_1103,In_115,In_993);
nor U1104 (N_1104,In_734,In_253);
nand U1105 (N_1105,In_639,In_860);
or U1106 (N_1106,In_835,In_715);
or U1107 (N_1107,In_631,In_360);
and U1108 (N_1108,In_289,In_368);
nand U1109 (N_1109,In_96,In_711);
nor U1110 (N_1110,In_692,In_328);
or U1111 (N_1111,In_527,In_993);
or U1112 (N_1112,In_888,In_596);
and U1113 (N_1113,In_811,In_576);
or U1114 (N_1114,In_993,In_966);
or U1115 (N_1115,In_274,In_223);
or U1116 (N_1116,In_282,In_817);
nand U1117 (N_1117,In_128,In_573);
nand U1118 (N_1118,In_802,In_708);
nand U1119 (N_1119,In_99,In_316);
or U1120 (N_1120,In_822,In_219);
nor U1121 (N_1121,In_643,In_234);
xnor U1122 (N_1122,In_593,In_199);
nor U1123 (N_1123,In_664,In_167);
nor U1124 (N_1124,In_383,In_884);
or U1125 (N_1125,In_662,In_30);
and U1126 (N_1126,In_720,In_232);
nand U1127 (N_1127,In_257,In_746);
or U1128 (N_1128,In_77,In_623);
xor U1129 (N_1129,In_762,In_664);
and U1130 (N_1130,In_307,In_684);
nand U1131 (N_1131,In_230,In_284);
or U1132 (N_1132,In_595,In_829);
nand U1133 (N_1133,In_933,In_82);
nor U1134 (N_1134,In_451,In_648);
or U1135 (N_1135,In_178,In_818);
or U1136 (N_1136,In_737,In_13);
nor U1137 (N_1137,In_646,In_174);
or U1138 (N_1138,In_588,In_32);
xnor U1139 (N_1139,In_474,In_392);
xnor U1140 (N_1140,In_287,In_526);
xor U1141 (N_1141,In_986,In_980);
and U1142 (N_1142,In_721,In_966);
and U1143 (N_1143,In_547,In_215);
xor U1144 (N_1144,In_474,In_704);
nor U1145 (N_1145,In_697,In_867);
xnor U1146 (N_1146,In_653,In_849);
xnor U1147 (N_1147,In_644,In_229);
xor U1148 (N_1148,In_480,In_795);
or U1149 (N_1149,In_347,In_916);
and U1150 (N_1150,In_94,In_142);
or U1151 (N_1151,In_404,In_942);
xor U1152 (N_1152,In_103,In_786);
and U1153 (N_1153,In_803,In_531);
and U1154 (N_1154,In_44,In_811);
nor U1155 (N_1155,In_500,In_38);
nor U1156 (N_1156,In_902,In_571);
or U1157 (N_1157,In_614,In_314);
nand U1158 (N_1158,In_847,In_84);
and U1159 (N_1159,In_689,In_747);
nand U1160 (N_1160,In_803,In_236);
nand U1161 (N_1161,In_764,In_852);
and U1162 (N_1162,In_366,In_626);
and U1163 (N_1163,In_692,In_520);
nand U1164 (N_1164,In_735,In_522);
xnor U1165 (N_1165,In_871,In_787);
and U1166 (N_1166,In_900,In_767);
xnor U1167 (N_1167,In_778,In_521);
xor U1168 (N_1168,In_68,In_351);
nor U1169 (N_1169,In_434,In_861);
and U1170 (N_1170,In_286,In_553);
or U1171 (N_1171,In_557,In_940);
and U1172 (N_1172,In_20,In_355);
or U1173 (N_1173,In_320,In_369);
nand U1174 (N_1174,In_420,In_851);
nand U1175 (N_1175,In_319,In_255);
or U1176 (N_1176,In_430,In_575);
nand U1177 (N_1177,In_380,In_181);
xnor U1178 (N_1178,In_234,In_720);
nor U1179 (N_1179,In_496,In_138);
or U1180 (N_1180,In_377,In_872);
and U1181 (N_1181,In_929,In_382);
and U1182 (N_1182,In_800,In_392);
nand U1183 (N_1183,In_783,In_647);
nor U1184 (N_1184,In_173,In_739);
or U1185 (N_1185,In_205,In_781);
xnor U1186 (N_1186,In_155,In_226);
and U1187 (N_1187,In_345,In_448);
xnor U1188 (N_1188,In_931,In_905);
xor U1189 (N_1189,In_109,In_449);
nor U1190 (N_1190,In_378,In_608);
or U1191 (N_1191,In_849,In_729);
or U1192 (N_1192,In_781,In_573);
nand U1193 (N_1193,In_764,In_527);
xor U1194 (N_1194,In_479,In_562);
nor U1195 (N_1195,In_268,In_117);
nand U1196 (N_1196,In_633,In_254);
and U1197 (N_1197,In_776,In_992);
nor U1198 (N_1198,In_80,In_617);
xnor U1199 (N_1199,In_133,In_55);
nor U1200 (N_1200,In_997,In_567);
xnor U1201 (N_1201,In_290,In_150);
and U1202 (N_1202,In_977,In_801);
or U1203 (N_1203,In_120,In_303);
and U1204 (N_1204,In_214,In_669);
xnor U1205 (N_1205,In_2,In_17);
nor U1206 (N_1206,In_73,In_725);
nor U1207 (N_1207,In_220,In_508);
and U1208 (N_1208,In_468,In_656);
nor U1209 (N_1209,In_212,In_327);
xor U1210 (N_1210,In_599,In_189);
and U1211 (N_1211,In_442,In_599);
nand U1212 (N_1212,In_784,In_623);
nand U1213 (N_1213,In_451,In_939);
and U1214 (N_1214,In_707,In_431);
and U1215 (N_1215,In_168,In_232);
and U1216 (N_1216,In_894,In_853);
nand U1217 (N_1217,In_362,In_390);
nand U1218 (N_1218,In_811,In_243);
or U1219 (N_1219,In_784,In_833);
nand U1220 (N_1220,In_61,In_533);
or U1221 (N_1221,In_911,In_572);
or U1222 (N_1222,In_660,In_896);
and U1223 (N_1223,In_521,In_924);
or U1224 (N_1224,In_718,In_33);
or U1225 (N_1225,In_315,In_41);
or U1226 (N_1226,In_563,In_4);
or U1227 (N_1227,In_769,In_996);
or U1228 (N_1228,In_852,In_178);
and U1229 (N_1229,In_955,In_527);
nor U1230 (N_1230,In_321,In_17);
and U1231 (N_1231,In_317,In_729);
nor U1232 (N_1232,In_58,In_968);
or U1233 (N_1233,In_886,In_106);
nand U1234 (N_1234,In_107,In_929);
nand U1235 (N_1235,In_524,In_744);
nor U1236 (N_1236,In_363,In_856);
or U1237 (N_1237,In_42,In_780);
xnor U1238 (N_1238,In_809,In_459);
or U1239 (N_1239,In_758,In_394);
xnor U1240 (N_1240,In_657,In_511);
and U1241 (N_1241,In_840,In_56);
nor U1242 (N_1242,In_416,In_926);
or U1243 (N_1243,In_962,In_613);
xnor U1244 (N_1244,In_824,In_121);
nor U1245 (N_1245,In_88,In_421);
and U1246 (N_1246,In_579,In_997);
or U1247 (N_1247,In_438,In_735);
nor U1248 (N_1248,In_398,In_38);
and U1249 (N_1249,In_172,In_731);
nand U1250 (N_1250,In_890,In_100);
xor U1251 (N_1251,In_582,In_5);
nor U1252 (N_1252,In_182,In_269);
or U1253 (N_1253,In_190,In_25);
nand U1254 (N_1254,In_508,In_35);
or U1255 (N_1255,In_774,In_792);
nand U1256 (N_1256,In_932,In_456);
nor U1257 (N_1257,In_154,In_554);
nor U1258 (N_1258,In_171,In_511);
xnor U1259 (N_1259,In_730,In_823);
or U1260 (N_1260,In_570,In_660);
xor U1261 (N_1261,In_193,In_814);
and U1262 (N_1262,In_112,In_11);
and U1263 (N_1263,In_641,In_98);
xnor U1264 (N_1264,In_977,In_463);
xnor U1265 (N_1265,In_488,In_819);
nand U1266 (N_1266,In_54,In_109);
xnor U1267 (N_1267,In_986,In_74);
nor U1268 (N_1268,In_455,In_918);
nand U1269 (N_1269,In_214,In_941);
nand U1270 (N_1270,In_323,In_534);
or U1271 (N_1271,In_189,In_880);
xor U1272 (N_1272,In_821,In_4);
nor U1273 (N_1273,In_528,In_746);
or U1274 (N_1274,In_784,In_584);
and U1275 (N_1275,In_964,In_182);
and U1276 (N_1276,In_587,In_823);
and U1277 (N_1277,In_475,In_248);
xnor U1278 (N_1278,In_525,In_621);
nand U1279 (N_1279,In_177,In_538);
nand U1280 (N_1280,In_50,In_175);
or U1281 (N_1281,In_623,In_249);
nand U1282 (N_1282,In_697,In_789);
and U1283 (N_1283,In_325,In_431);
or U1284 (N_1284,In_725,In_254);
or U1285 (N_1285,In_894,In_62);
or U1286 (N_1286,In_944,In_703);
nand U1287 (N_1287,In_965,In_345);
or U1288 (N_1288,In_277,In_618);
nor U1289 (N_1289,In_489,In_555);
nand U1290 (N_1290,In_891,In_382);
nand U1291 (N_1291,In_963,In_263);
or U1292 (N_1292,In_564,In_383);
and U1293 (N_1293,In_227,In_283);
nor U1294 (N_1294,In_513,In_284);
nand U1295 (N_1295,In_74,In_793);
xor U1296 (N_1296,In_148,In_829);
and U1297 (N_1297,In_272,In_335);
or U1298 (N_1298,In_288,In_542);
nand U1299 (N_1299,In_904,In_885);
and U1300 (N_1300,In_952,In_119);
nor U1301 (N_1301,In_991,In_787);
nand U1302 (N_1302,In_185,In_413);
or U1303 (N_1303,In_582,In_344);
nor U1304 (N_1304,In_477,In_319);
and U1305 (N_1305,In_798,In_656);
and U1306 (N_1306,In_883,In_55);
and U1307 (N_1307,In_109,In_97);
nand U1308 (N_1308,In_325,In_201);
nor U1309 (N_1309,In_675,In_422);
nand U1310 (N_1310,In_597,In_986);
xnor U1311 (N_1311,In_75,In_965);
and U1312 (N_1312,In_707,In_786);
nand U1313 (N_1313,In_68,In_899);
and U1314 (N_1314,In_36,In_212);
nor U1315 (N_1315,In_64,In_185);
xor U1316 (N_1316,In_793,In_216);
nor U1317 (N_1317,In_251,In_822);
nand U1318 (N_1318,In_837,In_43);
and U1319 (N_1319,In_651,In_186);
nand U1320 (N_1320,In_727,In_426);
or U1321 (N_1321,In_857,In_644);
nand U1322 (N_1322,In_695,In_524);
xnor U1323 (N_1323,In_719,In_864);
and U1324 (N_1324,In_961,In_185);
and U1325 (N_1325,In_796,In_379);
and U1326 (N_1326,In_8,In_246);
xor U1327 (N_1327,In_387,In_316);
xnor U1328 (N_1328,In_662,In_780);
nor U1329 (N_1329,In_16,In_27);
or U1330 (N_1330,In_80,In_889);
nor U1331 (N_1331,In_227,In_584);
or U1332 (N_1332,In_898,In_895);
nand U1333 (N_1333,In_604,In_338);
nand U1334 (N_1334,In_694,In_99);
and U1335 (N_1335,In_389,In_998);
xnor U1336 (N_1336,In_321,In_162);
nor U1337 (N_1337,In_675,In_103);
and U1338 (N_1338,In_598,In_828);
or U1339 (N_1339,In_815,In_156);
or U1340 (N_1340,In_348,In_706);
nor U1341 (N_1341,In_92,In_110);
nand U1342 (N_1342,In_935,In_393);
and U1343 (N_1343,In_750,In_310);
nand U1344 (N_1344,In_907,In_957);
nor U1345 (N_1345,In_182,In_566);
xnor U1346 (N_1346,In_381,In_472);
or U1347 (N_1347,In_489,In_990);
xor U1348 (N_1348,In_886,In_578);
nand U1349 (N_1349,In_87,In_903);
nand U1350 (N_1350,In_675,In_471);
and U1351 (N_1351,In_360,In_293);
or U1352 (N_1352,In_735,In_215);
nand U1353 (N_1353,In_696,In_178);
nor U1354 (N_1354,In_181,In_165);
xor U1355 (N_1355,In_921,In_949);
or U1356 (N_1356,In_755,In_388);
nor U1357 (N_1357,In_15,In_723);
xor U1358 (N_1358,In_556,In_672);
xnor U1359 (N_1359,In_456,In_291);
xnor U1360 (N_1360,In_787,In_317);
xnor U1361 (N_1361,In_575,In_817);
nor U1362 (N_1362,In_860,In_1);
nand U1363 (N_1363,In_698,In_687);
and U1364 (N_1364,In_548,In_288);
xnor U1365 (N_1365,In_393,In_743);
nand U1366 (N_1366,In_227,In_247);
nand U1367 (N_1367,In_21,In_973);
xor U1368 (N_1368,In_511,In_996);
nor U1369 (N_1369,In_514,In_566);
and U1370 (N_1370,In_638,In_167);
nand U1371 (N_1371,In_201,In_333);
and U1372 (N_1372,In_123,In_175);
or U1373 (N_1373,In_202,In_15);
or U1374 (N_1374,In_537,In_447);
nor U1375 (N_1375,In_851,In_27);
or U1376 (N_1376,In_304,In_119);
nor U1377 (N_1377,In_219,In_253);
xnor U1378 (N_1378,In_505,In_856);
nand U1379 (N_1379,In_701,In_993);
xor U1380 (N_1380,In_603,In_615);
or U1381 (N_1381,In_138,In_338);
or U1382 (N_1382,In_576,In_958);
nor U1383 (N_1383,In_977,In_508);
or U1384 (N_1384,In_959,In_992);
and U1385 (N_1385,In_161,In_631);
nand U1386 (N_1386,In_399,In_963);
nand U1387 (N_1387,In_203,In_546);
xor U1388 (N_1388,In_451,In_847);
xnor U1389 (N_1389,In_447,In_453);
or U1390 (N_1390,In_762,In_414);
xor U1391 (N_1391,In_2,In_499);
nor U1392 (N_1392,In_254,In_406);
xnor U1393 (N_1393,In_267,In_977);
or U1394 (N_1394,In_642,In_927);
or U1395 (N_1395,In_271,In_858);
or U1396 (N_1396,In_154,In_784);
or U1397 (N_1397,In_685,In_968);
and U1398 (N_1398,In_371,In_574);
xnor U1399 (N_1399,In_725,In_865);
nor U1400 (N_1400,In_377,In_974);
and U1401 (N_1401,In_45,In_798);
xor U1402 (N_1402,In_964,In_160);
nand U1403 (N_1403,In_757,In_794);
nor U1404 (N_1404,In_31,In_353);
nand U1405 (N_1405,In_750,In_864);
and U1406 (N_1406,In_186,In_216);
or U1407 (N_1407,In_659,In_412);
nand U1408 (N_1408,In_918,In_1);
xnor U1409 (N_1409,In_505,In_87);
nand U1410 (N_1410,In_826,In_795);
nand U1411 (N_1411,In_626,In_772);
nor U1412 (N_1412,In_533,In_767);
and U1413 (N_1413,In_560,In_792);
or U1414 (N_1414,In_21,In_62);
and U1415 (N_1415,In_471,In_720);
nand U1416 (N_1416,In_240,In_604);
nand U1417 (N_1417,In_801,In_280);
or U1418 (N_1418,In_491,In_484);
xor U1419 (N_1419,In_878,In_372);
or U1420 (N_1420,In_763,In_420);
xor U1421 (N_1421,In_82,In_315);
or U1422 (N_1422,In_673,In_854);
and U1423 (N_1423,In_20,In_194);
nand U1424 (N_1424,In_94,In_574);
nand U1425 (N_1425,In_701,In_566);
nand U1426 (N_1426,In_837,In_789);
and U1427 (N_1427,In_715,In_459);
and U1428 (N_1428,In_188,In_10);
xnor U1429 (N_1429,In_28,In_226);
nand U1430 (N_1430,In_769,In_983);
nand U1431 (N_1431,In_960,In_841);
and U1432 (N_1432,In_354,In_683);
xor U1433 (N_1433,In_585,In_898);
nand U1434 (N_1434,In_773,In_893);
and U1435 (N_1435,In_827,In_598);
and U1436 (N_1436,In_32,In_694);
or U1437 (N_1437,In_738,In_544);
and U1438 (N_1438,In_224,In_24);
or U1439 (N_1439,In_209,In_883);
or U1440 (N_1440,In_53,In_967);
xor U1441 (N_1441,In_756,In_903);
xor U1442 (N_1442,In_537,In_162);
xnor U1443 (N_1443,In_725,In_645);
or U1444 (N_1444,In_531,In_1);
nand U1445 (N_1445,In_69,In_612);
xor U1446 (N_1446,In_874,In_828);
nor U1447 (N_1447,In_833,In_35);
or U1448 (N_1448,In_215,In_153);
nor U1449 (N_1449,In_305,In_785);
xnor U1450 (N_1450,In_501,In_613);
and U1451 (N_1451,In_70,In_160);
and U1452 (N_1452,In_82,In_640);
nor U1453 (N_1453,In_923,In_727);
or U1454 (N_1454,In_288,In_14);
nor U1455 (N_1455,In_956,In_647);
nor U1456 (N_1456,In_568,In_884);
nor U1457 (N_1457,In_287,In_489);
or U1458 (N_1458,In_946,In_735);
nand U1459 (N_1459,In_326,In_740);
or U1460 (N_1460,In_764,In_323);
or U1461 (N_1461,In_661,In_433);
or U1462 (N_1462,In_454,In_743);
or U1463 (N_1463,In_714,In_382);
nand U1464 (N_1464,In_184,In_887);
or U1465 (N_1465,In_197,In_547);
nand U1466 (N_1466,In_311,In_194);
or U1467 (N_1467,In_184,In_292);
or U1468 (N_1468,In_443,In_460);
nand U1469 (N_1469,In_161,In_199);
and U1470 (N_1470,In_407,In_517);
and U1471 (N_1471,In_823,In_496);
nand U1472 (N_1472,In_377,In_944);
nor U1473 (N_1473,In_686,In_154);
xor U1474 (N_1474,In_802,In_376);
nand U1475 (N_1475,In_256,In_81);
nand U1476 (N_1476,In_298,In_825);
nand U1477 (N_1477,In_356,In_200);
nand U1478 (N_1478,In_290,In_845);
and U1479 (N_1479,In_919,In_930);
nor U1480 (N_1480,In_584,In_666);
nand U1481 (N_1481,In_429,In_603);
or U1482 (N_1482,In_227,In_332);
nand U1483 (N_1483,In_683,In_801);
xor U1484 (N_1484,In_486,In_283);
and U1485 (N_1485,In_122,In_474);
or U1486 (N_1486,In_475,In_741);
and U1487 (N_1487,In_800,In_719);
nor U1488 (N_1488,In_214,In_180);
nor U1489 (N_1489,In_870,In_793);
and U1490 (N_1490,In_751,In_358);
xor U1491 (N_1491,In_91,In_168);
and U1492 (N_1492,In_126,In_799);
or U1493 (N_1493,In_190,In_284);
and U1494 (N_1494,In_216,In_293);
xor U1495 (N_1495,In_276,In_745);
nand U1496 (N_1496,In_556,In_834);
and U1497 (N_1497,In_992,In_424);
xor U1498 (N_1498,In_863,In_239);
or U1499 (N_1499,In_649,In_744);
xor U1500 (N_1500,In_496,In_44);
nand U1501 (N_1501,In_992,In_292);
xor U1502 (N_1502,In_130,In_894);
nand U1503 (N_1503,In_14,In_120);
nor U1504 (N_1504,In_929,In_39);
or U1505 (N_1505,In_784,In_414);
nand U1506 (N_1506,In_135,In_215);
xor U1507 (N_1507,In_155,In_629);
and U1508 (N_1508,In_943,In_346);
xnor U1509 (N_1509,In_449,In_73);
xnor U1510 (N_1510,In_911,In_463);
and U1511 (N_1511,In_188,In_892);
nor U1512 (N_1512,In_52,In_188);
xor U1513 (N_1513,In_661,In_868);
or U1514 (N_1514,In_280,In_829);
xnor U1515 (N_1515,In_801,In_723);
xor U1516 (N_1516,In_395,In_486);
nand U1517 (N_1517,In_556,In_414);
or U1518 (N_1518,In_372,In_62);
xnor U1519 (N_1519,In_713,In_126);
or U1520 (N_1520,In_422,In_279);
or U1521 (N_1521,In_699,In_30);
xor U1522 (N_1522,In_668,In_504);
or U1523 (N_1523,In_90,In_185);
nand U1524 (N_1524,In_306,In_395);
or U1525 (N_1525,In_710,In_169);
nor U1526 (N_1526,In_108,In_710);
and U1527 (N_1527,In_99,In_296);
and U1528 (N_1528,In_435,In_240);
nor U1529 (N_1529,In_769,In_165);
or U1530 (N_1530,In_243,In_954);
nand U1531 (N_1531,In_629,In_592);
xnor U1532 (N_1532,In_897,In_164);
or U1533 (N_1533,In_493,In_380);
xnor U1534 (N_1534,In_241,In_501);
and U1535 (N_1535,In_484,In_620);
nand U1536 (N_1536,In_553,In_467);
or U1537 (N_1537,In_654,In_266);
nor U1538 (N_1538,In_629,In_640);
and U1539 (N_1539,In_742,In_108);
nor U1540 (N_1540,In_7,In_461);
nand U1541 (N_1541,In_896,In_766);
nor U1542 (N_1542,In_128,In_996);
and U1543 (N_1543,In_52,In_605);
or U1544 (N_1544,In_443,In_553);
or U1545 (N_1545,In_97,In_687);
nand U1546 (N_1546,In_538,In_730);
nor U1547 (N_1547,In_598,In_469);
or U1548 (N_1548,In_762,In_775);
nor U1549 (N_1549,In_989,In_276);
nor U1550 (N_1550,In_436,In_872);
or U1551 (N_1551,In_52,In_788);
nand U1552 (N_1552,In_155,In_909);
xor U1553 (N_1553,In_844,In_825);
xnor U1554 (N_1554,In_554,In_381);
nand U1555 (N_1555,In_13,In_536);
and U1556 (N_1556,In_488,In_503);
nor U1557 (N_1557,In_976,In_727);
nand U1558 (N_1558,In_140,In_330);
and U1559 (N_1559,In_233,In_558);
and U1560 (N_1560,In_256,In_770);
or U1561 (N_1561,In_795,In_745);
nand U1562 (N_1562,In_456,In_785);
or U1563 (N_1563,In_11,In_628);
or U1564 (N_1564,In_188,In_915);
xnor U1565 (N_1565,In_334,In_521);
nor U1566 (N_1566,In_890,In_877);
nor U1567 (N_1567,In_538,In_281);
xor U1568 (N_1568,In_538,In_124);
nand U1569 (N_1569,In_936,In_458);
and U1570 (N_1570,In_480,In_390);
nor U1571 (N_1571,In_260,In_747);
nand U1572 (N_1572,In_0,In_952);
or U1573 (N_1573,In_579,In_749);
nor U1574 (N_1574,In_266,In_255);
or U1575 (N_1575,In_505,In_109);
xor U1576 (N_1576,In_919,In_541);
xnor U1577 (N_1577,In_525,In_696);
xnor U1578 (N_1578,In_718,In_748);
xnor U1579 (N_1579,In_190,In_954);
and U1580 (N_1580,In_420,In_327);
nor U1581 (N_1581,In_802,In_152);
xnor U1582 (N_1582,In_281,In_408);
nand U1583 (N_1583,In_852,In_253);
nand U1584 (N_1584,In_602,In_938);
or U1585 (N_1585,In_371,In_529);
and U1586 (N_1586,In_836,In_411);
nand U1587 (N_1587,In_259,In_519);
and U1588 (N_1588,In_490,In_103);
xor U1589 (N_1589,In_338,In_297);
and U1590 (N_1590,In_404,In_844);
xnor U1591 (N_1591,In_348,In_535);
or U1592 (N_1592,In_500,In_982);
or U1593 (N_1593,In_80,In_372);
xor U1594 (N_1594,In_82,In_91);
nor U1595 (N_1595,In_944,In_478);
or U1596 (N_1596,In_453,In_765);
xnor U1597 (N_1597,In_64,In_45);
xnor U1598 (N_1598,In_258,In_569);
and U1599 (N_1599,In_307,In_198);
xnor U1600 (N_1600,In_697,In_514);
nand U1601 (N_1601,In_598,In_399);
xnor U1602 (N_1602,In_145,In_890);
nor U1603 (N_1603,In_2,In_61);
xor U1604 (N_1604,In_424,In_574);
or U1605 (N_1605,In_612,In_353);
and U1606 (N_1606,In_720,In_899);
or U1607 (N_1607,In_764,In_986);
xor U1608 (N_1608,In_309,In_149);
and U1609 (N_1609,In_369,In_249);
nand U1610 (N_1610,In_896,In_0);
nor U1611 (N_1611,In_891,In_538);
and U1612 (N_1612,In_672,In_110);
nand U1613 (N_1613,In_719,In_162);
nand U1614 (N_1614,In_327,In_530);
xor U1615 (N_1615,In_890,In_456);
nand U1616 (N_1616,In_9,In_357);
and U1617 (N_1617,In_271,In_181);
or U1618 (N_1618,In_299,In_288);
and U1619 (N_1619,In_229,In_868);
nor U1620 (N_1620,In_689,In_108);
nand U1621 (N_1621,In_750,In_853);
nor U1622 (N_1622,In_173,In_568);
nor U1623 (N_1623,In_186,In_100);
and U1624 (N_1624,In_35,In_511);
or U1625 (N_1625,In_985,In_184);
nand U1626 (N_1626,In_940,In_726);
xor U1627 (N_1627,In_55,In_864);
nand U1628 (N_1628,In_105,In_317);
xor U1629 (N_1629,In_58,In_771);
xnor U1630 (N_1630,In_292,In_860);
or U1631 (N_1631,In_948,In_747);
or U1632 (N_1632,In_57,In_534);
nand U1633 (N_1633,In_500,In_563);
nor U1634 (N_1634,In_999,In_605);
or U1635 (N_1635,In_648,In_288);
xor U1636 (N_1636,In_778,In_306);
nor U1637 (N_1637,In_437,In_851);
nor U1638 (N_1638,In_188,In_755);
or U1639 (N_1639,In_178,In_793);
nand U1640 (N_1640,In_754,In_811);
nand U1641 (N_1641,In_786,In_863);
xor U1642 (N_1642,In_223,In_901);
nor U1643 (N_1643,In_897,In_491);
or U1644 (N_1644,In_818,In_558);
or U1645 (N_1645,In_587,In_151);
xnor U1646 (N_1646,In_780,In_314);
nor U1647 (N_1647,In_854,In_33);
and U1648 (N_1648,In_898,In_304);
nor U1649 (N_1649,In_473,In_749);
xnor U1650 (N_1650,In_493,In_668);
and U1651 (N_1651,In_736,In_76);
xor U1652 (N_1652,In_641,In_288);
or U1653 (N_1653,In_355,In_303);
xor U1654 (N_1654,In_694,In_735);
nor U1655 (N_1655,In_465,In_65);
xnor U1656 (N_1656,In_36,In_602);
and U1657 (N_1657,In_917,In_988);
xor U1658 (N_1658,In_634,In_459);
and U1659 (N_1659,In_200,In_628);
nand U1660 (N_1660,In_275,In_536);
nand U1661 (N_1661,In_329,In_874);
and U1662 (N_1662,In_450,In_946);
and U1663 (N_1663,In_529,In_346);
xnor U1664 (N_1664,In_21,In_3);
nor U1665 (N_1665,In_761,In_803);
or U1666 (N_1666,In_962,In_688);
xnor U1667 (N_1667,In_508,In_491);
xor U1668 (N_1668,In_816,In_814);
nor U1669 (N_1669,In_126,In_581);
xor U1670 (N_1670,In_213,In_408);
nand U1671 (N_1671,In_88,In_309);
nand U1672 (N_1672,In_383,In_810);
nor U1673 (N_1673,In_276,In_458);
or U1674 (N_1674,In_269,In_903);
xnor U1675 (N_1675,In_30,In_540);
nand U1676 (N_1676,In_533,In_812);
nand U1677 (N_1677,In_397,In_338);
nor U1678 (N_1678,In_905,In_179);
and U1679 (N_1679,In_739,In_709);
nor U1680 (N_1680,In_200,In_497);
or U1681 (N_1681,In_828,In_28);
nor U1682 (N_1682,In_856,In_106);
nor U1683 (N_1683,In_317,In_767);
xnor U1684 (N_1684,In_777,In_283);
nand U1685 (N_1685,In_573,In_45);
nand U1686 (N_1686,In_99,In_149);
nor U1687 (N_1687,In_785,In_340);
nand U1688 (N_1688,In_511,In_587);
xnor U1689 (N_1689,In_751,In_659);
or U1690 (N_1690,In_391,In_835);
nor U1691 (N_1691,In_240,In_756);
xnor U1692 (N_1692,In_685,In_221);
nor U1693 (N_1693,In_734,In_398);
nand U1694 (N_1694,In_391,In_149);
or U1695 (N_1695,In_199,In_953);
and U1696 (N_1696,In_68,In_589);
nor U1697 (N_1697,In_41,In_745);
xnor U1698 (N_1698,In_734,In_847);
and U1699 (N_1699,In_954,In_225);
or U1700 (N_1700,In_294,In_462);
xor U1701 (N_1701,In_922,In_411);
xnor U1702 (N_1702,In_777,In_730);
and U1703 (N_1703,In_811,In_664);
and U1704 (N_1704,In_367,In_679);
xor U1705 (N_1705,In_158,In_590);
nand U1706 (N_1706,In_818,In_713);
nand U1707 (N_1707,In_553,In_496);
or U1708 (N_1708,In_628,In_455);
xor U1709 (N_1709,In_207,In_615);
nand U1710 (N_1710,In_478,In_2);
nor U1711 (N_1711,In_867,In_828);
nor U1712 (N_1712,In_541,In_78);
and U1713 (N_1713,In_503,In_956);
xnor U1714 (N_1714,In_87,In_336);
and U1715 (N_1715,In_5,In_23);
xnor U1716 (N_1716,In_890,In_983);
nor U1717 (N_1717,In_131,In_402);
or U1718 (N_1718,In_707,In_773);
or U1719 (N_1719,In_179,In_263);
or U1720 (N_1720,In_313,In_438);
xnor U1721 (N_1721,In_176,In_863);
nor U1722 (N_1722,In_213,In_987);
or U1723 (N_1723,In_40,In_570);
and U1724 (N_1724,In_230,In_176);
nand U1725 (N_1725,In_93,In_249);
xnor U1726 (N_1726,In_420,In_496);
or U1727 (N_1727,In_208,In_453);
nor U1728 (N_1728,In_976,In_323);
and U1729 (N_1729,In_407,In_571);
and U1730 (N_1730,In_526,In_495);
nand U1731 (N_1731,In_543,In_265);
xor U1732 (N_1732,In_629,In_311);
nand U1733 (N_1733,In_174,In_673);
nand U1734 (N_1734,In_323,In_896);
and U1735 (N_1735,In_403,In_755);
or U1736 (N_1736,In_283,In_45);
xnor U1737 (N_1737,In_516,In_935);
or U1738 (N_1738,In_840,In_674);
nand U1739 (N_1739,In_290,In_438);
xnor U1740 (N_1740,In_124,In_682);
and U1741 (N_1741,In_472,In_226);
or U1742 (N_1742,In_205,In_94);
and U1743 (N_1743,In_747,In_113);
or U1744 (N_1744,In_203,In_127);
nor U1745 (N_1745,In_807,In_114);
and U1746 (N_1746,In_93,In_773);
xor U1747 (N_1747,In_755,In_669);
nor U1748 (N_1748,In_851,In_269);
nor U1749 (N_1749,In_277,In_556);
or U1750 (N_1750,In_136,In_150);
or U1751 (N_1751,In_429,In_370);
and U1752 (N_1752,In_410,In_280);
xor U1753 (N_1753,In_147,In_882);
or U1754 (N_1754,In_671,In_732);
nor U1755 (N_1755,In_797,In_381);
or U1756 (N_1756,In_95,In_683);
nor U1757 (N_1757,In_893,In_77);
nor U1758 (N_1758,In_941,In_274);
or U1759 (N_1759,In_93,In_99);
nand U1760 (N_1760,In_732,In_986);
xnor U1761 (N_1761,In_616,In_20);
nand U1762 (N_1762,In_482,In_623);
xnor U1763 (N_1763,In_563,In_3);
xor U1764 (N_1764,In_453,In_235);
nor U1765 (N_1765,In_128,In_316);
and U1766 (N_1766,In_223,In_624);
xnor U1767 (N_1767,In_975,In_488);
and U1768 (N_1768,In_880,In_550);
xnor U1769 (N_1769,In_377,In_169);
nor U1770 (N_1770,In_117,In_272);
nor U1771 (N_1771,In_729,In_239);
or U1772 (N_1772,In_15,In_545);
or U1773 (N_1773,In_148,In_201);
xnor U1774 (N_1774,In_611,In_841);
and U1775 (N_1775,In_981,In_884);
or U1776 (N_1776,In_25,In_412);
xnor U1777 (N_1777,In_429,In_889);
or U1778 (N_1778,In_959,In_770);
nand U1779 (N_1779,In_52,In_428);
nand U1780 (N_1780,In_629,In_120);
xor U1781 (N_1781,In_152,In_46);
xnor U1782 (N_1782,In_310,In_153);
xor U1783 (N_1783,In_469,In_76);
and U1784 (N_1784,In_427,In_528);
nand U1785 (N_1785,In_827,In_211);
nor U1786 (N_1786,In_126,In_715);
or U1787 (N_1787,In_835,In_520);
nor U1788 (N_1788,In_280,In_151);
or U1789 (N_1789,In_86,In_650);
nor U1790 (N_1790,In_990,In_553);
nor U1791 (N_1791,In_223,In_683);
and U1792 (N_1792,In_878,In_765);
and U1793 (N_1793,In_280,In_919);
nand U1794 (N_1794,In_516,In_375);
nor U1795 (N_1795,In_631,In_978);
xnor U1796 (N_1796,In_644,In_501);
and U1797 (N_1797,In_21,In_587);
or U1798 (N_1798,In_384,In_625);
nor U1799 (N_1799,In_135,In_372);
nor U1800 (N_1800,In_835,In_142);
or U1801 (N_1801,In_921,In_342);
nor U1802 (N_1802,In_202,In_513);
and U1803 (N_1803,In_578,In_607);
and U1804 (N_1804,In_486,In_893);
xor U1805 (N_1805,In_701,In_480);
and U1806 (N_1806,In_27,In_891);
or U1807 (N_1807,In_783,In_348);
nand U1808 (N_1808,In_83,In_680);
and U1809 (N_1809,In_839,In_429);
nand U1810 (N_1810,In_127,In_270);
nor U1811 (N_1811,In_551,In_500);
or U1812 (N_1812,In_747,In_188);
or U1813 (N_1813,In_989,In_551);
or U1814 (N_1814,In_845,In_198);
nor U1815 (N_1815,In_401,In_701);
or U1816 (N_1816,In_17,In_604);
or U1817 (N_1817,In_426,In_510);
and U1818 (N_1818,In_418,In_256);
and U1819 (N_1819,In_120,In_732);
nor U1820 (N_1820,In_214,In_250);
nor U1821 (N_1821,In_739,In_496);
nand U1822 (N_1822,In_33,In_327);
or U1823 (N_1823,In_248,In_596);
nor U1824 (N_1824,In_332,In_516);
and U1825 (N_1825,In_515,In_684);
or U1826 (N_1826,In_440,In_436);
nand U1827 (N_1827,In_330,In_918);
nor U1828 (N_1828,In_18,In_564);
nand U1829 (N_1829,In_465,In_289);
xor U1830 (N_1830,In_563,In_456);
nand U1831 (N_1831,In_474,In_712);
nand U1832 (N_1832,In_660,In_796);
and U1833 (N_1833,In_289,In_280);
and U1834 (N_1834,In_902,In_312);
or U1835 (N_1835,In_712,In_546);
and U1836 (N_1836,In_163,In_40);
nor U1837 (N_1837,In_917,In_49);
nand U1838 (N_1838,In_478,In_311);
nor U1839 (N_1839,In_130,In_191);
and U1840 (N_1840,In_885,In_196);
nor U1841 (N_1841,In_480,In_393);
or U1842 (N_1842,In_19,In_963);
nor U1843 (N_1843,In_620,In_17);
xor U1844 (N_1844,In_242,In_179);
or U1845 (N_1845,In_503,In_374);
nand U1846 (N_1846,In_699,In_302);
nor U1847 (N_1847,In_315,In_296);
or U1848 (N_1848,In_386,In_497);
xnor U1849 (N_1849,In_168,In_620);
xnor U1850 (N_1850,In_578,In_203);
or U1851 (N_1851,In_844,In_483);
nor U1852 (N_1852,In_14,In_950);
nand U1853 (N_1853,In_657,In_949);
nor U1854 (N_1854,In_268,In_575);
nand U1855 (N_1855,In_867,In_308);
xnor U1856 (N_1856,In_231,In_741);
or U1857 (N_1857,In_713,In_379);
nand U1858 (N_1858,In_928,In_494);
or U1859 (N_1859,In_568,In_408);
nand U1860 (N_1860,In_49,In_264);
nand U1861 (N_1861,In_889,In_690);
and U1862 (N_1862,In_290,In_305);
xnor U1863 (N_1863,In_443,In_717);
or U1864 (N_1864,In_326,In_290);
nor U1865 (N_1865,In_381,In_225);
xnor U1866 (N_1866,In_543,In_254);
nor U1867 (N_1867,In_947,In_43);
or U1868 (N_1868,In_827,In_453);
or U1869 (N_1869,In_744,In_955);
xnor U1870 (N_1870,In_161,In_344);
nand U1871 (N_1871,In_213,In_300);
nor U1872 (N_1872,In_580,In_320);
nor U1873 (N_1873,In_589,In_801);
xor U1874 (N_1874,In_914,In_481);
nor U1875 (N_1875,In_505,In_687);
and U1876 (N_1876,In_369,In_985);
xor U1877 (N_1877,In_318,In_427);
and U1878 (N_1878,In_936,In_256);
or U1879 (N_1879,In_683,In_856);
or U1880 (N_1880,In_324,In_806);
xor U1881 (N_1881,In_318,In_957);
or U1882 (N_1882,In_797,In_271);
or U1883 (N_1883,In_72,In_895);
nand U1884 (N_1884,In_896,In_139);
or U1885 (N_1885,In_713,In_994);
nand U1886 (N_1886,In_862,In_735);
and U1887 (N_1887,In_747,In_371);
xor U1888 (N_1888,In_249,In_733);
or U1889 (N_1889,In_363,In_447);
or U1890 (N_1890,In_390,In_570);
or U1891 (N_1891,In_510,In_631);
nor U1892 (N_1892,In_837,In_987);
nor U1893 (N_1893,In_42,In_629);
nand U1894 (N_1894,In_762,In_780);
nand U1895 (N_1895,In_224,In_510);
nor U1896 (N_1896,In_364,In_735);
nor U1897 (N_1897,In_963,In_994);
and U1898 (N_1898,In_944,In_421);
nand U1899 (N_1899,In_134,In_330);
nand U1900 (N_1900,In_462,In_539);
nand U1901 (N_1901,In_97,In_117);
nor U1902 (N_1902,In_199,In_852);
xor U1903 (N_1903,In_147,In_788);
xnor U1904 (N_1904,In_703,In_553);
nand U1905 (N_1905,In_551,In_353);
or U1906 (N_1906,In_390,In_415);
nand U1907 (N_1907,In_990,In_788);
xor U1908 (N_1908,In_736,In_302);
nor U1909 (N_1909,In_228,In_427);
xnor U1910 (N_1910,In_142,In_561);
or U1911 (N_1911,In_346,In_474);
nand U1912 (N_1912,In_911,In_929);
and U1913 (N_1913,In_795,In_849);
xnor U1914 (N_1914,In_658,In_520);
nor U1915 (N_1915,In_172,In_353);
nand U1916 (N_1916,In_651,In_537);
and U1917 (N_1917,In_945,In_243);
xor U1918 (N_1918,In_968,In_71);
and U1919 (N_1919,In_392,In_142);
nor U1920 (N_1920,In_158,In_639);
and U1921 (N_1921,In_19,In_918);
and U1922 (N_1922,In_678,In_489);
nand U1923 (N_1923,In_70,In_867);
xor U1924 (N_1924,In_233,In_436);
or U1925 (N_1925,In_431,In_918);
or U1926 (N_1926,In_575,In_255);
nand U1927 (N_1927,In_526,In_428);
nand U1928 (N_1928,In_75,In_882);
xor U1929 (N_1929,In_33,In_499);
nand U1930 (N_1930,In_985,In_78);
nand U1931 (N_1931,In_46,In_632);
nand U1932 (N_1932,In_814,In_738);
and U1933 (N_1933,In_669,In_44);
or U1934 (N_1934,In_36,In_607);
nand U1935 (N_1935,In_291,In_949);
or U1936 (N_1936,In_65,In_208);
xor U1937 (N_1937,In_69,In_321);
nor U1938 (N_1938,In_581,In_425);
nor U1939 (N_1939,In_850,In_678);
nor U1940 (N_1940,In_151,In_692);
nor U1941 (N_1941,In_471,In_759);
and U1942 (N_1942,In_22,In_23);
xor U1943 (N_1943,In_223,In_784);
or U1944 (N_1944,In_973,In_194);
and U1945 (N_1945,In_783,In_986);
nand U1946 (N_1946,In_941,In_891);
and U1947 (N_1947,In_636,In_934);
or U1948 (N_1948,In_438,In_743);
nand U1949 (N_1949,In_712,In_176);
nand U1950 (N_1950,In_955,In_923);
nor U1951 (N_1951,In_124,In_100);
xor U1952 (N_1952,In_744,In_992);
and U1953 (N_1953,In_198,In_151);
or U1954 (N_1954,In_481,In_493);
nor U1955 (N_1955,In_888,In_79);
or U1956 (N_1956,In_131,In_696);
xor U1957 (N_1957,In_278,In_814);
or U1958 (N_1958,In_356,In_220);
nor U1959 (N_1959,In_916,In_310);
nor U1960 (N_1960,In_702,In_147);
nand U1961 (N_1961,In_51,In_83);
or U1962 (N_1962,In_839,In_417);
nand U1963 (N_1963,In_538,In_887);
xnor U1964 (N_1964,In_311,In_734);
xnor U1965 (N_1965,In_27,In_769);
and U1966 (N_1966,In_108,In_926);
and U1967 (N_1967,In_894,In_607);
nand U1968 (N_1968,In_705,In_373);
nor U1969 (N_1969,In_884,In_918);
or U1970 (N_1970,In_470,In_81);
and U1971 (N_1971,In_463,In_479);
nand U1972 (N_1972,In_917,In_417);
nor U1973 (N_1973,In_572,In_103);
nor U1974 (N_1974,In_558,In_971);
nor U1975 (N_1975,In_932,In_897);
and U1976 (N_1976,In_818,In_290);
nand U1977 (N_1977,In_670,In_815);
xnor U1978 (N_1978,In_388,In_144);
and U1979 (N_1979,In_945,In_141);
nand U1980 (N_1980,In_959,In_895);
xnor U1981 (N_1981,In_18,In_750);
and U1982 (N_1982,In_305,In_486);
and U1983 (N_1983,In_37,In_187);
xor U1984 (N_1984,In_985,In_165);
and U1985 (N_1985,In_378,In_554);
xor U1986 (N_1986,In_115,In_94);
and U1987 (N_1987,In_141,In_793);
nor U1988 (N_1988,In_777,In_646);
and U1989 (N_1989,In_52,In_589);
xnor U1990 (N_1990,In_343,In_862);
nor U1991 (N_1991,In_909,In_921);
nand U1992 (N_1992,In_996,In_292);
nand U1993 (N_1993,In_736,In_951);
and U1994 (N_1994,In_55,In_98);
xor U1995 (N_1995,In_321,In_135);
xor U1996 (N_1996,In_109,In_251);
and U1997 (N_1997,In_600,In_570);
or U1998 (N_1998,In_894,In_710);
nor U1999 (N_1999,In_325,In_429);
nor U2000 (N_2000,In_269,In_147);
nor U2001 (N_2001,In_460,In_52);
and U2002 (N_2002,In_966,In_765);
nand U2003 (N_2003,In_487,In_407);
and U2004 (N_2004,In_75,In_964);
xnor U2005 (N_2005,In_181,In_924);
and U2006 (N_2006,In_802,In_912);
or U2007 (N_2007,In_360,In_412);
and U2008 (N_2008,In_54,In_331);
and U2009 (N_2009,In_195,In_436);
nand U2010 (N_2010,In_696,In_997);
xor U2011 (N_2011,In_802,In_202);
xor U2012 (N_2012,In_458,In_644);
xnor U2013 (N_2013,In_639,In_748);
nor U2014 (N_2014,In_923,In_720);
or U2015 (N_2015,In_606,In_123);
xnor U2016 (N_2016,In_520,In_341);
or U2017 (N_2017,In_293,In_656);
xnor U2018 (N_2018,In_457,In_80);
nand U2019 (N_2019,In_362,In_65);
and U2020 (N_2020,In_915,In_385);
xnor U2021 (N_2021,In_716,In_866);
xor U2022 (N_2022,In_749,In_373);
nor U2023 (N_2023,In_221,In_156);
nor U2024 (N_2024,In_3,In_931);
xnor U2025 (N_2025,In_488,In_221);
xnor U2026 (N_2026,In_429,In_101);
xor U2027 (N_2027,In_719,In_650);
nor U2028 (N_2028,In_187,In_512);
xor U2029 (N_2029,In_540,In_777);
xor U2030 (N_2030,In_823,In_613);
nor U2031 (N_2031,In_679,In_615);
and U2032 (N_2032,In_291,In_630);
xor U2033 (N_2033,In_471,In_890);
and U2034 (N_2034,In_290,In_834);
nand U2035 (N_2035,In_841,In_185);
and U2036 (N_2036,In_482,In_496);
nand U2037 (N_2037,In_748,In_83);
nor U2038 (N_2038,In_823,In_114);
nor U2039 (N_2039,In_792,In_892);
nand U2040 (N_2040,In_677,In_138);
and U2041 (N_2041,In_277,In_30);
xnor U2042 (N_2042,In_420,In_60);
nor U2043 (N_2043,In_746,In_236);
nand U2044 (N_2044,In_112,In_204);
or U2045 (N_2045,In_974,In_957);
nand U2046 (N_2046,In_817,In_360);
nand U2047 (N_2047,In_100,In_235);
nand U2048 (N_2048,In_879,In_448);
nor U2049 (N_2049,In_295,In_631);
and U2050 (N_2050,In_223,In_857);
and U2051 (N_2051,In_245,In_93);
or U2052 (N_2052,In_606,In_259);
nor U2053 (N_2053,In_114,In_124);
nand U2054 (N_2054,In_945,In_651);
nor U2055 (N_2055,In_885,In_698);
nor U2056 (N_2056,In_274,In_338);
nor U2057 (N_2057,In_645,In_482);
and U2058 (N_2058,In_477,In_788);
xor U2059 (N_2059,In_527,In_650);
or U2060 (N_2060,In_24,In_491);
nand U2061 (N_2061,In_912,In_326);
and U2062 (N_2062,In_284,In_113);
nor U2063 (N_2063,In_715,In_39);
xnor U2064 (N_2064,In_525,In_695);
nor U2065 (N_2065,In_484,In_371);
nand U2066 (N_2066,In_175,In_310);
nand U2067 (N_2067,In_889,In_417);
nand U2068 (N_2068,In_80,In_770);
xnor U2069 (N_2069,In_246,In_870);
and U2070 (N_2070,In_723,In_168);
nor U2071 (N_2071,In_792,In_990);
nand U2072 (N_2072,In_933,In_757);
and U2073 (N_2073,In_37,In_633);
xor U2074 (N_2074,In_458,In_438);
nand U2075 (N_2075,In_340,In_571);
xor U2076 (N_2076,In_991,In_561);
xor U2077 (N_2077,In_108,In_370);
and U2078 (N_2078,In_548,In_332);
and U2079 (N_2079,In_332,In_426);
nor U2080 (N_2080,In_788,In_55);
or U2081 (N_2081,In_578,In_966);
nor U2082 (N_2082,In_729,In_715);
nor U2083 (N_2083,In_573,In_475);
xor U2084 (N_2084,In_315,In_126);
xnor U2085 (N_2085,In_877,In_511);
nand U2086 (N_2086,In_127,In_271);
nand U2087 (N_2087,In_965,In_751);
xnor U2088 (N_2088,In_286,In_134);
nor U2089 (N_2089,In_409,In_269);
xor U2090 (N_2090,In_531,In_676);
and U2091 (N_2091,In_113,In_37);
nor U2092 (N_2092,In_691,In_315);
nand U2093 (N_2093,In_739,In_399);
and U2094 (N_2094,In_382,In_308);
xnor U2095 (N_2095,In_584,In_421);
and U2096 (N_2096,In_459,In_783);
or U2097 (N_2097,In_96,In_557);
xor U2098 (N_2098,In_449,In_741);
nand U2099 (N_2099,In_439,In_56);
xor U2100 (N_2100,In_224,In_796);
xor U2101 (N_2101,In_903,In_751);
xnor U2102 (N_2102,In_838,In_41);
xor U2103 (N_2103,In_318,In_434);
and U2104 (N_2104,In_362,In_71);
nor U2105 (N_2105,In_575,In_498);
and U2106 (N_2106,In_730,In_407);
nor U2107 (N_2107,In_828,In_3);
xor U2108 (N_2108,In_709,In_289);
xor U2109 (N_2109,In_634,In_870);
nor U2110 (N_2110,In_955,In_19);
nand U2111 (N_2111,In_71,In_789);
nand U2112 (N_2112,In_736,In_567);
and U2113 (N_2113,In_181,In_91);
nand U2114 (N_2114,In_699,In_968);
nand U2115 (N_2115,In_277,In_648);
nor U2116 (N_2116,In_203,In_681);
nor U2117 (N_2117,In_90,In_197);
or U2118 (N_2118,In_285,In_318);
nand U2119 (N_2119,In_903,In_647);
nor U2120 (N_2120,In_396,In_321);
nor U2121 (N_2121,In_750,In_521);
nor U2122 (N_2122,In_28,In_273);
and U2123 (N_2123,In_648,In_503);
nand U2124 (N_2124,In_600,In_13);
and U2125 (N_2125,In_455,In_782);
nand U2126 (N_2126,In_332,In_645);
nand U2127 (N_2127,In_634,In_756);
and U2128 (N_2128,In_547,In_295);
xnor U2129 (N_2129,In_424,In_903);
nand U2130 (N_2130,In_197,In_14);
nand U2131 (N_2131,In_385,In_989);
nor U2132 (N_2132,In_953,In_243);
and U2133 (N_2133,In_723,In_145);
xnor U2134 (N_2134,In_226,In_435);
nor U2135 (N_2135,In_442,In_276);
or U2136 (N_2136,In_665,In_69);
nor U2137 (N_2137,In_717,In_709);
or U2138 (N_2138,In_977,In_539);
nand U2139 (N_2139,In_664,In_12);
or U2140 (N_2140,In_41,In_994);
or U2141 (N_2141,In_807,In_847);
nand U2142 (N_2142,In_735,In_632);
or U2143 (N_2143,In_470,In_365);
nand U2144 (N_2144,In_600,In_64);
nor U2145 (N_2145,In_167,In_625);
nand U2146 (N_2146,In_725,In_465);
and U2147 (N_2147,In_327,In_496);
or U2148 (N_2148,In_425,In_762);
nand U2149 (N_2149,In_601,In_937);
nand U2150 (N_2150,In_714,In_699);
nand U2151 (N_2151,In_809,In_178);
and U2152 (N_2152,In_647,In_19);
nor U2153 (N_2153,In_119,In_260);
nor U2154 (N_2154,In_195,In_321);
and U2155 (N_2155,In_602,In_252);
xnor U2156 (N_2156,In_824,In_185);
or U2157 (N_2157,In_699,In_356);
and U2158 (N_2158,In_906,In_980);
or U2159 (N_2159,In_562,In_971);
nor U2160 (N_2160,In_537,In_348);
and U2161 (N_2161,In_237,In_481);
and U2162 (N_2162,In_951,In_706);
nand U2163 (N_2163,In_185,In_687);
nor U2164 (N_2164,In_546,In_671);
nor U2165 (N_2165,In_345,In_138);
xor U2166 (N_2166,In_10,In_396);
and U2167 (N_2167,In_649,In_220);
nor U2168 (N_2168,In_872,In_475);
nor U2169 (N_2169,In_412,In_509);
nor U2170 (N_2170,In_613,In_870);
nor U2171 (N_2171,In_392,In_135);
and U2172 (N_2172,In_291,In_182);
and U2173 (N_2173,In_699,In_814);
xnor U2174 (N_2174,In_544,In_347);
nand U2175 (N_2175,In_858,In_758);
xnor U2176 (N_2176,In_229,In_227);
and U2177 (N_2177,In_294,In_794);
nor U2178 (N_2178,In_927,In_437);
and U2179 (N_2179,In_268,In_519);
xor U2180 (N_2180,In_675,In_68);
nand U2181 (N_2181,In_988,In_634);
nand U2182 (N_2182,In_34,In_356);
and U2183 (N_2183,In_290,In_541);
nand U2184 (N_2184,In_963,In_296);
and U2185 (N_2185,In_740,In_354);
or U2186 (N_2186,In_865,In_917);
xnor U2187 (N_2187,In_237,In_312);
xor U2188 (N_2188,In_640,In_896);
or U2189 (N_2189,In_992,In_129);
nand U2190 (N_2190,In_511,In_308);
nand U2191 (N_2191,In_881,In_715);
nand U2192 (N_2192,In_774,In_991);
or U2193 (N_2193,In_97,In_785);
or U2194 (N_2194,In_451,In_291);
nand U2195 (N_2195,In_101,In_713);
or U2196 (N_2196,In_619,In_831);
or U2197 (N_2197,In_438,In_541);
xor U2198 (N_2198,In_782,In_300);
xnor U2199 (N_2199,In_325,In_48);
nor U2200 (N_2200,In_895,In_564);
or U2201 (N_2201,In_649,In_432);
xor U2202 (N_2202,In_468,In_803);
nor U2203 (N_2203,In_239,In_644);
nor U2204 (N_2204,In_506,In_810);
and U2205 (N_2205,In_952,In_753);
nand U2206 (N_2206,In_956,In_482);
xor U2207 (N_2207,In_143,In_560);
or U2208 (N_2208,In_43,In_222);
and U2209 (N_2209,In_357,In_551);
or U2210 (N_2210,In_969,In_295);
or U2211 (N_2211,In_408,In_660);
and U2212 (N_2212,In_347,In_323);
xnor U2213 (N_2213,In_152,In_567);
nor U2214 (N_2214,In_259,In_121);
or U2215 (N_2215,In_283,In_221);
or U2216 (N_2216,In_263,In_964);
nor U2217 (N_2217,In_648,In_530);
or U2218 (N_2218,In_773,In_708);
nand U2219 (N_2219,In_56,In_781);
and U2220 (N_2220,In_17,In_36);
nand U2221 (N_2221,In_465,In_292);
nor U2222 (N_2222,In_859,In_160);
nor U2223 (N_2223,In_125,In_838);
or U2224 (N_2224,In_806,In_227);
nand U2225 (N_2225,In_350,In_693);
or U2226 (N_2226,In_996,In_153);
and U2227 (N_2227,In_643,In_559);
nand U2228 (N_2228,In_734,In_552);
xnor U2229 (N_2229,In_856,In_869);
nor U2230 (N_2230,In_300,In_947);
xnor U2231 (N_2231,In_527,In_880);
or U2232 (N_2232,In_736,In_354);
xnor U2233 (N_2233,In_320,In_903);
nand U2234 (N_2234,In_104,In_332);
nor U2235 (N_2235,In_786,In_119);
nor U2236 (N_2236,In_138,In_741);
nand U2237 (N_2237,In_494,In_874);
xnor U2238 (N_2238,In_57,In_772);
and U2239 (N_2239,In_189,In_7);
xor U2240 (N_2240,In_682,In_681);
or U2241 (N_2241,In_529,In_261);
nor U2242 (N_2242,In_636,In_89);
nor U2243 (N_2243,In_134,In_844);
or U2244 (N_2244,In_548,In_704);
or U2245 (N_2245,In_314,In_969);
or U2246 (N_2246,In_178,In_420);
xor U2247 (N_2247,In_196,In_895);
and U2248 (N_2248,In_836,In_557);
or U2249 (N_2249,In_256,In_893);
xor U2250 (N_2250,In_489,In_997);
and U2251 (N_2251,In_34,In_560);
nand U2252 (N_2252,In_183,In_637);
or U2253 (N_2253,In_35,In_732);
and U2254 (N_2254,In_767,In_381);
nand U2255 (N_2255,In_749,In_453);
xnor U2256 (N_2256,In_916,In_263);
and U2257 (N_2257,In_283,In_66);
nor U2258 (N_2258,In_733,In_908);
xor U2259 (N_2259,In_184,In_400);
nand U2260 (N_2260,In_740,In_231);
or U2261 (N_2261,In_957,In_172);
or U2262 (N_2262,In_418,In_570);
xnor U2263 (N_2263,In_952,In_904);
nand U2264 (N_2264,In_777,In_395);
or U2265 (N_2265,In_36,In_233);
nor U2266 (N_2266,In_588,In_895);
nor U2267 (N_2267,In_211,In_516);
xor U2268 (N_2268,In_761,In_328);
xor U2269 (N_2269,In_215,In_892);
nand U2270 (N_2270,In_442,In_593);
nor U2271 (N_2271,In_333,In_812);
xnor U2272 (N_2272,In_51,In_768);
or U2273 (N_2273,In_401,In_900);
nor U2274 (N_2274,In_270,In_967);
nor U2275 (N_2275,In_298,In_7);
nand U2276 (N_2276,In_805,In_978);
xor U2277 (N_2277,In_833,In_143);
nand U2278 (N_2278,In_483,In_755);
xnor U2279 (N_2279,In_258,In_401);
and U2280 (N_2280,In_902,In_636);
and U2281 (N_2281,In_753,In_862);
and U2282 (N_2282,In_257,In_581);
nor U2283 (N_2283,In_969,In_764);
xor U2284 (N_2284,In_221,In_486);
xor U2285 (N_2285,In_826,In_692);
xnor U2286 (N_2286,In_618,In_945);
and U2287 (N_2287,In_545,In_532);
and U2288 (N_2288,In_600,In_488);
or U2289 (N_2289,In_399,In_206);
or U2290 (N_2290,In_413,In_725);
and U2291 (N_2291,In_260,In_562);
nor U2292 (N_2292,In_680,In_978);
xor U2293 (N_2293,In_859,In_13);
nor U2294 (N_2294,In_788,In_593);
nor U2295 (N_2295,In_761,In_305);
xor U2296 (N_2296,In_331,In_285);
or U2297 (N_2297,In_707,In_610);
and U2298 (N_2298,In_881,In_272);
nand U2299 (N_2299,In_757,In_390);
or U2300 (N_2300,In_985,In_665);
nand U2301 (N_2301,In_662,In_275);
nor U2302 (N_2302,In_311,In_242);
and U2303 (N_2303,In_719,In_153);
nand U2304 (N_2304,In_909,In_947);
and U2305 (N_2305,In_53,In_981);
nor U2306 (N_2306,In_213,In_782);
or U2307 (N_2307,In_293,In_937);
xnor U2308 (N_2308,In_960,In_838);
nand U2309 (N_2309,In_638,In_745);
and U2310 (N_2310,In_79,In_533);
xnor U2311 (N_2311,In_220,In_294);
nor U2312 (N_2312,In_288,In_251);
nor U2313 (N_2313,In_526,In_99);
and U2314 (N_2314,In_383,In_892);
and U2315 (N_2315,In_648,In_249);
nor U2316 (N_2316,In_63,In_768);
xnor U2317 (N_2317,In_105,In_364);
and U2318 (N_2318,In_325,In_981);
xor U2319 (N_2319,In_257,In_223);
nor U2320 (N_2320,In_658,In_437);
or U2321 (N_2321,In_536,In_861);
xor U2322 (N_2322,In_172,In_571);
or U2323 (N_2323,In_906,In_451);
nor U2324 (N_2324,In_610,In_158);
xor U2325 (N_2325,In_134,In_343);
xnor U2326 (N_2326,In_47,In_976);
and U2327 (N_2327,In_255,In_431);
nand U2328 (N_2328,In_406,In_929);
nor U2329 (N_2329,In_240,In_611);
or U2330 (N_2330,In_369,In_921);
nand U2331 (N_2331,In_265,In_753);
xnor U2332 (N_2332,In_200,In_339);
and U2333 (N_2333,In_974,In_308);
nand U2334 (N_2334,In_374,In_493);
or U2335 (N_2335,In_515,In_498);
xor U2336 (N_2336,In_740,In_992);
nor U2337 (N_2337,In_748,In_658);
xor U2338 (N_2338,In_608,In_136);
nor U2339 (N_2339,In_902,In_957);
xnor U2340 (N_2340,In_752,In_337);
or U2341 (N_2341,In_693,In_311);
nor U2342 (N_2342,In_858,In_995);
nand U2343 (N_2343,In_333,In_5);
xnor U2344 (N_2344,In_27,In_337);
nand U2345 (N_2345,In_996,In_921);
nand U2346 (N_2346,In_471,In_908);
nor U2347 (N_2347,In_175,In_825);
nand U2348 (N_2348,In_583,In_862);
nand U2349 (N_2349,In_292,In_197);
nor U2350 (N_2350,In_476,In_665);
xnor U2351 (N_2351,In_217,In_126);
xnor U2352 (N_2352,In_829,In_866);
nand U2353 (N_2353,In_603,In_722);
nand U2354 (N_2354,In_744,In_963);
xor U2355 (N_2355,In_79,In_467);
and U2356 (N_2356,In_523,In_654);
and U2357 (N_2357,In_353,In_554);
nor U2358 (N_2358,In_818,In_907);
nor U2359 (N_2359,In_812,In_264);
nand U2360 (N_2360,In_982,In_99);
xor U2361 (N_2361,In_884,In_449);
xor U2362 (N_2362,In_493,In_962);
or U2363 (N_2363,In_312,In_191);
or U2364 (N_2364,In_772,In_320);
and U2365 (N_2365,In_231,In_516);
and U2366 (N_2366,In_407,In_154);
nor U2367 (N_2367,In_21,In_658);
nor U2368 (N_2368,In_135,In_756);
or U2369 (N_2369,In_297,In_710);
nand U2370 (N_2370,In_932,In_636);
nand U2371 (N_2371,In_309,In_324);
and U2372 (N_2372,In_601,In_198);
nand U2373 (N_2373,In_683,In_803);
or U2374 (N_2374,In_505,In_168);
nand U2375 (N_2375,In_440,In_710);
and U2376 (N_2376,In_56,In_569);
or U2377 (N_2377,In_635,In_666);
and U2378 (N_2378,In_911,In_899);
nor U2379 (N_2379,In_758,In_97);
and U2380 (N_2380,In_446,In_488);
and U2381 (N_2381,In_231,In_405);
nor U2382 (N_2382,In_478,In_846);
or U2383 (N_2383,In_363,In_612);
or U2384 (N_2384,In_592,In_852);
nor U2385 (N_2385,In_18,In_666);
and U2386 (N_2386,In_724,In_835);
and U2387 (N_2387,In_362,In_74);
xor U2388 (N_2388,In_724,In_709);
xnor U2389 (N_2389,In_619,In_345);
nand U2390 (N_2390,In_82,In_26);
nand U2391 (N_2391,In_80,In_682);
nand U2392 (N_2392,In_156,In_842);
or U2393 (N_2393,In_221,In_718);
or U2394 (N_2394,In_469,In_158);
nor U2395 (N_2395,In_948,In_289);
nand U2396 (N_2396,In_577,In_488);
and U2397 (N_2397,In_965,In_739);
or U2398 (N_2398,In_544,In_483);
and U2399 (N_2399,In_645,In_721);
or U2400 (N_2400,In_807,In_302);
and U2401 (N_2401,In_827,In_252);
and U2402 (N_2402,In_80,In_225);
or U2403 (N_2403,In_925,In_597);
nor U2404 (N_2404,In_249,In_33);
nand U2405 (N_2405,In_118,In_710);
or U2406 (N_2406,In_889,In_612);
nor U2407 (N_2407,In_688,In_415);
or U2408 (N_2408,In_689,In_902);
xor U2409 (N_2409,In_321,In_20);
or U2410 (N_2410,In_576,In_574);
nor U2411 (N_2411,In_527,In_90);
and U2412 (N_2412,In_995,In_553);
nor U2413 (N_2413,In_551,In_470);
or U2414 (N_2414,In_702,In_369);
or U2415 (N_2415,In_1,In_588);
xnor U2416 (N_2416,In_344,In_144);
or U2417 (N_2417,In_414,In_727);
and U2418 (N_2418,In_878,In_876);
nor U2419 (N_2419,In_527,In_909);
nand U2420 (N_2420,In_326,In_996);
nand U2421 (N_2421,In_344,In_318);
xnor U2422 (N_2422,In_408,In_822);
xor U2423 (N_2423,In_351,In_504);
or U2424 (N_2424,In_271,In_517);
nand U2425 (N_2425,In_971,In_103);
and U2426 (N_2426,In_368,In_962);
and U2427 (N_2427,In_22,In_622);
and U2428 (N_2428,In_456,In_845);
nand U2429 (N_2429,In_131,In_57);
nor U2430 (N_2430,In_714,In_862);
or U2431 (N_2431,In_29,In_315);
xor U2432 (N_2432,In_930,In_474);
and U2433 (N_2433,In_899,In_130);
xor U2434 (N_2434,In_494,In_210);
nand U2435 (N_2435,In_965,In_681);
nand U2436 (N_2436,In_772,In_795);
nand U2437 (N_2437,In_281,In_694);
and U2438 (N_2438,In_999,In_395);
nor U2439 (N_2439,In_831,In_895);
xnor U2440 (N_2440,In_16,In_962);
nand U2441 (N_2441,In_205,In_372);
and U2442 (N_2442,In_166,In_83);
or U2443 (N_2443,In_842,In_256);
xnor U2444 (N_2444,In_835,In_172);
nor U2445 (N_2445,In_178,In_814);
nand U2446 (N_2446,In_122,In_187);
and U2447 (N_2447,In_603,In_982);
nand U2448 (N_2448,In_957,In_55);
nor U2449 (N_2449,In_384,In_557);
or U2450 (N_2450,In_100,In_243);
or U2451 (N_2451,In_718,In_12);
or U2452 (N_2452,In_891,In_722);
or U2453 (N_2453,In_42,In_680);
xor U2454 (N_2454,In_388,In_392);
nand U2455 (N_2455,In_254,In_228);
or U2456 (N_2456,In_157,In_368);
and U2457 (N_2457,In_937,In_345);
nor U2458 (N_2458,In_995,In_269);
xor U2459 (N_2459,In_162,In_63);
and U2460 (N_2460,In_103,In_760);
xor U2461 (N_2461,In_407,In_618);
nor U2462 (N_2462,In_696,In_991);
nor U2463 (N_2463,In_255,In_203);
nor U2464 (N_2464,In_496,In_48);
nand U2465 (N_2465,In_110,In_690);
nand U2466 (N_2466,In_982,In_512);
nand U2467 (N_2467,In_84,In_250);
nand U2468 (N_2468,In_666,In_805);
and U2469 (N_2469,In_710,In_331);
nand U2470 (N_2470,In_61,In_509);
nand U2471 (N_2471,In_248,In_452);
nand U2472 (N_2472,In_313,In_862);
nor U2473 (N_2473,In_904,In_911);
nor U2474 (N_2474,In_609,In_62);
or U2475 (N_2475,In_718,In_958);
or U2476 (N_2476,In_872,In_805);
nand U2477 (N_2477,In_599,In_673);
or U2478 (N_2478,In_278,In_901);
nand U2479 (N_2479,In_531,In_450);
nand U2480 (N_2480,In_701,In_749);
nand U2481 (N_2481,In_590,In_367);
nand U2482 (N_2482,In_730,In_875);
and U2483 (N_2483,In_58,In_751);
and U2484 (N_2484,In_293,In_55);
xnor U2485 (N_2485,In_17,In_626);
or U2486 (N_2486,In_52,In_310);
and U2487 (N_2487,In_97,In_370);
and U2488 (N_2488,In_568,In_486);
nand U2489 (N_2489,In_980,In_593);
or U2490 (N_2490,In_584,In_13);
and U2491 (N_2491,In_669,In_410);
xnor U2492 (N_2492,In_156,In_691);
xnor U2493 (N_2493,In_34,In_659);
nor U2494 (N_2494,In_650,In_681);
or U2495 (N_2495,In_629,In_283);
nor U2496 (N_2496,In_330,In_635);
nor U2497 (N_2497,In_114,In_668);
or U2498 (N_2498,In_279,In_375);
and U2499 (N_2499,In_665,In_593);
or U2500 (N_2500,In_216,In_498);
and U2501 (N_2501,In_67,In_378);
and U2502 (N_2502,In_155,In_700);
xnor U2503 (N_2503,In_837,In_154);
nor U2504 (N_2504,In_237,In_59);
or U2505 (N_2505,In_639,In_602);
nand U2506 (N_2506,In_438,In_197);
nor U2507 (N_2507,In_235,In_813);
and U2508 (N_2508,In_29,In_428);
xor U2509 (N_2509,In_738,In_700);
nor U2510 (N_2510,In_715,In_577);
and U2511 (N_2511,In_261,In_847);
or U2512 (N_2512,In_404,In_194);
or U2513 (N_2513,In_765,In_460);
nor U2514 (N_2514,In_63,In_585);
or U2515 (N_2515,In_884,In_516);
nor U2516 (N_2516,In_937,In_691);
or U2517 (N_2517,In_946,In_50);
nor U2518 (N_2518,In_312,In_243);
or U2519 (N_2519,In_189,In_911);
nor U2520 (N_2520,In_538,In_379);
or U2521 (N_2521,In_386,In_993);
nor U2522 (N_2522,In_88,In_593);
xor U2523 (N_2523,In_620,In_118);
xor U2524 (N_2524,In_866,In_235);
or U2525 (N_2525,In_563,In_397);
nand U2526 (N_2526,In_399,In_608);
xnor U2527 (N_2527,In_746,In_426);
xnor U2528 (N_2528,In_793,In_658);
or U2529 (N_2529,In_733,In_871);
nand U2530 (N_2530,In_976,In_486);
nor U2531 (N_2531,In_166,In_947);
nand U2532 (N_2532,In_673,In_675);
or U2533 (N_2533,In_191,In_521);
xor U2534 (N_2534,In_188,In_314);
and U2535 (N_2535,In_604,In_885);
nor U2536 (N_2536,In_650,In_453);
and U2537 (N_2537,In_890,In_632);
xnor U2538 (N_2538,In_163,In_967);
nor U2539 (N_2539,In_305,In_413);
or U2540 (N_2540,In_463,In_828);
nand U2541 (N_2541,In_955,In_118);
xor U2542 (N_2542,In_991,In_898);
and U2543 (N_2543,In_268,In_380);
nor U2544 (N_2544,In_341,In_614);
or U2545 (N_2545,In_163,In_247);
nor U2546 (N_2546,In_618,In_971);
and U2547 (N_2547,In_413,In_544);
xnor U2548 (N_2548,In_736,In_103);
xor U2549 (N_2549,In_250,In_139);
nor U2550 (N_2550,In_231,In_364);
nor U2551 (N_2551,In_714,In_837);
nand U2552 (N_2552,In_68,In_19);
xnor U2553 (N_2553,In_705,In_676);
nand U2554 (N_2554,In_508,In_773);
or U2555 (N_2555,In_554,In_597);
and U2556 (N_2556,In_782,In_429);
xor U2557 (N_2557,In_92,In_623);
nor U2558 (N_2558,In_292,In_573);
nand U2559 (N_2559,In_533,In_680);
and U2560 (N_2560,In_907,In_873);
or U2561 (N_2561,In_652,In_887);
nand U2562 (N_2562,In_192,In_481);
nor U2563 (N_2563,In_50,In_761);
xor U2564 (N_2564,In_860,In_686);
xnor U2565 (N_2565,In_679,In_603);
xnor U2566 (N_2566,In_777,In_350);
nor U2567 (N_2567,In_998,In_554);
nor U2568 (N_2568,In_559,In_564);
and U2569 (N_2569,In_234,In_180);
or U2570 (N_2570,In_754,In_208);
and U2571 (N_2571,In_945,In_706);
and U2572 (N_2572,In_953,In_453);
and U2573 (N_2573,In_477,In_628);
or U2574 (N_2574,In_218,In_370);
nor U2575 (N_2575,In_217,In_686);
and U2576 (N_2576,In_136,In_105);
nand U2577 (N_2577,In_702,In_996);
xnor U2578 (N_2578,In_882,In_173);
nor U2579 (N_2579,In_70,In_521);
xnor U2580 (N_2580,In_371,In_852);
nand U2581 (N_2581,In_898,In_446);
or U2582 (N_2582,In_324,In_788);
nor U2583 (N_2583,In_503,In_789);
nand U2584 (N_2584,In_487,In_139);
or U2585 (N_2585,In_840,In_588);
and U2586 (N_2586,In_721,In_548);
or U2587 (N_2587,In_165,In_122);
or U2588 (N_2588,In_743,In_279);
xor U2589 (N_2589,In_483,In_961);
xnor U2590 (N_2590,In_834,In_565);
nor U2591 (N_2591,In_998,In_261);
nand U2592 (N_2592,In_621,In_282);
or U2593 (N_2593,In_140,In_615);
and U2594 (N_2594,In_221,In_751);
and U2595 (N_2595,In_553,In_266);
and U2596 (N_2596,In_371,In_183);
or U2597 (N_2597,In_369,In_980);
nor U2598 (N_2598,In_587,In_849);
and U2599 (N_2599,In_119,In_371);
nor U2600 (N_2600,In_551,In_736);
nor U2601 (N_2601,In_517,In_937);
nor U2602 (N_2602,In_724,In_368);
nor U2603 (N_2603,In_135,In_723);
or U2604 (N_2604,In_94,In_753);
nor U2605 (N_2605,In_330,In_562);
or U2606 (N_2606,In_889,In_900);
xor U2607 (N_2607,In_758,In_919);
nor U2608 (N_2608,In_662,In_919);
or U2609 (N_2609,In_154,In_75);
nand U2610 (N_2610,In_860,In_785);
nor U2611 (N_2611,In_451,In_350);
and U2612 (N_2612,In_211,In_505);
xnor U2613 (N_2613,In_754,In_55);
nand U2614 (N_2614,In_403,In_375);
and U2615 (N_2615,In_299,In_331);
nand U2616 (N_2616,In_133,In_528);
or U2617 (N_2617,In_946,In_82);
xnor U2618 (N_2618,In_314,In_808);
nand U2619 (N_2619,In_53,In_806);
nand U2620 (N_2620,In_458,In_205);
xnor U2621 (N_2621,In_243,In_816);
xor U2622 (N_2622,In_14,In_167);
or U2623 (N_2623,In_70,In_43);
nand U2624 (N_2624,In_598,In_286);
or U2625 (N_2625,In_806,In_407);
and U2626 (N_2626,In_764,In_205);
and U2627 (N_2627,In_584,In_61);
nor U2628 (N_2628,In_489,In_341);
xor U2629 (N_2629,In_766,In_699);
or U2630 (N_2630,In_291,In_328);
nor U2631 (N_2631,In_376,In_689);
and U2632 (N_2632,In_182,In_655);
nor U2633 (N_2633,In_936,In_97);
nor U2634 (N_2634,In_225,In_812);
or U2635 (N_2635,In_284,In_330);
xnor U2636 (N_2636,In_763,In_919);
xor U2637 (N_2637,In_252,In_720);
xnor U2638 (N_2638,In_26,In_45);
xnor U2639 (N_2639,In_562,In_736);
nor U2640 (N_2640,In_41,In_629);
nand U2641 (N_2641,In_128,In_455);
and U2642 (N_2642,In_131,In_757);
or U2643 (N_2643,In_266,In_681);
xnor U2644 (N_2644,In_295,In_231);
or U2645 (N_2645,In_431,In_241);
or U2646 (N_2646,In_25,In_407);
or U2647 (N_2647,In_868,In_983);
nor U2648 (N_2648,In_499,In_95);
xor U2649 (N_2649,In_205,In_924);
xor U2650 (N_2650,In_920,In_335);
nand U2651 (N_2651,In_750,In_821);
and U2652 (N_2652,In_606,In_434);
xnor U2653 (N_2653,In_16,In_532);
and U2654 (N_2654,In_507,In_128);
nand U2655 (N_2655,In_401,In_277);
nor U2656 (N_2656,In_586,In_313);
xnor U2657 (N_2657,In_813,In_645);
xnor U2658 (N_2658,In_538,In_74);
xnor U2659 (N_2659,In_453,In_830);
or U2660 (N_2660,In_705,In_683);
xnor U2661 (N_2661,In_535,In_632);
and U2662 (N_2662,In_695,In_744);
xnor U2663 (N_2663,In_706,In_808);
and U2664 (N_2664,In_357,In_869);
nor U2665 (N_2665,In_114,In_621);
or U2666 (N_2666,In_503,In_108);
nand U2667 (N_2667,In_976,In_992);
and U2668 (N_2668,In_739,In_743);
and U2669 (N_2669,In_715,In_857);
nor U2670 (N_2670,In_550,In_972);
or U2671 (N_2671,In_822,In_69);
xnor U2672 (N_2672,In_721,In_207);
or U2673 (N_2673,In_99,In_123);
and U2674 (N_2674,In_616,In_940);
or U2675 (N_2675,In_82,In_273);
nand U2676 (N_2676,In_24,In_927);
and U2677 (N_2677,In_693,In_155);
nor U2678 (N_2678,In_495,In_302);
and U2679 (N_2679,In_209,In_850);
nor U2680 (N_2680,In_600,In_755);
nand U2681 (N_2681,In_178,In_466);
and U2682 (N_2682,In_427,In_729);
or U2683 (N_2683,In_972,In_167);
or U2684 (N_2684,In_374,In_45);
nor U2685 (N_2685,In_786,In_509);
nand U2686 (N_2686,In_119,In_243);
nor U2687 (N_2687,In_845,In_332);
or U2688 (N_2688,In_175,In_78);
nor U2689 (N_2689,In_192,In_592);
or U2690 (N_2690,In_1,In_234);
nor U2691 (N_2691,In_187,In_510);
nor U2692 (N_2692,In_19,In_355);
xnor U2693 (N_2693,In_291,In_82);
nor U2694 (N_2694,In_243,In_14);
and U2695 (N_2695,In_97,In_452);
nand U2696 (N_2696,In_817,In_864);
nor U2697 (N_2697,In_539,In_831);
or U2698 (N_2698,In_874,In_132);
nand U2699 (N_2699,In_194,In_633);
nor U2700 (N_2700,In_694,In_889);
xor U2701 (N_2701,In_938,In_171);
nor U2702 (N_2702,In_142,In_566);
and U2703 (N_2703,In_331,In_553);
nand U2704 (N_2704,In_316,In_425);
or U2705 (N_2705,In_455,In_461);
nand U2706 (N_2706,In_322,In_243);
nor U2707 (N_2707,In_666,In_718);
and U2708 (N_2708,In_890,In_712);
xnor U2709 (N_2709,In_139,In_526);
nand U2710 (N_2710,In_260,In_354);
and U2711 (N_2711,In_530,In_206);
xnor U2712 (N_2712,In_279,In_468);
and U2713 (N_2713,In_867,In_744);
and U2714 (N_2714,In_532,In_881);
nor U2715 (N_2715,In_880,In_306);
xnor U2716 (N_2716,In_696,In_546);
xor U2717 (N_2717,In_72,In_579);
xnor U2718 (N_2718,In_914,In_897);
or U2719 (N_2719,In_447,In_451);
nand U2720 (N_2720,In_419,In_204);
nand U2721 (N_2721,In_443,In_185);
nor U2722 (N_2722,In_454,In_994);
nand U2723 (N_2723,In_424,In_588);
xnor U2724 (N_2724,In_969,In_361);
and U2725 (N_2725,In_484,In_729);
and U2726 (N_2726,In_831,In_736);
xor U2727 (N_2727,In_158,In_730);
and U2728 (N_2728,In_900,In_61);
and U2729 (N_2729,In_34,In_332);
nand U2730 (N_2730,In_320,In_689);
nor U2731 (N_2731,In_763,In_246);
xnor U2732 (N_2732,In_252,In_559);
nand U2733 (N_2733,In_576,In_246);
or U2734 (N_2734,In_325,In_933);
or U2735 (N_2735,In_546,In_466);
or U2736 (N_2736,In_730,In_376);
and U2737 (N_2737,In_195,In_337);
and U2738 (N_2738,In_313,In_231);
and U2739 (N_2739,In_56,In_263);
and U2740 (N_2740,In_472,In_982);
nand U2741 (N_2741,In_32,In_492);
nor U2742 (N_2742,In_731,In_809);
nand U2743 (N_2743,In_537,In_5);
nand U2744 (N_2744,In_58,In_213);
nor U2745 (N_2745,In_583,In_296);
and U2746 (N_2746,In_910,In_820);
and U2747 (N_2747,In_325,In_301);
nor U2748 (N_2748,In_48,In_386);
or U2749 (N_2749,In_436,In_864);
or U2750 (N_2750,In_961,In_926);
nor U2751 (N_2751,In_877,In_661);
xnor U2752 (N_2752,In_572,In_46);
xnor U2753 (N_2753,In_686,In_269);
or U2754 (N_2754,In_917,In_113);
nor U2755 (N_2755,In_135,In_518);
nand U2756 (N_2756,In_340,In_135);
and U2757 (N_2757,In_797,In_938);
or U2758 (N_2758,In_250,In_647);
or U2759 (N_2759,In_943,In_563);
and U2760 (N_2760,In_729,In_587);
and U2761 (N_2761,In_664,In_919);
nand U2762 (N_2762,In_680,In_905);
and U2763 (N_2763,In_553,In_435);
nand U2764 (N_2764,In_109,In_385);
nand U2765 (N_2765,In_850,In_84);
or U2766 (N_2766,In_518,In_506);
or U2767 (N_2767,In_251,In_391);
nand U2768 (N_2768,In_940,In_841);
xor U2769 (N_2769,In_877,In_803);
and U2770 (N_2770,In_645,In_466);
xor U2771 (N_2771,In_104,In_463);
nand U2772 (N_2772,In_134,In_175);
nor U2773 (N_2773,In_289,In_178);
and U2774 (N_2774,In_506,In_653);
xnor U2775 (N_2775,In_301,In_493);
and U2776 (N_2776,In_805,In_66);
xor U2777 (N_2777,In_338,In_891);
or U2778 (N_2778,In_249,In_8);
and U2779 (N_2779,In_538,In_641);
or U2780 (N_2780,In_649,In_247);
nor U2781 (N_2781,In_55,In_103);
nand U2782 (N_2782,In_383,In_586);
and U2783 (N_2783,In_858,In_651);
nor U2784 (N_2784,In_540,In_280);
xor U2785 (N_2785,In_955,In_264);
or U2786 (N_2786,In_271,In_840);
xnor U2787 (N_2787,In_594,In_336);
nand U2788 (N_2788,In_164,In_611);
xor U2789 (N_2789,In_568,In_411);
and U2790 (N_2790,In_230,In_240);
nor U2791 (N_2791,In_224,In_364);
or U2792 (N_2792,In_857,In_123);
nand U2793 (N_2793,In_771,In_540);
xnor U2794 (N_2794,In_374,In_436);
nand U2795 (N_2795,In_353,In_875);
or U2796 (N_2796,In_530,In_832);
xnor U2797 (N_2797,In_953,In_404);
and U2798 (N_2798,In_158,In_668);
and U2799 (N_2799,In_908,In_989);
and U2800 (N_2800,In_358,In_383);
nor U2801 (N_2801,In_985,In_307);
nand U2802 (N_2802,In_956,In_879);
or U2803 (N_2803,In_328,In_938);
or U2804 (N_2804,In_666,In_227);
xor U2805 (N_2805,In_290,In_796);
or U2806 (N_2806,In_470,In_182);
nor U2807 (N_2807,In_788,In_175);
and U2808 (N_2808,In_191,In_824);
nand U2809 (N_2809,In_606,In_3);
nor U2810 (N_2810,In_158,In_744);
nand U2811 (N_2811,In_438,In_979);
xnor U2812 (N_2812,In_786,In_944);
and U2813 (N_2813,In_627,In_953);
nand U2814 (N_2814,In_164,In_867);
nor U2815 (N_2815,In_452,In_523);
and U2816 (N_2816,In_173,In_895);
nand U2817 (N_2817,In_760,In_448);
and U2818 (N_2818,In_139,In_123);
xor U2819 (N_2819,In_947,In_599);
and U2820 (N_2820,In_254,In_168);
xnor U2821 (N_2821,In_997,In_649);
nor U2822 (N_2822,In_185,In_662);
nor U2823 (N_2823,In_221,In_225);
and U2824 (N_2824,In_31,In_968);
or U2825 (N_2825,In_59,In_959);
or U2826 (N_2826,In_270,In_469);
nand U2827 (N_2827,In_529,In_508);
or U2828 (N_2828,In_643,In_427);
nor U2829 (N_2829,In_788,In_607);
nand U2830 (N_2830,In_509,In_378);
and U2831 (N_2831,In_15,In_895);
and U2832 (N_2832,In_763,In_532);
or U2833 (N_2833,In_585,In_739);
xnor U2834 (N_2834,In_323,In_126);
and U2835 (N_2835,In_755,In_579);
nor U2836 (N_2836,In_936,In_674);
nor U2837 (N_2837,In_335,In_485);
nor U2838 (N_2838,In_959,In_585);
or U2839 (N_2839,In_877,In_946);
or U2840 (N_2840,In_242,In_40);
xor U2841 (N_2841,In_176,In_164);
or U2842 (N_2842,In_785,In_909);
and U2843 (N_2843,In_474,In_789);
xor U2844 (N_2844,In_387,In_50);
nor U2845 (N_2845,In_568,In_450);
nor U2846 (N_2846,In_551,In_393);
and U2847 (N_2847,In_901,In_293);
or U2848 (N_2848,In_70,In_448);
xor U2849 (N_2849,In_421,In_770);
or U2850 (N_2850,In_288,In_449);
nor U2851 (N_2851,In_905,In_438);
nand U2852 (N_2852,In_835,In_555);
nand U2853 (N_2853,In_17,In_162);
nor U2854 (N_2854,In_915,In_935);
and U2855 (N_2855,In_394,In_122);
and U2856 (N_2856,In_999,In_464);
nand U2857 (N_2857,In_508,In_63);
nor U2858 (N_2858,In_147,In_212);
nor U2859 (N_2859,In_945,In_413);
nor U2860 (N_2860,In_549,In_741);
nor U2861 (N_2861,In_570,In_89);
or U2862 (N_2862,In_755,In_200);
or U2863 (N_2863,In_307,In_808);
xnor U2864 (N_2864,In_878,In_850);
nand U2865 (N_2865,In_801,In_90);
nand U2866 (N_2866,In_468,In_3);
or U2867 (N_2867,In_741,In_361);
nand U2868 (N_2868,In_494,In_490);
nor U2869 (N_2869,In_4,In_512);
and U2870 (N_2870,In_718,In_862);
and U2871 (N_2871,In_291,In_516);
xnor U2872 (N_2872,In_692,In_745);
and U2873 (N_2873,In_933,In_513);
xor U2874 (N_2874,In_746,In_10);
xor U2875 (N_2875,In_626,In_462);
or U2876 (N_2876,In_124,In_434);
and U2877 (N_2877,In_140,In_884);
nor U2878 (N_2878,In_49,In_704);
xor U2879 (N_2879,In_383,In_815);
or U2880 (N_2880,In_617,In_440);
nor U2881 (N_2881,In_325,In_502);
xor U2882 (N_2882,In_651,In_26);
xnor U2883 (N_2883,In_648,In_872);
and U2884 (N_2884,In_539,In_435);
or U2885 (N_2885,In_942,In_585);
xor U2886 (N_2886,In_662,In_199);
nand U2887 (N_2887,In_916,In_387);
or U2888 (N_2888,In_592,In_445);
xnor U2889 (N_2889,In_199,In_565);
xor U2890 (N_2890,In_659,In_646);
and U2891 (N_2891,In_276,In_638);
or U2892 (N_2892,In_574,In_611);
nor U2893 (N_2893,In_270,In_506);
nand U2894 (N_2894,In_309,In_750);
nor U2895 (N_2895,In_379,In_81);
or U2896 (N_2896,In_337,In_287);
xnor U2897 (N_2897,In_111,In_152);
or U2898 (N_2898,In_255,In_720);
nand U2899 (N_2899,In_116,In_516);
xnor U2900 (N_2900,In_557,In_881);
nand U2901 (N_2901,In_150,In_186);
xor U2902 (N_2902,In_683,In_996);
nor U2903 (N_2903,In_552,In_612);
nand U2904 (N_2904,In_981,In_274);
and U2905 (N_2905,In_444,In_851);
and U2906 (N_2906,In_391,In_264);
nand U2907 (N_2907,In_194,In_265);
nand U2908 (N_2908,In_568,In_210);
xnor U2909 (N_2909,In_11,In_201);
or U2910 (N_2910,In_394,In_370);
nor U2911 (N_2911,In_17,In_515);
nor U2912 (N_2912,In_310,In_873);
or U2913 (N_2913,In_620,In_9);
and U2914 (N_2914,In_936,In_116);
or U2915 (N_2915,In_833,In_245);
and U2916 (N_2916,In_198,In_501);
nand U2917 (N_2917,In_422,In_68);
nor U2918 (N_2918,In_968,In_482);
or U2919 (N_2919,In_62,In_778);
nand U2920 (N_2920,In_462,In_810);
or U2921 (N_2921,In_524,In_225);
or U2922 (N_2922,In_870,In_891);
and U2923 (N_2923,In_194,In_543);
or U2924 (N_2924,In_698,In_833);
xor U2925 (N_2925,In_806,In_554);
and U2926 (N_2926,In_386,In_230);
and U2927 (N_2927,In_290,In_513);
nor U2928 (N_2928,In_757,In_661);
nor U2929 (N_2929,In_691,In_538);
nand U2930 (N_2930,In_963,In_176);
or U2931 (N_2931,In_723,In_777);
xnor U2932 (N_2932,In_29,In_79);
and U2933 (N_2933,In_73,In_694);
and U2934 (N_2934,In_687,In_245);
nor U2935 (N_2935,In_859,In_947);
or U2936 (N_2936,In_569,In_626);
nor U2937 (N_2937,In_594,In_487);
nand U2938 (N_2938,In_411,In_34);
nand U2939 (N_2939,In_884,In_674);
nand U2940 (N_2940,In_492,In_217);
nand U2941 (N_2941,In_995,In_618);
nor U2942 (N_2942,In_141,In_460);
xor U2943 (N_2943,In_786,In_94);
nor U2944 (N_2944,In_606,In_670);
nor U2945 (N_2945,In_408,In_512);
and U2946 (N_2946,In_634,In_235);
nand U2947 (N_2947,In_185,In_155);
xnor U2948 (N_2948,In_395,In_673);
or U2949 (N_2949,In_497,In_631);
xor U2950 (N_2950,In_257,In_999);
xnor U2951 (N_2951,In_652,In_979);
nand U2952 (N_2952,In_330,In_902);
nand U2953 (N_2953,In_711,In_312);
and U2954 (N_2954,In_485,In_136);
xor U2955 (N_2955,In_83,In_695);
xor U2956 (N_2956,In_514,In_617);
and U2957 (N_2957,In_906,In_859);
nand U2958 (N_2958,In_466,In_563);
xor U2959 (N_2959,In_136,In_754);
or U2960 (N_2960,In_153,In_931);
nor U2961 (N_2961,In_518,In_552);
nor U2962 (N_2962,In_189,In_438);
nand U2963 (N_2963,In_489,In_527);
and U2964 (N_2964,In_316,In_276);
nor U2965 (N_2965,In_669,In_460);
or U2966 (N_2966,In_279,In_842);
and U2967 (N_2967,In_595,In_89);
and U2968 (N_2968,In_565,In_305);
nand U2969 (N_2969,In_118,In_301);
nand U2970 (N_2970,In_256,In_244);
nand U2971 (N_2971,In_805,In_443);
nand U2972 (N_2972,In_424,In_649);
nor U2973 (N_2973,In_565,In_537);
nor U2974 (N_2974,In_602,In_879);
and U2975 (N_2975,In_501,In_532);
xnor U2976 (N_2976,In_635,In_31);
xnor U2977 (N_2977,In_516,In_473);
nand U2978 (N_2978,In_506,In_413);
or U2979 (N_2979,In_738,In_375);
nor U2980 (N_2980,In_937,In_582);
or U2981 (N_2981,In_40,In_418);
nand U2982 (N_2982,In_5,In_187);
and U2983 (N_2983,In_304,In_302);
xnor U2984 (N_2984,In_319,In_962);
or U2985 (N_2985,In_240,In_271);
nand U2986 (N_2986,In_66,In_859);
nand U2987 (N_2987,In_435,In_805);
xnor U2988 (N_2988,In_416,In_292);
xor U2989 (N_2989,In_400,In_541);
nand U2990 (N_2990,In_764,In_815);
nand U2991 (N_2991,In_984,In_837);
nand U2992 (N_2992,In_930,In_584);
nand U2993 (N_2993,In_920,In_890);
and U2994 (N_2994,In_949,In_56);
or U2995 (N_2995,In_64,In_299);
or U2996 (N_2996,In_71,In_368);
xnor U2997 (N_2997,In_866,In_153);
or U2998 (N_2998,In_181,In_417);
nand U2999 (N_2999,In_782,In_937);
and U3000 (N_3000,In_150,In_638);
or U3001 (N_3001,In_957,In_849);
nor U3002 (N_3002,In_702,In_626);
and U3003 (N_3003,In_423,In_978);
and U3004 (N_3004,In_703,In_715);
or U3005 (N_3005,In_271,In_686);
nand U3006 (N_3006,In_781,In_994);
nor U3007 (N_3007,In_378,In_737);
and U3008 (N_3008,In_510,In_614);
xor U3009 (N_3009,In_57,In_138);
nor U3010 (N_3010,In_189,In_136);
nand U3011 (N_3011,In_877,In_220);
and U3012 (N_3012,In_462,In_149);
or U3013 (N_3013,In_212,In_380);
nor U3014 (N_3014,In_969,In_898);
xnor U3015 (N_3015,In_287,In_181);
xor U3016 (N_3016,In_215,In_973);
nor U3017 (N_3017,In_290,In_820);
xor U3018 (N_3018,In_8,In_971);
nor U3019 (N_3019,In_797,In_654);
nand U3020 (N_3020,In_390,In_722);
nand U3021 (N_3021,In_252,In_668);
xnor U3022 (N_3022,In_502,In_916);
and U3023 (N_3023,In_740,In_897);
nor U3024 (N_3024,In_781,In_505);
xnor U3025 (N_3025,In_454,In_261);
nor U3026 (N_3026,In_225,In_206);
or U3027 (N_3027,In_363,In_208);
or U3028 (N_3028,In_87,In_683);
nand U3029 (N_3029,In_361,In_125);
nand U3030 (N_3030,In_291,In_61);
xnor U3031 (N_3031,In_561,In_645);
and U3032 (N_3032,In_64,In_81);
or U3033 (N_3033,In_263,In_952);
and U3034 (N_3034,In_483,In_579);
xor U3035 (N_3035,In_319,In_181);
nor U3036 (N_3036,In_646,In_920);
or U3037 (N_3037,In_789,In_584);
xor U3038 (N_3038,In_393,In_518);
nor U3039 (N_3039,In_0,In_965);
nor U3040 (N_3040,In_491,In_347);
nor U3041 (N_3041,In_774,In_630);
xor U3042 (N_3042,In_61,In_646);
nor U3043 (N_3043,In_145,In_734);
and U3044 (N_3044,In_392,In_580);
nand U3045 (N_3045,In_531,In_649);
or U3046 (N_3046,In_591,In_706);
and U3047 (N_3047,In_83,In_167);
or U3048 (N_3048,In_461,In_955);
or U3049 (N_3049,In_528,In_350);
nor U3050 (N_3050,In_378,In_450);
xnor U3051 (N_3051,In_96,In_654);
and U3052 (N_3052,In_737,In_776);
xor U3053 (N_3053,In_351,In_206);
or U3054 (N_3054,In_470,In_390);
or U3055 (N_3055,In_270,In_752);
xnor U3056 (N_3056,In_989,In_765);
nand U3057 (N_3057,In_139,In_97);
or U3058 (N_3058,In_252,In_850);
nor U3059 (N_3059,In_684,In_525);
and U3060 (N_3060,In_505,In_622);
or U3061 (N_3061,In_812,In_637);
nor U3062 (N_3062,In_119,In_84);
and U3063 (N_3063,In_476,In_116);
or U3064 (N_3064,In_980,In_243);
or U3065 (N_3065,In_863,In_64);
nand U3066 (N_3066,In_158,In_587);
xor U3067 (N_3067,In_757,In_438);
xor U3068 (N_3068,In_676,In_101);
nand U3069 (N_3069,In_1,In_600);
and U3070 (N_3070,In_245,In_639);
or U3071 (N_3071,In_596,In_250);
xor U3072 (N_3072,In_687,In_385);
or U3073 (N_3073,In_429,In_903);
or U3074 (N_3074,In_667,In_200);
xnor U3075 (N_3075,In_233,In_570);
or U3076 (N_3076,In_542,In_366);
or U3077 (N_3077,In_446,In_721);
nand U3078 (N_3078,In_978,In_544);
xor U3079 (N_3079,In_789,In_513);
xor U3080 (N_3080,In_313,In_934);
and U3081 (N_3081,In_867,In_661);
xnor U3082 (N_3082,In_192,In_221);
or U3083 (N_3083,In_390,In_567);
or U3084 (N_3084,In_491,In_262);
xor U3085 (N_3085,In_523,In_941);
xor U3086 (N_3086,In_24,In_546);
and U3087 (N_3087,In_22,In_204);
and U3088 (N_3088,In_858,In_647);
and U3089 (N_3089,In_59,In_917);
xor U3090 (N_3090,In_641,In_328);
nor U3091 (N_3091,In_794,In_94);
nor U3092 (N_3092,In_752,In_322);
nand U3093 (N_3093,In_239,In_987);
or U3094 (N_3094,In_439,In_272);
nand U3095 (N_3095,In_30,In_1);
nand U3096 (N_3096,In_472,In_179);
nand U3097 (N_3097,In_250,In_577);
or U3098 (N_3098,In_921,In_314);
xor U3099 (N_3099,In_635,In_42);
nand U3100 (N_3100,In_964,In_739);
nor U3101 (N_3101,In_582,In_51);
nand U3102 (N_3102,In_195,In_733);
and U3103 (N_3103,In_404,In_760);
nand U3104 (N_3104,In_371,In_809);
nand U3105 (N_3105,In_603,In_923);
xor U3106 (N_3106,In_574,In_678);
nand U3107 (N_3107,In_909,In_524);
or U3108 (N_3108,In_973,In_51);
nor U3109 (N_3109,In_657,In_995);
and U3110 (N_3110,In_718,In_275);
nor U3111 (N_3111,In_937,In_677);
and U3112 (N_3112,In_331,In_793);
xnor U3113 (N_3113,In_966,In_664);
nor U3114 (N_3114,In_803,In_961);
nand U3115 (N_3115,In_704,In_159);
and U3116 (N_3116,In_661,In_410);
xor U3117 (N_3117,In_154,In_159);
or U3118 (N_3118,In_303,In_683);
nor U3119 (N_3119,In_434,In_657);
and U3120 (N_3120,In_969,In_272);
nor U3121 (N_3121,In_462,In_575);
and U3122 (N_3122,In_937,In_386);
nand U3123 (N_3123,In_842,In_154);
xor U3124 (N_3124,In_957,In_266);
nor U3125 (N_3125,In_722,In_42);
nor U3126 (N_3126,In_659,In_718);
and U3127 (N_3127,In_182,In_272);
and U3128 (N_3128,In_198,In_826);
xor U3129 (N_3129,In_525,In_223);
nor U3130 (N_3130,In_937,In_149);
nand U3131 (N_3131,In_524,In_696);
and U3132 (N_3132,In_609,In_487);
nand U3133 (N_3133,In_599,In_431);
xnor U3134 (N_3134,In_719,In_212);
nand U3135 (N_3135,In_715,In_104);
xnor U3136 (N_3136,In_390,In_169);
and U3137 (N_3137,In_185,In_480);
xor U3138 (N_3138,In_868,In_801);
and U3139 (N_3139,In_721,In_646);
xnor U3140 (N_3140,In_389,In_185);
or U3141 (N_3141,In_385,In_264);
and U3142 (N_3142,In_12,In_626);
nand U3143 (N_3143,In_684,In_133);
xor U3144 (N_3144,In_25,In_880);
xor U3145 (N_3145,In_52,In_282);
xnor U3146 (N_3146,In_419,In_751);
nor U3147 (N_3147,In_718,In_923);
and U3148 (N_3148,In_532,In_524);
nand U3149 (N_3149,In_358,In_17);
nand U3150 (N_3150,In_109,In_34);
or U3151 (N_3151,In_277,In_760);
xnor U3152 (N_3152,In_803,In_138);
or U3153 (N_3153,In_446,In_90);
xor U3154 (N_3154,In_679,In_307);
or U3155 (N_3155,In_70,In_298);
nand U3156 (N_3156,In_17,In_622);
xnor U3157 (N_3157,In_579,In_346);
and U3158 (N_3158,In_652,In_606);
nand U3159 (N_3159,In_719,In_234);
xnor U3160 (N_3160,In_263,In_287);
nand U3161 (N_3161,In_846,In_228);
nand U3162 (N_3162,In_817,In_538);
xor U3163 (N_3163,In_951,In_158);
nor U3164 (N_3164,In_854,In_344);
xor U3165 (N_3165,In_109,In_655);
or U3166 (N_3166,In_620,In_1);
nand U3167 (N_3167,In_97,In_665);
and U3168 (N_3168,In_534,In_487);
or U3169 (N_3169,In_755,In_787);
xor U3170 (N_3170,In_0,In_801);
and U3171 (N_3171,In_917,In_373);
or U3172 (N_3172,In_145,In_43);
and U3173 (N_3173,In_789,In_480);
nor U3174 (N_3174,In_460,In_758);
nand U3175 (N_3175,In_966,In_791);
xnor U3176 (N_3176,In_187,In_354);
nand U3177 (N_3177,In_533,In_258);
xor U3178 (N_3178,In_208,In_215);
xor U3179 (N_3179,In_454,In_450);
nor U3180 (N_3180,In_768,In_46);
and U3181 (N_3181,In_748,In_589);
nor U3182 (N_3182,In_440,In_392);
or U3183 (N_3183,In_734,In_336);
and U3184 (N_3184,In_583,In_265);
nor U3185 (N_3185,In_56,In_66);
and U3186 (N_3186,In_572,In_724);
and U3187 (N_3187,In_461,In_568);
and U3188 (N_3188,In_317,In_566);
nor U3189 (N_3189,In_983,In_589);
or U3190 (N_3190,In_55,In_101);
or U3191 (N_3191,In_402,In_133);
nand U3192 (N_3192,In_650,In_140);
xor U3193 (N_3193,In_508,In_745);
xor U3194 (N_3194,In_818,In_260);
nand U3195 (N_3195,In_353,In_52);
and U3196 (N_3196,In_866,In_72);
nor U3197 (N_3197,In_594,In_712);
nand U3198 (N_3198,In_798,In_58);
and U3199 (N_3199,In_770,In_862);
nor U3200 (N_3200,In_532,In_716);
nor U3201 (N_3201,In_111,In_18);
or U3202 (N_3202,In_289,In_398);
nor U3203 (N_3203,In_299,In_149);
nor U3204 (N_3204,In_504,In_27);
nand U3205 (N_3205,In_372,In_987);
and U3206 (N_3206,In_145,In_544);
or U3207 (N_3207,In_916,In_443);
xnor U3208 (N_3208,In_337,In_317);
and U3209 (N_3209,In_763,In_729);
or U3210 (N_3210,In_28,In_367);
or U3211 (N_3211,In_354,In_355);
or U3212 (N_3212,In_833,In_415);
xnor U3213 (N_3213,In_411,In_180);
or U3214 (N_3214,In_694,In_434);
xnor U3215 (N_3215,In_827,In_133);
and U3216 (N_3216,In_625,In_491);
or U3217 (N_3217,In_341,In_816);
nor U3218 (N_3218,In_440,In_198);
nand U3219 (N_3219,In_967,In_808);
or U3220 (N_3220,In_178,In_205);
xnor U3221 (N_3221,In_197,In_162);
or U3222 (N_3222,In_307,In_975);
nand U3223 (N_3223,In_779,In_65);
or U3224 (N_3224,In_182,In_810);
and U3225 (N_3225,In_862,In_49);
or U3226 (N_3226,In_347,In_620);
xor U3227 (N_3227,In_804,In_486);
xnor U3228 (N_3228,In_754,In_810);
or U3229 (N_3229,In_814,In_635);
nor U3230 (N_3230,In_964,In_836);
nor U3231 (N_3231,In_665,In_218);
xnor U3232 (N_3232,In_126,In_48);
or U3233 (N_3233,In_549,In_738);
or U3234 (N_3234,In_491,In_917);
xnor U3235 (N_3235,In_555,In_646);
nor U3236 (N_3236,In_921,In_429);
xor U3237 (N_3237,In_64,In_543);
and U3238 (N_3238,In_216,In_647);
xor U3239 (N_3239,In_761,In_257);
nor U3240 (N_3240,In_139,In_201);
xor U3241 (N_3241,In_803,In_293);
and U3242 (N_3242,In_587,In_339);
nand U3243 (N_3243,In_9,In_930);
xor U3244 (N_3244,In_41,In_351);
nor U3245 (N_3245,In_292,In_300);
xor U3246 (N_3246,In_432,In_299);
and U3247 (N_3247,In_875,In_919);
or U3248 (N_3248,In_612,In_745);
and U3249 (N_3249,In_630,In_488);
or U3250 (N_3250,In_833,In_350);
nor U3251 (N_3251,In_542,In_210);
xnor U3252 (N_3252,In_580,In_72);
nand U3253 (N_3253,In_887,In_902);
and U3254 (N_3254,In_988,In_43);
nor U3255 (N_3255,In_746,In_17);
and U3256 (N_3256,In_343,In_36);
xor U3257 (N_3257,In_722,In_546);
nand U3258 (N_3258,In_294,In_203);
and U3259 (N_3259,In_188,In_767);
xor U3260 (N_3260,In_254,In_900);
or U3261 (N_3261,In_395,In_411);
xor U3262 (N_3262,In_874,In_124);
xor U3263 (N_3263,In_856,In_412);
nor U3264 (N_3264,In_109,In_730);
xor U3265 (N_3265,In_896,In_767);
nor U3266 (N_3266,In_312,In_826);
xor U3267 (N_3267,In_215,In_928);
xor U3268 (N_3268,In_473,In_457);
xor U3269 (N_3269,In_117,In_962);
nor U3270 (N_3270,In_101,In_968);
xor U3271 (N_3271,In_475,In_756);
nor U3272 (N_3272,In_534,In_888);
and U3273 (N_3273,In_985,In_660);
nor U3274 (N_3274,In_694,In_882);
xnor U3275 (N_3275,In_383,In_949);
nor U3276 (N_3276,In_1,In_410);
nor U3277 (N_3277,In_582,In_195);
and U3278 (N_3278,In_434,In_349);
and U3279 (N_3279,In_402,In_743);
or U3280 (N_3280,In_992,In_118);
or U3281 (N_3281,In_536,In_876);
xor U3282 (N_3282,In_960,In_940);
xnor U3283 (N_3283,In_894,In_435);
or U3284 (N_3284,In_279,In_831);
or U3285 (N_3285,In_816,In_343);
or U3286 (N_3286,In_328,In_717);
or U3287 (N_3287,In_797,In_535);
xor U3288 (N_3288,In_912,In_103);
nor U3289 (N_3289,In_823,In_345);
xor U3290 (N_3290,In_512,In_92);
nor U3291 (N_3291,In_256,In_148);
nand U3292 (N_3292,In_218,In_483);
nand U3293 (N_3293,In_26,In_961);
or U3294 (N_3294,In_501,In_652);
and U3295 (N_3295,In_270,In_176);
and U3296 (N_3296,In_320,In_721);
and U3297 (N_3297,In_432,In_628);
and U3298 (N_3298,In_823,In_379);
nor U3299 (N_3299,In_238,In_679);
and U3300 (N_3300,In_834,In_732);
or U3301 (N_3301,In_242,In_979);
xor U3302 (N_3302,In_603,In_79);
and U3303 (N_3303,In_535,In_437);
or U3304 (N_3304,In_46,In_751);
and U3305 (N_3305,In_166,In_772);
xnor U3306 (N_3306,In_443,In_859);
nor U3307 (N_3307,In_896,In_525);
nor U3308 (N_3308,In_240,In_408);
or U3309 (N_3309,In_559,In_305);
and U3310 (N_3310,In_868,In_57);
or U3311 (N_3311,In_603,In_378);
nor U3312 (N_3312,In_213,In_979);
nor U3313 (N_3313,In_64,In_176);
nor U3314 (N_3314,In_672,In_581);
or U3315 (N_3315,In_529,In_12);
or U3316 (N_3316,In_510,In_145);
nand U3317 (N_3317,In_244,In_705);
or U3318 (N_3318,In_213,In_231);
and U3319 (N_3319,In_218,In_973);
or U3320 (N_3320,In_914,In_636);
xor U3321 (N_3321,In_39,In_319);
xnor U3322 (N_3322,In_975,In_895);
nor U3323 (N_3323,In_977,In_963);
and U3324 (N_3324,In_263,In_205);
xor U3325 (N_3325,In_389,In_567);
nor U3326 (N_3326,In_546,In_822);
xor U3327 (N_3327,In_657,In_970);
nand U3328 (N_3328,In_516,In_152);
and U3329 (N_3329,In_98,In_674);
or U3330 (N_3330,In_18,In_301);
xor U3331 (N_3331,In_176,In_18);
nand U3332 (N_3332,In_429,In_706);
nand U3333 (N_3333,In_389,In_603);
and U3334 (N_3334,In_527,In_878);
or U3335 (N_3335,In_363,In_844);
and U3336 (N_3336,In_719,In_930);
nand U3337 (N_3337,In_325,In_427);
nor U3338 (N_3338,In_403,In_163);
nor U3339 (N_3339,In_11,In_987);
and U3340 (N_3340,In_736,In_807);
xor U3341 (N_3341,In_987,In_260);
nand U3342 (N_3342,In_734,In_981);
nor U3343 (N_3343,In_626,In_470);
nand U3344 (N_3344,In_216,In_825);
and U3345 (N_3345,In_339,In_612);
and U3346 (N_3346,In_556,In_887);
xnor U3347 (N_3347,In_295,In_926);
nor U3348 (N_3348,In_746,In_344);
and U3349 (N_3349,In_98,In_193);
and U3350 (N_3350,In_961,In_413);
and U3351 (N_3351,In_726,In_540);
nor U3352 (N_3352,In_756,In_697);
nand U3353 (N_3353,In_583,In_184);
and U3354 (N_3354,In_799,In_757);
nand U3355 (N_3355,In_460,In_550);
and U3356 (N_3356,In_992,In_900);
nand U3357 (N_3357,In_880,In_965);
xor U3358 (N_3358,In_36,In_46);
xor U3359 (N_3359,In_937,In_741);
xor U3360 (N_3360,In_1,In_462);
nand U3361 (N_3361,In_421,In_158);
nand U3362 (N_3362,In_835,In_711);
xor U3363 (N_3363,In_430,In_690);
xnor U3364 (N_3364,In_998,In_999);
or U3365 (N_3365,In_243,In_899);
nand U3366 (N_3366,In_2,In_859);
nand U3367 (N_3367,In_52,In_372);
nand U3368 (N_3368,In_899,In_410);
xnor U3369 (N_3369,In_950,In_703);
nand U3370 (N_3370,In_173,In_962);
nand U3371 (N_3371,In_110,In_528);
and U3372 (N_3372,In_51,In_178);
nand U3373 (N_3373,In_858,In_529);
or U3374 (N_3374,In_991,In_811);
and U3375 (N_3375,In_875,In_414);
nor U3376 (N_3376,In_481,In_669);
nor U3377 (N_3377,In_562,In_527);
nand U3378 (N_3378,In_313,In_891);
or U3379 (N_3379,In_138,In_220);
nor U3380 (N_3380,In_409,In_575);
and U3381 (N_3381,In_35,In_503);
or U3382 (N_3382,In_755,In_614);
and U3383 (N_3383,In_432,In_331);
nor U3384 (N_3384,In_901,In_53);
xnor U3385 (N_3385,In_409,In_24);
nand U3386 (N_3386,In_642,In_225);
nand U3387 (N_3387,In_748,In_909);
nor U3388 (N_3388,In_7,In_536);
or U3389 (N_3389,In_854,In_369);
nor U3390 (N_3390,In_480,In_193);
nor U3391 (N_3391,In_602,In_10);
or U3392 (N_3392,In_67,In_698);
or U3393 (N_3393,In_120,In_604);
nand U3394 (N_3394,In_9,In_904);
and U3395 (N_3395,In_567,In_850);
xor U3396 (N_3396,In_281,In_479);
or U3397 (N_3397,In_775,In_898);
and U3398 (N_3398,In_410,In_131);
nor U3399 (N_3399,In_530,In_201);
nor U3400 (N_3400,In_814,In_700);
and U3401 (N_3401,In_778,In_702);
nand U3402 (N_3402,In_364,In_569);
nor U3403 (N_3403,In_828,In_863);
and U3404 (N_3404,In_734,In_834);
xnor U3405 (N_3405,In_865,In_80);
nand U3406 (N_3406,In_106,In_566);
nand U3407 (N_3407,In_168,In_140);
xor U3408 (N_3408,In_721,In_732);
nor U3409 (N_3409,In_700,In_553);
nor U3410 (N_3410,In_579,In_849);
and U3411 (N_3411,In_842,In_97);
nor U3412 (N_3412,In_858,In_818);
nand U3413 (N_3413,In_28,In_705);
nand U3414 (N_3414,In_808,In_770);
xnor U3415 (N_3415,In_741,In_210);
and U3416 (N_3416,In_232,In_516);
and U3417 (N_3417,In_467,In_511);
and U3418 (N_3418,In_76,In_995);
xnor U3419 (N_3419,In_38,In_809);
xor U3420 (N_3420,In_668,In_941);
and U3421 (N_3421,In_781,In_837);
nand U3422 (N_3422,In_389,In_961);
xnor U3423 (N_3423,In_563,In_71);
or U3424 (N_3424,In_613,In_57);
or U3425 (N_3425,In_954,In_493);
nand U3426 (N_3426,In_565,In_24);
and U3427 (N_3427,In_39,In_246);
nor U3428 (N_3428,In_879,In_286);
or U3429 (N_3429,In_45,In_130);
and U3430 (N_3430,In_313,In_451);
nor U3431 (N_3431,In_956,In_670);
or U3432 (N_3432,In_88,In_669);
xnor U3433 (N_3433,In_10,In_663);
nor U3434 (N_3434,In_225,In_515);
or U3435 (N_3435,In_648,In_502);
nand U3436 (N_3436,In_430,In_836);
or U3437 (N_3437,In_379,In_380);
or U3438 (N_3438,In_218,In_415);
and U3439 (N_3439,In_154,In_10);
xnor U3440 (N_3440,In_578,In_340);
nor U3441 (N_3441,In_790,In_707);
and U3442 (N_3442,In_482,In_959);
and U3443 (N_3443,In_304,In_742);
xnor U3444 (N_3444,In_571,In_391);
nand U3445 (N_3445,In_300,In_247);
nor U3446 (N_3446,In_576,In_567);
and U3447 (N_3447,In_829,In_128);
xor U3448 (N_3448,In_494,In_533);
or U3449 (N_3449,In_269,In_646);
and U3450 (N_3450,In_247,In_174);
nand U3451 (N_3451,In_965,In_695);
xor U3452 (N_3452,In_459,In_676);
nand U3453 (N_3453,In_511,In_245);
xor U3454 (N_3454,In_478,In_355);
nand U3455 (N_3455,In_80,In_869);
xnor U3456 (N_3456,In_850,In_653);
or U3457 (N_3457,In_363,In_803);
nor U3458 (N_3458,In_533,In_275);
and U3459 (N_3459,In_84,In_532);
nor U3460 (N_3460,In_191,In_354);
nor U3461 (N_3461,In_889,In_282);
or U3462 (N_3462,In_201,In_351);
nand U3463 (N_3463,In_784,In_574);
nand U3464 (N_3464,In_54,In_174);
nand U3465 (N_3465,In_6,In_739);
xnor U3466 (N_3466,In_687,In_325);
nand U3467 (N_3467,In_853,In_994);
or U3468 (N_3468,In_239,In_667);
or U3469 (N_3469,In_902,In_934);
nor U3470 (N_3470,In_16,In_303);
and U3471 (N_3471,In_384,In_388);
xnor U3472 (N_3472,In_441,In_605);
xnor U3473 (N_3473,In_777,In_941);
nand U3474 (N_3474,In_919,In_229);
xor U3475 (N_3475,In_474,In_434);
nand U3476 (N_3476,In_481,In_584);
or U3477 (N_3477,In_222,In_513);
or U3478 (N_3478,In_303,In_276);
and U3479 (N_3479,In_301,In_887);
nor U3480 (N_3480,In_466,In_293);
nand U3481 (N_3481,In_85,In_543);
nor U3482 (N_3482,In_986,In_968);
or U3483 (N_3483,In_92,In_53);
and U3484 (N_3484,In_443,In_41);
nor U3485 (N_3485,In_264,In_799);
or U3486 (N_3486,In_964,In_954);
xor U3487 (N_3487,In_859,In_453);
and U3488 (N_3488,In_628,In_842);
nor U3489 (N_3489,In_411,In_636);
and U3490 (N_3490,In_359,In_283);
nand U3491 (N_3491,In_312,In_253);
nor U3492 (N_3492,In_429,In_806);
and U3493 (N_3493,In_775,In_709);
or U3494 (N_3494,In_778,In_630);
or U3495 (N_3495,In_625,In_922);
nor U3496 (N_3496,In_917,In_628);
and U3497 (N_3497,In_920,In_170);
xnor U3498 (N_3498,In_895,In_330);
nand U3499 (N_3499,In_767,In_126);
nor U3500 (N_3500,In_132,In_481);
or U3501 (N_3501,In_269,In_393);
xor U3502 (N_3502,In_514,In_345);
nand U3503 (N_3503,In_768,In_285);
nor U3504 (N_3504,In_985,In_662);
nor U3505 (N_3505,In_753,In_726);
nand U3506 (N_3506,In_80,In_723);
and U3507 (N_3507,In_830,In_990);
or U3508 (N_3508,In_57,In_750);
or U3509 (N_3509,In_822,In_308);
nand U3510 (N_3510,In_561,In_122);
nand U3511 (N_3511,In_859,In_479);
and U3512 (N_3512,In_775,In_652);
xnor U3513 (N_3513,In_565,In_789);
nand U3514 (N_3514,In_223,In_238);
xnor U3515 (N_3515,In_504,In_666);
nand U3516 (N_3516,In_851,In_736);
or U3517 (N_3517,In_663,In_986);
or U3518 (N_3518,In_907,In_382);
or U3519 (N_3519,In_165,In_750);
xor U3520 (N_3520,In_242,In_55);
and U3521 (N_3521,In_174,In_914);
xnor U3522 (N_3522,In_559,In_70);
or U3523 (N_3523,In_862,In_636);
nor U3524 (N_3524,In_345,In_89);
nand U3525 (N_3525,In_362,In_55);
xor U3526 (N_3526,In_364,In_868);
and U3527 (N_3527,In_305,In_188);
nand U3528 (N_3528,In_922,In_547);
nor U3529 (N_3529,In_555,In_817);
or U3530 (N_3530,In_950,In_469);
and U3531 (N_3531,In_874,In_138);
nand U3532 (N_3532,In_472,In_69);
xor U3533 (N_3533,In_983,In_30);
nand U3534 (N_3534,In_998,In_600);
xnor U3535 (N_3535,In_648,In_993);
and U3536 (N_3536,In_994,In_239);
and U3537 (N_3537,In_129,In_46);
nor U3538 (N_3538,In_342,In_118);
and U3539 (N_3539,In_814,In_323);
xor U3540 (N_3540,In_297,In_435);
nor U3541 (N_3541,In_623,In_708);
nand U3542 (N_3542,In_650,In_588);
nand U3543 (N_3543,In_443,In_950);
nand U3544 (N_3544,In_822,In_652);
and U3545 (N_3545,In_11,In_365);
xnor U3546 (N_3546,In_991,In_858);
nor U3547 (N_3547,In_458,In_407);
or U3548 (N_3548,In_457,In_972);
or U3549 (N_3549,In_45,In_745);
and U3550 (N_3550,In_42,In_351);
nand U3551 (N_3551,In_519,In_345);
or U3552 (N_3552,In_372,In_522);
xnor U3553 (N_3553,In_97,In_326);
nor U3554 (N_3554,In_666,In_989);
nand U3555 (N_3555,In_9,In_228);
and U3556 (N_3556,In_323,In_760);
nand U3557 (N_3557,In_845,In_296);
nand U3558 (N_3558,In_441,In_326);
and U3559 (N_3559,In_74,In_996);
or U3560 (N_3560,In_3,In_544);
or U3561 (N_3561,In_459,In_192);
nand U3562 (N_3562,In_647,In_856);
nand U3563 (N_3563,In_336,In_986);
xor U3564 (N_3564,In_699,In_420);
or U3565 (N_3565,In_554,In_790);
nor U3566 (N_3566,In_518,In_111);
or U3567 (N_3567,In_466,In_885);
or U3568 (N_3568,In_629,In_891);
nand U3569 (N_3569,In_132,In_202);
nand U3570 (N_3570,In_226,In_76);
nand U3571 (N_3571,In_985,In_498);
nand U3572 (N_3572,In_404,In_158);
xnor U3573 (N_3573,In_620,In_234);
and U3574 (N_3574,In_225,In_527);
or U3575 (N_3575,In_143,In_858);
or U3576 (N_3576,In_153,In_344);
nor U3577 (N_3577,In_523,In_435);
nor U3578 (N_3578,In_724,In_118);
nor U3579 (N_3579,In_604,In_263);
and U3580 (N_3580,In_751,In_414);
xor U3581 (N_3581,In_889,In_953);
and U3582 (N_3582,In_422,In_933);
and U3583 (N_3583,In_929,In_583);
xnor U3584 (N_3584,In_613,In_487);
and U3585 (N_3585,In_972,In_981);
nor U3586 (N_3586,In_105,In_981);
and U3587 (N_3587,In_737,In_437);
xnor U3588 (N_3588,In_398,In_60);
xnor U3589 (N_3589,In_643,In_839);
xor U3590 (N_3590,In_780,In_755);
nor U3591 (N_3591,In_672,In_490);
and U3592 (N_3592,In_693,In_984);
or U3593 (N_3593,In_496,In_300);
nor U3594 (N_3594,In_489,In_469);
and U3595 (N_3595,In_871,In_583);
nor U3596 (N_3596,In_479,In_911);
xor U3597 (N_3597,In_220,In_23);
or U3598 (N_3598,In_524,In_901);
and U3599 (N_3599,In_340,In_479);
nand U3600 (N_3600,In_656,In_380);
or U3601 (N_3601,In_378,In_309);
xor U3602 (N_3602,In_891,In_108);
and U3603 (N_3603,In_379,In_25);
or U3604 (N_3604,In_806,In_386);
and U3605 (N_3605,In_912,In_93);
nand U3606 (N_3606,In_349,In_445);
nand U3607 (N_3607,In_142,In_391);
and U3608 (N_3608,In_497,In_213);
nor U3609 (N_3609,In_621,In_863);
and U3610 (N_3610,In_846,In_897);
nor U3611 (N_3611,In_591,In_522);
or U3612 (N_3612,In_752,In_812);
nor U3613 (N_3613,In_85,In_549);
or U3614 (N_3614,In_545,In_908);
or U3615 (N_3615,In_171,In_228);
or U3616 (N_3616,In_37,In_490);
nand U3617 (N_3617,In_253,In_132);
nor U3618 (N_3618,In_461,In_856);
nor U3619 (N_3619,In_750,In_119);
or U3620 (N_3620,In_321,In_843);
nand U3621 (N_3621,In_263,In_560);
and U3622 (N_3622,In_475,In_979);
and U3623 (N_3623,In_169,In_171);
xnor U3624 (N_3624,In_4,In_218);
nand U3625 (N_3625,In_838,In_715);
nand U3626 (N_3626,In_0,In_883);
xnor U3627 (N_3627,In_496,In_763);
and U3628 (N_3628,In_873,In_621);
nand U3629 (N_3629,In_325,In_664);
nand U3630 (N_3630,In_233,In_666);
or U3631 (N_3631,In_464,In_391);
nand U3632 (N_3632,In_851,In_504);
or U3633 (N_3633,In_685,In_383);
xnor U3634 (N_3634,In_804,In_829);
nor U3635 (N_3635,In_543,In_975);
xnor U3636 (N_3636,In_181,In_81);
xnor U3637 (N_3637,In_705,In_485);
nor U3638 (N_3638,In_687,In_216);
or U3639 (N_3639,In_89,In_29);
xor U3640 (N_3640,In_531,In_103);
or U3641 (N_3641,In_875,In_348);
and U3642 (N_3642,In_177,In_381);
xor U3643 (N_3643,In_150,In_163);
or U3644 (N_3644,In_643,In_818);
and U3645 (N_3645,In_47,In_372);
nand U3646 (N_3646,In_84,In_699);
nand U3647 (N_3647,In_543,In_462);
and U3648 (N_3648,In_403,In_121);
or U3649 (N_3649,In_635,In_665);
nor U3650 (N_3650,In_635,In_7);
and U3651 (N_3651,In_963,In_244);
xnor U3652 (N_3652,In_683,In_202);
or U3653 (N_3653,In_718,In_317);
and U3654 (N_3654,In_242,In_531);
nand U3655 (N_3655,In_378,In_984);
xor U3656 (N_3656,In_196,In_479);
nor U3657 (N_3657,In_994,In_964);
nor U3658 (N_3658,In_139,In_173);
and U3659 (N_3659,In_751,In_247);
nor U3660 (N_3660,In_787,In_183);
nor U3661 (N_3661,In_449,In_70);
xor U3662 (N_3662,In_714,In_991);
nand U3663 (N_3663,In_606,In_820);
nand U3664 (N_3664,In_198,In_484);
nor U3665 (N_3665,In_994,In_110);
nor U3666 (N_3666,In_446,In_654);
nor U3667 (N_3667,In_459,In_531);
nand U3668 (N_3668,In_310,In_879);
nor U3669 (N_3669,In_602,In_984);
nor U3670 (N_3670,In_87,In_826);
nor U3671 (N_3671,In_803,In_890);
nand U3672 (N_3672,In_659,In_942);
or U3673 (N_3673,In_263,In_593);
nor U3674 (N_3674,In_567,In_354);
or U3675 (N_3675,In_151,In_725);
or U3676 (N_3676,In_607,In_573);
or U3677 (N_3677,In_571,In_809);
xnor U3678 (N_3678,In_158,In_326);
and U3679 (N_3679,In_116,In_249);
and U3680 (N_3680,In_504,In_299);
or U3681 (N_3681,In_338,In_377);
and U3682 (N_3682,In_225,In_999);
and U3683 (N_3683,In_664,In_133);
nor U3684 (N_3684,In_190,In_467);
nor U3685 (N_3685,In_561,In_883);
xnor U3686 (N_3686,In_84,In_827);
nand U3687 (N_3687,In_25,In_382);
nand U3688 (N_3688,In_562,In_118);
or U3689 (N_3689,In_924,In_266);
xor U3690 (N_3690,In_396,In_604);
and U3691 (N_3691,In_347,In_707);
nor U3692 (N_3692,In_942,In_262);
nand U3693 (N_3693,In_287,In_321);
and U3694 (N_3694,In_283,In_447);
and U3695 (N_3695,In_771,In_716);
and U3696 (N_3696,In_184,In_697);
xnor U3697 (N_3697,In_821,In_436);
or U3698 (N_3698,In_53,In_117);
nor U3699 (N_3699,In_792,In_717);
nand U3700 (N_3700,In_127,In_643);
and U3701 (N_3701,In_439,In_670);
and U3702 (N_3702,In_966,In_209);
nor U3703 (N_3703,In_290,In_277);
xnor U3704 (N_3704,In_144,In_42);
xor U3705 (N_3705,In_154,In_311);
nand U3706 (N_3706,In_24,In_406);
and U3707 (N_3707,In_210,In_582);
or U3708 (N_3708,In_582,In_211);
nand U3709 (N_3709,In_859,In_478);
and U3710 (N_3710,In_42,In_330);
nand U3711 (N_3711,In_941,In_885);
xor U3712 (N_3712,In_591,In_178);
nand U3713 (N_3713,In_690,In_974);
xor U3714 (N_3714,In_155,In_655);
xor U3715 (N_3715,In_701,In_30);
or U3716 (N_3716,In_416,In_307);
and U3717 (N_3717,In_280,In_854);
and U3718 (N_3718,In_112,In_969);
nand U3719 (N_3719,In_269,In_443);
xnor U3720 (N_3720,In_92,In_136);
or U3721 (N_3721,In_747,In_663);
and U3722 (N_3722,In_574,In_995);
xor U3723 (N_3723,In_48,In_40);
nand U3724 (N_3724,In_25,In_805);
xnor U3725 (N_3725,In_140,In_31);
nand U3726 (N_3726,In_866,In_296);
and U3727 (N_3727,In_304,In_449);
and U3728 (N_3728,In_135,In_485);
nand U3729 (N_3729,In_943,In_629);
or U3730 (N_3730,In_598,In_563);
or U3731 (N_3731,In_952,In_592);
nand U3732 (N_3732,In_96,In_994);
or U3733 (N_3733,In_976,In_682);
nand U3734 (N_3734,In_615,In_395);
xor U3735 (N_3735,In_985,In_410);
nand U3736 (N_3736,In_505,In_571);
or U3737 (N_3737,In_225,In_4);
and U3738 (N_3738,In_965,In_461);
or U3739 (N_3739,In_291,In_767);
xor U3740 (N_3740,In_862,In_575);
nor U3741 (N_3741,In_939,In_290);
nor U3742 (N_3742,In_709,In_372);
and U3743 (N_3743,In_377,In_503);
or U3744 (N_3744,In_218,In_322);
or U3745 (N_3745,In_937,In_247);
xor U3746 (N_3746,In_10,In_743);
nand U3747 (N_3747,In_39,In_420);
nand U3748 (N_3748,In_208,In_787);
xor U3749 (N_3749,In_674,In_857);
nor U3750 (N_3750,In_123,In_855);
xnor U3751 (N_3751,In_551,In_975);
nand U3752 (N_3752,In_613,In_754);
nor U3753 (N_3753,In_29,In_748);
xnor U3754 (N_3754,In_532,In_241);
nor U3755 (N_3755,In_430,In_367);
xor U3756 (N_3756,In_540,In_435);
and U3757 (N_3757,In_696,In_647);
xor U3758 (N_3758,In_382,In_811);
nand U3759 (N_3759,In_336,In_518);
nand U3760 (N_3760,In_575,In_707);
nor U3761 (N_3761,In_38,In_68);
nand U3762 (N_3762,In_19,In_119);
nor U3763 (N_3763,In_923,In_588);
nand U3764 (N_3764,In_784,In_554);
nor U3765 (N_3765,In_186,In_732);
or U3766 (N_3766,In_779,In_347);
xnor U3767 (N_3767,In_914,In_928);
or U3768 (N_3768,In_30,In_497);
and U3769 (N_3769,In_721,In_854);
nand U3770 (N_3770,In_481,In_981);
or U3771 (N_3771,In_237,In_964);
or U3772 (N_3772,In_306,In_866);
nor U3773 (N_3773,In_346,In_712);
or U3774 (N_3774,In_952,In_494);
xnor U3775 (N_3775,In_789,In_233);
nor U3776 (N_3776,In_433,In_724);
xnor U3777 (N_3777,In_685,In_45);
nor U3778 (N_3778,In_23,In_505);
or U3779 (N_3779,In_270,In_525);
and U3780 (N_3780,In_757,In_555);
nand U3781 (N_3781,In_349,In_628);
nor U3782 (N_3782,In_599,In_778);
xor U3783 (N_3783,In_556,In_603);
nand U3784 (N_3784,In_523,In_105);
or U3785 (N_3785,In_290,In_370);
and U3786 (N_3786,In_723,In_282);
and U3787 (N_3787,In_883,In_573);
nand U3788 (N_3788,In_663,In_755);
or U3789 (N_3789,In_745,In_139);
nand U3790 (N_3790,In_601,In_160);
nor U3791 (N_3791,In_292,In_569);
xor U3792 (N_3792,In_524,In_847);
nand U3793 (N_3793,In_738,In_450);
and U3794 (N_3794,In_708,In_306);
or U3795 (N_3795,In_156,In_444);
and U3796 (N_3796,In_497,In_215);
nand U3797 (N_3797,In_54,In_560);
and U3798 (N_3798,In_171,In_57);
nand U3799 (N_3799,In_573,In_917);
nor U3800 (N_3800,In_798,In_394);
or U3801 (N_3801,In_151,In_734);
nor U3802 (N_3802,In_370,In_887);
or U3803 (N_3803,In_275,In_55);
nand U3804 (N_3804,In_507,In_783);
nand U3805 (N_3805,In_321,In_770);
xnor U3806 (N_3806,In_432,In_931);
or U3807 (N_3807,In_602,In_4);
nor U3808 (N_3808,In_252,In_355);
xnor U3809 (N_3809,In_305,In_726);
or U3810 (N_3810,In_803,In_401);
or U3811 (N_3811,In_546,In_248);
nand U3812 (N_3812,In_323,In_223);
or U3813 (N_3813,In_405,In_38);
nand U3814 (N_3814,In_475,In_179);
xnor U3815 (N_3815,In_446,In_322);
nand U3816 (N_3816,In_175,In_694);
or U3817 (N_3817,In_897,In_516);
nand U3818 (N_3818,In_243,In_385);
xnor U3819 (N_3819,In_845,In_702);
xnor U3820 (N_3820,In_374,In_340);
nor U3821 (N_3821,In_282,In_756);
xnor U3822 (N_3822,In_528,In_688);
nor U3823 (N_3823,In_195,In_465);
and U3824 (N_3824,In_7,In_418);
nand U3825 (N_3825,In_980,In_761);
and U3826 (N_3826,In_969,In_51);
xnor U3827 (N_3827,In_907,In_934);
nand U3828 (N_3828,In_446,In_993);
nand U3829 (N_3829,In_334,In_198);
or U3830 (N_3830,In_9,In_798);
nor U3831 (N_3831,In_547,In_67);
nand U3832 (N_3832,In_57,In_98);
nand U3833 (N_3833,In_784,In_825);
or U3834 (N_3834,In_477,In_687);
xor U3835 (N_3835,In_101,In_690);
and U3836 (N_3836,In_521,In_951);
xor U3837 (N_3837,In_671,In_350);
and U3838 (N_3838,In_854,In_407);
or U3839 (N_3839,In_462,In_485);
or U3840 (N_3840,In_479,In_798);
and U3841 (N_3841,In_52,In_41);
nand U3842 (N_3842,In_177,In_671);
nor U3843 (N_3843,In_513,In_381);
nor U3844 (N_3844,In_344,In_922);
nand U3845 (N_3845,In_741,In_129);
and U3846 (N_3846,In_136,In_889);
or U3847 (N_3847,In_66,In_435);
nand U3848 (N_3848,In_297,In_31);
or U3849 (N_3849,In_115,In_785);
nand U3850 (N_3850,In_342,In_719);
and U3851 (N_3851,In_443,In_772);
nor U3852 (N_3852,In_184,In_946);
and U3853 (N_3853,In_299,In_296);
or U3854 (N_3854,In_262,In_366);
xor U3855 (N_3855,In_762,In_942);
and U3856 (N_3856,In_555,In_703);
or U3857 (N_3857,In_401,In_929);
nand U3858 (N_3858,In_557,In_837);
xor U3859 (N_3859,In_799,In_77);
nand U3860 (N_3860,In_372,In_195);
and U3861 (N_3861,In_676,In_791);
nand U3862 (N_3862,In_279,In_479);
xnor U3863 (N_3863,In_427,In_476);
nand U3864 (N_3864,In_474,In_941);
and U3865 (N_3865,In_967,In_118);
nand U3866 (N_3866,In_900,In_222);
xor U3867 (N_3867,In_192,In_148);
or U3868 (N_3868,In_395,In_71);
or U3869 (N_3869,In_506,In_488);
xor U3870 (N_3870,In_46,In_577);
nand U3871 (N_3871,In_168,In_944);
nand U3872 (N_3872,In_56,In_648);
nand U3873 (N_3873,In_779,In_248);
or U3874 (N_3874,In_445,In_518);
nor U3875 (N_3875,In_633,In_301);
nand U3876 (N_3876,In_190,In_668);
nand U3877 (N_3877,In_773,In_807);
nand U3878 (N_3878,In_850,In_229);
or U3879 (N_3879,In_589,In_221);
nand U3880 (N_3880,In_655,In_428);
xnor U3881 (N_3881,In_296,In_927);
nand U3882 (N_3882,In_430,In_2);
nor U3883 (N_3883,In_402,In_211);
and U3884 (N_3884,In_26,In_335);
xor U3885 (N_3885,In_26,In_176);
nor U3886 (N_3886,In_773,In_657);
or U3887 (N_3887,In_532,In_681);
nor U3888 (N_3888,In_334,In_151);
nand U3889 (N_3889,In_772,In_822);
nand U3890 (N_3890,In_42,In_347);
nor U3891 (N_3891,In_179,In_194);
nand U3892 (N_3892,In_159,In_836);
nand U3893 (N_3893,In_440,In_574);
or U3894 (N_3894,In_251,In_103);
or U3895 (N_3895,In_966,In_490);
xnor U3896 (N_3896,In_874,In_456);
nand U3897 (N_3897,In_5,In_1);
nor U3898 (N_3898,In_416,In_73);
xnor U3899 (N_3899,In_70,In_248);
nor U3900 (N_3900,In_439,In_730);
or U3901 (N_3901,In_225,In_26);
nand U3902 (N_3902,In_164,In_913);
nor U3903 (N_3903,In_0,In_752);
and U3904 (N_3904,In_408,In_195);
or U3905 (N_3905,In_330,In_101);
or U3906 (N_3906,In_570,In_539);
or U3907 (N_3907,In_625,In_636);
and U3908 (N_3908,In_311,In_331);
nor U3909 (N_3909,In_789,In_384);
xor U3910 (N_3910,In_490,In_922);
nand U3911 (N_3911,In_206,In_774);
nor U3912 (N_3912,In_175,In_103);
and U3913 (N_3913,In_305,In_708);
xor U3914 (N_3914,In_902,In_154);
xor U3915 (N_3915,In_225,In_601);
and U3916 (N_3916,In_611,In_234);
nand U3917 (N_3917,In_457,In_78);
nor U3918 (N_3918,In_294,In_433);
xor U3919 (N_3919,In_66,In_249);
nor U3920 (N_3920,In_928,In_150);
or U3921 (N_3921,In_421,In_886);
and U3922 (N_3922,In_406,In_469);
xor U3923 (N_3923,In_131,In_43);
xor U3924 (N_3924,In_425,In_291);
and U3925 (N_3925,In_361,In_992);
and U3926 (N_3926,In_540,In_475);
nor U3927 (N_3927,In_100,In_475);
nor U3928 (N_3928,In_622,In_684);
or U3929 (N_3929,In_95,In_733);
xnor U3930 (N_3930,In_646,In_978);
nand U3931 (N_3931,In_463,In_750);
nand U3932 (N_3932,In_94,In_283);
and U3933 (N_3933,In_913,In_21);
nor U3934 (N_3934,In_73,In_600);
and U3935 (N_3935,In_251,In_769);
nor U3936 (N_3936,In_524,In_320);
nand U3937 (N_3937,In_815,In_340);
nand U3938 (N_3938,In_236,In_214);
and U3939 (N_3939,In_552,In_927);
or U3940 (N_3940,In_582,In_869);
or U3941 (N_3941,In_550,In_462);
and U3942 (N_3942,In_949,In_829);
xnor U3943 (N_3943,In_10,In_796);
or U3944 (N_3944,In_197,In_993);
and U3945 (N_3945,In_839,In_836);
or U3946 (N_3946,In_608,In_471);
xor U3947 (N_3947,In_111,In_663);
or U3948 (N_3948,In_334,In_384);
nand U3949 (N_3949,In_602,In_821);
or U3950 (N_3950,In_613,In_158);
nor U3951 (N_3951,In_723,In_24);
or U3952 (N_3952,In_612,In_447);
and U3953 (N_3953,In_479,In_404);
and U3954 (N_3954,In_370,In_641);
and U3955 (N_3955,In_762,In_963);
nand U3956 (N_3956,In_247,In_944);
nand U3957 (N_3957,In_415,In_488);
nor U3958 (N_3958,In_241,In_23);
nand U3959 (N_3959,In_125,In_638);
and U3960 (N_3960,In_660,In_441);
and U3961 (N_3961,In_681,In_904);
or U3962 (N_3962,In_503,In_456);
nor U3963 (N_3963,In_125,In_995);
and U3964 (N_3964,In_302,In_776);
or U3965 (N_3965,In_447,In_122);
xnor U3966 (N_3966,In_864,In_780);
xnor U3967 (N_3967,In_494,In_960);
nor U3968 (N_3968,In_522,In_317);
nand U3969 (N_3969,In_637,In_623);
nor U3970 (N_3970,In_937,In_112);
and U3971 (N_3971,In_851,In_350);
xor U3972 (N_3972,In_936,In_932);
or U3973 (N_3973,In_952,In_172);
and U3974 (N_3974,In_477,In_499);
nand U3975 (N_3975,In_360,In_306);
or U3976 (N_3976,In_874,In_393);
and U3977 (N_3977,In_856,In_671);
nand U3978 (N_3978,In_717,In_812);
xnor U3979 (N_3979,In_281,In_994);
or U3980 (N_3980,In_945,In_747);
xnor U3981 (N_3981,In_241,In_746);
or U3982 (N_3982,In_28,In_885);
nor U3983 (N_3983,In_657,In_106);
nand U3984 (N_3984,In_802,In_686);
and U3985 (N_3985,In_833,In_293);
or U3986 (N_3986,In_516,In_722);
xnor U3987 (N_3987,In_579,In_76);
and U3988 (N_3988,In_986,In_974);
or U3989 (N_3989,In_807,In_531);
or U3990 (N_3990,In_759,In_4);
nand U3991 (N_3991,In_695,In_670);
or U3992 (N_3992,In_286,In_456);
and U3993 (N_3993,In_120,In_383);
or U3994 (N_3994,In_322,In_658);
or U3995 (N_3995,In_279,In_598);
and U3996 (N_3996,In_952,In_176);
or U3997 (N_3997,In_666,In_44);
nand U3998 (N_3998,In_728,In_61);
or U3999 (N_3999,In_877,In_718);
nor U4000 (N_4000,In_616,In_75);
xor U4001 (N_4001,In_897,In_57);
and U4002 (N_4002,In_66,In_770);
nor U4003 (N_4003,In_934,In_151);
or U4004 (N_4004,In_301,In_245);
nand U4005 (N_4005,In_987,In_608);
nand U4006 (N_4006,In_209,In_301);
nand U4007 (N_4007,In_759,In_679);
or U4008 (N_4008,In_558,In_433);
nor U4009 (N_4009,In_328,In_704);
and U4010 (N_4010,In_435,In_521);
nor U4011 (N_4011,In_63,In_11);
xnor U4012 (N_4012,In_455,In_37);
nand U4013 (N_4013,In_552,In_588);
or U4014 (N_4014,In_407,In_462);
nor U4015 (N_4015,In_849,In_922);
nor U4016 (N_4016,In_86,In_309);
nor U4017 (N_4017,In_461,In_660);
or U4018 (N_4018,In_469,In_313);
and U4019 (N_4019,In_702,In_93);
and U4020 (N_4020,In_921,In_945);
and U4021 (N_4021,In_465,In_991);
or U4022 (N_4022,In_432,In_476);
and U4023 (N_4023,In_432,In_698);
nor U4024 (N_4024,In_585,In_676);
and U4025 (N_4025,In_317,In_891);
nor U4026 (N_4026,In_874,In_879);
nand U4027 (N_4027,In_342,In_807);
xor U4028 (N_4028,In_979,In_726);
nor U4029 (N_4029,In_384,In_931);
xor U4030 (N_4030,In_637,In_495);
or U4031 (N_4031,In_10,In_626);
nand U4032 (N_4032,In_358,In_893);
nor U4033 (N_4033,In_628,In_392);
xnor U4034 (N_4034,In_66,In_261);
and U4035 (N_4035,In_870,In_590);
nand U4036 (N_4036,In_362,In_475);
xnor U4037 (N_4037,In_376,In_970);
nor U4038 (N_4038,In_656,In_341);
or U4039 (N_4039,In_613,In_447);
and U4040 (N_4040,In_215,In_654);
nor U4041 (N_4041,In_264,In_675);
xor U4042 (N_4042,In_500,In_260);
xor U4043 (N_4043,In_824,In_285);
or U4044 (N_4044,In_681,In_491);
nor U4045 (N_4045,In_778,In_556);
xor U4046 (N_4046,In_420,In_677);
nor U4047 (N_4047,In_635,In_706);
or U4048 (N_4048,In_543,In_203);
xnor U4049 (N_4049,In_15,In_104);
xnor U4050 (N_4050,In_178,In_39);
and U4051 (N_4051,In_884,In_50);
nor U4052 (N_4052,In_585,In_671);
and U4053 (N_4053,In_764,In_274);
or U4054 (N_4054,In_561,In_812);
nor U4055 (N_4055,In_602,In_51);
nor U4056 (N_4056,In_988,In_452);
or U4057 (N_4057,In_330,In_106);
and U4058 (N_4058,In_457,In_376);
or U4059 (N_4059,In_694,In_204);
nand U4060 (N_4060,In_909,In_500);
nand U4061 (N_4061,In_550,In_962);
nand U4062 (N_4062,In_825,In_960);
nor U4063 (N_4063,In_819,In_385);
xor U4064 (N_4064,In_208,In_841);
xor U4065 (N_4065,In_95,In_516);
and U4066 (N_4066,In_915,In_85);
nor U4067 (N_4067,In_464,In_661);
nor U4068 (N_4068,In_518,In_946);
and U4069 (N_4069,In_522,In_104);
or U4070 (N_4070,In_785,In_829);
and U4071 (N_4071,In_551,In_125);
nor U4072 (N_4072,In_736,In_573);
nor U4073 (N_4073,In_238,In_720);
xor U4074 (N_4074,In_988,In_441);
xor U4075 (N_4075,In_558,In_426);
or U4076 (N_4076,In_187,In_382);
nor U4077 (N_4077,In_273,In_286);
xor U4078 (N_4078,In_368,In_889);
or U4079 (N_4079,In_112,In_840);
xor U4080 (N_4080,In_148,In_488);
nand U4081 (N_4081,In_196,In_896);
and U4082 (N_4082,In_235,In_810);
or U4083 (N_4083,In_660,In_540);
nand U4084 (N_4084,In_545,In_128);
or U4085 (N_4085,In_33,In_802);
xnor U4086 (N_4086,In_432,In_294);
nor U4087 (N_4087,In_600,In_976);
and U4088 (N_4088,In_246,In_506);
and U4089 (N_4089,In_381,In_25);
and U4090 (N_4090,In_61,In_659);
nand U4091 (N_4091,In_822,In_252);
or U4092 (N_4092,In_783,In_823);
xnor U4093 (N_4093,In_473,In_994);
and U4094 (N_4094,In_937,In_68);
and U4095 (N_4095,In_745,In_144);
nor U4096 (N_4096,In_393,In_733);
and U4097 (N_4097,In_921,In_135);
nand U4098 (N_4098,In_532,In_599);
or U4099 (N_4099,In_595,In_866);
xnor U4100 (N_4100,In_875,In_963);
nand U4101 (N_4101,In_109,In_784);
or U4102 (N_4102,In_353,In_80);
nor U4103 (N_4103,In_59,In_833);
or U4104 (N_4104,In_94,In_488);
and U4105 (N_4105,In_909,In_430);
and U4106 (N_4106,In_721,In_339);
nand U4107 (N_4107,In_83,In_667);
nor U4108 (N_4108,In_111,In_775);
or U4109 (N_4109,In_682,In_173);
and U4110 (N_4110,In_62,In_36);
or U4111 (N_4111,In_288,In_131);
nor U4112 (N_4112,In_923,In_550);
nor U4113 (N_4113,In_256,In_796);
nand U4114 (N_4114,In_446,In_873);
xor U4115 (N_4115,In_949,In_21);
and U4116 (N_4116,In_557,In_812);
nand U4117 (N_4117,In_301,In_986);
and U4118 (N_4118,In_109,In_376);
nor U4119 (N_4119,In_856,In_694);
and U4120 (N_4120,In_651,In_304);
nor U4121 (N_4121,In_824,In_630);
nand U4122 (N_4122,In_217,In_78);
nor U4123 (N_4123,In_341,In_989);
nor U4124 (N_4124,In_102,In_200);
and U4125 (N_4125,In_417,In_53);
xnor U4126 (N_4126,In_558,In_295);
nand U4127 (N_4127,In_566,In_513);
or U4128 (N_4128,In_743,In_990);
xor U4129 (N_4129,In_219,In_182);
xor U4130 (N_4130,In_461,In_251);
or U4131 (N_4131,In_335,In_579);
nand U4132 (N_4132,In_881,In_841);
nand U4133 (N_4133,In_595,In_739);
nand U4134 (N_4134,In_906,In_552);
or U4135 (N_4135,In_219,In_433);
xor U4136 (N_4136,In_319,In_973);
nand U4137 (N_4137,In_947,In_30);
nand U4138 (N_4138,In_922,In_396);
xor U4139 (N_4139,In_536,In_263);
nand U4140 (N_4140,In_437,In_909);
nand U4141 (N_4141,In_736,In_954);
nand U4142 (N_4142,In_161,In_794);
and U4143 (N_4143,In_411,In_805);
or U4144 (N_4144,In_867,In_437);
nor U4145 (N_4145,In_885,In_598);
and U4146 (N_4146,In_398,In_959);
and U4147 (N_4147,In_927,In_511);
or U4148 (N_4148,In_658,In_248);
xnor U4149 (N_4149,In_941,In_575);
and U4150 (N_4150,In_613,In_640);
nor U4151 (N_4151,In_126,In_752);
xor U4152 (N_4152,In_605,In_328);
nor U4153 (N_4153,In_539,In_249);
and U4154 (N_4154,In_263,In_289);
nor U4155 (N_4155,In_602,In_565);
and U4156 (N_4156,In_268,In_932);
and U4157 (N_4157,In_270,In_129);
xnor U4158 (N_4158,In_908,In_140);
nand U4159 (N_4159,In_743,In_341);
xor U4160 (N_4160,In_337,In_649);
nand U4161 (N_4161,In_816,In_730);
nand U4162 (N_4162,In_997,In_264);
or U4163 (N_4163,In_73,In_554);
or U4164 (N_4164,In_197,In_408);
and U4165 (N_4165,In_79,In_766);
xnor U4166 (N_4166,In_727,In_228);
nand U4167 (N_4167,In_21,In_733);
nand U4168 (N_4168,In_150,In_708);
nand U4169 (N_4169,In_40,In_935);
or U4170 (N_4170,In_675,In_881);
and U4171 (N_4171,In_128,In_220);
or U4172 (N_4172,In_524,In_572);
nand U4173 (N_4173,In_11,In_342);
or U4174 (N_4174,In_203,In_312);
and U4175 (N_4175,In_12,In_526);
xor U4176 (N_4176,In_23,In_586);
nand U4177 (N_4177,In_367,In_524);
or U4178 (N_4178,In_713,In_895);
nand U4179 (N_4179,In_273,In_174);
xor U4180 (N_4180,In_602,In_905);
and U4181 (N_4181,In_12,In_624);
nand U4182 (N_4182,In_764,In_633);
xor U4183 (N_4183,In_267,In_298);
or U4184 (N_4184,In_841,In_568);
nand U4185 (N_4185,In_658,In_591);
xor U4186 (N_4186,In_689,In_343);
and U4187 (N_4187,In_240,In_366);
or U4188 (N_4188,In_703,In_683);
and U4189 (N_4189,In_186,In_177);
xnor U4190 (N_4190,In_392,In_55);
nor U4191 (N_4191,In_359,In_979);
xnor U4192 (N_4192,In_958,In_241);
nor U4193 (N_4193,In_631,In_763);
and U4194 (N_4194,In_781,In_248);
and U4195 (N_4195,In_119,In_93);
nor U4196 (N_4196,In_487,In_896);
and U4197 (N_4197,In_491,In_679);
nand U4198 (N_4198,In_433,In_993);
nor U4199 (N_4199,In_438,In_275);
and U4200 (N_4200,In_701,In_948);
xor U4201 (N_4201,In_375,In_340);
nor U4202 (N_4202,In_153,In_51);
or U4203 (N_4203,In_514,In_102);
or U4204 (N_4204,In_914,In_521);
or U4205 (N_4205,In_140,In_896);
nor U4206 (N_4206,In_331,In_567);
xnor U4207 (N_4207,In_851,In_608);
or U4208 (N_4208,In_741,In_958);
or U4209 (N_4209,In_999,In_154);
and U4210 (N_4210,In_104,In_679);
or U4211 (N_4211,In_715,In_740);
or U4212 (N_4212,In_131,In_628);
nand U4213 (N_4213,In_463,In_336);
or U4214 (N_4214,In_336,In_400);
or U4215 (N_4215,In_952,In_791);
or U4216 (N_4216,In_357,In_241);
xnor U4217 (N_4217,In_956,In_850);
xnor U4218 (N_4218,In_275,In_741);
or U4219 (N_4219,In_392,In_26);
nor U4220 (N_4220,In_135,In_750);
and U4221 (N_4221,In_25,In_102);
and U4222 (N_4222,In_68,In_421);
xnor U4223 (N_4223,In_653,In_909);
nor U4224 (N_4224,In_204,In_413);
xnor U4225 (N_4225,In_24,In_309);
xor U4226 (N_4226,In_688,In_391);
or U4227 (N_4227,In_206,In_185);
or U4228 (N_4228,In_144,In_83);
and U4229 (N_4229,In_955,In_533);
or U4230 (N_4230,In_396,In_672);
or U4231 (N_4231,In_6,In_487);
nand U4232 (N_4232,In_999,In_427);
and U4233 (N_4233,In_103,In_92);
and U4234 (N_4234,In_618,In_773);
nor U4235 (N_4235,In_583,In_19);
and U4236 (N_4236,In_889,In_310);
nor U4237 (N_4237,In_983,In_10);
xnor U4238 (N_4238,In_178,In_146);
nor U4239 (N_4239,In_681,In_237);
xor U4240 (N_4240,In_883,In_233);
xor U4241 (N_4241,In_616,In_304);
nand U4242 (N_4242,In_909,In_873);
and U4243 (N_4243,In_419,In_922);
nand U4244 (N_4244,In_252,In_130);
nor U4245 (N_4245,In_189,In_61);
xor U4246 (N_4246,In_563,In_477);
xor U4247 (N_4247,In_726,In_999);
xor U4248 (N_4248,In_435,In_312);
or U4249 (N_4249,In_622,In_948);
nand U4250 (N_4250,In_713,In_698);
nor U4251 (N_4251,In_371,In_496);
or U4252 (N_4252,In_189,In_406);
or U4253 (N_4253,In_654,In_479);
nor U4254 (N_4254,In_812,In_70);
nor U4255 (N_4255,In_983,In_70);
or U4256 (N_4256,In_713,In_800);
and U4257 (N_4257,In_354,In_824);
xor U4258 (N_4258,In_332,In_401);
or U4259 (N_4259,In_305,In_949);
and U4260 (N_4260,In_975,In_778);
or U4261 (N_4261,In_251,In_963);
nor U4262 (N_4262,In_672,In_887);
nor U4263 (N_4263,In_709,In_634);
nor U4264 (N_4264,In_119,In_150);
nand U4265 (N_4265,In_618,In_843);
nor U4266 (N_4266,In_941,In_636);
or U4267 (N_4267,In_909,In_539);
nand U4268 (N_4268,In_121,In_702);
xnor U4269 (N_4269,In_859,In_451);
nand U4270 (N_4270,In_364,In_585);
xnor U4271 (N_4271,In_109,In_887);
or U4272 (N_4272,In_926,In_471);
nor U4273 (N_4273,In_299,In_307);
and U4274 (N_4274,In_61,In_182);
and U4275 (N_4275,In_11,In_405);
xnor U4276 (N_4276,In_237,In_818);
or U4277 (N_4277,In_83,In_980);
xor U4278 (N_4278,In_523,In_199);
and U4279 (N_4279,In_485,In_849);
and U4280 (N_4280,In_132,In_941);
or U4281 (N_4281,In_187,In_124);
or U4282 (N_4282,In_315,In_800);
nor U4283 (N_4283,In_371,In_788);
nor U4284 (N_4284,In_840,In_27);
nor U4285 (N_4285,In_127,In_285);
xor U4286 (N_4286,In_145,In_138);
and U4287 (N_4287,In_247,In_326);
nand U4288 (N_4288,In_979,In_757);
or U4289 (N_4289,In_647,In_301);
xnor U4290 (N_4290,In_929,In_747);
nor U4291 (N_4291,In_954,In_774);
nor U4292 (N_4292,In_1,In_217);
and U4293 (N_4293,In_901,In_104);
nand U4294 (N_4294,In_259,In_370);
or U4295 (N_4295,In_122,In_466);
and U4296 (N_4296,In_359,In_869);
or U4297 (N_4297,In_304,In_990);
nor U4298 (N_4298,In_527,In_123);
xnor U4299 (N_4299,In_320,In_498);
nand U4300 (N_4300,In_413,In_767);
nand U4301 (N_4301,In_648,In_490);
nand U4302 (N_4302,In_728,In_154);
or U4303 (N_4303,In_859,In_998);
nand U4304 (N_4304,In_384,In_240);
nand U4305 (N_4305,In_396,In_897);
nand U4306 (N_4306,In_873,In_443);
and U4307 (N_4307,In_839,In_473);
or U4308 (N_4308,In_666,In_537);
and U4309 (N_4309,In_407,In_721);
xnor U4310 (N_4310,In_130,In_580);
and U4311 (N_4311,In_168,In_509);
and U4312 (N_4312,In_207,In_128);
or U4313 (N_4313,In_838,In_678);
nor U4314 (N_4314,In_908,In_337);
nand U4315 (N_4315,In_373,In_241);
xnor U4316 (N_4316,In_722,In_760);
or U4317 (N_4317,In_736,In_533);
nand U4318 (N_4318,In_177,In_255);
nand U4319 (N_4319,In_349,In_50);
or U4320 (N_4320,In_658,In_674);
nor U4321 (N_4321,In_679,In_276);
nand U4322 (N_4322,In_257,In_784);
nor U4323 (N_4323,In_265,In_792);
nand U4324 (N_4324,In_848,In_17);
and U4325 (N_4325,In_502,In_580);
or U4326 (N_4326,In_35,In_994);
nor U4327 (N_4327,In_281,In_288);
or U4328 (N_4328,In_239,In_643);
and U4329 (N_4329,In_942,In_862);
nand U4330 (N_4330,In_897,In_198);
nor U4331 (N_4331,In_700,In_419);
nor U4332 (N_4332,In_391,In_964);
or U4333 (N_4333,In_16,In_14);
nand U4334 (N_4334,In_818,In_249);
nor U4335 (N_4335,In_545,In_470);
and U4336 (N_4336,In_205,In_403);
xnor U4337 (N_4337,In_238,In_294);
and U4338 (N_4338,In_96,In_112);
and U4339 (N_4339,In_28,In_928);
or U4340 (N_4340,In_11,In_847);
nand U4341 (N_4341,In_257,In_964);
or U4342 (N_4342,In_729,In_675);
xnor U4343 (N_4343,In_936,In_629);
or U4344 (N_4344,In_563,In_131);
nor U4345 (N_4345,In_510,In_751);
nor U4346 (N_4346,In_60,In_630);
nand U4347 (N_4347,In_698,In_595);
or U4348 (N_4348,In_317,In_490);
and U4349 (N_4349,In_792,In_236);
and U4350 (N_4350,In_185,In_28);
and U4351 (N_4351,In_637,In_223);
xor U4352 (N_4352,In_256,In_583);
xor U4353 (N_4353,In_527,In_746);
nor U4354 (N_4354,In_727,In_811);
nor U4355 (N_4355,In_438,In_966);
or U4356 (N_4356,In_127,In_423);
xnor U4357 (N_4357,In_87,In_842);
xor U4358 (N_4358,In_871,In_521);
or U4359 (N_4359,In_441,In_286);
or U4360 (N_4360,In_16,In_409);
nor U4361 (N_4361,In_923,In_817);
nand U4362 (N_4362,In_197,In_223);
nand U4363 (N_4363,In_311,In_845);
nand U4364 (N_4364,In_375,In_608);
and U4365 (N_4365,In_96,In_592);
or U4366 (N_4366,In_539,In_602);
or U4367 (N_4367,In_465,In_826);
xnor U4368 (N_4368,In_950,In_118);
nand U4369 (N_4369,In_56,In_800);
xnor U4370 (N_4370,In_163,In_677);
and U4371 (N_4371,In_989,In_262);
or U4372 (N_4372,In_238,In_306);
nand U4373 (N_4373,In_51,In_516);
nor U4374 (N_4374,In_999,In_495);
or U4375 (N_4375,In_418,In_239);
or U4376 (N_4376,In_202,In_753);
nor U4377 (N_4377,In_110,In_15);
or U4378 (N_4378,In_837,In_388);
or U4379 (N_4379,In_734,In_659);
xnor U4380 (N_4380,In_260,In_604);
nor U4381 (N_4381,In_987,In_218);
or U4382 (N_4382,In_587,In_515);
xor U4383 (N_4383,In_631,In_444);
nor U4384 (N_4384,In_84,In_679);
or U4385 (N_4385,In_548,In_832);
and U4386 (N_4386,In_126,In_840);
and U4387 (N_4387,In_487,In_92);
xnor U4388 (N_4388,In_626,In_963);
nand U4389 (N_4389,In_983,In_114);
nand U4390 (N_4390,In_112,In_381);
or U4391 (N_4391,In_370,In_515);
nand U4392 (N_4392,In_34,In_50);
nand U4393 (N_4393,In_623,In_419);
xor U4394 (N_4394,In_179,In_422);
nor U4395 (N_4395,In_434,In_490);
xnor U4396 (N_4396,In_590,In_28);
or U4397 (N_4397,In_253,In_699);
and U4398 (N_4398,In_48,In_309);
or U4399 (N_4399,In_202,In_603);
nand U4400 (N_4400,In_589,In_807);
xnor U4401 (N_4401,In_538,In_19);
nor U4402 (N_4402,In_59,In_54);
and U4403 (N_4403,In_671,In_918);
xor U4404 (N_4404,In_305,In_594);
or U4405 (N_4405,In_632,In_774);
nand U4406 (N_4406,In_800,In_216);
xor U4407 (N_4407,In_581,In_522);
nand U4408 (N_4408,In_119,In_231);
nor U4409 (N_4409,In_244,In_643);
and U4410 (N_4410,In_714,In_961);
xnor U4411 (N_4411,In_331,In_368);
nand U4412 (N_4412,In_702,In_704);
xnor U4413 (N_4413,In_223,In_309);
nand U4414 (N_4414,In_944,In_236);
xnor U4415 (N_4415,In_37,In_971);
nand U4416 (N_4416,In_347,In_363);
and U4417 (N_4417,In_355,In_575);
xor U4418 (N_4418,In_667,In_50);
or U4419 (N_4419,In_156,In_652);
nand U4420 (N_4420,In_765,In_537);
and U4421 (N_4421,In_576,In_312);
xnor U4422 (N_4422,In_11,In_161);
or U4423 (N_4423,In_462,In_536);
nand U4424 (N_4424,In_63,In_35);
and U4425 (N_4425,In_93,In_532);
nor U4426 (N_4426,In_367,In_869);
or U4427 (N_4427,In_906,In_265);
or U4428 (N_4428,In_849,In_363);
nor U4429 (N_4429,In_198,In_835);
nand U4430 (N_4430,In_816,In_978);
and U4431 (N_4431,In_819,In_162);
nor U4432 (N_4432,In_287,In_512);
xnor U4433 (N_4433,In_411,In_471);
nand U4434 (N_4434,In_873,In_236);
nand U4435 (N_4435,In_335,In_692);
and U4436 (N_4436,In_828,In_689);
nor U4437 (N_4437,In_626,In_236);
xnor U4438 (N_4438,In_435,In_785);
and U4439 (N_4439,In_558,In_283);
or U4440 (N_4440,In_709,In_271);
nor U4441 (N_4441,In_621,In_657);
nor U4442 (N_4442,In_68,In_159);
nand U4443 (N_4443,In_911,In_60);
nand U4444 (N_4444,In_658,In_638);
and U4445 (N_4445,In_905,In_47);
nand U4446 (N_4446,In_822,In_224);
and U4447 (N_4447,In_972,In_352);
xnor U4448 (N_4448,In_416,In_531);
or U4449 (N_4449,In_970,In_374);
nor U4450 (N_4450,In_76,In_216);
and U4451 (N_4451,In_127,In_933);
nand U4452 (N_4452,In_740,In_606);
nand U4453 (N_4453,In_621,In_615);
xnor U4454 (N_4454,In_964,In_909);
and U4455 (N_4455,In_385,In_764);
or U4456 (N_4456,In_452,In_208);
or U4457 (N_4457,In_3,In_306);
xnor U4458 (N_4458,In_368,In_770);
and U4459 (N_4459,In_243,In_551);
nand U4460 (N_4460,In_920,In_793);
and U4461 (N_4461,In_209,In_655);
nand U4462 (N_4462,In_285,In_169);
nor U4463 (N_4463,In_612,In_281);
nor U4464 (N_4464,In_731,In_708);
or U4465 (N_4465,In_985,In_661);
nor U4466 (N_4466,In_190,In_215);
xor U4467 (N_4467,In_407,In_91);
nor U4468 (N_4468,In_8,In_170);
nor U4469 (N_4469,In_844,In_834);
and U4470 (N_4470,In_625,In_571);
nand U4471 (N_4471,In_596,In_326);
or U4472 (N_4472,In_213,In_689);
or U4473 (N_4473,In_737,In_326);
and U4474 (N_4474,In_121,In_632);
nand U4475 (N_4475,In_859,In_609);
or U4476 (N_4476,In_728,In_58);
xor U4477 (N_4477,In_54,In_896);
or U4478 (N_4478,In_615,In_637);
or U4479 (N_4479,In_567,In_398);
and U4480 (N_4480,In_174,In_804);
xnor U4481 (N_4481,In_326,In_749);
or U4482 (N_4482,In_394,In_286);
or U4483 (N_4483,In_78,In_741);
nand U4484 (N_4484,In_645,In_394);
xor U4485 (N_4485,In_217,In_91);
or U4486 (N_4486,In_699,In_334);
and U4487 (N_4487,In_896,In_437);
xor U4488 (N_4488,In_693,In_471);
nor U4489 (N_4489,In_121,In_593);
and U4490 (N_4490,In_193,In_391);
nand U4491 (N_4491,In_799,In_884);
or U4492 (N_4492,In_129,In_736);
and U4493 (N_4493,In_884,In_670);
xnor U4494 (N_4494,In_132,In_423);
xnor U4495 (N_4495,In_51,In_172);
and U4496 (N_4496,In_705,In_393);
nor U4497 (N_4497,In_378,In_874);
nor U4498 (N_4498,In_246,In_346);
and U4499 (N_4499,In_244,In_98);
and U4500 (N_4500,In_410,In_933);
xnor U4501 (N_4501,In_231,In_200);
nor U4502 (N_4502,In_91,In_108);
or U4503 (N_4503,In_727,In_350);
nor U4504 (N_4504,In_411,In_4);
and U4505 (N_4505,In_24,In_534);
nand U4506 (N_4506,In_833,In_843);
or U4507 (N_4507,In_830,In_471);
or U4508 (N_4508,In_345,In_101);
nand U4509 (N_4509,In_828,In_190);
nand U4510 (N_4510,In_810,In_443);
xnor U4511 (N_4511,In_335,In_477);
nor U4512 (N_4512,In_917,In_630);
and U4513 (N_4513,In_276,In_824);
nand U4514 (N_4514,In_936,In_217);
xnor U4515 (N_4515,In_669,In_46);
xnor U4516 (N_4516,In_765,In_762);
and U4517 (N_4517,In_728,In_396);
and U4518 (N_4518,In_721,In_545);
or U4519 (N_4519,In_160,In_920);
xor U4520 (N_4520,In_160,In_517);
xor U4521 (N_4521,In_487,In_875);
and U4522 (N_4522,In_147,In_528);
and U4523 (N_4523,In_473,In_174);
nand U4524 (N_4524,In_918,In_143);
or U4525 (N_4525,In_94,In_649);
and U4526 (N_4526,In_23,In_773);
nand U4527 (N_4527,In_817,In_976);
nor U4528 (N_4528,In_848,In_751);
nand U4529 (N_4529,In_207,In_602);
nand U4530 (N_4530,In_898,In_974);
nand U4531 (N_4531,In_548,In_741);
or U4532 (N_4532,In_942,In_619);
and U4533 (N_4533,In_211,In_927);
nand U4534 (N_4534,In_1,In_53);
or U4535 (N_4535,In_612,In_426);
and U4536 (N_4536,In_468,In_150);
or U4537 (N_4537,In_610,In_587);
nor U4538 (N_4538,In_0,In_278);
or U4539 (N_4539,In_825,In_470);
and U4540 (N_4540,In_717,In_705);
nand U4541 (N_4541,In_174,In_228);
or U4542 (N_4542,In_740,In_53);
nor U4543 (N_4543,In_205,In_771);
nor U4544 (N_4544,In_512,In_452);
and U4545 (N_4545,In_559,In_642);
nor U4546 (N_4546,In_953,In_877);
xor U4547 (N_4547,In_823,In_407);
nand U4548 (N_4548,In_181,In_667);
nor U4549 (N_4549,In_867,In_845);
nor U4550 (N_4550,In_234,In_5);
nor U4551 (N_4551,In_125,In_718);
nand U4552 (N_4552,In_507,In_319);
or U4553 (N_4553,In_422,In_99);
and U4554 (N_4554,In_214,In_660);
or U4555 (N_4555,In_100,In_156);
xnor U4556 (N_4556,In_705,In_216);
xor U4557 (N_4557,In_727,In_181);
nor U4558 (N_4558,In_830,In_673);
nor U4559 (N_4559,In_590,In_105);
and U4560 (N_4560,In_347,In_840);
or U4561 (N_4561,In_293,In_439);
and U4562 (N_4562,In_618,In_613);
and U4563 (N_4563,In_203,In_233);
xor U4564 (N_4564,In_372,In_958);
or U4565 (N_4565,In_103,In_57);
or U4566 (N_4566,In_894,In_162);
nor U4567 (N_4567,In_598,In_161);
nor U4568 (N_4568,In_920,In_957);
xnor U4569 (N_4569,In_198,In_566);
nand U4570 (N_4570,In_215,In_981);
and U4571 (N_4571,In_257,In_649);
xor U4572 (N_4572,In_245,In_815);
xnor U4573 (N_4573,In_875,In_580);
xor U4574 (N_4574,In_598,In_817);
xor U4575 (N_4575,In_234,In_212);
xor U4576 (N_4576,In_330,In_351);
xnor U4577 (N_4577,In_87,In_802);
nand U4578 (N_4578,In_63,In_680);
and U4579 (N_4579,In_442,In_75);
nand U4580 (N_4580,In_114,In_348);
xnor U4581 (N_4581,In_489,In_99);
nor U4582 (N_4582,In_119,In_254);
nor U4583 (N_4583,In_306,In_312);
nor U4584 (N_4584,In_0,In_185);
nand U4585 (N_4585,In_771,In_286);
or U4586 (N_4586,In_530,In_942);
or U4587 (N_4587,In_396,In_223);
xor U4588 (N_4588,In_384,In_230);
and U4589 (N_4589,In_651,In_461);
and U4590 (N_4590,In_968,In_416);
nor U4591 (N_4591,In_13,In_26);
or U4592 (N_4592,In_699,In_817);
or U4593 (N_4593,In_991,In_574);
and U4594 (N_4594,In_401,In_195);
and U4595 (N_4595,In_5,In_157);
nor U4596 (N_4596,In_40,In_291);
and U4597 (N_4597,In_555,In_130);
xnor U4598 (N_4598,In_111,In_422);
or U4599 (N_4599,In_431,In_317);
nand U4600 (N_4600,In_220,In_243);
nor U4601 (N_4601,In_714,In_445);
and U4602 (N_4602,In_26,In_418);
xnor U4603 (N_4603,In_617,In_819);
or U4604 (N_4604,In_997,In_736);
or U4605 (N_4605,In_661,In_172);
or U4606 (N_4606,In_469,In_394);
xnor U4607 (N_4607,In_691,In_735);
xnor U4608 (N_4608,In_609,In_774);
and U4609 (N_4609,In_319,In_281);
nand U4610 (N_4610,In_4,In_680);
and U4611 (N_4611,In_971,In_450);
and U4612 (N_4612,In_702,In_48);
nor U4613 (N_4613,In_402,In_176);
nor U4614 (N_4614,In_227,In_981);
nor U4615 (N_4615,In_489,In_510);
or U4616 (N_4616,In_547,In_916);
or U4617 (N_4617,In_794,In_786);
or U4618 (N_4618,In_672,In_92);
nand U4619 (N_4619,In_290,In_564);
and U4620 (N_4620,In_458,In_487);
and U4621 (N_4621,In_18,In_347);
nand U4622 (N_4622,In_530,In_947);
or U4623 (N_4623,In_68,In_757);
xor U4624 (N_4624,In_962,In_202);
xor U4625 (N_4625,In_750,In_802);
and U4626 (N_4626,In_578,In_839);
nand U4627 (N_4627,In_353,In_784);
and U4628 (N_4628,In_42,In_618);
nand U4629 (N_4629,In_117,In_979);
xnor U4630 (N_4630,In_927,In_256);
nor U4631 (N_4631,In_454,In_1);
nand U4632 (N_4632,In_662,In_529);
or U4633 (N_4633,In_300,In_194);
nand U4634 (N_4634,In_329,In_737);
nand U4635 (N_4635,In_757,In_650);
nor U4636 (N_4636,In_758,In_914);
nand U4637 (N_4637,In_486,In_612);
or U4638 (N_4638,In_788,In_59);
or U4639 (N_4639,In_705,In_291);
and U4640 (N_4640,In_207,In_386);
xor U4641 (N_4641,In_701,In_121);
and U4642 (N_4642,In_489,In_403);
and U4643 (N_4643,In_995,In_938);
or U4644 (N_4644,In_875,In_25);
xor U4645 (N_4645,In_287,In_580);
nand U4646 (N_4646,In_51,In_535);
nor U4647 (N_4647,In_907,In_893);
nor U4648 (N_4648,In_383,In_601);
nand U4649 (N_4649,In_619,In_54);
xor U4650 (N_4650,In_294,In_837);
xor U4651 (N_4651,In_567,In_643);
and U4652 (N_4652,In_920,In_112);
or U4653 (N_4653,In_207,In_423);
or U4654 (N_4654,In_358,In_135);
xnor U4655 (N_4655,In_299,In_412);
or U4656 (N_4656,In_425,In_795);
nand U4657 (N_4657,In_936,In_608);
xnor U4658 (N_4658,In_844,In_879);
and U4659 (N_4659,In_131,In_172);
nor U4660 (N_4660,In_4,In_170);
and U4661 (N_4661,In_500,In_590);
xnor U4662 (N_4662,In_616,In_396);
nor U4663 (N_4663,In_300,In_104);
and U4664 (N_4664,In_526,In_869);
nand U4665 (N_4665,In_106,In_368);
nand U4666 (N_4666,In_965,In_877);
xor U4667 (N_4667,In_163,In_867);
nand U4668 (N_4668,In_63,In_684);
and U4669 (N_4669,In_999,In_56);
and U4670 (N_4670,In_86,In_548);
and U4671 (N_4671,In_88,In_544);
xnor U4672 (N_4672,In_63,In_107);
nor U4673 (N_4673,In_270,In_676);
xnor U4674 (N_4674,In_236,In_606);
nand U4675 (N_4675,In_708,In_413);
nand U4676 (N_4676,In_441,In_671);
xnor U4677 (N_4677,In_545,In_845);
nand U4678 (N_4678,In_226,In_378);
xnor U4679 (N_4679,In_47,In_798);
or U4680 (N_4680,In_837,In_794);
or U4681 (N_4681,In_195,In_21);
nand U4682 (N_4682,In_166,In_507);
xnor U4683 (N_4683,In_179,In_335);
nand U4684 (N_4684,In_393,In_923);
nand U4685 (N_4685,In_895,In_845);
nand U4686 (N_4686,In_748,In_645);
nor U4687 (N_4687,In_777,In_372);
or U4688 (N_4688,In_217,In_177);
or U4689 (N_4689,In_117,In_455);
or U4690 (N_4690,In_495,In_192);
and U4691 (N_4691,In_931,In_862);
and U4692 (N_4692,In_229,In_597);
xnor U4693 (N_4693,In_953,In_709);
nand U4694 (N_4694,In_650,In_807);
xor U4695 (N_4695,In_608,In_954);
nand U4696 (N_4696,In_731,In_365);
nand U4697 (N_4697,In_568,In_687);
xnor U4698 (N_4698,In_810,In_704);
xor U4699 (N_4699,In_222,In_202);
nor U4700 (N_4700,In_58,In_759);
and U4701 (N_4701,In_973,In_222);
nand U4702 (N_4702,In_77,In_192);
nand U4703 (N_4703,In_874,In_160);
nor U4704 (N_4704,In_419,In_737);
xnor U4705 (N_4705,In_717,In_982);
and U4706 (N_4706,In_468,In_263);
nand U4707 (N_4707,In_748,In_18);
xnor U4708 (N_4708,In_358,In_582);
or U4709 (N_4709,In_987,In_206);
and U4710 (N_4710,In_801,In_67);
and U4711 (N_4711,In_104,In_426);
or U4712 (N_4712,In_118,In_668);
xor U4713 (N_4713,In_334,In_380);
and U4714 (N_4714,In_884,In_632);
xnor U4715 (N_4715,In_206,In_803);
nor U4716 (N_4716,In_94,In_715);
nor U4717 (N_4717,In_581,In_41);
or U4718 (N_4718,In_839,In_368);
or U4719 (N_4719,In_92,In_360);
nand U4720 (N_4720,In_380,In_847);
or U4721 (N_4721,In_957,In_353);
and U4722 (N_4722,In_140,In_208);
and U4723 (N_4723,In_664,In_785);
nand U4724 (N_4724,In_262,In_558);
and U4725 (N_4725,In_850,In_140);
xor U4726 (N_4726,In_39,In_736);
nor U4727 (N_4727,In_583,In_928);
nor U4728 (N_4728,In_985,In_844);
or U4729 (N_4729,In_360,In_518);
nand U4730 (N_4730,In_194,In_28);
or U4731 (N_4731,In_327,In_804);
xnor U4732 (N_4732,In_597,In_510);
nor U4733 (N_4733,In_608,In_515);
nor U4734 (N_4734,In_321,In_735);
and U4735 (N_4735,In_430,In_369);
or U4736 (N_4736,In_489,In_834);
xnor U4737 (N_4737,In_510,In_720);
xnor U4738 (N_4738,In_511,In_946);
and U4739 (N_4739,In_574,In_971);
xor U4740 (N_4740,In_408,In_960);
nor U4741 (N_4741,In_257,In_117);
and U4742 (N_4742,In_595,In_954);
or U4743 (N_4743,In_227,In_923);
nor U4744 (N_4744,In_348,In_291);
xnor U4745 (N_4745,In_331,In_805);
and U4746 (N_4746,In_372,In_256);
nand U4747 (N_4747,In_570,In_783);
nand U4748 (N_4748,In_678,In_485);
nand U4749 (N_4749,In_949,In_797);
nor U4750 (N_4750,In_949,In_454);
nor U4751 (N_4751,In_549,In_354);
nand U4752 (N_4752,In_732,In_740);
nand U4753 (N_4753,In_502,In_352);
and U4754 (N_4754,In_128,In_214);
xor U4755 (N_4755,In_151,In_382);
or U4756 (N_4756,In_649,In_122);
xnor U4757 (N_4757,In_52,In_513);
xor U4758 (N_4758,In_657,In_965);
and U4759 (N_4759,In_119,In_865);
or U4760 (N_4760,In_662,In_430);
nor U4761 (N_4761,In_567,In_191);
xnor U4762 (N_4762,In_154,In_279);
xor U4763 (N_4763,In_119,In_576);
xnor U4764 (N_4764,In_666,In_899);
nor U4765 (N_4765,In_33,In_490);
xnor U4766 (N_4766,In_138,In_35);
and U4767 (N_4767,In_306,In_982);
nand U4768 (N_4768,In_592,In_418);
or U4769 (N_4769,In_131,In_797);
and U4770 (N_4770,In_729,In_585);
nor U4771 (N_4771,In_85,In_786);
and U4772 (N_4772,In_691,In_41);
nand U4773 (N_4773,In_465,In_173);
and U4774 (N_4774,In_751,In_34);
or U4775 (N_4775,In_128,In_163);
or U4776 (N_4776,In_576,In_716);
nor U4777 (N_4777,In_793,In_598);
nor U4778 (N_4778,In_540,In_219);
xor U4779 (N_4779,In_710,In_937);
and U4780 (N_4780,In_708,In_987);
nor U4781 (N_4781,In_852,In_211);
and U4782 (N_4782,In_1,In_536);
xor U4783 (N_4783,In_550,In_455);
or U4784 (N_4784,In_857,In_564);
nor U4785 (N_4785,In_45,In_974);
and U4786 (N_4786,In_737,In_114);
nor U4787 (N_4787,In_591,In_228);
nand U4788 (N_4788,In_453,In_38);
nor U4789 (N_4789,In_599,In_350);
nor U4790 (N_4790,In_883,In_885);
nand U4791 (N_4791,In_962,In_618);
and U4792 (N_4792,In_889,In_991);
xnor U4793 (N_4793,In_957,In_799);
nand U4794 (N_4794,In_217,In_21);
xnor U4795 (N_4795,In_236,In_643);
nor U4796 (N_4796,In_439,In_585);
or U4797 (N_4797,In_669,In_640);
nand U4798 (N_4798,In_272,In_485);
xor U4799 (N_4799,In_56,In_524);
nand U4800 (N_4800,In_960,In_606);
or U4801 (N_4801,In_658,In_536);
xnor U4802 (N_4802,In_5,In_287);
xor U4803 (N_4803,In_27,In_792);
and U4804 (N_4804,In_672,In_175);
or U4805 (N_4805,In_499,In_945);
nor U4806 (N_4806,In_844,In_230);
nor U4807 (N_4807,In_179,In_464);
nand U4808 (N_4808,In_106,In_963);
and U4809 (N_4809,In_86,In_606);
nor U4810 (N_4810,In_480,In_167);
or U4811 (N_4811,In_388,In_61);
xor U4812 (N_4812,In_811,In_669);
and U4813 (N_4813,In_328,In_756);
or U4814 (N_4814,In_515,In_314);
xnor U4815 (N_4815,In_933,In_309);
xnor U4816 (N_4816,In_282,In_279);
nor U4817 (N_4817,In_262,In_195);
nand U4818 (N_4818,In_744,In_308);
or U4819 (N_4819,In_209,In_11);
and U4820 (N_4820,In_778,In_928);
xor U4821 (N_4821,In_819,In_898);
nor U4822 (N_4822,In_705,In_703);
nand U4823 (N_4823,In_124,In_33);
and U4824 (N_4824,In_963,In_87);
nand U4825 (N_4825,In_842,In_63);
or U4826 (N_4826,In_811,In_495);
nor U4827 (N_4827,In_765,In_323);
xor U4828 (N_4828,In_762,In_968);
nand U4829 (N_4829,In_756,In_155);
nand U4830 (N_4830,In_451,In_204);
nand U4831 (N_4831,In_833,In_535);
or U4832 (N_4832,In_180,In_279);
nor U4833 (N_4833,In_671,In_110);
and U4834 (N_4834,In_650,In_74);
or U4835 (N_4835,In_391,In_601);
nand U4836 (N_4836,In_128,In_413);
nand U4837 (N_4837,In_894,In_135);
nor U4838 (N_4838,In_166,In_452);
nand U4839 (N_4839,In_2,In_672);
and U4840 (N_4840,In_592,In_314);
nand U4841 (N_4841,In_730,In_39);
nand U4842 (N_4842,In_103,In_331);
or U4843 (N_4843,In_652,In_295);
xnor U4844 (N_4844,In_763,In_618);
or U4845 (N_4845,In_269,In_904);
nor U4846 (N_4846,In_546,In_610);
xnor U4847 (N_4847,In_661,In_369);
and U4848 (N_4848,In_839,In_122);
or U4849 (N_4849,In_400,In_171);
or U4850 (N_4850,In_386,In_805);
nor U4851 (N_4851,In_192,In_786);
nand U4852 (N_4852,In_502,In_328);
and U4853 (N_4853,In_12,In_41);
or U4854 (N_4854,In_548,In_788);
nand U4855 (N_4855,In_348,In_190);
xnor U4856 (N_4856,In_235,In_735);
nand U4857 (N_4857,In_427,In_100);
or U4858 (N_4858,In_611,In_393);
nand U4859 (N_4859,In_78,In_345);
xor U4860 (N_4860,In_581,In_984);
xnor U4861 (N_4861,In_172,In_246);
xnor U4862 (N_4862,In_185,In_215);
xor U4863 (N_4863,In_402,In_31);
xor U4864 (N_4864,In_757,In_106);
or U4865 (N_4865,In_153,In_940);
or U4866 (N_4866,In_73,In_293);
and U4867 (N_4867,In_778,In_42);
nand U4868 (N_4868,In_377,In_939);
and U4869 (N_4869,In_74,In_439);
xor U4870 (N_4870,In_393,In_823);
and U4871 (N_4871,In_69,In_601);
or U4872 (N_4872,In_519,In_803);
and U4873 (N_4873,In_741,In_992);
nor U4874 (N_4874,In_656,In_353);
nor U4875 (N_4875,In_847,In_132);
and U4876 (N_4876,In_260,In_713);
and U4877 (N_4877,In_876,In_534);
and U4878 (N_4878,In_538,In_349);
or U4879 (N_4879,In_125,In_79);
or U4880 (N_4880,In_956,In_140);
xnor U4881 (N_4881,In_899,In_913);
and U4882 (N_4882,In_412,In_641);
or U4883 (N_4883,In_91,In_678);
nor U4884 (N_4884,In_990,In_525);
or U4885 (N_4885,In_59,In_696);
or U4886 (N_4886,In_267,In_299);
and U4887 (N_4887,In_202,In_578);
nand U4888 (N_4888,In_565,In_771);
nor U4889 (N_4889,In_692,In_372);
and U4890 (N_4890,In_267,In_505);
and U4891 (N_4891,In_631,In_761);
nor U4892 (N_4892,In_675,In_481);
and U4893 (N_4893,In_3,In_626);
or U4894 (N_4894,In_91,In_65);
and U4895 (N_4895,In_645,In_744);
nand U4896 (N_4896,In_340,In_368);
nor U4897 (N_4897,In_508,In_178);
xor U4898 (N_4898,In_108,In_810);
xnor U4899 (N_4899,In_224,In_250);
xor U4900 (N_4900,In_837,In_969);
or U4901 (N_4901,In_743,In_947);
xnor U4902 (N_4902,In_321,In_58);
or U4903 (N_4903,In_779,In_5);
nand U4904 (N_4904,In_23,In_862);
and U4905 (N_4905,In_109,In_401);
xnor U4906 (N_4906,In_906,In_995);
xnor U4907 (N_4907,In_324,In_43);
xnor U4908 (N_4908,In_74,In_477);
and U4909 (N_4909,In_838,In_469);
and U4910 (N_4910,In_139,In_719);
or U4911 (N_4911,In_313,In_415);
and U4912 (N_4912,In_505,In_289);
nor U4913 (N_4913,In_665,In_688);
nand U4914 (N_4914,In_351,In_252);
or U4915 (N_4915,In_514,In_4);
and U4916 (N_4916,In_558,In_931);
xnor U4917 (N_4917,In_389,In_351);
nor U4918 (N_4918,In_768,In_885);
and U4919 (N_4919,In_305,In_916);
and U4920 (N_4920,In_800,In_462);
or U4921 (N_4921,In_235,In_809);
or U4922 (N_4922,In_540,In_50);
nand U4923 (N_4923,In_216,In_301);
nand U4924 (N_4924,In_489,In_172);
nor U4925 (N_4925,In_225,In_602);
xnor U4926 (N_4926,In_5,In_846);
nand U4927 (N_4927,In_207,In_766);
nor U4928 (N_4928,In_353,In_917);
nand U4929 (N_4929,In_12,In_336);
nor U4930 (N_4930,In_416,In_579);
and U4931 (N_4931,In_670,In_140);
nand U4932 (N_4932,In_878,In_482);
nand U4933 (N_4933,In_877,In_125);
or U4934 (N_4934,In_333,In_530);
nor U4935 (N_4935,In_825,In_288);
or U4936 (N_4936,In_223,In_839);
or U4937 (N_4937,In_107,In_527);
nand U4938 (N_4938,In_513,In_45);
and U4939 (N_4939,In_797,In_725);
nor U4940 (N_4940,In_797,In_469);
or U4941 (N_4941,In_876,In_649);
or U4942 (N_4942,In_598,In_490);
nor U4943 (N_4943,In_7,In_370);
xnor U4944 (N_4944,In_974,In_755);
or U4945 (N_4945,In_652,In_314);
nor U4946 (N_4946,In_201,In_496);
and U4947 (N_4947,In_702,In_522);
and U4948 (N_4948,In_120,In_770);
nand U4949 (N_4949,In_889,In_908);
nand U4950 (N_4950,In_947,In_807);
nand U4951 (N_4951,In_598,In_284);
nor U4952 (N_4952,In_278,In_88);
nor U4953 (N_4953,In_586,In_25);
nand U4954 (N_4954,In_704,In_15);
nand U4955 (N_4955,In_201,In_780);
xor U4956 (N_4956,In_44,In_776);
nor U4957 (N_4957,In_298,In_857);
xnor U4958 (N_4958,In_674,In_870);
nor U4959 (N_4959,In_388,In_387);
and U4960 (N_4960,In_718,In_330);
nand U4961 (N_4961,In_739,In_937);
and U4962 (N_4962,In_848,In_309);
nand U4963 (N_4963,In_406,In_202);
and U4964 (N_4964,In_276,In_610);
and U4965 (N_4965,In_283,In_104);
nor U4966 (N_4966,In_775,In_93);
nor U4967 (N_4967,In_586,In_135);
and U4968 (N_4968,In_699,In_14);
nand U4969 (N_4969,In_268,In_57);
or U4970 (N_4970,In_942,In_600);
and U4971 (N_4971,In_734,In_165);
xor U4972 (N_4972,In_996,In_800);
nand U4973 (N_4973,In_673,In_851);
nand U4974 (N_4974,In_642,In_358);
nor U4975 (N_4975,In_65,In_770);
nor U4976 (N_4976,In_384,In_423);
nor U4977 (N_4977,In_461,In_192);
xnor U4978 (N_4978,In_349,In_925);
and U4979 (N_4979,In_336,In_691);
nor U4980 (N_4980,In_459,In_919);
nand U4981 (N_4981,In_803,In_841);
and U4982 (N_4982,In_607,In_611);
nand U4983 (N_4983,In_91,In_901);
nand U4984 (N_4984,In_698,In_596);
nor U4985 (N_4985,In_50,In_638);
and U4986 (N_4986,In_999,In_364);
nand U4987 (N_4987,In_424,In_517);
and U4988 (N_4988,In_991,In_746);
nand U4989 (N_4989,In_326,In_729);
nor U4990 (N_4990,In_685,In_737);
nor U4991 (N_4991,In_986,In_509);
and U4992 (N_4992,In_999,In_836);
and U4993 (N_4993,In_957,In_110);
nor U4994 (N_4994,In_638,In_643);
nand U4995 (N_4995,In_306,In_101);
nand U4996 (N_4996,In_103,In_605);
nand U4997 (N_4997,In_463,In_379);
nand U4998 (N_4998,In_777,In_665);
nor U4999 (N_4999,In_619,In_829);
nand U5000 (N_5000,N_4320,N_2511);
xor U5001 (N_5001,N_1586,N_233);
nor U5002 (N_5002,N_4077,N_4983);
or U5003 (N_5003,N_2611,N_1181);
xnor U5004 (N_5004,N_1458,N_2161);
or U5005 (N_5005,N_4907,N_1476);
or U5006 (N_5006,N_4158,N_495);
and U5007 (N_5007,N_2565,N_2683);
nand U5008 (N_5008,N_4156,N_4899);
and U5009 (N_5009,N_129,N_4345);
nand U5010 (N_5010,N_2996,N_447);
nand U5011 (N_5011,N_4238,N_2489);
or U5012 (N_5012,N_1621,N_2931);
or U5013 (N_5013,N_2838,N_382);
nor U5014 (N_5014,N_2098,N_1987);
nor U5015 (N_5015,N_2004,N_4691);
nor U5016 (N_5016,N_836,N_1677);
xnor U5017 (N_5017,N_2736,N_1413);
or U5018 (N_5018,N_3140,N_2227);
and U5019 (N_5019,N_4117,N_1789);
and U5020 (N_5020,N_3828,N_1409);
or U5021 (N_5021,N_4218,N_1399);
nor U5022 (N_5022,N_2497,N_2969);
and U5023 (N_5023,N_973,N_2705);
and U5024 (N_5024,N_1917,N_2492);
and U5025 (N_5025,N_4129,N_4217);
or U5026 (N_5026,N_4414,N_328);
and U5027 (N_5027,N_907,N_1781);
nor U5028 (N_5028,N_3535,N_3826);
or U5029 (N_5029,N_192,N_372);
and U5030 (N_5030,N_3138,N_4222);
or U5031 (N_5031,N_2772,N_1152);
and U5032 (N_5032,N_3960,N_865);
and U5033 (N_5033,N_3029,N_3507);
xor U5034 (N_5034,N_2314,N_3266);
and U5035 (N_5035,N_3817,N_2695);
nand U5036 (N_5036,N_3556,N_2206);
xor U5037 (N_5037,N_3359,N_648);
and U5038 (N_5038,N_1473,N_3179);
and U5039 (N_5039,N_4670,N_1821);
and U5040 (N_5040,N_755,N_736);
nand U5041 (N_5041,N_1211,N_1900);
or U5042 (N_5042,N_433,N_1784);
or U5043 (N_5043,N_2093,N_4245);
nor U5044 (N_5044,N_3791,N_4493);
nand U5045 (N_5045,N_2403,N_831);
or U5046 (N_5046,N_339,N_3715);
and U5047 (N_5047,N_1297,N_4554);
xor U5048 (N_5048,N_4177,N_4745);
xnor U5049 (N_5049,N_2071,N_3422);
nand U5050 (N_5050,N_4364,N_4005);
nand U5051 (N_5051,N_843,N_1353);
xor U5052 (N_5052,N_1188,N_3753);
or U5053 (N_5053,N_3433,N_2443);
nand U5054 (N_5054,N_596,N_1623);
xnor U5055 (N_5055,N_1847,N_987);
nand U5056 (N_5056,N_1991,N_2711);
or U5057 (N_5057,N_2134,N_717);
and U5058 (N_5058,N_4172,N_2876);
nand U5059 (N_5059,N_1651,N_2635);
nor U5060 (N_5060,N_4694,N_370);
or U5061 (N_5061,N_2391,N_3161);
xnor U5062 (N_5062,N_1788,N_2961);
xor U5063 (N_5063,N_1942,N_4291);
or U5064 (N_5064,N_4531,N_4242);
nand U5065 (N_5065,N_2785,N_4311);
or U5066 (N_5066,N_3302,N_799);
nand U5067 (N_5067,N_4638,N_4254);
xnor U5068 (N_5068,N_1906,N_36);
or U5069 (N_5069,N_3132,N_4346);
nor U5070 (N_5070,N_4572,N_4332);
nand U5071 (N_5071,N_475,N_179);
nor U5072 (N_5072,N_4934,N_2681);
and U5073 (N_5073,N_2327,N_4995);
xor U5074 (N_5074,N_1134,N_3597);
xor U5075 (N_5075,N_3989,N_4279);
nor U5076 (N_5076,N_1713,N_3530);
and U5077 (N_5077,N_1149,N_1450);
and U5078 (N_5078,N_636,N_943);
nor U5079 (N_5079,N_884,N_2294);
or U5080 (N_5080,N_2908,N_4573);
xor U5081 (N_5081,N_441,N_1962);
nand U5082 (N_5082,N_1873,N_692);
and U5083 (N_5083,N_1195,N_3965);
or U5084 (N_5084,N_3122,N_2460);
nand U5085 (N_5085,N_307,N_2075);
xnor U5086 (N_5086,N_3014,N_3956);
nand U5087 (N_5087,N_3457,N_1384);
nand U5088 (N_5088,N_4943,N_2);
or U5089 (N_5089,N_3400,N_2377);
xor U5090 (N_5090,N_1637,N_1056);
nand U5091 (N_5091,N_1835,N_3631);
and U5092 (N_5092,N_4268,N_4593);
nand U5093 (N_5093,N_1456,N_891);
and U5094 (N_5094,N_2439,N_1461);
nor U5095 (N_5095,N_1357,N_2648);
nor U5096 (N_5096,N_4062,N_2257);
or U5097 (N_5097,N_2577,N_2551);
nor U5098 (N_5098,N_1554,N_3235);
or U5099 (N_5099,N_440,N_1051);
or U5100 (N_5100,N_2018,N_2633);
nor U5101 (N_5101,N_4930,N_2625);
nor U5102 (N_5102,N_694,N_1485);
and U5103 (N_5103,N_4210,N_3057);
nor U5104 (N_5104,N_1958,N_4180);
nand U5105 (N_5105,N_2643,N_3314);
nor U5106 (N_5106,N_1592,N_2433);
nor U5107 (N_5107,N_2038,N_404);
nor U5108 (N_5108,N_3026,N_4952);
nor U5109 (N_5109,N_4626,N_1338);
or U5110 (N_5110,N_3009,N_3573);
nor U5111 (N_5111,N_641,N_199);
xnor U5112 (N_5112,N_3567,N_2613);
xor U5113 (N_5113,N_3577,N_4483);
or U5114 (N_5114,N_2766,N_4266);
nand U5115 (N_5115,N_3024,N_3875);
nand U5116 (N_5116,N_29,N_1408);
nor U5117 (N_5117,N_376,N_3462);
xor U5118 (N_5118,N_1214,N_1633);
and U5119 (N_5119,N_1773,N_1909);
nand U5120 (N_5120,N_640,N_163);
and U5121 (N_5121,N_2500,N_3624);
or U5122 (N_5122,N_1032,N_4886);
and U5123 (N_5123,N_128,N_3155);
and U5124 (N_5124,N_2234,N_3861);
nand U5125 (N_5125,N_4825,N_4119);
nor U5126 (N_5126,N_2941,N_945);
nand U5127 (N_5127,N_3156,N_1916);
nor U5128 (N_5128,N_750,N_4806);
nand U5129 (N_5129,N_2560,N_2680);
nand U5130 (N_5130,N_1889,N_558);
nor U5131 (N_5131,N_1972,N_2097);
or U5132 (N_5132,N_1982,N_3969);
nor U5133 (N_5133,N_1508,N_3690);
nor U5134 (N_5134,N_487,N_2900);
or U5135 (N_5135,N_4824,N_40);
and U5136 (N_5136,N_4153,N_2179);
nand U5137 (N_5137,N_291,N_2122);
nand U5138 (N_5138,N_1698,N_4956);
nand U5139 (N_5139,N_1726,N_2849);
and U5140 (N_5140,N_2697,N_707);
nor U5141 (N_5141,N_3851,N_3315);
nand U5142 (N_5142,N_2444,N_71);
nand U5143 (N_5143,N_2786,N_539);
or U5144 (N_5144,N_4081,N_2325);
xor U5145 (N_5145,N_691,N_1884);
nor U5146 (N_5146,N_1128,N_3526);
nor U5147 (N_5147,N_4082,N_4797);
nor U5148 (N_5148,N_1778,N_4073);
and U5149 (N_5149,N_1915,N_3193);
and U5150 (N_5150,N_2916,N_2525);
xnor U5151 (N_5151,N_3761,N_20);
xor U5152 (N_5152,N_4911,N_643);
or U5153 (N_5153,N_48,N_1209);
nand U5154 (N_5154,N_2707,N_1660);
or U5155 (N_5155,N_967,N_3815);
or U5156 (N_5156,N_4220,N_4025);
or U5157 (N_5157,N_4067,N_3525);
nor U5158 (N_5158,N_2652,N_826);
and U5159 (N_5159,N_503,N_4722);
and U5160 (N_5160,N_269,N_3395);
nor U5161 (N_5161,N_2535,N_480);
or U5162 (N_5162,N_2152,N_2569);
and U5163 (N_5163,N_602,N_3948);
and U5164 (N_5164,N_767,N_1393);
nor U5165 (N_5165,N_3063,N_258);
or U5166 (N_5166,N_4046,N_1995);
xnor U5167 (N_5167,N_3221,N_3819);
nand U5168 (N_5168,N_1268,N_4852);
and U5169 (N_5169,N_3432,N_2504);
nand U5170 (N_5170,N_1392,N_2163);
xnor U5171 (N_5171,N_4955,N_900);
nor U5172 (N_5172,N_3354,N_895);
nand U5173 (N_5173,N_4361,N_4446);
or U5174 (N_5174,N_2642,N_2666);
and U5175 (N_5175,N_3677,N_1434);
nand U5176 (N_5176,N_1684,N_1863);
and U5177 (N_5177,N_1832,N_2870);
nand U5178 (N_5178,N_1599,N_2480);
xor U5179 (N_5179,N_3284,N_2675);
nand U5180 (N_5180,N_2236,N_1208);
nand U5181 (N_5181,N_397,N_3553);
or U5182 (N_5182,N_2452,N_1736);
xnor U5183 (N_5183,N_4494,N_1729);
nand U5184 (N_5184,N_2396,N_4602);
and U5185 (N_5185,N_4862,N_458);
nor U5186 (N_5186,N_612,N_1078);
nor U5187 (N_5187,N_120,N_2842);
xor U5188 (N_5188,N_2253,N_4668);
or U5189 (N_5189,N_1182,N_1823);
and U5190 (N_5190,N_4275,N_2235);
nor U5191 (N_5191,N_570,N_1335);
nand U5192 (N_5192,N_52,N_1272);
and U5193 (N_5193,N_3520,N_1624);
nand U5194 (N_5194,N_74,N_3166);
xor U5195 (N_5195,N_578,N_1381);
nand U5196 (N_5196,N_1363,N_2077);
nor U5197 (N_5197,N_561,N_3532);
and U5198 (N_5198,N_1530,N_3318);
xnor U5199 (N_5199,N_4566,N_1154);
nor U5200 (N_5200,N_243,N_2266);
or U5201 (N_5201,N_3145,N_2508);
and U5202 (N_5202,N_91,N_2717);
or U5203 (N_5203,N_3726,N_2388);
nor U5204 (N_5204,N_4505,N_3979);
nor U5205 (N_5205,N_3511,N_2486);
xnor U5206 (N_5206,N_103,N_2171);
xor U5207 (N_5207,N_2986,N_4561);
nand U5208 (N_5208,N_1721,N_716);
and U5209 (N_5209,N_13,N_4834);
and U5210 (N_5210,N_183,N_2751);
and U5211 (N_5211,N_2410,N_4054);
nor U5212 (N_5212,N_1148,N_2364);
nand U5213 (N_5213,N_231,N_572);
or U5214 (N_5214,N_2767,N_2108);
nand U5215 (N_5215,N_4810,N_2856);
nand U5216 (N_5216,N_2954,N_1250);
or U5217 (N_5217,N_1885,N_2076);
nand U5218 (N_5218,N_2885,N_4926);
nor U5219 (N_5219,N_1864,N_4385);
nand U5220 (N_5220,N_950,N_2774);
nor U5221 (N_5221,N_4695,N_1059);
or U5222 (N_5222,N_3737,N_2868);
or U5223 (N_5223,N_1442,N_340);
nand U5224 (N_5224,N_4041,N_1316);
xor U5225 (N_5225,N_4632,N_400);
and U5226 (N_5226,N_3353,N_881);
nor U5227 (N_5227,N_3886,N_3419);
and U5228 (N_5228,N_1914,N_1750);
and U5229 (N_5229,N_4753,N_1119);
xor U5230 (N_5230,N_3574,N_76);
xor U5231 (N_5231,N_2835,N_19);
nor U5232 (N_5232,N_2553,N_3922);
or U5233 (N_5233,N_421,N_1082);
or U5234 (N_5234,N_903,N_2115);
nor U5235 (N_5235,N_4265,N_3191);
nor U5236 (N_5236,N_412,N_1463);
xor U5237 (N_5237,N_980,N_3021);
xor U5238 (N_5238,N_3152,N_4271);
xor U5239 (N_5239,N_2998,N_3163);
or U5240 (N_5240,N_537,N_361);
nand U5241 (N_5241,N_3608,N_952);
nor U5242 (N_5242,N_3966,N_2730);
nor U5243 (N_5243,N_4498,N_1678);
and U5244 (N_5244,N_3583,N_4109);
and U5245 (N_5245,N_3504,N_4288);
nor U5246 (N_5246,N_1039,N_1243);
xnor U5247 (N_5247,N_941,N_1782);
and U5248 (N_5248,N_2562,N_1327);
nor U5249 (N_5249,N_323,N_968);
and U5250 (N_5250,N_2753,N_657);
xor U5251 (N_5251,N_1030,N_478);
and U5252 (N_5252,N_3903,N_416);
or U5253 (N_5253,N_4149,N_921);
nand U5254 (N_5254,N_4200,N_301);
nand U5255 (N_5255,N_655,N_2459);
nand U5256 (N_5256,N_1371,N_3406);
nand U5257 (N_5257,N_186,N_4380);
nand U5258 (N_5258,N_3236,N_3897);
and U5259 (N_5259,N_1169,N_3928);
xnor U5260 (N_5260,N_4251,N_1764);
and U5261 (N_5261,N_2321,N_3135);
or U5262 (N_5262,N_2241,N_3131);
and U5263 (N_5263,N_3371,N_2369);
or U5264 (N_5264,N_852,N_3591);
or U5265 (N_5265,N_1761,N_2863);
nand U5266 (N_5266,N_3151,N_4140);
or U5267 (N_5267,N_3653,N_4545);
xnor U5268 (N_5268,N_1076,N_4103);
and U5269 (N_5269,N_3463,N_4391);
nand U5270 (N_5270,N_4548,N_4004);
and U5271 (N_5271,N_2043,N_2796);
nand U5272 (N_5272,N_2541,N_1616);
nor U5273 (N_5273,N_3051,N_2703);
xnor U5274 (N_5274,N_1215,N_4713);
and U5275 (N_5275,N_4307,N_3141);
nand U5276 (N_5276,N_2476,N_4428);
nand U5277 (N_5277,N_3823,N_234);
nor U5278 (N_5278,N_1440,N_402);
nand U5279 (N_5279,N_2570,N_4124);
nand U5280 (N_5280,N_4106,N_4927);
xnor U5281 (N_5281,N_4522,N_4565);
and U5282 (N_5282,N_3027,N_345);
and U5283 (N_5283,N_2877,N_4305);
nand U5284 (N_5284,N_3083,N_352);
and U5285 (N_5285,N_4725,N_2977);
nor U5286 (N_5286,N_113,N_1439);
nand U5287 (N_5287,N_2380,N_4151);
nand U5288 (N_5288,N_2336,N_2923);
and U5289 (N_5289,N_1446,N_2081);
and U5290 (N_5290,N_2805,N_3249);
or U5291 (N_5291,N_2907,N_1412);
nor U5292 (N_5292,N_310,N_1976);
nor U5293 (N_5293,N_3127,N_2381);
and U5294 (N_5294,N_2278,N_2400);
nor U5295 (N_5295,N_2568,N_2329);
nand U5296 (N_5296,N_204,N_971);
and U5297 (N_5297,N_3539,N_1825);
or U5298 (N_5298,N_357,N_1480);
and U5299 (N_5299,N_3290,N_835);
nor U5300 (N_5300,N_4032,N_418);
and U5301 (N_5301,N_3985,N_2563);
nand U5302 (N_5302,N_1610,N_4370);
xnor U5303 (N_5303,N_4030,N_1737);
nor U5304 (N_5304,N_2139,N_3037);
xnor U5305 (N_5305,N_1601,N_1718);
nand U5306 (N_5306,N_4134,N_442);
xor U5307 (N_5307,N_4343,N_333);
and U5308 (N_5308,N_4748,N_4451);
nor U5309 (N_5309,N_2376,N_955);
nor U5310 (N_5310,N_3736,N_4823);
nor U5311 (N_5311,N_1164,N_3208);
or U5312 (N_5312,N_4113,N_2337);
nand U5313 (N_5313,N_2123,N_781);
xor U5314 (N_5314,N_171,N_1303);
nand U5315 (N_5315,N_4513,N_3622);
and U5316 (N_5316,N_2888,N_894);
nand U5317 (N_5317,N_1000,N_689);
xor U5318 (N_5318,N_2995,N_2890);
or U5319 (N_5319,N_4201,N_346);
xor U5320 (N_5320,N_697,N_4272);
xor U5321 (N_5321,N_2769,N_906);
nor U5322 (N_5322,N_4604,N_2290);
nor U5323 (N_5323,N_3376,N_431);
and U5324 (N_5324,N_3411,N_735);
nor U5325 (N_5325,N_1329,N_2297);
or U5326 (N_5326,N_896,N_4707);
nor U5327 (N_5327,N_4719,N_4252);
nand U5328 (N_5328,N_94,N_518);
xor U5329 (N_5329,N_4693,N_2373);
or U5330 (N_5330,N_381,N_460);
or U5331 (N_5331,N_658,N_947);
or U5332 (N_5332,N_2678,N_4453);
xnor U5333 (N_5333,N_1288,N_2646);
or U5334 (N_5334,N_2917,N_2946);
xnor U5335 (N_5335,N_801,N_564);
xnor U5336 (N_5336,N_1562,N_2526);
nor U5337 (N_5337,N_4019,N_613);
and U5338 (N_5338,N_3987,N_1204);
nor U5339 (N_5339,N_1100,N_2318);
nand U5340 (N_5340,N_4649,N_3170);
xor U5341 (N_5341,N_2001,N_4068);
nor U5342 (N_5342,N_4469,N_1820);
nand U5343 (N_5343,N_4102,N_4865);
nand U5344 (N_5344,N_4987,N_4317);
or U5345 (N_5345,N_3202,N_146);
nor U5346 (N_5346,N_3201,N_4162);
nand U5347 (N_5347,N_321,N_3118);
nor U5348 (N_5348,N_58,N_3261);
nor U5349 (N_5349,N_4809,N_2363);
nand U5350 (N_5350,N_512,N_4860);
or U5351 (N_5351,N_4192,N_4904);
xor U5352 (N_5352,N_4829,N_1258);
nor U5353 (N_5353,N_814,N_2100);
and U5354 (N_5354,N_4142,N_2467);
and U5355 (N_5355,N_2855,N_1509);
and U5356 (N_5356,N_4518,N_2319);
nor U5357 (N_5357,N_4209,N_1053);
and U5358 (N_5358,N_805,N_4440);
and U5359 (N_5359,N_3452,N_3540);
or U5360 (N_5360,N_2105,N_1580);
xor U5361 (N_5361,N_3824,N_4061);
and U5362 (N_5362,N_4646,N_1373);
nor U5363 (N_5363,N_1519,N_848);
nand U5364 (N_5364,N_1992,N_545);
xor U5365 (N_5365,N_318,N_3307);
nor U5366 (N_5366,N_1939,N_10);
or U5367 (N_5367,N_700,N_1213);
nand U5368 (N_5368,N_4620,N_1938);
and U5369 (N_5369,N_4056,N_3555);
and U5370 (N_5370,N_1342,N_4340);
nor U5371 (N_5371,N_549,N_2713);
or U5372 (N_5372,N_2824,N_229);
and U5373 (N_5373,N_1683,N_723);
xor U5374 (N_5374,N_4957,N_872);
nand U5375 (N_5375,N_1499,N_1414);
xor U5376 (N_5376,N_294,N_514);
nor U5377 (N_5377,N_1240,N_3281);
nand U5378 (N_5378,N_3446,N_708);
nor U5379 (N_5379,N_1046,N_182);
nor U5380 (N_5380,N_4017,N_3086);
nor U5381 (N_5381,N_661,N_2596);
or U5382 (N_5382,N_4144,N_2477);
xnor U5383 (N_5383,N_1404,N_3588);
or U5384 (N_5384,N_2405,N_2884);
xnor U5385 (N_5385,N_353,N_2850);
nand U5386 (N_5386,N_759,N_1415);
and U5387 (N_5387,N_3469,N_3374);
xnor U5388 (N_5388,N_4114,N_119);
nor U5389 (N_5389,N_3080,N_2734);
or U5390 (N_5390,N_3932,N_4922);
nand U5391 (N_5391,N_3774,N_3659);
and U5392 (N_5392,N_1957,N_1091);
xor U5393 (N_5393,N_2335,N_1799);
and U5394 (N_5394,N_1850,N_30);
or U5395 (N_5395,N_3909,N_1115);
nand U5396 (N_5396,N_4267,N_2782);
nor U5397 (N_5397,N_3267,N_1090);
nor U5398 (N_5398,N_220,N_377);
nor U5399 (N_5399,N_213,N_3786);
nor U5400 (N_5400,N_4878,N_1098);
nand U5401 (N_5401,N_1732,N_4212);
xor U5402 (N_5402,N_299,N_4948);
nor U5403 (N_5403,N_3679,N_4325);
nand U5404 (N_5404,N_3045,N_2064);
nor U5405 (N_5405,N_4961,N_2677);
or U5406 (N_5406,N_3565,N_1937);
or U5407 (N_5407,N_1378,N_4419);
or U5408 (N_5408,N_962,N_2273);
xnor U5409 (N_5409,N_2160,N_4615);
and U5410 (N_5410,N_2758,N_2067);
and U5411 (N_5411,N_1614,N_2127);
and U5412 (N_5412,N_3172,N_3343);
nor U5413 (N_5413,N_1919,N_430);
and U5414 (N_5414,N_3076,N_4243);
or U5415 (N_5415,N_3,N_2042);
or U5416 (N_5416,N_1407,N_960);
xor U5417 (N_5417,N_3005,N_1487);
nand U5418 (N_5418,N_3330,N_1037);
nand U5419 (N_5419,N_1336,N_2402);
nor U5420 (N_5420,N_1930,N_1590);
nand U5421 (N_5421,N_1769,N_3164);
xnor U5422 (N_5422,N_4882,N_2660);
and U5423 (N_5423,N_2939,N_1679);
nor U5424 (N_5424,N_4590,N_2536);
and U5425 (N_5425,N_652,N_2600);
xor U5426 (N_5426,N_350,N_3943);
nand U5427 (N_5427,N_2033,N_4587);
nor U5428 (N_5428,N_3304,N_4913);
nand U5429 (N_5429,N_1777,N_1973);
nor U5430 (N_5430,N_3351,N_1179);
nand U5431 (N_5431,N_4971,N_4240);
nand U5432 (N_5432,N_916,N_2865);
nor U5433 (N_5433,N_1066,N_3377);
and U5434 (N_5434,N_4552,N_2968);
or U5435 (N_5435,N_1298,N_3490);
nor U5436 (N_5436,N_4476,N_2566);
xor U5437 (N_5437,N_2878,N_1131);
and U5438 (N_5438,N_4319,N_2136);
xor U5439 (N_5439,N_3919,N_4323);
nand U5440 (N_5440,N_2119,N_3185);
xor U5441 (N_5441,N_3258,N_4206);
or U5442 (N_5442,N_847,N_1072);
xnor U5443 (N_5443,N_4224,N_4534);
nor U5444 (N_5444,N_2869,N_3606);
or U5445 (N_5445,N_533,N_4020);
or U5446 (N_5446,N_4146,N_2817);
or U5447 (N_5447,N_276,N_148);
nand U5448 (N_5448,N_4094,N_4427);
nor U5449 (N_5449,N_2547,N_1125);
xnor U5450 (N_5450,N_2787,N_142);
nand U5451 (N_5451,N_4550,N_2924);
and U5452 (N_5452,N_2807,N_4975);
xnor U5453 (N_5453,N_3513,N_3289);
or U5454 (N_5454,N_2074,N_4504);
nand U5455 (N_5455,N_2762,N_147);
and U5456 (N_5456,N_2429,N_3356);
nor U5457 (N_5457,N_3571,N_1688);
xor U5458 (N_5458,N_4839,N_1954);
xor U5459 (N_5459,N_2187,N_4468);
and U5460 (N_5460,N_1712,N_2634);
nand U5461 (N_5461,N_1063,N_3380);
xor U5462 (N_5462,N_1663,N_1753);
and U5463 (N_5463,N_4635,N_378);
nand U5464 (N_5464,N_1576,N_2005);
or U5465 (N_5465,N_2035,N_2353);
nand U5466 (N_5466,N_2742,N_4411);
xnor U5467 (N_5467,N_2498,N_1305);
and U5468 (N_5468,N_926,N_4235);
nor U5469 (N_5469,N_3596,N_3551);
xnor U5470 (N_5470,N_2361,N_2034);
or U5471 (N_5471,N_2027,N_948);
nor U5472 (N_5472,N_1062,N_4136);
nand U5473 (N_5473,N_2904,N_1794);
nor U5474 (N_5474,N_870,N_172);
nor U5475 (N_5475,N_1,N_312);
xor U5476 (N_5476,N_3471,N_1490);
nor U5477 (N_5477,N_33,N_1959);
nand U5478 (N_5478,N_4169,N_200);
nor U5479 (N_5479,N_3101,N_1691);
and U5480 (N_5480,N_1568,N_4197);
nand U5481 (N_5481,N_4679,N_3742);
and U5482 (N_5482,N_557,N_997);
xor U5483 (N_5483,N_3843,N_3667);
nand U5484 (N_5484,N_2638,N_4811);
and U5485 (N_5485,N_490,N_3647);
nor U5486 (N_5486,N_3651,N_897);
xnor U5487 (N_5487,N_1935,N_3755);
and U5488 (N_5488,N_1245,N_1246);
and U5489 (N_5489,N_679,N_4612);
and U5490 (N_5490,N_1324,N_684);
nand U5491 (N_5491,N_249,N_3697);
and U5492 (N_5492,N_2999,N_2814);
or U5493 (N_5493,N_2862,N_3756);
nor U5494 (N_5494,N_4458,N_3382);
nand U5495 (N_5495,N_2340,N_3113);
xnor U5496 (N_5496,N_3747,N_1671);
nor U5497 (N_5497,N_4295,N_3088);
nor U5498 (N_5498,N_2506,N_3323);
nand U5499 (N_5499,N_1711,N_4953);
nor U5500 (N_5500,N_1536,N_667);
nor U5501 (N_5501,N_1061,N_1301);
nor U5502 (N_5502,N_783,N_178);
and U5503 (N_5503,N_2475,N_1704);
xnor U5504 (N_5504,N_3117,N_817);
nand U5505 (N_5505,N_2207,N_1418);
and U5506 (N_5506,N_3675,N_2260);
and U5507 (N_5507,N_263,N_3771);
or U5508 (N_5508,N_3413,N_3077);
or U5509 (N_5509,N_2723,N_2987);
or U5510 (N_5510,N_3870,N_4215);
nor U5511 (N_5511,N_1622,N_562);
nand U5512 (N_5512,N_793,N_515);
nand U5513 (N_5513,N_4365,N_3436);
nand U5514 (N_5514,N_1641,N_3552);
nor U5515 (N_5515,N_3183,N_283);
or U5516 (N_5516,N_4651,N_4426);
or U5517 (N_5517,N_1852,N_1129);
xor U5518 (N_5518,N_180,N_1812);
nor U5519 (N_5519,N_4059,N_4840);
or U5520 (N_5520,N_3831,N_1609);
or U5521 (N_5521,N_2054,N_3657);
nand U5522 (N_5522,N_4881,N_2158);
xnor U5523 (N_5523,N_1990,N_4647);
nor U5524 (N_5524,N_3326,N_575);
or U5525 (N_5525,N_1766,N_886);
nor U5526 (N_5526,N_1451,N_4991);
or U5527 (N_5527,N_1114,N_11);
xnor U5528 (N_5528,N_3981,N_3873);
and U5529 (N_5529,N_4799,N_526);
and U5530 (N_5530,N_3259,N_813);
or U5531 (N_5531,N_3912,N_4400);
xor U5532 (N_5532,N_4,N_3309);
or U5533 (N_5533,N_725,N_32);
nand U5534 (N_5534,N_1494,N_2072);
and U5535 (N_5535,N_1822,N_488);
and U5536 (N_5536,N_3311,N_4290);
and U5537 (N_5537,N_1876,N_395);
nor U5538 (N_5538,N_1547,N_3477);
nor U5539 (N_5539,N_1923,N_2167);
or U5540 (N_5540,N_3369,N_3623);
or U5541 (N_5541,N_3977,N_2513);
nor U5542 (N_5542,N_2932,N_4432);
xor U5543 (N_5543,N_3669,N_983);
xnor U5544 (N_5544,N_1024,N_3611);
nor U5545 (N_5545,N_2617,N_2407);
xor U5546 (N_5546,N_54,N_1296);
nor U5547 (N_5547,N_3194,N_1127);
nor U5548 (N_5548,N_2567,N_4621);
and U5549 (N_5549,N_2431,N_4076);
nand U5550 (N_5550,N_3052,N_938);
nand U5551 (N_5551,N_2331,N_2934);
or U5552 (N_5552,N_4591,N_3303);
and U5553 (N_5553,N_4071,N_1887);
nand U5554 (N_5554,N_2674,N_2531);
and U5555 (N_5555,N_216,N_110);
nand U5556 (N_5556,N_3114,N_1797);
or U5557 (N_5557,N_4619,N_2820);
xnor U5558 (N_5558,N_2385,N_2910);
or U5559 (N_5559,N_2546,N_3075);
nor U5560 (N_5560,N_2375,N_4521);
or U5561 (N_5561,N_827,N_389);
nor U5562 (N_5562,N_2441,N_1955);
nand U5563 (N_5563,N_401,N_3054);
nand U5564 (N_5564,N_1033,N_4013);
and U5565 (N_5565,N_4460,N_672);
nor U5566 (N_5566,N_494,N_1174);
and U5567 (N_5567,N_2529,N_35);
nor U5568 (N_5568,N_2585,N_3709);
xnor U5569 (N_5569,N_1844,N_292);
and U5570 (N_5570,N_571,N_550);
nand U5571 (N_5571,N_2857,N_1364);
and U5572 (N_5572,N_173,N_1271);
xor U5573 (N_5573,N_3096,N_624);
nand U5574 (N_5574,N_4894,N_1307);
and U5575 (N_5575,N_1467,N_4624);
nor U5576 (N_5576,N_2898,N_2030);
nand U5577 (N_5577,N_3847,N_4408);
nor U5578 (N_5578,N_227,N_1286);
and U5579 (N_5579,N_194,N_3724);
and U5580 (N_5580,N_2533,N_1138);
xor U5581 (N_5581,N_863,N_1459);
or U5582 (N_5582,N_3630,N_595);
nand U5583 (N_5583,N_3039,N_2197);
or U5584 (N_5584,N_2080,N_588);
nor U5585 (N_5585,N_3150,N_777);
nor U5586 (N_5586,N_1714,N_4161);
or U5587 (N_5587,N_4821,N_3740);
xnor U5588 (N_5588,N_2502,N_3779);
and U5589 (N_5589,N_3850,N_1354);
and U5590 (N_5590,N_3934,N_840);
xor U5591 (N_5591,N_4526,N_3357);
or U5592 (N_5592,N_2130,N_3569);
nor U5593 (N_5593,N_862,N_4613);
and U5594 (N_5594,N_1848,N_922);
xnor U5595 (N_5595,N_2082,N_738);
nor U5596 (N_5596,N_1178,N_1517);
nand U5597 (N_5597,N_390,N_3735);
or U5598 (N_5598,N_3256,N_189);
xnor U5599 (N_5599,N_4598,N_1981);
xnor U5600 (N_5600,N_2689,N_14);
nand U5601 (N_5601,N_3278,N_4564);
nor U5602 (N_5602,N_944,N_1465);
nand U5603 (N_5603,N_4807,N_996);
or U5604 (N_5604,N_3338,N_1310);
nand U5605 (N_5605,N_3798,N_465);
nor U5606 (N_5606,N_4445,N_807);
nor U5607 (N_5607,N_4687,N_4802);
and U5608 (N_5608,N_721,N_1612);
or U5609 (N_5609,N_427,N_3160);
nand U5610 (N_5610,N_4492,N_3033);
nand U5611 (N_5611,N_2155,N_4812);
or U5612 (N_5612,N_1493,N_702);
and U5613 (N_5613,N_3860,N_4321);
xnor U5614 (N_5614,N_2378,N_600);
nor U5615 (N_5615,N_874,N_3046);
or U5616 (N_5616,N_3955,N_3957);
nand U5617 (N_5617,N_3908,N_4401);
nor U5618 (N_5618,N_685,N_4569);
or U5619 (N_5619,N_456,N_844);
or U5620 (N_5620,N_753,N_464);
nor U5621 (N_5621,N_4586,N_3426);
and U5622 (N_5622,N_2653,N_2322);
nand U5623 (N_5623,N_651,N_3272);
xnor U5624 (N_5624,N_1484,N_3661);
and U5625 (N_5625,N_1333,N_1725);
nor U5626 (N_5626,N_2631,N_4297);
or U5627 (N_5627,N_4258,N_4376);
xnor U5628 (N_5628,N_241,N_4091);
nor U5629 (N_5629,N_1249,N_3696);
nor U5630 (N_5630,N_2292,N_107);
xnor U5631 (N_5631,N_4389,N_553);
xor U5632 (N_5632,N_2582,N_1360);
nand U5633 (N_5633,N_1960,N_3243);
nor U5634 (N_5634,N_136,N_4510);
nor U5635 (N_5635,N_3116,N_4417);
and U5636 (N_5636,N_2503,N_2958);
and U5637 (N_5637,N_4292,N_2561);
or U5638 (N_5638,N_4853,N_4628);
and U5639 (N_5639,N_3693,N_3910);
nand U5640 (N_5640,N_3125,N_1096);
nor U5641 (N_5641,N_1223,N_743);
nand U5642 (N_5642,N_1142,N_210);
xor U5643 (N_5643,N_4798,N_4373);
or U5644 (N_5644,N_914,N_3881);
xor U5645 (N_5645,N_2428,N_2825);
nor U5646 (N_5646,N_4801,N_3173);
or U5647 (N_5647,N_3857,N_4560);
nand U5648 (N_5648,N_3512,N_4008);
and U5649 (N_5649,N_4982,N_654);
or U5650 (N_5650,N_2593,N_4764);
nor U5651 (N_5651,N_4937,N_165);
xnor U5652 (N_5652,N_105,N_2099);
nor U5653 (N_5653,N_1170,N_206);
nand U5654 (N_5654,N_4783,N_3949);
or U5655 (N_5655,N_969,N_2181);
or U5656 (N_5656,N_4214,N_4633);
or U5657 (N_5657,N_569,N_2162);
and U5658 (N_5658,N_2779,N_3188);
or U5659 (N_5659,N_4037,N_4507);
nor U5660 (N_5660,N_3950,N_3022);
xor U5661 (N_5661,N_3600,N_1137);
nand U5662 (N_5662,N_829,N_3334);
xor U5663 (N_5663,N_4085,N_2735);
nor U5664 (N_5664,N_540,N_1105);
or U5665 (N_5665,N_3107,N_3074);
and U5666 (N_5666,N_4776,N_3386);
and U5667 (N_5667,N_1425,N_3402);
xor U5668 (N_5668,N_3047,N_625);
nor U5669 (N_5669,N_3120,N_1495);
xnor U5670 (N_5670,N_2921,N_2285);
and U5671 (N_5671,N_4578,N_145);
and U5672 (N_5672,N_4571,N_3638);
xnor U5673 (N_5673,N_4107,N_3929);
nand U5674 (N_5674,N_4732,N_379);
nor U5675 (N_5675,N_2471,N_168);
nand U5676 (N_5676,N_4111,N_2426);
nor U5677 (N_5677,N_4164,N_3136);
nand U5678 (N_5678,N_4589,N_158);
xor U5679 (N_5679,N_2223,N_4497);
or U5680 (N_5680,N_4580,N_3734);
and U5681 (N_5681,N_4850,N_1899);
nand U5682 (N_5682,N_711,N_267);
xor U5683 (N_5683,N_797,N_1748);
and U5684 (N_5684,N_1005,N_3953);
or U5685 (N_5685,N_605,N_1731);
xor U5686 (N_5686,N_3181,N_2926);
or U5687 (N_5687,N_3836,N_3020);
or U5688 (N_5688,N_3285,N_4864);
xor U5689 (N_5689,N_4599,N_3153);
nand U5690 (N_5690,N_2423,N_2221);
nand U5691 (N_5691,N_1543,N_3168);
xnor U5692 (N_5692,N_751,N_4897);
nor U5693 (N_5693,N_156,N_4167);
and U5694 (N_5694,N_1673,N_1719);
xor U5695 (N_5695,N_4880,N_2248);
or U5696 (N_5696,N_1374,N_1901);
xnor U5697 (N_5697,N_3582,N_593);
and U5698 (N_5698,N_3654,N_3222);
xor U5699 (N_5699,N_883,N_4181);
xnor U5700 (N_5700,N_4835,N_935);
or U5701 (N_5701,N_4883,N_1575);
or U5702 (N_5702,N_3104,N_4785);
nor U5703 (N_5703,N_2313,N_4846);
nand U5704 (N_5704,N_2457,N_4516);
xor U5705 (N_5705,N_3292,N_3633);
and U5706 (N_5706,N_2803,N_1248);
nor U5707 (N_5707,N_905,N_2626);
and U5708 (N_5708,N_2965,N_3723);
or U5709 (N_5709,N_3685,N_4353);
nor U5710 (N_5710,N_4143,N_3924);
nor U5711 (N_5711,N_140,N_270);
or U5712 (N_5712,N_804,N_2590);
and U5713 (N_5713,N_1537,N_47);
nand U5714 (N_5714,N_909,N_3058);
nor U5715 (N_5715,N_875,N_3684);
and U5716 (N_5716,N_1111,N_1696);
nor U5717 (N_5717,N_4448,N_2679);
and U5718 (N_5718,N_1055,N_3365);
nand U5719 (N_5719,N_756,N_1687);
and U5720 (N_5720,N_159,N_3337);
nand U5721 (N_5721,N_4318,N_2894);
nand U5722 (N_5722,N_3970,N_251);
or U5723 (N_5723,N_1735,N_4372);
or U5724 (N_5724,N_3094,N_3417);
nand U5725 (N_5725,N_3036,N_4641);
xor U5726 (N_5726,N_936,N_4780);
xor U5727 (N_5727,N_1201,N_92);
or U5728 (N_5728,N_1339,N_4538);
or U5729 (N_5729,N_4796,N_508);
or U5730 (N_5730,N_1155,N_3475);
nor U5731 (N_5731,N_4666,N_4771);
nor U5732 (N_5732,N_443,N_788);
nor U5733 (N_5733,N_1952,N_167);
or U5734 (N_5734,N_2843,N_1692);
or U5735 (N_5735,N_3344,N_4932);
or U5736 (N_5736,N_1967,N_2883);
and U5737 (N_5737,N_2947,N_4000);
or U5738 (N_5738,N_1838,N_4387);
nand U5739 (N_5739,N_4847,N_55);
nor U5740 (N_5740,N_3485,N_1452);
xor U5741 (N_5741,N_604,N_3673);
nand U5742 (N_5742,N_1833,N_3961);
or U5743 (N_5743,N_2367,N_911);
nor U5744 (N_5744,N_1561,N_2720);
and U5745 (N_5745,N_384,N_188);
and U5746 (N_5746,N_3862,N_842);
nand U5747 (N_5747,N_4470,N_3035);
or U5748 (N_5748,N_4191,N_4053);
xnor U5749 (N_5749,N_1931,N_1603);
nand U5750 (N_5750,N_3672,N_24);
nand U5751 (N_5751,N_4029,N_3942);
nor U5752 (N_5752,N_2818,N_3974);
nor U5753 (N_5753,N_1816,N_3549);
and U5754 (N_5754,N_2303,N_2086);
and U5755 (N_5755,N_2644,N_3066);
nor U5756 (N_5756,N_749,N_1573);
xnor U5757 (N_5757,N_499,N_1685);
xor U5758 (N_5758,N_4152,N_741);
and U5759 (N_5759,N_4959,N_1658);
nor U5760 (N_5760,N_4962,N_919);
nor U5761 (N_5761,N_1348,N_3274);
or U5762 (N_5762,N_4173,N_1380);
and U5763 (N_5763,N_762,N_3738);
or U5764 (N_5764,N_4770,N_297);
or U5765 (N_5765,N_3533,N_1104);
xor U5766 (N_5766,N_536,N_295);
and U5767 (N_5767,N_3766,N_2574);
xor U5768 (N_5768,N_3603,N_681);
and U5769 (N_5769,N_1965,N_1650);
or U5770 (N_5770,N_3430,N_2589);
or U5771 (N_5771,N_3496,N_362);
or U5772 (N_5772,N_1770,N_4452);
or U5773 (N_5773,N_4188,N_1600);
nor U5774 (N_5774,N_3822,N_2748);
nor U5775 (N_5775,N_1045,N_3182);
or U5776 (N_5776,N_77,N_2261);
or U5777 (N_5777,N_4540,N_585);
xnor U5778 (N_5778,N_4179,N_2112);
nor U5779 (N_5779,N_1968,N_1502);
xnor U5780 (N_5780,N_2584,N_1861);
and U5781 (N_5781,N_2090,N_437);
and U5782 (N_5782,N_3637,N_3649);
xor U5783 (N_5783,N_1740,N_2284);
nor U5784 (N_5784,N_4756,N_4758);
or U5785 (N_5785,N_4471,N_2619);
or U5786 (N_5786,N_2578,N_1186);
or U5787 (N_5787,N_1701,N_3867);
and U5788 (N_5788,N_3174,N_2740);
and U5789 (N_5789,N_4092,N_4872);
nor U5790 (N_5790,N_4097,N_611);
and U5791 (N_5791,N_3872,N_2682);
or U5792 (N_5792,N_2458,N_732);
nand U5793 (N_5793,N_819,N_890);
nand U5794 (N_5794,N_2316,N_4190);
nand U5795 (N_5795,N_4833,N_4450);
xor U5796 (N_5796,N_918,N_1429);
nor U5797 (N_5797,N_1080,N_828);
nor U5798 (N_5798,N_2434,N_2069);
nand U5799 (N_5799,N_4227,N_4938);
or U5800 (N_5800,N_2406,N_265);
and U5801 (N_5801,N_365,N_4575);
and U5802 (N_5802,N_311,N_1047);
and U5803 (N_5803,N_3620,N_2860);
or U5804 (N_5804,N_2832,N_1160);
nand U5805 (N_5805,N_3626,N_2627);
nand U5806 (N_5806,N_338,N_2046);
nor U5807 (N_5807,N_771,N_3682);
or U5808 (N_5808,N_1513,N_4648);
nand U5809 (N_5809,N_4449,N_4981);
nor U5810 (N_5810,N_4754,N_4875);
and U5811 (N_5811,N_4402,N_4123);
or U5812 (N_5812,N_740,N_425);
nor U5813 (N_5813,N_2466,N_2073);
or U5814 (N_5814,N_4558,N_4247);
xor U5815 (N_5815,N_2214,N_4437);
xnor U5816 (N_5816,N_1269,N_3087);
or U5817 (N_5817,N_2956,N_2810);
nand U5818 (N_5818,N_3340,N_1936);
or U5819 (N_5819,N_1744,N_1087);
or U5820 (N_5820,N_2366,N_3370);
xor U5821 (N_5821,N_4597,N_4502);
and U5822 (N_5822,N_1267,N_4351);
nand U5823 (N_5823,N_3293,N_3902);
and U5824 (N_5824,N_3341,N_977);
xor U5825 (N_5825,N_3882,N_326);
nor U5826 (N_5826,N_2281,N_322);
or U5827 (N_5827,N_4737,N_1225);
nor U5828 (N_5828,N_4639,N_4300);
xor U5829 (N_5829,N_4259,N_581);
nand U5830 (N_5830,N_3228,N_1292);
and U5831 (N_5831,N_4170,N_3784);
and U5832 (N_5832,N_4063,N_2556);
and U5833 (N_5833,N_1321,N_3536);
nand U5834 (N_5834,N_1121,N_38);
xnor U5835 (N_5835,N_4919,N_4306);
nand U5836 (N_5836,N_4489,N_2488);
nand U5837 (N_5837,N_1520,N_4176);
and U5838 (N_5838,N_3598,N_3945);
or U5839 (N_5839,N_4070,N_2135);
or U5840 (N_5840,N_3414,N_1198);
or U5841 (N_5841,N_1587,N_1387);
or U5842 (N_5842,N_3716,N_4583);
xor U5843 (N_5843,N_628,N_3200);
xnor U5844 (N_5844,N_925,N_4461);
xor U5845 (N_5845,N_929,N_117);
nand U5846 (N_5846,N_4233,N_794);
xor U5847 (N_5847,N_411,N_3473);
nor U5848 (N_5848,N_2836,N_3159);
or U5849 (N_5849,N_284,N_3097);
or U5850 (N_5850,N_3119,N_1771);
xor U5851 (N_5851,N_724,N_616);
nor U5852 (N_5852,N_329,N_2952);
nand U5853 (N_5853,N_1477,N_2328);
and U5854 (N_5854,N_1680,N_3946);
xor U5855 (N_5855,N_649,N_4577);
xor U5856 (N_5856,N_3849,N_3901);
xor U5857 (N_5857,N_4478,N_580);
or U5858 (N_5858,N_4339,N_1664);
nor U5859 (N_5859,N_3423,N_3524);
or U5860 (N_5860,N_3363,N_2776);
nand U5861 (N_5861,N_4918,N_151);
xor U5862 (N_5862,N_1318,N_4429);
xor U5863 (N_5863,N_1447,N_2002);
nand U5864 (N_5864,N_4965,N_2895);
nand U5865 (N_5865,N_1212,N_4423);
nor U5866 (N_5866,N_4939,N_275);
and U5867 (N_5867,N_2709,N_3387);
or U5868 (N_5868,N_3959,N_2985);
xor U5869 (N_5869,N_2399,N_1312);
xnor U5870 (N_5870,N_4706,N_1535);
nand U5871 (N_5871,N_876,N_4915);
nor U5872 (N_5872,N_4198,N_2804);
nand U5873 (N_5873,N_1430,N_1290);
xor U5874 (N_5874,N_1229,N_3299);
nand U5875 (N_5875,N_4250,N_152);
xnor U5876 (N_5876,N_3545,N_4363);
nor U5877 (N_5877,N_2791,N_223);
nor U5878 (N_5878,N_4087,N_3312);
nand U5879 (N_5879,N_3879,N_1988);
nand U5880 (N_5880,N_2936,N_885);
nor U5881 (N_5881,N_1829,N_867);
nand U5882 (N_5882,N_2382,N_731);
and U5883 (N_5883,N_2358,N_4685);
nand U5884 (N_5884,N_1308,N_1359);
nand U5885 (N_5885,N_1314,N_718);
xor U5886 (N_5886,N_1879,N_4277);
nand U5887 (N_5887,N_3488,N_2790);
xor U5888 (N_5888,N_3676,N_3322);
nor U5889 (N_5889,N_4889,N_1064);
xnor U5890 (N_5890,N_4728,N_2530);
and U5891 (N_5891,N_791,N_420);
and U5892 (N_5892,N_1774,N_3237);
or U5893 (N_5893,N_1264,N_56);
and U5894 (N_5894,N_2238,N_3493);
and U5895 (N_5895,N_3449,N_1686);
xor U5896 (N_5896,N_2903,N_2120);
xor U5897 (N_5897,N_4724,N_4038);
or U5898 (N_5898,N_45,N_2131);
or U5899 (N_5899,N_3245,N_2094);
and U5900 (N_5900,N_1021,N_2510);
and U5901 (N_5901,N_4236,N_4867);
or U5902 (N_5902,N_2386,N_1709);
and U5903 (N_5903,N_4110,N_3925);
or U5904 (N_5904,N_2811,N_3518);
nand U5905 (N_5905,N_3800,N_1849);
and U5906 (N_5906,N_2409,N_3345);
xnor U5907 (N_5907,N_1368,N_4584);
nand U5908 (N_5908,N_4131,N_3564);
or U5909 (N_5909,N_3489,N_4089);
nor U5910 (N_5910,N_4064,N_3613);
or U5911 (N_5911,N_4529,N_1143);
nand U5912 (N_5912,N_3165,N_2771);
nand U5913 (N_5913,N_1880,N_3453);
nand U5914 (N_5914,N_2819,N_4547);
nand U5915 (N_5915,N_4178,N_821);
or U5916 (N_5916,N_1488,N_1023);
nand U5917 (N_5917,N_2185,N_792);
or U5918 (N_5918,N_81,N_3899);
nor U5919 (N_5919,N_3324,N_99);
xnor U5920 (N_5920,N_2822,N_315);
nor U5921 (N_5921,N_2216,N_1504);
xnor U5922 (N_5922,N_1874,N_457);
xor U5923 (N_5923,N_3585,N_2516);
and U5924 (N_5924,N_705,N_3572);
nor U5925 (N_5925,N_3464,N_541);
and U5926 (N_5926,N_1001,N_877);
and U5927 (N_5927,N_592,N_4700);
and U5928 (N_5928,N_2527,N_4125);
xor U5929 (N_5929,N_769,N_4608);
and U5930 (N_5930,N_2494,N_3346);
and U5931 (N_5931,N_2539,N_3558);
or U5932 (N_5932,N_3578,N_3632);
nor U5933 (N_5933,N_1491,N_822);
xnor U5934 (N_5934,N_4137,N_4093);
xor U5935 (N_5935,N_1551,N_462);
xnor U5936 (N_5936,N_2087,N_97);
nor U5937 (N_5937,N_3364,N_3541);
nand U5938 (N_5938,N_2096,N_1428);
nand U5939 (N_5939,N_825,N_4132);
or U5940 (N_5940,N_3913,N_4863);
and U5941 (N_5941,N_1745,N_3032);
or U5942 (N_5942,N_271,N_2334);
xor U5943 (N_5943,N_1896,N_3438);
nand U5944 (N_5944,N_2177,N_261);
nand U5945 (N_5945,N_4711,N_3355);
and U5946 (N_5946,N_2983,N_2070);
nor U5947 (N_5947,N_4431,N_976);
or U5948 (N_5948,N_1516,N_931);
and U5949 (N_5949,N_4051,N_187);
nor U5950 (N_5950,N_2538,N_1557);
xnor U5951 (N_5951,N_4356,N_2295);
or U5952 (N_5952,N_4231,N_3093);
xor U5953 (N_5953,N_502,N_4344);
or U5954 (N_5954,N_1185,N_2960);
and U5955 (N_5955,N_4095,N_1907);
xor U5956 (N_5956,N_6,N_4893);
and U5957 (N_5957,N_1120,N_3189);
or U5958 (N_5958,N_2780,N_3980);
nor U5959 (N_5959,N_1817,N_3124);
or U5960 (N_5960,N_1941,N_1898);
or U5961 (N_5961,N_4264,N_2347);
or U5962 (N_5962,N_3884,N_1256);
and U5963 (N_5963,N_1943,N_4870);
or U5964 (N_5964,N_3764,N_25);
or U5965 (N_5965,N_367,N_214);
nor U5966 (N_5966,N_4308,N_1815);
xnor U5967 (N_5967,N_3550,N_3466);
and U5968 (N_5968,N_185,N_380);
or U5969 (N_5969,N_599,N_4759);
xor U5970 (N_5970,N_4968,N_90);
xnor U5971 (N_5971,N_286,N_4031);
or U5972 (N_5972,N_4794,N_3399);
xor U5973 (N_5973,N_4528,N_2011);
or U5974 (N_5974,N_4992,N_2036);
nor U5975 (N_5975,N_2057,N_956);
or U5976 (N_5976,N_1894,N_752);
and U5977 (N_5977,N_3759,N_1016);
nand U5978 (N_5978,N_3834,N_4644);
nor U5979 (N_5979,N_39,N_1401);
nor U5980 (N_5980,N_2521,N_3793);
or U5981 (N_5981,N_4042,N_4443);
xor U5982 (N_5982,N_1765,N_4393);
xnor U5983 (N_5983,N_520,N_3123);
xnor U5984 (N_5984,N_3431,N_1945);
or U5985 (N_5985,N_4990,N_3061);
or U5986 (N_5986,N_3412,N_4773);
or U5987 (N_5987,N_1132,N_4629);
and U5988 (N_5988,N_3481,N_4527);
or U5989 (N_5989,N_2866,N_4696);
nand U5990 (N_5990,N_810,N_4984);
nand U5991 (N_5991,N_2315,N_979);
xnor U5992 (N_5992,N_1122,N_1280);
nor U5993 (N_5993,N_2639,N_282);
nand U5994 (N_5994,N_4326,N_2685);
or U5995 (N_5995,N_3621,N_4741);
nor U5996 (N_5996,N_1964,N_3320);
or U5997 (N_5997,N_1085,N_4740);
or U5998 (N_5998,N_2514,N_3972);
and U5999 (N_5999,N_3440,N_1042);
xnor U6000 (N_6000,N_1629,N_860);
or U6001 (N_6001,N_3814,N_2710);
and U6002 (N_6002,N_3492,N_2276);
or U6003 (N_6003,N_2023,N_787);
and U6004 (N_6004,N_3805,N_313);
xor U6005 (N_6005,N_3589,N_1747);
nor U6006 (N_6006,N_2834,N_745);
xnor U6007 (N_6007,N_1156,N_4542);
and U6008 (N_6008,N_1693,N_3192);
xor U6009 (N_6009,N_3880,N_4281);
nor U6010 (N_6010,N_2540,N_642);
nor U6011 (N_6011,N_501,N_1558);
nand U6012 (N_6012,N_3770,N_1388);
and U6013 (N_6013,N_1167,N_4084);
xor U6014 (N_6014,N_789,N_4946);
xor U6015 (N_6015,N_3305,N_507);
xor U6016 (N_6016,N_160,N_3332);
xnor U6017 (N_6017,N_88,N_3067);
xor U6018 (N_6018,N_4665,N_3068);
and U6019 (N_6019,N_2031,N_1674);
nand U6020 (N_6020,N_1826,N_4327);
and U6021 (N_6021,N_4677,N_2125);
nor U6022 (N_6022,N_2274,N_4963);
or U6023 (N_6023,N_4012,N_760);
and U6024 (N_6024,N_4350,N_1094);
and U6025 (N_6025,N_1496,N_4256);
or U6026 (N_6026,N_3757,N_2874);
nand U6027 (N_6027,N_3646,N_1191);
nand U6028 (N_6028,N_4302,N_4331);
nor U6029 (N_6029,N_2247,N_3333);
and U6030 (N_6030,N_2305,N_853);
nand U6031 (N_6031,N_2201,N_647);
nor U6032 (N_6032,N_2195,N_4390);
nand U6033 (N_6033,N_4337,N_121);
nand U6034 (N_6034,N_2548,N_1503);
or U6035 (N_6035,N_4477,N_554);
xnor U6036 (N_6036,N_1870,N_746);
xnor U6037 (N_6037,N_4384,N_1541);
xor U6038 (N_6038,N_4723,N_1411);
nor U6039 (N_6039,N_2726,N_4827);
and U6040 (N_6040,N_511,N_2752);
and U6041 (N_6041,N_784,N_522);
nor U6042 (N_6042,N_28,N_4699);
nand U6043 (N_6043,N_2913,N_419);
nand U6044 (N_6044,N_3978,N_3405);
and U6045 (N_6045,N_1625,N_2594);
or U6046 (N_6046,N_3089,N_257);
or U6047 (N_6047,N_504,N_166);
xor U6048 (N_6048,N_1802,N_2792);
xnor U6049 (N_6049,N_4710,N_4822);
nor U6050 (N_6050,N_4007,N_770);
nor U6051 (N_6051,N_1630,N_2747);
and U6052 (N_6052,N_1486,N_4034);
or U6053 (N_6053,N_4793,N_1385);
nor U6054 (N_6054,N_1828,N_4887);
or U6055 (N_6055,N_2588,N_2264);
or U6056 (N_6056,N_3134,N_1095);
and U6057 (N_6057,N_4742,N_2823);
nor U6058 (N_6058,N_3996,N_932);
xor U6059 (N_6059,N_790,N_18);
and U6060 (N_6060,N_4681,N_3206);
and U6061 (N_6061,N_1836,N_4970);
and U6062 (N_6062,N_719,N_577);
nand U6063 (N_6063,N_765,N_3888);
or U6064 (N_6064,N_4455,N_3744);
nand U6065 (N_6065,N_871,N_3855);
and U6066 (N_6066,N_4592,N_2308);
nor U6067 (N_6067,N_290,N_2920);
nand U6068 (N_6068,N_3121,N_902);
or U6069 (N_6069,N_2432,N_324);
nand U6070 (N_6070,N_4733,N_0);
nand U6071 (N_6071,N_1845,N_3904);
nor U6072 (N_6072,N_4315,N_1207);
nand U6073 (N_6073,N_2465,N_2249);
xnor U6074 (N_6074,N_274,N_2343);
nand U6075 (N_6075,N_3282,N_2727);
nor U6076 (N_6076,N_4368,N_4856);
nand U6077 (N_6077,N_832,N_2905);
or U6078 (N_6078,N_631,N_1379);
and U6079 (N_6079,N_3210,N_4509);
nor U6080 (N_6080,N_2575,N_3832);
and U6081 (N_6081,N_3775,N_3732);
xor U6082 (N_6082,N_1730,N_115);
nor U6083 (N_6083,N_3283,N_4352);
or U6084 (N_6084,N_1257,N_1437);
nor U6085 (N_6085,N_2229,N_2354);
and U6086 (N_6086,N_2263,N_1092);
xor U6087 (N_6087,N_4817,N_64);
nor U6088 (N_6088,N_839,N_2887);
nand U6089 (N_6089,N_3958,N_3990);
nand U6090 (N_6090,N_1350,N_4406);
xnor U6091 (N_6091,N_706,N_1153);
and U6092 (N_6092,N_2269,N_2601);
xnor U6093 (N_6093,N_4023,N_1109);
xnor U6094 (N_6094,N_3725,N_4298);
xor U6095 (N_6095,N_1468,N_484);
or U6096 (N_6096,N_1749,N_2079);
and U6097 (N_6097,N_958,N_3802);
nand U6098 (N_6098,N_1700,N_3982);
and U6099 (N_6099,N_1500,N_1266);
and U6100 (N_6100,N_3917,N_3812);
nand U6101 (N_6101,N_1322,N_242);
xnor U6102 (N_6102,N_3636,N_207);
or U6103 (N_6103,N_618,N_2453);
nand U6104 (N_6104,N_1634,N_768);
nand U6105 (N_6105,N_1017,N_3947);
and U6106 (N_6106,N_970,N_1666);
nand U6107 (N_6107,N_1739,N_3617);
or U6108 (N_6108,N_2992,N_3537);
xor U6109 (N_6109,N_3914,N_3220);
nor U6110 (N_6110,N_3092,N_3758);
and U6111 (N_6111,N_2688,N_1947);
nand U6112 (N_6112,N_4533,N_2418);
nor U6113 (N_6113,N_1022,N_3710);
xnor U6114 (N_6114,N_2270,N_4467);
nand U6115 (N_6115,N_474,N_2006);
and U6116 (N_6116,N_3421,N_1159);
nor U6117 (N_6117,N_4322,N_4525);
xor U6118 (N_6118,N_2129,N_3671);
and U6119 (N_6119,N_2394,N_3391);
and U6120 (N_6120,N_3642,N_3239);
nor U6121 (N_6121,N_2957,N_4462);
and U6122 (N_6122,N_1997,N_2591);
xor U6123 (N_6123,N_632,N_3522);
nor U6124 (N_6124,N_1217,N_1706);
nand U6125 (N_6125,N_4814,N_3993);
nand U6126 (N_6126,N_4769,N_2048);
or U6127 (N_6127,N_1552,N_3226);
xor U6128 (N_6128,N_2667,N_4006);
or U6129 (N_6129,N_1840,N_1103);
or U6130 (N_6130,N_3681,N_4342);
or U6131 (N_6131,N_164,N_818);
nor U6132 (N_6132,N_3169,N_1346);
nand U6133 (N_6133,N_2580,N_211);
nor U6134 (N_6134,N_3048,N_1088);
nor U6135 (N_6135,N_3874,N_394);
xor U6136 (N_6136,N_656,N_2012);
and U6137 (N_6137,N_2641,N_2937);
nand U6138 (N_6138,N_3273,N_3794);
nor U6139 (N_6139,N_4757,N_3790);
and U6140 (N_6140,N_2473,N_302);
nor U6141 (N_6141,N_2332,N_1426);
nand U6142 (N_6142,N_1948,N_2848);
or U6143 (N_6143,N_2103,N_4441);
or U6144 (N_6144,N_2333,N_3689);
nand U6145 (N_6145,N_3410,N_75);
xor U6146 (N_6146,N_3845,N_1038);
or U6147 (N_6147,N_737,N_3017);
or U6148 (N_6148,N_209,N_1875);
and U6149 (N_6149,N_615,N_2722);
nor U6150 (N_6150,N_2745,N_2280);
and U6151 (N_6151,N_1998,N_305);
or U6152 (N_6152,N_1979,N_2456);
nor U6153 (N_6153,N_1668,N_4481);
xor U6154 (N_6154,N_3527,N_3085);
or U6155 (N_6155,N_3634,N_4253);
nor U6156 (N_6156,N_3129,N_4015);
xor U6157 (N_6157,N_990,N_3031);
nand U6158 (N_6158,N_4168,N_2217);
nand U6159 (N_6159,N_4775,N_2670);
and U6160 (N_6160,N_3801,N_3906);
or U6161 (N_6161,N_3865,N_1851);
nor U6162 (N_6162,N_1130,N_415);
and U6163 (N_6163,N_2341,N_3404);
xor U6164 (N_6164,N_1089,N_137);
and U6165 (N_6165,N_565,N_957);
nand U6166 (N_6166,N_2300,N_3988);
nand U6167 (N_6167,N_4148,N_2554);
nor U6168 (N_6168,N_4194,N_811);
nor U6169 (N_6169,N_806,N_2157);
or U6170 (N_6170,N_2559,N_3719);
or U6171 (N_6171,N_3976,N_703);
or U6172 (N_6172,N_964,N_1171);
nor U6173 (N_6173,N_4126,N_4692);
and U6174 (N_6174,N_1925,N_4303);
and U6175 (N_6175,N_1431,N_2760);
or U6176 (N_6176,N_3499,N_2552);
nor U6177 (N_6177,N_4186,N_1922);
or U6178 (N_6178,N_3263,N_601);
xor U6179 (N_6179,N_3219,N_3663);
and U6180 (N_6180,N_1273,N_2981);
nor U6181 (N_6181,N_3519,N_4357);
nor U6182 (N_6182,N_4645,N_497);
xnor U6183 (N_6183,N_3099,N_2398);
and U6184 (N_6184,N_1135,N_1112);
nor U6185 (N_6185,N_4977,N_2464);
nand U6186 (N_6186,N_4280,N_3434);
or U6187 (N_6187,N_1187,N_4313);
nand U6188 (N_6188,N_1795,N_1471);
or U6189 (N_6189,N_16,N_3717);
nor U6190 (N_6190,N_2668,N_622);
or U6191 (N_6191,N_4790,N_913);
xnor U6192 (N_6192,N_1351,N_3319);
or U6193 (N_6193,N_1511,N_1282);
nand U6194 (N_6194,N_534,N_1563);
xor U6195 (N_6195,N_1694,N_674);
nand U6196 (N_6196,N_3853,N_4689);
nor U6197 (N_6197,N_3408,N_4682);
xnor U6198 (N_6198,N_3425,N_175);
nor U6199 (N_6199,N_772,N_3390);
or U6200 (N_6200,N_4334,N_4819);
nand U6201 (N_6201,N_2873,N_1806);
and U6202 (N_6202,N_1866,N_3264);
or U6203 (N_6203,N_1604,N_2078);
or U6204 (N_6204,N_2982,N_4359);
or U6205 (N_6205,N_3664,N_4816);
xor U6206 (N_6206,N_161,N_4196);
and U6207 (N_6207,N_4697,N_3389);
or U6208 (N_6208,N_3983,N_2993);
nor U6209 (N_6209,N_3859,N_2794);
and U6210 (N_6210,N_1798,N_1386);
or U6211 (N_6211,N_2397,N_3521);
xnor U6212 (N_6212,N_608,N_4456);
or U6213 (N_6213,N_959,N_1259);
nor U6214 (N_6214,N_3543,N_2778);
and U6215 (N_6215,N_374,N_2872);
nand U6216 (N_6216,N_3604,N_4789);
nor U6217 (N_6217,N_620,N_2777);
or U6218 (N_6218,N_363,N_1905);
and U6219 (N_6219,N_715,N_3497);
xor U6220 (N_6220,N_1481,N_4581);
or U6221 (N_6221,N_388,N_590);
nor U6222 (N_6222,N_4782,N_3268);
nor U6223 (N_6223,N_4788,N_2528);
xor U6224 (N_6224,N_3100,N_131);
xnor U6225 (N_6225,N_1779,N_483);
and U6226 (N_6226,N_2708,N_4762);
or U6227 (N_6227,N_2192,N_3451);
xor U6228 (N_6228,N_359,N_664);
and U6229 (N_6229,N_2507,N_1315);
and U6230 (N_6230,N_435,N_4415);
nor U6231 (N_6231,N_1349,N_757);
and U6232 (N_6232,N_67,N_4674);
xor U6233 (N_6233,N_4289,N_1514);
xnor U6234 (N_6234,N_2938,N_4100);
and U6235 (N_6235,N_4001,N_4255);
nand U6236 (N_6236,N_4296,N_864);
xnor U6237 (N_6237,N_3176,N_1980);
or U6238 (N_6238,N_3378,N_3528);
and U6239 (N_6239,N_1270,N_334);
and U6240 (N_6240,N_1172,N_4036);
or U6241 (N_6241,N_4381,N_1515);
xor U6242 (N_6242,N_744,N_4690);
nand U6243 (N_6243,N_4083,N_3409);
and U6244 (N_6244,N_4969,N_1218);
nor U6245 (N_6245,N_177,N_1827);
and U6246 (N_6246,N_4014,N_422);
or U6247 (N_6247,N_3180,N_4655);
and U6248 (N_6248,N_1406,N_1971);
nor U6249 (N_6249,N_1260,N_4596);
or U6250 (N_6250,N_3625,N_2442);
nor U6251 (N_6251,N_2324,N_118);
nor U6252 (N_6252,N_3837,N_4743);
nand U6253 (N_6253,N_473,N_2694);
or U6254 (N_6254,N_4299,N_1041);
nand U6255 (N_6255,N_3907,N_3645);
nor U6256 (N_6256,N_3602,N_2637);
xnor U6257 (N_6257,N_3688,N_1065);
nor U6258 (N_6258,N_933,N_3297);
or U6259 (N_6259,N_3242,N_93);
and U6260 (N_6260,N_2630,N_2259);
xnor U6261 (N_6261,N_2016,N_135);
xor U6262 (N_6262,N_4211,N_3829);
nand U6263 (N_6263,N_1695,N_1608);
nand U6264 (N_6264,N_2288,N_1638);
xor U6265 (N_6265,N_2509,N_2040);
and U6266 (N_6266,N_2940,N_1009);
xor U6267 (N_6267,N_3487,N_2534);
or U6268 (N_6268,N_3939,N_1464);
nand U6269 (N_6269,N_2244,N_89);
xor U6270 (N_6270,N_2156,N_4338);
and U6271 (N_6271,N_680,N_3936);
nor U6272 (N_6272,N_4912,N_1710);
nand U6273 (N_6273,N_4066,N_4226);
nand U6274 (N_6274,N_834,N_3701);
nor U6275 (N_6275,N_1057,N_3640);
nor U6276 (N_6276,N_3575,N_303);
and U6277 (N_6277,N_2629,N_4228);
and U6278 (N_6278,N_1189,N_2422);
and U6279 (N_6279,N_2725,N_4563);
xnor U6280 (N_6280,N_2788,N_2154);
xnor U6281 (N_6281,N_408,N_3656);
and U6282 (N_6282,N_2911,N_639);
xor U6283 (N_6283,N_27,N_3167);
nand U6284 (N_6284,N_975,N_3509);
nor U6285 (N_6285,N_4057,N_445);
xor U6286 (N_6286,N_3702,N_477);
nand U6287 (N_6287,N_1631,N_2871);
nand U6288 (N_6288,N_1886,N_1811);
nor U6289 (N_6289,N_4716,N_476);
nand U6290 (N_6290,N_1441,N_4541);
and U6291 (N_6291,N_2623,N_1531);
or U6292 (N_6292,N_645,N_2770);
nand U6293 (N_6293,N_4354,N_1391);
xor U6294 (N_6294,N_403,N_453);
xor U6295 (N_6295,N_413,N_1818);
nand U6296 (N_6296,N_2286,N_3244);
nor U6297 (N_6297,N_1662,N_1983);
and U6298 (N_6298,N_4055,N_3327);
xor U6299 (N_6299,N_398,N_4739);
nand U6300 (N_6300,N_1665,N_237);
and U6301 (N_6301,N_2133,N_1803);
nor U6302 (N_6302,N_2505,N_4786);
and U6303 (N_6303,N_4928,N_3429);
nand U6304 (N_6304,N_4225,N_3310);
or U6305 (N_6305,N_1596,N_2949);
xor U6306 (N_6306,N_1556,N_523);
or U6307 (N_6307,N_4858,N_2893);
and U6308 (N_6308,N_1890,N_3162);
and U6309 (N_6309,N_3938,N_79);
and U6310 (N_6310,N_2598,N_621);
nor U6311 (N_6311,N_1723,N_2291);
or U6312 (N_6312,N_1398,N_3231);
nand U6313 (N_6313,N_2404,N_2809);
or U6314 (N_6314,N_2557,N_3601);
or U6315 (N_6315,N_3276,N_1843);
nor U6316 (N_6316,N_1859,N_2827);
nor U6317 (N_6317,N_469,N_858);
or U6318 (N_6318,N_892,N_2066);
nand U6319 (N_6319,N_4549,N_1521);
nor U6320 (N_6320,N_992,N_795);
nand U6321 (N_6321,N_1347,N_1708);
xnor U6322 (N_6322,N_4903,N_2959);
nor U6323 (N_6323,N_3300,N_1767);
nor U6324 (N_6324,N_1317,N_4329);
nor U6325 (N_6325,N_2656,N_1299);
nand U6326 (N_6326,N_287,N_4876);
nand U6327 (N_6327,N_434,N_1358);
nand U6328 (N_6328,N_535,N_4909);
nand U6329 (N_6329,N_3079,N_663);
nand U6330 (N_6330,N_898,N_4924);
or U6331 (N_6331,N_2789,N_3381);
nand U6332 (N_6332,N_4901,N_2242);
nand U6333 (N_6333,N_3441,N_4239);
or U6334 (N_6334,N_3373,N_3778);
and U6335 (N_6335,N_4708,N_3830);
xor U6336 (N_6336,N_496,N_1498);
nor U6337 (N_6337,N_3876,N_3858);
xnor U6338 (N_6338,N_2299,N_108);
and U6339 (N_6339,N_3041,N_1036);
xnor U6340 (N_6340,N_3643,N_2532);
and U6341 (N_6341,N_1251,N_70);
nand U6342 (N_6342,N_917,N_2049);
and U6343 (N_6343,N_3401,N_2669);
nor U6344 (N_6344,N_1157,N_4712);
xnor U6345 (N_6345,N_4026,N_4230);
and U6346 (N_6346,N_2395,N_314);
and U6347 (N_6347,N_4269,N_2013);
and U6348 (N_6348,N_4120,N_517);
or U6349 (N_6349,N_3705,N_2607);
nor U6350 (N_6350,N_2483,N_2765);
nor U6351 (N_6351,N_4438,N_4024);
or U6352 (N_6352,N_4219,N_3568);
nor U6353 (N_6353,N_3271,N_4556);
xor U6354 (N_6354,N_686,N_1435);
nor U6355 (N_6355,N_3502,N_57);
nand U6356 (N_6356,N_4394,N_3825);
nand U6357 (N_6357,N_2953,N_1893);
nand U6358 (N_6358,N_285,N_999);
xnor U6359 (N_6359,N_1117,N_1274);
nor U6360 (N_6360,N_3962,N_4703);
or U6361 (N_6361,N_1512,N_4848);
or U6362 (N_6362,N_1233,N_951);
nand U6363 (N_6363,N_2047,N_3820);
and U6364 (N_6364,N_190,N_3931);
or U6365 (N_6365,N_3000,N_4787);
and U6366 (N_6366,N_4282,N_279);
or U6367 (N_6367,N_355,N_3984);
nand U6368 (N_6368,N_4263,N_1567);
nor U6369 (N_6369,N_2440,N_141);
nor U6370 (N_6370,N_327,N_2706);
xnor U6371 (N_6371,N_1328,N_1661);
or U6372 (N_6372,N_984,N_2137);
nor U6373 (N_6373,N_2370,N_4382);
xor U6374 (N_6374,N_1448,N_1011);
nor U6375 (N_6375,N_4154,N_780);
nor U6376 (N_6376,N_138,N_4486);
nand U6377 (N_6377,N_4766,N_2237);
xor U6378 (N_6378,N_734,N_665);
nor U6379 (N_6379,N_4678,N_1015);
or U6380 (N_6380,N_3538,N_4261);
and U6381 (N_6381,N_1570,N_666);
and U6382 (N_6382,N_4543,N_2222);
xnor U6383 (N_6383,N_2293,N_2107);
or U6384 (N_6384,N_3721,N_3561);
or U6385 (N_6385,N_802,N_3028);
nor U6386 (N_6386,N_1052,N_1265);
or U6387 (N_6387,N_4993,N_455);
xor U6388 (N_6388,N_3842,N_3448);
or U6389 (N_6389,N_4676,N_3839);
nand U6390 (N_6390,N_2632,N_4998);
nor U6391 (N_6391,N_966,N_775);
or U6392 (N_6392,N_2188,N_915);
nor U6393 (N_6393,N_722,N_4294);
and U6394 (N_6394,N_1760,N_272);
xnor U6395 (N_6395,N_1449,N_2882);
xnor U6396 (N_6396,N_2915,N_2833);
xor U6397 (N_6397,N_2062,N_1654);
or U6398 (N_6398,N_529,N_2106);
and U6399 (N_6399,N_4844,N_2148);
nor U6400 (N_6400,N_3627,N_4940);
nand U6401 (N_6401,N_1332,N_341);
or U6402 (N_6402,N_2351,N_325);
and U6403 (N_6403,N_4967,N_4398);
xor U6404 (N_6404,N_2889,N_4491);
or U6405 (N_6405,N_2496,N_773);
xor U6406 (N_6406,N_4588,N_2199);
and U6407 (N_6407,N_1027,N_3251);
nor U6408 (N_6408,N_3797,N_4976);
xnor U6409 (N_6409,N_4159,N_256);
nor U6410 (N_6410,N_4675,N_2950);
and U6411 (N_6411,N_985,N_3480);
or U6412 (N_6412,N_3078,N_1984);
or U6413 (N_6413,N_3225,N_1460);
and U6414 (N_6414,N_3010,N_4673);
and U6415 (N_6415,N_4480,N_1985);
or U6416 (N_6416,N_2240,N_2852);
or U6417 (N_6417,N_972,N_1762);
nand U6418 (N_6418,N_1553,N_3652);
xor U6419 (N_6419,N_2693,N_4916);
or U6420 (N_6420,N_2925,N_551);
nor U6421 (N_6421,N_3298,N_1647);
xor U6422 (N_6422,N_3358,N_888);
and U6423 (N_6423,N_1615,N_3016);
or U6424 (N_6424,N_3209,N_308);
nor U6425 (N_6425,N_942,N_1158);
or U6426 (N_6426,N_2194,N_3787);
or U6427 (N_6427,N_669,N_693);
or U6428 (N_6428,N_3772,N_3069);
and U6429 (N_6429,N_86,N_2844);
or U6430 (N_6430,N_2014,N_1003);
or U6431 (N_6431,N_3933,N_4815);
or U6432 (N_6432,N_396,N_954);
nand U6433 (N_6433,N_3699,N_1040);
xnor U6434 (N_6434,N_3788,N_603);
nor U6435 (N_6435,N_4336,N_2124);
xor U6436 (N_6436,N_2845,N_833);
or U6437 (N_6437,N_619,N_1722);
nor U6438 (N_6438,N_3780,N_3040);
nand U6439 (N_6439,N_3687,N_4664);
nand U6440 (N_6440,N_3091,N_116);
xnor U6441 (N_6441,N_4435,N_4482);
and U6442 (N_6442,N_3070,N_489);
or U6443 (N_6443,N_2955,N_4433);
or U6444 (N_6444,N_61,N_1994);
nor U6445 (N_6445,N_1034,N_4958);
nor U6446 (N_6446,N_995,N_2190);
and U6447 (N_6447,N_4630,N_4841);
and U6448 (N_6448,N_1236,N_298);
nor U6449 (N_6449,N_4127,N_1655);
and U6450 (N_6450,N_2116,N_3607);
and U6451 (N_6451,N_2951,N_317);
or U6452 (N_6452,N_627,N_3644);
nand U6453 (N_6453,N_300,N_2861);
nand U6454 (N_6454,N_66,N_4669);
nand U6455 (N_6455,N_2914,N_238);
xor U6456 (N_6456,N_236,N_2928);
nor U6457 (N_6457,N_4283,N_3941);
nor U6458 (N_6458,N_144,N_4625);
nand U6459 (N_6459,N_4052,N_98);
nand U6460 (N_6460,N_4035,N_1474);
or U6461 (N_6461,N_2144,N_4642);
nand U6462 (N_6462,N_3692,N_1466);
nand U6463 (N_6463,N_3878,N_1320);
nand U6464 (N_6464,N_4738,N_1070);
nor U6465 (N_6465,N_2454,N_3951);
and U6466 (N_6466,N_3665,N_2826);
and U6467 (N_6467,N_1402,N_2211);
nand U6468 (N_6468,N_635,N_1597);
nor U6469 (N_6469,N_3178,N_3618);
or U6470 (N_6470,N_2696,N_4270);
xnor U6471 (N_6471,N_4420,N_2041);
or U6472 (N_6472,N_3612,N_436);
and U6473 (N_6473,N_53,N_2359);
xor U6474 (N_6474,N_132,N_2360);
and U6475 (N_6475,N_3864,N_1999);
or U6476 (N_6476,N_259,N_3306);
and U6477 (N_6477,N_2121,N_3385);
nand U6478 (N_6478,N_815,N_3223);
nand U6479 (N_6479,N_1455,N_4849);
nor U6480 (N_6480,N_4704,N_1403);
nor U6481 (N_6481,N_219,N_1895);
xor U6482 (N_6482,N_4512,N_2021);
or U6483 (N_6483,N_4058,N_106);
xor U6484 (N_6484,N_2383,N_579);
or U6485 (N_6485,N_2603,N_101);
and U6486 (N_6486,N_3655,N_4892);
nor U6487 (N_6487,N_678,N_2616);
nand U6488 (N_6488,N_4559,N_1145);
nor U6489 (N_6489,N_1702,N_1792);
xnor U6490 (N_6490,N_1809,N_899);
or U6491 (N_6491,N_4611,N_2829);
and U6492 (N_6492,N_1438,N_1139);
nand U6493 (N_6493,N_444,N_3238);
xnor U6494 (N_6494,N_1649,N_1813);
nand U6495 (N_6495,N_1892,N_1911);
nor U6496 (N_6496,N_2919,N_1934);
xnor U6497 (N_6497,N_215,N_2311);
xor U6498 (N_6498,N_2991,N_3280);
and U6499 (N_6499,N_470,N_3483);
or U6500 (N_6500,N_1203,N_1028);
or U6501 (N_6501,N_2017,N_981);
xor U6502 (N_6502,N_3691,N_1639);
nor U6503 (N_6503,N_4501,N_73);
nor U6504 (N_6504,N_3019,N_4618);
or U6505 (N_6505,N_1926,N_1309);
nand U6506 (N_6506,N_356,N_2853);
nor U6507 (N_6507,N_2277,N_2262);
and U6508 (N_6508,N_4260,N_3397);
and U6509 (N_6509,N_2387,N_4216);
nor U6510 (N_6510,N_2699,N_901);
nand U6511 (N_6511,N_4439,N_1196);
or U6512 (N_6512,N_2698,N_4405);
and U6513 (N_6513,N_3994,N_2573);
and U6514 (N_6514,N_3811,N_2478);
xor U6515 (N_6515,N_1302,N_4418);
nor U6516 (N_6516,N_3517,N_850);
nand U6517 (N_6517,N_2610,N_3683);
and U6518 (N_6518,N_3025,N_3050);
and U6519 (N_6519,N_2645,N_1933);
and U6520 (N_6520,N_3217,N_386);
nor U6521 (N_6521,N_1390,N_4908);
xnor U6522 (N_6522,N_4021,N_1489);
nor U6523 (N_6523,N_4424,N_4213);
nor U6524 (N_6524,N_2501,N_3501);
nor U6525 (N_6525,N_4906,N_21);
or U6526 (N_6526,N_3479,N_2114);
nand U6527 (N_6527,N_3392,N_1644);
or U6528 (N_6528,N_1165,N_1928);
xnor U6529 (N_6529,N_2150,N_3722);
or U6530 (N_6530,N_4221,N_587);
and U6531 (N_6531,N_1325,N_912);
and U6532 (N_6532,N_2372,N_638);
nand U6533 (N_6533,N_1397,N_3126);
and U6534 (N_6534,N_2859,N_670);
nand U6535 (N_6535,N_4508,N_2126);
xnor U6536 (N_6536,N_1940,N_1422);
nand U6537 (N_6537,N_4465,N_887);
nand U6538 (N_6538,N_3926,N_4377);
and U6539 (N_6539,N_254,N_3889);
xnor U6540 (N_6540,N_4779,N_2738);
nor U6541 (N_6541,N_4910,N_574);
nand U6542 (N_6542,N_3890,N_3731);
xnor U6543 (N_6543,N_1808,N_3854);
xor U6544 (N_6544,N_2320,N_406);
nor U6545 (N_6545,N_4944,N_4663);
xor U6546 (N_6546,N_986,N_2029);
or U6547 (N_6547,N_1073,N_3467);
xnor U6548 (N_6548,N_998,N_4086);
xnor U6549 (N_6549,N_3291,N_1986);
nor U6550 (N_6550,N_3954,N_4686);
nand U6551 (N_6551,N_1010,N_454);
xnor U6552 (N_6552,N_2555,N_3203);
and U6553 (N_6553,N_4749,N_85);
xnor U6554 (N_6554,N_2929,N_4601);
xnor U6555 (N_6555,N_1118,N_450);
xor U6556 (N_6556,N_2654,N_4274);
nor U6557 (N_6557,N_3255,N_2182);
nand U6558 (N_6558,N_2973,N_4900);
and U6559 (N_6559,N_1344,N_3891);
nor U6560 (N_6560,N_4472,N_764);
and U6561 (N_6561,N_4184,N_2858);
nor U6562 (N_6562,N_266,N_383);
xnor U6563 (N_6563,N_1846,N_4729);
or U6564 (N_6564,N_1014,N_3082);
and U6565 (N_6565,N_3523,N_4658);
or U6566 (N_6566,N_3767,N_2356);
nand U6567 (N_6567,N_3777,N_4003);
and U6568 (N_6568,N_472,N_4832);
and U6569 (N_6569,N_709,N_991);
and U6570 (N_6570,N_3614,N_598);
nand U6571 (N_6571,N_1528,N_176);
or U6572 (N_6572,N_4972,N_264);
or U6573 (N_6573,N_889,N_4047);
or U6574 (N_6574,N_3739,N_3930);
or U6575 (N_6575,N_4640,N_127);
or U6576 (N_6576,N_2323,N_2446);
nor U6577 (N_6577,N_2650,N_4804);
or U6578 (N_6578,N_2417,N_4488);
nand U6579 (N_6579,N_4203,N_4301);
nand U6580 (N_6580,N_4412,N_633);
or U6581 (N_6581,N_26,N_1362);
nor U6582 (N_6582,N_994,N_3852);
xnor U6583 (N_6583,N_4688,N_4183);
nor U6584 (N_6584,N_910,N_1842);
or U6585 (N_6585,N_920,N_124);
xor U6586 (N_6586,N_3102,N_3366);
xnor U6587 (N_6587,N_4135,N_4404);
nand U6588 (N_6588,N_861,N_471);
or U6589 (N_6589,N_584,N_617);
nor U6590 (N_6590,N_4079,N_452);
nor U6591 (N_6591,N_934,N_4347);
nand U6592 (N_6592,N_225,N_4333);
nand U6593 (N_6593,N_80,N_1205);
and U6594 (N_6594,N_2979,N_4199);
or U6595 (N_6595,N_205,N_1707);
and U6596 (N_6596,N_4396,N_2371);
nor U6597 (N_6597,N_1506,N_2519);
and U6598 (N_6598,N_1151,N_3090);
xor U6599 (N_6599,N_1370,N_1670);
or U6600 (N_6600,N_3648,N_4755);
nand U6601 (N_6601,N_2379,N_1462);
xor U6602 (N_6602,N_2028,N_2350);
nor U6603 (N_6603,N_1839,N_342);
nor U6604 (N_6604,N_4631,N_3595);
and U6605 (N_6605,N_695,N_268);
xor U6606 (N_6606,N_3379,N_3720);
or U6607 (N_6607,N_181,N_3435);
or U6608 (N_6608,N_1176,N_4293);
and U6609 (N_6609,N_1944,N_1433);
and U6610 (N_6610,N_2798,N_360);
nand U6611 (N_6611,N_2664,N_2007);
nor U6612 (N_6612,N_217,N_2719);
or U6613 (N_6613,N_1331,N_247);
nand U6614 (N_6614,N_2672,N_576);
nor U6615 (N_6615,N_3081,N_3205);
and U6616 (N_6616,N_2518,N_482);
or U6617 (N_6617,N_1689,N_3544);
xnor U6618 (N_6618,N_4582,N_463);
xnor U6619 (N_6619,N_347,N_3224);
nor U6620 (N_6620,N_3059,N_1239);
and U6621 (N_6621,N_1163,N_2055);
nor U6622 (N_6622,N_3804,N_3670);
nor U6623 (N_6623,N_1084,N_3918);
and U6624 (N_6624,N_246,N_3474);
nand U6625 (N_6625,N_4623,N_385);
xnor U6626 (N_6626,N_1841,N_191);
nor U6627 (N_6627,N_4609,N_3916);
and U6628 (N_6628,N_1527,N_3214);
nor U6629 (N_6629,N_1144,N_1234);
or U6630 (N_6630,N_1482,N_1444);
and U6631 (N_6631,N_4078,N_3746);
nand U6632 (N_6632,N_634,N_426);
xor U6633 (N_6633,N_193,N_4923);
xor U6634 (N_6634,N_37,N_660);
nor U6635 (N_6635,N_4232,N_713);
nor U6636 (N_6636,N_525,N_3175);
nand U6637 (N_6637,N_392,N_3895);
or U6638 (N_6638,N_459,N_1559);
nor U6639 (N_6639,N_2219,N_3084);
and U6640 (N_6640,N_428,N_332);
nand U6641 (N_6641,N_2168,N_506);
or U6642 (N_6642,N_3514,N_3807);
xnor U6643 (N_6643,N_432,N_1790);
and U6644 (N_6644,N_49,N_2737);
xor U6645 (N_6645,N_3971,N_730);
nand U6646 (N_6646,N_3973,N_4033);
and U6647 (N_6647,N_4284,N_4027);
nand U6648 (N_6648,N_2692,N_368);
nor U6649 (N_6649,N_841,N_1620);
nor U6650 (N_6650,N_1281,N_1475);
xor U6651 (N_6651,N_2839,N_493);
or U6652 (N_6652,N_3294,N_1221);
nor U6653 (N_6653,N_4312,N_3730);
or U6654 (N_6654,N_3986,N_1311);
nand U6655 (N_6655,N_3186,N_4935);
or U6656 (N_6656,N_3782,N_2146);
nor U6657 (N_6657,N_1247,N_3197);
nand U6658 (N_6658,N_3130,N_4425);
nand U6659 (N_6659,N_2272,N_1356);
nor U6660 (N_6660,N_316,N_2448);
nor U6661 (N_6661,N_609,N_2224);
and U6662 (N_6662,N_1510,N_2469);
nor U6663 (N_6663,N_1652,N_375);
xnor U6664 (N_6664,N_1220,N_1029);
or U6665 (N_6665,N_4671,N_4484);
xnor U6666 (N_6666,N_3011,N_3002);
xor U6667 (N_6667,N_72,N_2512);
and U6668 (N_6668,N_4422,N_3952);
and U6669 (N_6669,N_46,N_1255);
nand U6670 (N_6670,N_878,N_309);
and U6671 (N_6671,N_3212,N_3629);
or U6672 (N_6672,N_1427,N_803);
xor U6673 (N_6673,N_2296,N_2537);
and U6674 (N_6674,N_2256,N_2602);
xor U6675 (N_6675,N_1479,N_4130);
and U6676 (N_6676,N_1912,N_2118);
xnor U6677 (N_6677,N_4768,N_4661);
and U6678 (N_6678,N_3034,N_1253);
and U6679 (N_6679,N_2658,N_2724);
nor U6680 (N_6680,N_4010,N_2608);
nor U6681 (N_6681,N_3133,N_3616);
and U6682 (N_6682,N_3743,N_1177);
nor U6683 (N_6683,N_2761,N_1946);
nor U6684 (N_6684,N_747,N_2189);
and U6685 (N_6685,N_2220,N_798);
nor U6686 (N_6686,N_505,N_1369);
xnor U6687 (N_6687,N_2716,N_4929);
nor U6688 (N_6688,N_1810,N_2111);
or U6689 (N_6689,N_1969,N_3044);
and U6690 (N_6690,N_446,N_1081);
or U6691 (N_6691,N_3896,N_4145);
and U6692 (N_6692,N_2606,N_4375);
nor U6693 (N_6693,N_3460,N_1237);
nor U6694 (N_6694,N_2718,N_184);
and U6695 (N_6695,N_4009,N_4781);
nand U6696 (N_6696,N_2104,N_4506);
xnor U6697 (N_6697,N_637,N_4045);
nand U6698 (N_6698,N_849,N_1244);
and U6699 (N_6699,N_3491,N_3361);
and U6700 (N_6700,N_1751,N_349);
and U6701 (N_6701,N_2550,N_3639);
nor U6702 (N_6702,N_1106,N_1754);
nand U6703 (N_6703,N_563,N_3171);
xnor U6704 (N_6704,N_2342,N_739);
xnor U6705 (N_6705,N_2053,N_857);
or U6706 (N_6706,N_3329,N_963);
and U6707 (N_6707,N_1853,N_1645);
nand U6708 (N_6708,N_1742,N_2032);
nor U6709 (N_6709,N_3442,N_4511);
or U6710 (N_6710,N_1180,N_3252);
nor U6711 (N_6711,N_3348,N_591);
nand U6712 (N_6712,N_3233,N_2178);
xnor U6713 (N_6713,N_3260,N_4653);
and U6714 (N_6714,N_344,N_1184);
and U6715 (N_6715,N_2044,N_928);
nand U6716 (N_6716,N_4720,N_4721);
nand U6717 (N_6717,N_4278,N_3546);
xor U6718 (N_6718,N_1913,N_823);
xor U6719 (N_6719,N_1101,N_2282);
nand U6720 (N_6720,N_527,N_1013);
xor U6721 (N_6721,N_3748,N_1263);
and U6722 (N_6722,N_485,N_893);
and U6723 (N_6723,N_1242,N_3576);
xnor U6724 (N_6724,N_776,N_2659);
nand U6725 (N_6725,N_1526,N_927);
and U6726 (N_6726,N_2271,N_1505);
nand U6727 (N_6727,N_3012,N_880);
and U6728 (N_6728,N_3641,N_2491);
or U6729 (N_6729,N_720,N_218);
nand U6730 (N_6730,N_623,N_1330);
and U6731 (N_6731,N_2462,N_1345);
or U6732 (N_6732,N_2944,N_4503);
nand U6733 (N_6733,N_2980,N_3773);
nand U6734 (N_6734,N_1400,N_2065);
nor U6735 (N_6735,N_4610,N_2967);
or U6736 (N_6736,N_1824,N_4257);
nor U6737 (N_6737,N_2800,N_3478);
xor U6738 (N_6738,N_4262,N_2592);
or U6739 (N_6739,N_4530,N_2743);
nand U6740 (N_6740,N_1855,N_1421);
or U6741 (N_6741,N_1283,N_1648);
nand U6742 (N_6742,N_2230,N_3240);
nand U6743 (N_6743,N_3461,N_417);
nand U6744 (N_6744,N_4171,N_4523);
nand U6745 (N_6745,N_904,N_1605);
nor U6746 (N_6746,N_4335,N_4553);
nor U6747 (N_6747,N_2056,N_2172);
xor U6748 (N_6748,N_2306,N_1524);
and U6749 (N_6749,N_1758,N_2039);
nand U6750 (N_6750,N_2875,N_34);
xor U6751 (N_6751,N_273,N_2628);
and U6752 (N_6752,N_3108,N_4603);
or U6753 (N_6753,N_1365,N_3383);
xor U6754 (N_6754,N_2420,N_949);
nor U6755 (N_6755,N_1478,N_1319);
and U6756 (N_6756,N_583,N_4410);
xor U6757 (N_6757,N_3795,N_4099);
nor U6758 (N_6758,N_882,N_4532);
xor U6759 (N_6759,N_1304,N_4515);
and U6760 (N_6760,N_2821,N_3557);
and U6761 (N_6761,N_3562,N_3455);
xnor U6762 (N_6762,N_4594,N_60);
or U6763 (N_6763,N_4367,N_4407);
or U6764 (N_6764,N_2355,N_1501);
nor U6765 (N_6765,N_331,N_1277);
or U6766 (N_6766,N_1924,N_3803);
or U6767 (N_6767,N_1295,N_556);
xor U6768 (N_6768,N_4403,N_2204);
or U6769 (N_6769,N_3137,N_4514);
and U6770 (N_6770,N_3055,N_2022);
or U6771 (N_6771,N_668,N_2251);
nand U6772 (N_6772,N_1564,N_170);
or U6773 (N_6773,N_2840,N_4985);
xnor U6774 (N_6774,N_513,N_250);
nand U6775 (N_6775,N_4495,N_2912);
xor U6776 (N_6776,N_1518,N_4122);
nor U6777 (N_6777,N_2357,N_3729);
nor U6778 (N_6778,N_939,N_3456);
nand U6779 (N_6779,N_2317,N_2326);
or U6780 (N_6780,N_2102,N_3868);
and U6781 (N_6781,N_4684,N_2218);
nand U6782 (N_6782,N_542,N_1417);
and U6783 (N_6783,N_978,N_1776);
nand U6784 (N_6784,N_1006,N_1068);
or U6785 (N_6785,N_3420,N_1436);
or U6786 (N_6786,N_2215,N_2597);
and U6787 (N_6787,N_4607,N_1595);
xnor U6788 (N_6788,N_2101,N_466);
nor U6789 (N_6789,N_4727,N_3148);
nor U6790 (N_6790,N_1050,N_2245);
nor U6791 (N_6791,N_3060,N_2205);
and U6792 (N_6792,N_629,N_3619);
nand U6793 (N_6793,N_1593,N_224);
nand U6794 (N_6794,N_1786,N_800);
xnor U6795 (N_6795,N_3465,N_424);
nand U6796 (N_6796,N_4155,N_4851);
and U6797 (N_6797,N_2348,N_4328);
xor U6798 (N_6798,N_3560,N_1598);
and U6799 (N_6799,N_498,N_2599);
nor U6800 (N_6800,N_351,N_1352);
xnor U6801 (N_6801,N_3418,N_1110);
or U6802 (N_6802,N_4874,N_4444);
nor U6803 (N_6803,N_2416,N_3900);
nor U6804 (N_6804,N_782,N_682);
xnor U6805 (N_6805,N_2997,N_4360);
nand U6806 (N_6806,N_2943,N_104);
and U6807 (N_6807,N_2289,N_2612);
or U6808 (N_6808,N_1012,N_4349);
and U6809 (N_6809,N_100,N_1200);
and U6810 (N_6810,N_1756,N_1007);
or U6811 (N_6811,N_467,N_4746);
nand U6812 (N_6812,N_677,N_2345);
nand U6813 (N_6813,N_2389,N_2933);
or U6814 (N_6814,N_4902,N_1416);
or U6815 (N_6815,N_2113,N_1019);
or U6816 (N_6816,N_3776,N_3559);
and U6817 (N_6817,N_330,N_4165);
nor U6818 (N_6818,N_2749,N_4535);
or U6819 (N_6819,N_946,N_4890);
and U6820 (N_6820,N_3424,N_544);
and U6821 (N_6821,N_2522,N_481);
nor U6822 (N_6822,N_3023,N_1703);
nand U6823 (N_6823,N_3840,N_2063);
and U6824 (N_6824,N_123,N_4831);
and U6825 (N_6825,N_2906,N_1591);
xnor U6826 (N_6826,N_3542,N_2994);
and U6827 (N_6827,N_1291,N_4395);
nor U6828 (N_6828,N_3073,N_1232);
nand U6829 (N_6829,N_4667,N_521);
and U6830 (N_6830,N_2781,N_387);
xor U6831 (N_6831,N_701,N_4941);
nand U6832 (N_6832,N_1830,N_3368);
xnor U6833 (N_6833,N_671,N_235);
and U6834 (N_6834,N_2058,N_114);
or U6835 (N_6835,N_1868,N_2020);
xnor U6836 (N_6836,N_2415,N_2145);
or U6837 (N_6837,N_1566,N_1252);
nor U6838 (N_6838,N_3018,N_1785);
xor U6839 (N_6839,N_1539,N_1636);
nor U6840 (N_6840,N_808,N_1571);
or U6841 (N_6841,N_2142,N_4830);
and U6842 (N_6842,N_4473,N_1949);
nor U6843 (N_6843,N_3362,N_4273);
xnor U6844 (N_6844,N_2413,N_4657);
nor U6845 (N_6845,N_2061,N_230);
and U6846 (N_6846,N_239,N_2891);
or U6847 (N_6847,N_1004,N_3342);
nor U6848 (N_6848,N_4717,N_3599);
or U6849 (N_6849,N_1044,N_2304);
or U6850 (N_6850,N_1183,N_2140);
nor U6851 (N_6851,N_2816,N_4752);
or U6852 (N_6852,N_4175,N_2312);
nor U6853 (N_6853,N_2759,N_3331);
xor U6854 (N_6854,N_2942,N_4820);
nand U6855 (N_6855,N_1231,N_754);
xor U6856 (N_6856,N_1454,N_3013);
and U6857 (N_6857,N_854,N_1602);
nand U6858 (N_6858,N_1676,N_4366);
or U6859 (N_6859,N_3177,N_4246);
xnor U6860 (N_6860,N_812,N_555);
nand U6861 (N_6861,N_4857,N_2754);
nor U6862 (N_6862,N_232,N_3940);
nor U6863 (N_6863,N_1675,N_1193);
nor U6864 (N_6864,N_3053,N_2989);
or U6865 (N_6865,N_1642,N_1060);
nand U6866 (N_6866,N_606,N_2019);
xnor U6867 (N_6867,N_1837,N_3254);
or U6868 (N_6868,N_2975,N_1079);
nor U6869 (N_6869,N_673,N_2517);
nand U6870 (N_6870,N_2815,N_1589);
nor U6871 (N_6871,N_2461,N_1289);
nor U6872 (N_6872,N_196,N_704);
nor U6873 (N_6873,N_3352,N_989);
nor U6874 (N_6874,N_149,N_1927);
nor U6875 (N_6875,N_1780,N_2793);
nor U6876 (N_6876,N_2026,N_4803);
nor U6877 (N_6877,N_364,N_552);
nand U6878 (N_6878,N_1613,N_4362);
xor U6879 (N_6879,N_779,N_2544);
or U6880 (N_6880,N_3968,N_2864);
nand U6881 (N_6881,N_1697,N_1049);
nor U6882 (N_6882,N_1857,N_4774);
and U6883 (N_6883,N_2586,N_139);
xor U6884 (N_6884,N_3711,N_3004);
or U6885 (N_6885,N_1293,N_4248);
and U6886 (N_6886,N_2200,N_2579);
xor U6887 (N_6887,N_1150,N_4871);
xnor U6888 (N_6888,N_4842,N_3590);
xor U6889 (N_6889,N_2808,N_3915);
nor U6890 (N_6890,N_2255,N_405);
nor U6891 (N_6891,N_2384,N_644);
and U6892 (N_6892,N_2750,N_1856);
xnor U6893 (N_6893,N_1801,N_4836);
or U6894 (N_6894,N_1669,N_3841);
xor U6895 (N_6895,N_1929,N_1545);
and U6896 (N_6896,N_1882,N_3666);
and U6897 (N_6897,N_1334,N_714);
and U6898 (N_6898,N_4868,N_2401);
nor U6899 (N_6899,N_2487,N_2060);
xor U6900 (N_6900,N_982,N_1560);
and U6901 (N_6901,N_4978,N_262);
xor U6902 (N_6902,N_1578,N_4795);
nor U6903 (N_6903,N_923,N_3321);
and U6904 (N_6904,N_4650,N_597);
xor U6905 (N_6905,N_4324,N_4421);
and U6906 (N_6906,N_1376,N_3944);
or U6907 (N_6907,N_924,N_4237);
xnor U6908 (N_6908,N_3190,N_3316);
and U6909 (N_6909,N_4979,N_4989);
nand U6910 (N_6910,N_2246,N_3216);
or U6911 (N_6911,N_4873,N_2000);
xor U6912 (N_6912,N_2721,N_3658);
xnor U6913 (N_6913,N_1420,N_2091);
nand U6914 (N_6914,N_4600,N_4997);
nor U6915 (N_6915,N_2089,N_2176);
or U6916 (N_6916,N_3704,N_1533);
or U6917 (N_6917,N_3887,N_2896);
or U6918 (N_6918,N_4388,N_1194);
nand U6919 (N_6919,N_4189,N_208);
and U6920 (N_6920,N_4659,N_4043);
nor U6921 (N_6921,N_2686,N_3043);
nand U6922 (N_6922,N_1254,N_559);
nand U6923 (N_6923,N_51,N_3008);
and U6924 (N_6924,N_4193,N_3447);
or U6925 (N_6925,N_4436,N_1667);
and U6926 (N_6926,N_1759,N_1396);
xnor U6927 (N_6927,N_155,N_3998);
xor U6928 (N_6928,N_4974,N_3927);
nor U6929 (N_6929,N_2427,N_4378);
and U6930 (N_6930,N_1523,N_2368);
nand U6931 (N_6931,N_851,N_1228);
xnor U6932 (N_6932,N_2231,N_84);
nor U6933 (N_6933,N_4735,N_69);
nand U6934 (N_6934,N_3110,N_2309);
or U6935 (N_6935,N_4778,N_2615);
nand U6936 (N_6936,N_614,N_1457);
nor U6937 (N_6937,N_277,N_1190);
nor U6938 (N_6938,N_1646,N_4072);
xnor U6939 (N_6939,N_3921,N_1126);
nand U6940 (N_6940,N_1872,N_4374);
xnor U6941 (N_6941,N_4947,N_244);
and U6942 (N_6942,N_1124,N_630);
nand U6943 (N_6943,N_4896,N_2184);
nand U6944 (N_6944,N_2886,N_414);
and U6945 (N_6945,N_1216,N_41);
nand U6946 (N_6946,N_2881,N_4044);
nand U6947 (N_6947,N_1951,N_3763);
and U6948 (N_6948,N_1978,N_3468);
or U6949 (N_6949,N_3813,N_4765);
xnor U6950 (N_6950,N_4118,N_1367);
nor U6951 (N_6951,N_3580,N_1377);
xor U6952 (N_6952,N_3336,N_1682);
nand U6953 (N_6953,N_1546,N_4702);
or U6954 (N_6954,N_4767,N_2558);
or U6955 (N_6955,N_2438,N_4517);
nor U6956 (N_6956,N_1226,N_4207);
and U6957 (N_6957,N_3554,N_448);
and U6958 (N_6958,N_4022,N_2050);
and U6959 (N_6959,N_4330,N_4920);
nor U6960 (N_6960,N_4701,N_1705);
nand U6961 (N_6961,N_1565,N_1550);
or U6962 (N_6962,N_2024,N_2283);
nand U6963 (N_6963,N_1389,N_1093);
nor U6964 (N_6964,N_1910,N_4519);
or U6965 (N_6965,N_2902,N_2545);
nor U6966 (N_6966,N_2180,N_2609);
and U6967 (N_6967,N_438,N_4726);
nand U6968 (N_6968,N_111,N_4348);
and U6969 (N_6969,N_3065,N_4905);
nor U6970 (N_6970,N_1542,N_2165);
and U6971 (N_6971,N_2258,N_3844);
nor U6972 (N_6972,N_2344,N_4018);
xnor U6973 (N_6973,N_153,N_62);
xnor U6974 (N_6974,N_3049,N_4074);
nor U6975 (N_6975,N_3563,N_1793);
or U6976 (N_6976,N_659,N_3277);
xor U6977 (N_6977,N_2147,N_4826);
nand U6978 (N_6978,N_3838,N_2618);
and U6979 (N_6979,N_4464,N_3246);
xnor U6980 (N_6980,N_1227,N_3752);
nor U6981 (N_6981,N_4546,N_486);
nand U6982 (N_6982,N_726,N_4371);
xor U6983 (N_6983,N_3495,N_3015);
nand U6984 (N_6984,N_4709,N_2159);
xor U6985 (N_6985,N_3253,N_710);
and U6986 (N_6986,N_3372,N_4105);
xnor U6987 (N_6987,N_3139,N_2421);
nand U6988 (N_6988,N_4539,N_2542);
nor U6989 (N_6989,N_4069,N_17);
or U6990 (N_6990,N_2649,N_1970);
nand U6991 (N_6991,N_2837,N_4195);
xor U6992 (N_6992,N_1532,N_2045);
or U6993 (N_6993,N_3001,N_1728);
or U6994 (N_6994,N_2768,N_2110);
xnor U6995 (N_6995,N_157,N_1611);
and U6996 (N_6996,N_1424,N_1932);
and U6997 (N_6997,N_3762,N_122);
nor U6998 (N_6998,N_3833,N_2455);
and U6999 (N_6999,N_202,N_1168);
nand U7000 (N_7000,N_3700,N_2198);
nand U7001 (N_7001,N_3071,N_2298);
and U7002 (N_7002,N_2414,N_2392);
nor U7003 (N_7003,N_1659,N_1903);
xor U7004 (N_7004,N_3105,N_1653);
xnor U7005 (N_7005,N_1443,N_1529);
nand U7006 (N_7006,N_449,N_3454);
nor U7007 (N_7007,N_2068,N_4986);
nor U7008 (N_7008,N_3816,N_2232);
and U7009 (N_7009,N_4808,N_610);
xor U7010 (N_7010,N_1720,N_2763);
nor U7011 (N_7011,N_4249,N_830);
and U7012 (N_7012,N_1626,N_4855);
nor U7013 (N_7013,N_4309,N_1819);
and U7014 (N_7014,N_2799,N_3650);
xor U7015 (N_7015,N_4459,N_1002);
and U7016 (N_7016,N_1888,N_2025);
and U7017 (N_7017,N_3678,N_4040);
and U7018 (N_7018,N_2922,N_369);
and U7019 (N_7019,N_582,N_2828);
nor U7020 (N_7020,N_4792,N_3885);
nor U7021 (N_7021,N_4744,N_2173);
xor U7022 (N_7022,N_2339,N_154);
and U7023 (N_7023,N_65,N_3713);
nand U7024 (N_7024,N_2009,N_2083);
xor U7025 (N_7025,N_1445,N_1724);
nand U7026 (N_7026,N_3609,N_3515);
xnor U7027 (N_7027,N_4244,N_1772);
xnor U7028 (N_7028,N_1146,N_3198);
or U7029 (N_7029,N_4652,N_134);
or U7030 (N_7030,N_2208,N_3187);
nand U7031 (N_7031,N_1279,N_1921);
or U7032 (N_7032,N_198,N_766);
nand U7033 (N_7033,N_1026,N_4654);
and U7034 (N_7034,N_1375,N_439);
and U7035 (N_7035,N_3103,N_3579);
and U7036 (N_7036,N_3584,N_1656);
nor U7037 (N_7037,N_2684,N_4843);
xor U7038 (N_7038,N_4204,N_203);
nand U7039 (N_7039,N_4660,N_1224);
xnor U7040 (N_7040,N_126,N_3360);
and U7041 (N_7041,N_1069,N_4936);
nor U7042 (N_7042,N_2411,N_3516);
and U7043 (N_7043,N_4121,N_3635);
nand U7044 (N_7044,N_2851,N_1787);
xor U7045 (N_7045,N_4656,N_1804);
and U7046 (N_7046,N_3792,N_2484);
and U7047 (N_7047,N_2812,N_2191);
and U7048 (N_7048,N_4098,N_2662);
nor U7049 (N_7049,N_809,N_3510);
nand U7050 (N_7050,N_1067,N_3999);
nand U7051 (N_7051,N_1419,N_4576);
nor U7052 (N_7052,N_4672,N_4705);
nor U7053 (N_7053,N_3494,N_2918);
xor U7054 (N_7054,N_4138,N_1699);
nor U7055 (N_7055,N_3476,N_516);
nor U7056 (N_7056,N_3269,N_524);
and U7057 (N_7057,N_63,N_1902);
or U7058 (N_7058,N_2897,N_1492);
nand U7059 (N_7059,N_3444,N_4524);
xnor U7060 (N_7060,N_2233,N_3375);
and U7061 (N_7061,N_2084,N_3547);
nand U7062 (N_7062,N_201,N_4537);
or U7063 (N_7063,N_2003,N_4606);
nor U7064 (N_7064,N_240,N_761);
and U7065 (N_7065,N_2715,N_3199);
nand U7066 (N_7066,N_393,N_2879);
xor U7067 (N_7067,N_1993,N_607);
nor U7068 (N_7068,N_1690,N_3992);
nor U7069 (N_7069,N_538,N_1854);
xor U7070 (N_7070,N_4933,N_1920);
or U7071 (N_7071,N_1054,N_4622);
nor U7072 (N_7072,N_3443,N_4454);
nand U7073 (N_7073,N_5,N_479);
and U7074 (N_7074,N_2795,N_3751);
xor U7075 (N_7075,N_2739,N_2117);
xor U7076 (N_7076,N_9,N_2757);
xor U7077 (N_7077,N_3712,N_3706);
or U7078 (N_7078,N_4185,N_343);
nor U7079 (N_7079,N_2604,N_2572);
or U7080 (N_7080,N_4866,N_1572);
xor U7081 (N_7081,N_3184,N_4434);
nor U7082 (N_7082,N_4960,N_280);
nand U7083 (N_7083,N_125,N_1337);
nor U7084 (N_7084,N_2728,N_4355);
and U7085 (N_7085,N_2481,N_2196);
nor U7086 (N_7086,N_4116,N_2978);
xnor U7087 (N_7087,N_4002,N_3768);
xnor U7088 (N_7088,N_1206,N_2265);
xnor U7089 (N_7089,N_3388,N_4141);
nand U7090 (N_7090,N_1235,N_2267);
nand U7091 (N_7091,N_4463,N_2657);
nor U7092 (N_7092,N_2437,N_1752);
and U7093 (N_7093,N_50,N_3967);
xor U7094 (N_7094,N_1738,N_3799);
and U7095 (N_7095,N_354,N_2687);
xor U7096 (N_7096,N_4090,N_3809);
xnor U7097 (N_7097,N_3296,N_195);
nand U7098 (N_7098,N_4413,N_1238);
xnor U7099 (N_7099,N_2784,N_2408);
nand U7100 (N_7100,N_3662,N_2250);
nand U7101 (N_7101,N_2702,N_2700);
nor U7102 (N_7102,N_712,N_1950);
nand U7103 (N_7103,N_4763,N_4187);
or U7104 (N_7104,N_3810,N_3241);
nand U7105 (N_7105,N_2520,N_528);
or U7106 (N_7106,N_1584,N_2203);
or U7107 (N_7107,N_3741,N_4585);
and U7108 (N_7108,N_4734,N_567);
nor U7109 (N_7109,N_2301,N_3095);
and U7110 (N_7110,N_4496,N_3458);
nor U7111 (N_7111,N_3218,N_859);
nor U7112 (N_7112,N_2287,N_2773);
nor U7113 (N_7113,N_2254,N_2008);
xnor U7114 (N_7114,N_3427,N_699);
nand U7115 (N_7115,N_130,N_1366);
and U7116 (N_7116,N_1025,N_2587);
xnor U7117 (N_7117,N_4891,N_1635);
xor U7118 (N_7118,N_4574,N_3498);
nand U7119 (N_7119,N_1606,N_1540);
nor U7120 (N_7120,N_4617,N_4579);
and U7121 (N_7121,N_4570,N_2349);
nor U7122 (N_7122,N_4223,N_3313);
and U7123 (N_7123,N_4286,N_1881);
or U7124 (N_7124,N_4828,N_293);
nand U7125 (N_7125,N_1974,N_3482);
nor U7126 (N_7126,N_594,N_174);
and U7127 (N_7127,N_729,N_1161);
and U7128 (N_7128,N_1099,N_83);
nor U7129 (N_7129,N_1768,N_2676);
nor U7130 (N_7130,N_1619,N_4544);
and U7131 (N_7131,N_2802,N_2151);
nand U7132 (N_7132,N_4888,N_2595);
nand U7133 (N_7133,N_1746,N_1618);
nand U7134 (N_7134,N_3154,N_2830);
xnor U7135 (N_7135,N_2088,N_3789);
xnor U7136 (N_7136,N_212,N_1020);
nand U7137 (N_7137,N_2445,N_4966);
nand U7138 (N_7138,N_1372,N_492);
nor U7139 (N_7139,N_4485,N_2605);
or U7140 (N_7140,N_3610,N_4877);
or U7141 (N_7141,N_4784,N_1800);
nor U7142 (N_7142,N_3007,N_1383);
and U7143 (N_7143,N_4147,N_2741);
nor U7144 (N_7144,N_626,N_3745);
xnor U7145 (N_7145,N_1136,N_4048);
nand U7146 (N_7146,N_2149,N_4202);
nand U7147 (N_7147,N_2948,N_4016);
xor U7148 (N_7148,N_2346,N_3301);
and U7149 (N_7149,N_2966,N_1294);
nor U7150 (N_7150,N_2164,N_796);
xor U7151 (N_7151,N_2412,N_4208);
nor U7152 (N_7152,N_4760,N_2963);
nand U7153 (N_7153,N_2624,N_733);
nand U7154 (N_7154,N_2801,N_2132);
xnor U7155 (N_7155,N_3531,N_3848);
xnor U7156 (N_7156,N_4379,N_568);
and U7157 (N_7157,N_3407,N_4101);
nor U7158 (N_7158,N_3350,N_22);
or U7159 (N_7159,N_3911,N_1607);
or U7160 (N_7160,N_728,N_1763);
and U7161 (N_7161,N_1361,N_4949);
xor U7162 (N_7162,N_1323,N_4341);
and U7163 (N_7163,N_3846,N_2109);
xnor U7164 (N_7164,N_4680,N_409);
and U7165 (N_7165,N_4241,N_2964);
nor U7166 (N_7166,N_3668,N_2275);
xnor U7167 (N_7167,N_150,N_255);
or U7168 (N_7168,N_1192,N_3109);
nor U7169 (N_7169,N_2059,N_3866);
or U7170 (N_7170,N_3470,N_468);
and U7171 (N_7171,N_1043,N_2972);
or U7172 (N_7172,N_4994,N_1031);
and U7173 (N_7173,N_4234,N_162);
nand U7174 (N_7174,N_1627,N_866);
or U7175 (N_7175,N_2671,N_3279);
or U7176 (N_7176,N_2186,N_3393);
xor U7177 (N_7177,N_4049,N_3275);
nand U7178 (N_7178,N_4160,N_4568);
nor U7179 (N_7179,N_2212,N_2733);
nand U7180 (N_7180,N_530,N_2210);
and U7181 (N_7181,N_1743,N_3566);
xnor U7182 (N_7182,N_3213,N_3581);
and U7183 (N_7183,N_3529,N_2797);
nand U7184 (N_7184,N_3149,N_1741);
nor U7185 (N_7185,N_1966,N_1805);
nand U7186 (N_7186,N_2153,N_2092);
or U7187 (N_7187,N_2338,N_3335);
and U7188 (N_7188,N_1102,N_87);
nand U7189 (N_7189,N_4304,N_1166);
nand U7190 (N_7190,N_2583,N_2927);
xor U7191 (N_7191,N_4791,N_1862);
or U7192 (N_7192,N_3628,N_3437);
or U7193 (N_7193,N_2499,N_500);
nand U7194 (N_7194,N_4205,N_953);
and U7195 (N_7195,N_78,N_4942);
xnor U7196 (N_7196,N_3827,N_260);
xor U7197 (N_7197,N_1640,N_2490);
nor U7198 (N_7198,N_3030,N_2174);
nor U7199 (N_7199,N_1113,N_2651);
nand U7200 (N_7200,N_252,N_3250);
nand U7201 (N_7201,N_824,N_1904);
and U7202 (N_7202,N_3898,N_2746);
nor U7203 (N_7203,N_2447,N_399);
nand U7204 (N_7204,N_2813,N_2846);
or U7205 (N_7205,N_4898,N_296);
xnor U7206 (N_7206,N_4557,N_3325);
nor U7207 (N_7207,N_2228,N_2690);
or U7208 (N_7208,N_2435,N_855);
or U7209 (N_7209,N_1538,N_2640);
or U7210 (N_7210,N_4999,N_4838);
nand U7211 (N_7211,N_2243,N_1577);
nand U7212 (N_7212,N_3038,N_4399);
nor U7213 (N_7213,N_1202,N_3905);
nor U7214 (N_7214,N_3112,N_3991);
or U7215 (N_7215,N_1643,N_4383);
or U7216 (N_7216,N_3821,N_3894);
nor U7217 (N_7217,N_3265,N_2166);
nor U7218 (N_7218,N_1075,N_1432);
and U7219 (N_7219,N_348,N_4945);
xor U7220 (N_7220,N_4643,N_2239);
or U7221 (N_7221,N_2661,N_4683);
nor U7222 (N_7222,N_2485,N_3733);
or U7223 (N_7223,N_2732,N_221);
nor U7224 (N_7224,N_1878,N_3660);
nor U7225 (N_7225,N_4627,N_8);
nor U7226 (N_7226,N_3143,N_2984);
or U7227 (N_7227,N_2193,N_391);
xor U7228 (N_7228,N_1222,N_698);
nor U7229 (N_7229,N_2621,N_1975);
or U7230 (N_7230,N_3703,N_1008);
nor U7231 (N_7231,N_4950,N_1275);
xnor U7232 (N_7232,N_2523,N_4595);
nor U7233 (N_7233,N_2701,N_3158);
or U7234 (N_7234,N_2620,N_3006);
nor U7235 (N_7235,N_2945,N_3935);
nor U7236 (N_7236,N_3196,N_3428);
nand U7237 (N_7237,N_1775,N_908);
nand U7238 (N_7238,N_3570,N_222);
nor U7239 (N_7239,N_4813,N_1116);
xor U7240 (N_7240,N_4805,N_1548);
and U7241 (N_7241,N_3750,N_3605);
xnor U7242 (N_7242,N_3234,N_1897);
nor U7243 (N_7243,N_4115,N_4369);
xnor U7244 (N_7244,N_2268,N_245);
xor U7245 (N_7245,N_42,N_4276);
or U7246 (N_7246,N_3871,N_3111);
nand U7247 (N_7247,N_1497,N_1230);
and U7248 (N_7248,N_4080,N_2756);
nor U7249 (N_7249,N_4715,N_2665);
nand U7250 (N_7250,N_2729,N_3749);
or U7251 (N_7251,N_1961,N_2549);
xor U7252 (N_7252,N_4818,N_3384);
nor U7253 (N_7253,N_1261,N_3963);
or U7254 (N_7254,N_96,N_4104);
nor U7255 (N_7255,N_2783,N_3339);
xor U7256 (N_7256,N_1058,N_2974);
and U7257 (N_7257,N_4567,N_1582);
and U7258 (N_7258,N_306,N_410);
nand U7259 (N_7259,N_4885,N_4914);
and U7260 (N_7260,N_3592,N_3144);
xor U7261 (N_7261,N_2390,N_4409);
xor U7262 (N_7262,N_1755,N_965);
xnor U7263 (N_7263,N_3367,N_1219);
nand U7264 (N_7264,N_988,N_3398);
or U7265 (N_7265,N_3754,N_3211);
nand U7266 (N_7266,N_1284,N_3818);
nor U7267 (N_7267,N_1276,N_4951);
or U7268 (N_7268,N_3714,N_3760);
nand U7269 (N_7269,N_1410,N_573);
xnor U7270 (N_7270,N_1783,N_2543);
nor U7271 (N_7271,N_1871,N_4011);
or U7272 (N_7272,N_1086,N_3796);
and U7273 (N_7273,N_4859,N_3106);
nand U7274 (N_7274,N_253,N_837);
and U7275 (N_7275,N_1588,N_281);
and U7276 (N_7276,N_4731,N_3257);
or U7277 (N_7277,N_2095,N_197);
or U7278 (N_7278,N_95,N_3459);
and U7279 (N_7279,N_1483,N_748);
nor U7280 (N_7280,N_2867,N_846);
xor U7281 (N_7281,N_461,N_4869);
or U7282 (N_7282,N_3785,N_4112);
or U7283 (N_7283,N_1147,N_2744);
nand U7284 (N_7284,N_763,N_337);
and U7285 (N_7285,N_3146,N_1472);
or U7286 (N_7286,N_4358,N_696);
or U7287 (N_7287,N_82,N_1757);
and U7288 (N_7288,N_4777,N_4392);
and U7289 (N_7289,N_2450,N_4285);
and U7290 (N_7290,N_1807,N_4964);
xor U7291 (N_7291,N_112,N_2209);
or U7292 (N_7292,N_993,N_2775);
or U7293 (N_7293,N_1469,N_4837);
nand U7294 (N_7294,N_2764,N_2252);
or U7295 (N_7295,N_3718,N_742);
nor U7296 (N_7296,N_2470,N_758);
xor U7297 (N_7297,N_589,N_1141);
nor U7298 (N_7298,N_3883,N_3923);
nor U7299 (N_7299,N_1908,N_4747);
nand U7300 (N_7300,N_429,N_3593);
or U7301 (N_7301,N_4761,N_2202);
nor U7302 (N_7302,N_4060,N_3615);
nor U7303 (N_7303,N_785,N_1534);
or U7304 (N_7304,N_23,N_44);
nand U7305 (N_7305,N_3808,N_727);
nor U7306 (N_7306,N_1173,N_2015);
or U7307 (N_7307,N_1672,N_3937);
and U7308 (N_7308,N_1883,N_2419);
and U7309 (N_7309,N_4490,N_1733);
or U7310 (N_7310,N_546,N_3877);
or U7311 (N_7311,N_3317,N_532);
nand U7312 (N_7312,N_1071,N_676);
nor U7313 (N_7313,N_1340,N_2128);
or U7314 (N_7314,N_4925,N_1869);
nand U7315 (N_7315,N_2138,N_662);
and U7316 (N_7316,N_12,N_4163);
xor U7317 (N_7317,N_3548,N_4988);
or U7318 (N_7318,N_2169,N_2425);
xor U7319 (N_7319,N_3229,N_566);
nand U7320 (N_7320,N_868,N_2970);
nand U7321 (N_7321,N_3500,N_358);
and U7322 (N_7322,N_2962,N_1077);
or U7323 (N_7323,N_4096,N_4751);
nor U7324 (N_7324,N_3765,N_2051);
nand U7325 (N_7325,N_4139,N_1197);
and U7326 (N_7326,N_4536,N_940);
or U7327 (N_7327,N_3230,N_3349);
nor U7328 (N_7328,N_1681,N_423);
nand U7329 (N_7329,N_2899,N_1996);
nand U7330 (N_7330,N_2170,N_1858);
nand U7331 (N_7331,N_2330,N_4736);
xor U7332 (N_7332,N_3503,N_4772);
and U7333 (N_7333,N_3586,N_3783);
or U7334 (N_7334,N_1953,N_3997);
nor U7335 (N_7335,N_2493,N_3396);
or U7336 (N_7336,N_3484,N_1048);
or U7337 (N_7337,N_690,N_3270);
and U7338 (N_7338,N_336,N_1657);
nor U7339 (N_7339,N_1507,N_2307);
xor U7340 (N_7340,N_2841,N_3445);
or U7341 (N_7341,N_2935,N_2622);
nand U7342 (N_7342,N_1326,N_4174);
nand U7343 (N_7343,N_1262,N_1108);
nor U7344 (N_7344,N_2141,N_3207);
or U7345 (N_7345,N_3286,N_3287);
nand U7346 (N_7346,N_491,N_3115);
xnor U7347 (N_7347,N_3892,N_3893);
nand U7348 (N_7348,N_68,N_3707);
or U7349 (N_7349,N_4718,N_2673);
or U7350 (N_7350,N_4520,N_4954);
and U7351 (N_7351,N_4150,N_1423);
xor U7352 (N_7352,N_1877,N_2663);
nor U7353 (N_7353,N_3308,N_407);
or U7354 (N_7354,N_1867,N_3227);
nor U7355 (N_7355,N_3248,N_879);
xnor U7356 (N_7356,N_778,N_4800);
xor U7357 (N_7357,N_4314,N_548);
xnor U7358 (N_7358,N_1581,N_3416);
nand U7359 (N_7359,N_4442,N_869);
xnor U7360 (N_7360,N_335,N_1544);
or U7361 (N_7361,N_4555,N_1341);
nor U7362 (N_7362,N_2468,N_3806);
xor U7363 (N_7363,N_873,N_3098);
nand U7364 (N_7364,N_2010,N_845);
or U7365 (N_7365,N_3147,N_2880);
xnor U7366 (N_7366,N_1278,N_4996);
or U7367 (N_7367,N_3064,N_2571);
nor U7368 (N_7368,N_2472,N_2712);
xor U7369 (N_7369,N_2495,N_3204);
nand U7370 (N_7370,N_675,N_650);
xor U7371 (N_7371,N_2430,N_2971);
xnor U7372 (N_7372,N_4479,N_1617);
or U7373 (N_7373,N_3698,N_1313);
xor U7374 (N_7374,N_1300,N_2424);
and U7375 (N_7375,N_1074,N_3262);
and U7376 (N_7376,N_4316,N_320);
or U7377 (N_7377,N_1734,N_4499);
or U7378 (N_7378,N_2085,N_451);
nor U7379 (N_7379,N_1715,N_3439);
xor U7380 (N_7380,N_2731,N_319);
and U7381 (N_7381,N_248,N_3856);
xnor U7382 (N_7382,N_2279,N_3594);
nor U7383 (N_7383,N_2636,N_1241);
nand U7384 (N_7384,N_1522,N_4730);
xor U7385 (N_7385,N_4562,N_1140);
or U7386 (N_7386,N_3727,N_3072);
xnor U7387 (N_7387,N_687,N_2310);
xor U7388 (N_7388,N_15,N_547);
nor U7389 (N_7389,N_3232,N_4614);
nor U7390 (N_7390,N_2614,N_1834);
xor U7391 (N_7391,N_2909,N_1977);
or U7392 (N_7392,N_4416,N_2479);
xor U7393 (N_7393,N_4065,N_2988);
and U7394 (N_7394,N_1287,N_937);
and U7395 (N_7395,N_1574,N_4500);
nor U7396 (N_7396,N_4931,N_3835);
and U7397 (N_7397,N_3295,N_510);
and U7398 (N_7398,N_2576,N_143);
xor U7399 (N_7399,N_4466,N_2436);
nand U7400 (N_7400,N_2806,N_4551);
nand U7401 (N_7401,N_2213,N_1814);
and U7402 (N_7402,N_1525,N_4884);
nand U7403 (N_7403,N_1717,N_59);
and U7404 (N_7404,N_2524,N_1405);
nor U7405 (N_7405,N_2901,N_43);
or U7406 (N_7406,N_169,N_774);
nor U7407 (N_7407,N_2482,N_4133);
xnor U7408 (N_7408,N_4075,N_1133);
or U7409 (N_7409,N_1035,N_1175);
nor U7410 (N_7410,N_2691,N_4616);
and U7411 (N_7411,N_4039,N_4854);
nor U7412 (N_7412,N_3450,N_109);
or U7413 (N_7413,N_3505,N_4917);
nand U7414 (N_7414,N_1470,N_519);
and U7415 (N_7415,N_4487,N_4845);
nand U7416 (N_7416,N_3769,N_2854);
nor U7417 (N_7417,N_3215,N_3328);
xor U7418 (N_7418,N_653,N_2714);
nand U7419 (N_7419,N_560,N_816);
or U7420 (N_7420,N_2655,N_4430);
nor U7421 (N_7421,N_4386,N_3686);
or U7422 (N_7422,N_4028,N_4636);
and U7423 (N_7423,N_4634,N_3472);
nor U7424 (N_7424,N_1989,N_4166);
nor U7425 (N_7425,N_3394,N_3486);
nand U7426 (N_7426,N_1918,N_1716);
nand U7427 (N_7427,N_1956,N_2564);
nand U7428 (N_7428,N_3042,N_1395);
nand U7429 (N_7429,N_2892,N_2365);
or U7430 (N_7430,N_2225,N_3708);
nand U7431 (N_7431,N_2183,N_4287);
nor U7432 (N_7432,N_228,N_1831);
xnor U7433 (N_7433,N_2449,N_1199);
or U7434 (N_7434,N_1865,N_2647);
xor U7435 (N_7435,N_1083,N_2704);
and U7436 (N_7436,N_4447,N_1343);
and U7437 (N_7437,N_1285,N_3347);
or U7438 (N_7438,N_4879,N_4921);
nand U7439 (N_7439,N_1549,N_3062);
or U7440 (N_7440,N_1891,N_2474);
nor U7441 (N_7441,N_2515,N_3964);
xnor U7442 (N_7442,N_2451,N_2990);
and U7443 (N_7443,N_1453,N_1585);
or U7444 (N_7444,N_4605,N_4088);
and U7445 (N_7445,N_3288,N_2302);
nor U7446 (N_7446,N_2930,N_683);
xnor U7447 (N_7447,N_4980,N_1579);
nand U7448 (N_7448,N_1355,N_930);
nand U7449 (N_7449,N_1123,N_586);
nand U7450 (N_7450,N_838,N_2362);
nor U7451 (N_7451,N_3781,N_3403);
xor U7452 (N_7452,N_304,N_1018);
or U7453 (N_7453,N_133,N_3415);
nand U7454 (N_7454,N_2831,N_820);
or U7455 (N_7455,N_4750,N_3587);
nor U7456 (N_7456,N_4157,N_1097);
nand U7457 (N_7457,N_7,N_278);
and U7458 (N_7458,N_1555,N_1306);
xor U7459 (N_7459,N_3920,N_1963);
nand U7460 (N_7460,N_3195,N_2175);
and U7461 (N_7461,N_4861,N_4895);
nor U7462 (N_7462,N_1628,N_1569);
nor U7463 (N_7463,N_3995,N_3003);
and U7464 (N_7464,N_856,N_3247);
nand U7465 (N_7465,N_1382,N_3157);
or U7466 (N_7466,N_3869,N_3674);
nand U7467 (N_7467,N_4182,N_2581);
nand U7468 (N_7468,N_4310,N_2847);
and U7469 (N_7469,N_1860,N_2352);
nand U7470 (N_7470,N_4714,N_543);
nor U7471 (N_7471,N_1394,N_3695);
or U7472 (N_7472,N_3128,N_2052);
nor U7473 (N_7473,N_3863,N_288);
or U7474 (N_7474,N_1594,N_1107);
nor U7475 (N_7475,N_2226,N_4474);
and U7476 (N_7476,N_4108,N_2755);
nor U7477 (N_7477,N_3506,N_102);
or U7478 (N_7478,N_2463,N_2374);
nor U7479 (N_7479,N_974,N_1632);
or U7480 (N_7480,N_3694,N_2143);
or U7481 (N_7481,N_4229,N_3508);
and U7482 (N_7482,N_4457,N_2037);
nand U7483 (N_7483,N_1791,N_4662);
or U7484 (N_7484,N_1210,N_1796);
nand U7485 (N_7485,N_3056,N_961);
nor U7486 (N_7486,N_4973,N_4128);
nand U7487 (N_7487,N_1583,N_509);
xnor U7488 (N_7488,N_4637,N_4050);
xnor U7489 (N_7489,N_3142,N_786);
nand U7490 (N_7490,N_31,N_1727);
or U7491 (N_7491,N_646,N_289);
or U7492 (N_7492,N_1162,N_2393);
nor U7493 (N_7493,N_4397,N_373);
and U7494 (N_7494,N_688,N_3728);
nor U7495 (N_7495,N_4698,N_371);
or U7496 (N_7496,N_3975,N_366);
nand U7497 (N_7497,N_3680,N_2976);
nor U7498 (N_7498,N_4475,N_226);
xnor U7499 (N_7499,N_3534,N_531);
and U7500 (N_7500,N_461,N_1825);
or U7501 (N_7501,N_870,N_2798);
and U7502 (N_7502,N_1422,N_1486);
nand U7503 (N_7503,N_4552,N_1096);
or U7504 (N_7504,N_1797,N_1020);
xor U7505 (N_7505,N_3851,N_4028);
xnor U7506 (N_7506,N_290,N_3951);
nor U7507 (N_7507,N_2406,N_2389);
or U7508 (N_7508,N_2149,N_3361);
and U7509 (N_7509,N_2101,N_1045);
and U7510 (N_7510,N_2514,N_2081);
nand U7511 (N_7511,N_1911,N_3140);
nor U7512 (N_7512,N_4571,N_348);
or U7513 (N_7513,N_2266,N_463);
nand U7514 (N_7514,N_25,N_3720);
or U7515 (N_7515,N_3533,N_1875);
nand U7516 (N_7516,N_1034,N_2981);
xor U7517 (N_7517,N_2088,N_924);
nor U7518 (N_7518,N_2210,N_50);
or U7519 (N_7519,N_4136,N_3726);
xnor U7520 (N_7520,N_4394,N_541);
or U7521 (N_7521,N_2905,N_146);
or U7522 (N_7522,N_3766,N_428);
or U7523 (N_7523,N_67,N_4619);
nor U7524 (N_7524,N_4070,N_1255);
and U7525 (N_7525,N_549,N_2278);
xnor U7526 (N_7526,N_4286,N_1269);
and U7527 (N_7527,N_0,N_4994);
nand U7528 (N_7528,N_613,N_2039);
nor U7529 (N_7529,N_4032,N_4892);
or U7530 (N_7530,N_1850,N_3077);
nor U7531 (N_7531,N_1455,N_4418);
nand U7532 (N_7532,N_4405,N_2125);
and U7533 (N_7533,N_4112,N_3644);
nand U7534 (N_7534,N_1973,N_2154);
and U7535 (N_7535,N_3380,N_147);
nand U7536 (N_7536,N_3163,N_1954);
nand U7537 (N_7537,N_1168,N_4612);
or U7538 (N_7538,N_1926,N_2264);
xnor U7539 (N_7539,N_2872,N_2502);
xnor U7540 (N_7540,N_2573,N_2620);
and U7541 (N_7541,N_4540,N_1026);
nand U7542 (N_7542,N_4685,N_626);
or U7543 (N_7543,N_3732,N_2980);
and U7544 (N_7544,N_1633,N_1742);
nand U7545 (N_7545,N_4100,N_4808);
xor U7546 (N_7546,N_600,N_2884);
and U7547 (N_7547,N_2920,N_4333);
or U7548 (N_7548,N_434,N_4497);
nand U7549 (N_7549,N_3834,N_1709);
nor U7550 (N_7550,N_854,N_2318);
or U7551 (N_7551,N_4828,N_4206);
nor U7552 (N_7552,N_1513,N_4733);
and U7553 (N_7553,N_4943,N_1492);
nand U7554 (N_7554,N_3380,N_4683);
and U7555 (N_7555,N_974,N_1818);
nor U7556 (N_7556,N_1100,N_2220);
or U7557 (N_7557,N_328,N_1886);
or U7558 (N_7558,N_2918,N_2804);
nand U7559 (N_7559,N_4295,N_921);
nor U7560 (N_7560,N_118,N_1077);
and U7561 (N_7561,N_4461,N_1743);
or U7562 (N_7562,N_3876,N_3922);
or U7563 (N_7563,N_2062,N_4503);
nand U7564 (N_7564,N_4897,N_3014);
xor U7565 (N_7565,N_855,N_2897);
xnor U7566 (N_7566,N_2239,N_2203);
or U7567 (N_7567,N_4048,N_2430);
xor U7568 (N_7568,N_1064,N_1193);
and U7569 (N_7569,N_850,N_505);
and U7570 (N_7570,N_1985,N_81);
nor U7571 (N_7571,N_1529,N_348);
nor U7572 (N_7572,N_710,N_3118);
nor U7573 (N_7573,N_3195,N_1174);
and U7574 (N_7574,N_30,N_4270);
nor U7575 (N_7575,N_413,N_2769);
nor U7576 (N_7576,N_392,N_2112);
nor U7577 (N_7577,N_1083,N_4490);
nand U7578 (N_7578,N_310,N_4693);
nor U7579 (N_7579,N_4939,N_4172);
and U7580 (N_7580,N_3988,N_3331);
or U7581 (N_7581,N_4569,N_3911);
and U7582 (N_7582,N_1489,N_1879);
xnor U7583 (N_7583,N_2442,N_651);
or U7584 (N_7584,N_2217,N_3484);
and U7585 (N_7585,N_911,N_4122);
nor U7586 (N_7586,N_3231,N_4373);
nand U7587 (N_7587,N_2387,N_709);
or U7588 (N_7588,N_1074,N_4531);
or U7589 (N_7589,N_878,N_3224);
nor U7590 (N_7590,N_3212,N_3330);
nand U7591 (N_7591,N_1787,N_2846);
or U7592 (N_7592,N_1995,N_850);
nand U7593 (N_7593,N_2602,N_2937);
or U7594 (N_7594,N_1333,N_3269);
xnor U7595 (N_7595,N_1884,N_3713);
and U7596 (N_7596,N_4167,N_1686);
xor U7597 (N_7597,N_1088,N_4185);
nor U7598 (N_7598,N_1543,N_2848);
nor U7599 (N_7599,N_4445,N_1572);
nand U7600 (N_7600,N_1172,N_2290);
and U7601 (N_7601,N_1213,N_1208);
xnor U7602 (N_7602,N_2306,N_421);
nor U7603 (N_7603,N_482,N_1199);
or U7604 (N_7604,N_965,N_7);
xnor U7605 (N_7605,N_522,N_253);
or U7606 (N_7606,N_2454,N_572);
nand U7607 (N_7607,N_200,N_2821);
or U7608 (N_7608,N_560,N_2251);
nand U7609 (N_7609,N_1013,N_1391);
and U7610 (N_7610,N_4546,N_3177);
nor U7611 (N_7611,N_4543,N_967);
nor U7612 (N_7612,N_1725,N_4877);
and U7613 (N_7613,N_1734,N_1857);
xnor U7614 (N_7614,N_470,N_2161);
nand U7615 (N_7615,N_2740,N_3676);
or U7616 (N_7616,N_2728,N_2616);
xor U7617 (N_7617,N_3316,N_4198);
xnor U7618 (N_7618,N_4776,N_4242);
xnor U7619 (N_7619,N_1984,N_4077);
xnor U7620 (N_7620,N_2538,N_1497);
xnor U7621 (N_7621,N_1972,N_19);
nand U7622 (N_7622,N_568,N_1725);
nor U7623 (N_7623,N_1934,N_699);
nor U7624 (N_7624,N_4416,N_532);
xnor U7625 (N_7625,N_1052,N_1189);
and U7626 (N_7626,N_3157,N_4122);
nor U7627 (N_7627,N_2962,N_3117);
xnor U7628 (N_7628,N_1670,N_2297);
or U7629 (N_7629,N_442,N_3603);
nor U7630 (N_7630,N_1174,N_2088);
nor U7631 (N_7631,N_2398,N_4169);
nor U7632 (N_7632,N_2483,N_1787);
nand U7633 (N_7633,N_1996,N_2043);
and U7634 (N_7634,N_206,N_2636);
nand U7635 (N_7635,N_3405,N_3324);
or U7636 (N_7636,N_1381,N_2731);
xor U7637 (N_7637,N_4834,N_746);
and U7638 (N_7638,N_3535,N_4941);
or U7639 (N_7639,N_745,N_3260);
nor U7640 (N_7640,N_808,N_799);
nor U7641 (N_7641,N_836,N_832);
xor U7642 (N_7642,N_4416,N_319);
xnor U7643 (N_7643,N_3748,N_642);
nor U7644 (N_7644,N_4612,N_471);
or U7645 (N_7645,N_4410,N_2783);
nand U7646 (N_7646,N_3824,N_1790);
or U7647 (N_7647,N_955,N_2749);
xnor U7648 (N_7648,N_1988,N_2865);
or U7649 (N_7649,N_3700,N_1637);
xnor U7650 (N_7650,N_3477,N_2236);
and U7651 (N_7651,N_2521,N_2044);
xnor U7652 (N_7652,N_1946,N_4631);
nor U7653 (N_7653,N_3055,N_4489);
or U7654 (N_7654,N_2738,N_4083);
nand U7655 (N_7655,N_4972,N_4640);
and U7656 (N_7656,N_2283,N_919);
nor U7657 (N_7657,N_3118,N_2);
nand U7658 (N_7658,N_464,N_2293);
xor U7659 (N_7659,N_2751,N_3623);
nor U7660 (N_7660,N_1026,N_2755);
nand U7661 (N_7661,N_4096,N_3954);
and U7662 (N_7662,N_3242,N_2679);
nand U7663 (N_7663,N_98,N_1238);
and U7664 (N_7664,N_352,N_2011);
or U7665 (N_7665,N_2388,N_2681);
xor U7666 (N_7666,N_732,N_1979);
nand U7667 (N_7667,N_785,N_1486);
and U7668 (N_7668,N_1485,N_4917);
and U7669 (N_7669,N_4031,N_1487);
and U7670 (N_7670,N_53,N_3264);
or U7671 (N_7671,N_4642,N_368);
nand U7672 (N_7672,N_463,N_2870);
and U7673 (N_7673,N_1515,N_3084);
and U7674 (N_7674,N_2745,N_1799);
or U7675 (N_7675,N_4920,N_389);
nand U7676 (N_7676,N_4754,N_3375);
nor U7677 (N_7677,N_1803,N_2125);
nand U7678 (N_7678,N_3854,N_3220);
and U7679 (N_7679,N_2279,N_3191);
nand U7680 (N_7680,N_2577,N_310);
and U7681 (N_7681,N_4949,N_4651);
nor U7682 (N_7682,N_4952,N_2170);
xnor U7683 (N_7683,N_1932,N_1191);
and U7684 (N_7684,N_1708,N_4223);
or U7685 (N_7685,N_199,N_1663);
xnor U7686 (N_7686,N_2851,N_1216);
nand U7687 (N_7687,N_3101,N_4158);
nand U7688 (N_7688,N_118,N_1068);
nor U7689 (N_7689,N_4298,N_450);
nor U7690 (N_7690,N_1049,N_899);
nor U7691 (N_7691,N_327,N_2860);
nand U7692 (N_7692,N_265,N_416);
nand U7693 (N_7693,N_1739,N_4694);
xnor U7694 (N_7694,N_2939,N_1220);
xnor U7695 (N_7695,N_43,N_4969);
nand U7696 (N_7696,N_3090,N_1703);
or U7697 (N_7697,N_2759,N_196);
xor U7698 (N_7698,N_4391,N_1008);
nand U7699 (N_7699,N_3876,N_2533);
xnor U7700 (N_7700,N_4824,N_2648);
and U7701 (N_7701,N_2793,N_880);
nor U7702 (N_7702,N_2927,N_2249);
nor U7703 (N_7703,N_553,N_2028);
nand U7704 (N_7704,N_431,N_4473);
or U7705 (N_7705,N_562,N_1663);
nand U7706 (N_7706,N_90,N_1442);
and U7707 (N_7707,N_2820,N_321);
nand U7708 (N_7708,N_742,N_2552);
nor U7709 (N_7709,N_105,N_4889);
and U7710 (N_7710,N_1386,N_379);
and U7711 (N_7711,N_780,N_747);
nor U7712 (N_7712,N_2105,N_439);
xor U7713 (N_7713,N_3119,N_2238);
nand U7714 (N_7714,N_4436,N_652);
nor U7715 (N_7715,N_2091,N_625);
or U7716 (N_7716,N_975,N_2094);
xnor U7717 (N_7717,N_1401,N_1122);
or U7718 (N_7718,N_1300,N_3742);
nor U7719 (N_7719,N_3490,N_3044);
nand U7720 (N_7720,N_1122,N_233);
xor U7721 (N_7721,N_4450,N_819);
nand U7722 (N_7722,N_127,N_1054);
nor U7723 (N_7723,N_3386,N_795);
and U7724 (N_7724,N_1972,N_878);
nor U7725 (N_7725,N_3832,N_2294);
nand U7726 (N_7726,N_950,N_4505);
or U7727 (N_7727,N_4012,N_1753);
xor U7728 (N_7728,N_1335,N_4321);
nor U7729 (N_7729,N_4497,N_2494);
xnor U7730 (N_7730,N_1953,N_2103);
or U7731 (N_7731,N_1432,N_232);
and U7732 (N_7732,N_1320,N_940);
xnor U7733 (N_7733,N_2605,N_817);
nand U7734 (N_7734,N_3884,N_1265);
nor U7735 (N_7735,N_2070,N_2093);
and U7736 (N_7736,N_4116,N_1663);
xor U7737 (N_7737,N_815,N_3614);
and U7738 (N_7738,N_420,N_3468);
or U7739 (N_7739,N_4633,N_3632);
or U7740 (N_7740,N_785,N_2269);
and U7741 (N_7741,N_662,N_4968);
nor U7742 (N_7742,N_4601,N_1237);
and U7743 (N_7743,N_1082,N_2386);
or U7744 (N_7744,N_4830,N_3175);
nand U7745 (N_7745,N_4749,N_4689);
xor U7746 (N_7746,N_346,N_950);
and U7747 (N_7747,N_2332,N_2141);
and U7748 (N_7748,N_3025,N_758);
and U7749 (N_7749,N_3188,N_2481);
nand U7750 (N_7750,N_50,N_4838);
nand U7751 (N_7751,N_4014,N_384);
nand U7752 (N_7752,N_3308,N_1698);
or U7753 (N_7753,N_1151,N_2385);
and U7754 (N_7754,N_2236,N_4548);
nand U7755 (N_7755,N_2779,N_3498);
and U7756 (N_7756,N_366,N_4712);
or U7757 (N_7757,N_2095,N_4752);
and U7758 (N_7758,N_3455,N_1362);
and U7759 (N_7759,N_1021,N_2449);
nand U7760 (N_7760,N_3891,N_2414);
xor U7761 (N_7761,N_3139,N_2168);
and U7762 (N_7762,N_4778,N_3099);
nor U7763 (N_7763,N_399,N_4425);
xnor U7764 (N_7764,N_1725,N_4111);
nor U7765 (N_7765,N_2377,N_3931);
and U7766 (N_7766,N_3540,N_2092);
and U7767 (N_7767,N_4768,N_2085);
or U7768 (N_7768,N_1260,N_1696);
xnor U7769 (N_7769,N_2744,N_1757);
xor U7770 (N_7770,N_3436,N_3866);
and U7771 (N_7771,N_2970,N_519);
nor U7772 (N_7772,N_2537,N_763);
xor U7773 (N_7773,N_791,N_2369);
xor U7774 (N_7774,N_1515,N_1592);
nor U7775 (N_7775,N_1107,N_810);
nor U7776 (N_7776,N_1988,N_1456);
xnor U7777 (N_7777,N_2144,N_4543);
xor U7778 (N_7778,N_4123,N_784);
and U7779 (N_7779,N_4750,N_3785);
or U7780 (N_7780,N_3422,N_2276);
or U7781 (N_7781,N_496,N_1729);
and U7782 (N_7782,N_2713,N_648);
nor U7783 (N_7783,N_374,N_2211);
xor U7784 (N_7784,N_3837,N_3723);
nor U7785 (N_7785,N_668,N_1977);
nand U7786 (N_7786,N_3030,N_4976);
nand U7787 (N_7787,N_2871,N_4198);
nand U7788 (N_7788,N_2936,N_3705);
nand U7789 (N_7789,N_3690,N_389);
and U7790 (N_7790,N_3774,N_532);
or U7791 (N_7791,N_845,N_2179);
or U7792 (N_7792,N_1879,N_805);
nor U7793 (N_7793,N_3650,N_3789);
or U7794 (N_7794,N_4003,N_4378);
and U7795 (N_7795,N_2499,N_4983);
xor U7796 (N_7796,N_3984,N_1000);
and U7797 (N_7797,N_107,N_397);
or U7798 (N_7798,N_1948,N_4116);
or U7799 (N_7799,N_1508,N_4347);
xnor U7800 (N_7800,N_4822,N_4602);
or U7801 (N_7801,N_3086,N_1931);
xor U7802 (N_7802,N_488,N_2823);
or U7803 (N_7803,N_4131,N_1843);
and U7804 (N_7804,N_2263,N_530);
or U7805 (N_7805,N_2889,N_3251);
and U7806 (N_7806,N_2338,N_2306);
or U7807 (N_7807,N_2187,N_1133);
xor U7808 (N_7808,N_2913,N_4811);
xor U7809 (N_7809,N_1697,N_4105);
nand U7810 (N_7810,N_2254,N_2575);
nor U7811 (N_7811,N_1735,N_3626);
and U7812 (N_7812,N_2932,N_1525);
nor U7813 (N_7813,N_1201,N_3855);
nand U7814 (N_7814,N_2863,N_1394);
nor U7815 (N_7815,N_1365,N_318);
xor U7816 (N_7816,N_586,N_4357);
xor U7817 (N_7817,N_1295,N_2390);
or U7818 (N_7818,N_4761,N_2167);
nand U7819 (N_7819,N_961,N_4273);
and U7820 (N_7820,N_3606,N_3398);
nor U7821 (N_7821,N_3767,N_541);
nand U7822 (N_7822,N_2453,N_377);
and U7823 (N_7823,N_4006,N_1697);
and U7824 (N_7824,N_2283,N_3186);
nand U7825 (N_7825,N_2848,N_1374);
nor U7826 (N_7826,N_1199,N_123);
or U7827 (N_7827,N_3516,N_722);
nor U7828 (N_7828,N_3417,N_4314);
nand U7829 (N_7829,N_4809,N_957);
xnor U7830 (N_7830,N_659,N_4015);
and U7831 (N_7831,N_4976,N_2692);
xnor U7832 (N_7832,N_1160,N_4621);
and U7833 (N_7833,N_3710,N_2509);
and U7834 (N_7834,N_3426,N_907);
xor U7835 (N_7835,N_1947,N_1437);
or U7836 (N_7836,N_668,N_4123);
and U7837 (N_7837,N_4775,N_1073);
or U7838 (N_7838,N_3858,N_2739);
nor U7839 (N_7839,N_351,N_2911);
or U7840 (N_7840,N_658,N_1302);
or U7841 (N_7841,N_647,N_3000);
or U7842 (N_7842,N_50,N_2878);
nand U7843 (N_7843,N_4217,N_3291);
nor U7844 (N_7844,N_349,N_2142);
and U7845 (N_7845,N_2084,N_238);
or U7846 (N_7846,N_756,N_2121);
xnor U7847 (N_7847,N_4157,N_1657);
or U7848 (N_7848,N_4837,N_1538);
and U7849 (N_7849,N_2361,N_3630);
nand U7850 (N_7850,N_3426,N_2188);
and U7851 (N_7851,N_1207,N_3305);
nand U7852 (N_7852,N_4211,N_1652);
nand U7853 (N_7853,N_1099,N_3616);
or U7854 (N_7854,N_4681,N_2810);
nand U7855 (N_7855,N_4496,N_2469);
nand U7856 (N_7856,N_637,N_1202);
and U7857 (N_7857,N_1308,N_3638);
or U7858 (N_7858,N_3737,N_3494);
nor U7859 (N_7859,N_3529,N_1410);
xnor U7860 (N_7860,N_985,N_1933);
and U7861 (N_7861,N_1320,N_2312);
nand U7862 (N_7862,N_1691,N_464);
nor U7863 (N_7863,N_2151,N_3386);
xnor U7864 (N_7864,N_2295,N_3225);
xnor U7865 (N_7865,N_4617,N_3702);
xor U7866 (N_7866,N_2108,N_2415);
xor U7867 (N_7867,N_2194,N_4688);
nand U7868 (N_7868,N_525,N_1779);
and U7869 (N_7869,N_1080,N_1782);
xnor U7870 (N_7870,N_342,N_3797);
or U7871 (N_7871,N_417,N_3360);
and U7872 (N_7872,N_4683,N_245);
xnor U7873 (N_7873,N_3146,N_984);
or U7874 (N_7874,N_1423,N_4927);
or U7875 (N_7875,N_1368,N_4744);
or U7876 (N_7876,N_1306,N_295);
nor U7877 (N_7877,N_2887,N_2816);
and U7878 (N_7878,N_2316,N_4783);
nor U7879 (N_7879,N_3026,N_2749);
xor U7880 (N_7880,N_2431,N_4624);
nand U7881 (N_7881,N_3261,N_1843);
nor U7882 (N_7882,N_4386,N_2332);
xnor U7883 (N_7883,N_669,N_2648);
nor U7884 (N_7884,N_760,N_1479);
and U7885 (N_7885,N_2878,N_2975);
and U7886 (N_7886,N_1918,N_2710);
xor U7887 (N_7887,N_2083,N_444);
or U7888 (N_7888,N_2926,N_3079);
and U7889 (N_7889,N_2696,N_2276);
nor U7890 (N_7890,N_2314,N_1495);
and U7891 (N_7891,N_1770,N_2691);
or U7892 (N_7892,N_4923,N_3826);
xnor U7893 (N_7893,N_3020,N_3390);
nor U7894 (N_7894,N_3020,N_3947);
nand U7895 (N_7895,N_4708,N_1350);
and U7896 (N_7896,N_583,N_473);
or U7897 (N_7897,N_3321,N_3279);
xnor U7898 (N_7898,N_2520,N_3033);
nand U7899 (N_7899,N_3697,N_4216);
or U7900 (N_7900,N_417,N_4610);
nor U7901 (N_7901,N_2852,N_3961);
or U7902 (N_7902,N_886,N_165);
or U7903 (N_7903,N_3404,N_2);
nor U7904 (N_7904,N_713,N_1017);
or U7905 (N_7905,N_1779,N_1497);
nand U7906 (N_7906,N_3219,N_1505);
and U7907 (N_7907,N_668,N_1232);
and U7908 (N_7908,N_1874,N_3486);
xnor U7909 (N_7909,N_963,N_1040);
nand U7910 (N_7910,N_2154,N_969);
xor U7911 (N_7911,N_3580,N_3008);
nor U7912 (N_7912,N_2618,N_1053);
nor U7913 (N_7913,N_1243,N_2909);
and U7914 (N_7914,N_3715,N_876);
nand U7915 (N_7915,N_2879,N_2721);
nand U7916 (N_7916,N_633,N_1737);
nand U7917 (N_7917,N_3917,N_336);
xor U7918 (N_7918,N_3815,N_1631);
nor U7919 (N_7919,N_4638,N_318);
nand U7920 (N_7920,N_2094,N_2259);
nor U7921 (N_7921,N_2306,N_3120);
and U7922 (N_7922,N_797,N_734);
or U7923 (N_7923,N_220,N_3527);
and U7924 (N_7924,N_3428,N_1946);
nor U7925 (N_7925,N_2674,N_771);
nor U7926 (N_7926,N_822,N_339);
and U7927 (N_7927,N_1456,N_3623);
and U7928 (N_7928,N_1187,N_219);
nand U7929 (N_7929,N_4230,N_2680);
and U7930 (N_7930,N_1580,N_3152);
or U7931 (N_7931,N_3905,N_556);
nor U7932 (N_7932,N_1360,N_2733);
nor U7933 (N_7933,N_572,N_1898);
and U7934 (N_7934,N_3849,N_2080);
or U7935 (N_7935,N_353,N_4804);
and U7936 (N_7936,N_768,N_4800);
nand U7937 (N_7937,N_1371,N_3246);
nor U7938 (N_7938,N_4616,N_4696);
or U7939 (N_7939,N_2729,N_3071);
nor U7940 (N_7940,N_3328,N_658);
xor U7941 (N_7941,N_4805,N_2883);
and U7942 (N_7942,N_1604,N_3164);
xnor U7943 (N_7943,N_859,N_210);
or U7944 (N_7944,N_1757,N_3564);
or U7945 (N_7945,N_3967,N_1595);
nor U7946 (N_7946,N_727,N_3354);
and U7947 (N_7947,N_1290,N_2185);
nand U7948 (N_7948,N_4150,N_1351);
and U7949 (N_7949,N_4691,N_1483);
xnor U7950 (N_7950,N_4933,N_647);
and U7951 (N_7951,N_2007,N_2584);
nor U7952 (N_7952,N_2598,N_3408);
and U7953 (N_7953,N_3200,N_1546);
and U7954 (N_7954,N_1753,N_2655);
nor U7955 (N_7955,N_1936,N_3740);
nor U7956 (N_7956,N_1544,N_3520);
and U7957 (N_7957,N_2282,N_4679);
nand U7958 (N_7958,N_854,N_3428);
and U7959 (N_7959,N_3218,N_2677);
nand U7960 (N_7960,N_3800,N_1008);
nor U7961 (N_7961,N_2481,N_2618);
xnor U7962 (N_7962,N_2039,N_4447);
nand U7963 (N_7963,N_2206,N_929);
nor U7964 (N_7964,N_3194,N_4921);
and U7965 (N_7965,N_4386,N_3938);
xnor U7966 (N_7966,N_944,N_2270);
xnor U7967 (N_7967,N_3065,N_709);
nand U7968 (N_7968,N_3651,N_784);
nor U7969 (N_7969,N_2024,N_3150);
and U7970 (N_7970,N_3897,N_263);
nor U7971 (N_7971,N_265,N_1139);
or U7972 (N_7972,N_2055,N_2989);
xor U7973 (N_7973,N_1173,N_2869);
nor U7974 (N_7974,N_3705,N_4969);
nand U7975 (N_7975,N_1460,N_2588);
nand U7976 (N_7976,N_3779,N_3024);
and U7977 (N_7977,N_1482,N_2691);
nor U7978 (N_7978,N_3338,N_285);
nand U7979 (N_7979,N_4521,N_307);
nor U7980 (N_7980,N_4635,N_1162);
or U7981 (N_7981,N_35,N_1064);
nand U7982 (N_7982,N_4416,N_1308);
nand U7983 (N_7983,N_2866,N_1331);
nor U7984 (N_7984,N_2840,N_952);
and U7985 (N_7985,N_3329,N_2831);
xnor U7986 (N_7986,N_3045,N_1333);
nand U7987 (N_7987,N_3256,N_1436);
nand U7988 (N_7988,N_713,N_2174);
nand U7989 (N_7989,N_4965,N_3919);
xor U7990 (N_7990,N_2855,N_905);
nand U7991 (N_7991,N_2088,N_3866);
nor U7992 (N_7992,N_4393,N_329);
nor U7993 (N_7993,N_3695,N_2201);
xnor U7994 (N_7994,N_2578,N_355);
nor U7995 (N_7995,N_2844,N_4942);
or U7996 (N_7996,N_1877,N_4875);
or U7997 (N_7997,N_2361,N_4125);
xor U7998 (N_7998,N_4946,N_3286);
nand U7999 (N_7999,N_2770,N_2437);
or U8000 (N_8000,N_4560,N_4010);
nor U8001 (N_8001,N_4244,N_4621);
xnor U8002 (N_8002,N_3201,N_1817);
or U8003 (N_8003,N_436,N_3873);
xnor U8004 (N_8004,N_2588,N_520);
xor U8005 (N_8005,N_1747,N_265);
or U8006 (N_8006,N_472,N_4423);
xor U8007 (N_8007,N_3733,N_3441);
or U8008 (N_8008,N_2290,N_3111);
xor U8009 (N_8009,N_2881,N_611);
and U8010 (N_8010,N_1375,N_2739);
or U8011 (N_8011,N_1089,N_3339);
nor U8012 (N_8012,N_3611,N_329);
xor U8013 (N_8013,N_2493,N_4734);
and U8014 (N_8014,N_3692,N_2402);
nor U8015 (N_8015,N_3345,N_2480);
nand U8016 (N_8016,N_2331,N_1520);
nor U8017 (N_8017,N_530,N_2593);
nor U8018 (N_8018,N_3028,N_2869);
or U8019 (N_8019,N_4793,N_1399);
nor U8020 (N_8020,N_1452,N_1523);
nor U8021 (N_8021,N_4154,N_4550);
xor U8022 (N_8022,N_1300,N_3503);
xnor U8023 (N_8023,N_4528,N_2256);
and U8024 (N_8024,N_1931,N_622);
or U8025 (N_8025,N_359,N_747);
nor U8026 (N_8026,N_3030,N_377);
and U8027 (N_8027,N_2179,N_4974);
xnor U8028 (N_8028,N_873,N_1982);
xnor U8029 (N_8029,N_2153,N_944);
xor U8030 (N_8030,N_3296,N_402);
and U8031 (N_8031,N_615,N_3654);
nor U8032 (N_8032,N_4707,N_4722);
or U8033 (N_8033,N_3580,N_30);
or U8034 (N_8034,N_2180,N_4616);
nor U8035 (N_8035,N_3649,N_2906);
xnor U8036 (N_8036,N_137,N_4295);
or U8037 (N_8037,N_2956,N_3696);
and U8038 (N_8038,N_3396,N_3131);
nand U8039 (N_8039,N_4308,N_1052);
nand U8040 (N_8040,N_3502,N_827);
or U8041 (N_8041,N_826,N_2252);
nor U8042 (N_8042,N_2681,N_1425);
and U8043 (N_8043,N_1525,N_1776);
or U8044 (N_8044,N_1841,N_2310);
nor U8045 (N_8045,N_6,N_4722);
nor U8046 (N_8046,N_2132,N_2564);
nor U8047 (N_8047,N_2138,N_2292);
or U8048 (N_8048,N_3613,N_3132);
xnor U8049 (N_8049,N_4792,N_629);
nor U8050 (N_8050,N_2369,N_3228);
nand U8051 (N_8051,N_1869,N_1996);
nand U8052 (N_8052,N_3326,N_2800);
and U8053 (N_8053,N_2475,N_1650);
and U8054 (N_8054,N_4062,N_775);
nor U8055 (N_8055,N_2098,N_2619);
xor U8056 (N_8056,N_571,N_3992);
or U8057 (N_8057,N_3751,N_162);
and U8058 (N_8058,N_4223,N_1781);
and U8059 (N_8059,N_2275,N_4500);
xor U8060 (N_8060,N_1823,N_4977);
nand U8061 (N_8061,N_3882,N_1316);
nor U8062 (N_8062,N_16,N_2979);
or U8063 (N_8063,N_1967,N_983);
nand U8064 (N_8064,N_3050,N_608);
nor U8065 (N_8065,N_2050,N_1982);
nor U8066 (N_8066,N_2665,N_4821);
and U8067 (N_8067,N_2778,N_3873);
nor U8068 (N_8068,N_4974,N_116);
nor U8069 (N_8069,N_4583,N_2841);
and U8070 (N_8070,N_4392,N_2219);
or U8071 (N_8071,N_4656,N_769);
nand U8072 (N_8072,N_3107,N_3077);
or U8073 (N_8073,N_326,N_2809);
nand U8074 (N_8074,N_4009,N_4343);
nor U8075 (N_8075,N_650,N_146);
or U8076 (N_8076,N_332,N_2864);
nand U8077 (N_8077,N_3336,N_719);
or U8078 (N_8078,N_1655,N_2387);
and U8079 (N_8079,N_4835,N_3430);
and U8080 (N_8080,N_4444,N_1713);
nand U8081 (N_8081,N_4682,N_2821);
xnor U8082 (N_8082,N_1891,N_3698);
nand U8083 (N_8083,N_567,N_2237);
and U8084 (N_8084,N_3247,N_977);
nand U8085 (N_8085,N_3618,N_767);
xnor U8086 (N_8086,N_1203,N_1213);
xnor U8087 (N_8087,N_4731,N_2133);
xnor U8088 (N_8088,N_1576,N_2740);
or U8089 (N_8089,N_4363,N_2023);
nor U8090 (N_8090,N_1940,N_3029);
nor U8091 (N_8091,N_4031,N_1897);
xnor U8092 (N_8092,N_4280,N_1108);
xnor U8093 (N_8093,N_2513,N_3506);
and U8094 (N_8094,N_3043,N_3680);
nand U8095 (N_8095,N_3656,N_2077);
xnor U8096 (N_8096,N_3188,N_4830);
nand U8097 (N_8097,N_2831,N_2294);
nor U8098 (N_8098,N_1202,N_3290);
and U8099 (N_8099,N_16,N_188);
nor U8100 (N_8100,N_3790,N_4663);
and U8101 (N_8101,N_3394,N_708);
nand U8102 (N_8102,N_224,N_3254);
or U8103 (N_8103,N_4137,N_4446);
and U8104 (N_8104,N_1987,N_2291);
nor U8105 (N_8105,N_503,N_1141);
and U8106 (N_8106,N_4220,N_1281);
nor U8107 (N_8107,N_2183,N_2687);
xor U8108 (N_8108,N_416,N_2888);
nor U8109 (N_8109,N_4373,N_3464);
nand U8110 (N_8110,N_502,N_3733);
nor U8111 (N_8111,N_1563,N_38);
or U8112 (N_8112,N_4850,N_2027);
and U8113 (N_8113,N_1936,N_4032);
and U8114 (N_8114,N_2135,N_2324);
nand U8115 (N_8115,N_3698,N_753);
or U8116 (N_8116,N_2365,N_4164);
nand U8117 (N_8117,N_4648,N_3913);
or U8118 (N_8118,N_2056,N_1836);
nor U8119 (N_8119,N_429,N_4161);
nor U8120 (N_8120,N_696,N_1391);
nand U8121 (N_8121,N_710,N_1641);
and U8122 (N_8122,N_1461,N_2845);
nand U8123 (N_8123,N_1074,N_168);
nand U8124 (N_8124,N_356,N_704);
and U8125 (N_8125,N_3947,N_3260);
nor U8126 (N_8126,N_4495,N_683);
and U8127 (N_8127,N_1299,N_974);
xor U8128 (N_8128,N_3472,N_4326);
or U8129 (N_8129,N_418,N_1606);
nor U8130 (N_8130,N_556,N_160);
nor U8131 (N_8131,N_66,N_1685);
nor U8132 (N_8132,N_3474,N_3197);
xnor U8133 (N_8133,N_952,N_4531);
or U8134 (N_8134,N_1605,N_4934);
nand U8135 (N_8135,N_792,N_372);
nor U8136 (N_8136,N_107,N_1889);
or U8137 (N_8137,N_3865,N_1560);
and U8138 (N_8138,N_466,N_1025);
nor U8139 (N_8139,N_438,N_1096);
nand U8140 (N_8140,N_607,N_731);
or U8141 (N_8141,N_1593,N_4100);
xor U8142 (N_8142,N_3881,N_1326);
and U8143 (N_8143,N_4243,N_1626);
or U8144 (N_8144,N_3220,N_493);
xnor U8145 (N_8145,N_2689,N_3870);
nand U8146 (N_8146,N_3495,N_1526);
nor U8147 (N_8147,N_2505,N_4132);
nand U8148 (N_8148,N_4795,N_2136);
xnor U8149 (N_8149,N_4352,N_774);
xnor U8150 (N_8150,N_3320,N_2273);
xor U8151 (N_8151,N_2014,N_154);
or U8152 (N_8152,N_4934,N_4085);
nand U8153 (N_8153,N_3423,N_1717);
or U8154 (N_8154,N_2750,N_3126);
and U8155 (N_8155,N_4288,N_4378);
nand U8156 (N_8156,N_3477,N_1053);
nand U8157 (N_8157,N_3616,N_2022);
xnor U8158 (N_8158,N_1449,N_3298);
and U8159 (N_8159,N_594,N_367);
nor U8160 (N_8160,N_3648,N_1477);
nor U8161 (N_8161,N_2830,N_1783);
xnor U8162 (N_8162,N_1131,N_1123);
nand U8163 (N_8163,N_3765,N_1098);
and U8164 (N_8164,N_2961,N_854);
nand U8165 (N_8165,N_173,N_523);
and U8166 (N_8166,N_4900,N_2388);
nor U8167 (N_8167,N_3801,N_813);
nor U8168 (N_8168,N_1695,N_1779);
xnor U8169 (N_8169,N_4608,N_3518);
nor U8170 (N_8170,N_1311,N_2303);
xnor U8171 (N_8171,N_1597,N_3589);
or U8172 (N_8172,N_1630,N_273);
or U8173 (N_8173,N_556,N_3100);
nor U8174 (N_8174,N_313,N_2415);
xnor U8175 (N_8175,N_963,N_1759);
nand U8176 (N_8176,N_4640,N_3793);
nor U8177 (N_8177,N_694,N_4215);
nand U8178 (N_8178,N_1420,N_2356);
and U8179 (N_8179,N_3624,N_480);
xor U8180 (N_8180,N_3027,N_3285);
or U8181 (N_8181,N_951,N_1990);
xor U8182 (N_8182,N_2546,N_4386);
xor U8183 (N_8183,N_445,N_4730);
nand U8184 (N_8184,N_1077,N_250);
nand U8185 (N_8185,N_4433,N_3542);
or U8186 (N_8186,N_1273,N_3160);
nor U8187 (N_8187,N_1643,N_1431);
nor U8188 (N_8188,N_3715,N_4786);
nor U8189 (N_8189,N_3801,N_3170);
nand U8190 (N_8190,N_1228,N_514);
nor U8191 (N_8191,N_3764,N_4114);
and U8192 (N_8192,N_3898,N_607);
xnor U8193 (N_8193,N_1586,N_4996);
nor U8194 (N_8194,N_3136,N_4185);
and U8195 (N_8195,N_3391,N_4116);
xnor U8196 (N_8196,N_4729,N_3782);
or U8197 (N_8197,N_1762,N_2965);
xnor U8198 (N_8198,N_1773,N_1522);
and U8199 (N_8199,N_250,N_1710);
xor U8200 (N_8200,N_4620,N_3923);
nor U8201 (N_8201,N_4293,N_2069);
and U8202 (N_8202,N_1483,N_1322);
or U8203 (N_8203,N_4422,N_390);
xor U8204 (N_8204,N_1641,N_1961);
or U8205 (N_8205,N_2769,N_2337);
xor U8206 (N_8206,N_4727,N_1174);
or U8207 (N_8207,N_369,N_2259);
xor U8208 (N_8208,N_4114,N_4638);
nand U8209 (N_8209,N_40,N_3825);
and U8210 (N_8210,N_2698,N_3612);
nor U8211 (N_8211,N_2501,N_4272);
nand U8212 (N_8212,N_2773,N_4444);
nor U8213 (N_8213,N_2530,N_2680);
or U8214 (N_8214,N_2398,N_192);
nand U8215 (N_8215,N_4352,N_2906);
xor U8216 (N_8216,N_449,N_2191);
nor U8217 (N_8217,N_669,N_4273);
xor U8218 (N_8218,N_3490,N_1902);
or U8219 (N_8219,N_4533,N_4390);
nor U8220 (N_8220,N_854,N_2340);
nand U8221 (N_8221,N_467,N_3572);
nand U8222 (N_8222,N_2943,N_2227);
and U8223 (N_8223,N_1160,N_1415);
or U8224 (N_8224,N_1653,N_2342);
nor U8225 (N_8225,N_264,N_2020);
nand U8226 (N_8226,N_1901,N_1624);
and U8227 (N_8227,N_930,N_2918);
nor U8228 (N_8228,N_1289,N_2997);
xnor U8229 (N_8229,N_1710,N_4033);
nand U8230 (N_8230,N_1745,N_3780);
nor U8231 (N_8231,N_4179,N_4183);
and U8232 (N_8232,N_2348,N_1530);
nor U8233 (N_8233,N_4993,N_200);
xnor U8234 (N_8234,N_4765,N_1910);
nor U8235 (N_8235,N_4824,N_2856);
xnor U8236 (N_8236,N_3160,N_4173);
xnor U8237 (N_8237,N_3254,N_2264);
nand U8238 (N_8238,N_3056,N_2610);
xnor U8239 (N_8239,N_318,N_3891);
nor U8240 (N_8240,N_601,N_3208);
nand U8241 (N_8241,N_1195,N_4761);
or U8242 (N_8242,N_132,N_2475);
or U8243 (N_8243,N_3215,N_1421);
nor U8244 (N_8244,N_3552,N_1919);
or U8245 (N_8245,N_26,N_1121);
and U8246 (N_8246,N_1149,N_1855);
xor U8247 (N_8247,N_2470,N_3814);
nand U8248 (N_8248,N_3732,N_1946);
and U8249 (N_8249,N_1944,N_93);
nor U8250 (N_8250,N_4643,N_640);
or U8251 (N_8251,N_4258,N_4340);
nand U8252 (N_8252,N_3695,N_383);
or U8253 (N_8253,N_4807,N_1835);
nor U8254 (N_8254,N_2077,N_279);
nor U8255 (N_8255,N_3386,N_3148);
nand U8256 (N_8256,N_1038,N_3);
nand U8257 (N_8257,N_3919,N_4791);
nor U8258 (N_8258,N_3726,N_4860);
and U8259 (N_8259,N_1287,N_2078);
and U8260 (N_8260,N_4528,N_2308);
or U8261 (N_8261,N_1460,N_2090);
nand U8262 (N_8262,N_3612,N_4680);
or U8263 (N_8263,N_659,N_2160);
xor U8264 (N_8264,N_2518,N_3691);
nor U8265 (N_8265,N_492,N_3490);
nor U8266 (N_8266,N_1558,N_2327);
nor U8267 (N_8267,N_4906,N_3818);
nor U8268 (N_8268,N_3237,N_617);
xor U8269 (N_8269,N_3885,N_2108);
and U8270 (N_8270,N_2179,N_4415);
xnor U8271 (N_8271,N_912,N_2989);
nor U8272 (N_8272,N_780,N_4781);
nand U8273 (N_8273,N_2968,N_4747);
and U8274 (N_8274,N_4909,N_2133);
or U8275 (N_8275,N_4329,N_2494);
or U8276 (N_8276,N_2923,N_2572);
or U8277 (N_8277,N_4301,N_2926);
or U8278 (N_8278,N_979,N_2054);
nor U8279 (N_8279,N_4276,N_2093);
or U8280 (N_8280,N_1962,N_4009);
or U8281 (N_8281,N_4542,N_1795);
nor U8282 (N_8282,N_1990,N_4492);
nor U8283 (N_8283,N_208,N_1642);
xor U8284 (N_8284,N_3963,N_676);
nor U8285 (N_8285,N_3586,N_2571);
or U8286 (N_8286,N_2728,N_3378);
nand U8287 (N_8287,N_297,N_1799);
and U8288 (N_8288,N_4343,N_2664);
nor U8289 (N_8289,N_2566,N_1935);
nand U8290 (N_8290,N_3663,N_4954);
xor U8291 (N_8291,N_3340,N_1841);
nor U8292 (N_8292,N_2519,N_4126);
or U8293 (N_8293,N_728,N_76);
or U8294 (N_8294,N_3447,N_3015);
and U8295 (N_8295,N_568,N_1223);
and U8296 (N_8296,N_4925,N_4241);
xnor U8297 (N_8297,N_3914,N_3536);
and U8298 (N_8298,N_2642,N_2212);
nand U8299 (N_8299,N_1287,N_816);
and U8300 (N_8300,N_4037,N_1328);
nand U8301 (N_8301,N_2880,N_293);
and U8302 (N_8302,N_1196,N_4451);
and U8303 (N_8303,N_1983,N_594);
and U8304 (N_8304,N_4153,N_213);
and U8305 (N_8305,N_1526,N_788);
or U8306 (N_8306,N_4900,N_3662);
and U8307 (N_8307,N_1430,N_3484);
and U8308 (N_8308,N_2543,N_4720);
or U8309 (N_8309,N_3656,N_3068);
and U8310 (N_8310,N_1189,N_2874);
and U8311 (N_8311,N_2111,N_3250);
xor U8312 (N_8312,N_4621,N_4633);
and U8313 (N_8313,N_1277,N_219);
nand U8314 (N_8314,N_2486,N_2270);
and U8315 (N_8315,N_1520,N_2357);
nor U8316 (N_8316,N_4389,N_613);
xor U8317 (N_8317,N_4384,N_902);
xnor U8318 (N_8318,N_2847,N_1729);
nor U8319 (N_8319,N_2597,N_331);
and U8320 (N_8320,N_324,N_1683);
or U8321 (N_8321,N_2500,N_4960);
xor U8322 (N_8322,N_1150,N_3472);
xnor U8323 (N_8323,N_3464,N_2525);
or U8324 (N_8324,N_1795,N_819);
nand U8325 (N_8325,N_3307,N_4997);
and U8326 (N_8326,N_3176,N_3647);
nor U8327 (N_8327,N_331,N_4744);
xnor U8328 (N_8328,N_4448,N_590);
nor U8329 (N_8329,N_3228,N_142);
xnor U8330 (N_8330,N_809,N_3374);
or U8331 (N_8331,N_3181,N_3158);
nand U8332 (N_8332,N_1249,N_2242);
nand U8333 (N_8333,N_3788,N_4347);
nor U8334 (N_8334,N_3574,N_1872);
and U8335 (N_8335,N_3759,N_3010);
nor U8336 (N_8336,N_836,N_1632);
or U8337 (N_8337,N_3771,N_4063);
nor U8338 (N_8338,N_4262,N_3620);
nand U8339 (N_8339,N_4819,N_2770);
and U8340 (N_8340,N_1059,N_198);
nand U8341 (N_8341,N_2254,N_2475);
nor U8342 (N_8342,N_1732,N_387);
nor U8343 (N_8343,N_590,N_562);
nor U8344 (N_8344,N_3915,N_4714);
and U8345 (N_8345,N_2210,N_649);
or U8346 (N_8346,N_3416,N_4078);
xnor U8347 (N_8347,N_2725,N_1633);
nand U8348 (N_8348,N_952,N_1170);
nor U8349 (N_8349,N_2258,N_4947);
or U8350 (N_8350,N_4619,N_405);
nand U8351 (N_8351,N_3502,N_2487);
or U8352 (N_8352,N_4683,N_1642);
nand U8353 (N_8353,N_354,N_2003);
xnor U8354 (N_8354,N_4003,N_3250);
and U8355 (N_8355,N_2874,N_3632);
nor U8356 (N_8356,N_3069,N_3536);
nand U8357 (N_8357,N_2463,N_4967);
xor U8358 (N_8358,N_1284,N_4216);
xor U8359 (N_8359,N_4335,N_2023);
xor U8360 (N_8360,N_1357,N_4554);
xor U8361 (N_8361,N_1630,N_1278);
or U8362 (N_8362,N_2245,N_2609);
xor U8363 (N_8363,N_4396,N_3318);
or U8364 (N_8364,N_3621,N_1079);
and U8365 (N_8365,N_492,N_3676);
nor U8366 (N_8366,N_4052,N_3420);
or U8367 (N_8367,N_2833,N_217);
and U8368 (N_8368,N_4845,N_23);
or U8369 (N_8369,N_2333,N_2630);
or U8370 (N_8370,N_1473,N_404);
xor U8371 (N_8371,N_151,N_4263);
and U8372 (N_8372,N_1894,N_2746);
or U8373 (N_8373,N_494,N_4432);
and U8374 (N_8374,N_499,N_4414);
nand U8375 (N_8375,N_838,N_688);
xnor U8376 (N_8376,N_1981,N_535);
nor U8377 (N_8377,N_1606,N_2746);
nand U8378 (N_8378,N_797,N_81);
and U8379 (N_8379,N_4373,N_4122);
nor U8380 (N_8380,N_4392,N_1550);
nor U8381 (N_8381,N_4925,N_936);
nor U8382 (N_8382,N_1510,N_2635);
and U8383 (N_8383,N_1583,N_4562);
and U8384 (N_8384,N_1864,N_3128);
nand U8385 (N_8385,N_2341,N_2769);
nand U8386 (N_8386,N_2468,N_4494);
nor U8387 (N_8387,N_2686,N_1122);
nor U8388 (N_8388,N_3723,N_4107);
nand U8389 (N_8389,N_1113,N_3438);
nor U8390 (N_8390,N_1540,N_827);
nand U8391 (N_8391,N_4262,N_326);
or U8392 (N_8392,N_3588,N_1142);
xnor U8393 (N_8393,N_2874,N_2734);
xor U8394 (N_8394,N_2610,N_1265);
nand U8395 (N_8395,N_4663,N_4859);
or U8396 (N_8396,N_1379,N_1754);
xor U8397 (N_8397,N_3186,N_1237);
nand U8398 (N_8398,N_9,N_1772);
nand U8399 (N_8399,N_4949,N_3501);
and U8400 (N_8400,N_4854,N_4822);
nor U8401 (N_8401,N_468,N_2128);
nor U8402 (N_8402,N_476,N_3506);
and U8403 (N_8403,N_2150,N_1041);
nand U8404 (N_8404,N_2145,N_3069);
or U8405 (N_8405,N_4866,N_2804);
xor U8406 (N_8406,N_3271,N_1892);
nand U8407 (N_8407,N_4759,N_4709);
nor U8408 (N_8408,N_417,N_4913);
or U8409 (N_8409,N_3316,N_4604);
and U8410 (N_8410,N_2728,N_4964);
nand U8411 (N_8411,N_979,N_633);
nand U8412 (N_8412,N_906,N_3898);
nor U8413 (N_8413,N_876,N_56);
or U8414 (N_8414,N_3778,N_1276);
nand U8415 (N_8415,N_539,N_2344);
and U8416 (N_8416,N_2681,N_2902);
or U8417 (N_8417,N_3475,N_2507);
nand U8418 (N_8418,N_3167,N_2389);
nor U8419 (N_8419,N_4223,N_1504);
nor U8420 (N_8420,N_4981,N_2370);
or U8421 (N_8421,N_956,N_4115);
nor U8422 (N_8422,N_719,N_1153);
and U8423 (N_8423,N_2175,N_1495);
nand U8424 (N_8424,N_4723,N_939);
nor U8425 (N_8425,N_2469,N_4066);
xor U8426 (N_8426,N_507,N_3060);
xnor U8427 (N_8427,N_3543,N_4547);
nor U8428 (N_8428,N_4560,N_3842);
or U8429 (N_8429,N_1336,N_3937);
xor U8430 (N_8430,N_2349,N_2552);
xor U8431 (N_8431,N_3850,N_119);
nand U8432 (N_8432,N_2214,N_1238);
nand U8433 (N_8433,N_715,N_1940);
nor U8434 (N_8434,N_211,N_4799);
nor U8435 (N_8435,N_4814,N_176);
or U8436 (N_8436,N_1600,N_833);
xor U8437 (N_8437,N_2926,N_2501);
or U8438 (N_8438,N_2039,N_2617);
nand U8439 (N_8439,N_767,N_3578);
or U8440 (N_8440,N_2404,N_2083);
or U8441 (N_8441,N_543,N_2326);
or U8442 (N_8442,N_3479,N_1450);
nand U8443 (N_8443,N_4825,N_1459);
or U8444 (N_8444,N_3195,N_2679);
nand U8445 (N_8445,N_1030,N_1319);
and U8446 (N_8446,N_4800,N_2);
nor U8447 (N_8447,N_4896,N_4148);
nand U8448 (N_8448,N_4759,N_2993);
nor U8449 (N_8449,N_3661,N_4056);
xor U8450 (N_8450,N_2149,N_4312);
xnor U8451 (N_8451,N_440,N_4033);
nand U8452 (N_8452,N_2730,N_2964);
xnor U8453 (N_8453,N_299,N_4164);
nand U8454 (N_8454,N_4282,N_3460);
nor U8455 (N_8455,N_1346,N_1026);
and U8456 (N_8456,N_1320,N_272);
xnor U8457 (N_8457,N_2319,N_3251);
and U8458 (N_8458,N_100,N_16);
and U8459 (N_8459,N_4846,N_3581);
and U8460 (N_8460,N_2287,N_241);
and U8461 (N_8461,N_4186,N_3334);
and U8462 (N_8462,N_4368,N_1988);
xnor U8463 (N_8463,N_4606,N_1313);
or U8464 (N_8464,N_4398,N_3189);
xnor U8465 (N_8465,N_1033,N_3745);
or U8466 (N_8466,N_4647,N_2884);
or U8467 (N_8467,N_170,N_2112);
and U8468 (N_8468,N_2798,N_365);
nand U8469 (N_8469,N_749,N_906);
or U8470 (N_8470,N_2185,N_1912);
or U8471 (N_8471,N_271,N_847);
xor U8472 (N_8472,N_3755,N_1152);
nor U8473 (N_8473,N_2354,N_2271);
and U8474 (N_8474,N_1859,N_589);
nor U8475 (N_8475,N_3545,N_4115);
nor U8476 (N_8476,N_56,N_787);
xnor U8477 (N_8477,N_169,N_3906);
xnor U8478 (N_8478,N_4944,N_184);
xor U8479 (N_8479,N_2599,N_4193);
or U8480 (N_8480,N_1593,N_482);
xor U8481 (N_8481,N_1741,N_1009);
xnor U8482 (N_8482,N_4345,N_2018);
or U8483 (N_8483,N_4746,N_2470);
xnor U8484 (N_8484,N_2078,N_4406);
and U8485 (N_8485,N_832,N_1269);
or U8486 (N_8486,N_1438,N_1255);
xnor U8487 (N_8487,N_392,N_1166);
xor U8488 (N_8488,N_4463,N_4113);
nand U8489 (N_8489,N_4359,N_4609);
nor U8490 (N_8490,N_2809,N_680);
and U8491 (N_8491,N_4088,N_3609);
nor U8492 (N_8492,N_478,N_4476);
xor U8493 (N_8493,N_1586,N_2748);
and U8494 (N_8494,N_526,N_3714);
and U8495 (N_8495,N_1262,N_4571);
nor U8496 (N_8496,N_2025,N_4638);
and U8497 (N_8497,N_2203,N_2778);
or U8498 (N_8498,N_1114,N_4163);
xor U8499 (N_8499,N_2347,N_4419);
or U8500 (N_8500,N_171,N_1656);
or U8501 (N_8501,N_781,N_134);
nor U8502 (N_8502,N_4030,N_4816);
and U8503 (N_8503,N_2978,N_4894);
and U8504 (N_8504,N_4199,N_2472);
nor U8505 (N_8505,N_895,N_363);
or U8506 (N_8506,N_4066,N_1866);
and U8507 (N_8507,N_1693,N_3379);
and U8508 (N_8508,N_4316,N_185);
nor U8509 (N_8509,N_1372,N_2046);
nand U8510 (N_8510,N_1549,N_4480);
xor U8511 (N_8511,N_2847,N_862);
xor U8512 (N_8512,N_1108,N_4493);
and U8513 (N_8513,N_4093,N_4548);
nand U8514 (N_8514,N_701,N_2556);
nand U8515 (N_8515,N_1782,N_973);
xnor U8516 (N_8516,N_4172,N_2196);
xor U8517 (N_8517,N_2147,N_2067);
nor U8518 (N_8518,N_4825,N_1094);
nand U8519 (N_8519,N_361,N_2919);
xor U8520 (N_8520,N_598,N_421);
and U8521 (N_8521,N_3270,N_483);
nor U8522 (N_8522,N_3376,N_2820);
nand U8523 (N_8523,N_4206,N_1387);
or U8524 (N_8524,N_986,N_3450);
xnor U8525 (N_8525,N_4650,N_4436);
and U8526 (N_8526,N_2496,N_949);
or U8527 (N_8527,N_632,N_2039);
or U8528 (N_8528,N_4682,N_3825);
or U8529 (N_8529,N_3428,N_2394);
and U8530 (N_8530,N_274,N_4138);
and U8531 (N_8531,N_1671,N_2609);
nor U8532 (N_8532,N_3940,N_4026);
xnor U8533 (N_8533,N_4514,N_3875);
nor U8534 (N_8534,N_491,N_4068);
xor U8535 (N_8535,N_3662,N_2648);
and U8536 (N_8536,N_4376,N_4292);
nand U8537 (N_8537,N_4239,N_3781);
nand U8538 (N_8538,N_2663,N_4856);
or U8539 (N_8539,N_1225,N_4408);
nor U8540 (N_8540,N_576,N_2545);
nand U8541 (N_8541,N_4770,N_1619);
nand U8542 (N_8542,N_3847,N_4738);
xnor U8543 (N_8543,N_4357,N_4373);
xnor U8544 (N_8544,N_4938,N_796);
and U8545 (N_8545,N_1506,N_1388);
and U8546 (N_8546,N_1064,N_2962);
or U8547 (N_8547,N_745,N_3665);
nor U8548 (N_8548,N_4239,N_1601);
nor U8549 (N_8549,N_253,N_382);
and U8550 (N_8550,N_2231,N_3047);
xor U8551 (N_8551,N_4539,N_3709);
xnor U8552 (N_8552,N_1760,N_4429);
nand U8553 (N_8553,N_4383,N_607);
and U8554 (N_8554,N_3877,N_2981);
and U8555 (N_8555,N_4958,N_3847);
nor U8556 (N_8556,N_1050,N_3976);
nor U8557 (N_8557,N_2870,N_4694);
or U8558 (N_8558,N_210,N_1285);
and U8559 (N_8559,N_2159,N_4149);
nand U8560 (N_8560,N_2072,N_1346);
or U8561 (N_8561,N_3339,N_2232);
xor U8562 (N_8562,N_1683,N_1577);
or U8563 (N_8563,N_4490,N_634);
or U8564 (N_8564,N_4587,N_3119);
and U8565 (N_8565,N_2002,N_2119);
and U8566 (N_8566,N_1122,N_1775);
xor U8567 (N_8567,N_2404,N_1173);
and U8568 (N_8568,N_3887,N_4305);
nand U8569 (N_8569,N_4433,N_3828);
nor U8570 (N_8570,N_1017,N_4674);
or U8571 (N_8571,N_4211,N_2831);
nand U8572 (N_8572,N_3819,N_2249);
nand U8573 (N_8573,N_3482,N_1493);
xnor U8574 (N_8574,N_3562,N_816);
and U8575 (N_8575,N_1910,N_615);
nand U8576 (N_8576,N_2160,N_1599);
or U8577 (N_8577,N_2958,N_3045);
or U8578 (N_8578,N_3844,N_2853);
or U8579 (N_8579,N_4813,N_179);
nand U8580 (N_8580,N_3821,N_2770);
and U8581 (N_8581,N_4168,N_2052);
or U8582 (N_8582,N_330,N_3595);
or U8583 (N_8583,N_1516,N_4929);
nor U8584 (N_8584,N_3370,N_732);
or U8585 (N_8585,N_822,N_4038);
and U8586 (N_8586,N_2363,N_2391);
and U8587 (N_8587,N_2311,N_4659);
xnor U8588 (N_8588,N_3960,N_2106);
and U8589 (N_8589,N_4752,N_751);
and U8590 (N_8590,N_3400,N_1398);
xor U8591 (N_8591,N_2268,N_4364);
nor U8592 (N_8592,N_4857,N_3147);
nor U8593 (N_8593,N_2547,N_1675);
and U8594 (N_8594,N_4134,N_2119);
xnor U8595 (N_8595,N_2145,N_4603);
xnor U8596 (N_8596,N_1114,N_135);
nand U8597 (N_8597,N_1793,N_3623);
and U8598 (N_8598,N_1162,N_2319);
or U8599 (N_8599,N_1639,N_3854);
xnor U8600 (N_8600,N_3474,N_385);
or U8601 (N_8601,N_2420,N_161);
nand U8602 (N_8602,N_2177,N_4973);
nor U8603 (N_8603,N_4263,N_4955);
xnor U8604 (N_8604,N_396,N_4407);
xor U8605 (N_8605,N_3002,N_3550);
nor U8606 (N_8606,N_1015,N_1103);
nand U8607 (N_8607,N_4886,N_3180);
nand U8608 (N_8608,N_4892,N_2793);
nand U8609 (N_8609,N_2930,N_3047);
nand U8610 (N_8610,N_3233,N_1863);
nor U8611 (N_8611,N_1430,N_930);
and U8612 (N_8612,N_1651,N_1629);
and U8613 (N_8613,N_762,N_334);
xor U8614 (N_8614,N_258,N_2691);
nand U8615 (N_8615,N_4485,N_1048);
nand U8616 (N_8616,N_1703,N_1768);
nor U8617 (N_8617,N_4733,N_3435);
nand U8618 (N_8618,N_1141,N_446);
and U8619 (N_8619,N_802,N_1424);
nor U8620 (N_8620,N_1398,N_4079);
nand U8621 (N_8621,N_1126,N_4737);
xor U8622 (N_8622,N_429,N_2032);
xnor U8623 (N_8623,N_914,N_1796);
xor U8624 (N_8624,N_1876,N_1995);
or U8625 (N_8625,N_2251,N_3703);
nor U8626 (N_8626,N_1092,N_1729);
nand U8627 (N_8627,N_1914,N_1629);
xnor U8628 (N_8628,N_1420,N_2850);
nor U8629 (N_8629,N_546,N_4471);
or U8630 (N_8630,N_151,N_2266);
xnor U8631 (N_8631,N_883,N_2779);
and U8632 (N_8632,N_3284,N_172);
or U8633 (N_8633,N_617,N_3683);
nor U8634 (N_8634,N_4124,N_3660);
nand U8635 (N_8635,N_3522,N_2982);
nor U8636 (N_8636,N_2678,N_1509);
nor U8637 (N_8637,N_1509,N_87);
nor U8638 (N_8638,N_134,N_4204);
nor U8639 (N_8639,N_2285,N_3160);
or U8640 (N_8640,N_4488,N_2458);
nor U8641 (N_8641,N_1413,N_4963);
xor U8642 (N_8642,N_3251,N_1519);
xor U8643 (N_8643,N_4536,N_2496);
nand U8644 (N_8644,N_3062,N_3157);
or U8645 (N_8645,N_1681,N_228);
nand U8646 (N_8646,N_782,N_197);
nor U8647 (N_8647,N_2450,N_2095);
and U8648 (N_8648,N_3940,N_3800);
xor U8649 (N_8649,N_3753,N_1963);
nor U8650 (N_8650,N_2952,N_379);
nand U8651 (N_8651,N_3273,N_98);
or U8652 (N_8652,N_211,N_1967);
nor U8653 (N_8653,N_3362,N_3363);
and U8654 (N_8654,N_4022,N_3667);
nor U8655 (N_8655,N_1802,N_1349);
or U8656 (N_8656,N_908,N_166);
and U8657 (N_8657,N_3144,N_4418);
and U8658 (N_8658,N_3263,N_2801);
nand U8659 (N_8659,N_2725,N_2475);
xnor U8660 (N_8660,N_2404,N_2517);
nor U8661 (N_8661,N_4205,N_4847);
xnor U8662 (N_8662,N_644,N_1148);
and U8663 (N_8663,N_4184,N_2308);
nand U8664 (N_8664,N_2190,N_2497);
xnor U8665 (N_8665,N_31,N_4054);
and U8666 (N_8666,N_4801,N_952);
and U8667 (N_8667,N_2888,N_2643);
nor U8668 (N_8668,N_4197,N_3624);
xnor U8669 (N_8669,N_3985,N_1320);
nor U8670 (N_8670,N_4080,N_1601);
and U8671 (N_8671,N_2015,N_3107);
xnor U8672 (N_8672,N_2368,N_3203);
nor U8673 (N_8673,N_1855,N_3812);
xor U8674 (N_8674,N_3399,N_3366);
nor U8675 (N_8675,N_513,N_3378);
or U8676 (N_8676,N_1656,N_2461);
or U8677 (N_8677,N_308,N_1643);
and U8678 (N_8678,N_2872,N_3586);
nor U8679 (N_8679,N_4172,N_4156);
nor U8680 (N_8680,N_718,N_635);
and U8681 (N_8681,N_2165,N_839);
or U8682 (N_8682,N_4543,N_2644);
xor U8683 (N_8683,N_2195,N_3523);
xor U8684 (N_8684,N_975,N_2032);
or U8685 (N_8685,N_2125,N_3380);
or U8686 (N_8686,N_1398,N_3410);
and U8687 (N_8687,N_3050,N_919);
or U8688 (N_8688,N_4853,N_4111);
xnor U8689 (N_8689,N_4734,N_3451);
nor U8690 (N_8690,N_3932,N_2585);
and U8691 (N_8691,N_229,N_3671);
nand U8692 (N_8692,N_3892,N_4259);
and U8693 (N_8693,N_3545,N_754);
xor U8694 (N_8694,N_2576,N_93);
or U8695 (N_8695,N_1734,N_2811);
xor U8696 (N_8696,N_2481,N_1835);
xor U8697 (N_8697,N_2034,N_1059);
nor U8698 (N_8698,N_4022,N_2059);
and U8699 (N_8699,N_1172,N_3691);
nand U8700 (N_8700,N_2938,N_409);
xor U8701 (N_8701,N_1753,N_4891);
xor U8702 (N_8702,N_2730,N_4826);
xnor U8703 (N_8703,N_1269,N_4232);
and U8704 (N_8704,N_369,N_2610);
xnor U8705 (N_8705,N_895,N_3501);
nand U8706 (N_8706,N_1,N_2801);
and U8707 (N_8707,N_4223,N_80);
or U8708 (N_8708,N_3428,N_1077);
nand U8709 (N_8709,N_2386,N_4211);
or U8710 (N_8710,N_2767,N_2660);
xor U8711 (N_8711,N_4756,N_2798);
xor U8712 (N_8712,N_2871,N_1619);
xor U8713 (N_8713,N_433,N_3764);
or U8714 (N_8714,N_4421,N_4622);
xor U8715 (N_8715,N_734,N_3559);
nand U8716 (N_8716,N_4921,N_4681);
or U8717 (N_8717,N_4273,N_2360);
nor U8718 (N_8718,N_3212,N_211);
nand U8719 (N_8719,N_1735,N_826);
nand U8720 (N_8720,N_85,N_4884);
or U8721 (N_8721,N_3373,N_2070);
nand U8722 (N_8722,N_141,N_619);
xor U8723 (N_8723,N_825,N_3714);
nor U8724 (N_8724,N_4578,N_858);
nor U8725 (N_8725,N_4141,N_4308);
and U8726 (N_8726,N_4482,N_2747);
and U8727 (N_8727,N_1085,N_3246);
xnor U8728 (N_8728,N_2089,N_2258);
or U8729 (N_8729,N_709,N_4123);
and U8730 (N_8730,N_4777,N_267);
xnor U8731 (N_8731,N_3546,N_4555);
nor U8732 (N_8732,N_4802,N_3967);
nor U8733 (N_8733,N_2063,N_3660);
xnor U8734 (N_8734,N_94,N_4692);
xnor U8735 (N_8735,N_409,N_4393);
nor U8736 (N_8736,N_468,N_1567);
nand U8737 (N_8737,N_4645,N_226);
or U8738 (N_8738,N_1130,N_3161);
xor U8739 (N_8739,N_185,N_707);
nor U8740 (N_8740,N_3736,N_3277);
xor U8741 (N_8741,N_854,N_2999);
nor U8742 (N_8742,N_2341,N_2111);
nor U8743 (N_8743,N_3566,N_4472);
and U8744 (N_8744,N_4828,N_2670);
nand U8745 (N_8745,N_1446,N_4629);
xnor U8746 (N_8746,N_4965,N_1602);
and U8747 (N_8747,N_2693,N_3392);
and U8748 (N_8748,N_2328,N_1279);
nand U8749 (N_8749,N_1815,N_2694);
nor U8750 (N_8750,N_887,N_2640);
or U8751 (N_8751,N_1795,N_4239);
xnor U8752 (N_8752,N_949,N_1770);
and U8753 (N_8753,N_1116,N_3235);
or U8754 (N_8754,N_1329,N_148);
nor U8755 (N_8755,N_3904,N_255);
or U8756 (N_8756,N_1895,N_4232);
xnor U8757 (N_8757,N_2147,N_349);
nor U8758 (N_8758,N_1742,N_2288);
xor U8759 (N_8759,N_3309,N_3368);
xor U8760 (N_8760,N_2489,N_2023);
or U8761 (N_8761,N_1393,N_980);
nor U8762 (N_8762,N_3386,N_4332);
nand U8763 (N_8763,N_3155,N_4538);
or U8764 (N_8764,N_4072,N_2638);
nor U8765 (N_8765,N_4164,N_4559);
and U8766 (N_8766,N_339,N_1576);
xor U8767 (N_8767,N_1528,N_1211);
xor U8768 (N_8768,N_1856,N_3428);
xor U8769 (N_8769,N_2161,N_3429);
nor U8770 (N_8770,N_3530,N_1379);
nor U8771 (N_8771,N_1317,N_3461);
and U8772 (N_8772,N_4380,N_2621);
or U8773 (N_8773,N_2821,N_2033);
xnor U8774 (N_8774,N_4364,N_367);
and U8775 (N_8775,N_4940,N_4215);
and U8776 (N_8776,N_4135,N_3191);
nand U8777 (N_8777,N_1489,N_1248);
nor U8778 (N_8778,N_565,N_1337);
nor U8779 (N_8779,N_4785,N_2273);
and U8780 (N_8780,N_2396,N_1392);
or U8781 (N_8781,N_68,N_1391);
xnor U8782 (N_8782,N_2155,N_2554);
and U8783 (N_8783,N_2256,N_3707);
nand U8784 (N_8784,N_4921,N_366);
and U8785 (N_8785,N_4945,N_479);
nor U8786 (N_8786,N_3791,N_4975);
or U8787 (N_8787,N_952,N_2972);
nand U8788 (N_8788,N_3379,N_4230);
nor U8789 (N_8789,N_3329,N_952);
or U8790 (N_8790,N_533,N_2950);
or U8791 (N_8791,N_2743,N_3262);
or U8792 (N_8792,N_3999,N_3718);
and U8793 (N_8793,N_39,N_2185);
nor U8794 (N_8794,N_3701,N_1897);
nor U8795 (N_8795,N_1251,N_294);
nor U8796 (N_8796,N_2886,N_2992);
or U8797 (N_8797,N_4655,N_4264);
xnor U8798 (N_8798,N_3540,N_4383);
nor U8799 (N_8799,N_4769,N_421);
and U8800 (N_8800,N_4555,N_3882);
nor U8801 (N_8801,N_2295,N_3881);
xor U8802 (N_8802,N_1573,N_1251);
nor U8803 (N_8803,N_3855,N_3259);
nor U8804 (N_8804,N_3804,N_1868);
xnor U8805 (N_8805,N_2294,N_390);
and U8806 (N_8806,N_1939,N_3565);
nand U8807 (N_8807,N_3616,N_2231);
and U8808 (N_8808,N_1323,N_3545);
nor U8809 (N_8809,N_1025,N_591);
xnor U8810 (N_8810,N_2916,N_2716);
nand U8811 (N_8811,N_180,N_4513);
xnor U8812 (N_8812,N_2162,N_3900);
nand U8813 (N_8813,N_4288,N_157);
xnor U8814 (N_8814,N_4576,N_4248);
xnor U8815 (N_8815,N_2751,N_3276);
nor U8816 (N_8816,N_3694,N_2341);
nor U8817 (N_8817,N_3971,N_3968);
xor U8818 (N_8818,N_605,N_209);
nor U8819 (N_8819,N_2817,N_3104);
and U8820 (N_8820,N_2599,N_4671);
nand U8821 (N_8821,N_2026,N_1125);
and U8822 (N_8822,N_4311,N_2314);
or U8823 (N_8823,N_4652,N_3889);
nand U8824 (N_8824,N_1116,N_931);
nor U8825 (N_8825,N_1236,N_2578);
nand U8826 (N_8826,N_2877,N_4104);
xnor U8827 (N_8827,N_562,N_4376);
nor U8828 (N_8828,N_1208,N_703);
and U8829 (N_8829,N_2222,N_2060);
xnor U8830 (N_8830,N_369,N_4030);
and U8831 (N_8831,N_3028,N_4102);
and U8832 (N_8832,N_2849,N_1482);
nor U8833 (N_8833,N_3349,N_3778);
nand U8834 (N_8834,N_710,N_4808);
or U8835 (N_8835,N_1496,N_1558);
or U8836 (N_8836,N_2725,N_3107);
nor U8837 (N_8837,N_3334,N_3896);
xnor U8838 (N_8838,N_2306,N_3609);
or U8839 (N_8839,N_2115,N_3592);
or U8840 (N_8840,N_4706,N_1032);
or U8841 (N_8841,N_2858,N_1842);
or U8842 (N_8842,N_3065,N_1770);
or U8843 (N_8843,N_870,N_1899);
nand U8844 (N_8844,N_3057,N_1313);
xor U8845 (N_8845,N_2536,N_2642);
or U8846 (N_8846,N_2698,N_2838);
xor U8847 (N_8847,N_1856,N_4091);
nor U8848 (N_8848,N_3326,N_2951);
or U8849 (N_8849,N_3972,N_1457);
and U8850 (N_8850,N_4097,N_4281);
and U8851 (N_8851,N_1394,N_4942);
nor U8852 (N_8852,N_1750,N_3387);
nand U8853 (N_8853,N_3009,N_4570);
nand U8854 (N_8854,N_3731,N_347);
or U8855 (N_8855,N_2375,N_4101);
nor U8856 (N_8856,N_3921,N_4655);
nand U8857 (N_8857,N_3562,N_3922);
and U8858 (N_8858,N_3008,N_1880);
or U8859 (N_8859,N_2604,N_100);
and U8860 (N_8860,N_3884,N_3853);
or U8861 (N_8861,N_3855,N_2876);
and U8862 (N_8862,N_2059,N_1660);
nor U8863 (N_8863,N_1860,N_2875);
xor U8864 (N_8864,N_4763,N_4275);
and U8865 (N_8865,N_4539,N_2467);
nor U8866 (N_8866,N_4329,N_544);
nand U8867 (N_8867,N_1382,N_493);
and U8868 (N_8868,N_3824,N_4247);
nand U8869 (N_8869,N_1415,N_317);
xnor U8870 (N_8870,N_4657,N_3203);
or U8871 (N_8871,N_1690,N_848);
xnor U8872 (N_8872,N_4496,N_745);
nand U8873 (N_8873,N_290,N_2001);
nand U8874 (N_8874,N_2140,N_3024);
and U8875 (N_8875,N_483,N_3006);
nor U8876 (N_8876,N_395,N_3650);
nand U8877 (N_8877,N_1668,N_1219);
and U8878 (N_8878,N_4943,N_1238);
or U8879 (N_8879,N_2787,N_271);
nand U8880 (N_8880,N_56,N_94);
nand U8881 (N_8881,N_4682,N_2204);
nor U8882 (N_8882,N_3470,N_4848);
xnor U8883 (N_8883,N_4326,N_2858);
nor U8884 (N_8884,N_3707,N_3449);
xnor U8885 (N_8885,N_4075,N_935);
xor U8886 (N_8886,N_1320,N_2448);
xnor U8887 (N_8887,N_4813,N_323);
nand U8888 (N_8888,N_2052,N_2551);
and U8889 (N_8889,N_3460,N_227);
xor U8890 (N_8890,N_1481,N_2148);
or U8891 (N_8891,N_4394,N_4918);
xnor U8892 (N_8892,N_42,N_4054);
nor U8893 (N_8893,N_4675,N_3309);
xnor U8894 (N_8894,N_575,N_4178);
or U8895 (N_8895,N_3578,N_3378);
and U8896 (N_8896,N_4167,N_2046);
and U8897 (N_8897,N_17,N_2573);
xnor U8898 (N_8898,N_2735,N_241);
and U8899 (N_8899,N_3684,N_360);
xor U8900 (N_8900,N_3880,N_838);
and U8901 (N_8901,N_4227,N_4709);
xor U8902 (N_8902,N_1834,N_2120);
xor U8903 (N_8903,N_3008,N_1750);
nand U8904 (N_8904,N_4251,N_2561);
nand U8905 (N_8905,N_1846,N_4244);
or U8906 (N_8906,N_1394,N_3861);
or U8907 (N_8907,N_4215,N_1819);
xnor U8908 (N_8908,N_1438,N_2300);
xnor U8909 (N_8909,N_721,N_1495);
xnor U8910 (N_8910,N_4281,N_4856);
nor U8911 (N_8911,N_4780,N_2920);
nand U8912 (N_8912,N_4597,N_549);
and U8913 (N_8913,N_2389,N_4052);
xor U8914 (N_8914,N_4388,N_2814);
or U8915 (N_8915,N_3843,N_1527);
and U8916 (N_8916,N_3374,N_1743);
or U8917 (N_8917,N_4510,N_796);
or U8918 (N_8918,N_501,N_430);
nor U8919 (N_8919,N_2663,N_2468);
xor U8920 (N_8920,N_4203,N_30);
nor U8921 (N_8921,N_669,N_4104);
or U8922 (N_8922,N_108,N_3282);
and U8923 (N_8923,N_3723,N_3879);
nor U8924 (N_8924,N_3390,N_1565);
or U8925 (N_8925,N_2631,N_284);
xnor U8926 (N_8926,N_2775,N_4570);
or U8927 (N_8927,N_3537,N_4105);
nand U8928 (N_8928,N_204,N_4963);
nand U8929 (N_8929,N_2665,N_389);
nand U8930 (N_8930,N_2964,N_2766);
and U8931 (N_8931,N_727,N_46);
and U8932 (N_8932,N_3864,N_3397);
or U8933 (N_8933,N_4834,N_4253);
nand U8934 (N_8934,N_3710,N_407);
or U8935 (N_8935,N_1308,N_693);
nor U8936 (N_8936,N_670,N_627);
nand U8937 (N_8937,N_3921,N_320);
nand U8938 (N_8938,N_2264,N_105);
nand U8939 (N_8939,N_3297,N_4873);
xor U8940 (N_8940,N_761,N_1099);
or U8941 (N_8941,N_933,N_2452);
or U8942 (N_8942,N_2422,N_173);
or U8943 (N_8943,N_1236,N_2070);
nor U8944 (N_8944,N_4997,N_4331);
or U8945 (N_8945,N_2516,N_4138);
or U8946 (N_8946,N_4040,N_4610);
nand U8947 (N_8947,N_4919,N_1193);
or U8948 (N_8948,N_4275,N_3673);
xnor U8949 (N_8949,N_4115,N_867);
xor U8950 (N_8950,N_3250,N_3116);
nor U8951 (N_8951,N_3662,N_3663);
and U8952 (N_8952,N_4039,N_1345);
nand U8953 (N_8953,N_3073,N_2979);
nor U8954 (N_8954,N_309,N_1967);
or U8955 (N_8955,N_1900,N_2794);
nand U8956 (N_8956,N_3887,N_2708);
nor U8957 (N_8957,N_3981,N_2309);
and U8958 (N_8958,N_1989,N_3127);
xor U8959 (N_8959,N_2006,N_4090);
nor U8960 (N_8960,N_1507,N_3193);
xor U8961 (N_8961,N_2475,N_337);
and U8962 (N_8962,N_2271,N_3839);
or U8963 (N_8963,N_1015,N_1380);
xor U8964 (N_8964,N_2031,N_2437);
xnor U8965 (N_8965,N_13,N_1908);
nand U8966 (N_8966,N_4075,N_1161);
and U8967 (N_8967,N_1773,N_1857);
and U8968 (N_8968,N_3945,N_3741);
or U8969 (N_8969,N_447,N_1747);
nor U8970 (N_8970,N_3371,N_4037);
and U8971 (N_8971,N_1623,N_506);
nand U8972 (N_8972,N_1435,N_2960);
xor U8973 (N_8973,N_3988,N_298);
nor U8974 (N_8974,N_471,N_3969);
nor U8975 (N_8975,N_2458,N_3510);
and U8976 (N_8976,N_3684,N_1324);
nand U8977 (N_8977,N_1898,N_563);
xnor U8978 (N_8978,N_4136,N_2626);
nor U8979 (N_8979,N_352,N_3115);
nand U8980 (N_8980,N_1819,N_3402);
or U8981 (N_8981,N_1056,N_1900);
xnor U8982 (N_8982,N_2071,N_1951);
or U8983 (N_8983,N_697,N_416);
nand U8984 (N_8984,N_3391,N_4475);
and U8985 (N_8985,N_4612,N_1001);
nor U8986 (N_8986,N_1993,N_3056);
nor U8987 (N_8987,N_201,N_317);
nand U8988 (N_8988,N_3662,N_2349);
and U8989 (N_8989,N_3152,N_2867);
xnor U8990 (N_8990,N_2325,N_2418);
nand U8991 (N_8991,N_1231,N_695);
nor U8992 (N_8992,N_492,N_661);
nor U8993 (N_8993,N_2362,N_2891);
nor U8994 (N_8994,N_4747,N_1354);
nand U8995 (N_8995,N_876,N_1973);
nand U8996 (N_8996,N_3816,N_49);
nor U8997 (N_8997,N_2266,N_3631);
nor U8998 (N_8998,N_477,N_137);
and U8999 (N_8999,N_3376,N_4559);
nand U9000 (N_9000,N_2955,N_1754);
xor U9001 (N_9001,N_1796,N_472);
or U9002 (N_9002,N_2007,N_2784);
or U9003 (N_9003,N_1313,N_4864);
nor U9004 (N_9004,N_2870,N_837);
xor U9005 (N_9005,N_2442,N_3939);
nand U9006 (N_9006,N_2049,N_3768);
nand U9007 (N_9007,N_4029,N_4045);
and U9008 (N_9008,N_469,N_1102);
xor U9009 (N_9009,N_2666,N_3510);
nor U9010 (N_9010,N_1454,N_358);
and U9011 (N_9011,N_4255,N_2899);
xor U9012 (N_9012,N_3954,N_3823);
or U9013 (N_9013,N_195,N_2816);
and U9014 (N_9014,N_1125,N_3650);
xor U9015 (N_9015,N_1369,N_3356);
and U9016 (N_9016,N_3964,N_311);
nand U9017 (N_9017,N_4736,N_784);
or U9018 (N_9018,N_1241,N_2958);
and U9019 (N_9019,N_974,N_3558);
nor U9020 (N_9020,N_2770,N_4204);
xnor U9021 (N_9021,N_923,N_2791);
nand U9022 (N_9022,N_4792,N_1512);
or U9023 (N_9023,N_3925,N_2578);
xor U9024 (N_9024,N_677,N_1517);
and U9025 (N_9025,N_2632,N_681);
nand U9026 (N_9026,N_1942,N_1584);
nand U9027 (N_9027,N_2000,N_1948);
nor U9028 (N_9028,N_3340,N_3194);
xor U9029 (N_9029,N_2623,N_417);
or U9030 (N_9030,N_9,N_4629);
xor U9031 (N_9031,N_233,N_635);
nand U9032 (N_9032,N_655,N_4816);
nor U9033 (N_9033,N_3119,N_1317);
and U9034 (N_9034,N_1618,N_2546);
and U9035 (N_9035,N_4474,N_3804);
xnor U9036 (N_9036,N_948,N_3689);
nor U9037 (N_9037,N_1946,N_745);
and U9038 (N_9038,N_3818,N_2707);
xor U9039 (N_9039,N_4286,N_3243);
xnor U9040 (N_9040,N_2729,N_4824);
xor U9041 (N_9041,N_2247,N_2895);
or U9042 (N_9042,N_2684,N_126);
and U9043 (N_9043,N_3288,N_383);
nor U9044 (N_9044,N_3231,N_4811);
nor U9045 (N_9045,N_2263,N_549);
nor U9046 (N_9046,N_2313,N_500);
and U9047 (N_9047,N_54,N_3744);
nor U9048 (N_9048,N_2843,N_49);
nand U9049 (N_9049,N_3804,N_4613);
xor U9050 (N_9050,N_4222,N_4088);
or U9051 (N_9051,N_2924,N_3755);
nor U9052 (N_9052,N_4625,N_1218);
and U9053 (N_9053,N_4459,N_1094);
or U9054 (N_9054,N_296,N_3591);
nand U9055 (N_9055,N_176,N_1515);
nor U9056 (N_9056,N_310,N_3009);
or U9057 (N_9057,N_1154,N_4362);
or U9058 (N_9058,N_3296,N_3210);
and U9059 (N_9059,N_180,N_4278);
nand U9060 (N_9060,N_1659,N_2987);
nand U9061 (N_9061,N_2499,N_3247);
nor U9062 (N_9062,N_4420,N_2061);
or U9063 (N_9063,N_2604,N_1751);
nor U9064 (N_9064,N_313,N_4741);
or U9065 (N_9065,N_1962,N_1047);
nand U9066 (N_9066,N_425,N_1088);
or U9067 (N_9067,N_1511,N_465);
nor U9068 (N_9068,N_1938,N_1149);
or U9069 (N_9069,N_4522,N_2087);
nor U9070 (N_9070,N_311,N_1312);
xnor U9071 (N_9071,N_4458,N_1314);
nor U9072 (N_9072,N_722,N_1809);
xnor U9073 (N_9073,N_3112,N_3909);
or U9074 (N_9074,N_3167,N_1634);
xnor U9075 (N_9075,N_758,N_1596);
and U9076 (N_9076,N_739,N_2728);
or U9077 (N_9077,N_180,N_1908);
nand U9078 (N_9078,N_1778,N_4784);
xnor U9079 (N_9079,N_1459,N_2827);
or U9080 (N_9080,N_4053,N_604);
nor U9081 (N_9081,N_3532,N_3682);
nor U9082 (N_9082,N_650,N_264);
nor U9083 (N_9083,N_1706,N_291);
xor U9084 (N_9084,N_3214,N_3885);
nand U9085 (N_9085,N_4573,N_2937);
xor U9086 (N_9086,N_3793,N_4992);
nor U9087 (N_9087,N_859,N_4360);
xor U9088 (N_9088,N_3136,N_4956);
xnor U9089 (N_9089,N_4706,N_4403);
and U9090 (N_9090,N_751,N_3562);
and U9091 (N_9091,N_3509,N_1102);
and U9092 (N_9092,N_1819,N_32);
nand U9093 (N_9093,N_3926,N_1323);
nor U9094 (N_9094,N_610,N_4953);
nor U9095 (N_9095,N_639,N_2678);
nand U9096 (N_9096,N_2196,N_3324);
nand U9097 (N_9097,N_1891,N_1138);
and U9098 (N_9098,N_491,N_3388);
and U9099 (N_9099,N_1025,N_1114);
nor U9100 (N_9100,N_3016,N_901);
xnor U9101 (N_9101,N_1713,N_1892);
nor U9102 (N_9102,N_3723,N_3937);
and U9103 (N_9103,N_1250,N_420);
and U9104 (N_9104,N_4386,N_4683);
xor U9105 (N_9105,N_2644,N_2487);
xnor U9106 (N_9106,N_752,N_2251);
nor U9107 (N_9107,N_4249,N_2524);
nand U9108 (N_9108,N_763,N_1328);
nor U9109 (N_9109,N_1392,N_3783);
nand U9110 (N_9110,N_1087,N_4905);
and U9111 (N_9111,N_1820,N_105);
and U9112 (N_9112,N_940,N_3352);
nor U9113 (N_9113,N_4684,N_477);
xnor U9114 (N_9114,N_141,N_838);
and U9115 (N_9115,N_4559,N_196);
or U9116 (N_9116,N_3591,N_564);
nor U9117 (N_9117,N_1769,N_2355);
xor U9118 (N_9118,N_4146,N_4613);
nor U9119 (N_9119,N_4612,N_3969);
xnor U9120 (N_9120,N_3518,N_2854);
xnor U9121 (N_9121,N_4036,N_1440);
nor U9122 (N_9122,N_2094,N_4764);
nand U9123 (N_9123,N_1521,N_663);
nand U9124 (N_9124,N_2991,N_871);
xor U9125 (N_9125,N_2183,N_2719);
nand U9126 (N_9126,N_1381,N_2640);
nand U9127 (N_9127,N_4239,N_4423);
xnor U9128 (N_9128,N_3181,N_457);
xnor U9129 (N_9129,N_4677,N_2671);
xor U9130 (N_9130,N_1382,N_969);
nor U9131 (N_9131,N_1393,N_1978);
and U9132 (N_9132,N_841,N_3274);
nand U9133 (N_9133,N_154,N_2268);
nor U9134 (N_9134,N_3209,N_711);
nor U9135 (N_9135,N_2245,N_3308);
nand U9136 (N_9136,N_3184,N_1327);
or U9137 (N_9137,N_3555,N_2298);
xnor U9138 (N_9138,N_696,N_317);
xnor U9139 (N_9139,N_1677,N_4954);
nand U9140 (N_9140,N_2903,N_3450);
or U9141 (N_9141,N_4774,N_1540);
nor U9142 (N_9142,N_4129,N_4471);
and U9143 (N_9143,N_3053,N_3207);
or U9144 (N_9144,N_3559,N_1605);
or U9145 (N_9145,N_3765,N_511);
nand U9146 (N_9146,N_142,N_3678);
nand U9147 (N_9147,N_155,N_1514);
or U9148 (N_9148,N_436,N_4251);
and U9149 (N_9149,N_2012,N_1995);
or U9150 (N_9150,N_4414,N_707);
nand U9151 (N_9151,N_3724,N_1531);
xor U9152 (N_9152,N_2582,N_2517);
nand U9153 (N_9153,N_3996,N_2094);
or U9154 (N_9154,N_1079,N_3661);
and U9155 (N_9155,N_1152,N_2950);
xor U9156 (N_9156,N_3483,N_971);
or U9157 (N_9157,N_50,N_2187);
and U9158 (N_9158,N_2910,N_3464);
xor U9159 (N_9159,N_3139,N_4490);
xor U9160 (N_9160,N_64,N_2131);
or U9161 (N_9161,N_2489,N_3750);
xnor U9162 (N_9162,N_906,N_3934);
nor U9163 (N_9163,N_2038,N_3575);
xor U9164 (N_9164,N_3129,N_1464);
and U9165 (N_9165,N_527,N_2353);
or U9166 (N_9166,N_196,N_105);
nand U9167 (N_9167,N_841,N_3095);
or U9168 (N_9168,N_4880,N_3804);
xor U9169 (N_9169,N_3022,N_642);
or U9170 (N_9170,N_3559,N_2414);
xnor U9171 (N_9171,N_2490,N_2926);
or U9172 (N_9172,N_4614,N_88);
or U9173 (N_9173,N_4935,N_4836);
xor U9174 (N_9174,N_2728,N_4942);
and U9175 (N_9175,N_1391,N_2160);
and U9176 (N_9176,N_4119,N_346);
xor U9177 (N_9177,N_457,N_971);
or U9178 (N_9178,N_2317,N_1851);
and U9179 (N_9179,N_2834,N_1345);
and U9180 (N_9180,N_387,N_1988);
nor U9181 (N_9181,N_1775,N_4552);
xnor U9182 (N_9182,N_3091,N_158);
nor U9183 (N_9183,N_2811,N_3540);
xor U9184 (N_9184,N_2316,N_461);
nor U9185 (N_9185,N_2453,N_4190);
nand U9186 (N_9186,N_4365,N_4077);
and U9187 (N_9187,N_669,N_4477);
xnor U9188 (N_9188,N_1633,N_3874);
and U9189 (N_9189,N_3840,N_4229);
nor U9190 (N_9190,N_4147,N_3473);
xnor U9191 (N_9191,N_935,N_729);
nor U9192 (N_9192,N_1561,N_1602);
xnor U9193 (N_9193,N_1599,N_3893);
nor U9194 (N_9194,N_1026,N_2441);
nor U9195 (N_9195,N_3286,N_3160);
or U9196 (N_9196,N_4802,N_1397);
xnor U9197 (N_9197,N_4240,N_3444);
nor U9198 (N_9198,N_68,N_8);
and U9199 (N_9199,N_3572,N_4448);
xnor U9200 (N_9200,N_3466,N_1036);
xnor U9201 (N_9201,N_2474,N_3794);
nor U9202 (N_9202,N_4480,N_1873);
and U9203 (N_9203,N_1330,N_4435);
and U9204 (N_9204,N_4502,N_3775);
nor U9205 (N_9205,N_4641,N_3882);
nor U9206 (N_9206,N_1904,N_376);
and U9207 (N_9207,N_1005,N_1632);
xnor U9208 (N_9208,N_4798,N_3293);
and U9209 (N_9209,N_4102,N_4928);
nor U9210 (N_9210,N_1706,N_2361);
and U9211 (N_9211,N_3381,N_4069);
and U9212 (N_9212,N_4678,N_1965);
nand U9213 (N_9213,N_2726,N_1988);
xor U9214 (N_9214,N_300,N_1157);
nand U9215 (N_9215,N_3075,N_3110);
xor U9216 (N_9216,N_4792,N_3227);
or U9217 (N_9217,N_4782,N_4212);
nor U9218 (N_9218,N_1776,N_1864);
xor U9219 (N_9219,N_1385,N_3212);
and U9220 (N_9220,N_838,N_1780);
xor U9221 (N_9221,N_1322,N_2810);
xor U9222 (N_9222,N_1800,N_2320);
xor U9223 (N_9223,N_1938,N_3372);
nand U9224 (N_9224,N_4250,N_675);
nor U9225 (N_9225,N_1795,N_1794);
nor U9226 (N_9226,N_669,N_2509);
xnor U9227 (N_9227,N_3845,N_4444);
xor U9228 (N_9228,N_306,N_1238);
xor U9229 (N_9229,N_4202,N_1450);
or U9230 (N_9230,N_121,N_2976);
and U9231 (N_9231,N_1916,N_4390);
nand U9232 (N_9232,N_718,N_2126);
nor U9233 (N_9233,N_4341,N_4854);
nor U9234 (N_9234,N_3726,N_4069);
nor U9235 (N_9235,N_3148,N_4493);
nor U9236 (N_9236,N_877,N_3069);
and U9237 (N_9237,N_1591,N_2595);
nand U9238 (N_9238,N_2136,N_4430);
nor U9239 (N_9239,N_4883,N_3515);
nand U9240 (N_9240,N_1588,N_1156);
xor U9241 (N_9241,N_3338,N_3028);
and U9242 (N_9242,N_1661,N_4908);
nor U9243 (N_9243,N_2006,N_3708);
nand U9244 (N_9244,N_890,N_1322);
nor U9245 (N_9245,N_2840,N_4261);
and U9246 (N_9246,N_1358,N_3821);
nand U9247 (N_9247,N_2175,N_763);
or U9248 (N_9248,N_3192,N_2981);
xnor U9249 (N_9249,N_3263,N_2749);
or U9250 (N_9250,N_212,N_2201);
nor U9251 (N_9251,N_4474,N_3375);
xor U9252 (N_9252,N_2657,N_2087);
xnor U9253 (N_9253,N_2794,N_19);
nor U9254 (N_9254,N_2520,N_2744);
nand U9255 (N_9255,N_3709,N_2175);
nand U9256 (N_9256,N_1858,N_9);
and U9257 (N_9257,N_3942,N_4461);
nor U9258 (N_9258,N_2206,N_511);
nor U9259 (N_9259,N_4954,N_939);
and U9260 (N_9260,N_2053,N_2869);
and U9261 (N_9261,N_1262,N_2373);
and U9262 (N_9262,N_852,N_3613);
or U9263 (N_9263,N_808,N_4761);
nor U9264 (N_9264,N_4260,N_1533);
nand U9265 (N_9265,N_4974,N_3494);
or U9266 (N_9266,N_492,N_1207);
nor U9267 (N_9267,N_1921,N_2524);
xnor U9268 (N_9268,N_822,N_2682);
and U9269 (N_9269,N_4274,N_1680);
and U9270 (N_9270,N_823,N_251);
nand U9271 (N_9271,N_518,N_2781);
nand U9272 (N_9272,N_4959,N_1262);
nand U9273 (N_9273,N_2938,N_1347);
xor U9274 (N_9274,N_4336,N_1318);
nor U9275 (N_9275,N_1283,N_4796);
xnor U9276 (N_9276,N_3984,N_1721);
and U9277 (N_9277,N_1955,N_3406);
nand U9278 (N_9278,N_4700,N_1509);
or U9279 (N_9279,N_1865,N_692);
nor U9280 (N_9280,N_1113,N_2538);
xnor U9281 (N_9281,N_4652,N_2347);
xnor U9282 (N_9282,N_3487,N_145);
or U9283 (N_9283,N_0,N_708);
xor U9284 (N_9284,N_2154,N_2323);
or U9285 (N_9285,N_161,N_2767);
nand U9286 (N_9286,N_3079,N_1022);
nor U9287 (N_9287,N_115,N_4676);
nor U9288 (N_9288,N_1278,N_4212);
or U9289 (N_9289,N_1457,N_4492);
xnor U9290 (N_9290,N_4256,N_1089);
xnor U9291 (N_9291,N_4630,N_1647);
xnor U9292 (N_9292,N_3261,N_4916);
xnor U9293 (N_9293,N_2004,N_4928);
nor U9294 (N_9294,N_3771,N_2554);
or U9295 (N_9295,N_557,N_2310);
and U9296 (N_9296,N_1520,N_4156);
nor U9297 (N_9297,N_1247,N_811);
xnor U9298 (N_9298,N_2101,N_30);
and U9299 (N_9299,N_1978,N_359);
or U9300 (N_9300,N_4007,N_1354);
or U9301 (N_9301,N_616,N_1296);
nor U9302 (N_9302,N_4856,N_1699);
nor U9303 (N_9303,N_3678,N_938);
and U9304 (N_9304,N_2015,N_4170);
nand U9305 (N_9305,N_2458,N_2246);
or U9306 (N_9306,N_1831,N_1799);
and U9307 (N_9307,N_2490,N_999);
nor U9308 (N_9308,N_514,N_1211);
and U9309 (N_9309,N_3040,N_2643);
nor U9310 (N_9310,N_4430,N_3673);
nor U9311 (N_9311,N_4837,N_4645);
or U9312 (N_9312,N_2438,N_2867);
nand U9313 (N_9313,N_113,N_4064);
xor U9314 (N_9314,N_1316,N_2743);
or U9315 (N_9315,N_4738,N_3866);
or U9316 (N_9316,N_1751,N_2736);
nand U9317 (N_9317,N_928,N_1087);
and U9318 (N_9318,N_3298,N_3980);
nand U9319 (N_9319,N_1025,N_2734);
nand U9320 (N_9320,N_3812,N_3460);
and U9321 (N_9321,N_4868,N_1153);
or U9322 (N_9322,N_2201,N_4540);
nand U9323 (N_9323,N_3073,N_1378);
nor U9324 (N_9324,N_1221,N_4407);
xor U9325 (N_9325,N_843,N_1114);
nor U9326 (N_9326,N_2328,N_3414);
nor U9327 (N_9327,N_4115,N_3797);
nand U9328 (N_9328,N_4836,N_4413);
xnor U9329 (N_9329,N_4586,N_3980);
xor U9330 (N_9330,N_1119,N_162);
nand U9331 (N_9331,N_2600,N_3525);
nand U9332 (N_9332,N_2894,N_2268);
or U9333 (N_9333,N_4954,N_1718);
nor U9334 (N_9334,N_2744,N_2498);
xor U9335 (N_9335,N_1306,N_262);
xnor U9336 (N_9336,N_257,N_1119);
nor U9337 (N_9337,N_1492,N_2490);
xnor U9338 (N_9338,N_4690,N_752);
nand U9339 (N_9339,N_1482,N_2048);
nor U9340 (N_9340,N_392,N_1556);
xnor U9341 (N_9341,N_3471,N_2712);
xnor U9342 (N_9342,N_521,N_3545);
nand U9343 (N_9343,N_1576,N_1325);
nor U9344 (N_9344,N_484,N_1850);
nor U9345 (N_9345,N_936,N_1235);
nor U9346 (N_9346,N_1520,N_2108);
xnor U9347 (N_9347,N_693,N_4251);
xor U9348 (N_9348,N_3769,N_3689);
nor U9349 (N_9349,N_1981,N_760);
nand U9350 (N_9350,N_1279,N_382);
or U9351 (N_9351,N_4810,N_1942);
nor U9352 (N_9352,N_2315,N_4064);
or U9353 (N_9353,N_2282,N_3757);
xnor U9354 (N_9354,N_190,N_3389);
and U9355 (N_9355,N_1287,N_2724);
nand U9356 (N_9356,N_2086,N_3388);
and U9357 (N_9357,N_661,N_3257);
nor U9358 (N_9358,N_2675,N_650);
and U9359 (N_9359,N_2254,N_2226);
xor U9360 (N_9360,N_483,N_2759);
or U9361 (N_9361,N_2703,N_3965);
and U9362 (N_9362,N_2333,N_545);
and U9363 (N_9363,N_1260,N_3508);
and U9364 (N_9364,N_2747,N_4338);
nand U9365 (N_9365,N_373,N_1151);
or U9366 (N_9366,N_830,N_4342);
nor U9367 (N_9367,N_2244,N_1533);
nor U9368 (N_9368,N_2529,N_3337);
nor U9369 (N_9369,N_1780,N_2444);
nor U9370 (N_9370,N_4747,N_3838);
nor U9371 (N_9371,N_2049,N_4738);
and U9372 (N_9372,N_2165,N_3971);
and U9373 (N_9373,N_2281,N_136);
xnor U9374 (N_9374,N_3685,N_4669);
nor U9375 (N_9375,N_1532,N_1970);
nand U9376 (N_9376,N_4951,N_4990);
xnor U9377 (N_9377,N_392,N_2191);
nand U9378 (N_9378,N_4292,N_1493);
or U9379 (N_9379,N_588,N_859);
xor U9380 (N_9380,N_1037,N_1528);
xor U9381 (N_9381,N_3039,N_3910);
and U9382 (N_9382,N_2830,N_4096);
or U9383 (N_9383,N_4503,N_2838);
or U9384 (N_9384,N_2323,N_4862);
or U9385 (N_9385,N_1088,N_199);
and U9386 (N_9386,N_2717,N_4013);
nand U9387 (N_9387,N_4893,N_4582);
nor U9388 (N_9388,N_2570,N_1741);
nor U9389 (N_9389,N_2598,N_3299);
or U9390 (N_9390,N_4565,N_1990);
nand U9391 (N_9391,N_4998,N_2351);
and U9392 (N_9392,N_1114,N_4475);
nand U9393 (N_9393,N_218,N_2944);
or U9394 (N_9394,N_1388,N_3512);
nor U9395 (N_9395,N_127,N_81);
or U9396 (N_9396,N_2569,N_2449);
nand U9397 (N_9397,N_3061,N_1936);
or U9398 (N_9398,N_728,N_403);
nor U9399 (N_9399,N_4336,N_3977);
or U9400 (N_9400,N_511,N_1555);
and U9401 (N_9401,N_4751,N_307);
nand U9402 (N_9402,N_1966,N_349);
or U9403 (N_9403,N_2888,N_3098);
and U9404 (N_9404,N_3235,N_3420);
nor U9405 (N_9405,N_2989,N_577);
or U9406 (N_9406,N_4778,N_4220);
or U9407 (N_9407,N_4011,N_2992);
nand U9408 (N_9408,N_1831,N_4723);
nand U9409 (N_9409,N_3900,N_2075);
xnor U9410 (N_9410,N_2905,N_1626);
xor U9411 (N_9411,N_1483,N_359);
nor U9412 (N_9412,N_1602,N_1091);
nor U9413 (N_9413,N_4232,N_2237);
nor U9414 (N_9414,N_445,N_1403);
xor U9415 (N_9415,N_1544,N_1615);
or U9416 (N_9416,N_3233,N_3609);
xnor U9417 (N_9417,N_2938,N_2139);
or U9418 (N_9418,N_2774,N_3648);
and U9419 (N_9419,N_1047,N_1076);
nand U9420 (N_9420,N_1915,N_284);
or U9421 (N_9421,N_3052,N_843);
nand U9422 (N_9422,N_3446,N_2045);
nand U9423 (N_9423,N_1914,N_1154);
and U9424 (N_9424,N_1059,N_4084);
nand U9425 (N_9425,N_1008,N_288);
xnor U9426 (N_9426,N_3488,N_1807);
and U9427 (N_9427,N_4513,N_4320);
nor U9428 (N_9428,N_3367,N_4993);
xnor U9429 (N_9429,N_4090,N_403);
nor U9430 (N_9430,N_212,N_3639);
or U9431 (N_9431,N_1559,N_1753);
or U9432 (N_9432,N_410,N_4647);
and U9433 (N_9433,N_2668,N_2340);
xnor U9434 (N_9434,N_3922,N_4797);
xnor U9435 (N_9435,N_4349,N_2212);
xor U9436 (N_9436,N_4272,N_1682);
xor U9437 (N_9437,N_2857,N_3155);
xnor U9438 (N_9438,N_2336,N_2889);
nor U9439 (N_9439,N_355,N_2213);
and U9440 (N_9440,N_1249,N_3044);
and U9441 (N_9441,N_1300,N_3121);
nand U9442 (N_9442,N_2915,N_3939);
or U9443 (N_9443,N_2140,N_837);
xor U9444 (N_9444,N_2153,N_1903);
or U9445 (N_9445,N_1273,N_2552);
xnor U9446 (N_9446,N_3551,N_231);
xor U9447 (N_9447,N_953,N_876);
or U9448 (N_9448,N_1078,N_3742);
or U9449 (N_9449,N_3038,N_35);
nand U9450 (N_9450,N_1489,N_2589);
and U9451 (N_9451,N_4722,N_3890);
and U9452 (N_9452,N_2062,N_2077);
and U9453 (N_9453,N_4013,N_1405);
nor U9454 (N_9454,N_2827,N_4310);
and U9455 (N_9455,N_956,N_2816);
and U9456 (N_9456,N_1154,N_2383);
and U9457 (N_9457,N_2074,N_22);
or U9458 (N_9458,N_2741,N_3646);
and U9459 (N_9459,N_2013,N_196);
nor U9460 (N_9460,N_726,N_1129);
nand U9461 (N_9461,N_1369,N_2313);
nor U9462 (N_9462,N_4934,N_1066);
nor U9463 (N_9463,N_2831,N_1357);
nor U9464 (N_9464,N_611,N_4543);
nor U9465 (N_9465,N_299,N_1626);
nor U9466 (N_9466,N_1621,N_1247);
nor U9467 (N_9467,N_4764,N_108);
or U9468 (N_9468,N_2165,N_969);
nor U9469 (N_9469,N_1142,N_4451);
and U9470 (N_9470,N_1109,N_338);
or U9471 (N_9471,N_3272,N_4013);
nand U9472 (N_9472,N_239,N_2744);
or U9473 (N_9473,N_1395,N_4030);
and U9474 (N_9474,N_921,N_2445);
and U9475 (N_9475,N_3149,N_246);
or U9476 (N_9476,N_3410,N_2987);
nor U9477 (N_9477,N_716,N_4540);
xor U9478 (N_9478,N_722,N_4825);
xor U9479 (N_9479,N_246,N_1904);
nor U9480 (N_9480,N_1978,N_1483);
nand U9481 (N_9481,N_2086,N_4734);
nand U9482 (N_9482,N_2021,N_467);
or U9483 (N_9483,N_1861,N_4674);
and U9484 (N_9484,N_4923,N_4151);
nand U9485 (N_9485,N_3281,N_700);
xor U9486 (N_9486,N_89,N_981);
and U9487 (N_9487,N_4667,N_3184);
or U9488 (N_9488,N_3295,N_1874);
or U9489 (N_9489,N_3320,N_4013);
or U9490 (N_9490,N_474,N_249);
and U9491 (N_9491,N_2209,N_1903);
xor U9492 (N_9492,N_1865,N_2653);
or U9493 (N_9493,N_1665,N_724);
nor U9494 (N_9494,N_2420,N_304);
nand U9495 (N_9495,N_156,N_338);
or U9496 (N_9496,N_4355,N_3776);
nor U9497 (N_9497,N_3263,N_784);
xor U9498 (N_9498,N_2484,N_554);
nand U9499 (N_9499,N_2397,N_1096);
xor U9500 (N_9500,N_2971,N_3691);
xnor U9501 (N_9501,N_4863,N_1926);
nand U9502 (N_9502,N_4276,N_1069);
nand U9503 (N_9503,N_4321,N_2216);
and U9504 (N_9504,N_4727,N_2249);
or U9505 (N_9505,N_1991,N_1158);
nor U9506 (N_9506,N_3757,N_1207);
nand U9507 (N_9507,N_4730,N_2605);
nor U9508 (N_9508,N_2095,N_3896);
nor U9509 (N_9509,N_4554,N_1596);
nand U9510 (N_9510,N_4857,N_3032);
nand U9511 (N_9511,N_722,N_4763);
nor U9512 (N_9512,N_4757,N_4836);
and U9513 (N_9513,N_2076,N_4786);
or U9514 (N_9514,N_4161,N_1149);
xor U9515 (N_9515,N_1318,N_750);
nor U9516 (N_9516,N_4318,N_1104);
and U9517 (N_9517,N_759,N_1446);
nand U9518 (N_9518,N_2190,N_4983);
xnor U9519 (N_9519,N_2352,N_2757);
nor U9520 (N_9520,N_3047,N_3549);
xnor U9521 (N_9521,N_3020,N_3719);
nor U9522 (N_9522,N_3749,N_2714);
nor U9523 (N_9523,N_3466,N_610);
xor U9524 (N_9524,N_2034,N_245);
nand U9525 (N_9525,N_1199,N_2198);
nand U9526 (N_9526,N_1061,N_4068);
xor U9527 (N_9527,N_192,N_301);
nor U9528 (N_9528,N_1557,N_611);
nand U9529 (N_9529,N_3965,N_4402);
and U9530 (N_9530,N_181,N_3409);
or U9531 (N_9531,N_640,N_1020);
and U9532 (N_9532,N_161,N_1605);
nand U9533 (N_9533,N_3129,N_4064);
xor U9534 (N_9534,N_1814,N_4924);
nand U9535 (N_9535,N_4809,N_3306);
xor U9536 (N_9536,N_1199,N_1575);
nand U9537 (N_9537,N_4505,N_3011);
or U9538 (N_9538,N_2699,N_2006);
nand U9539 (N_9539,N_733,N_4852);
nor U9540 (N_9540,N_342,N_1436);
and U9541 (N_9541,N_1828,N_2931);
nand U9542 (N_9542,N_4113,N_4467);
and U9543 (N_9543,N_3571,N_602);
nand U9544 (N_9544,N_4415,N_3557);
or U9545 (N_9545,N_4242,N_821);
xnor U9546 (N_9546,N_3971,N_4833);
or U9547 (N_9547,N_4576,N_801);
and U9548 (N_9548,N_4846,N_144);
nand U9549 (N_9549,N_2539,N_3151);
xor U9550 (N_9550,N_1796,N_4225);
or U9551 (N_9551,N_979,N_3960);
and U9552 (N_9552,N_1393,N_1572);
and U9553 (N_9553,N_4168,N_676);
nand U9554 (N_9554,N_4252,N_2426);
xor U9555 (N_9555,N_133,N_2907);
nand U9556 (N_9556,N_924,N_295);
nand U9557 (N_9557,N_2192,N_4847);
or U9558 (N_9558,N_4428,N_4778);
and U9559 (N_9559,N_2271,N_3373);
and U9560 (N_9560,N_2997,N_4554);
or U9561 (N_9561,N_108,N_4740);
or U9562 (N_9562,N_1659,N_2832);
nor U9563 (N_9563,N_4361,N_3640);
nand U9564 (N_9564,N_4947,N_3835);
nand U9565 (N_9565,N_2904,N_1299);
xor U9566 (N_9566,N_3144,N_625);
xnor U9567 (N_9567,N_3238,N_1966);
nand U9568 (N_9568,N_335,N_3633);
nand U9569 (N_9569,N_1375,N_961);
nand U9570 (N_9570,N_168,N_346);
xor U9571 (N_9571,N_3946,N_2432);
and U9572 (N_9572,N_765,N_4101);
and U9573 (N_9573,N_3814,N_1072);
nand U9574 (N_9574,N_3582,N_3222);
xor U9575 (N_9575,N_3442,N_1398);
nor U9576 (N_9576,N_1996,N_4057);
or U9577 (N_9577,N_750,N_812);
and U9578 (N_9578,N_1685,N_828);
nand U9579 (N_9579,N_4170,N_600);
nand U9580 (N_9580,N_2450,N_4315);
and U9581 (N_9581,N_3354,N_4629);
xnor U9582 (N_9582,N_2663,N_552);
or U9583 (N_9583,N_3956,N_1609);
nand U9584 (N_9584,N_1016,N_2456);
and U9585 (N_9585,N_3528,N_3694);
nand U9586 (N_9586,N_4258,N_903);
and U9587 (N_9587,N_2356,N_4974);
and U9588 (N_9588,N_3259,N_1787);
or U9589 (N_9589,N_4040,N_714);
nor U9590 (N_9590,N_2959,N_2622);
nand U9591 (N_9591,N_3055,N_3592);
and U9592 (N_9592,N_230,N_1638);
or U9593 (N_9593,N_4064,N_4503);
nor U9594 (N_9594,N_3196,N_4621);
and U9595 (N_9595,N_1438,N_2507);
or U9596 (N_9596,N_3418,N_1770);
or U9597 (N_9597,N_3806,N_4473);
xnor U9598 (N_9598,N_4995,N_2370);
nor U9599 (N_9599,N_526,N_48);
nand U9600 (N_9600,N_2997,N_3631);
nand U9601 (N_9601,N_3955,N_3875);
xnor U9602 (N_9602,N_4708,N_2566);
nor U9603 (N_9603,N_1832,N_2489);
nand U9604 (N_9604,N_90,N_2917);
or U9605 (N_9605,N_422,N_582);
xnor U9606 (N_9606,N_2395,N_642);
xor U9607 (N_9607,N_4727,N_802);
or U9608 (N_9608,N_2588,N_2042);
xnor U9609 (N_9609,N_1004,N_3939);
and U9610 (N_9610,N_3221,N_2026);
and U9611 (N_9611,N_3862,N_2012);
or U9612 (N_9612,N_2290,N_3560);
or U9613 (N_9613,N_2247,N_3668);
nand U9614 (N_9614,N_1191,N_4887);
or U9615 (N_9615,N_3907,N_1811);
nor U9616 (N_9616,N_1546,N_1291);
nand U9617 (N_9617,N_1073,N_750);
and U9618 (N_9618,N_3559,N_2782);
nor U9619 (N_9619,N_2660,N_924);
and U9620 (N_9620,N_4029,N_2973);
nand U9621 (N_9621,N_3089,N_573);
nand U9622 (N_9622,N_2189,N_1019);
xor U9623 (N_9623,N_2003,N_3795);
nor U9624 (N_9624,N_4610,N_1809);
nand U9625 (N_9625,N_1609,N_726);
or U9626 (N_9626,N_1367,N_3099);
nand U9627 (N_9627,N_3129,N_1101);
nand U9628 (N_9628,N_1195,N_1124);
xor U9629 (N_9629,N_3212,N_3049);
xor U9630 (N_9630,N_835,N_704);
nand U9631 (N_9631,N_435,N_2300);
xnor U9632 (N_9632,N_3265,N_1467);
nand U9633 (N_9633,N_1562,N_4087);
nor U9634 (N_9634,N_597,N_2503);
or U9635 (N_9635,N_3032,N_3621);
nor U9636 (N_9636,N_60,N_1237);
nand U9637 (N_9637,N_1975,N_3567);
and U9638 (N_9638,N_3335,N_3919);
xor U9639 (N_9639,N_4546,N_1604);
nor U9640 (N_9640,N_4280,N_2969);
nor U9641 (N_9641,N_1420,N_754);
nand U9642 (N_9642,N_4353,N_771);
nand U9643 (N_9643,N_4000,N_482);
xnor U9644 (N_9644,N_1786,N_1950);
nor U9645 (N_9645,N_2245,N_4062);
nor U9646 (N_9646,N_2371,N_316);
nor U9647 (N_9647,N_4071,N_2601);
nor U9648 (N_9648,N_3360,N_2198);
or U9649 (N_9649,N_1399,N_4613);
nor U9650 (N_9650,N_899,N_3641);
nor U9651 (N_9651,N_2056,N_2832);
nor U9652 (N_9652,N_1642,N_1676);
xor U9653 (N_9653,N_1756,N_185);
nor U9654 (N_9654,N_1125,N_3710);
xor U9655 (N_9655,N_1303,N_4716);
nand U9656 (N_9656,N_111,N_1351);
xor U9657 (N_9657,N_3004,N_3708);
or U9658 (N_9658,N_2656,N_1019);
nor U9659 (N_9659,N_326,N_1919);
nor U9660 (N_9660,N_1452,N_4794);
nand U9661 (N_9661,N_1439,N_4632);
and U9662 (N_9662,N_3901,N_377);
and U9663 (N_9663,N_1963,N_2491);
xor U9664 (N_9664,N_2324,N_1886);
xor U9665 (N_9665,N_2899,N_1116);
and U9666 (N_9666,N_2392,N_4911);
xnor U9667 (N_9667,N_4576,N_4231);
or U9668 (N_9668,N_644,N_2098);
or U9669 (N_9669,N_513,N_4986);
nand U9670 (N_9670,N_3638,N_1574);
xor U9671 (N_9671,N_4219,N_1787);
nor U9672 (N_9672,N_4362,N_4332);
nor U9673 (N_9673,N_1730,N_62);
and U9674 (N_9674,N_4965,N_3208);
or U9675 (N_9675,N_4790,N_574);
nor U9676 (N_9676,N_1410,N_4942);
nor U9677 (N_9677,N_3752,N_4506);
nand U9678 (N_9678,N_4412,N_1740);
and U9679 (N_9679,N_919,N_4776);
or U9680 (N_9680,N_2790,N_2345);
or U9681 (N_9681,N_3360,N_4346);
nor U9682 (N_9682,N_3275,N_83);
xor U9683 (N_9683,N_4712,N_3971);
nor U9684 (N_9684,N_4191,N_4013);
nand U9685 (N_9685,N_2353,N_1123);
and U9686 (N_9686,N_2913,N_4168);
or U9687 (N_9687,N_2299,N_233);
xor U9688 (N_9688,N_4365,N_384);
nand U9689 (N_9689,N_1401,N_3704);
and U9690 (N_9690,N_4070,N_1767);
xnor U9691 (N_9691,N_4184,N_3550);
and U9692 (N_9692,N_373,N_3441);
nand U9693 (N_9693,N_1361,N_1272);
nor U9694 (N_9694,N_3913,N_2202);
or U9695 (N_9695,N_1371,N_4917);
and U9696 (N_9696,N_1188,N_3969);
xnor U9697 (N_9697,N_3559,N_1354);
and U9698 (N_9698,N_3032,N_1792);
nor U9699 (N_9699,N_2426,N_971);
xnor U9700 (N_9700,N_969,N_3224);
xor U9701 (N_9701,N_4741,N_2981);
nor U9702 (N_9702,N_347,N_4734);
or U9703 (N_9703,N_617,N_2277);
or U9704 (N_9704,N_4169,N_1637);
nor U9705 (N_9705,N_2376,N_1646);
nor U9706 (N_9706,N_1205,N_4078);
or U9707 (N_9707,N_1777,N_1137);
nor U9708 (N_9708,N_4900,N_37);
or U9709 (N_9709,N_3435,N_1483);
xnor U9710 (N_9710,N_2574,N_396);
xor U9711 (N_9711,N_74,N_552);
xor U9712 (N_9712,N_3916,N_1213);
xor U9713 (N_9713,N_2558,N_2668);
nor U9714 (N_9714,N_4235,N_109);
and U9715 (N_9715,N_594,N_550);
xor U9716 (N_9716,N_3345,N_3309);
or U9717 (N_9717,N_1220,N_3485);
and U9718 (N_9718,N_2443,N_379);
xnor U9719 (N_9719,N_3413,N_4655);
nand U9720 (N_9720,N_3820,N_850);
nand U9721 (N_9721,N_4302,N_2237);
nand U9722 (N_9722,N_3603,N_2935);
xnor U9723 (N_9723,N_1084,N_4774);
xor U9724 (N_9724,N_69,N_505);
xor U9725 (N_9725,N_4489,N_3831);
nor U9726 (N_9726,N_1851,N_2730);
and U9727 (N_9727,N_1769,N_625);
or U9728 (N_9728,N_407,N_3168);
and U9729 (N_9729,N_2413,N_724);
or U9730 (N_9730,N_2534,N_418);
or U9731 (N_9731,N_1519,N_3762);
or U9732 (N_9732,N_202,N_2242);
or U9733 (N_9733,N_1190,N_4813);
nor U9734 (N_9734,N_3457,N_1155);
and U9735 (N_9735,N_3941,N_3433);
xor U9736 (N_9736,N_3928,N_1512);
nor U9737 (N_9737,N_1586,N_2829);
nand U9738 (N_9738,N_3573,N_1133);
or U9739 (N_9739,N_4162,N_147);
xnor U9740 (N_9740,N_2917,N_4946);
xor U9741 (N_9741,N_326,N_3481);
and U9742 (N_9742,N_19,N_1253);
nor U9743 (N_9743,N_4753,N_4934);
nor U9744 (N_9744,N_4486,N_896);
or U9745 (N_9745,N_678,N_2947);
nand U9746 (N_9746,N_747,N_437);
and U9747 (N_9747,N_712,N_3006);
nand U9748 (N_9748,N_1775,N_2803);
or U9749 (N_9749,N_3983,N_2699);
nand U9750 (N_9750,N_1016,N_2142);
nand U9751 (N_9751,N_3667,N_3547);
nor U9752 (N_9752,N_2976,N_842);
and U9753 (N_9753,N_1820,N_1922);
nor U9754 (N_9754,N_4348,N_3463);
nor U9755 (N_9755,N_2844,N_3582);
and U9756 (N_9756,N_2324,N_474);
xor U9757 (N_9757,N_1879,N_4176);
and U9758 (N_9758,N_355,N_604);
nor U9759 (N_9759,N_4415,N_1808);
xor U9760 (N_9760,N_3536,N_230);
xor U9761 (N_9761,N_4074,N_2393);
nand U9762 (N_9762,N_26,N_1199);
nor U9763 (N_9763,N_3334,N_504);
and U9764 (N_9764,N_4563,N_4630);
nand U9765 (N_9765,N_3785,N_2867);
xnor U9766 (N_9766,N_4491,N_4768);
xnor U9767 (N_9767,N_917,N_1965);
nor U9768 (N_9768,N_3780,N_841);
nand U9769 (N_9769,N_1812,N_3710);
nand U9770 (N_9770,N_1409,N_4095);
and U9771 (N_9771,N_2759,N_3520);
xor U9772 (N_9772,N_3,N_1182);
nand U9773 (N_9773,N_4703,N_2354);
or U9774 (N_9774,N_4891,N_292);
nand U9775 (N_9775,N_2786,N_1251);
xnor U9776 (N_9776,N_1892,N_1346);
xnor U9777 (N_9777,N_3409,N_4948);
and U9778 (N_9778,N_1370,N_3654);
and U9779 (N_9779,N_2475,N_532);
nor U9780 (N_9780,N_4627,N_3840);
or U9781 (N_9781,N_381,N_2423);
nand U9782 (N_9782,N_1262,N_79);
nand U9783 (N_9783,N_845,N_1831);
and U9784 (N_9784,N_3140,N_1005);
and U9785 (N_9785,N_1755,N_1679);
nand U9786 (N_9786,N_2567,N_3846);
and U9787 (N_9787,N_4627,N_439);
or U9788 (N_9788,N_4921,N_3667);
or U9789 (N_9789,N_227,N_3585);
xor U9790 (N_9790,N_3180,N_2929);
nand U9791 (N_9791,N_614,N_1856);
nor U9792 (N_9792,N_1075,N_4233);
or U9793 (N_9793,N_4424,N_3904);
nand U9794 (N_9794,N_2294,N_3131);
and U9795 (N_9795,N_2352,N_485);
nor U9796 (N_9796,N_2370,N_1155);
nor U9797 (N_9797,N_2533,N_2741);
or U9798 (N_9798,N_3209,N_1449);
nand U9799 (N_9799,N_1430,N_2661);
and U9800 (N_9800,N_925,N_3535);
or U9801 (N_9801,N_1103,N_3965);
xor U9802 (N_9802,N_1692,N_778);
xnor U9803 (N_9803,N_3304,N_2033);
nand U9804 (N_9804,N_1354,N_2611);
nor U9805 (N_9805,N_2838,N_2992);
nand U9806 (N_9806,N_2027,N_3151);
or U9807 (N_9807,N_1193,N_4175);
nor U9808 (N_9808,N_3887,N_1249);
nor U9809 (N_9809,N_1343,N_791);
nor U9810 (N_9810,N_3175,N_1230);
or U9811 (N_9811,N_3460,N_164);
and U9812 (N_9812,N_2942,N_303);
or U9813 (N_9813,N_3553,N_4295);
or U9814 (N_9814,N_2232,N_3112);
nand U9815 (N_9815,N_3125,N_4310);
or U9816 (N_9816,N_2808,N_1135);
or U9817 (N_9817,N_987,N_3776);
or U9818 (N_9818,N_3986,N_1332);
nand U9819 (N_9819,N_3133,N_4797);
nor U9820 (N_9820,N_4228,N_485);
nand U9821 (N_9821,N_2654,N_834);
or U9822 (N_9822,N_1635,N_3598);
and U9823 (N_9823,N_3916,N_3022);
or U9824 (N_9824,N_3408,N_1522);
xor U9825 (N_9825,N_516,N_3187);
or U9826 (N_9826,N_1425,N_4646);
nand U9827 (N_9827,N_637,N_4056);
nand U9828 (N_9828,N_1552,N_1310);
xnor U9829 (N_9829,N_1022,N_2531);
and U9830 (N_9830,N_3316,N_4548);
and U9831 (N_9831,N_395,N_3238);
nor U9832 (N_9832,N_4686,N_1271);
xnor U9833 (N_9833,N_3973,N_4688);
nor U9834 (N_9834,N_1013,N_160);
nor U9835 (N_9835,N_645,N_1861);
or U9836 (N_9836,N_1237,N_529);
nand U9837 (N_9837,N_2654,N_53);
and U9838 (N_9838,N_4730,N_3345);
nand U9839 (N_9839,N_3125,N_3049);
nand U9840 (N_9840,N_2850,N_3484);
and U9841 (N_9841,N_2524,N_3569);
nand U9842 (N_9842,N_2123,N_3280);
nand U9843 (N_9843,N_3511,N_752);
nor U9844 (N_9844,N_1091,N_4431);
nand U9845 (N_9845,N_362,N_2418);
or U9846 (N_9846,N_3967,N_2504);
and U9847 (N_9847,N_4908,N_3231);
nor U9848 (N_9848,N_750,N_2106);
xnor U9849 (N_9849,N_1882,N_2189);
and U9850 (N_9850,N_917,N_3564);
or U9851 (N_9851,N_3777,N_3839);
nand U9852 (N_9852,N_4081,N_3443);
xor U9853 (N_9853,N_4493,N_2588);
xnor U9854 (N_9854,N_677,N_3140);
nand U9855 (N_9855,N_2792,N_1646);
nand U9856 (N_9856,N_3178,N_2650);
nand U9857 (N_9857,N_1695,N_1838);
nand U9858 (N_9858,N_2867,N_3816);
nor U9859 (N_9859,N_360,N_2056);
nor U9860 (N_9860,N_1845,N_1876);
xor U9861 (N_9861,N_3984,N_353);
or U9862 (N_9862,N_973,N_1688);
xor U9863 (N_9863,N_2957,N_4475);
nor U9864 (N_9864,N_4062,N_4240);
or U9865 (N_9865,N_963,N_1324);
nand U9866 (N_9866,N_4443,N_2620);
or U9867 (N_9867,N_4980,N_800);
xnor U9868 (N_9868,N_4544,N_2978);
nand U9869 (N_9869,N_2321,N_2565);
nor U9870 (N_9870,N_58,N_4126);
and U9871 (N_9871,N_4298,N_4226);
and U9872 (N_9872,N_1179,N_1741);
or U9873 (N_9873,N_383,N_4586);
or U9874 (N_9874,N_3846,N_1475);
xor U9875 (N_9875,N_3826,N_3904);
xor U9876 (N_9876,N_656,N_4382);
and U9877 (N_9877,N_4850,N_1362);
nand U9878 (N_9878,N_2594,N_1662);
nor U9879 (N_9879,N_3218,N_2272);
xnor U9880 (N_9880,N_1495,N_4727);
xnor U9881 (N_9881,N_2530,N_1422);
xnor U9882 (N_9882,N_1653,N_4696);
or U9883 (N_9883,N_2886,N_3789);
and U9884 (N_9884,N_1735,N_1218);
xnor U9885 (N_9885,N_4990,N_4721);
and U9886 (N_9886,N_1968,N_3432);
and U9887 (N_9887,N_210,N_2899);
and U9888 (N_9888,N_2205,N_2736);
and U9889 (N_9889,N_3601,N_2815);
nor U9890 (N_9890,N_4095,N_2057);
and U9891 (N_9891,N_3462,N_3261);
or U9892 (N_9892,N_1425,N_3496);
and U9893 (N_9893,N_3619,N_1342);
xnor U9894 (N_9894,N_4256,N_2445);
nor U9895 (N_9895,N_4704,N_2221);
and U9896 (N_9896,N_563,N_4097);
xor U9897 (N_9897,N_3014,N_4922);
or U9898 (N_9898,N_4850,N_4242);
xor U9899 (N_9899,N_1742,N_1033);
xor U9900 (N_9900,N_2946,N_3628);
xnor U9901 (N_9901,N_4761,N_1798);
nand U9902 (N_9902,N_4828,N_4305);
and U9903 (N_9903,N_3012,N_3906);
nor U9904 (N_9904,N_4719,N_2578);
xnor U9905 (N_9905,N_1284,N_3352);
or U9906 (N_9906,N_4303,N_2195);
or U9907 (N_9907,N_4919,N_3294);
and U9908 (N_9908,N_2669,N_2515);
nand U9909 (N_9909,N_4128,N_3236);
nand U9910 (N_9910,N_3169,N_2606);
or U9911 (N_9911,N_3682,N_4826);
xor U9912 (N_9912,N_3402,N_1941);
nor U9913 (N_9913,N_4285,N_328);
xnor U9914 (N_9914,N_2699,N_2104);
nand U9915 (N_9915,N_1946,N_4719);
or U9916 (N_9916,N_1553,N_456);
nand U9917 (N_9917,N_950,N_1412);
or U9918 (N_9918,N_2558,N_1249);
and U9919 (N_9919,N_667,N_4467);
nand U9920 (N_9920,N_4454,N_2754);
nand U9921 (N_9921,N_3089,N_3588);
nor U9922 (N_9922,N_4244,N_2003);
or U9923 (N_9923,N_4650,N_870);
and U9924 (N_9924,N_40,N_2872);
nand U9925 (N_9925,N_2937,N_3839);
xor U9926 (N_9926,N_3283,N_1658);
and U9927 (N_9927,N_2754,N_4586);
nor U9928 (N_9928,N_273,N_4236);
xor U9929 (N_9929,N_199,N_51);
nand U9930 (N_9930,N_1268,N_1587);
or U9931 (N_9931,N_399,N_2760);
nand U9932 (N_9932,N_3113,N_447);
nand U9933 (N_9933,N_3475,N_1379);
or U9934 (N_9934,N_4476,N_4559);
xnor U9935 (N_9935,N_352,N_405);
and U9936 (N_9936,N_117,N_1092);
nand U9937 (N_9937,N_2413,N_4902);
xor U9938 (N_9938,N_3962,N_4093);
nand U9939 (N_9939,N_2050,N_3962);
or U9940 (N_9940,N_1205,N_4088);
nand U9941 (N_9941,N_1577,N_2407);
xnor U9942 (N_9942,N_4805,N_3065);
or U9943 (N_9943,N_2376,N_29);
nand U9944 (N_9944,N_3928,N_1790);
xnor U9945 (N_9945,N_2408,N_451);
nor U9946 (N_9946,N_4518,N_3778);
or U9947 (N_9947,N_1853,N_1280);
xnor U9948 (N_9948,N_3849,N_2848);
and U9949 (N_9949,N_250,N_704);
xor U9950 (N_9950,N_2023,N_1893);
or U9951 (N_9951,N_861,N_491);
nand U9952 (N_9952,N_689,N_3198);
xor U9953 (N_9953,N_4729,N_456);
nand U9954 (N_9954,N_3813,N_43);
xnor U9955 (N_9955,N_3066,N_902);
nand U9956 (N_9956,N_2415,N_815);
nand U9957 (N_9957,N_2493,N_4898);
xor U9958 (N_9958,N_3455,N_1181);
nand U9959 (N_9959,N_3533,N_829);
and U9960 (N_9960,N_1914,N_2038);
or U9961 (N_9961,N_1658,N_361);
nand U9962 (N_9962,N_729,N_3207);
xnor U9963 (N_9963,N_2488,N_2764);
and U9964 (N_9964,N_3674,N_427);
or U9965 (N_9965,N_1098,N_2844);
nand U9966 (N_9966,N_2334,N_129);
xnor U9967 (N_9967,N_2991,N_4017);
xor U9968 (N_9968,N_4621,N_1825);
xor U9969 (N_9969,N_1002,N_1913);
nand U9970 (N_9970,N_1587,N_3981);
nand U9971 (N_9971,N_3021,N_2527);
nand U9972 (N_9972,N_2628,N_4988);
xor U9973 (N_9973,N_349,N_4822);
or U9974 (N_9974,N_3694,N_2202);
xnor U9975 (N_9975,N_3674,N_1799);
nand U9976 (N_9976,N_2867,N_4400);
xnor U9977 (N_9977,N_3832,N_857);
nand U9978 (N_9978,N_1829,N_948);
nand U9979 (N_9979,N_1625,N_2011);
xnor U9980 (N_9980,N_2696,N_1443);
nand U9981 (N_9981,N_3621,N_3862);
and U9982 (N_9982,N_2783,N_712);
nand U9983 (N_9983,N_1145,N_927);
and U9984 (N_9984,N_2181,N_533);
nor U9985 (N_9985,N_620,N_1350);
xnor U9986 (N_9986,N_4601,N_4357);
or U9987 (N_9987,N_3604,N_884);
or U9988 (N_9988,N_4170,N_1628);
nor U9989 (N_9989,N_1395,N_2628);
nand U9990 (N_9990,N_984,N_1258);
and U9991 (N_9991,N_3168,N_4995);
and U9992 (N_9992,N_4189,N_2507);
and U9993 (N_9993,N_2894,N_4210);
and U9994 (N_9994,N_642,N_4396);
nand U9995 (N_9995,N_4944,N_3680);
or U9996 (N_9996,N_1125,N_3858);
xnor U9997 (N_9997,N_4902,N_2230);
xnor U9998 (N_9998,N_481,N_4047);
xor U9999 (N_9999,N_1915,N_4177);
and UO_0 (O_0,N_5383,N_9392);
and UO_1 (O_1,N_6653,N_7824);
nor UO_2 (O_2,N_5124,N_5300);
and UO_3 (O_3,N_6328,N_9575);
or UO_4 (O_4,N_5287,N_7508);
nand UO_5 (O_5,N_8535,N_5115);
nor UO_6 (O_6,N_7855,N_8459);
or UO_7 (O_7,N_7341,N_5946);
nand UO_8 (O_8,N_6683,N_6048);
nand UO_9 (O_9,N_9219,N_7889);
or UO_10 (O_10,N_9080,N_8261);
xor UO_11 (O_11,N_6200,N_8643);
nand UO_12 (O_12,N_6910,N_8205);
or UO_13 (O_13,N_5725,N_8406);
nand UO_14 (O_14,N_9083,N_5748);
nor UO_15 (O_15,N_6180,N_8597);
nor UO_16 (O_16,N_6838,N_7481);
nor UO_17 (O_17,N_6172,N_9253);
or UO_18 (O_18,N_8218,N_9853);
or UO_19 (O_19,N_6492,N_7790);
nor UO_20 (O_20,N_9633,N_9876);
nand UO_21 (O_21,N_6089,N_7154);
or UO_22 (O_22,N_5928,N_6562);
nor UO_23 (O_23,N_6296,N_5102);
nand UO_24 (O_24,N_8384,N_7800);
or UO_25 (O_25,N_9895,N_7608);
nand UO_26 (O_26,N_7787,N_9005);
nand UO_27 (O_27,N_8972,N_7666);
or UO_28 (O_28,N_8166,N_6763);
nand UO_29 (O_29,N_8347,N_9963);
or UO_30 (O_30,N_5910,N_7046);
nand UO_31 (O_31,N_6270,N_8054);
nand UO_32 (O_32,N_9798,N_9280);
or UO_33 (O_33,N_9590,N_5376);
xnor UO_34 (O_34,N_9707,N_7335);
or UO_35 (O_35,N_8161,N_9938);
xor UO_36 (O_36,N_8387,N_9685);
or UO_37 (O_37,N_9731,N_6050);
and UO_38 (O_38,N_7484,N_6025);
and UO_39 (O_39,N_9556,N_7865);
nor UO_40 (O_40,N_5540,N_9243);
or UO_41 (O_41,N_7580,N_5924);
and UO_42 (O_42,N_6835,N_6948);
nor UO_43 (O_43,N_8721,N_6475);
and UO_44 (O_44,N_5225,N_9235);
nor UO_45 (O_45,N_8173,N_8504);
xor UO_46 (O_46,N_9053,N_5932);
nand UO_47 (O_47,N_7297,N_8712);
and UO_48 (O_48,N_7428,N_8354);
xor UO_49 (O_49,N_6103,N_8016);
nor UO_50 (O_50,N_6801,N_5415);
nor UO_51 (O_51,N_6239,N_8555);
xor UO_52 (O_52,N_9472,N_5914);
nand UO_53 (O_53,N_7109,N_7725);
nor UO_54 (O_54,N_7300,N_6657);
nor UO_55 (O_55,N_8037,N_6153);
nand UO_56 (O_56,N_8999,N_8239);
xnor UO_57 (O_57,N_8415,N_5696);
nor UO_58 (O_58,N_7007,N_9056);
nor UO_59 (O_59,N_6952,N_5286);
xor UO_60 (O_60,N_5877,N_7543);
and UO_61 (O_61,N_7353,N_9484);
or UO_62 (O_62,N_5943,N_9749);
nor UO_63 (O_63,N_9730,N_6781);
and UO_64 (O_64,N_6419,N_6264);
and UO_65 (O_65,N_6217,N_8002);
xor UO_66 (O_66,N_5330,N_5260);
xor UO_67 (O_67,N_6031,N_7799);
and UO_68 (O_68,N_6257,N_5270);
xnor UO_69 (O_69,N_6412,N_6017);
and UO_70 (O_70,N_8063,N_6918);
xnor UO_71 (O_71,N_5476,N_5094);
xor UO_72 (O_72,N_9022,N_8596);
nor UO_73 (O_73,N_6615,N_9642);
or UO_74 (O_74,N_9382,N_9206);
nor UO_75 (O_75,N_9105,N_5487);
or UO_76 (O_76,N_6084,N_9769);
nand UO_77 (O_77,N_9334,N_8025);
or UO_78 (O_78,N_8466,N_7929);
or UO_79 (O_79,N_7697,N_6875);
and UO_80 (O_80,N_6881,N_5907);
xnor UO_81 (O_81,N_6920,N_6927);
nor UO_82 (O_82,N_5817,N_8508);
and UO_83 (O_83,N_6957,N_5159);
or UO_84 (O_84,N_6446,N_9782);
xnor UO_85 (O_85,N_8775,N_8823);
or UO_86 (O_86,N_9221,N_8518);
or UO_87 (O_87,N_7258,N_7517);
nor UO_88 (O_88,N_8579,N_7145);
nand UO_89 (O_89,N_8921,N_7304);
or UO_90 (O_90,N_6038,N_7094);
and UO_91 (O_91,N_8912,N_9130);
and UO_92 (O_92,N_8305,N_9273);
nand UO_93 (O_93,N_9409,N_9679);
xor UO_94 (O_94,N_6860,N_5746);
or UO_95 (O_95,N_5742,N_7177);
and UO_96 (O_96,N_9658,N_8815);
xor UO_97 (O_97,N_7207,N_7350);
nor UO_98 (O_98,N_8551,N_6851);
nor UO_99 (O_99,N_9848,N_7795);
or UO_100 (O_100,N_9626,N_8672);
nor UO_101 (O_101,N_8020,N_6441);
or UO_102 (O_102,N_7721,N_7354);
nor UO_103 (O_103,N_9586,N_9378);
and UO_104 (O_104,N_8625,N_8671);
nand UO_105 (O_105,N_6388,N_5846);
xor UO_106 (O_106,N_7936,N_7158);
xor UO_107 (O_107,N_8810,N_5788);
xor UO_108 (O_108,N_5876,N_5543);
nand UO_109 (O_109,N_8074,N_9996);
or UO_110 (O_110,N_6076,N_5478);
xor UO_111 (O_111,N_9281,N_7488);
xor UO_112 (O_112,N_7871,N_7456);
nand UO_113 (O_113,N_7609,N_9690);
or UO_114 (O_114,N_7429,N_8249);
xor UO_115 (O_115,N_6599,N_6995);
xor UO_116 (O_116,N_7647,N_9947);
nor UO_117 (O_117,N_6255,N_6712);
xor UO_118 (O_118,N_8482,N_6720);
nand UO_119 (O_119,N_8373,N_5289);
or UO_120 (O_120,N_9496,N_5654);
nand UO_121 (O_121,N_7486,N_5911);
nor UO_122 (O_122,N_9775,N_5798);
nand UO_123 (O_123,N_6322,N_7404);
nand UO_124 (O_124,N_8907,N_6786);
xor UO_125 (O_125,N_6049,N_9810);
nand UO_126 (O_126,N_9014,N_9192);
nand UO_127 (O_127,N_9912,N_9716);
or UO_128 (O_128,N_7271,N_8862);
or UO_129 (O_129,N_9249,N_7844);
nor UO_130 (O_130,N_5926,N_8960);
nor UO_131 (O_131,N_6061,N_5940);
or UO_132 (O_132,N_8766,N_9814);
nand UO_133 (O_133,N_6013,N_8315);
xor UO_134 (O_134,N_9141,N_9118);
xnor UO_135 (O_135,N_6895,N_7920);
or UO_136 (O_136,N_9024,N_9910);
and UO_137 (O_137,N_9131,N_8374);
nand UO_138 (O_138,N_7877,N_9041);
and UO_139 (O_139,N_6384,N_9615);
and UO_140 (O_140,N_8527,N_5023);
nand UO_141 (O_141,N_9121,N_9238);
and UO_142 (O_142,N_8969,N_8195);
or UO_143 (O_143,N_8920,N_5028);
xor UO_144 (O_144,N_5900,N_8348);
xnor UO_145 (O_145,N_6314,N_7381);
nand UO_146 (O_146,N_7050,N_7575);
and UO_147 (O_147,N_9453,N_8887);
or UO_148 (O_148,N_9874,N_8244);
and UO_149 (O_149,N_8091,N_8233);
or UO_150 (O_150,N_6627,N_6776);
xnor UO_151 (O_151,N_6744,N_8117);
xor UO_152 (O_152,N_6624,N_8515);
nand UO_153 (O_153,N_8139,N_5643);
and UO_154 (O_154,N_5887,N_5141);
nor UO_155 (O_155,N_8397,N_7657);
and UO_156 (O_156,N_5325,N_9518);
and UO_157 (O_157,N_6566,N_6277);
xnor UO_158 (O_158,N_8946,N_7991);
or UO_159 (O_159,N_5347,N_9352);
and UO_160 (O_160,N_5304,N_7351);
nor UO_161 (O_161,N_6392,N_9669);
and UO_162 (O_162,N_8719,N_8270);
and UO_163 (O_163,N_8351,N_5252);
nor UO_164 (O_164,N_5355,N_5675);
nand UO_165 (O_165,N_6090,N_8036);
nand UO_166 (O_166,N_9795,N_9369);
and UO_167 (O_167,N_9919,N_9506);
or UO_168 (O_168,N_7103,N_6959);
nand UO_169 (O_169,N_9266,N_8171);
or UO_170 (O_170,N_9728,N_9138);
nor UO_171 (O_171,N_5828,N_8359);
and UO_172 (O_172,N_5063,N_7166);
xor UO_173 (O_173,N_8404,N_8795);
nor UO_174 (O_174,N_6752,N_6261);
xnor UO_175 (O_175,N_8984,N_8248);
nor UO_176 (O_176,N_5606,N_5024);
nand UO_177 (O_177,N_9272,N_6308);
nor UO_178 (O_178,N_9201,N_6638);
and UO_179 (O_179,N_8039,N_8140);
and UO_180 (O_180,N_5973,N_7691);
nor UO_181 (O_181,N_7226,N_6142);
nor UO_182 (O_182,N_9406,N_7495);
or UO_183 (O_183,N_5871,N_6931);
and UO_184 (O_184,N_9787,N_5259);
xor UO_185 (O_185,N_8170,N_6430);
and UO_186 (O_186,N_7533,N_8104);
nor UO_187 (O_187,N_8027,N_6855);
nor UO_188 (O_188,N_7031,N_6577);
nand UO_189 (O_189,N_5802,N_9086);
nor UO_190 (O_190,N_9666,N_6782);
nand UO_191 (O_191,N_6745,N_8990);
or UO_192 (O_192,N_8340,N_9701);
nand UO_193 (O_193,N_7810,N_7966);
xnor UO_194 (O_194,N_9262,N_6067);
or UO_195 (O_195,N_6495,N_5823);
and UO_196 (O_196,N_5727,N_9144);
or UO_197 (O_197,N_7449,N_6625);
nand UO_198 (O_198,N_6483,N_6827);
nand UO_199 (O_199,N_9288,N_8350);
nand UO_200 (O_200,N_5935,N_7767);
nor UO_201 (O_201,N_6568,N_6055);
nor UO_202 (O_202,N_8476,N_8335);
nor UO_203 (O_203,N_9977,N_6333);
xnor UO_204 (O_204,N_5938,N_7834);
nand UO_205 (O_205,N_6821,N_5886);
xor UO_206 (O_206,N_8917,N_7274);
and UO_207 (O_207,N_9514,N_5966);
and UO_208 (O_208,N_9360,N_6532);
or UO_209 (O_209,N_5396,N_9002);
nand UO_210 (O_210,N_7487,N_5197);
or UO_211 (O_211,N_8809,N_5482);
xor UO_212 (O_212,N_8980,N_6734);
xnor UO_213 (O_213,N_8456,N_6858);
nor UO_214 (O_214,N_6916,N_6263);
nor UO_215 (O_215,N_7127,N_6068);
nand UO_216 (O_216,N_8971,N_5567);
and UO_217 (O_217,N_9199,N_7706);
nor UO_218 (O_218,N_5872,N_6166);
nand UO_219 (O_219,N_6907,N_7314);
nor UO_220 (O_220,N_9515,N_7163);
or UO_221 (O_221,N_9873,N_9137);
or UO_222 (O_222,N_7136,N_7831);
xor UO_223 (O_223,N_6424,N_7123);
nand UO_224 (O_224,N_8651,N_5029);
nand UO_225 (O_225,N_6613,N_7470);
and UO_226 (O_226,N_9686,N_6941);
xor UO_227 (O_227,N_7038,N_9058);
nand UO_228 (O_228,N_9610,N_8863);
nand UO_229 (O_229,N_7282,N_9309);
xnor UO_230 (O_230,N_9574,N_8026);
or UO_231 (O_231,N_9100,N_7345);
nor UO_232 (O_232,N_8873,N_9725);
nor UO_233 (O_233,N_7310,N_5048);
and UO_234 (O_234,N_8094,N_8928);
xor UO_235 (O_235,N_6199,N_6099);
xor UO_236 (O_236,N_6843,N_9720);
and UO_237 (O_237,N_5160,N_7108);
xor UO_238 (O_238,N_9306,N_8126);
and UO_239 (O_239,N_7930,N_7147);
xnor UO_240 (O_240,N_5394,N_5954);
nand UO_241 (O_241,N_9552,N_7707);
and UO_242 (O_242,N_7534,N_5890);
xor UO_243 (O_243,N_6640,N_6518);
nand UO_244 (O_244,N_7540,N_9345);
nand UO_245 (O_245,N_7067,N_7524);
or UO_246 (O_246,N_8732,N_5263);
and UO_247 (O_247,N_8461,N_6332);
or UO_248 (O_248,N_7248,N_9638);
or UO_249 (O_249,N_6220,N_9601);
or UO_250 (O_250,N_6592,N_7121);
and UO_251 (O_251,N_5255,N_5456);
or UO_252 (O_252,N_9129,N_7705);
nand UO_253 (O_253,N_6859,N_9632);
nor UO_254 (O_254,N_8297,N_6380);
nand UO_255 (O_255,N_9989,N_6487);
and UO_256 (O_256,N_5152,N_6623);
xor UO_257 (O_257,N_7757,N_7100);
nand UO_258 (O_258,N_7016,N_6012);
and UO_259 (O_259,N_9755,N_9186);
nor UO_260 (O_260,N_7285,N_9452);
or UO_261 (O_261,N_6191,N_8017);
or UO_262 (O_262,N_7909,N_5363);
and UO_263 (O_263,N_7188,N_8635);
xor UO_264 (O_264,N_8578,N_7840);
and UO_265 (O_265,N_9148,N_5208);
nand UO_266 (O_266,N_8449,N_8993);
nor UO_267 (O_267,N_9511,N_6579);
nand UO_268 (O_268,N_9381,N_8536);
nand UO_269 (O_269,N_8634,N_9331);
and UO_270 (O_270,N_5318,N_8167);
or UO_271 (O_271,N_5529,N_8163);
xor UO_272 (O_272,N_6349,N_8981);
nand UO_273 (O_273,N_6982,N_8637);
nand UO_274 (O_274,N_5971,N_9258);
xor UO_275 (O_275,N_8469,N_6452);
xnor UO_276 (O_276,N_5856,N_9940);
nand UO_277 (O_277,N_9204,N_6066);
xnor UO_278 (O_278,N_5571,N_7677);
nor UO_279 (O_279,N_9803,N_9477);
or UO_280 (O_280,N_7015,N_6706);
or UO_281 (O_281,N_5088,N_8533);
and UO_282 (O_282,N_6134,N_8839);
and UO_283 (O_283,N_6058,N_5013);
or UO_284 (O_284,N_8370,N_7489);
and UO_285 (O_285,N_8629,N_9478);
or UO_286 (O_286,N_5620,N_8944);
xnor UO_287 (O_287,N_8780,N_7415);
xnor UO_288 (O_288,N_6347,N_9962);
or UO_289 (O_289,N_7106,N_5694);
or UO_290 (O_290,N_5070,N_7416);
and UO_291 (O_291,N_8023,N_8910);
nand UO_292 (O_292,N_5261,N_8573);
and UO_293 (O_293,N_6659,N_7162);
or UO_294 (O_294,N_5575,N_9493);
xnor UO_295 (O_295,N_6963,N_5453);
nand UO_296 (O_296,N_9580,N_8070);
and UO_297 (O_297,N_8264,N_7443);
nor UO_298 (O_298,N_8072,N_7809);
and UO_299 (O_299,N_8287,N_8758);
or UO_300 (O_300,N_9924,N_6644);
and UO_301 (O_301,N_6691,N_9189);
nand UO_302 (O_302,N_5982,N_7634);
or UO_303 (O_303,N_8232,N_5142);
and UO_304 (O_304,N_7637,N_9741);
or UO_305 (O_305,N_6383,N_9342);
xnor UO_306 (O_306,N_6095,N_7664);
xor UO_307 (O_307,N_9095,N_5499);
nand UO_308 (O_308,N_9579,N_8301);
or UO_309 (O_309,N_9628,N_6197);
xnor UO_310 (O_310,N_5017,N_9625);
xnor UO_311 (O_311,N_6272,N_7122);
nor UO_312 (O_312,N_5831,N_9743);
and UO_313 (O_313,N_6366,N_5189);
and UO_314 (O_314,N_8029,N_8379);
nor UO_315 (O_315,N_6558,N_8567);
and UO_316 (O_316,N_9011,N_8836);
nand UO_317 (O_317,N_5812,N_8561);
nor UO_318 (O_318,N_7835,N_8737);
or UO_319 (O_319,N_6561,N_6081);
nor UO_320 (O_320,N_8694,N_6958);
or UO_321 (O_321,N_7217,N_8558);
and UO_322 (O_322,N_9930,N_9415);
and UO_323 (O_323,N_9285,N_6276);
xnor UO_324 (O_324,N_7990,N_9176);
or UO_325 (O_325,N_7763,N_7394);
xnor UO_326 (O_326,N_7696,N_7425);
nor UO_327 (O_327,N_6775,N_9844);
and UO_328 (O_328,N_6665,N_7048);
nand UO_329 (O_329,N_5146,N_7280);
nor UO_330 (O_330,N_8989,N_6321);
and UO_331 (O_331,N_7598,N_5918);
and UO_332 (O_332,N_9420,N_6862);
or UO_333 (O_333,N_5651,N_9291);
or UO_334 (O_334,N_5494,N_7471);
xor UO_335 (O_335,N_5648,N_9953);
or UO_336 (O_336,N_7985,N_8254);
nand UO_337 (O_337,N_9525,N_6467);
xor UO_338 (O_338,N_6671,N_6127);
xnor UO_339 (O_339,N_6517,N_6553);
and UO_340 (O_340,N_8222,N_8768);
and UO_341 (O_341,N_5011,N_9896);
or UO_342 (O_342,N_7729,N_5655);
nor UO_343 (O_343,N_7652,N_7595);
or UO_344 (O_344,N_6619,N_9356);
nor UO_345 (O_345,N_8058,N_8563);
or UO_346 (O_346,N_9832,N_5544);
or UO_347 (O_347,N_8271,N_8975);
or UO_348 (O_348,N_9967,N_5150);
nor UO_349 (O_349,N_9635,N_6667);
and UO_350 (O_350,N_8257,N_7435);
nand UO_351 (O_351,N_6030,N_6468);
xnor UO_352 (O_352,N_7700,N_5685);
nand UO_353 (O_353,N_9905,N_7545);
or UO_354 (O_354,N_8941,N_5776);
and UO_355 (O_355,N_7753,N_6954);
or UO_356 (O_356,N_5125,N_7538);
xnor UO_357 (O_357,N_6426,N_8088);
nor UO_358 (O_358,N_9470,N_8826);
nor UO_359 (O_359,N_6177,N_5615);
nand UO_360 (O_360,N_5163,N_8342);
nand UO_361 (O_361,N_7260,N_9319);
nand UO_362 (O_362,N_7252,N_6319);
xnor UO_363 (O_363,N_7837,N_7027);
xnor UO_364 (O_364,N_9046,N_8736);
nor UO_365 (O_365,N_8243,N_8229);
xnor UO_366 (O_366,N_8692,N_9605);
and UO_367 (O_367,N_8425,N_7165);
and UO_368 (O_368,N_9069,N_5006);
nor UO_369 (O_369,N_8753,N_8353);
nand UO_370 (O_370,N_9060,N_5408);
nor UO_371 (O_371,N_9950,N_8876);
and UO_372 (O_372,N_8879,N_6567);
nor UO_373 (O_373,N_7861,N_8827);
nor UO_374 (O_374,N_8467,N_5662);
xor UO_375 (O_375,N_6032,N_6373);
nor UO_376 (O_376,N_5783,N_6425);
nor UO_377 (O_377,N_6078,N_7363);
or UO_378 (O_378,N_9300,N_8548);
xnor UO_379 (O_379,N_8119,N_8645);
or UO_380 (O_380,N_9152,N_7685);
or UO_381 (O_381,N_7190,N_7602);
and UO_382 (O_382,N_8582,N_6400);
or UO_383 (O_383,N_8979,N_6991);
nand UO_384 (O_384,N_9732,N_5036);
and UO_385 (O_385,N_6148,N_7748);
or UO_386 (O_386,N_8849,N_8018);
nor UO_387 (O_387,N_7235,N_5749);
nand UO_388 (O_388,N_9321,N_6118);
xor UO_389 (O_389,N_5338,N_6139);
or UO_390 (O_390,N_7051,N_6416);
xnor UO_391 (O_391,N_6337,N_9538);
xnor UO_392 (O_392,N_8372,N_9000);
or UO_393 (O_393,N_8821,N_6541);
nand UO_394 (O_394,N_7958,N_7389);
and UO_395 (O_395,N_9191,N_7037);
and UO_396 (O_396,N_6795,N_8831);
xor UO_397 (O_397,N_6654,N_6225);
nand UO_398 (O_398,N_7793,N_8046);
nor UO_399 (O_399,N_8691,N_5485);
xor UO_400 (O_400,N_9859,N_6538);
nand UO_401 (O_401,N_7069,N_5782);
nor UO_402 (O_402,N_8794,N_7961);
nor UO_403 (O_403,N_8089,N_8857);
xnor UO_404 (O_404,N_6731,N_8465);
xor UO_405 (O_405,N_5795,N_8365);
and UO_406 (O_406,N_6814,N_9160);
nor UO_407 (O_407,N_8899,N_9978);
and UO_408 (O_408,N_5271,N_7829);
nor UO_409 (O_409,N_7539,N_9724);
and UO_410 (O_410,N_8601,N_8951);
nor UO_411 (O_411,N_8130,N_6304);
nor UO_412 (O_412,N_5730,N_7189);
xor UO_413 (O_413,N_6829,N_6486);
xnor UO_414 (O_414,N_6489,N_7380);
or UO_415 (O_415,N_8600,N_7656);
nor UO_416 (O_416,N_6988,N_5555);
or UO_417 (O_417,N_7611,N_5228);
nand UO_418 (O_418,N_7060,N_8141);
xor UO_419 (O_419,N_6074,N_8961);
nand UO_420 (O_420,N_9587,N_8165);
xor UO_421 (O_421,N_9866,N_7233);
xor UO_422 (O_422,N_9033,N_6464);
and UO_423 (O_423,N_5824,N_6621);
nor UO_424 (O_424,N_6603,N_6609);
nor UO_425 (O_425,N_5451,N_9861);
and UO_426 (O_426,N_5406,N_9405);
xnor UO_427 (O_427,N_8302,N_5869);
xnor UO_428 (O_428,N_7373,N_5254);
and UO_429 (O_429,N_5213,N_9901);
nand UO_430 (O_430,N_9278,N_8235);
and UO_431 (O_431,N_5238,N_6945);
nand UO_432 (O_432,N_7243,N_5467);
or UO_433 (O_433,N_5086,N_7014);
and UO_434 (O_434,N_6705,N_6813);
nor UO_435 (O_435,N_8355,N_9825);
nor UO_436 (O_436,N_7057,N_6122);
and UO_437 (O_437,N_9040,N_8848);
or UO_438 (O_438,N_7528,N_9098);
nor UO_439 (O_439,N_7374,N_8164);
or UO_440 (O_440,N_8904,N_5267);
and UO_441 (O_441,N_7934,N_7291);
nand UO_442 (O_442,N_5722,N_8090);
and UO_443 (O_443,N_8053,N_6800);
or UO_444 (O_444,N_7307,N_7720);
xor UO_445 (O_445,N_5805,N_7234);
nand UO_446 (O_446,N_6409,N_6062);
or UO_447 (O_447,N_5033,N_9816);
nand UO_448 (O_448,N_5671,N_6531);
and UO_449 (O_449,N_8953,N_9872);
or UO_450 (O_450,N_8591,N_7510);
nor UO_451 (O_451,N_6188,N_8564);
or UO_452 (O_452,N_9739,N_8633);
nand UO_453 (O_453,N_8933,N_5118);
nand UO_454 (O_454,N_7437,N_5777);
or UO_455 (O_455,N_8502,N_5358);
and UO_456 (O_456,N_6451,N_7526);
and UO_457 (O_457,N_9528,N_6933);
or UO_458 (O_458,N_9293,N_6759);
xor UO_459 (O_459,N_6072,N_9471);
nor UO_460 (O_460,N_6928,N_9893);
nand UO_461 (O_461,N_9554,N_9432);
xnor UO_462 (O_462,N_5888,N_9805);
and UO_463 (O_463,N_5131,N_8915);
and UO_464 (O_464,N_9490,N_9294);
nor UO_465 (O_465,N_9675,N_9088);
and UO_466 (O_466,N_5528,N_7943);
xor UO_467 (O_467,N_8819,N_5106);
nand UO_468 (O_468,N_6350,N_6890);
nor UO_469 (O_469,N_8291,N_7605);
nor UO_470 (O_470,N_6980,N_6309);
xor UO_471 (O_471,N_7496,N_5965);
xor UO_472 (O_472,N_6051,N_5458);
nand UO_473 (O_473,N_9208,N_8686);
and UO_474 (O_474,N_8890,N_7887);
nor UO_475 (O_475,N_9326,N_7971);
and UO_476 (O_476,N_9788,N_7976);
nand UO_477 (O_477,N_5019,N_7750);
nor UO_478 (O_478,N_7995,N_8763);
xnor UO_479 (O_479,N_6007,N_5616);
nand UO_480 (O_480,N_8032,N_9400);
and UO_481 (O_481,N_7424,N_6241);
xnor UO_482 (O_482,N_8797,N_5369);
or UO_483 (O_483,N_9316,N_5042);
and UO_484 (O_484,N_7775,N_7529);
and UO_485 (O_485,N_9617,N_9376);
nand UO_486 (O_486,N_9299,N_6693);
xor UO_487 (O_487,N_6879,N_8991);
and UO_488 (O_488,N_9951,N_7823);
or UO_489 (O_489,N_6470,N_5686);
nor UO_490 (O_490,N_5078,N_7279);
or UO_491 (O_491,N_9619,N_5021);
nand UO_492 (O_492,N_8224,N_9548);
xor UO_493 (O_493,N_6923,N_9702);
nand UO_494 (O_494,N_7076,N_5153);
nand UO_495 (O_495,N_6196,N_8662);
nand UO_496 (O_496,N_6970,N_9327);
nor UO_497 (O_497,N_5372,N_6227);
nand UO_498 (O_498,N_6125,N_5865);
or UO_499 (O_499,N_5765,N_8722);
nor UO_500 (O_500,N_7982,N_5420);
xor UO_501 (O_501,N_7808,N_8396);
and UO_502 (O_502,N_9116,N_6646);
and UO_503 (O_503,N_7925,N_6990);
and UO_504 (O_504,N_9494,N_9412);
xor UO_505 (O_505,N_9536,N_8192);
nor UO_506 (O_506,N_7328,N_9877);
and UO_507 (O_507,N_6240,N_6819);
or UO_508 (O_508,N_8419,N_8022);
and UO_509 (O_509,N_9786,N_9437);
xor UO_510 (O_510,N_9240,N_5829);
and UO_511 (O_511,N_8896,N_6676);
and UO_512 (O_512,N_7391,N_9667);
and UO_513 (O_513,N_8252,N_5491);
nand UO_514 (O_514,N_6584,N_8893);
nand UO_515 (O_515,N_5060,N_9178);
nand UO_516 (O_516,N_7139,N_6629);
and UO_517 (O_517,N_6323,N_7713);
nor UO_518 (O_518,N_9665,N_9001);
xor UO_519 (O_519,N_7588,N_7392);
nor UO_520 (O_520,N_9142,N_7161);
and UO_521 (O_521,N_7789,N_7056);
and UO_522 (O_522,N_6466,N_5979);
and UO_523 (O_523,N_7138,N_7267);
and UO_524 (O_524,N_5364,N_5666);
or UO_525 (O_525,N_9467,N_5596);
or UO_526 (O_526,N_6407,N_7500);
nand UO_527 (O_527,N_6938,N_8512);
or UO_528 (O_528,N_8604,N_7878);
nor UO_529 (O_529,N_6649,N_9197);
nand UO_530 (O_530,N_6773,N_5915);
or UO_531 (O_531,N_8854,N_9195);
nor UO_532 (O_532,N_8735,N_9236);
nor UO_533 (O_533,N_7583,N_5995);
and UO_534 (O_534,N_8044,N_7679);
nor UO_535 (O_535,N_5322,N_5859);
nand UO_536 (O_536,N_5706,N_5903);
and UO_537 (O_537,N_8174,N_8781);
or UO_538 (O_538,N_6060,N_8695);
nor UO_539 (O_539,N_6126,N_6340);
nor UO_540 (O_540,N_7535,N_5658);
xor UO_541 (O_541,N_5145,N_6986);
nor UO_542 (O_542,N_8380,N_9964);
xor UO_543 (O_543,N_9245,N_9268);
and UO_544 (O_544,N_9337,N_7079);
and UO_545 (O_545,N_7115,N_7370);
xnor UO_546 (O_546,N_9408,N_8534);
xor UO_547 (O_547,N_6867,N_5941);
xnor UO_548 (O_548,N_7357,N_8615);
xor UO_549 (O_549,N_8138,N_5379);
xor UO_550 (O_550,N_9710,N_9547);
nand UO_551 (O_551,N_6436,N_6202);
or UO_552 (O_552,N_9827,N_9427);
xnor UO_553 (O_553,N_9431,N_9802);
and UO_554 (O_554,N_6248,N_5366);
xnor UO_555 (O_555,N_9763,N_7506);
nand UO_556 (O_556,N_7276,N_8358);
nand UO_557 (O_557,N_7615,N_8496);
xor UO_558 (O_558,N_9062,N_7197);
nor UO_559 (O_559,N_6936,N_7883);
nand UO_560 (O_560,N_5969,N_6144);
nor UO_561 (O_561,N_7743,N_9362);
nand UO_562 (O_562,N_6794,N_8111);
nand UO_563 (O_563,N_6785,N_5361);
or UO_564 (O_564,N_7585,N_6826);
and UO_565 (O_565,N_7680,N_7515);
nand UO_566 (O_566,N_9850,N_9015);
or UO_567 (O_567,N_6024,N_9247);
nor UO_568 (O_568,N_8443,N_9530);
or UO_569 (O_569,N_8450,N_7176);
nand UO_570 (O_570,N_7549,N_9124);
or UO_571 (O_571,N_8842,N_9516);
nor UO_572 (O_572,N_6902,N_7548);
or UO_573 (O_573,N_6901,N_9045);
nor UO_574 (O_574,N_8143,N_9597);
nand UO_575 (O_575,N_8718,N_5122);
nor UO_576 (O_576,N_8930,N_5623);
and UO_577 (O_577,N_7850,N_9147);
xnor UO_578 (O_578,N_9009,N_6668);
nand UO_579 (O_579,N_8332,N_9609);
xnor UO_580 (O_580,N_6290,N_5414);
xnor UO_581 (O_581,N_6765,N_9837);
and UO_582 (O_582,N_7408,N_9394);
or UO_583 (O_583,N_6360,N_6585);
nand UO_584 (O_584,N_6563,N_8491);
nand UO_585 (O_585,N_7420,N_8471);
nor UO_586 (O_586,N_8986,N_8409);
xnor UO_587 (O_587,N_5594,N_9153);
nand UO_588 (O_588,N_6680,N_7811);
and UO_589 (O_589,N_8505,N_9187);
and UO_590 (O_590,N_8782,N_6506);
nor UO_591 (O_591,N_5084,N_6056);
nand UO_592 (O_592,N_9593,N_8363);
and UO_593 (O_593,N_6565,N_6445);
nor UO_594 (O_594,N_6684,N_8872);
or UO_595 (O_595,N_7036,N_6278);
and UO_596 (O_596,N_5904,N_5690);
and UO_597 (O_597,N_9375,N_5100);
nand UO_598 (O_598,N_9101,N_7324);
nand UO_599 (O_599,N_5522,N_9090);
or UO_600 (O_600,N_6317,N_6658);
and UO_601 (O_601,N_8460,N_8773);
nand UO_602 (O_602,N_9821,N_9372);
nor UO_603 (O_603,N_8865,N_8431);
and UO_604 (O_604,N_6774,N_8874);
nor UO_605 (O_605,N_9689,N_9073);
and UO_606 (O_606,N_6273,N_9289);
xor UO_607 (O_607,N_5558,N_8376);
nand UO_608 (O_608,N_7536,N_7501);
and UO_609 (O_609,N_6942,N_6458);
nor UO_610 (O_610,N_7815,N_8446);
and UO_611 (O_611,N_6992,N_5315);
xor UO_612 (O_612,N_7625,N_8339);
and UO_613 (O_613,N_9296,N_8092);
xnor UO_614 (O_614,N_7011,N_5077);
nand UO_615 (O_615,N_8177,N_7229);
or UO_616 (O_616,N_5986,N_7941);
and UO_617 (O_617,N_5492,N_8660);
xor UO_618 (O_618,N_7021,N_7562);
and UO_619 (O_619,N_9984,N_9995);
and UO_620 (O_620,N_9966,N_6973);
or UO_621 (O_621,N_6453,N_7343);
nor UO_622 (O_622,N_5840,N_6414);
and UO_623 (O_623,N_9361,N_8976);
xor UO_624 (O_624,N_7546,N_9719);
and UO_625 (O_625,N_9329,N_5939);
nor UO_626 (O_626,N_8537,N_6488);
nor UO_627 (O_627,N_9834,N_6431);
nand UO_628 (O_628,N_5500,N_9807);
nor UO_629 (O_629,N_9421,N_5292);
and UO_630 (O_630,N_7827,N_8648);
and UO_631 (O_631,N_5429,N_6463);
xor UO_632 (O_632,N_8647,N_8522);
nand UO_633 (O_633,N_5661,N_5665);
and UO_634 (O_634,N_8010,N_6303);
and UO_635 (O_635,N_5839,N_6546);
nand UO_636 (O_636,N_9343,N_6913);
xnor UO_637 (O_637,N_7622,N_9469);
nor UO_638 (O_638,N_8843,N_7892);
xnor UO_639 (O_639,N_5851,N_6145);
and UO_640 (O_640,N_6543,N_6187);
xor UO_641 (O_641,N_5386,N_6642);
nand UO_642 (O_642,N_6305,N_6357);
nand UO_643 (O_643,N_6828,N_5072);
and UO_644 (O_644,N_7296,N_9527);
nor UO_645 (O_645,N_9799,N_9026);
nand UO_646 (O_646,N_6703,N_7204);
xnor UO_647 (O_647,N_9505,N_5919);
and UO_648 (O_648,N_6138,N_9384);
and UO_649 (O_649,N_6355,N_5297);
nor UO_650 (O_650,N_8544,N_7938);
nor UO_651 (O_651,N_7120,N_5912);
and UO_652 (O_652,N_6494,N_5906);
nand UO_653 (O_653,N_8470,N_8656);
xnor UO_654 (O_654,N_8030,N_5760);
nor UO_655 (O_655,N_6209,N_6628);
or UO_656 (O_656,N_6904,N_6677);
nand UO_657 (O_657,N_5639,N_8116);
nand UO_658 (O_658,N_5819,N_5521);
nand UO_659 (O_659,N_7186,N_7075);
and UO_660 (O_660,N_8383,N_9900);
or UO_661 (O_661,N_6442,N_7777);
or UO_662 (O_662,N_6964,N_9125);
nor UO_663 (O_663,N_7203,N_5027);
xor UO_664 (O_664,N_5232,N_5274);
or UO_665 (O_665,N_8549,N_7346);
or UO_666 (O_666,N_9314,N_5387);
nor UO_667 (O_667,N_5020,N_7978);
nand UO_668 (O_668,N_7187,N_8269);
nor UO_669 (O_669,N_8784,N_5466);
xor UO_670 (O_670,N_5180,N_9284);
nand UO_671 (O_671,N_8859,N_5642);
nor UO_672 (O_672,N_8760,N_7205);
nor UO_673 (O_673,N_9433,N_9926);
and UO_674 (O_674,N_7749,N_7091);
nor UO_675 (O_675,N_9793,N_5293);
nor UO_676 (O_676,N_6233,N_9123);
nand UO_677 (O_677,N_7505,N_6271);
and UO_678 (O_678,N_5673,N_5380);
or UO_679 (O_679,N_9760,N_8041);
and UO_680 (O_680,N_7755,N_8151);
nand UO_681 (O_681,N_5385,N_9332);
nand UO_682 (O_682,N_8182,N_9465);
nor UO_683 (O_683,N_6528,N_6015);
or UO_684 (O_684,N_8125,N_8565);
xnor UO_685 (O_685,N_8097,N_6783);
nand UO_686 (O_686,N_6950,N_6358);
nand UO_687 (O_687,N_9885,N_6674);
xnor UO_688 (O_688,N_9081,N_5656);
xnor UO_689 (O_689,N_6435,N_8272);
and UO_690 (O_690,N_5923,N_6112);
and UO_691 (O_691,N_7269,N_7485);
xor UO_692 (O_692,N_7928,N_8369);
xor UO_693 (O_693,N_5687,N_5857);
xnor UO_694 (O_694,N_5498,N_9082);
or UO_695 (O_695,N_7308,N_8318);
and UO_696 (O_696,N_5603,N_8429);
and UO_697 (O_697,N_5844,N_6632);
or UO_698 (O_698,N_7741,N_6096);
xnor UO_699 (O_699,N_6014,N_8381);
xnor UO_700 (O_700,N_6354,N_8853);
nand UO_701 (O_701,N_6313,N_8328);
or UO_702 (O_702,N_6169,N_9766);
nand UO_703 (O_703,N_7237,N_5958);
or UO_704 (O_704,N_6912,N_9255);
nor UO_705 (O_705,N_5509,N_9581);
nand UO_706 (O_706,N_7955,N_8199);
xor UO_707 (O_707,N_9570,N_6178);
nor UO_708 (O_708,N_6190,N_9648);
nand UO_709 (O_709,N_7239,N_6154);
and UO_710 (O_710,N_6438,N_9945);
and UO_711 (O_711,N_8223,N_6527);
nor UO_712 (O_712,N_8987,N_5963);
nand UO_713 (O_713,N_8813,N_9904);
or UO_714 (O_714,N_5542,N_7125);
nor UO_715 (O_715,N_9154,N_7295);
and UO_716 (O_716,N_6755,N_8108);
or UO_717 (O_717,N_7368,N_7316);
xnor UO_718 (O_718,N_6878,N_8581);
nand UO_719 (O_719,N_9179,N_8569);
or UO_720 (O_720,N_8674,N_5893);
nand UO_721 (O_721,N_7012,N_7689);
nor UO_722 (O_722,N_6523,N_7760);
nand UO_723 (O_723,N_7098,N_8666);
or UO_724 (O_724,N_8411,N_8957);
or UO_725 (O_725,N_8623,N_7250);
nand UO_726 (O_726,N_6105,N_7025);
and UO_727 (O_727,N_6189,N_9757);
xnor UO_728 (O_728,N_6165,N_5400);
xor UO_729 (O_729,N_8416,N_9998);
nand UO_730 (O_730,N_5479,N_5207);
nor UO_731 (O_731,N_6777,N_6281);
xnor UO_732 (O_732,N_7309,N_5244);
nand UO_733 (O_733,N_9474,N_9210);
and UO_734 (O_734,N_7445,N_9429);
and UO_735 (O_735,N_7593,N_8178);
xnor UO_736 (O_736,N_5113,N_8599);
or UO_737 (O_737,N_6097,N_6764);
nand UO_738 (O_738,N_5809,N_8321);
nor UO_739 (O_739,N_7004,N_6883);
xor UO_740 (O_740,N_5157,N_6806);
nor UO_741 (O_741,N_7899,N_8285);
xnor UO_742 (O_742,N_8064,N_6131);
xnor UO_743 (O_743,N_5878,N_5920);
nor UO_744 (O_744,N_6919,N_5524);
xnor UO_745 (O_745,N_6413,N_9908);
or UO_746 (O_746,N_6588,N_9907);
nand UO_747 (O_747,N_6472,N_5961);
and UO_748 (O_748,N_6971,N_5663);
nor UO_749 (O_749,N_9407,N_8407);
or UO_750 (O_750,N_6293,N_7774);
nor UO_751 (O_751,N_9091,N_6885);
or UO_752 (O_752,N_6591,N_9035);
and UO_753 (O_753,N_9884,N_7433);
xor UO_754 (O_754,N_8377,N_9705);
nand UO_755 (O_755,N_6481,N_7044);
or UO_756 (O_756,N_6020,N_6326);
nor UO_757 (O_757,N_6622,N_8447);
and UO_758 (O_758,N_9535,N_8811);
xnor UO_759 (O_759,N_5638,N_7240);
nor UO_760 (O_760,N_5459,N_5032);
or UO_761 (O_761,N_8298,N_9959);
nand UO_762 (O_762,N_7013,N_7169);
nor UO_763 (O_763,N_6737,N_5179);
nor UO_764 (O_764,N_5576,N_8209);
nor UO_765 (O_765,N_8659,N_7151);
xor UO_766 (O_766,N_5947,N_5336);
nand UO_767 (O_767,N_8220,N_9796);
nand UO_768 (O_768,N_8822,N_5195);
nand UO_769 (O_769,N_7465,N_8451);
nand UO_770 (O_770,N_7918,N_8142);
and UO_771 (O_771,N_7731,N_8307);
nand UO_772 (O_772,N_9899,N_5371);
nor UO_773 (O_773,N_6456,N_9991);
or UO_774 (O_774,N_9468,N_6685);
nand UO_775 (O_775,N_7080,N_8366);
or UO_776 (O_776,N_9445,N_8640);
or UO_777 (O_777,N_9287,N_9096);
and UO_778 (O_778,N_7020,N_7178);
or UO_779 (O_779,N_8242,N_9983);
and UO_780 (O_780,N_8898,N_7215);
nand UO_781 (O_781,N_9230,N_8770);
nor UO_782 (O_782,N_5121,N_8619);
and UO_783 (O_783,N_6484,N_9423);
and UO_784 (O_784,N_7028,N_9158);
and UO_785 (O_785,N_7356,N_5635);
nor UO_786 (O_786,N_7492,N_9340);
and UO_787 (O_787,N_9676,N_5584);
nand UO_788 (O_788,N_6849,N_9368);
xnor UO_789 (O_789,N_9704,N_9157);
and UO_790 (O_790,N_6497,N_8817);
nand UO_791 (O_791,N_9170,N_8576);
or UO_792 (O_792,N_7254,N_8186);
nor UO_793 (O_793,N_9244,N_9887);
nor UO_794 (O_794,N_8776,N_6534);
and UO_795 (O_795,N_7135,N_5800);
and UO_796 (O_796,N_8851,N_9055);
or UO_797 (O_797,N_7002,N_7641);
xnor UO_798 (O_798,N_5810,N_8480);
or UO_799 (O_799,N_6042,N_8901);
nor UO_800 (O_800,N_5018,N_7643);
nand UO_801 (O_801,N_6824,N_9031);
and UO_802 (O_802,N_9233,N_7676);
or UO_803 (O_803,N_7218,N_8925);
and UO_804 (O_804,N_5341,N_8762);
xor UO_805 (O_805,N_5841,N_9561);
nand UO_806 (O_806,N_5423,N_6286);
or UO_807 (O_807,N_8791,N_7618);
nor UO_808 (O_808,N_6837,N_9583);
nor UO_809 (O_809,N_8115,N_9475);
nand UO_810 (O_810,N_7502,N_8630);
and UO_811 (O_811,N_8121,N_7804);
xor UO_812 (O_812,N_5047,N_8977);
nand UO_813 (O_813,N_8861,N_6465);
nor UO_814 (O_814,N_5419,N_8803);
or UO_815 (O_815,N_5041,N_7005);
or UO_816 (O_816,N_5595,N_7576);
and UO_817 (O_817,N_9146,N_5230);
or UO_818 (O_818,N_9085,N_8334);
nor UO_819 (O_819,N_9512,N_7419);
nand UO_820 (O_820,N_8316,N_8913);
xnor UO_821 (O_821,N_5570,N_9566);
and UO_822 (O_822,N_7994,N_5123);
or UO_823 (O_823,N_6274,N_8047);
or UO_824 (O_824,N_8942,N_7390);
xor UO_825 (O_825,N_9792,N_8278);
xnor UO_826 (O_826,N_6510,N_5010);
nor UO_827 (O_827,N_8789,N_6678);
nand UO_828 (O_828,N_7491,N_6767);
and UO_829 (O_829,N_8183,N_6002);
xor UO_830 (O_830,N_7323,N_6093);
or UO_831 (O_831,N_5452,N_8344);
or UO_832 (O_832,N_8389,N_9502);
or UO_833 (O_833,N_8325,N_6194);
nand UO_834 (O_834,N_8948,N_8294);
nand UO_835 (O_835,N_9008,N_5715);
and UO_836 (O_836,N_7146,N_5791);
xnor UO_837 (O_837,N_6892,N_7710);
nor UO_838 (O_838,N_6738,N_6932);
nand UO_839 (O_839,N_7065,N_8102);
and UO_840 (O_840,N_5870,N_6069);
nand UO_841 (O_841,N_7574,N_6573);
xor UO_842 (O_842,N_9975,N_9770);
and UO_843 (O_843,N_7772,N_7360);
nand UO_844 (O_844,N_7838,N_6833);
or UO_845 (O_845,N_6841,N_7460);
nand UO_846 (O_846,N_7040,N_5064);
and UO_847 (O_847,N_6161,N_7423);
or UO_848 (O_848,N_5416,N_5203);
nand UO_849 (O_849,N_6922,N_5176);
nor UO_850 (O_850,N_8994,N_7265);
nand UO_851 (O_851,N_6836,N_9181);
xnor UO_852 (O_852,N_9135,N_7009);
nand UO_853 (O_853,N_8992,N_9499);
nand UO_854 (O_854,N_9365,N_5204);
nand UO_855 (O_855,N_5889,N_7338);
or UO_856 (O_856,N_5849,N_7305);
and UO_857 (O_857,N_5470,N_5786);
or UO_858 (O_858,N_9611,N_7654);
or UO_859 (O_859,N_8727,N_9023);
or UO_860 (O_860,N_7072,N_6756);
or UO_861 (O_861,N_8498,N_7780);
xor UO_862 (O_862,N_6823,N_6717);
or UO_863 (O_863,N_9169,N_6533);
xnor UO_864 (O_864,N_7054,N_7355);
nand UO_865 (O_865,N_7184,N_5196);
nor UO_866 (O_866,N_8949,N_8752);
xnor UO_867 (O_867,N_8066,N_8492);
nand UO_868 (O_868,N_7975,N_8414);
nand UO_869 (O_869,N_8556,N_6618);
nor UO_870 (O_870,N_6474,N_7452);
xor UO_871 (O_871,N_7915,N_7728);
nor UO_872 (O_872,N_6586,N_7552);
nor UO_873 (O_873,N_7140,N_8681);
nand UO_874 (O_874,N_7172,N_8568);
nand UO_875 (O_875,N_6761,N_7256);
and UO_876 (O_876,N_6063,N_7983);
xor UO_877 (O_877,N_7418,N_8965);
nor UO_878 (O_878,N_8168,N_8250);
nand UO_879 (O_879,N_9596,N_5014);
nor UO_880 (O_880,N_7225,N_8448);
xnor UO_881 (O_881,N_8005,N_5688);
nor UO_882 (O_882,N_9852,N_8324);
xor UO_883 (O_883,N_7723,N_6500);
nand UO_884 (O_884,N_8059,N_6559);
xor UO_885 (O_885,N_5449,N_5758);
and UO_886 (O_886,N_5375,N_5793);
xnor UO_887 (O_887,N_7348,N_6847);
nand UO_888 (O_888,N_7693,N_7523);
nand UO_889 (O_889,N_6955,N_9892);
xor UO_890 (O_890,N_9205,N_9673);
nand UO_891 (O_891,N_5922,N_9303);
nor UO_892 (O_892,N_6036,N_8276);
nor UO_893 (O_893,N_9781,N_5188);
nor UO_894 (O_894,N_7347,N_7459);
xnor UO_895 (O_895,N_6411,N_7367);
nor UO_896 (O_896,N_8333,N_9745);
xor UO_897 (O_897,N_5587,N_7066);
nor UO_898 (O_898,N_5333,N_6427);
nor UO_899 (O_899,N_6236,N_9275);
and UO_900 (O_900,N_9497,N_7766);
or UO_901 (O_901,N_5578,N_7074);
nand UO_902 (O_902,N_5737,N_8685);
xor UO_903 (O_903,N_7261,N_8043);
nand UO_904 (O_904,N_5426,N_9217);
nor UO_905 (O_905,N_5564,N_8306);
nor UO_906 (O_906,N_7655,N_5311);
and UO_907 (O_907,N_5512,N_8517);
and UO_908 (O_908,N_9140,N_5373);
xnor UO_909 (O_909,N_6865,N_7765);
or UO_910 (O_910,N_5069,N_8131);
and UO_911 (O_911,N_6218,N_9212);
xnor UO_912 (O_912,N_5883,N_8349);
and UO_913 (O_913,N_9006,N_5327);
nand UO_914 (O_914,N_7601,N_7263);
xnor UO_915 (O_915,N_5306,N_7722);
xor UO_916 (O_916,N_8189,N_8922);
and UO_917 (O_917,N_6011,N_7128);
or UO_918 (O_918,N_9168,N_7438);
nand UO_919 (O_919,N_8057,N_6643);
nor UO_920 (O_920,N_8546,N_9111);
xor UO_921 (O_921,N_9336,N_7541);
or UO_922 (O_922,N_7849,N_9777);
xor UO_923 (O_923,N_5148,N_7033);
and UO_924 (O_924,N_7483,N_6551);
nor UO_925 (O_925,N_7716,N_5993);
nand UO_926 (O_926,N_7940,N_6079);
nor UO_927 (O_927,N_9371,N_7686);
nor UO_928 (O_928,N_9092,N_5181);
or UO_929 (O_929,N_5510,N_6539);
nor UO_930 (O_930,N_5736,N_8884);
or UO_931 (O_931,N_9177,N_5505);
nor UO_932 (O_932,N_9209,N_8663);
xor UO_933 (O_933,N_6348,N_6318);
or UO_934 (O_934,N_8201,N_7587);
and UO_935 (O_935,N_9416,N_5956);
nand UO_936 (O_936,N_7195,N_8012);
nand UO_937 (O_937,N_7668,N_8764);
nand UO_938 (O_938,N_6804,N_8742);
or UO_939 (O_939,N_7732,N_5465);
and UO_940 (O_940,N_8850,N_9434);
and UO_941 (O_941,N_8045,N_6336);
and UO_942 (O_942,N_6193,N_9762);
nand UO_943 (O_943,N_7714,N_9183);
nor UO_944 (O_944,N_6370,N_8750);
nor UO_945 (O_945,N_6873,N_8497);
nand UO_946 (O_946,N_6460,N_9753);
xor UO_947 (O_947,N_9678,N_6812);
nor UO_948 (O_948,N_7385,N_6171);
and UO_949 (O_949,N_7862,N_6108);
nand UO_950 (O_950,N_9824,N_5626);
and UO_951 (O_951,N_7783,N_9634);
xnor UO_952 (O_952,N_6136,N_9537);
or UO_953 (O_953,N_9703,N_5360);
nand UO_954 (O_954,N_8364,N_5562);
and UO_955 (O_955,N_8771,N_5137);
nor UO_956 (O_956,N_8627,N_5609);
and UO_957 (O_957,N_9915,N_8641);
xnor UO_958 (O_958,N_8609,N_9569);
and UO_959 (O_959,N_9629,N_9027);
and UO_960 (O_960,N_8122,N_8124);
or UO_961 (O_961,N_6147,N_6092);
and UO_962 (O_962,N_8690,N_7671);
nand UO_963 (O_963,N_6772,N_6476);
nor UO_964 (O_964,N_6159,N_8711);
xor UO_965 (O_965,N_6167,N_9565);
xor UO_966 (O_966,N_7673,N_7984);
nor UO_967 (O_967,N_5182,N_7785);
nand UO_968 (O_968,N_5796,N_8606);
and UO_969 (O_969,N_6265,N_8019);
nor UO_970 (O_970,N_6876,N_5699);
nand UO_971 (O_971,N_5237,N_6351);
or UO_972 (O_972,N_7378,N_9606);
xor UO_973 (O_973,N_7908,N_6793);
or UO_974 (O_974,N_5134,N_9656);
nor UO_975 (O_975,N_5934,N_6226);
nand UO_976 (O_976,N_7532,N_5640);
nor UO_977 (O_977,N_9539,N_6201);
or UO_978 (O_978,N_9681,N_8009);
nor UO_979 (O_979,N_5071,N_7053);
nor UO_980 (O_980,N_5607,N_5161);
nand UO_981 (O_981,N_8513,N_8593);
xnor UO_982 (O_982,N_7320,N_7858);
and UO_983 (O_983,N_5110,N_8799);
and UO_984 (O_984,N_7628,N_6001);
and UO_985 (O_985,N_7665,N_6447);
nor UO_986 (O_986,N_8083,N_5475);
or UO_987 (O_987,N_7997,N_5343);
or UO_988 (O_988,N_5837,N_8346);
xnor UO_989 (O_989,N_6617,N_9458);
xnor UO_990 (O_990,N_9122,N_6287);
xor UO_991 (O_991,N_5972,N_6330);
and UO_992 (O_992,N_7633,N_7474);
and UO_993 (O_993,N_9584,N_9234);
and UO_994 (O_994,N_5395,N_5632);
nor UO_995 (O_995,N_7432,N_6082);
nand UO_996 (O_996,N_7064,N_6604);
and UO_997 (O_997,N_9145,N_6537);
nor UO_998 (O_998,N_8268,N_8612);
and UO_999 (O_999,N_6284,N_9349);
nor UO_1000 (O_1000,N_9668,N_6754);
nand UO_1001 (O_1001,N_9222,N_5533);
and UO_1002 (O_1002,N_5461,N_7068);
nand UO_1003 (O_1003,N_9748,N_5210);
xor UO_1004 (O_1004,N_8203,N_5556);
nand UO_1005 (O_1005,N_8883,N_5814);
nand UO_1006 (O_1006,N_7825,N_8824);
nand UO_1007 (O_1007,N_7259,N_5245);
nand UO_1008 (O_1008,N_5762,N_9460);
xor UO_1009 (O_1009,N_8237,N_5701);
or UO_1010 (O_1010,N_7859,N_9733);
xor UO_1011 (O_1011,N_5480,N_5281);
nand UO_1012 (O_1012,N_6418,N_9010);
xor UO_1013 (O_1013,N_8368,N_8231);
xnor UO_1014 (O_1014,N_9845,N_7442);
or UO_1015 (O_1015,N_5774,N_7856);
nor UO_1016 (O_1016,N_7084,N_6041);
and UO_1017 (O_1017,N_9974,N_6769);
xor UO_1018 (O_1018,N_8962,N_7898);
xnor UO_1019 (O_1019,N_6949,N_7644);
or UO_1020 (O_1020,N_9598,N_9698);
and UO_1021 (O_1021,N_8006,N_5726);
or UO_1022 (O_1022,N_6505,N_7318);
and UO_1023 (O_1023,N_8705,N_9374);
nand UO_1024 (O_1024,N_9050,N_6450);
nor UO_1025 (O_1025,N_9216,N_8828);
nor UO_1026 (O_1026,N_5104,N_6119);
or UO_1027 (O_1027,N_7864,N_6729);
nor UO_1028 (O_1028,N_8145,N_6224);
nand UO_1029 (O_1029,N_7382,N_6548);
or UO_1030 (O_1030,N_6046,N_9932);
nor UO_1031 (O_1031,N_5342,N_7950);
nor UO_1032 (O_1032,N_6880,N_7393);
and UO_1033 (O_1033,N_6212,N_9075);
nor UO_1034 (O_1034,N_9047,N_7022);
xnor UO_1035 (O_1035,N_6730,N_5202);
nor UO_1036 (O_1036,N_8382,N_7779);
nor UO_1037 (O_1037,N_7302,N_7126);
nor UO_1038 (O_1038,N_5874,N_7876);
nor UO_1039 (O_1039,N_9671,N_5664);
and UO_1040 (O_1040,N_6675,N_6779);
xnor UO_1041 (O_1041,N_8300,N_7979);
or UO_1042 (O_1042,N_8392,N_6387);
nand UO_1043 (O_1043,N_9627,N_7704);
nand UO_1044 (O_1044,N_5155,N_6057);
xnor UO_1045 (O_1045,N_9970,N_9127);
nor UO_1046 (O_1046,N_9099,N_9851);
nand UO_1047 (O_1047,N_9456,N_6267);
xnor UO_1048 (O_1048,N_5206,N_5566);
or UO_1049 (O_1049,N_7262,N_7264);
nor UO_1050 (O_1050,N_6019,N_5092);
and UO_1051 (O_1051,N_8547,N_6960);
nand UO_1052 (O_1052,N_8557,N_7600);
and UO_1053 (O_1053,N_8914,N_8806);
and UO_1054 (O_1054,N_9902,N_9647);
nor UO_1055 (O_1055,N_5240,N_6893);
or UO_1056 (O_1056,N_6389,N_5848);
xnor UO_1057 (O_1057,N_7361,N_6698);
or UO_1058 (O_1058,N_7843,N_9533);
or UO_1059 (O_1059,N_5862,N_5641);
and UO_1060 (O_1060,N_7284,N_5720);
nand UO_1061 (O_1061,N_9811,N_6173);
xnor UO_1062 (O_1062,N_8749,N_5425);
and UO_1063 (O_1063,N_6367,N_6975);
nand UO_1064 (O_1064,N_5707,N_5215);
and UO_1065 (O_1065,N_6029,N_5231);
or UO_1066 (O_1066,N_9736,N_7414);
or UO_1067 (O_1067,N_7451,N_9226);
nor UO_1068 (O_1068,N_9004,N_5393);
nand UO_1069 (O_1069,N_9398,N_5354);
xnor UO_1070 (O_1070,N_8918,N_5272);
or UO_1071 (O_1071,N_6040,N_5243);
or UO_1072 (O_1072,N_7377,N_9504);
or UO_1073 (O_1073,N_9640,N_8729);
and UO_1074 (O_1074,N_8160,N_9495);
nand UO_1075 (O_1075,N_8048,N_6612);
or UO_1076 (O_1076,N_8440,N_7095);
nand UO_1077 (O_1077,N_6116,N_7339);
nor UO_1078 (O_1078,N_8463,N_8653);
and UO_1079 (O_1079,N_7559,N_5346);
or UO_1080 (O_1080,N_6143,N_9359);
xnor UO_1081 (O_1081,N_9879,N_7819);
and UO_1082 (O_1082,N_9113,N_9304);
or UO_1083 (O_1083,N_5834,N_8273);
and UO_1084 (O_1084,N_7399,N_5477);
xnor UO_1085 (O_1085,N_9858,N_9322);
nand UO_1086 (O_1086,N_7088,N_5660);
and UO_1087 (O_1087,N_8716,N_6291);
xor UO_1088 (O_1088,N_8128,N_7872);
nor UO_1089 (O_1089,N_5807,N_8553);
xor UO_1090 (O_1090,N_5066,N_8683);
nand UO_1091 (O_1091,N_8858,N_6520);
xnor UO_1092 (O_1092,N_8710,N_9986);
xnor UO_1093 (O_1093,N_5627,N_8731);
and UO_1094 (O_1094,N_5296,N_7581);
nand UO_1095 (O_1095,N_7337,N_9200);
nor UO_1096 (O_1096,N_9190,N_9607);
xnor UO_1097 (O_1097,N_8702,N_5119);
xnor UO_1098 (O_1098,N_8162,N_9891);
and UO_1099 (O_1099,N_9225,N_5835);
xor UO_1100 (O_1100,N_9500,N_6521);
nor UO_1101 (O_1101,N_8255,N_6983);
and UO_1102 (O_1102,N_6170,N_8200);
or UO_1103 (O_1103,N_6182,N_5326);
nor UO_1104 (O_1104,N_9328,N_9357);
xor UO_1105 (O_1105,N_8055,N_5605);
or UO_1106 (O_1106,N_7077,N_7556);
and UO_1107 (O_1107,N_8357,N_9729);
nor UO_1108 (O_1108,N_7822,N_7427);
xor UO_1109 (O_1109,N_6149,N_7761);
or UO_1110 (O_1110,N_6672,N_9363);
nand UO_1111 (O_1111,N_8947,N_7651);
nand UO_1112 (O_1112,N_5317,N_5483);
xor UO_1113 (O_1113,N_5044,N_5813);
and UO_1114 (O_1114,N_6669,N_9061);
and UO_1115 (O_1115,N_7071,N_8696);
and UO_1116 (O_1116,N_5140,N_5209);
nor UO_1117 (O_1117,N_5710,N_6150);
nor UO_1118 (O_1118,N_6331,N_9425);
and UO_1119 (O_1119,N_7518,N_6498);
nand UO_1120 (O_1120,N_5403,N_5672);
nand UO_1121 (O_1121,N_8526,N_5917);
nor UO_1122 (O_1122,N_9623,N_9740);
and UO_1123 (O_1123,N_8759,N_8970);
nor UO_1124 (O_1124,N_8792,N_5775);
nor UO_1125 (O_1125,N_8830,N_8472);
or UO_1126 (O_1126,N_9509,N_5549);
xor UO_1127 (O_1127,N_5407,N_8275);
xnor UO_1128 (O_1128,N_6750,N_5678);
and UO_1129 (O_1129,N_9052,N_7913);
xor UO_1130 (O_1130,N_6564,N_7582);
nor UO_1131 (O_1131,N_8462,N_8926);
or UO_1132 (O_1132,N_6701,N_6587);
xnor UO_1133 (O_1133,N_6047,N_9411);
nor UO_1134 (O_1134,N_5413,N_9889);
and UO_1135 (O_1135,N_6035,N_5205);
or UO_1136 (O_1136,N_8499,N_8588);
and UO_1137 (O_1137,N_5953,N_6993);
nor UO_1138 (O_1138,N_7813,N_8421);
nand UO_1139 (O_1139,N_9038,N_9708);
nor UO_1140 (O_1140,N_6803,N_5321);
nand UO_1141 (O_1141,N_9659,N_8326);
nor UO_1142 (O_1142,N_6021,N_9695);
nand UO_1143 (O_1143,N_5096,N_6059);
xor UO_1144 (O_1144,N_7584,N_9418);
nor UO_1145 (O_1145,N_9660,N_9301);
and UO_1146 (O_1146,N_8998,N_7327);
xor UO_1147 (O_1147,N_5691,N_7507);
nor UO_1148 (O_1148,N_5553,N_7124);
xor UO_1149 (O_1149,N_6788,N_7244);
nand UO_1150 (O_1150,N_8113,N_7242);
xor UO_1151 (O_1151,N_9688,N_8153);
and UO_1152 (O_1152,N_7214,N_6850);
nor UO_1153 (O_1153,N_7703,N_7439);
nand UO_1154 (O_1154,N_8511,N_7578);
nand UO_1155 (O_1155,N_6616,N_7059);
and UO_1156 (O_1156,N_7631,N_5511);
nor UO_1157 (O_1157,N_6485,N_6000);
xor UO_1158 (O_1158,N_8441,N_6098);
nor UO_1159 (O_1159,N_5370,N_5535);
or UO_1160 (O_1160,N_5674,N_7062);
nand UO_1161 (O_1161,N_7567,N_6114);
xnor UO_1162 (O_1162,N_5863,N_9602);
and UO_1163 (O_1163,N_5186,N_9917);
and UO_1164 (O_1164,N_7616,N_7089);
nand UO_1165 (O_1165,N_8251,N_7087);
and UO_1166 (O_1166,N_6449,N_6863);
xnor UO_1167 (O_1167,N_9573,N_7592);
nor UO_1168 (O_1168,N_7156,N_6866);
and UO_1169 (O_1169,N_9928,N_9849);
nand UO_1170 (O_1170,N_9488,N_8093);
xnor UO_1171 (O_1171,N_9198,N_9311);
xnor UO_1172 (O_1172,N_9150,N_9347);
and UO_1173 (O_1173,N_5200,N_5832);
nand UO_1174 (O_1174,N_9612,N_7773);
or UO_1175 (O_1175,N_5242,N_6661);
nand UO_1176 (O_1176,N_8428,N_5046);
nand UO_1177 (O_1177,N_7897,N_8973);
or UO_1178 (O_1178,N_9639,N_6915);
or UO_1179 (O_1179,N_5569,N_6018);
nand UO_1180 (O_1180,N_5950,N_6371);
xnor UO_1181 (O_1181,N_7213,N_7682);
or UO_1182 (O_1182,N_5985,N_7255);
nand UO_1183 (O_1183,N_7194,N_5352);
nor UO_1184 (O_1184,N_7134,N_9613);
xnor UO_1185 (O_1185,N_5411,N_7695);
nand UO_1186 (O_1186,N_8631,N_9990);
xnor UO_1187 (O_1187,N_6306,N_6719);
nand UO_1188 (O_1188,N_9591,N_6977);
nand UO_1189 (O_1189,N_9106,N_9202);
or UO_1190 (O_1190,N_5994,N_6502);
xor UO_1191 (O_1191,N_6816,N_9631);
xnor UO_1192 (O_1192,N_8709,N_8479);
nand UO_1193 (O_1193,N_5942,N_7379);
or UO_1194 (O_1194,N_6213,N_6423);
nor UO_1195 (O_1195,N_9750,N_5531);
or UO_1196 (O_1196,N_8510,N_9641);
nand UO_1197 (O_1197,N_8919,N_6569);
and UO_1198 (O_1198,N_6937,N_6999);
nand UO_1199 (O_1199,N_7446,N_6647);
nand UO_1200 (O_1200,N_6796,N_9758);
or UO_1201 (O_1201,N_9399,N_9937);
and UO_1202 (O_1202,N_8283,N_6530);
xor UO_1203 (O_1203,N_8408,N_6243);
or UO_1204 (O_1204,N_5450,N_8777);
or UO_1205 (O_1205,N_7604,N_8889);
nor UO_1206 (O_1206,N_8060,N_5220);
xnor UO_1207 (O_1207,N_9034,N_9697);
xor UO_1208 (O_1208,N_6989,N_8995);
xor UO_1209 (O_1209,N_5258,N_9655);
nand UO_1210 (O_1210,N_5009,N_8495);
nor UO_1211 (O_1211,N_9325,N_8983);
nand UO_1212 (O_1212,N_5581,N_9355);
xor UO_1213 (O_1213,N_8337,N_9097);
xnor UO_1214 (O_1214,N_8613,N_5412);
or UO_1215 (O_1215,N_6168,N_9388);
nor UO_1216 (O_1216,N_8678,N_8187);
nor UO_1217 (O_1217,N_7894,N_9167);
nand UO_1218 (O_1218,N_9454,N_6259);
xor UO_1219 (O_1219,N_5990,N_5653);
nor UO_1220 (O_1220,N_5645,N_9976);
and UO_1221 (O_1221,N_7768,N_8520);
and UO_1222 (O_1222,N_9549,N_9324);
nand UO_1223 (O_1223,N_7922,N_5432);
nand UO_1224 (O_1224,N_7035,N_8708);
xnor UO_1225 (O_1225,N_9507,N_5057);
nor UO_1226 (O_1226,N_7649,N_6655);
xnor UO_1227 (O_1227,N_8587,N_6924);
and UO_1228 (O_1228,N_7290,N_5294);
or UO_1229 (O_1229,N_5693,N_8477);
and UO_1230 (O_1230,N_6298,N_8410);
nand UO_1231 (O_1231,N_8436,N_8210);
nor UO_1232 (O_1232,N_7164,N_6686);
xor UO_1233 (O_1233,N_7826,N_7464);
or UO_1234 (O_1234,N_9229,N_5767);
xnor UO_1235 (O_1235,N_7674,N_6815);
nand UO_1236 (O_1236,N_8552,N_7150);
nand UO_1237 (O_1237,N_5392,N_8723);
nor UO_1238 (O_1238,N_8049,N_8490);
nand UO_1239 (O_1239,N_8675,N_8042);
nand UO_1240 (O_1240,N_5136,N_8234);
nor UO_1241 (O_1241,N_9608,N_6401);
nor UO_1242 (O_1242,N_7667,N_6842);
nand UO_1243 (O_1243,N_8101,N_5264);
or UO_1244 (O_1244,N_7561,N_6529);
nand UO_1245 (O_1245,N_9483,N_5502);
or UO_1246 (O_1246,N_8402,N_6909);
or UO_1247 (O_1247,N_8266,N_8265);
or UO_1248 (O_1248,N_5448,N_5167);
or UO_1249 (O_1249,N_5288,N_8611);
nand UO_1250 (O_1250,N_5440,N_9077);
nor UO_1251 (O_1251,N_7413,N_5808);
xnor UO_1252 (O_1252,N_5646,N_5740);
and UO_1253 (O_1253,N_7398,N_6799);
xor UO_1254 (O_1254,N_7981,N_7210);
nand UO_1255 (O_1255,N_5496,N_5446);
and UO_1256 (O_1256,N_9264,N_8751);
nor UO_1257 (O_1257,N_6723,N_7266);
xnor UO_1258 (O_1258,N_8745,N_8855);
xnor UO_1259 (O_1259,N_5580,N_6802);
nand UO_1260 (O_1260,N_7833,N_6162);
or UO_1261 (O_1261,N_5780,N_5175);
or UO_1262 (O_1262,N_5211,N_5614);
and UO_1263 (O_1263,N_5039,N_5820);
xnor UO_1264 (O_1264,N_8481,N_6889);
and UO_1265 (O_1265,N_7684,N_9519);
nor UO_1266 (O_1266,N_9016,N_8007);
nor UO_1267 (O_1267,N_6361,N_7694);
or UO_1268 (O_1268,N_8118,N_5224);
nor UO_1269 (O_1269,N_7426,N_8693);
nor UO_1270 (O_1270,N_6714,N_8227);
nor UO_1271 (O_1271,N_9076,N_8069);
and UO_1272 (O_1272,N_7560,N_6378);
and UO_1273 (O_1273,N_8021,N_5348);
or UO_1274 (O_1274,N_6593,N_7692);
nor UO_1275 (O_1275,N_9276,N_6976);
nor UO_1276 (O_1276,N_5040,N_6262);
or UO_1277 (O_1277,N_9931,N_5026);
xor UO_1278 (O_1278,N_6770,N_5015);
and UO_1279 (O_1279,N_8607,N_7143);
or UO_1280 (O_1280,N_7854,N_7101);
xnor UO_1281 (O_1281,N_9290,N_6727);
nor UO_1282 (O_1282,N_9335,N_7881);
xnor UO_1283 (O_1283,N_9295,N_6176);
or UO_1284 (O_1284,N_5866,N_8592);
nor UO_1285 (O_1285,N_8159,N_5967);
nor UO_1286 (O_1286,N_9459,N_8881);
nor UO_1287 (O_1287,N_6130,N_7907);
xor UO_1288 (O_1288,N_5171,N_6094);
nand UO_1289 (O_1289,N_5778,N_8602);
nor UO_1290 (O_1290,N_5053,N_5381);
xnor UO_1291 (O_1291,N_9109,N_7191);
nor UO_1292 (O_1292,N_8963,N_8500);
nand UO_1293 (O_1293,N_9112,N_7784);
nor UO_1294 (O_1294,N_7457,N_8703);
nand UO_1295 (O_1295,N_6258,N_9481);
and UO_1296 (O_1296,N_8541,N_7231);
and UO_1297 (O_1297,N_8620,N_8514);
and UO_1298 (O_1298,N_9529,N_9155);
nor UO_1299 (O_1299,N_8923,N_5668);
and UO_1300 (O_1300,N_6549,N_6778);
and UO_1301 (O_1301,N_5250,N_6984);
xnor UO_1302 (O_1302,N_6222,N_6575);
and UO_1303 (O_1303,N_8288,N_6376);
nor UO_1304 (O_1304,N_5650,N_7998);
or UO_1305 (O_1305,N_5838,N_6757);
xnor UO_1306 (O_1306,N_8575,N_6395);
xnor UO_1307 (O_1307,N_8524,N_7959);
nor UO_1308 (O_1308,N_6299,N_8096);
nor UO_1309 (O_1309,N_8099,N_5649);
nand UO_1310 (O_1310,N_8430,N_6461);
nand UO_1311 (O_1311,N_7717,N_6065);
nand UO_1312 (O_1312,N_6728,N_5061);
or UO_1313 (O_1313,N_7181,N_7951);
and UO_1314 (O_1314,N_5409,N_6997);
nor UO_1315 (O_1315,N_7802,N_9320);
or UO_1316 (O_1316,N_8725,N_7882);
xor UO_1317 (O_1317,N_7935,N_9119);
nor UO_1318 (O_1318,N_5998,N_6557);
nor UO_1319 (O_1319,N_8157,N_5977);
nor UO_1320 (O_1320,N_8062,N_7275);
and UO_1321 (O_1321,N_7117,N_7762);
and UO_1322 (O_1322,N_5850,N_9084);
xor UO_1323 (O_1323,N_7709,N_5323);
or UO_1324 (O_1324,N_8621,N_7431);
or UO_1325 (O_1325,N_5144,N_5750);
nor UO_1326 (O_1326,N_6028,N_5068);
or UO_1327 (O_1327,N_7230,N_9032);
nor UO_1328 (O_1328,N_7253,N_8309);
or UO_1329 (O_1329,N_9890,N_9649);
or UO_1330 (O_1330,N_5582,N_9674);
nand UO_1331 (O_1331,N_8832,N_7494);
nor UO_1332 (O_1332,N_6353,N_5797);
xnor UO_1333 (O_1333,N_6739,N_6064);
or UO_1334 (O_1334,N_9385,N_6379);
and UO_1335 (O_1335,N_9078,N_9231);
nand UO_1336 (O_1336,N_5621,N_6252);
and UO_1337 (O_1337,N_7669,N_7454);
nand UO_1338 (O_1338,N_5227,N_6219);
and UO_1339 (O_1339,N_9828,N_7544);
and UO_1340 (O_1340,N_7550,N_8106);
or UO_1341 (O_1341,N_5534,N_7663);
nor UO_1342 (O_1342,N_9117,N_5779);
and UO_1343 (O_1343,N_5248,N_5708);
and UO_1344 (O_1344,N_5825,N_7006);
xnor UO_1345 (O_1345,N_8454,N_9797);
and UO_1346 (O_1346,N_6972,N_5065);
and UO_1347 (O_1347,N_7639,N_8540);
nor UO_1348 (O_1348,N_8198,N_5852);
and UO_1349 (O_1349,N_5390,N_9094);
nor UO_1350 (O_1350,N_6343,N_6688);
or UO_1351 (O_1351,N_9867,N_7568);
nor UO_1352 (O_1352,N_9927,N_9207);
xor UO_1353 (O_1353,N_9971,N_9110);
nor UO_1354 (O_1354,N_8743,N_9903);
and UO_1355 (O_1355,N_9833,N_5629);
xnor UO_1356 (O_1356,N_8968,N_5855);
and UO_1357 (O_1357,N_7209,N_8532);
nand UO_1358 (O_1358,N_9270,N_7839);
nand UO_1359 (O_1359,N_6552,N_6320);
or UO_1360 (O_1360,N_5804,N_8082);
nor UO_1361 (O_1361,N_6285,N_5111);
nand UO_1362 (O_1362,N_9897,N_5310);
or UO_1363 (O_1363,N_7565,N_8911);
or UO_1364 (O_1364,N_5340,N_6480);
xnor UO_1365 (O_1365,N_6874,N_9341);
and UO_1366 (O_1366,N_8078,N_7278);
and UO_1367 (O_1367,N_6792,N_7530);
nor UO_1368 (O_1368,N_5151,N_5612);
xnor UO_1369 (O_1369,N_8714,N_5218);
nor UO_1370 (O_1370,N_6344,N_7814);
or UO_1371 (O_1371,N_5992,N_6550);
or UO_1372 (O_1372,N_8658,N_6341);
nor UO_1373 (O_1373,N_7281,N_7514);
xnor UO_1374 (O_1374,N_6133,N_6386);
nand UO_1375 (O_1375,N_7270,N_7821);
and UO_1376 (O_1376,N_5335,N_8147);
nor UO_1377 (O_1377,N_8452,N_5283);
or UO_1378 (O_1378,N_9274,N_5217);
xor UO_1379 (O_1379,N_5617,N_5826);
nand UO_1380 (O_1380,N_8152,N_7436);
xnor UO_1381 (O_1381,N_9692,N_6639);
nand UO_1382 (O_1382,N_6985,N_7642);
nor UO_1383 (O_1383,N_6522,N_8804);
nand UO_1384 (O_1384,N_5368,N_9269);
nor UO_1385 (O_1385,N_6968,N_9922);
or UO_1386 (O_1386,N_9396,N_8772);
and UO_1387 (O_1387,N_9439,N_6185);
xor UO_1388 (O_1388,N_9841,N_6715);
or UO_1389 (O_1389,N_7756,N_9577);
or UO_1390 (O_1390,N_9560,N_8172);
and UO_1391 (O_1391,N_5249,N_9523);
or UO_1392 (O_1392,N_8473,N_8475);
or UO_1393 (O_1393,N_5388,N_5921);
nor UO_1394 (O_1394,N_7232,N_9817);
xor UO_1395 (O_1395,N_5875,N_8765);
nor UO_1396 (O_1396,N_8726,N_5328);
and UO_1397 (O_1397,N_8281,N_7475);
nor UO_1398 (O_1398,N_8852,N_6288);
or UO_1399 (O_1399,N_7952,N_8673);
nand UO_1400 (O_1400,N_9451,N_9875);
nand UO_1401 (O_1401,N_7715,N_7055);
nor UO_1402 (O_1402,N_7358,N_6831);
nand UO_1403 (O_1403,N_7180,N_8903);
nand UO_1404 (O_1404,N_9012,N_7073);
nor UO_1405 (O_1405,N_8085,N_8225);
and UO_1406 (O_1406,N_5105,N_8566);
and UO_1407 (O_1407,N_7142,N_7104);
and UO_1408 (O_1408,N_7171,N_5759);
nor UO_1409 (O_1409,N_9260,N_6369);
nor UO_1410 (O_1410,N_5464,N_6888);
xor UO_1411 (O_1411,N_5389,N_8538);
nor UO_1412 (O_1412,N_8013,N_7236);
nand UO_1413 (O_1413,N_8181,N_8412);
nor UO_1414 (O_1414,N_5625,N_8323);
and UO_1415 (O_1415,N_5214,N_8156);
nand UO_1416 (O_1416,N_6073,N_6512);
nor UO_1417 (O_1417,N_6961,N_8507);
and UO_1418 (O_1418,N_7573,N_6109);
and UO_1419 (O_1419,N_8489,N_8240);
xor UO_1420 (O_1420,N_5541,N_6610);
xor UO_1421 (O_1421,N_5295,N_9920);
xnor UO_1422 (O_1422,N_6808,N_7557);
and UO_1423 (O_1423,N_8877,N_9436);
nand UO_1424 (O_1424,N_6987,N_5002);
and UO_1425 (O_1425,N_7890,N_9042);
nor UO_1426 (O_1426,N_9184,N_6282);
or UO_1427 (O_1427,N_7086,N_8570);
nand UO_1428 (O_1428,N_7321,N_6429);
and UO_1429 (O_1429,N_7434,N_5784);
nor UO_1430 (O_1430,N_9888,N_7462);
xor UO_1431 (O_1431,N_6375,N_9949);
or UO_1432 (O_1432,N_6682,N_6307);
nand UO_1433 (O_1433,N_8788,N_5703);
and UO_1434 (O_1434,N_7551,N_8338);
and UO_1435 (O_1435,N_5572,N_8149);
or UO_1436 (O_1436,N_5892,N_6006);
nand UO_1437 (O_1437,N_8632,N_8668);
nor UO_1438 (O_1438,N_7078,N_8864);
and UO_1439 (O_1439,N_7919,N_5622);
xor UO_1440 (O_1440,N_5827,N_9691);
nor UO_1441 (O_1441,N_9174,N_5593);
xnor UO_1442 (O_1442,N_5754,N_5091);
nand UO_1443 (O_1443,N_5976,N_9636);
xnor UO_1444 (O_1444,N_5443,N_6229);
nor UO_1445 (O_1445,N_6052,N_8964);
nor UO_1446 (O_1446,N_5980,N_8783);
xnor UO_1447 (O_1447,N_7241,N_8583);
nand UO_1448 (O_1448,N_9139,N_5978);
or UO_1449 (O_1449,N_5035,N_7085);
xnor UO_1450 (O_1450,N_9585,N_8395);
nand UO_1451 (O_1451,N_7817,N_6141);
nor UO_1452 (O_1452,N_5418,N_7553);
nor UO_1453 (O_1453,N_7148,N_9994);
or UO_1454 (O_1454,N_5516,N_6335);
or UO_1455 (O_1455,N_9578,N_9466);
or UO_1456 (O_1456,N_7102,N_5517);
and UO_1457 (O_1457,N_7946,N_9312);
nand UO_1458 (O_1458,N_7157,N_6325);
or UO_1459 (O_1459,N_8038,N_5854);
or UO_1460 (O_1460,N_6235,N_6540);
xor UO_1461 (O_1461,N_8313,N_7322);
nor UO_1462 (O_1462,N_5016,N_8988);
xnor UO_1463 (O_1463,N_7554,N_5551);
nand UO_1464 (O_1464,N_8644,N_5899);
or UO_1465 (O_1465,N_6477,N_6524);
nor UO_1466 (O_1466,N_9868,N_9043);
nor UO_1467 (O_1467,N_7497,N_7764);
and UO_1468 (O_1468,N_7000,N_5716);
nand UO_1469 (O_1469,N_6820,N_8399);
or UO_1470 (O_1470,N_8929,N_9256);
and UO_1471 (O_1471,N_7083,N_7917);
xnor UO_1472 (O_1472,N_8779,N_7853);
and UO_1473 (O_1473,N_5495,N_5331);
and UO_1474 (O_1474,N_9108,N_9404);
and UO_1475 (O_1475,N_7400,N_7092);
nand UO_1476 (O_1476,N_7885,N_9323);
xor UO_1477 (O_1477,N_5052,N_5677);
or UO_1478 (O_1478,N_7520,N_5695);
and UO_1479 (O_1479,N_7944,N_8746);
nor UO_1480 (O_1480,N_7504,N_9603);
nand UO_1481 (O_1481,N_8503,N_9227);
or UO_1482 (O_1482,N_5669,N_7522);
or UO_1483 (O_1483,N_7746,N_5437);
nand UO_1484 (O_1484,N_9070,N_9934);
nor UO_1485 (O_1485,N_5178,N_5473);
nor UO_1486 (O_1486,N_7277,N_8068);
or UO_1487 (O_1487,N_7168,N_7223);
xnor UO_1488 (O_1488,N_6751,N_5506);
and UO_1489 (O_1489,N_5265,N_5515);
nor UO_1490 (O_1490,N_6311,N_6010);
and UO_1491 (O_1491,N_5391,N_6210);
nand UO_1492 (O_1492,N_8571,N_6117);
and UO_1493 (O_1493,N_6886,N_9487);
nand UO_1494 (O_1494,N_7963,N_9401);
xor UO_1495 (O_1495,N_8439,N_7558);
and UO_1496 (O_1496,N_9840,N_5868);
nand UO_1497 (O_1497,N_6023,N_6711);
nor UO_1498 (O_1498,N_5357,N_5733);
and UO_1499 (O_1499,N_7132,N_5345);
endmodule